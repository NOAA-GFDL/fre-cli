netcdf \20030101.atmos_static_cmip.tile3 {
dimensions:
	grid_xt = 96 ;
	grid_yt = 96 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:associated_files = "area: 20030101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 time = 0 ;

 orog =
  1.957085, 182.3516, 345.853, 566.5532, 583.9197, 703.0031, 841.8619, 
    930.701, 1327.418, 1866.999, 2029.211, 1998.469, 1606.435, 2058.914, 
    894.809, 267.2261, 1038.635, 95.99315, -29, -29, -14.74468, 50.54665, 
    131.9456, 149.8255, 180.3951, 144.0376, 117.0449, 65.4011, 47.57902, 
    52.56764, 62.57636, 88.29622, 103.0397, 116.2788, 146.1452, 149.0459, 
    260.9405, 209.8252, 240.3782, 305.7633, 380.0433, 410.2039, 401.1645, 
    344.6812, 350.6726, 420.6497, 639.9168, 1359.416, 1773.189, 1596.877, 
    1193.995, 945.0976, 478.8944, 313.0052, 364.5321, 544.9355, 728.1349, 
    913.1708, 1094.162, 1205.655, 1103.695, 1186.761, 1181.66, 1198.702, 
    1409.169, 1265.896, 1273.084, 1305.134, 1441.755, 1591.454, 1519.917, 
    1441.886, 1330.869, 1070.649, 1189.587, 1315.408, 1415.29, 1531.97, 
    1529.214, 1473.449, 1430.014, 1306.896, 1270.828, 872.1915, 165.6583, 
    2.112291, 1.155395, 0.02070807, 0.08559992, 13.39372, 105.9956, 72.41502, 
    2.817191, 0, 0, 0.04834903,
  0.02893994, 4.580082, 170.3799, 581.9701, 947.2767, 1071.069, 1146.666, 
    1154.808, 1640.017, 1900.844, 1998.073, 1884.909, 1641.079, 1859.79, 
    780.6656, 620.8061, 1727.327, 225.5852, -29, -29, -29, 38.14354, 
    126.9196, 155.8592, 184.8903, 179.1412, 129.6505, 97.10344, 37.13656, 
    33.23013, 51.04347, 71.70508, 91.74311, 103.1298, 126.9913, 145.6968, 
    179.7494, 230.5837, 298.0778, 375.3928, 434.7722, 459.8557, 350.7677, 
    343.3709, 347.6726, 356.1186, 381.6495, 446.8376, 603.9845, 758.576, 
    881.1244, 1095.882, 904.9011, 568.9519, 433.0408, 654.4484, 862.9261, 
    1147.874, 1391.479, 1546.497, 1694.146, 1655.956, 1846.877, 1863.535, 
    1773.414, 1861.801, 1658.115, 1432.014, 1446.591, 1505.779, 1598.366, 
    1639.378, 1501.092, 1183.134, 1002.323, 1205.448, 1280.397, 1347.836, 
    1565.089, 1583.707, 1551.659, 1326.685, 1098.686, 688.5358, 124.0418, 
    3.131963, 2.67241, 0, 0, 0.3741298, 0, 14.65283, 0, 0, 0, 0.08931515,
  735.5396, 867.0506, 660.6748, 924.9462, 1301.789, 1480.976, 1317.01, 
    1341.343, 1806.828, 2025.722, 2183.452, 2051.318, 1930.586, 1732.126, 
    665.5182, 1034.291, 2036.85, 544.5954, -29, -29, -28.76467, 38.63471, 
    172.218, 155.2569, 183.3024, 142.7022, 156.3304, 131.9387, 71.52921, 
    29.83442, 38.42982, 63.1153, 82.10826, 123.0225, 117.6491, 159.6424, 
    210.2419, 265.2799, 324.6303, 429.2385, 526.7354, 552.8436, 445.1412, 
    408.4677, 410.2799, 482.5757, 457.1882, 425.4275, 467.3434, 724.1971, 
    978.342, 1341.993, 1428.619, 1158.37, 714.2965, 634.1248, 1100.511, 
    1729.557, 2079.457, 2205.601, 2096.228, 1923.082, 2023.244, 2032.364, 
    2087.194, 1819.859, 1741.359, 1652.907, 1411.046, 1353.822, 1332.2, 
    1373.966, 1373.264, 1169.126, 951.4221, 1059.032, 1129.511, 1144.062, 
    1270.443, 1435.999, 1450.52, 1447.836, 1236.854, 758.832, 350.9756, 
    181.3987, 25.64147, 0, 7.676435, 3.285792, 0, 0, 0, 0, 4.333813, 55.45658,
  1304.387, 1437.602, 1376.26, 1494.452, 1659.236, 1723.898, 1639.994, 
    1657.578, 1850.001, 2092.416, 1922.954, 1856.68, 1913.263, 1612.252, 
    1244.188, 1688.415, 1823.349, 597.8655, -28.95335, -29, -29, 36.93167, 
    126.3385, 56.37119, 89.7822, 66.37797, 91.53525, 123.4684, 92.97884, 
    64.8284, 57.79882, 59.7579, 86.7978, 105.0893, 148.6383, 195.5772, 
    329.0817, 307.0089, 342.0926, 436.9752, 591.1713, 694.5746, 679.3177, 
    636.2111, 632.0756, 646.1209, 669.288, 648.6287, 782.5434, 883.3128, 
    793.3741, 676.8798, 926.3399, 801.6874, 746.4554, 1202.792, 1920.346, 
    2443.33, 2322.053, 1982.287, 1837.848, 1673.851, 1988.25, 2200.716, 
    1986.238, 1899.81, 1884.782, 1790.649, 1548.873, 1296.591, 1256.828, 
    1255.077, 1205.229, 1093.803, 927.5923, 972.8065, 1059.568, 1028.104, 
    1103.09, 1202.041, 1344.654, 1430.761, 1304.095, 857.4107, 614.5168, 
    408.0826, 142.5798, 1.184603, 40.65562, 3.480806, 0, 1.402507, 22.73934, 
    1.869505, 22.95708, 208.0578,
  1176.996, 1274.15, 1167.862, 1260.973, 1305.267, 1444.57, 1547.88, 
    1561.639, 1724.48, 1392.404, 542.0779, 297.3251, 709.7617, 908.8043, 
    1689.685, 1619.551, 990.7944, 115.7064, -24.46063, -28.99723, -29, 11.77, 
    -18.20284, -18.30782, -26.05886, -15.76914, 55.73129, 98.28559, 125.4715, 
    138.3384, 126.8703, 111.3977, 77.0961, 90.02938, 117.3675, 253.6755, 
    387.6956, 435.0849, 377.246, 411.8622, 531.7675, 673.597, 770.8846, 
    853.8765, 854.3976, 850.265, 792.6041, 745.4413, 733.783, 735.1926, 
    603.2223, 591.2675, 993.4567, 1367.18, 1860.522, 2238.518, 2511.91, 
    2284.058, 1663.224, 1322.216, 1438.35, 1776.375, 2169.013, 2455.426, 
    2488.388, 2387.191, 2351.167, 2100.744, 1704.273, 1439.597, 1375.393, 
    1281.368, 1147.538, 1084.584, 931.0007, 951.1368, 1033.676, 1018.033, 
    1023.891, 1108.402, 1268.471, 1365.725, 1364.301, 974.9635, 739.7955, 
    399.5302, 73.64684, 12.84806, 147.529, 5.471954, 0, 24.00544, 116.3721, 
    114.7116, 240.0056, 341.1817,
  1120.788, 1306.315, 1094.511, 1054.712, 1080.561, 1158.717, 1213.522, 
    1205.066, 948.7064, 166.4328, 0, 0, 7.011492, 766.0705, 1910.302, 
    1318.522, 220.8738, 20.13437, -22.87948, -28.96292, -28.99967, -28.96005, 
    -28.95333, -28.95845, -28.27328, -19.16533, 25.35257, 78.57539, 126.1784, 
    178.1593, 206.8317, 152.6626, 97.64114, 76.05511, 110.28, 209.1862, 
    385.8008, 487.759, 490.3545, 435.6064, 477.5195, 573.1337, 679.9717, 
    815.3858, 863.851, 795.056, 638.4842, 521.1765, 490.9408, 599.1897, 
    654.6764, 994.7811, 1491.828, 2086.955, 2473.281, 2589.081, 2203.682, 
    1937.777, 1327.908, 1322.338, 1643.389, 1980.04, 2347.152, 2586.005, 
    2474.671, 2249.25, 1973.765, 1742.107, 1577.967, 1488.696, 1454.051, 
    1334.462, 1222.04, 1055.741, 975.7679, 973.0269, 1098.012, 1137.429, 
    1093.573, 1125.746, 1300.224, 1360.541, 1194.296, 881.052, 581.177, 
    281.8254, 19.61534, 84.07046, 212.6468, 69.3125, 29.19267, 158.5775, 
    304.7471, 402.8232, 454.9509, 428.1056,
  1187.477, 1316.139, 1129.726, 991.171, 1030.374, 1016.187, 1020.988, 
    818.59, 381.7968, 0, 0, 0, 0, 1129.767, 1979.666, 998.5098, 264.3186, 
    59.78041, -4.723167, -24.42554, -28.50731, -28.65225, -28.92911, -29, 
    -28.607, -24.37205, 20.2152, 104.2612, 164.2149, 231.1236, 260.2584, 
    221.0597, 141.5681, 105.8174, 115.9729, 151.8276, 274.3087, 439.8468, 
    448.8825, 399.3673, 408.2239, 453.6656, 569.141, 609.5902, 626.4427, 
    521.6019, 365.9188, 284.7949, 285.1086, 423.1974, 846.5926, 1237.006, 
    1726.326, 2102.346, 2434.645, 2372.822, 2198.263, 1666.205, 1424.405, 
    1409.403, 1744.127, 2013.176, 2073.452, 2140.749, 2030.338, 1827.267, 
    1580.342, 1325.149, 1298.67, 1349.97, 1428.83, 1395.826, 1250.978, 
    1179.868, 1037.025, 1015.187, 1152.761, 1271.608, 1141.957, 1128.437, 
    1250.247, 1118.777, 820.3528, 513.1799, 459.0807, 201.0253, 50.98212, 
    173.3005, 353.3956, 272.952, 377.204, 340.7662, 338.8821, 282.7307, 
    42.52118, 0,
  911.2604, 1162.884, 1137.084, 979.4952, 1010.004, 1126.895, 1059.642, 
    869.5664, 252.7621, 0, 0, 0, 0, 1150.678, 1275, 595.7617, 273.573, 
    133.9935, 32.51972, -16.08583, -22.48619, -23.88273, -23.75681, 
    -24.06026, -24.22806, -20.21073, 10.21312, 100.5829, 164.7874, 248.1127, 
    306.6323, 287.0247, 220.7695, 169.7234, 135.2546, 137.2507, 172.6728, 
    311.0542, 341.0001, 327.2497, 348.4995, 425.6412, 463.1763, 447.4398, 
    353.7435, 252.8357, 186.9208, 193.5265, 269.0485, 416.4105, 833.4974, 
    1255.776, 1478.953, 1658.504, 2096.166, 2288.637, 1723.026, 1429.502, 
    949.519, 1162.872, 1667.993, 1924.058, 2051.646, 1868.885, 1679.083, 
    1502.363, 1410.3, 1248.582, 1158.49, 1393.645, 1598.457, 1420.972, 
    1293.249, 1159.699, 1133.274, 1037.51, 1155.602, 1250.937, 1090.242, 
    1007.832, 1146.141, 923.0365, 519.2554, 340.7791, 297.567, 152.0113, 
    84.55415, 319.1597, 474.4228, 619.5093, 846.3072, 366.6542, 0.09596219, 
    0, 0, 0,
  612.0165, 1024.829, 1129.861, 947.5595, 1080.557, 1194.547, 1150.219, 
    904.1955, 156.9333, 0, 0, 0, 0, 583.678, 439.6959, 309.7408, 232.4993, 
    133.5744, 75.71014, -1.082752, -7.73104, -16.27212, -16.11549, -15.90899, 
    -15.91451, -10.86247, 4.381418, 61.24113, 156.1658, 234.102, 316.4874, 
    335.1181, 275.5302, 255.234, 212.9649, 181.6552, 180.8939, 256.1131, 
    302.8167, 311.314, 343.6282, 353.8376, 353.0165, 257.5091, 195.26, 
    136.4342, 132.6939, 165.401, 204.5192, 263.7407, 417.9625, 651.0251, 
    757.1484, 1176.346, 1630.802, 1775.998, 1641.073, 1216.329, 1179.213, 
    1361.391, 1647.038, 1987.515, 2015.377, 1927.813, 1564.168, 1375.637, 
    1276.543, 1056.094, 1081.178, 1433.004, 1697.667, 1528.249, 1249.511, 
    1163.054, 1084.624, 1005.993, 992.0644, 1018.707, 950.4731, 940.6085, 
    1033.09, 798.034, 387.972, 229.6093, 197.4241, 132.7397, 211.0327, 
    408.1602, 644.9759, 902.4259, 1280.562, 421.0834, 0, 0, 0, 0,
  358.6493, 740.4105, 851.3992, 682.4423, 613.3671, 561.9201, 439.3097, 
    284.2988, 0, 0, 0, 0, 0, 164.7004, 99.19429, 101.628, 107.9559, 74.77886, 
    89.1244, 63.77163, 1.608809, -6.549558, -9.00685, -8.677175, -9.026371, 
    -3.706912, 1.230656, 51.11661, 139.9139, 209.1897, 282.7745, 328.7339, 
    305.7128, 303.4295, 269.2504, 220.6103, 194.5171, 252.9004, 301.2274, 
    362.1626, 362.2566, 319.3198, 217.928, 137.8181, 105.979, 105.6061, 
    114.0887, 135.0031, 185.067, 190.351, 191.2327, 234.4863, 323.938, 
    543.4288, 1060.478, 1268.447, 1192.681, 1328.727, 1228.022, 1216.701, 
    1586.167, 1872.411, 2054.413, 1874.194, 1613.623, 1458.215, 1250.402, 
    935.8388, 937.23, 1296.085, 1562.618, 1421.365, 1164.499, 1045.977, 
    969.0322, 885.1325, 801.2127, 811.7344, 891.5575, 953.3035, 938.8203, 
    644.8547, 285.5817, 157.9158, 154.0628, 172.5158, 282.7875, 469.8745, 
    706.7769, 1102.511, 1230.183, 277.3174, 0, 0, 0, 0,
  132.9001, 385.4105, 339.2654, 181.7644, 142.398, 0.8909621, 0, 0, 0, 0, 0, 
    0, 4.920471, 45.10483, 8.741613, 47.47253, 68.29308, 52.40722, 93.38539, 
    77.34655, 43.84061, 4.212869, 4.007848, 10.19131, 4.169814, 0.9422171, 
    9.296235, 56.39237, 118.7264, 170.1291, 210.7619, 320.4744, 331.2771, 
    318.584, 273.9849, 219.1942, 178.2944, 198.5368, 260.3773, 310.2903, 
    314.4893, 238.4738, 144.5557, 99.9539, 97.97208, 100.8626, 114.6869, 
    130.8342, 169.4516, 185.3304, 185.0731, 235.592, 278.8924, 478.6136, 
    764.5692, 685.5565, 811.843, 974.8875, 1184.866, 1309.973, 1492.49, 
    1975.901, 2111.276, 1920.701, 1584.152, 1393.754, 1227.47, 867.7672, 
    863.7648, 1180.989, 1434.811, 1408.729, 1119.982, 937.4036, 832.1047, 
    725.7586, 654.3876, 681.5729, 879.4352, 1001.297, 813.8375, 472.1414, 
    186.7852, 145.5977, 173.9421, 209.2027, 326.0379, 476.7007, 804.9005, 
    1109.927, 922.321, 75.55848, 0, 0, 0, 0,
  55.06753, 268.7123, 117.1969, 34.0993, 31.63307, 0, 0, 0, 0, 0, 75.30566, 
    123.2075, 25.73137, 4.677011, 0.4355646, 21.74989, 39.51146, 59.60038, 
    56.39664, 83.5396, 72.77475, 42.05199, 25.05266, 18.50826, 21.90979, 
    18.97606, 32.88521, 52.70894, 108.0705, 133.6327, 212.1806, 346.0227, 
    454.2986, 381.998, 286.2616, 211.4252, 172.9534, 157.5838, 173.7746, 
    195.4111, 173.0165, 139.0157, 104.9335, 99.12243, 103.3306, 100.5489, 
    103.4557, 134.8257, 162.8266, 185.8695, 232.4137, 269.2041, 308.7599, 
    614.8231, 747.6427, 544.698, 422.7588, 738.6674, 1183.856, 1471.337, 
    1606.683, 1839.523, 1757.208, 1367.475, 928.4243, 840.8771, 759.8136, 
    793.3425, 873.0726, 1079.337, 1313.67, 1351.702, 1047.42, 866.4039, 
    745.4284, 686.4276, 600.6986, 676.6058, 942.1893, 1006.475, 678.2116, 
    313.3897, 146.0503, 136.1638, 173.3874, 203.2215, 423.4491, 556.2217, 
    687.7593, 707.8784, 130.9646, 0, 0, 0, 0, 0,
  7.121133, 32.15426, 84.65013, 100.6684, 128.3299, 0, 0, 0, 0, 0, 37.53299, 
    141.1044, 20.04803, 0.0226125, 4.211974, 29.80108, 80.3756, 118.8334, 
    109.4529, 114.3332, 124.4319, 101.2349, 79.91515, 62.1116, 42.87167, 
    62.06577, 74.78121, 105.4743, 125.4183, 177.7379, 223.2901, 362.0724, 
    497.8951, 520.5967, 347.3084, 218.1198, 160.7832, 142.836, 141.2242, 
    142.3133, 130.3157, 119.2133, 114.2978, 107.0357, 102.9367, 104.6058, 
    110.6453, 123.0354, 142.3407, 155.8816, 175.0349, 218.0002, 336.6488, 
    481.0204, 622.3756, 464.2339, 567.8765, 821.3962, 1203.486, 1431.367, 
    1332.833, 1153.785, 908.6243, 652.9219, 598.5366, 569.8493, 665.6304, 
    778.8425, 895.4351, 980.2097, 1137.299, 1139.964, 917.5201, 727.8011, 
    697.3036, 645.4094, 611.8453, 750.6511, 997.3835, 898.4934, 452.9046, 
    187.9874, 131.9667, 132.1604, 162.3042, 257.2846, 519.6144, 578.7543, 
    534.0048, 299.177, 10.42934, 0, 0, 0, 0, 0,
  29.01102, 22.0339, 235.5383, 205.7878, 202.3339, 34.00895, 0, 0, 0, 0, 
    0.7499724, 39.96126, 8.142411, 27.61915, 77.46246, 141.4588, 165.7684, 
    167.3914, 132.9326, 131.5184, 138.1546, 130.3924, 147.073, 128.6659, 
    88.82133, 71.90593, 79.99207, 93.95091, 122.2475, 174.1009, 224.5994, 
    264.6025, 432.1731, 552.0823, 489.6333, 281.8752, 171.4949, 136.2069, 
    133.1193, 125.4225, 126.965, 120.7626, 111.4299, 101.8144, 99.97607, 
    113.2573, 118.6737, 130.7982, 136.456, 127.7007, 138.2258, 178.1324, 
    196.5107, 345.3022, 326.9236, 389.049, 456.8989, 544.9363, 644.9791, 
    795.9853, 714.1006, 626.2784, 512.6625, 545.9469, 686.3776, 774.8943, 
    722.8535, 808.6535, 999.6533, 978.3033, 988.0608, 965.1602, 774.5897, 
    743.5015, 720.1992, 658.6784, 645.7189, 780.3297, 934.1503, 668.8269, 
    269.4187, 138.0441, 142.1439, 151.7155, 169.5889, 303.9595, 540.4365, 
    608.5374, 528.3405, 294.674, 2.237589, 0, 0, 0, 0, 0,
  111.4144, 193.5326, 681.5145, 360.9993, 352.8302, 226.3572, 174.55, 
    37.86699, 0.2644904, 0.002788612, 0, 3.079878, 23.88782, 46.11481, 
    80.04777, 123.263, 147.1195, 144.2522, 130.5605, 152.2023, 141.6269, 
    132.931, 157.0246, 184.9375, 164.1916, 154.953, 124.2921, 92.66442, 
    103.1418, 164.1006, 233.3318, 178.8902, 210.3269, 409.1046, 418.7644, 
    336.8872, 189.2744, 130.1919, 111.7867, 105.783, 110.7427, 102.534, 
    94.83035, 91.60812, 107.021, 117.6856, 130.0774, 128.3777, 127.6499, 
    111.2988, 106.9357, 137.1521, 166.8579, 176.284, 241.0266, 287.8779, 
    322.1338, 316.6681, 333.3232, 405.2602, 465.2554, 453.8713, 526.2246, 
    631.4445, 775.7401, 794.0515, 706.1703, 873.7288, 1141.089, 1067.214, 
    1009.558, 878.1597, 765.5309, 814.0995, 825.5641, 682.4036, 688.0043, 
    821.9866, 793.0577, 482.589, 210.6379, 172.7338, 171.0665, 163.2869, 
    239.3744, 290.9917, 518.2194, 476.0343, 344.188, 253.0163, 199.3618, 
    0.09988576, 0, 0, 0, 0,
  396.4076, 461.4612, 931.6284, 727.4689, 459.6009, 316.0923, 161.0612, 
    61.08897, 39.84538, 14.21865, 16.21696, 14.69456, 42.59837, 83.79881, 
    96.42057, 106.7112, 127.726, 139.3746, 149.1176, 158.2953, 146.0142, 
    133.0698, 149.0564, 185.547, 219.5478, 236.7041, 204.2428, 142.1788, 
    111.0571, 152.1457, 197.096, 162.3448, 145.3164, 257.3849, 359.7718, 
    344.883, 231.0725, 134.1741, 96.72655, 77.17216, 67.97431, 71.95205, 
    78.97033, 92.42341, 106.5057, 121.7666, 113.3711, 112.7681, 100.1774, 
    90.3449, 93.89151, 126.1822, 144.4522, 167.8977, 184.3656, 222.1504, 
    216.4159, 276.5192, 273.3236, 330.4809, 405.03, 466.5895, 519.9902, 
    669.0401, 778.4682, 755.4747, 760.0569, 995.1483, 1292.865, 1133.658, 
    1035.321, 891.3419, 745.2759, 794.439, 820.8765, 731.4034, 825.5676, 
    816.8707, 654.7597, 365.2853, 254.1914, 241.2478, 251.6084, 300.0577, 
    283.1929, 314.035, 356.0846, 297.13, 224.8416, 403.2619, 439.1473, 
    0.3467962, 0, 0, 0, 0,
  855.1598, 709.2625, 1002.592, 837.1132, 519.1252, 130.5939, 71.12158, 
    81.11422, 142.1018, 51.00807, 96.93317, 79.51467, 95.48483, 129.0423, 
    140.4562, 103.5044, 126.4621, 151.7047, 177.8282, 174.2761, 156.9096, 
    144.2187, 154.5808, 180.015, 203.6465, 223.6183, 210.2678, 151.1036, 
    112.8854, 117.9561, 134.9364, 127.8695, 129.1225, 218.7797, 270.9187, 
    350.6521, 238.6366, 134.1218, 93.92628, 66.70253, 59.81225, 64.58974, 
    83.67481, 91.74277, 99.39961, 97.78426, 98.12943, 79.38904, 76.33865, 
    79.66943, 96.24992, 117.7307, 139.8467, 146.7351, 147.0995, 206.1468, 
    254.7715, 275.4333, 300.4858, 331.8605, 412.4602, 458.4528, 508.2016, 
    647.9883, 697.1085, 851.0264, 924.2222, 1209.887, 1389.744, 1105.53, 
    981.9774, 946.9201, 772.724, 746.0531, 774.8968, 822.0195, 896.6089, 
    762.1265, 469.3407, 356.1171, 319.8726, 356.8423, 393.546, 402.3568, 
    300.6212, 214.0752, 218.7073, 138.1364, 184.7563, 493.152, 362.86, 0, 0, 
    0, 0, 0,
  886.0403, 899.0963, 842.0179, 772.5779, 432.9344, 92.04449, 177.5087, 
    546.1584, 477.8832, 337.027, 119.8037, 133.9722, 151.3862, 176.6996, 
    157.914, 107.5661, 123.6268, 163.6318, 191.2482, 207.9477, 183.4089, 
    166.7186, 150.5348, 152.3792, 164.6893, 178.3489, 177.4384, 146.3247, 
    116.5272, 132.4336, 138.0589, 139.9558, 167.7014, 180.2253, 221.528, 
    303.055, 258.0195, 122.0804, 91.42705, 76.97997, 52.65008, 55.3461, 
    72.29636, 81.25592, 81.83448, 87.9664, 75.1608, 69.10935, 76.35617, 
    101.0703, 128.3883, 140.7466, 138.2242, 132.6284, 251.6389, 360.3346, 
    363.8312, 345.4504, 282.5562, 300.7509, 352.1882, 428.2724, 480.032, 
    508.1172, 638.3249, 969.0288, 1175.973, 1303.747, 1379.587, 1075.456, 
    939.7833, 971.2458, 876.7556, 679.537, 703.0974, 840.0677, 888.4769, 
    685.1582, 465.5422, 392.8445, 362.4918, 364.3657, 413.9269, 386.9064, 
    151.63, 102.4381, 140.1844, 97.34532, 357.6024, 508.7825, 100.0093, 0, 0, 
    0, 0.4358488, 0,
  377.0912, 777.9293, 847.1389, 613.7839, 347.3856, 183.928, 503.8705, 
    767.5604, 736.3063, 591.572, 261.3434, 142.1519, 203.053, 216.3297, 
    177.3449, 117.8392, 131.8621, 155.6192, 186.6643, 210.5387, 213.1024, 
    198.3484, 171.8902, 133.9252, 133.7206, 147.76, 149.0784, 123.2078, 
    117.5802, 128.9419, 142.8373, 162.3329, 190.3584, 196.8235, 191.6556, 
    277.8559, 336.0329, 136.4615, 78.44816, 67.13183, 57.19013, 45.63347, 
    56.64672, 62.35668, 62.41399, 58.50655, 64.08222, 61.68793, 82.98176, 
    109.022, 132.2926, 141.4133, 130.0148, 202.6298, 352.5894, 478.8041, 
    483.1053, 383.9174, 324.0171, 288.2619, 333.3291, 429.6476, 498.3948, 
    476.5586, 511.4784, 972.3265, 1117.176, 1333.446, 1231.988, 1100.885, 
    955.795, 961.8926, 865.2928, 707.8149, 605.3251, 700.6523, 739.4321, 
    558.5131, 402.4283, 297.584, 211.9652, 189.1523, 300.2366, 262.1036, 
    80.62009, 63.98812, 122.1838, 218.2967, 512.9334, 462.9636, 1.060671, 0, 
    0, 0, 37.38868, 81.3967,
  0, 594.21, 1018.811, 745.1058, 412.2401, 385.4236, 638.6064, 788.1194, 
    668.9521, 749.03, 562.7498, 197.1136, 243.5414, 257.3966, 197.9897, 
    130.8538, 123.876, 145.1576, 174.6566, 198.9581, 214.8165, 215.6441, 
    189.8338, 139.6603, 120.3094, 124.8503, 116.1674, 109.7017, 110.3707, 
    135.235, 142.0241, 170.4792, 213.9434, 209.5347, 167.4813, 264.8561, 
    348.0725, 240.3373, 75.87767, 79.91491, 71.83314, 45.36616, 48.33675, 
    52.77137, 49.97958, 59.72789, 63.37616, 71.72295, 88.81493, 109.8572, 
    136.8765, 144.6113, 151.7365, 193.6578, 319.4838, 403.0927, 398.4877, 
    411.3876, 349.0669, 324.9615, 351.6237, 448.8545, 494.1817, 457.7076, 
    444.8627, 679.2474, 972.8405, 1012.391, 1150.945, 1145.6, 1127.534, 
    944.8821, 822.8835, 703.0647, 531.0294, 464.5009, 428.4065, 363.7079, 
    263.4396, 211.7635, 198.9796, 267.8853, 350.3128, 264.7803, 65.758, 
    59.44502, 199.1785, 430.2982, 657.9562, 212.0221, 0, 0, 0, 97.63541, 
    113.3308, 41.61473,
  0, 399.1143, 1120.441, 820.4569, 297.3376, 195.9688, 434.3469, 519.7678, 
    533.1642, 758.1817, 711.3763, 342.4791, 278.5041, 278.4136, 214.2995, 
    149.314, 124.3232, 138.1995, 163.2455, 188.7315, 200.2267, 205.1242, 
    191.2654, 153.1303, 140.5527, 120.2366, 117.1466, 119.59, 127.6191, 
    134.2686, 149.6515, 164.0252, 186.4469, 196.4661, 161.6761, 177.2666, 
    334.9556, 307.35, 143.2057, 109.0354, 87.71973, 79.37965, 65.37148, 
    76.016, 76.0844, 78.8138, 85.20406, 92.65923, 120.6024, 124.1407, 
    141.3281, 120.2449, 152.1772, 252.603, 380.783, 423.7603, 464.9473, 
    420.7524, 383.9003, 365.9595, 382.3451, 404.967, 427.5276, 426.6728, 
    395.3827, 540.5605, 755.1957, 952.8699, 1084.376, 1365.629, 1383.233, 
    963.2598, 743.7776, 748.3361, 583.3853, 439.8699, 330.5274, 274.6473, 
    239.082, 218.2501, 375.178, 416.6259, 488.4598, 300.3638, 65.87481, 
    54.1222, 354.7472, 673.2607, 622.6516, 29.62266, 0, 0, 0, 206.3307, 
    149.5761, 0,
  0.003310259, 133.1911, 940.6332, 781.675, 248.0849, 90.08338, 116.6424, 
    220.5476, 304.2039, 419.5131, 703.8474, 411.9249, 301.6213, 267.3719, 
    209.3017, 160.7548, 131.8181, 134.4422, 157.0661, 185.6122, 207.0094, 
    210.453, 201.0542, 179.5661, 159.3497, 148.5723, 124.2159, 138.4398, 
    148.6608, 162.3591, 173.3146, 175.035, 184.1364, 181.5239, 173.0168, 
    157.8075, 250.5602, 304.8704, 179.2655, 67.08978, 85.99716, 73.47701, 
    103.1553, 107.7299, 100.9882, 96.31065, 80.26945, 83.55797, 94.24591, 
    113.5028, 87.01515, 83.67673, 216.3896, 356.1998, 462.2934, 496.7366, 
    464.9568, 424.9034, 395.8524, 405.8656, 396.2522, 369.3352, 362.0952, 
    392.2811, 403.4277, 532.8717, 897.1837, 937.3101, 997.2128, 1238.674, 
    1234.297, 916.9507, 798.6755, 785.5186, 683.3135, 527.7955, 404.3859, 
    329.3802, 251.766, 331.9852, 519.2047, 603.6315, 693.9681, 306.4999, 
    50.3644, 206.1701, 627.575, 741.8391, 292.8152, 0, 0, 0.002287545, 
    47.08162, 366.3271, 345.8133, 140.5091,
  0.1355318, 54.76622, 752.4495, 779.2272, 233.4452, 90.45777, 81.94717, 
    83.38457, 113.8429, 180.5548, 517.6541, 398.6514, 294.062, 222.6104, 
    177.3117, 146.8111, 135.3791, 142.748, 161.5963, 189.4258, 213.6966, 
    218.6755, 216.248, 169.9221, 153.2071, 133.3895, 136.4664, 149.2455, 
    169.6985, 177.9319, 169.0834, 158.8819, 153.8374, 154.3419, 155.6863, 
    159.3348, 168.2593, 263.9666, 210.4024, 63.44218, 42.57559, 53.28033, 
    74.75113, 94.46678, 84.90047, 77.8112, 56.29344, 41.15648, 64.81905, 
    77.03599, 86.15321, 102.1669, 314.0604, 390.679, 394.7146, 406.8066, 
    419.1735, 403.4146, 401.5237, 394.1876, 379.7701, 337.2509, 349.9233, 
    401.1396, 396.1155, 511.2408, 755.8575, 709.9775, 686.9054, 793.6512, 
    1004.453, 980.0493, 971.1741, 917.5543, 726.7474, 512.3557, 394.0262, 
    441.8013, 404.3204, 456.4452, 727.2965, 845.9907, 812.4409, 408.3134, 
    83.84931, 448.7415, 730.8319, 467.4902, 0.9863583, 0, 1.720724, 35.83591, 
    297.3234, 472.4654, 318.6473, 2.667824,
  2.786609, 2.644013, 504.1062, 684.3657, 243.8393, 124.4904, 120.2434, 
    118.8162, 136.5323, 274.2844, 459.7988, 323.3001, 252.3182, 197.7955, 
    158.2456, 143.8349, 155.14, 171.036, 179.7861, 181.361, 194.9534, 
    211.9559, 228.9097, 199.0386, 153.3901, 145.1039, 136.1797, 149.812, 
    166.3282, 157.6181, 154.2063, 126.907, 146.2792, 140.0006, 147.5358, 
    162.919, 152.3721, 222.5984, 246.1506, 256.06, 62.73549, 34.49001, 
    46.63019, 67.38826, 49.56528, 57.15746, 51.01564, 36.49106, 33.8912, 
    64.45266, 63.10199, 144.3528, 351.2276, 400.1565, 401.1474, 439.6917, 
    469.2003, 431.5126, 411.8654, 369.9917, 321.8169, 323.1301, 326.4559, 
    382.4082, 378.7637, 344.4705, 461.5488, 414.4735, 376.186, 542.0886, 
    713.6682, 832.4791, 967.1309, 1007.369, 852.7335, 704.9957, 550.9443, 
    581.854, 539.4864, 852.6191, 1003.918, 778.0033, 665.1097, 266.5093, 
    311.5761, 683.8643, 705.9689, 96.01817, 0, 1.189999, 8.842051, 47.33828, 
    140.6496, 324.6157, 137.269, 0,
  276.4731, 0, 179.3712, 525.0765, 251.7486, 132.691, 157.0414, 154.7416, 
    302.1239, 580.2548, 583.1707, 323.0918, 206.9382, 174.8136, 156.9467, 
    158.7047, 172.3876, 199.9602, 184.0974, 164.6234, 165.0962, 185.8372, 
    203.0004, 193.7835, 175.1679, 146.9807, 142.3714, 150.1652, 157.6037, 
    163.3478, 129.6109, 129.2951, 159.414, 161.3647, 162.9705, 181.9612, 
    128.0042, 147.4346, 353.2044, 345.6928, 272.2606, 81.65241, 31.30544, 
    29.65827, 24.55814, 44.82172, 50.73238, 36.99446, 29.24441, 45.64774, 
    56.69508, 147.8097, 350.2406, 446.015, 517.4972, 568.1435, 509.0543, 
    480.6918, 464.3664, 407.0969, 359.9652, 325.3537, 336.1723, 338.7549, 
    334.156, 299.1234, 313.2734, 332.2038, 383.9116, 472.8965, 632.2615, 
    813.0618, 1026.41, 1103.619, 1136.821, 1031.338, 975.8419, 689.2612, 
    568.7227, 943.745, 852.9982, 485.5357, 236.3455, 271.7433, 463.5656, 
    614.2126, 345.1251, 0, 16.48282, 105.6186, 7.521848, 0, 0, 87.10019, 
    40.73374, 0,
  508.8716, 70.13601, 6.784113, 372.3694, 322.6259, 293.2125, 242.353, 
    173.0082, 268.3181, 591.1161, 536.0643, 296.8539, 202.5906, 164.5604, 
    144.654, 150.5097, 161.7568, 165.6213, 170.2032, 147.5072, 145.3487, 
    118.8593, 111.2818, 111.6931, 136.4204, 155.4414, 171.5328, 140.8391, 
    169.3844, 138.0114, 124.348, 104.4207, 145.8794, 164.8125, 186.8414, 
    188.481, 126.0499, 90.26923, 110.4248, 252.1565, 185.2361, 152.9825, 
    177.3863, 27.33101, 14.74302, 22.59383, 32.78283, 24.52886, 36.56748, 
    50.80676, 80.63863, 201.0317, 398.6272, 570.3611, 631.2753, 643.4182, 
    537.705, 514.1293, 540.4216, 502.6988, 444.1647, 409.5107, 358.6469, 
    313.3456, 229.5331, 227.212, 262.0572, 326.5652, 403.6352, 469.1498, 
    543.0381, 673.6775, 820.8776, 1047.744, 949.5495, 1148.552, 1111.228, 
    855.2848, 484.6896, 661.6188, 513.8441, 249.184, 299.0674, 415.421, 
    493.6745, 252.4404, 5.99207, 59.10885, 97.5045, 79.21317, 10.46941, 0, 0, 
    43.29576, 3.355622, 0,
  443.5912, 255.1915, 0.09644534, 195.873, 487.8073, 735.0255, 695.2324, 
    348.3268, 280.6532, 412.6371, 385.954, 220.2776, 204.6375, 127.3774, 
    125.8829, 139.0522, 124.0497, 124.0424, 125.5306, 122.1397, 132.0455, 
    96.83639, 60.97416, 63.26183, 70.19158, 96.56532, 138.9745, 127.6716, 
    134.1593, 150.0386, 90.46266, 84.52273, 112.2292, 121.4295, 151.5019, 
    166.1176, 108.1869, 79.91405, 92.42285, 97.96801, 124.7679, 221.8664, 
    228.2843, 115.3288, 24.56494, 14.8802, 20.65261, 31.73664, 49.24442, 
    60.99174, 105.08, 244.0706, 521.9723, 723.241, 767.3787, 664.4177, 
    487.5122, 513.0247, 515.0753, 538.3448, 511.0675, 463.2043, 376.3399, 
    264.3518, 201.9225, 193.3568, 293.2623, 334.261, 373.6343, 439.8721, 
    490.5887, 493.9969, 600.4854, 755.9476, 924.3199, 950.3077, 1052.388, 
    779.1483, 183.5563, 265.7245, 179.8311, 213.6126, 282.3783, 202.5462, 
    128.2361, 30.74742, 219.925, 102.526, 0, 0, 0, 0, 0, 16.26684, 0.6956787, 0,
  260.7036, 393.7766, 11.27141, 23.8249, 678.2915, 1205.305, 983.3217, 
    600.5497, 405.7943, 426.7081, 384.4165, 217.486, 141.1087, 113.0105, 
    118.703, 126.1676, 90.83533, 74.9175, 85.22266, 86.1847, 108.5499, 
    97.74491, 85.57736, 64.07814, 40.13272, 24.09916, 78.24743, 80.76043, 
    124.5104, 132.6886, 90.25305, 50.69267, 81.38572, 64.80839, 89.60198, 
    115.1036, 102.3747, 89.09599, 91.98434, 106.8285, 90.62163, 137.0851, 
    183.7695, 40.38134, 27.67106, 11.31515, 23.2658, 37.70986, 46.24703, 
    62.2045, 86.09678, 336.5412, 717.0566, 919.0491, 854.2428, 596.1452, 
    380.2888, 384.9098, 468.5178, 498.7417, 522.8006, 451.6152, 351.5222, 
    233.9609, 161.0052, 184.1114, 234.4022, 294.4582, 302.137, 342.4128, 
    411.9693, 392.7577, 351.6703, 590.9839, 653.2507, 725.2677, 801.4582, 
    656.3619, 55.66471, 28.70166, 97.66091, 137.6178, 146.7572, 75.24693, 
    99.51981, 291.1764, 193.6622, 6.543282, 0, 0, 0, 0, 10.53877, 52.14492, 
    0, 0,
  43.77597, 464.1584, 56.89383, 468.3003, 1272.138, 1580.384, 1018.172, 
    560.8243, 492.4376, 414.2195, 387.2528, 175.9947, 96.38813, 88.09875, 
    109.2793, 71.96533, 25.01822, 58.2986, 73.01802, 38.57325, 49.70271, 
    62.90857, 57.06133, 27.90662, 27.32676, 23.32841, 78.08787, 112.5397, 
    118.9064, 113.533, 66.1688, 38.50869, 78.81353, 50.76294, 38.3057, 
    62.43602, 80.58298, 45.74772, 40.23263, 38.5184, 22.24349, 97.94888, 
    42.41491, 12.44253, 28.08678, 14.85801, 30.86785, 37.11079, 35.73439, 
    33.91776, 124.3871, 381.5867, 780.6381, 921.0138, 807.3401, 514.1893, 
    283.6758, 323.1736, 314.6895, 374.642, 395.0815, 392.9985, 310.7736, 
    226.0156, 184.2313, 147.4343, 164.883, 202.6225, 252.7558, 260.424, 
    307.9431, 309.5395, 311.4832, 401.2553, 517.3415, 550.1964, 679.3637, 
    525.896, 1.616105, 2.896513, 88.79086, 59.5556, 70.75466, 69.71838, 
    122.3319, 154.2911, 15.59744, 0, 0, 0, 0, 0, 27.71455, 6.569491, 0, 0,
  0, 439.4178, 195.6855, 907.5368, 1805.264, 1501.639, 712.643, 483.2295, 
    497.7593, 420.5321, 315.0768, 136.8431, 80.70911, 102.5947, 110.8975, 
    56.06786, 0.2648131, 3.387826, 36.63493, 22.48626, 4.213938, 32.13628, 
    34.12004, 9.394886, 55.34244, 71.22887, 124.1325, 164.2337, 141.1722, 
    73.3173, 29.08077, 2.917876, 50.12897, 16.72008, 8.767165, 20.09276, 
    6.12492, 9.995467, 2.303684, 0.02967453, 7.202766, 15.59999, 0, 4.923676, 
    28.76822, 14.64493, 19.81721, 22.2378, 29.72172, 55.51414, 46.22926, 
    135.3196, 311.9851, 389.0701, 426.3514, 394.7778, 346.0056, 381.4013, 
    311.8159, 286.077, 316.2218, 321.0644, 306.4557, 227.0812, 163.6294, 
    111.7403, 127.4932, 171.2171, 128.8476, 186.4454, 234.3389, 277.8444, 
    263.8623, 387.7439, 507.9923, 593.5289, 671.5868, 151.9244, 0, 0, 
    0.1526855, 11.12141, 27.27045, 5.642293, 0, 0, 0, 0, 0, 0, 0, 0, 
    29.69389, 0, 0, 0,
  336.1212, 283.2744, 280.2505, 1349.746, 1791.143, 1240.253, 581.5303, 
    454.5894, 529.9597, 451.9621, 271.3024, 88.98106, 65.69213, 79.26176, 
    83.76402, 15.86282, 0, 0, 0, 0.01159282, 3.559813, 3.361201, 26.5549, 
    78.995, 104.8708, 111.296, 123.7502, 183.7094, 170.4765, 96.75568, 
    18.82452, 36.92904, 173.0009, 147.0736, 0.6561724, 40.09827, 1.400087, 
    18.67419, 0, 4.921213, 17.68606, 0.02064603, 0, 0.5728964, 18.75198, 
    13.3812, 8.656983, 8.488718, 38.44683, 61.09453, 51.83106, 52.62397, 
    58.6014, 59.39347, 165.6035, 290.221, 454.3603, 531.7468, 356.0366, 
    250.5548, 230.6507, 267.4886, 263.0035, 170.9993, 101.3395, 226.0812, 
    405.6003, 438.8228, 243.4076, 140.5213, 194.1314, 222.0123, 325.5292, 
    476.0626, 621.8958, 708.6229, 614.3857, 5.007009, 0, 0, 0.5131387, 
    10.68596, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.96639, 0, 0, 0,
  1014.961, 1059.676, 999.4585, 1486.217, 1353.48, 822.1008, 483.4728, 
    423.429, 432.9811, 400.1913, 184.7545, 59.76541, 51.08024, 32.45238, 
    3.397727, 1.339373, 0.5192116, 1.949396, 6.878533, 0.8359628, 0, 
    0.4469217, 32.46057, 94.17204, 138.7826, 139.0123, 142.075, 170.2651, 
    199.8437, 156.3874, 66.95568, 99.59976, 214.9215, 163.2938, 0, 
    0.00557197, 0, 0, 0, 37.75103, 85.04147, 0, 0, 0, 2.593199, 6.704577, 
    0.9132928, 2.0938, 109.5198, 89.66087, 71.78169, 61.52934, 55.7276, 
    50.0367, 66.96713, 204.8958, 385.6734, 415.6871, 273.868, 163.4537, 
    185.3572, 235.6016, 183.325, 121.5506, 331.4378, 656.7086, 973.7778, 
    936.9366, 698.6102, 315.4651, 158.0312, 304.8352, 599.1711, 767.9793, 
    739.1931, 587.2299, 272.567, 0, 0, 0.0005063568, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.3449626, 0.8638448, 0, 0, 0,
  1276.519, 1596.647, 1710.525, 1532.737, 942.0485, 525.4172, 468.8974, 
    340.8898, 335.7376, 367.5742, 202.7082, 87.97628, 47.15509, 23.6611, 
    2.109894, 16.11546, 63.89506, 99.67946, 35.14595, 6.804534, 11.33926, 
    3.489694, 4.426375, 51.48684, 116.296, 132.7959, 119.1194, 141.0041, 
    206.496, 213.7981, 189.8233, 189.694, 225.2005, 137.5171, 0, 0, 0, 0, 0, 
    51.36637, 209.3645, 35.64569, 0, 0, 0, 0.1678525, 0, 0, 2.154153, 
    17.08876, 89.85088, 131.7713, 127.0772, 66.14963, 54.64122, 98.0938, 
    154.5197, 216.6144, 122.0288, 144.2869, 194.6717, 195.0684, 113.4059, 
    305.1859, 773.1769, 944.6837, 944.9396, 1041.262, 1010.897, 714.8572, 
    441.2517, 615.52, 994.8956, 1017.131, 735.3895, 398.553, 39.48136, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.48005, 0, 0, 0, 0,
  576.1854, 931.6247, 906.6362, 782.9591, 492.1016, 465.3861, 284.8566, 
    247.166, 278.3712, 328.5902, 197.9191, 70.77742, 37.59184, 12.53315, 
    7.181137, 43.26176, 121.2297, 201.0618, 133.2232, 65.32127, 50.51119, 
    18.33489, 0, 0.11232, 20.32129, 27.82987, 23.76683, 29.30825, 141.2721, 
    243.3896, 253.101, 230.2507, 183.3705, 51.35647, 0, 0, 0, 0, 0, 0, 
    70.44017, 221.9524, 66.5798, 0, 0, 0, 0, 0, 0.3017679, 8.757327, 
    127.2703, 222.3685, 176.8489, 129.8425, 56.31729, 30.53881, 53.13721, 
    56.63842, 85.90793, 110.0528, 170.028, 155.7422, 181.1576, 658.582, 
    891.925, 765.0097, 566.7166, 683.1484, 938.3599, 946.0663, 950.6962, 
    1152.784, 1400.864, 1190.112, 699.8245, 303.8513, 1.38781, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.373055, 0.3063857, 0, 0, 0, 0,
  645.5978, 651.4741, 348.0461, 338.1821, 333.729, 297.324, 274.5483, 
    329.6071, 320.4292, 242.4523, 142.7768, 33.2918, 19.17206, 13.50416, 
    14.204, 8.873847, 37.03663, 147.5774, 138.1909, 116.1385, 174.9569, 
    163.6211, 73.71962, 29.18241, 51.88186, 92.01063, 38.92251, 26.84706, 
    114.0117, 203.6541, 270.5715, 215.7726, 151.7382, 14.68677, 0, 0, 0, 0, 
    0, 0, 0, 40.54074, 369.3293, 317.3165, 114.3371, 3.862887, 0, 0, 0.11153, 
    0.006048144, 19.55387, 142.5781, 154.5665, 123.9076, 179.1985, 79.16, 
    14.5393, 34.07465, 42.74265, 97.64807, 169.0159, 219.1613, 396.9012, 
    642.2534, 732.5916, 397.1309, 377.0508, 643.4995, 985.1297, 1109.908, 
    1146.201, 1363.316, 1434.265, 1369.427, 928.765, 436.3409, 111.6556, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.772016, 0.006933623, 0, 0, 0, 0, 0,
  832.0802, 796.4195, 452.5931, 305.7719, 293.3802, 263.662, 251.0075, 
    350.6158, 214.3606, 118.4772, 23.99523, 9.823727, 0.9374197, 9.133391, 
    30.28316, 31.31364, 7.673902, 30.12636, 73.6406, 163.2412, 282.5515, 
    383.3724, 343.9316, 270.9898, 269.3295, 315.7319, 274.4701, 208.2753, 
    218.7913, 263.5744, 306.8953, 271.2532, 182.3894, 67.36945, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.676641, 71.09753, 100.5261, 93.03223, 0, 0, 0, 0.029983, 
    0.2834589, 5.7791, 29.0103, 202.0174, 299.2979, 245.8783, 10.45641, 
    3.441845, 9.227307, 65.13091, 143.5608, 212.5292, 258.0329, 406.613, 
    314.3367, 276.2676, 445.5888, 781.3271, 1096.255, 1218.235, 1079.923, 
    998.8617, 1214.761, 1232.076, 1011.277, 597.6057, 136.1366, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.308824, 17.42456, 0, 0, 0, 0, 0, 0,
  522.8505, 646.8199, 434.2559, 254.1983, 198.1381, 141.3106, 157.4017, 
    202.436, 98.83956, 4.720938, 5.80146, 1.222248, 0.002537446, 0, 6.751021, 
    16.09051, 4.110047, 0, 67.87675, 217.9813, 406.6455, 577.1392, 615.5616, 
    464.1506, 415.4912, 491.5859, 515.1653, 499.5445, 526.2872, 472.2782, 
    484.1233, 346.7195, 209.6823, 28.12877, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.04541712, 0.1208085, 35.22072, 93.14128, 169.8435, 
    92.35309, 0, 0, 0.01013316, 4.865694, 16.84927, 23.22182, 27.02969, 
    119.0616, 246.3213, 518.4421, 657.4585, 736.8021, 1052.213, 1052.852, 
    1112.684, 1157.132, 1119.51, 1128.288, 975.9925, 711.0227, 271.4639, 
    11.86194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20065, 51.1852, 0, 0, 0, 0, 0, 0, 0,
  189.5987, 372.6584, 272.8972, 153.0684, 129.0797, 107.2802, 101.2548, 
    98.52764, 13.1368, 0.6186931, -0.0932398, 0.01887309, 0, 0, 0, 0, 
    5.934471, 249.3546, 496.3241, 641.0406, 712.6684, 883.3423, 769.7581, 
    568.9565, 546.6921, 654.5696, 742.6288, 773.7735, 770.8872, 664.8349, 
    517.9086, 240.3035, 48.13427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 25.80465, 75.88532, 127.7064, 5.597481, 0.01321575, 0.01744381, 
    0, 0, 0, 0.008600875, 0.2463465, 0, 3.196367, 26.82889, 218.4336, 
    438.3653, 500.2625, 445.5697, 536.2654, 907.6587, 1133.265, 1245.885, 
    1148.132, 918.5613, 905.1179, 873.1757, 565.6349, 139.6936, 9.307497, 0, 
    0, 0, 0, 0, 0, 0, 5.973339, 51.01183, 18.53154, 0, 0, 0, 0, 0, 0, 0,
  66.53913, 126.0707, 158.3924, 101.3495, 129.9872, 153.1423, 111.0585, 
    69.88337, 5.909921, 0, 0, 0, 0, 0, 0, 0, 6.110831, 443.8941, 822.0618, 
    1065.257, 1147.54, 1026.579, 615.9289, 217.0476, 161.5421, 240.8548, 
    308.3307, 226.1226, 224.5132, 167.3122, 91.86687, 2.702835, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.687579, 0, 0, 0, 0, 2.009178, 150.2296, 
    137.6718, 53.3191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01111945, 8.059679, 
    76.88058, 223.2468, 192.0626, 54.48991, 351.7439, 523.5924, 854.4131, 
    841.848, 774.7855, 709.6036, 701.8489, 900.449, 776.0449, 283.2952, 
    20.40456, 0, 0, 3.21502, 41.93052, 145.8842, 257.1946, 238.5102, 
    233.1759, 92.08567, 0, 0, 0, 0, 0, 0, 0, 0,
  10.54719, 38.52236, 89.41316, 88.45621, 129.8748, 140.0378, 1.758609, 
    3.622372, 20.79722, 16.84281, 3.764497, 0, 0, 0, 0, 0, 0, 9.974582, 
    203.0671, 552.9215, 723.358, 628.1764, 114.8102, 1.827135, 0, 0, 
    0.02597354, 4.145141, 11.91014, 1.813728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.070437, 19.12915, 65.26246, 40.89855, 0, 1.946335, 0.4316256, 
    4.962647, 138.3129, 0, 0, 0, 0, 0, 0, 0, 0, 0.7391827, 0.9985219, 
    0.398542, 4.360011, 16.71775, 12.17988, 71.93053, 79.30731, 98.12679, 
    133.4162, 234.3277, 244.6326, 294.9109, 406.4966, 458.4559, 607.9581, 
    806.5295, 651.6235, 97.59635, 26.42796, 0, 11.91634, 142.9294, 523.1003, 
    623.8453, 728.3721, 414.541, 179.0205, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.2375568, 35.22453, 45.78533, 100.8335, 98.73385, 0, 19.24257, 
    69.95895, 49.19936, 14.10529, 0.5963095, 0, 0, 0, 0, 0, 0, 0, 14.52876, 
    100.917, 29.60974, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.002305, 0, 0, 
    0.049075, 0, 0, 0, 0, 10.97873, 31.62269, 20.17602, 8.189528, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24.33025, 35.88162, 3.392136, 8.202249, 
    9.667623, 4.784458, 29.97687, 95.48793, 70.86581, 107.1511, 47.01993, 
    186.0479, 250.5408, 327.3635, 495.9941, 663.1337, 707.337, 343.3452, 0, 
    0, 12.89661, 177.2778, 526.8167, 650.3031, 730.8545, 475.256, 140.5307, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.1563355, 32.96153, 93.6973, 8.055909, 7.271522, 46.84789, 107.1797, 
    96.87433, 65.0823, 5.47474, 1.638984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46.7029, 45.70561, 2.701415, 
    1.950268, 1.063997, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.490511, 10.38847, 0.8451264, 0, 0.1427283, 5.747555, 26.19526, 
    79.84738, 54.79946, 32.89713, 97.37908, 252.4611, 375.3538, 398.1776, 
    596.9442, 749.3185, 517.8513, 3.130794, 0, 0, 92.81933, 348.3482, 
    500.1969, 715.4668, 515.3165, 78.95136, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 23.82193, 117.2348, 1.692671, 2.966081, 75.61375, 119.2401, 
    156.9432, 150.2247, 187.7098, 168.4926, 20.22646, 0, 0, 0, 0, 
    0.008525716, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112.4393, 
    187.7537, 277.7043, 196.2434, 63.29765, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.6239529, 13.39494, 0, 0, 0, 1.266546, 41.70436, 
    25.22967, 28.20456, 109.732, 279.7055, 394.6047, 507.9118, 776.3243, 
    775.1523, 364.5099, 50.67634, 5.433064, 185.3506, 421.2495, 414.1049, 
    393.2517, 297.5771, 294.7875, 7.586363, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 2.931184, 22.6025, 0, 26.93795, 109.4093, 139.878, 177.1416, 
    88.31774, 86.30247, 174.0245, 163.1162, 240.8645, 75.69065, 3.21588, 
    0.5801046, 6.936382, 0.1045908, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.200257, 139.026, 418.142, 149.2554, 1.2402, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.164914, 0.7948571, 0, 0, 0, 
    0.001168255, 16.67364, 19.89136, 43.50631, 130.2915, 266.5667, 415.8081, 
    554.9022, 713.0673, 638.9822, 273.1252, 216.0703, 123.0732, 400.6276, 
    240.1565, 113.1827, 94.77327, 41.31813, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 12.43825, 0.1656403, 16.24762, 3.12718, 2.06611, 
    13.84467, 122.0781, 227.2487, 363.1719, 217.4649, 58.97001, 0.598401, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.693333, 86.21237, 
    0.054159, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.497975e-05, 0, 0, 0, 0, 0, 4.237197, 6.721555, 63.53002, 114.1027, 
    265.6567, 554.0557, 724.3539, 712.1773, 539.7785, 160.6944, 68.24227, 
    103.9293, 73.31152, 28.09826, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0.03340246, 0, 4.537661, 95.45872, 73.8838, 90.62366, 
    59.25259, 54.20035, 152.8858, 94.76863, 8.248804, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1057689, 19.82886, 
    233.0814, 269.9969, 373.4673, 617.0306, 770.7498, 660.8774, 426.0227, 
    199.58, 211.4468, 198.4001, 14.72842, 0, 0, 0, 0, 15.84741, 3.091941, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 68.96684, 105.0802, 102.1657, 102.4648, 46.12123, 
    0.1862036, 4.137225, 14.37615, 0, 0, 0, 5.570907, 19.88484, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1777319, 
    320.2881, 508.4323, 575.6027, 669.407, 672.3879, 490.291, 289.8031, 
    238.265, 313.8378, 200.7386, 9.265935, 0, 0, 0, 0, 0.1091187, 4.402359, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1957944, 113.7033, 75.3949, 52.71202, 37.44812, 
    0.2004635, 0, 0, 0.123569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13.78675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.807943, 138.4678, 
    425.4565, 693.1362, 582.7962, 419.3349, 270.5754, 275.724, 489.4667, 
    545.7513, 206.3423, 1.7709, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 20.8598, 0.006193054, 2.341495, 0.4137827, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4644903, 19.146, 0.3230906, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76.46013, 93.74072, 366.0079, 
    496.2035, 424.2791, 175.4117, 154.8367, 347.1221, 670.9517, 666.6006, 
    261.9197, 13.65668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.259748, 
    120.2423, 2.125335, 0, 0, 0, 0, 0, 0, 0, 0, 0.5916959, 0, 2.078349, 
    11.29419, 52.72276, 269.5899, 324.7525, 54.04507, 40.68792, 0.01734185, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27.23831, 326.5949, 448.5767, 470.8265, 265.0998, 97.36693, 175.0721, 
    356.4594, 464.9758, 296.394, 24.18855, 0, 0, 0, 0, 0, 0, 0, 0, 6.498864, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 434.9876, 
    549.625, 194.8289, 0, 0, 0, 0, 0, 0, 0, 49.79148, 229.9053, 270.3666, 
    218.3152, 435.0714, 763.8671, 711.7297, 577.2573, 432.7135, 282.8728, 
    35.13057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 9.57939, 23.93509, 458.746, 758.4965, 540.113, 253.5558, 102.6653, 
    138.8913, 305.0443, 234.599, 15.73475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.66078, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.860931, 
    705.9603, 764.272, 264.1802, 0.009830754, 0, 0, 0, 26.49382, 30.51307, 
    107.7551, 497.813, 1169.735, 1488.845, 1487.634, 1470.97, 1528.288, 
    1292.458, 1079.739, 876.5819, 425.0653, 38.33871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.993676, 78.49228, 0, 
    302.9012, 626.1432, 557.4089, 253.4888, 65.42033, 56.02234, 195.751, 
    71.06109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04533782, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39.38756, 
    486.9271, 529.4836, 132.7024, 0, 0, 0, 188.4812, 192.5964, 498.543, 
    708.6475, 1124.227, 1743.003, 2079.127, 2174.609, 2030.333, 2037.837, 
    1968.742, 1794.981, 1306.613, 536.4325, 38.71229, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2987449, 0.9965169, 0, 
    24.91258, 299.2193, 349.5217, 135.9241, 25.71449, 1.858234, 83.3325, 
    37.25776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5446421, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008149051, 
    79.37028, 181.9968, 190.1527, 16.7675, 0, 13.55061, 980.6506, 768.5872, 
    1105.977, 1530.174, 1995.253, 2289.703, 2406.146, 2417.229, 2295.283, 
    2278.623, 2349.081, 2062.894, 1572.461, 794.2656, 199.4317, 65.12003, 
    90.86436, 1.968355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 58.45197, 215.2836, 156.8912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.912825, 3.799026, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10.55764, 11.55569, 0, 0, 140.3663, 1585.396, 1665.679, 1860.954, 
    2327.909, 2685.942, 2719.711, 2651.773, 2599.41, 2509.09, 2444.553, 
    2411.1, 2231.088, 1777.786, 1073.075, 389.2512, 394.257, 742.5377, 
    431.4628, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.323763, 161.9636, 163.3663, 42.97362, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2813061, 5.751188, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 162.3825, 1830.881, 2420.234, 2799.512, 2933.921, 3054.115, 
    3021.108, 2897.282, 2813.163, 2631.317, 2454.22, 2377.28, 2253.893, 
    1763.675, 967.3515, 294.468, 567.5514, 896.8688, 723.8139, 165.1352, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22.55821, 
    205.1908, 176.4454, 100.5338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.576109, 1.351869, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 224.3244, 1715.302, 2661.883, 3042.112, 3078.042, 3083.966, 
    3056.699, 2966.114, 2775.983, 2461.252, 2203.078, 2069.804, 2055.312, 
    1617.411, 858.8635, 63.53865, 565.2546, 820.6309, 464.1451, 208.9816, 
    21.89472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.308722, 
    41.45142, 0, 0, 39.56498, 1.861557, 0.9454954, 8.430882, 0, 0, 0.2580895, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 15.21186, 1.925179, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 69.28409, 1442.782, 2432.051, 3022.305, 3064.017, 2982.046, 2920.952, 
    2867.871, 2768.787, 2520.354, 2211.113, 1641.312, 1364.499, 1291.194, 
    1387.434, 845.2209, 244.3112, 296.0118, 614.2589, 358.0775, 523.442, 
    111.5307, 0.1241507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.110101, 52.63713, 243.9889, 184.6683, 0.4007951, 7.643325, 46.26271, 
    0.01746987, 11.53573, 9.214417, 0, 0, 2.880076, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 20.27884, 0.2822629, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 388.4866, 1897.231, 2823.74, 3016.014, 2869.568, 2752.483, 2647.189, 
    2529.865, 2443.268, 2159.798, 1604.969, 955.6561, 423.3286, 422.3328, 
    778.8141, 553.3457, 156.9905, 464.2124, 635.9963, 351.1034, 437.6381, 
    20.91868, 26.49133, 1.27366, 1.299142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.944896, 32.97338, 270.1112, 460.1797, 328.6203, 29.76436, 98.42758, 
    162.2669, 21.47914, 0.01439463, 0.09217066, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01224168, 16.85926, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 220.2471, 1591.738, 2466.678, 2747.279, 2660.819, 2426.795, 2163.563, 
    1904.25, 1726.834, 1309.499, 717.4695, 72.1908, 0.01969476, 0, 139.6303, 
    56.38565, 0.01733694, 280.8316, 373.5753, 88.71832, 60.37281, 22.64031, 
    35.58979, 1.627476, 11.44019, 3.820878, 2.149208, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01889744, 6.854713, 95.4062, 415.7192, 609.9531, 237.4828, 87.95111, 
    174.6365, 179.5905, 1.821839, 0.4608677, 1.038414, 1.955436, 0, 0, 0, 0, 
    0.4032466, 0, 0, 0, 0, 0, 23.75265, 6.992056, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 344.95, 1579.479, 2305.747, 2500.39, 2205.512, 1810.193, 1200.209, 
    851.3199, 495.871, 307.6716, 18.7188, 0, 0, 0, 0, 0, 0.007190464, 
    328.6132, 334.6894, 151.1666, 47.72522, 19.96992, 2.669097, 2.000999, 
    5.087904, 39.56742, 29.48166, 1.290598, 0, 0, 0, 0, 0, 0, 0, 0, 7.210662, 
    34.74933, 341.6028, 763.1323, 677.7067, 334.8472, 120.0849, 233.7542, 
    94.9697, 21.47264, 47.76735, 13.35156, 8.629306, 32.41949, 2.232151, 0, 
    0, 0, 1.06906, 0, 0, 0, 0, 12.63473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    220.6236, 1349.775, 2132.709, 2395.235, 2048.53, 1480.806, 855.7775, 
    314.9611, 477.5641, 130.0667, 3.648897, 0, 0, 0, 0, 0, 0, 10.08162, 
    642.4855, 281.7012, 101.1102, 60.59174, 61.11189, 54.33709, 36.61767, 
    64.51082, 191.8937, 50.27359, 0.1158935, 0.7644691, 0, 0, 0, 0, 0, 0, 0, 
    127.1192, 404.733, 737.6123, 874.3842, 641.8504, 235.5844, 192.8914, 
    214.4153, 206.9348, 198.1494, 125.9625, 26.56938, 2.941694, 5.601278, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.25005, 1.223589, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    123.0767, 1440.606, 2345.219, 2595.379, 2201.878, 1579.878, 765.6243, 
    263.2791, 17.18813, 95.84882, 0, 0, 0, 0, 0, 0, 0, 18.90151, 14.24182, 
    240.224, 244.171, 170.7711, 72.88946, 36.88171, 3.688538, 30.90802, 
    42.64079, 82.76118, 41.20324, 110.692, 64.07503, 0, 0, 0, 0, 0, 0, 
    116.6442, 851.2905, 1040.522, 1011.616, 761.973, 391.5457, 285.8691, 
    222.6031, 231.2289, 132.9321, 127.5657, 79.20253, 79.93398, 60.85431, 
    7.069205, 0, 0, 0, 0, 0, 0, 0.002840273, 31.90177, 12.23519, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    113.4006, 1133.138, 2195.308, 2608.468, 2239.793, 1572.94, 1003.211, 
    518.9925, 189.4889, 0.6126093, 0, 0, 0, 0, 0, 0, 0.1651795, 133.9569, 
    417.8274, 384.9297, 215.625, 141.7358, 90.05803, 79.19399, 29.33371, 
    2.240706, 12.30619, 0.2534847, 0, 94.7438, 162.481, 149.9046, 37.89026, 
    0, 0, 0, 0, 5.356696, 552.9598, 964.9863, 891.923, 640.1644, 439.5914, 
    361.2435, 278.5941, 283.0451, 244.8269, 280.0539, 219.772, 241.4119, 
    332.4167, 319.8716, 147.7597, 7.835948, 0, 0, 0, 0, 0.3774112, 84.49905, 
    37.25802, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30.39107, 
    914.6385, 1832.73, 2461.096, 2238.884, 1490.557, 718.7988, 432.395, 
    372.0842, 0.9015442, 0, 0, 0, 0, 0, 105.8306, 357.3896, 523.8076, 
    521.7178, 440.9008, 328.9724, 202.1082, 166.6164, 82.55063, 126.2423, 
    70.6189, 12.28226, 42.67114, 60.72597, 91.16128, 142.8304, 148.7395, 
    152.2123, 97.86357, 0, 0.3341298, 0.6432131, 4.719822, 37.05452, 468.78, 
    599.9188, 399.7013, 211.5083, 353.3973, 316.7687, 280.8083, 341.3538, 
    511.3751, 442.6859, 504.624, 253.1497, 250.1017, 213.2764, 67.04365, 
    3.304585, 0, 0, 0.1683532, 53.87643, 48.47186, 10.75609, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89.8662, 
    469.3024, 1154.713, 1449.781, 1272.478, 681.3491, 128.84, 4.544834, 0, 0, 
    0, 0, 0, 5.419511, 61.07015, 489.1122, 578.3217, 527.3911, 395.0327, 
    218.0269, 167.6713, 137.974, 115.5373, 0.6435879, 88.33016, 45.21404, 
    6.509036, 44.30594, 115.2863, 242.208, 245.5465, 151.2771, 0.4254271, 
    11.1162, 1.786039, 48.14689, 37.55202, 70.14665, 156.7791, 498.9786, 
    523.2408, 473.1295, 354.968, 545.134, 489.5596, 703.8699, 925.6036, 
    986.3214, 886.7418, 869.757, 604.8533, 197.4831, 113.1076, 12.6825, 0, 
    0.02486209, 6.962315, 96.1065, 54.04581, 0.01545697, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1216824, 0.9288862, 134.0087, 201.5549, 60.90172, 0.3555474, 0, 0, 0, 
    0, 0, 355.5598, 602.0829, 651.0312, 450.9958, 386.381, 256.653, 158.6886, 
    43.34907, 61.85168, 159.5036, 113.3953, 25.31179, 87.31884, 165.2257, 
    4.966446, 0.1061549, 45.43877, 108.6841, 188.0823, 174.495, 113.4314, 
    0.01686891, 145.4191, 132.487, 172.8789, 193.6581, 150.9564, 166.1918, 
    400.6677, 583.3967, 722.2389, 745.6167, 800.6808, 849.4872, 1009.411, 
    1053.753, 947.8483, 415.5219, 584.1187, 491.2827, 259.1023, 215.041, 
    112.3413, 76.86075, 134.8813, 221.4578, 45.61331, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.875198, 477.9095, 533.1882, 461.8639, 235.7978, 
    111.7738, 22.34331, 6.797899, 1.574463, 51.39446, 134.1712, 4.203103, 
    6.980784, 108.1984, 118.4102, 3.881124, 11.86376, 72.39351, 102.465, 
    159.5778, 156.6727, 107.9339, 109.4576, 488.6499, 418.6319, 300.2693, 
    237.9754, 185.1014, 104.7926, 403.3925, 659.502, 1010.157, 881.0416, 
    936.1367, 774.4136, 1186.745, 1002.815, 1015.139, 535.5046, 386.2178, 
    179.3871, 69.36623, 267.0681, 111.3501, 67.82533, 6.994944, 1.526611, 
    3.172025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.725166, 102.8057, 111.4602, 125.5778, 65.69091, 
    11.31183, 6.297175, 5.844241, 2.358717, 171.9062, 167.7866, 43.11033, 
    79.99084, 74.58493, 27.5016, 14.16823, 6.523846, 31.63298, 63.06898, 
    67.15324, 85.22324, 67.61577, 224.0022, 476.0859, 396.943, 309.3507, 
    246.142, 132.8316, 335.7784, 784.7097, 1053.235, 1127.867, 967.6097, 
    771.317, 924.9985, 1333.487, 1034.066, 789.8601, 234.963, 249.6979, 
    81.2932, 14.26598, 163.186, 164.9658, 5.164979, 1.026154, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.19746, 170.4447, 463.7712, 416.7452, 239.2617, 
    79.01589, 6.674962, 0, 0, 49.56345, 226.9828, 192.8199, 164.6065, 
    182.8128, 118.2701, 17.30331, 8.986745, 3.3333, 23.55511, 61.35153, 
    53.04255, 132.2586, 229.133, 315.2996, 329.1717, 262.2387, 250.0072, 
    217.4491, 311.0166, 854.7855, 1325.855, 1237.892, 1063.641, 815.3153, 
    855.515, 1043.939, 1759.73, 1143.116, 371.2457, 14.33288, 2.286062, 0, 0, 
    0.1220521, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 13.13908, 199.9922, 369.35, 332.041, 183.8263, 
    84.41653, 28.31347, 5.11356, 0, 3.346521, 94.1303, 145.3444, 260.3771, 
    308.1046, 216.5467, 65.93798, 66.89045, 91.82342, 129.8517, 169.2161, 
    212.0327, 380.3462, 430.9281, 398.8634, 271.8267, 213.1764, 198.3177, 
    260.7658, 507.0705, 1261.594, 1556.329, 1201.677, 977.4053, 903.3651, 
    1023.128, 1437.7, 2083.172, 1221.35, 86.26831, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.492808, 28.12763, 241.1122, 312.6933, 227.4316, 
    40.73929, 3.901017, 60.77868, 29.63254, 0, 37.46666, 47.92201, 90.67201, 
    252.6916, 297.8447, 250.6762, 146.2321, 137.6703, 164.451, 210.1363, 
    267.7924, 336.6427, 471.1196, 486.8597, 425.3645, 315.1228, 279.0462, 
    273.7747, 290.0505, 636.9206, 1410.759, 1544.152, 1250.766, 1127.925, 
    1065.812, 1110.734, 1416.591, 1600.496, 408.8422, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 8.41072, 11.77269, 0, 0, 1.62508, 8.022939, 6.219764, 0, 
    20.28673, 0.6057806, 40.99087, 150.5031, 84.34249, 84.26646, 195.8636, 
    227.4629, 190.5297, 136.6387, 154.2375, 176.6017, 216.4878, 304.6136, 
    374.8836, 462.7287, 472.5354, 402.6108, 307.9417, 327.0253, 306.5867, 
    373.0538, 668.3615, 1415.796, 1557.029, 1306.125, 1279.073, 1162.341, 
    1153.206, 1149.406, 1078.977, 41.16324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.901734, 217.5294, 284.0266, 9.755486, 12.21576, 30.38478, 
    126.8581, 295.4576, 261.4576, 148.2994, 19.41799, 0.001383794, 4.122153, 
    25.35506, 13.69719, 14.41783, 64.17224, 71.70509, 82.17438, 88.62575, 
    143.002, 168.497, 227.1901, 295.2106, 377.9786, 424.9349, 434.2556, 
    359.2029, 243.9208, 256.3825, 320.5891, 276.9689, 544.5539, 1255.969, 
    1424.041, 1287.706, 1179.742, 1196.443, 1053.201, 1167.506, 829.4473, 
    18.81178, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3367717, 55.36858, 332.4312, 482.9248, 279.4982, 0, 4.759403, 138.2639, 
    246.2088, 336.8652, 256.5343, 116.4693, 7.490035, 1.586183, 5.608893, 
    0.125523, 0.02205558, 0, 18.84512, 43.35651, 73.8119, 134.7575, 190.767, 
    245.426, 262.851, 321.6095, 350.954, 368.8531, 361.5361, 275.9557, 
    193.2714, 264.4291, 287.2755, 295.1925, 454.3226, 894.5059, 1154.717, 
    973.0314, 1099.105, 1148.796, 1120.024, 862.0306, 375.9889, 12.88452, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2140546, 
    0.1701733, 26.3982, 16.54789, 11.51096, 64.69183, 320.2927, 487.4863, 
    486.2169, 178.1183, 52.80968, 111.4205, 188.5571, 226.6747, 194.1454, 
    121.9309, 19.68636, 0, 0, 0, 0, 0, 0, 0.08443239, 12.21449, 77.40128, 
    139.2317, 232.2935, 274.8673, 306.887, 328.7855, 366.2649, 352.3075, 
    297.598, 212.2141, 162.9654, 161.8156, 294.4319, 331.9783, 424.2078, 
    668.4012, 775.5222, 991.9241, 1072.528, 1282.538, 1139.612, 931.2537, 
    216.4193, 62.45685, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.731169, 
    99.69241, 145.8221, 164.5461, 190.2277, 222.6298, 352.1655, 453.9755, 
    483.7257, 366.7473, 201.0961, 195.8921, 224.278, 247.8174, 199.336, 
    145.5127, 58.51702, 0.01620398, 1.724691, 0, 0, 0, 0, 0, 0, 3.441099, 
    66.59528, 167.6643, 266.4513, 312.1495, 332.5176, 373.2896, 422.7214, 
    417.7817, 331.4211, 227.7531, 191.2091, 276.8271, 346.7453, 491.9813, 
    515.8571, 477.7105, 837.2191, 1215.665, 1373.787, 1364.735, 1284.096, 
    957.2903, 218.0976, 83.97918, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.299129, 134.0267, 
    294.2319, 344.9782, 270.6827, 318.7709, 384.5544, 494.1917, 494.657, 
    473.3284, 365.3275, 308.8357, 293.0063, 310.0292, 272.0663, 223.5598, 
    135.7657, 49.15474, 0.05388123, 0.2981069, 0, 0, 0, 0, 0, 0, 0.2216611, 
    69.87698, 190.6432, 286.7062, 330.1897, 367.8758, 406.1044, 450.1877, 
    427.9415, 330.3656, 250.8139, 289.5048, 447.8335, 462.0058, 478.6495, 
    494.2013, 530.5643, 958.8607, 1535.851, 1566.941, 1493.999, 1267.836, 
    1004.899, 187.0762, 37.84942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2778322, 1.216981, 0.320554, 
    82.15788, 124.0773, 328.814, 414.2038, 370.9027, 408.5572, 474.0244, 
    515.583, 504.9358, 517.7888, 478.3085, 405.8519, 390.0446, 340.6481, 
    284.1749, 193.1102, 63.77376, 0.2711483, 0.001171568, 0, 0, 0, 0, 0, 0, 
    0, 0.01659026, 97.79198, 225.3099, 301.7682, 358.1664, 393.5924, 
    409.4816, 387.7672, 372.0033, 279.7969, 234.8109, 369.993, 486.2102, 
    487.3097, 453.6224, 565.4487, 638.8194, 1025.565, 1495.267, 1465.116, 
    1353.271, 1132.2, 829.127, 232.6918, 86.18745, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03872748, 20.11839, 53.78059, 
    33.44499, 88.68514, 177.8256, 19.69762, 253.2851, 404.7767, 437.9373, 
    469.3643, 499.6412, 501.7674, 551.6224, 574.769, 536.6869, 488.521, 
    416.7465, 350.7989, 264.6436, 127.1555, 0.415809, 0.4254224, 0, 0, 0, 0, 
    0, 0, 0, 0.6914847, 19.04652, 131.946, 247.1787, 306.9858, 363.0714, 
    397.9942, 400.0674, 409.7594, 398.0919, 355.8009, 291.4016, 333.1392, 
    498.2859, 440.002, 539.7181, 723.6176, 765.5291, 965.6453, 1312.768, 
    1339.947, 1188.61, 996.9376, 753.3426, 184.1582, 17.82256, 30.13374, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.789168, 70.13921, 107.3934, 180.0283, 
    234.5805, 241.1893, 107.9595, 15.09211, 188.5137, 368.2224, 514.8614, 
    566.2856, 554.1669, 566.897, 608.2187, 604.4344, 543.1758, 479.5136, 
    420.2968, 358.7137, 272.7408, 113.1928, 4.518106, 5.010964, 0, 0, 0, 0, 
    0, 0, 0.7098004, 13.29282, 97.01318, 193.7101, 286.6924, 317.051, 
    366.6038, 397.0652, 432.3381, 481.5545, 519.4891, 467.0329, 436.6177, 
    526.4904, 556.9227, 596.2275, 609.3391, 692.4142, 720.394, 862.9467, 
    1120.028, 1117.907, 1092.196, 985.4866, 917.553, 349.6905, 24.9056, 
    102.5677, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.45255, 45.57545, 90.12004, 208.861, 
    326.2532, 247.4885, 3.031927, 0.8162752, 62.72859, 240.1284, 478.4014, 
    642.7585, 624.4623, 612.9011, 633.5761, 635.511, 540.0829, 464.6622, 
    389.1842, 327.2373, 250.5822, 128.0566, 4.151914, 0.01724564, 0, 0, 0, 
    0.06221788, 16.14303, 56.51927, 60.10637, 63.71621, 129.8515, 214.7995, 
    265.7689, 302.5134, 336.1973, 365.2288, 442.3849, 504.6011, 502.0141, 
    480.3363, 467.8888, 553.1976, 593.0986, 637.1354, 629.6438, 659.4634, 
    735.4026, 1028.44, 1056.044, 946.681, 926.314, 1064.744, 949.1011, 
    392.1784, 18.68724, 70.3578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.13205, 81.59405, 283.5952, 
    99.12554, 0, 2.600603, 22.27865, 40.11892, 259.8885, 493.662, 624.6654, 
    578.1021, 631.7147, 627.2502, 560.2089, 436.4544, 359.2498, 263.4945, 
    198.2276, 96.85187, 8.224985, 0.006419148, 10.41262, 28.47488, 33.42284, 
    63.55798, 89.37606, 117.4287, 123.5775, 113.715, 153.6499, 198.5007, 
    238.3534, 277.4305, 321.2411, 352.9605, 414.103, 455.9593, 452.3423, 
    458.7655, 565.2747, 608.5494, 639.5411, 687.265, 764.0191, 736.5245, 
    987.5319, 1266.858, 1113.241, 848.986, 966.5779, 1123.773, 1059.529, 
    375.9788, 5.606318, 11.23915, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50.03308, 18.7767, 0, 
    1.26797, 38.3414, 37.16248, 6.458248, 236.8902, 463.1305, 562.8348, 
    578.8032, 630.9438, 520.6262, 426.2543, 325.3188, 244.9647, 138.4487, 
    36.07342, 0.5078325, 2.94648, 57.33051, 95.80891, 105.8, 111.6879, 
    121.1859, 142.7138, 152.8308, 160.8624, 182.531, 201.2338, 222.661, 
    264.4805, 303.7233, 333.4624, 371.3336, 438.1491, 455.2211, 496.9004, 
    597.2755, 643.8214, 617.1034, 691.8447, 823.0101, 988.5286, 1358.407, 
    1648.078, 1373.022, 979.8769, 1118.349, 1293.235, 1281.518, 524.8214, 
    12.07863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.53168, 7.44618, 
    0.2774768, 0, 35.85915, 285.9109, 179.5872, 150.5524, 421.4404, 514.148, 
    569.3135, 533.7565, 453.5545, 348.8341, 297.6014, 196.2376, 72.14723, 
    1.141348, 3.445107, 14.83014, 68.87897, 118.991, 129.5745, 158.0152, 
    182.8073, 209.6761, 221.1556, 222.757, 222.7252, 225.1968, 215.3978, 
    252.5812, 274.6012, 313.8231, 378.8444, 483.5266, 526.6315, 559.9622, 
    581.9632, 617.732, 638.4788, 691.2427, 829.9338, 1126.817, 1687.072, 
    1798.549, 1466.908, 1100.552, 1091.336, 1508.885, 1401.512, 703.5411, 
    81.51077, 0.2449444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.97898, 137.8128, 2.629696, 
    0.1815157, 0, 28.15523, 299.744, 311.1771, 79.97313, 377.6644, 488.9033, 
    461.6871, 486.7418, 409.492, 350.8954, 279.0941, 180.3749, 25.7736, 
    3.397881, 18.72686, 43.95182, 103.1606, 144.6976, 190.1044, 222.457, 
    259.2217, 285.7209, 287.2361, 281.1645, 272.6286, 249.3425, 225.9028, 
    238.7993, 272.0008, 332.6962, 384.1511, 468.3911, 546.1947, 577.4488, 
    627.5869, 635.5259, 700.1279, 776.9152, 929.8552, 1510.917, 1895.887, 
    1799.537, 1355.943, 1119.573, 1392.253, 1618.039, 1311.142, 575.1276, 
    257.3511, 0.8315546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.894205, 72.59029, 14.85453, 
    7.508962, 13.51235, 142.9096, 296.0406, 327.9227, 156.2393, 437.1971, 
    388.5025, 385.3842, 401.033, 394.5582, 335.838, 280.1766, 193.5683, 
    96.386, 35.52516, 58.84515, 86.79417, 122.0659, 181.4595, 237.5804, 
    289.2039, 326.9966, 354.348, 356.1935, 336.6149, 307.5397, 253.4356, 
    225.7552, 236.1096, 334.7573, 444.7771, 494.1808, 514.2294, 524.8425, 
    587.1181, 631.0831, 694.0496, 751.4611, 825.4266, 1097.83, 1658.775, 
    2006.745, 1602.702, 1223.444, 1127.629, 1333.478, 1458.12, 871.0525, 
    466.6771, 267.9041, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01038057, 0, 6.643703, 101.4879, 
    82.98901, 51.23274, 85.14922, 210.2779, 283.6747, 309.324, 233.2301, 
    492.1425, 371.6667, 362.65, 444.5501, 397.6977, 330.4786, 280.92, 
    273.9966, 219.3448, 153.7401, 126.073, 117.5657, 150.8828, 219.6838, 
    283.4588, 333.4008, 374.8239, 400.1253, 395.6437, 375.5026, 312.2456, 
    243.2001, 227.2077, 279.3844, 409.5839, 514.515, 561.0614, 561.6627, 
    541.6973, 592.7158, 646.3815, 705.6855, 755.9585, 820.3306, 1077.465, 
    1725.695, 1795.541, 1577.446, 1249.411, 1148.976, 1319.127, 995.0981, 
    382.848, 349.3625, 65.2517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.50258, 104.9451, 82.473, 
    92.12851, 176.1149, 268.6027, 316.0862, 341.2645, 486.9077, 443.9214, 
    441.7123, 453.1961, 411.6028, 339.4975, 305.282, 294.3625, 287.3364, 
    230.1652, 207.584, 207.6316, 229.0633, 299.8941, 320.3898, 366.2971, 
    403.0446, 399.9144, 400.9593, 372.4525, 306.9135, 239.632, 240.6821, 
    343.6025, 474.4823, 553.2586, 592.0007, 575.3657, 602.5383, 624.6992, 
    700.6254, 727.1317, 764.283, 781.6901, 1065.684, 1631.907, 1692.728, 
    1571.499, 1298.507, 1313.886, 1286.554, 934.9397, 106.3758, 289.6695, 
    15.00103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.55675, 115.867, 
    22.48811, 65.3556, 149.1486, 286.7424, 407.3988, 236.5376, 274.9689, 
    357.7444, 443.3862, 421.6057, 401.2734, 343.1813, 298.683, 307.432, 
    300.7722, 291.2484, 308.8382, 334.8492, 323.8983, 337.6805, 341.7525, 
    399.8321, 429.9846, 410.5637, 382.6377, 354.2699, 306.8083, 234.6121, 
    282.1734, 378.2628, 513.45, 570.4268, 609.7987, 630.7244, 657.3438, 
    763.2346, 822.8828, 897.2252, 876.2137, 902.7307, 1085.887, 1506.075, 
    1453.561, 1306.629, 1103.886, 1026.492, 1225.022, 985.5616, 402.682, 
    411.0314, 92.16769, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.036347, 62.52849, 
    3.547037, 32.43497, 104.1824, 329.8143, 462.2404, 251.2797, 109.8259, 
    300.0777, 382.1133, 340.6129, 357.1865, 326.0741, 305.6071, 339.9389, 
    372.1312, 391.5172, 407.5522, 352.1345, 293.8417, 268.1846, 292.7089, 
    444.7627, 466.584, 417.2143, 374.3411, 349.6299, 313.55, 266.888, 
    336.9229, 432.6651, 484.9139, 546.2026, 630.8204, 650.4514, 755.9393, 
    824.0303, 861.4523, 911.7997, 958.1385, 976.4166, 1254.706, 1563.365, 
    1293.88, 1170.993, 864.0294, 700.7004, 757.6398, 917.2304, 682.3601, 
    402.354, 43.28111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05915249, 0.08011421, 0, 
    6.02283, 76.62966, 347.7174, 469.9626, 235.3439, 100.1177, 160.2919, 
    227.011, 263.368, 336.6925, 322.0186, 290.6877, 363.0302, 432.0052, 
    448.0348, 357.6713, 268.9411, 179.2584, 179, 233.9073, 359.2671, 
    464.7566, 411.7307, 372.834, 358.2526, 326.1168, 293.7316, 402.5888, 
    470.521, 497.5835, 578.8224, 635.5013, 674.5109, 734.5461, 763.5286, 
    810.0879, 885.3263, 939.2901, 1104.282, 1317.147, 1582.151, 1373.822, 
    1213.066, 873.9077, 635.079, 382.4486, 656.3605, 884.5526, 664.905, 
    217.4573, 32.62277, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.014362, 
    61.41228, 327.5756, 417.7493, 328.8751, 249.4016, 131.7789, 157.5266, 
    287.179, 367.0403, 311.7421, 237.5124, 263.4082, 315.4411, 318.5938, 
    269.0101, 179.5965, 192.4013, 228.7823, 193.9452, 278.2494, 363.2266, 
    430.6738, 408.0237, 404.8087, 350.7692, 302.6519, 419.8691, 508.0556, 
    530.116, 605.4689, 677.9661, 698.0052, 724.3315, 784.8451, 801.787, 
    928.4433, 1166.382, 1351.242, 1463.7, 1691.588, 1541.213, 1399.71, 
    1026.168, 717.6241, 512.4301, 377.8375, 697.6708, 594.645, 397.4904, 
    142.8448, 0.532489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2053152, 
    67.53915, 303.6299, 379.2345, 436.3914, 423.1708, 180.6438, 155.2336, 
    276.7622, 326.9408, 266.7624, 175.7495, 176.1388, 195.9187, 226.1668, 
    186.327, 215.0712, 291.8131, 416.8516, 394.0894, 300.8634, 340.7516, 
    360.322, 408.5583, 425.7607, 360.9985, 326.2549, 435.8652, 544.7354, 
    572.8199, 653.0318, 746.2729, 793.1929, 824.189, 828.2086, 914.1102, 
    1028.284, 1346.432, 1671.313, 1678.606, 1814.529, 1881.197, 1709.896, 
    1406.109, 1219.147, 1059.282, 948.7432, 834.345, 919.3475, 724.296, 
    356.6761, 76.5276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8787696, 13.35174, 
    137.5124, 287.6332, 345.7241, 417.4199, 379.3897, 131.3522, 106.2649, 
    169.0464, 272.2558, 288.1475, 201.0602, 176.5896, 223.6827, 266.1863, 
    218.2081, 176.9505, 269.0522, 436.2097, 486.094, 402.9827, 347.54, 
    334.3905, 365.894, 393.4282, 347.4721, 379.8949, 443.5723, 566.2279, 
    602.1741, 676.5858, 812.3363, 900.5889, 908.915, 931.9954, 944.5102, 
    1117.414, 1304.28, 1882.296, 1832.433, 1976.871, 2069.233, 2070.061, 
    1899.477, 1551.457, 1340.278, 1386.592, 1314.673, 1244.868, 1230.34, 
    806.1844, 287.225, 40.42369, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.817714, 35.69061, 
    138.5443, 281.9023, 361.2498, 453.4521, 359.1906, 222.1722, 156.6933, 
    136.975, 236.7071, 325.3279, 228.1469, 196.3775, 242.6227, 329.216, 
    249.9151, 180.1256, 229.7955, 351.343, 390.6742, 362.7199, 313.2054, 
    299.3227, 315.3665, 337.3273, 403.3815, 440.4469, 459.0341, 544.0665, 
    574.6163, 685.2004, 805.9506, 978.1014, 1079.502, 1060.385, 1335.979, 
    1386.026, 1736.179, 2369.993, 2377.097, 2108.683, 2192.729, 2248.685, 
    2160.981, 1428.064, 1097.215, 1308.715, 1435.482, 1437.344, 1562.363, 
    1290.539, 805.3401, 441.8997, 16.92101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
