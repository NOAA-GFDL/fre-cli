netcdf atmos_scalar.185001-185412.ch4global {
dimensions:
	time = UNLIMITED ; // (60 currently)
	nv = 2 ;
variables:
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	float ch4global(time) ;
		ch4global:long_name = "Global Mean Mole Fraction of CH4" ;
		ch4global:units = "1e-09" ;
		ch4global:missing_value = 1.e+20f ;
		ch4global:_FillValue = 1.e+20f ;
		ch4global:cell_methods = "time: mean" ;
		ch4global:time_avg_info = "average_T1,average_T2,average_DT" ;
		ch4global:standard_name = "mole_fraction_of_methane_in_air" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;

// global attributes:
		:filename = "atmos_scalar.185001-185412.ch4global.nc" ;
		:title = "ESM4_historical_D1" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 
    30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 
    396, 424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 
    820, 850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 
    1215, 1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 
    1580, 1611, 1641, 1672, 1703, 1733, 1764, 1794 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 
    424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 
    850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 1215, 
    1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 1580, 
    1611, 1641, 1672, 1703, 1733, 1764, 1794, 1825 ;

 ch4global = 785.6929, 785.4942, 785.5226, 785.7922, 786.0576, 786.2314, 
    786.1946, 786.1538, 786.2097, 786.2639, 786.2376, 786.0377, 785.7965, 
    785.6385, 785.6697, 785.9232, 786.2079, 786.3453, 786.3303, 786.3425, 
    786.4296, 786.4482, 786.4036, 786.2725, 786.0201, 785.8631, 785.9703, 
    786.3475, 786.7098, 786.9166, 787.0101, 787.1331, 787.2822, 787.4207, 
    787.3549, 787.2523, 787.0323, 786.9629, 787.1694, 787.539, 787.8179, 
    788.0863, 788.2224, 788.3068, 788.4232, 788.5469, 788.66, 788.5295, 
    788.2682, 788.2153, 788.4113, 788.8005, 789.1882, 789.4916, 789.6053, 
    789.6478, 789.7908, 789.9327, 789.9973, 789.9347 ;

 nv = 1, 2 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825 ;
}
