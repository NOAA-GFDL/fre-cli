netcdf \20030101.atmos_static_cmip.tile4 {
dimensions:
	grid_xt = 96 ;
	grid_yt = 96 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:associated_files = "area: 20030101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 time = 0 ;

 orog =
  0.05263353, 0.9425675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.210776, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.252779, 74.21071, 95.69428, 
    40.84037, 37.33909, 173.0547, 413.3694, 558.9451, 332.2694, 351.5737, 
    71.52609, 0.03417388, 1.300127, 17.79588, 8.458535, 18.73478, 17.63159, 
    0, 0, 0, 24.16101, 0, 0, 0, 0, 0, 0, 0, 1.372658, 299.2773, 291.463, 0, 
    0, 0, 0, 0, 0.0248737, 34.27986, 188.9342, 329.4237, 350.9251, 251.6835, 
    165.8015, 165.6417, 201.2802, 268.5535, 314.2737, 338.9506, 356.3144, 
    377.6248, 410.6694, 439.9049, 453.2951, 445.0014, 438.5307, 407.9247, 
    339.9653, 265.3149, 224.8092, 190.4008, 158.7892, 103.6094, 19.02374, 0, 
    0, 0,
  9.158454, 18.90683, 3.012916, 53.90588, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2984579, 4.255527, 
    84.79544, 147.7691, 233.7292, 347.7168, 36.84171, 0, 0, 0, 0, 0, 0, 
    0.4999831, 0, 0, 0, 25.2615, 9.891716, 381.2982, 0.7240577, 0, 0, 0, 0, 
    147.3826, 251.5665, 17.10577, 0, 0, 0, 0, 0, 12.48063, 173.854, 367.2847, 
    472.174, 458.6521, 325.3309, 227.1559, 236.9397, 249.4832, 296.6798, 
    348.9885, 370.6396, 368.1631, 393.7355, 411.4686, 451.679, 461.741, 
    457.9003, 439.6093, 391.6231, 291.6416, 227.3665, 205.8765, 180.0435, 
    108.2699, 20.55778, 0, 0, 0, 0,
  146.5898, 178.415, 28.03686, 31.16747, 0, 0, 0, 0, 0, 0, 0, 0, 0.03837012, 
    1.052421, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.03251622, 0.6342183, 0, 0.003365346, 0.1732605, 15.05509, 
    0.627657, 0, 0, 5.064898, 0.5615213, 22.54741, 2.144348, 0, 0, 255.0734, 
    8.867086, 0, 0, 0.008958309, 1.017161, 28.21741, 115.5201, 0, 0, 0, 0, 0, 
    0, 66.54465, 223.7023, 341.7935, 467.8122, 479.3343, 405.95, 344.1333, 
    317.8734, 316.412, 353.7882, 397.7623, 399.601, 410.1562, 420.6944, 
    456.795, 491.1674, 486.9185, 461.8076, 437.4255, 366.8581, 265.5489, 
    220.6245, 207.5233, 145.059, 52.48993, 0.02635965, 0, 0, 0, 0,
  312.5654, 332.0361, 48.98602, 0.01820307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2560336, 10.64937, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6525263, 85.40112, 154.1216, 
    145.2693, 104.7963, 68.44398, 59.66086, 5.658707, 51.90486, 0, 
    0.0002234011, 0.002236324, 0, 4.058273, 2.615149, 0, 0, 0, 0, 0, 0, 0, 
    45.61565, 143.503, 253.2654, 347.6613, 440.0746, 419.2403, 373.5648, 
    356.8692, 343.2001, 372.7208, 395.3455, 415.5849, 430.8153, 461.9744, 
    506.336, 526.5826, 478.6951, 428.0603, 393.4123, 322.4732, 237.9073, 
    211.1528, 175.5259, 95.53486, 5.59942, 0, 0, 0, 0, 0,
  277.1137, 216.7668, 65.78798, 0.01913495, 0, 6.423023, 0.05600383, 0, 0, 0, 
    0.008824782, 0.03805306, 5.421787, 6.542611, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.47252, 
    50.65664, 159.9921, 46.69725, 1.587591, 2.254171, 0.6875598, 155.2946, 
    109.7841, 0, 0, 0, 0, 6.335535, 1.460464, 0, 0, 0, 0, 0, 0, 0, 
    0.001764559, 51.18093, 107.6214, 220.6243, 313.7549, 357.301, 394.333, 
    380.0004, 369.1454, 378.0013, 370.4623, 409.9088, 457.2517, 510.6886, 
    598.5809, 591.0898, 488.7568, 418.8461, 368.6212, 287.8756, 211.7777, 
    183.3996, 128.3429, 26.55859, 0, 0, 0, 0, 0, 0,
  212.3771, 135.9476, 49.42075, 12.49728, 1.597956, 29.35641, 0.7934011, 
    2.107809, 0.008830293, 0.1460706, 1.322528, 19.1708, 1.042597, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1036084, 1.6234, 0.4369082, 1.249874, 151.7508, 
    165.1876, 0.1203202, 0, 0, 0.966633, 12.21299, 9.954236, 0, 0, 0, 0, 0, 
    0, 3.324982, 15.32631, 53.0812, 144.7708, 241.6709, 340.8276, 409.1607, 
    415.9962, 398.8717, 383.6034, 399.2011, 408.1645, 448.2938, 490.6762, 
    554.4016, 678.0546, 651.3043, 520.1175, 420.8705, 346.4621, 250.8538, 
    183.0857, 142.4498, 71.22203, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.2228342, 92.88892, 92.60233, 105.3637, 26.52375, 48.40273, 
    0.01253158, 0.2781332, 0.141384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2986155, 
    21.97212, 8.348226, 29.30048, 39.99499, 130.1351, 0.8950866, 0.01966914, 
    0.1630157, 0, 1.952829, 0.5040591, 0, 0, 0.01611275, 9.610229, 1.459349, 
    12.85996, 65.72018, 116.1776, 128.0019, 182.2513, 290.8639, 369.8836, 
    386.0753, 385.8762, 379.3724, 393.9282, 482.3826, 500.4763, 549.5696, 
    534.1202, 548.6902, 680.6912, 636.6417, 504.3287, 394.722, 296.3079, 
    208.9966, 140.6372, 97.57526, 13.33891, 0, 0, 0, 0, 0, 0, 0,
  3.996322, 0, 0, 0, 50.35525, 185.5548, 442.7651, 434.7867, 141.749, 
    8.424508, 0, 0, 0, 0, 0, 0.1385595, 0, 0.002443571, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001546636, 0, 
    0.01753371, 0.1784294, 55.34111, 40.54953, 0.06547624, 0, 18.5789, 
    0.6467119, 0, 0, 0.177912, 16.41363, 1.020464, 0, 0, 0.602079, 19.27653, 
    21.5851, 68.39326, 126.2266, 171.0694, 149.9013, 169.6777, 212.8275, 
    259.4587, 299.9385, 330.8089, 379.1569, 457.7391, 561.8567, 588.5029, 
    657.3253, 569.2491, 539.7734, 651.1829, 576.2408, 456.6287, 351.4606, 
    268.712, 186.3495, 104.8361, 52.63164, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0005410447, 0, 0, 217.2333, 150.0148, 147.8175, 59.43842, 0.09743718, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.004347128, 0.0005053915, 0, 0, 0, 0, 0, 
    108.7065, 172.8124, 10.6465, 39.72498, 0, 0.7019937, 0.6240747, 
    0.03666175, 3.923619, 11.28015, 0, 0, 0, 3.333197, 1.626409, 22.94781, 
    129.1699, 146.3097, 179.6523, 197.7332, 215.7947, 216.2458, 233.5067, 
    262.7396, 313.8624, 413.2129, 513.4584, 611.7216, 655.2258, 697.314, 
    587.9772, 544.4241, 623.3768, 528.1633, 394.2646, 303.2613, 223.6158, 
    176.0974, 98.5352, 40.67016, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.232757, 299.1098, 203.6477, 310.9305, 75.55457, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.001199378, 0, 0, 0, 0, 0, 424.0066, 651.8306, 74.5641, 
    110.6031, 137.6324, 0, 13.58554, 3.612053, 0, 0, 0, 0, 0, 4.653972, 
    12.98408, 132.1312, 225.6729, 202.1573, 187.3596, 223.9869, 245.0216, 
    232.7687, 241.0014, 265.6889, 318.4467, 431.9607, 541.9741, 643.3138, 
    668.8045, 639.2117, 512.8416, 507.6131, 530.3688, 426.9925, 321.1112, 
    237.3463, 202.2683, 173.7212, 111.4122, 27.88606, 0.0005438055, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 7.312272, 276.3273, 222.199, 363.1713, 12.21931, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90.08727, 874.5997, 248.2439, 134.9055, 
    106.5157, 0.7966748, 0.7750768, 0, 0, 0, 0, 0, 0, 0.2795637, 82.28407, 
    222.2338, 273.5854, 174.7247, 157.3741, 226.9098, 240.163, 230.1125, 
    254.5082, 294.148, 347.3311, 423.4855, 534.6428, 652.4855, 646.5594, 
    522.6107, 419.5539, 415.7138, 385.7757, 312.2747, 240.9982, 187.6149, 
    173.349, 160.6252, 114.4855, 27.0409, 0.0163472, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 160.1758, 213.3217, 235.5445, 48.00871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1112008, 2.781888, 0, 0, 0, 0, 0, 0, 0.003032611, 0.002118202, 
    0.5433614, 129.5313, 49.79841, 273.5827, 358.0385, 0.1867804, 9.040846, 
    16.79832, 2.512043, 0, 0, 0, 0, 0, 35.23597, 159.6615, 147.6077, 
    74.15279, 137.9986, 222.0329, 251.3415, 221.7983, 254.7236, 313.5164, 
    386.5862, 445.4337, 529.6935, 615.8958, 546.6193, 383.2585, 296.0247, 
    296.5038, 254.086, 225.9015, 197.0486, 177.1107, 159.7694, 143.3112, 
    134.4598, 60.69848, 9.276337, 0.07938728, 0.01935789, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 27.43061, 219.741, 182.4642, 145.6093, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14.73238, 8.035018, 0.002533916, 53.32179, 
    714.6627, 33.22498, 0, 0.08153576, 0, 0, 0, 0, 0, 0.1116458, 37.3478, 
    87.57549, 65.60155, 24.98499, 84.27135, 185.5645, 240.6545, 223.1828, 
    218.4679, 277.7992, 354.8269, 407.7614, 464.1208, 475.2428, 366.5284, 
    234.6922, 185.0667, 166.5074, 146.0874, 128.0777, 140.4522, 156.122, 
    159.8683, 152.9146, 170.7601, 142.2226, 55.40218, 25.69629, 0.2789844, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 118.9879, 364.7967, 262.5878, 200.3751, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0001877957, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.174198, 31.60677, 64.70731, 426.1732, 
    1363.807, 80.13299, 0, 0, 0, 0, 0, 0, 0.001290981, 2.815794, 26.87397, 
    19.16058, 8.644664, 1.876151, 39.90991, 143.068, 242.9099, 243.2124, 
    226.8486, 243.0945, 292.6472, 323.9382, 340.012, 310.8246, 220.8903, 
    156.6606, 105.6535, 84.0586, 78.32101, 71.50745, 87.09168, 128.866, 
    135.5459, 129.0692, 191.9514, 186.9409, 94.13192, 30.83496, 1.997563, 0, 
    0, 0, 0, 0,
  0, 0, 0.001936688, 46.618, 536.6373, 662.6491, 249.3386, 9.803163, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0001813781, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.459199, 103.5565, 
    661.9141, 1840.713, 219.5788, 0, 0, 0, 0, 0, 0, 0.1876374, 0.1116077, 
    4.196786, 0.6972661, 4.548798, 0.01515518, 19.67255, 135.7905, 257.0113, 
    277.3361, 253.3402, 236.5977, 238.597, 251.8898, 254.7406, 193.7241, 
    141.234, 99.71603, 61.99655, 29.32073, 13.64046, -0.03668842, 26.70518, 
    81.82543, 91.48897, 122.1683, 146.8756, 124.3265, 10.31211, 9.660895, 
    54.39833, 0.2762197, 0, 0, 0, 0,
  0, 0, 9.334058, 13.71354, 852.7475, 1096.084, 774.6525, 27.61173, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3280411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.112605, 141.024, 
    649.2419, 1983.348, 335.0366, 8.158025, 0.01285483, 1.803418, 2.566564, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.23637, 88.12022, 180.32, 243.7138, 259.6231, 
    232.9355, 205.8438, 203.9321, 192.951, 139.2836, 88.90681, 58.0747, 
    29.76662, 21.18993, 11.34657, 5.685978, 55.80595, 145.4924, 131.7599, 
    161.3288, 202.1818, 105.8592, 47.85705, 21.31422, 9.101623, 0, 0, 0, 0, 0,
  0, 0, 8.083728, 68.44715, 763.899, 819.9758, 573.8215, 67.20765, 0.8818858, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7558494, 202.6879, 
    672.795, 1732.209, 589.0763, 7.808373, 5.980556, 7.959057, 2.644362, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.5032064, 14.71771, 71.34007, 168.8776, 270.6567, 
    303.8179, 249.176, 188.3204, 150.6268, 103.42, 72.58722, 47.76024, 
    32.59775, 32.64248, 32.45184, 44.43424, 191.6641, 289.115, 320.5233, 
    411.2173, 393.0303, 296.0738, 190.0115, 73.94491, 0, 0, 0, 0, 0, 0,
  66.48343, 32.72926, 167.2516, 442.8591, 671.6302, 377.1797, 87.32704, 
    19.9507, 2.892875, 2.136357, 0.122568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003015865, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 80.25523, 370.7058, 1206.437, 775.0638, 72.39935, 
    11.08876, 20.55738, 1.923679, 0, 0, 0, 0, 0, 0, 0, 0, 0.7043098, 
    1.508858, 23.05793, 109.5643, 245.116, 339.6685, 319.9632, 211.4899, 
    138.8699, 98.34061, 73.37244, 64.12723, 38.16045, 37.41049, 28.51176, 
    38.78846, 65.09164, 118.0438, 185.5842, 257.3457, 215.2173, 108.8992, 
    78.36304, 35.72548, 8.264409, 4.238366, 0, 0, 0, 0,
  239.6041, 383.8715, 385.9552, 312.772, 354.1241, 158.2608, 13.44928, 
    4.439478, 0, 0, 0, 0, 0, 0.09766659, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004302262, 0.0009284276, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 65.84852, 257.2979, 725.2047, 976.9874, 203.7428, 
    26.53415, 26.40429, 12.97825, 0.3968416, 0, 0, 0, 0, 0, 0, 0, 0.2833899, 
    4.319847, 22.68953, 64.89889, 145.0534, 252.3569, 284.3854, 198.8476, 
    134.2758, 109.1641, 94.01095, 84.8871, 77.70658, 60.97504, 74.0986, 
    72.99908, 65.58603, 81.69981, 146.6016, 168.7964, 71.73798, 47.58058, 
    76.26965, 85.34253, 80.94412, 51.16417, 1.088907, 0, 0, 0,
  35.46908, 312.2523, 343.7193, 52.41047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1450596, 0.2184766, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.563134, 211.3301, 
    384.9349, 1012.969, 418.6268, 39.3827, 21.14776, 22.11357, 1.319225, 
    0.0001826946, 0.325497, 7.54947, 17.82139, 17.77085, 7.49655, 7.957342, 
    17.79939, 33.27032, 62.76324, 85.09935, 112.5088, 181.6462, 216.9371, 
    186.2492, 155.3895, 145.2876, 116.1752, 123.2312, 99.18019, 108.5044, 
    122.6949, 130.1461, 147.0177, 165.934, 161.3787, 95.41556, 49.94404, 
    50.94572, 86.07488, 121.9567, 174.7541, 113.5709, 7.699672, 0, 0, 0,
  0, 0, 0.5505809, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001916892, 
    0.488546, 0.3526058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01420734, 0, 156.4859, 171.2163, 
    1219.024, 1056.763, 227.3387, 20.19563, 22.60979, 1.255557, 6.144281, 
    45.4059, 62.7279, 97.57623, 101.1371, 78.44479, 56.55574, 70.73415, 
    121.4387, 190.2598, 228.6013, 167.1219, 186.6875, 214.2366, 206.5289, 
    194.4333, 173.067, 148.9911, 138.2063, 137.0002, 114.045, 110.0555, 
    138.2256, 143.1514, 155.9583, 107.2437, 61.62659, 60.00345, 62.52522, 
    75.2979, 158.1422, 252.193, 158.513, 1.751702, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002090689, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.008890191, 0, 67.49846, 202.0233, 1369.146, 1749.797, 
    579.0088, 20.74646, 6.495084, 0.0398635, 0, 0.4435986, 33.07759, 
    104.0203, 126.4093, 121.4114, 170.4067, 174.3627, 297.59, 418.0954, 
    490.278, 321.4501, 244.4302, 235.4262, 221.5576, 202.6546, 203.2396, 
    181.423, 183.7679, 160.8642, 143.6052, 126.7736, 119.1805, 123.6257, 
    103.5322, 71.23041, 75.24308, 72.00915, 65.68742, 95.67825, 220.7509, 
    320.3375, 166.0607, 14.94885, 1.212338, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3.35338, 0, 0, 0, 0, 0.0004769792, 0, 
    0.002373848, 0, 0, 0, 0, 0, 0, 0, 0, 0.01198174, 0, 1.170512, 26.17266, 
    920.9006, 1707.259, 548.358, 20.86545, 0, 0.02919498, 0, 8.295179e-05, 0, 
    0, 35.60873, 140.6726, 286.2187, 453.8871, 521.0576, 613.5406, 659.2684, 
    461.6195, 300.6107, 239.819, 229.6721, 231.9149, 274.6986, 262.3438, 
    217.9245, 185.6427, 156.8371, 124.7931, 111.6993, 114.7953, 105.9933, 
    95.67621, 83.49066, 78.79841, 74.49798, 111.6916, 266.0449, 268.2371, 
    42.25449, 0.02493712, 6.948849, 14.83968, 1.402666,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02394337, 0.2515746, 1.703864, 0.6291896, 0, 0.9544802, 1.295154, 
    1.900995, 1.829548, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003334169, 0.03683696, 0, 0, 61.67533, 497.1606, 1393.26, 921.786, 
    59.75617, 0, 0, 0, 0, 0, 0, 6.670186, 82.0864, 333.7366, 541.2671, 
    570.7663, 536.9034, 532.7047, 394.265, 316.7436, 281.2391, 283.4858, 
    317.4317, 337.6651, 311.4881, 252.3808, 196.0773, 158.135, 125.2839, 
    134.8932, 179.5908, 192.6594, 129.4154, 113.4966, 95.49207, 84.65179, 
    142.4767, 365.9221, 196.9136, 16.26885, 0, 0.993293, 210.9197, 320.5146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02792097, 0.3531507, 0.003153964, 0.09298629, 0, 0, 0, 0, 0, 
    0, 0, 0.0001550621, 0.0009271714, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007608135, 
    3.504901, 0.001191585, 14.31241, 84.53024, 1429.565, 1028.788, 570.2425, 
    25.71225, 0, 0, 0, 0, 0, 0, 0, 0.09222035, 52.24155, 104.2645, 261.9759, 
    312.8363, 286.0649, 269.9135, 332.5363, 391.7218, 436.5949, 425.3459, 
    349.5745, 251.7458, 185.8572, 143.547, 127.1319, 162.576, 240.0095, 
    253.7423, 196.6642, 167.1082, 130.5137, 139.8822, 425.961, 584.0701, 
    310.1891, 38.10512, 0.02188468, 0, 361.8489, 634.4559,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001512036, 0.001056419, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15.89228, 0.001179482, 0, 21.14887, 913.0068, 
    631.769, 1033.281, 837.3952, 31.48905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40.69078, 178.1973, 265.3913, 266.2013, 311.1905, 385.2721, 539.8588, 
    509.8239, 403.6374, 271.508, 176.3666, 138.3279, 123.0365, 145.8404, 
    203.9677, 254.9663, 219.4427, 240.7227, 267.1184, 484.1792, 681.328, 
    560.1155, 64.38747, 0.4352941, 0.003382807, 21.7661, 322.7632, 527.2258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7188078, 0, 0, 61.33807, 32.43402, 0.02485147, 145.2208, 627.1351, 
    287.4496, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.030678, 173.7331, 291.2982, 
    273.0661, 228.335, 327.7041, 474.7168, 494.3539, 377.0089, 256.2113, 
    177.9035, 140.8263, 131.356, 217.1942, 248.0046, 340.0473, 375.9899, 
    423.7958, 646.5859, 890.8132, 866.5603, 245.1126, 0, 0.05396707, 
    15.20921, 54.39197, 211.3136, 100.6684,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004543338, 0.003639919, 0, 
    0, 0, 0, 0, 0, 0, 3.531564, 0, 0, 0.7084563, 78.24866, 42.92502, 0, 0, 
    190.1828, 388.3742, 0, 0, 0, 0, 0, 0, 0.0004599308, 0, 0, 0, 13.8153, 
    130.9336, 144.9227, 177.9052, 219.8537, 376.9983, 361.93, 311.2201, 
    244.8839, 182.8421, 166.0394, 252.0663, 336.3086, 451.3323, 625.0237, 
    672.2084, 702.3406, 778.5399, 890.1186, 667.5145, 73.84701, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005854287, 0.00247674, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.313361, 16.38288, 0, 0, 147.3413, 142.4732, 0, 
    0.01397031, 50.75145, 186.9594, 0.1209901, 0, 0, 0, 0, 0, 0.000225285, 0, 
    0, 0, 0.01659336, 0.8779683, 47.25842, 88.2861, 235.9072, 276.3875, 
    324.9, 309.995, 270.1249, 234.3954, 347.3555, 412.644, 514.5791, 
    475.2197, 635.9094, 686.1741, 527.5653, 319.2344, 137.6655, 58.22589, 
    0.5826872, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001475661, 0.08985677, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0006000945, 5.420241, 14.74992, 9.866526, 369.6528, 
    31.99669, 0, 0.6211213, 22.01926, 26.09454, 0.01676102, 0, 0, 0, 0, 0, 
    0.0003724534, 0.0007511377, 0, 0, 0, 0.01054211, 4.9378, 35.11487, 
    209.5712, 293.8589, 365.6923, 371.3261, 394.2154, 492.1788, 710.024, 
    811.8054, 617.807, 343.5852, 201.6402, 88.6078, 33.18766, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002061675, 0.3639224, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.565544, 67.44887, 210.6318, 174.2347, 0, 0, 
    0.02026485, 0.5374939, 1.169389, 0.06065548, 0, 0, 0, 0, 0, 0.0005888037, 
    0, 0, 0, 0, 0, 0, 0.1444359, 50.93018, 158.3956, 294.5731, 366.2896, 
    503.3458, 626.3784, 834.7375, 746.9637, 477.1703, 102.5894, 2.179536, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0016285, 0.005161504, 
    0, 0, 0, 0, 0, 0, 0, 0.1744462, 11.87143, 189.9295, 0, 0, 0, 0, 3.378064, 
    2.925041, 6.432992, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001116622, 
    2.862813, 19.07391, 72.97668, 86.10835, 181.0871, 146.8998, 161.6484, 
    63.05329, 18.52388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.587682e-05, 0.0007486434, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003512555, 0, 0, 0.004746107, 0, 0, 0, 0, 0, 0, 0, 0, 0.001910802, 
    1.540883, 1.139802, 0, 0, 0, 0.00339965, 0, 5.067101, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7.394003e-05, 0, 0, 0, 0, 0, 0, 0, 0.1596736, 0.01119117, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002488717, 0, 0, 0, 
    0.00192382, 0, 0.0008238192, 0, 0, 0, 0, 0.004534618, 0.01042992, 
    128.6895, 111.6004, 0.9109875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 51.51996, 6.180326, 1.820795, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001911541, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009544371, 0, 24.92486, 51.07422, 23.80963, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.353347, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.248243, 20.32495, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.077861e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.002998321, 0.00326913, 0, 30.07554, 20.11271, 3.618359, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1637487, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001798506, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.00186227, 0, 0.03316185, 16.06968, 162.5954, 0, 
    3.422852, 0, 0, 0, 0, 0, 0, 0, 0.01038289, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001204468, 0, 0, 0.002527093, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66.34259, 22.89227, 15.44103, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001601016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06553058, 0.5628351, 51.22266, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9606495, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002309131, 
    0.6115905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.192964, 73.24959, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00447468, 0, 0, 0.001755983, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002103772, 1.21489, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 87.1916, 75.72276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.003544959, 0, 0, 0, 0, 0, 0, 0.0002654338, 0.001121242, 
    0.004204868, 0.001509032, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.04547353, 5.79191, 1.342976, 0.6890895, 0.2234796, 61.70195, 
    24.68652, 0, 0, 0, 0, 1.058887, 146.1155, 5.113419, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001511727, 0.00117502, 0.001633006, 
    0.007605216, 0, 0, 0, 0, 0, 0, 0, 0, 0.04061029, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1014451, 0, 1.253367, 0.0007692035, 16.09134, 27.76863, 48.46694, 
    11.74502, 0, 0, 0, 4.819854, 6.666916, 2.695935, 0, 0, 0, 0, 0, 0, 
    0.01972353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202.3895,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0006035659, 0, 0, 0, 0, 0, 0, 0.01408904, 0, 
    0.003578367, 0.004032353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03354037, 0, 0, 7.591219, 30.95796, 10.42947, 11.57776, 0, 0, 0, 
    2.446361, 0.008315299, 0, 0, 0, 0, 0, 0, 0.5451445, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 120.6041, 854.0955,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001588834, 0, 0, 0, 0.005239161, 0.009033938, 
    0.0005203752, 0.001356567, 0.001431737, 0.006111554, 0, 0, 0, 0, 0, 
    0.02182276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007873155, 0, 0, 0, 0, 0, 0, 
    18.8254, 15.31145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.272007, 709.054, 928.3032,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002614032, 0, 0.007351434, 
    0.003707968, 6.454103e-05, 0.001235135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0002616841, 0, 0, 0, 0, 0, 0, 0, 0.2473145, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    463.5101, 849.1191, 684.9581,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004843049, 0.002349587, 
    0.01799333, 0.00371025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004212329, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.004271484, 0, 0, 0, 0, 0, 0, 0, 0, 57.22657, 460.95, 639.7565, 
    519.5239, 33.79907,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001354043, 0, 
    0.006613636, 0.007528742, 0.02743311, 0.01341464, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003410095, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05400946, 4.694293, 0.3870355, 0, 0, 0, 0, 0, 141.1749, 
    601.933, 831.244, 543.7769, 58.66973, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01415738, 0.04210776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.679655, 
    105.733, 8.447727, 0, 0, 27.24204, 24.39606, 7.753161, 352.5742, 
    608.2495, 37.65978, 0.09178872, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01123114, 0.01882986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29.1145, 27.4687, 
    38.2424, 74.43308, 193.5007, 196.5712, 7.365326, 66.00092, 2.113855, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01327394, 0.003187717, 0, 0, 0.002941251, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.80582, 
    74.16306, 226.1258, 582.3444, 525.9813, 293.4045, 129.4705, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0153161, 0.005200402, 0, 0, 0, 0.003570459, 0.002388353, 0, 0, 0, 0, 
    0.1976552, 0, 0, 0, 0.1872808, 0.7276393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3034186, 214.9815, 492.9658, 326.6951, 
    73.56389, 0.05476749, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002162333, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9388899, 
    193.1229, 6.378803, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 258.6678, 289.7753, 3.976977, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.009249282, 0.001536941, 0, 0, 0, 0, 0, 0, 0, 40.0586, 
    32.99025, 2.803985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.30081, 1.451902, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0009401445, 0.0004037078, 0, 0, 0, 0, 
    0.1391184, 50.75321, 3.125369, 1.116508, 0.2084151, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933637, 0.05200977, 
    1.095076, 0.4746633, 0, 0.0152259, 0.00121065, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003794074, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.873821, 0, 0, 0, 
    0.0909774, 0.106935, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04739007, 0.5167308, 
    0.02355359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005289078, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0004078763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.796603,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.600741e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008196245, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2539265, 0, 
    0.1848694, 0, 0, 0, 0, 0, 0, 0.02119472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.612157,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009860342, 0, 0, 0, 
    0.5821458, 1.014729, 1.475074, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007580966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00020889, 0.003413063, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.08453731, 0, 0.6124651, 0.0904895, 0.04531468, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.060883, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006160314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0004963353, 0, 0.002697561, 0, 0, 0, 
    0.002501344, 0.003084639, 0, 0, 0, 60.34301, 23.29774, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001295554, 0.002088146, 0, 0, 0, 0, 0.003850434, 0, 0.003216584, 
    0, 0, 6.297387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2759891, 0, 0, 0, 0, 1.456678, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002685973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.603688, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.042054e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003275427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001260254, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004184085, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001634963, 0, 0, 0, 0, 
    0.00182365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004781314, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002623971, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1032847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02264775, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01294437, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45.58595, 
    19.94605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01843011, 0, 0, 0, 0, 0.0006814443, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05284531, 0, 0.2416257, 0.6087035, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01169867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009131898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006104111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002335767, 39.18405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0105723, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01319931, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1318502, 0, 0, 0.3468482, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45.02456, 0.7059237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0927918, 0.01668262, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0472814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    140.8308, 155.7868, 125.8311, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02154752, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    749.9999, 457.7867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.01483413, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.498203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002601753, 
    0.002704989, 0, 0, 0, 0, 0, 0, 0.001969324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003557655, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02448131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00550229, 0, 0, 0, 0, 0.0046798, 
    1.793624, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.448954, 0, 
    0.00866163, 0, 0, 0, 0, 0.4479904, 0.01966327, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005507405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.460738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03048245, 
    61.25506, 0, 0, 0, 0, 0, 0, 0.3824942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02183831, 
    0.2123545, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04637172, 
    0.008339238, 0, 0, 0.03448581, 0, 0, 0, 0, 0, 0, 0, 0.196157, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005239569, 
    0.0212123, 0.0003524371, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02602657, 
    0.02576878, 0.0369913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01774269, 
    0.006849611, 0.01812511, 0.007378699, 0.04169989, 0, 0, 0, 0.0002408772, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
