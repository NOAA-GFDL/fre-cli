netcdf atmos_tracer.bk {
dimensions:
	phalf = 50 ;
variables:
	float bk(phalf) ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:missing_value = 1.e+20f ;
		bk:_FillValue = 1.e+20f ;
		bk:cell_methods = "time: point" ;
	double phalf(phalf) ;
		phalf:long_name = "ref half pressure level" ;
		phalf:units = "mb" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;

// global attributes:
		:filename = "00080101.atmos_tracer.tile1.nc" ;
		:title = "ESM4_piClim-NTCF" ;
		:associated_files = "area: 00080101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "19.1" ;
		:git_hash = "5a324f5f5c98dbb620b25cd98a6add9da8861ee5" ;
		:creationtime = "Mon Jun  6 22:26:34 2022" ;
		:hostname = "pp212" ;
		:history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /xtmp/Luis.Sal-bey/ptmp/archive/oar.gfdl.bgrp-account/CMIP6/ESM4/AerChemMIP/ESM4_piClim-NTCF/gfdl.ncrc4-intel16-prod-openmp/history/00080101.nc --input_file 00080101.atmos_tracer --associated_file_dir /xtmp/Luis.Sal-bey/ptmp/archive/oar.gfdl.bgrp-account/CMIP6/ESM4/AerChemMIP/ESM4_piClim-NTCF/gfdl.ncrc4-intel16-prod-openmp/history/00080101.nc --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 00080101.atmos_tracer.nc" ;
data:

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;
}
