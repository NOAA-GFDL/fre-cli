netcdf atmos.1980-1981.aliq.04 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:18 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.04.nc reduced/atmos.1980-1981.aliq.04.nc\n",
			"Mon Aug 25 14:40:36 2025: cdo -O -s -select,month=4 merged_output.nc monthly_nc_files/all_years.4.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.491454e-05, -7.42517e-10, 0, 
    0, 0, 0, 0, 0, 0, 0, -1.623246e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -5.380911e-06, 1.278162e-05, 0, 0, -7.943193e-07, 
    0, -4.283098e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.757685e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.569328e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0003642836, 0, 0, 0, 0, 0, 0, 0, 0, -1.69733e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 2.499794e-05, 0, 0, -2.274656e-06, 0, 3.802678e-05, 0.0001548736, 0, 
    0, 0.0001461148, -3.910648e-05, 2.177815e-05, -5.702183e-06, 
    -1.807615e-05, 0, 0, 0, 0, 0, 0, 0, 0, -2.275796e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.438848e-05, 1.689035e-05, 0, 0, 0.0002735912, 
    4.110739e-06, -1.390127e-05, 0, 0, 0, 0, 0, 0, 0, 0, -3.504308e-06, 
    1.096253e-05, 0, 0, -3.188327e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.663719e-05, 0, -0.0001160957, 0, 0, 
    -4.58973e-07, 0, 0, 0, 0, 0, 0.000520047, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.566732e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.000994088, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.001996772, 0, -1.41573e-06, 0, 0, 0, 0, 0, 0, 
    0.0002055478, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.001046785, 0, 0.0005786567, -2.205904e-05, -3.797931e-05, 
    0.0005172273, 0.0006732095, 3.613427e-06, 0.001016858, 0.0006698571, 
    -0.0001283127, 0.0005283724, 0.001088517, -5.611428e-05, -2.28383e-06, 
    -2.673986e-06, 0, 0, 0, 0, 0, 0, 1.808198e-05, 0, 0, 0, 0,
  -6.411175e-06, 0, 0, 0, 0, 0, 0, 0, -1.760994e-05, 0.0007558836, 0, 0, 
    0.0007850931, 0.001337464, -1.795857e-05, 0, -5.497652e-06, 0, 0, 0, 0, 
    0, 0, -4.60356e-05, -1.135319e-05, 0, -8.360386e-06, -7.647077e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009899436, -2.690378e-05, -0.0001637936, 0, 
    -3.246882e-06, -4.819216e-06, -1.987635e-05, 0, 0, 0, 0, 0.001630046, 
    -3.776023e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.465536e-05, -6.841548e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.002605347, -3.649575e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -1.173088e-05, 0.003185465, 8.58631e-05, -3.112825e-05, 0, 0, 
    0, 0, 0, 0, 0.001077973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0006149225, 0.001077429, -2.17681e-05, 0.00138015, 4.679416e-06, 
    -0.0001548638, 0.0008132799, 0.002071628, 3.613427e-06, 0.001285653, 
    0.0008365569, 0.002655819, 0.0007053604, 0.001757712, -9.617e-05, 
    -1.154116e-05, -2.134986e-05, 0, 0, 0, -1.064672e-05, 0, -1.689933e-06, 
    0.0001522377, 0, 0, 0, 0,
  0.0005156765, 0.001432193, 0, 0, -6.294744e-06, 0, 0, 0, -1.802302e-06, 
    0.001536814, 7.243992e-06, 0, 0.0025377, 0.002892897, -2.900702e-05, 0, 
    -1.924178e-05, 0, 0, 0, 0, 1.588386e-05, 0, -0.0001186017, 0.0003889729, 
    0, -4.197845e-05, 1.213552e-05, -6.110913e-06,
  0, 0, 0, 0, 0, 0, -8.336983e-11, 0, 0, 0.003217523, -6.000705e-05, 
    0.000242894, -2.107283e-05, 0.001804488, -1.800736e-05, -5.503559e-05, 0, 
    -1.504726e-06, 0, 0, 0.002724583, -1.107371e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005358429, 0.0001516947, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 5.833304e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.575363e-05, 0, 
    0, 0, 0, 0, 0, 0, -1.745593e-05, 0, -4.414261e-06, 0, 0,
  0, 0, 0, 0, 0.004662332, 0.0002130163, 0.0003465379, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.134476e-09, 0, 0,
  0, 0, 0, 0, -2.644633e-05, 0.005483839, 0.001623294, -8.212028e-05, 
    -8.522567e-06, 0, 0, 0, 0, 0, 0.002235443, -1.962075e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.003859847, 0.001907267, -7.480653e-05, 0.00231231, 0.0004022267, 
    0.0002508449, 0.0009777647, 0.00686786, 3.613427e-06, 0.006852584, 
    0.001136127, 0.007399492, 0.002124379, 0.003945623, 0.0001527504, 
    -2.431104e-05, 4.151184e-05, 0, 0, 0, -1.419562e-05, 0, -5.154955e-05, 
    0.002099497, 0, 0.0001051962, 0, 0,
  0.0007842905, 0.001902923, 0, 0, -1.318253e-05, 0, 0, 0, 3.42615e-05, 
    0.004389359, 1.938693e-05, 0, 0.00495671, 0.007157575, 0.006136442, 0, 
    -5.095648e-06, 0, -2.242613e-05, 0, 0, 4.425204e-05, 6.048206e-05, 
    0.0005204447, 0.001314361, -5.744832e-06, 9.52542e-05, 4.258166e-06, 
    -2.095241e-05,
  0, 0, 0, 0, 0, 0, -1.500803e-05, 0, 0, 0.00707751, -9.208797e-05, 
    0.0004784295, -4.028161e-05, 0.005351774, 0.000549168, 0.001479737, 0, 
    -7.523631e-06, 0, -1.221895e-05, 0.004230457, -4.365374e-05, 0, 0, 
    -1.132373e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003892925, 0.0004622074, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 3.203591e-08, 0, 0, 0, 0, 0.0001087251, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.682603e-09, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0001876883, -1.332305e-05, 5.765285e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001294324, 0.0001907234, 0, 0, 6.24918e-05, -2.381428e-05, 0, 0, 
    9.300435e-06, 0.0005589972, 4.707368e-05, 0.0001594924, 0,
  0, 0, 0, 0, 0.006868374, 0.00192549, 0.002955829, 0, 0, -5.222852e-07, 0, 
    0, 0, 0, 0, -5.564366e-05, 0, 0, 0.001114702, 3.201319e-05, 0, 0, 0, 0, 
    0, 0.000234695, 0.0002750984, 0, 0,
  0, 0, 0, 0, 0.0003488423, 0.01261893, 0.003577997, -0.0001163299, 
    -4.141931e-05, 0, 0, 0, 0, -2.119976e-05, 0.007225475, 0.0001300664, 
    -8.592877e-06, -7.868065e-06, 0, -1.14644e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.005589811, 0.001925518, -0.0001303516, 0.002903703, 0.001546603, 
    0.001966262, 0.001200846, 0.01157992, -1.238554e-05, 0.01207376, 
    0.002713095, 0.01196643, 0.003341474, 0.009034036, 0.002254359, 
    -5.587597e-05, 5.367091e-05, 0, 0, 0, -2.839124e-05, 0, -0.0001189737, 
    0.004112622, 0, 0.001406834, 0, 0,
  0.00278799, 0.004873573, 0.0002497894, 0, -2.791e-05, 0, 0, 0, 
    0.0002077292, 0.009022266, 3.132122e-05, -1.040581e-05, 0.01014631, 
    0.01081318, 0.007707291, -2.63244e-06, 0.0002155673, -1.54071e-05, 
    -2.110991e-05, -1.414244e-06, 0, 0.0002191612, 0.00154495, 0.003197913, 
    0.003582189, 2.150391e-05, 0.002518157, 0.0005397978, 0.0002066073,
  0, 0, 0, -3.233098e-07, 0, 0, -5.645521e-05, -6.306695e-06, 0, 0.01165058, 
    -1.243701e-05, 0.004787448, 0.000782471, 0.00941091, 0.001938012, 
    0.004375837, 8.291355e-05, -4.878383e-05, 0, -2.129218e-05, 0.00930408, 
    -9.034853e-05, 0, -1.076161e-06, -2.499942e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01026602, 0.0006212945, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -7.576209e-06, 0.0001190188, 0, 0, 0, 0, 0.002951967, 
    0.0006933585, 0.0003159647, -2.831442e-06, -3.472732e-06, 0, 0, 0, 0, 0, 
    0, 0, -8.847248e-05, 0.0004063143, -2.902503e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.027991e-05, 0.0002107099, 0, 0, 
    -9.255886e-07, 0, 0, 0, 0, 0, 0, 0, -5.078373e-06, -1.084497e-06, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -7.828256e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.529753e-07, 0, -2.242147e-06, 0, 0, 0, 0, 0, 0, 0, -2.47863e-06, 0,
  -5.074226e-06, 0, 0, 0.001928769, 0.0004548107, 0.0001352988, 
    -1.494515e-05, 0.0006633236, 0, 0, -1.205303e-05, 0, 0, 0, 0, 
    -2.705473e-05, 0.00366916, 0.001011363, -9.43768e-05, -4.022543e-06, 
    0.001950041, 0.0009456906, 0, 0, 0.000733631, 0.00226802, 0.003018287, 
    0.002470974, 0,
  0, 0, -5.000813e-06, 1.135406e-05, 0.009534401, 0.00508503, 0.006239862, 0, 
    0, -7.581871e-06, 0, 0, -1.009456e-06, -1.463257e-06, 0.001182371, 
    4.877614e-05, 0, 0.0001333763, 0.003985526, 0.0005832363, 0, 0, 0, 0, 
    -1.50352e-05, 0.002109442, 0.00085243, 0, 0,
  0, 0, 0, -3.309896e-06, 0.001619932, 0.01844303, 0.004832704, 
    -7.262955e-06, 2.456336e-05, 0, 0, 0, 0, 0.0003570672, 0.01799121, 
    0.0004436375, -2.356659e-05, -4.422884e-05, 0.0008480866, -2.392332e-05, 
    0, 0, 0, 0, -3.124979e-06, 0, 0, 0, 0,
  0, 0.01052948, 0.004833025, -3.377893e-05, 0.004089096, 0.002627531, 
    0.006272356, 0.00290825, 0.02198784, -4.226273e-05, 0.01940807, 
    0.003578624, 0.01981042, 0.006678916, 0.01637574, 0.008166454, 
    -0.0001522252, 0.0002130977, 0, 0, 0, -9.529444e-05, 0, 0.0004123174, 
    0.005842687, 0, 0.002019091, -2.457303e-06, 0,
  0.007472226, 0.008393236, 0.0002841359, 0, 6.999153e-06, 0, 0, 
    -4.685812e-06, 0.000199888, 0.01451165, 0.000573453, 1.983681e-05, 
    0.01674252, 0.01945648, 0.01211298, -1.410554e-05, 0.0003982597, 
    -7.526905e-05, -3.108837e-05, -5.790953e-06, 4.669968e-06, 0.002500871, 
    0.002842449, 0.009286767, 0.004978022, 0.0001263523, 0.006852439, 
    0.001078604, 0.0001796783,
  1.31076e-05, 0, 0, 0.0001408459, 0, 0, -0.0001788377, -1.446967e-05, 
    -9.604384e-06, 0.01895422, 0.0009125306, 0.008728663, 0.005251018, 
    0.01645689, 0.003659393, 0.009950889, 0.0002918026, 9.227057e-05, 
    -4.384368e-09, 8.903802e-05, 0.01495959, -0.000171036, 0, -1.346336e-05, 
    -2.101217e-05, -4.484164e-05, 0, -6.976731e-08, -1.548109e-05,
  0, 0, 0, -1.073558e-06, 0, 0, 0, 0, 0, 0, 0.01567508, 0.001158472, 0, 0, 0, 
    0, 0, 3.39215e-05, -4.17804e-05, 0, 3.929247e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0003099985, 0.001199072, 0, 0, 0, -1.688197e-05, 0.01052241, 
    0.003622914, 0.001217157, 0.0008773331, 0.0004311634, 0, -1.283096e-05, 
    0, 0, 0, 0, 0, -0.0001387145, 0.0008069857, 0.0002007712, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -5.914002e-05, 0, 0, 0, 0, 0.0004674458, 0.002199156, 
    -2.879489e-05, 0.0002346341, 0.000580367, 0, 0, 0, 0, 0, 0, 
    -8.314475e-06, 7.933458e-05, 0.0001059995, 0.0001394932, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -4.411895e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.0004972162, -4.177029e-06, 0, 0, 7.565386e-07, 2.000182e-06, 0, 0, 0, 0, 
    0, -4.293656e-05, 0, 0, 0, 0.0001368033, -1.135146e-05, 6.597902e-05, 0, 
    0.0007693438, 0, 0.0007502539, 0.0001446547, 0, 0, -4.535804e-06, 
    -7.464055e-05, 0.0006559961, 6.037592e-06,
  -7.764473e-05, -4.136783e-05, 0, 0.004354771, 0.003927932, 0.002664308, 
    0.0004612252, 0.001963196, 0, 0.000221878, 0.0001911389, -5.458668e-06, 
    0, 0, -6.372472e-06, -0.0001067267, 0.009868866, 0.003217478, 
    0.001828405, 3.200834e-05, 0.009757398, 0.002510887, 0.001920741, 0, 
    0.001436873, 0.007871232, 0.007197787, 0.005716342, -2.95619e-05,
  0, 0, -5.317535e-05, 0.0004757857, 0.01436587, 0.006831999, 0.01521513, 0, 
    -1.080237e-06, 0.0004932195, 0, 0, -3.550604e-05, -0.0001079512, 
    0.004563219, 0.002258532, 0.0005844879, 0.002153908, 0.01054172, 
    0.002715355, 0.0006383528, -1.915427e-05, 0, 0, -3.369949e-05, 
    0.005763242, 0.002947228, 0.0001549959, 0,
  0, -2.861145e-06, 0, 4.616937e-05, 0.002286192, 0.0266669, 0.006066591, 
    0.0004690945, 0.001326711, 0, 0, 0, -8.357472e-08, 0.002474369, 
    0.03699875, 0.003912547, 2.831163e-05, 0.0004916746, 0.002016373, 
    1.257728e-05, -1.445641e-05, 0, 0, 7.39199e-10, 0.000513415, 0, 0, 0, 0,
  0, 0.02163761, 0.007860693, 0.003283771, 0.00727579, 0.008611652, 
    0.01381181, 0.005830721, 0.03901272, -2.97053e-05, 0.03307065, 
    0.01096453, 0.0310764, 0.01334757, 0.0280898, 0.01908761, -9.178442e-05, 
    0.0007839008, 0, 0, 0, -0.000121879, 0, 0.002008767, 0.01422437, 
    -4.750718e-06, 0.002700516, -3.417532e-05, 0,
  0.01348752, 0.01132821, 0.001372766, -4.88781e-06, 0.0004541487, 0, 
    3.80037e-07, 0.0001030796, 0.002520174, 0.02317044, 0.004021117, 
    0.001429878, 0.02228298, 0.03991046, 0.01811255, 9.536427e-06, 
    0.0006511107, 6.362843e-06, 0.0009632052, -3.579992e-05, -2.81774e-05, 
    0.006194804, 0.004484865, 0.01971339, 0.01145012, 0.0005314135, 
    0.01259552, 0.004564326, 0.003044491,
  0.0002280543, 0, -2.621183e-06, 0.0002721685, -1.156804e-05, 2.727015e-06, 
    -0.0001502463, -5.597451e-05, -0.0001003223, 0.02738216, 0.00375611, 
    0.02096477, 0.01336415, 0.03370394, 0.00689099, 0.01746084, 0.002682174, 
    0.0008691497, -6.009182e-06, 0.000898248, 0.02936874, 9.284841e-05, 
    9.569001e-06, 0.000157177, 0.0007103127, 8.768556e-05, 0, -2.935927e-05, 
    6.196614e-05,
  0, 0, 0, -2.374204e-06, 0, 0, 1.999305e-05, -4.45869e-06, 1.422038e-05, 0, 
    0.01843735, 0.003909592, -2.119132e-08, -5.995446e-08, 0, 0, 0, 
    0.0007746479, 0.0005437859, 9.90978e-05, 0.0001632224, 0, -3.091452e-06, 
    0, 0, -4.116079e-07, 0, -7.221708e-06, 0,
  0, 0, 0.0001858546, 0.0005392072, 0.002510902, -6.205758e-06, 0, 0, 
    -7.802156e-05, 0.01740222, 0.0147756, 0.002100166, 0.008555703, 
    0.001089604, 0, -2.566192e-05, 0, 5.701632e-05, 0, 8.271483e-08, 0, 
    0.0002977923, 0.001397395, 0.002236206, 1.270653e-05, 0, 0.002822629, 0, 0,
  0, 0, 0, -7.945695e-08, -6.442765e-06, -0.0001433952, 0, 0, 0, 0, 
    0.002823514, 0.00740031, 0.00297608, 0.00217304, 0.001806598, 0, 0, 0, 0, 
    0, 0, -5.007606e-05, 0.002512247, 0.0009075514, 0.0001604763, 
    1.673711e-05, 1.762324e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.227725e-08, 0, -1.106044e-05, -5.307126e-06, 0.0005439058, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.407148e-05, 0, -2.671451e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001442577, -3.581564e-05, 2.466236e-06, -5.149006e-06, 0.00114023, 
    0.0005350551, 0.00283247, 0, 4.717573e-06, 0, 0, 5.722572e-05, 
    2.526887e-05, 0, 0, 0.002889021, 0.002062971, 0.0005350773, 
    -1.342586e-06, 0.002875091, 0.003342555, 0.003393662, 0.003418272, 0, 0, 
    -6.466973e-05, 0.0001743541, 0.002046425, 0.003507502,
  0.0001983751, 0.0006449107, -1.237124e-07, 0.008674694, 0.009876116, 
    0.005556751, 0.003658874, 0.007389686, 0, 0.002758604, 0.003249267, 
    6.191082e-05, 0, 0, 0.00132201, 0.000927712, 0.01862156, 0.01065552, 
    0.02254722, 0.005238884, 0.02087396, 0.00916325, 0.007216358, 
    7.383194e-05, 0.004698929, 0.0188625, 0.01081587, 0.01492762, 
    -9.082178e-05,
  0, 0, -9.894543e-05, 0.004114062, 0.01805696, 0.01041333, 0.02615705, 0, 
    7.409535e-05, 0.004236687, 0.0006293466, 0.000151343, 0.00148058, 
    0.0001259119, 0.01036354, 0.01247216, 0.009298552, 0.008163625, 
    0.02531325, 0.01210521, 0.004162816, -7.797184e-05, 0, 9.863328e-10, 
    0.0001822864, 0.01342179, 0.009828911, 0.004166414, -2.924362e-06,
  0, -5.265978e-06, 0, 0.0003669831, 0.003658637, 0.0383542, 0.009437636, 
    0.001979597, 0.005212538, -4.174819e-06, 2.941233e-07, 3.751951e-05, 
    -3.977748e-05, 0.006707096, 0.05376659, 0.01530904, 0.004063819, 
    0.003780467, 0.007635097, 0.0001102606, -3.079184e-05, 0, -1.928892e-06, 
    2.347466e-06, 0.001558148, -3.135047e-06, -7.063603e-06, 0, 0,
  -1.182634e-06, 0.03594533, 0.0122608, 0.01289341, 0.01605295, 0.04273182, 
    0.04306468, 0.01852708, 0.06131133, 0.005856971, 0.05572088, 0.02531866, 
    0.05277481, 0.03421669, 0.05045089, 0.0471512, 0.002830253, 0.005968896, 
    0.0007564849, 0, -5.267756e-05, 0.0001913319, 2.66285e-09, 0.02011007, 
    0.02239512, 0.0001442251, 0.002544225, -0.000106737, 0,
  0.02685762, 0.0247549, 0.01375556, 0.0002372659, 0.003531081, 
    -7.272451e-06, -3.798152e-06, 0.001923183, 0.02452391, 0.05011558, 
    0.01603531, 0.007660755, 0.05184422, 0.068996, 0.03418409, 0.0003761837, 
    0.005179048, 0.001480526, 0.001637603, -3.25254e-05, 0.001408137, 
    0.01177338, 0.009961901, 0.06205924, 0.02451012, 0.001578942, 0.01879061, 
    0.009185145, 0.02212088,
  0.0006093006, -9.541009e-06, 0.0002650397, 0.0002827398, 0.0004172557, 
    0.001110117, 0.008041818, 0.0008351723, 0.0006184375, 0.03999509, 
    0.006500979, 0.03692949, 0.03418479, 0.06272755, 0.0114199, 0.03811093, 
    0.01126776, 0.004654341, 0.0004940925, 0.001523318, 0.04640736, 
    0.0009221823, 0.0006724049, 0.001527683, 0.00269022, 0.00409588, 0, 
    0.0002343433, 0.005392967,
  0, 1.249611e-09, 0, -3.640317e-06, 0.000129821, -3.650191e-07, 
    5.662848e-07, -9.119181e-06, 0.000299128, 1.586972e-06, 0.01859375, 
    0.01163955, 0.0005018564, 0.0002834735, 0.0002985634, -3.8642e-07, 
    -1.656451e-05, 0.007540185, 0.003989493, 0.004451464, 0.001840052, 
    0.0001742595, -1.518862e-05, 0.0002088635, 0, -5.246706e-05, 
    -7.123144e-07, 6.358651e-05, -1.548429e-07,
  0, 0, 0.001404856, 0.0008360329, 0.006244997, 0.000268502, 0, 0, 
    -0.0001236775, 0.03068572, 0.03084579, 0.009689393, 0.01826579, 
    0.004449766, -0.0001195728, -7.371244e-05, 0, 0.002410072, -6.954794e-06, 
    0.000249935, 0, 0.0004111118, 0.003594545, 0.00532771, 0.001775716, 
    0.0002392867, 0.005818154, 0, 0,
  0, -9.498573e-07, 0, 0.000825148, 0.0003941018, -0.000177877, -7.37441e-06, 
    -3.056434e-06, 0, -7.511301e-07, 0.003672027, 0.01339498, 0.007030529, 
    0.005144287, 0.004285551, -1.064683e-05, -4.255997e-06, 0, 0, 0, 0, 
    7.855817e-05, 0.005645757, 0.005530584, 0.0009744738, 0.002068321, 
    0.0009228333, 0, 0,
  2.414833e-05, 0.0002841261, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.027439e-07, 
    0.0009008424, 0, 0, 0, 0, 0, 0, -3.59729e-05, -6.844438e-05, 
    9.684405e-05, 6.391647e-05, 0.002936711, 0, 1.079128e-05, 0,
  -1.617908e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.702844e-06, 0, 0, 0, 0.0004453365,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0002522005, -2.247072e-06, 0, 0, 0, 0, 0, 1.47345e-05, 0, -2.423798e-05, 
    0, 0.0003990116, 0, 0, 0.0005342606, 0, 0.0001612779, 0.000372072, 
    0.0002400089, 3.367454e-05, 0.0004392044, 0, 0.0002620507, -5.280185e-06, 
    0, 0, 0.0001109412, 0, 0,
  0.005576322, 0.0002794621, 0.0002675778, -6.341986e-05, 0.005297206, 
    0.00324636, 0.008232424, 0.001617305, 0.002433467, -7.507878e-06, 
    -1.043455e-06, 0.003023901, 0.000219521, 0, -2.129266e-05, 0.006517626, 
    0.006667995, 0.002706252, 0.003820525, 0.007529317, 0.009444403, 
    0.01121165, 0.005976076, 0.001302878, 6.86115e-06, 0.002041047, 
    0.00132925, 0.00692712, 0.008373136,
  0.0006935495, 0.009147828, -3.32046e-05, 0.01674148, 0.01820531, 0.0118909, 
    0.008446326, 0.01248446, 0.0002720151, 0.003937592, 0.006477838, 
    0.00572979, -5.023821e-06, 0.001520924, 0.007055642, 0.005453921, 
    0.0327118, 0.0201158, 0.04639982, 0.02535388, 0.03687948, 0.01301998, 
    0.01842825, 0.002576421, 0.01064909, 0.03677243, 0.01731, 0.02851814, 
    0.006651564,
  0, -5.172476e-10, -9.414079e-05, 0.0123117, 0.02620292, 0.01275172, 
    0.04327111, -3.684309e-05, 0.00669751, 0.01025461, 0.002768069, 
    -1.772222e-05, 0.002167874, 0.005142277, 0.01953855, 0.04210574, 
    0.04114295, 0.0253464, 0.05762763, 0.0275469, 0.01908223, 0.001129474, 
    0.001836617, 0.005752801, 0.001057932, 0.02085812, 0.03526727, 
    0.008416151, -2.038748e-05,
  2.717696e-06, -1.811449e-05, 1.016564e-05, 0.01902519, 0.02358592, 
    0.04848856, 0.03143353, 0.007308553, 0.009937748, 0.0003521577, 
    0.0005561498, 0.0005004022, -0.0001458338, 0.0121445, 0.09655283, 
    0.06362545, 0.0512509, 0.01417659, 0.01883638, 0.001318056, 0.001153563, 
    -1.350519e-05, 0.0001562403, 0.007587147, 0.009174534, 9.96564e-05, 
    0.001657727, 6.567999e-05, -7.845222e-07,
  0.0005052452, 0.08847712, 0.03404428, 0.02767816, 0.03436262, 0.1487399, 
    0.1098908, 0.08681655, 0.1835693, 0.06293926, 0.09471174, 0.1139151, 
    0.1293776, 0.1726562, 0.1525193, 0.1485561, 0.05280983, 0.03651834, 
    0.007976235, 0.0001119396, 0.0002837158, 0.003322546, -3.727746e-06, 
    0.1088159, 0.07431468, 0.001580229, 0.005221626, 0.0001326601, 
    -1.784836e-05,
  0.1572473, 0.05810659, 0.07694396, 0.001064661, 0.02574665, 0.0011934, 
    0.0002562602, 0.01671107, 0.09186775, 0.1253297, 0.1266666, 0.06626648, 
    0.2428613, 0.1572765, 0.1270841, 0.01412432, 0.03948822, 0.01421602, 
    0.00649651, 0.004120219, 0.006796407, 0.02117123, 0.02104316, 0.2051055, 
    0.09907945, 0.009440914, 0.03862416, 0.02845775, 0.09859881,
  0.01038733, 0.00091257, 0.001898157, 0.001590122, 0.00306428, 0.004889197, 
    0.0630345, 0.01067113, 0.03509293, 0.06057941, 0.01901019, 0.08058169, 
    0.1586755, 0.1463615, 0.05298297, 0.07789488, 0.0394448, 0.01614474, 
    0.00279192, 0.006688526, 0.07264683, 0.01900184, 0.003886075, 0.02901433, 
    0.01810978, 0.01165206, 0.0002324437, 0.004362506, 0.04019536,
  4.754078e-05, -3.298251e-05, -6.657329e-06, 0.002583808, 0.0003682612, 
    0.0008407414, 0.0001456683, 0.0004063809, 0.002485442, 0.001218168, 
    0.02033383, 0.01953494, 0.01508819, 0.002145129, 0.003737099, 
    -6.417435e-05, 0.0005310623, 0.01711768, 0.01520583, 0.009990924, 
    0.0127094, 0.009134078, 0.000111505, 0.0007651256, -6.300424e-06, 
    0.0001638254, -0.0001192056, 0.001817033, -2.792222e-05,
  -4.084643e-07, -2.389517e-05, 0.006365528, 0.002070297, 0.01055547, 
    0.002928699, -5.694179e-06, 0, 0.001482127, 0.04914257, 0.05869124, 
    0.02562248, 0.0284487, 0.01471958, 0.004071401, 0.001460544, 
    0.0008170248, 0.007677023, 0.0001140214, 0.001175365, 8.464894e-05, 
    0.001275508, 0.005045796, 0.01008879, 0.007483672, 0.003740189, 
    0.009524593, -2.037937e-05, -1.352177e-08,
  -1.621419e-05, -1.133434e-05, -6.881189e-06, 0.002858071, 0.003168149, 
    0.0008924926, 0.0009118941, 0.0001666294, -5.987918e-06, -2.173157e-05, 
    0.005603558, 0.01810292, 0.01348075, 0.01232538, 0.0139086, 0.001374731, 
    0.0004243643, 0.0004595391, 2.369049e-06, -7.330621e-06, -5.328278e-06, 
    0.001645947, 0.0131389, 0.02013713, 0.004770944, 0.004033249, 
    0.001802408, 0, -6.622121e-07,
  0.004387329, 0.003368664, 0, 0.0002554704, 0, 0, 0, 0, 0, 0, 0, 
    -2.065767e-05, -4.433612e-05, 0.002522482, 0.003608047, -2.415365e-06, 
    0.0004525514, 0, -1.84719e-06, -3.809379e-05, -9.369237e-09, 0.001014984, 
    0.001794819, 0.004272254, 0.005563183, 0.005276019, 0.0006507075, 
    0.001865777, -4.1775e-05,
  0.0008749968, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9.068722e-05, 0, 0.001312271, -3.021142e-05, 0, 0, 0.001994224,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.285752e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.813935e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.233009e-05, 0, 0, 0, 
    0, -1.193859e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0008598578, 0.0002118149, -1.246055e-06, 6.009593e-05, 3.937063e-05, 
    -3.989117e-06, -3.488182e-06, 0.001049157, 0.0007887626, 0.0002048453, 
    -6.115402e-05, 0.0014557, 4.656583e-05, 0, 0.002359928, 0.001287896, 
    0.001127868, 0.00267175, 0.003853398, 9.738717e-05, 0.001500666, 
    -5.744387e-06, 0.002165671, 0.0005524001, 0, 0, 0.001516371, 
    -5.077414e-08, -5.211796e-05,
  0.01802603, 0.003222716, 0.002772301, -0.0002832846, 0.02139496, 
    0.01418134, 0.01562177, 0.008011462, 0.0062793, 0.0002826859, 
    0.0005440438, 0.007586235, 0.006907345, 0.002287542, 0.0005415068, 
    0.01125008, 0.01671, 0.01203276, 0.02834287, 0.013315, 0.01633989, 
    0.02063385, 0.009325545, 0.006225373, 0.001577938, 0.005428615, 
    0.004615878, 0.01200472, 0.02059864,
  0.01441101, 0.01587774, 0.00127951, 0.0289654, 0.02966128, 0.03065563, 
    0.01771018, 0.02589743, 0.003569285, 0.01557544, 0.01187045, 0.01342114, 
    0.001160824, 0.00635492, 0.02252874, 0.01517284, 0.05992096, 0.03976076, 
    0.08536835, 0.06433271, 0.07178305, 0.02604397, 0.02801156, 0.01291968, 
    0.01936715, 0.05533365, 0.02748248, 0.05270895, 0.02407063,
  0.002155503, 0.0007194297, 0.0004223525, 0.01916109, 0.03799945, 
    0.03034197, 0.09110881, 0.02459867, 0.05574779, 0.07045493, 0.01612849, 
    0.006664012, 0.004399883, 0.01286168, 0.04121006, 0.07939554, 0.1231794, 
    0.08056039, 0.1572583, 0.09554803, 0.04609235, 0.01491449, 0.005308593, 
    0.01582219, 0.01513339, 0.07290553, 0.0898235, 0.04675785, 0.0108138,
  1.425175e-05, 0.001078778, 0.03354124, 0.02952283, 0.09447181, 0.1161886, 
    0.08961155, 0.04776238, 0.05330282, 0.08540305, 0.01026809, 0.009741148, 
    0.008169742, 0.02749744, 0.126524, 0.1280289, 0.1148354, 0.1057081, 
    0.134578, 0.0507433, 0.03295251, 0.01726805, 0.01452242, 0.08067702, 
    0.0747288, 0.0475114, 0.06456658, 0.06297016, 0.01785705,
  0.0004112616, 0.1525034, 0.2346409, 0.08361483, 0.06585366, 0.1634444, 
    0.1340253, 0.09495728, 0.196488, 0.07601138, 0.1135797, 0.1203536, 
    0.1115207, 0.1459716, 0.1312523, 0.1426809, 0.09605721, 0.09396327, 
    0.05516383, 0.02574601, 0.02423145, 0.02647091, 0.01443983, 0.3000356, 
    0.1432807, 0.03511335, 0.03599962, 0.1002918, 0.001832095,
  0.1616823, 0.3019328, 0.3435864, 0.01708334, 0.06590933, 0.00894744, 
    0.01018984, 0.08323085, 0.3112293, 0.3260133, 0.1238312, 0.07813545, 
    0.2262603, 0.1444559, 0.09463473, 0.01683686, 0.03310531, 0.02479324, 
    0.02794179, 0.006912905, 0.01888026, 0.03639244, 0.05047566, 0.3241073, 
    0.2248655, 0.05379739, 0.09968653, 0.06394408, 0.1104555,
  0.07045685, 0.06785729, 0.01848816, 0.007625975, 0.04475805, 0.01846652, 
    0.09917049, 0.03788755, 0.04511814, 0.06929328, 0.02041598, 0.08012542, 
    0.141518, 0.1286289, 0.0771604, 0.1679843, 0.0918604, 0.05749995, 
    0.08549228, 0.08994025, 0.1596747, 0.06319625, 0.02814263, 0.09178723, 
    0.07414001, 0.04329398, 0.04351415, 0.03673127, 0.2514997,
  0.07218632, 0.02578668, 0.0003694522, 0.01667546, 0.04006175, 0.03600772, 
    0.03190547, 0.03427129, 0.04805852, 0.01981375, 0.04779333, 0.02476003, 
    0.03923632, 0.006720876, 0.02704398, 0.008844566, 0.007884413, 
    0.04315515, 0.1071033, 0.1056579, 0.152309, 0.07889364, 0.01607878, 
    0.03609123, 0.02084346, 0.05449631, 0.03748744, 0.03016616, 0.02061039,
  -9.165614e-05, 2.346068e-05, 0.009276429, 0.005071433, 0.02213768, 
    0.008725902, 5.980855e-05, -1.243692e-05, 0.00784322, 0.08936253, 
    0.1249918, 0.08550607, 0.07316715, 0.04248028, 0.02789451, 0.0110717, 
    0.009953491, 0.03367642, 0.003370366, 0.006328038, 0.002429805, 
    0.01086196, 0.01502078, 0.02569432, 0.01789072, 0.01651777, 0.02531509, 
    0.01399357, -1.295008e-05,
  -2.87146e-05, 0.0006997294, 0.0002239916, 0.00589778, 0.008703843, 
    0.001990754, 0.001899412, 0.0003280184, -2.906148e-05, 0.0005057696, 
    0.007914551, 0.02447568, 0.02936332, 0.032799, 0.03283951, 0.005617675, 
    0.002440743, 0.003165247, 0.001480019, -9.612379e-05, -1.440066e-05, 
    0.004893979, 0.02584517, 0.04727215, 0.01840731, 0.01260982, 0.002580352, 
    -4.640461e-06, -1.493962e-05,
  0.006850681, 0.004189451, -1.987647e-06, 0.0008004915, 0, 0, 0, 0, 0, 0, 0, 
    -6.274196e-05, 0.0006294323, 0.003713248, 0.005413662, -2.574777e-05, 
    0.002770097, 3.530944e-06, -1.297969e-05, -5.560969e-05, 0.0004519042, 
    0.001438871, 0.0047474, 0.01546658, 0.01602821, 0.01111825, 0.002032418, 
    0.004388527, 0.003190549,
  0.003919531, 0.0005012352, 0.001549352, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0001960316, 0.00219082, -1.84868e-06, 0.002373964, 
    -6.107322e-05, 0, 0.001457678, 0.001902784,
  0, -3.816521e-07, 6.974581e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0006908094, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -2.621954e-05, 1.402279e-05, 0, 0, 0, 0, 0, 0, 0, 0, -4.683275e-05, 
    -8.63993e-05, 0, 0, 0, -5.556822e-05, 0.001439648, 0.001367684, 
    0.0002351381, -1.384138e-05, 0, 0, 5.682087e-07, 0, 0, 0, 0,
  0.003662103, 0.003729818, 0.0003142728, 0.002439686, 0.001774873, 
    0.00020646, 5.591798e-05, 0.00106285, 0.002966222, 0.001152613, 
    0.0001901503, 0.003259576, 0.003093052, 0.0004542375, 0.003029374, 
    0.003574045, 0.004546427, 0.006293789, 0.01009993, 0.00552104, 
    0.009217199, 0.005258034, 0.003464399, 0.002688324, 0, -3.791618e-05, 
    0.002383025, 0.0006970049, 0.00117796,
  0.03617413, 0.02799691, 0.02469856, 0.005926077, 0.03675839, 0.03551292, 
    0.02994923, 0.02824465, 0.01995876, 0.009051225, 0.006785082, 0.01534737, 
    0.01461243, 0.009930166, 0.01159581, 0.02452728, 0.04409729, 0.04066772, 
    0.03700583, 0.05017201, 0.05934445, 0.06470793, 0.0303119, 0.01321737, 
    0.005780133, 0.01106401, 0.01631978, 0.02764385, 0.04264176,
  0.04901861, 0.03869605, 0.01646822, 0.05321, 0.08334974, 0.0645653, 
    0.04384543, 0.06466835, 0.03495675, 0.04235876, 0.06117768, 0.07723302, 
    0.02131275, 0.01497316, 0.04538783, 0.04503328, 0.1058308, 0.08666706, 
    0.1009761, 0.1591183, 0.1568961, 0.06971914, 0.05876435, 0.03563115, 
    0.05555293, 0.08218879, 0.05777111, 0.1150287, 0.1063688,
  0.03069807, 0.02368079, 0.00296962, 0.07613741, 0.08468609, 0.08101831, 
    0.1525958, 0.07351388, 0.1030944, 0.1542472, 0.1344111, 0.06991319, 
    0.02618793, 0.04557733, 0.05799118, 0.1386018, 0.1457658, 0.1204602, 
    0.1884815, 0.1679114, 0.1476625, 0.06272128, 0.04232416, 0.0409239, 
    0.03308434, 0.1119712, 0.159785, 0.119295, 0.07643252,
  7.447425e-05, 0.0004606042, 0.06621651, 0.02554412, 0.07656628, 0.09203835, 
    0.07933812, 0.04202002, 0.07492198, 0.0824717, 0.01284756, 0.00686333, 
    0.01005347, 0.04243711, 0.1273729, 0.1101542, 0.08906562, 0.07982165, 
    0.1156549, 0.03937917, 0.03472117, 0.005630614, 0.003369405, 0.06770586, 
    0.05445731, 0.06066421, 0.06166093, 0.07844345, 0.01436995,
  4.593549e-05, 0.1324287, 0.2103156, 0.06210005, 0.04591116, 0.1157728, 
    0.1115985, 0.06752247, 0.1596639, 0.05506615, 0.1026123, 0.09604623, 
    0.09288177, 0.1190105, 0.109585, 0.1134987, 0.05819171, 0.06800999, 
    0.02779501, 0.01278504, 0.0128997, 0.01863138, 0.002932573, 0.2522859, 
    0.1186847, 0.02116061, 0.02270885, 0.06575664, 0.0001273598,
  0.1261645, 0.2669976, 0.2676799, 0.01119198, 0.04665364, 0.005519452, 
    0.004249617, 0.05859095, 0.2485062, 0.2769687, 0.08088003, 0.05812607, 
    0.1751328, 0.1258941, 0.07208088, 0.007555767, 0.02131409, 0.0173195, 
    0.01979837, 0.00565938, 0.01003705, 0.02658389, 0.03872982, 0.2869126, 
    0.1863892, 0.04238757, 0.07685268, 0.04313807, 0.07759038,
  0.07394002, 0.0417702, 0.01241424, 0.05960302, 0.04683331, 0.0117051, 
    0.06463608, 0.0201904, 0.03075587, 0.05769339, 0.01389626, 0.06548169, 
    0.1241801, 0.112757, 0.05601109, 0.1409365, 0.1082187, 0.03993607, 
    0.046778, 0.05433396, 0.1278474, 0.04340062, 0.01145879, 0.04547648, 
    0.05919601, 0.02392115, 0.03388042, 0.009546474, 0.2048365,
  0.1069665, 0.07130566, 0.008711325, 0.0260953, 0.09699723, 0.0430594, 
    0.03213011, 0.01889715, 0.0383121, 0.01385989, 0.04265089, 0.02149414, 
    0.03654125, 0.003647734, 0.03624353, 0.01125079, 0.0121669, 0.04750925, 
    0.1175659, 0.1024248, 0.1259386, 0.07361891, 0.01969893, 0.05210729, 
    0.02146421, 0.1045635, 0.08117174, 0.04400752, 0.06701629,
  0.04258741, 0.01028168, 0.02616165, 0.01176761, 0.03985922, 0.04864455, 
    0.0285735, -2.633716e-05, 0.01869087, 0.124505, 0.1664373, 0.1511077, 
    0.1357538, 0.122386, 0.09905556, 0.06779496, 0.05264474, 0.04638656, 
    0.02224161, 0.02856429, 0.01510948, 0.08087128, 0.1357952, 0.09086291, 
    0.09042382, 0.1024, 0.0597954, 0.008148427, 0.02550464,
  0.0003451664, 0.003247032, 0.005292085, 0.01244049, 0.02109139, 0.02620025, 
    0.005624806, 0.0009321817, 0.008708064, 0.002655856, 0.02312013, 
    0.03790405, 0.0576249, 0.115062, 0.114229, 0.09729771, 0.04213079, 
    0.03961658, 0.02584709, 3.159266e-05, -1.080654e-05, 0.01151263, 
    0.04276345, 0.08371002, 0.04470561, 0.04144188, 0.01289521, 0.008534426, 
    0.00164175,
  0.01030426, 0.006199013, -6.011095e-05, 0.0007827983, -1.734332e-05, 
    -1.784961e-05, 0, 0, 0, -9.546335e-06, -1.229165e-06, 0.0007408118, 
    0.006602448, 0.009175678, 0.0107321, 0.00285424, 0.01609035, 0.008102822, 
    0.00345383, 0.001528113, 0.001803233, 0.002661985, 0.00756729, 
    0.02705367, 0.04218666, 0.03259712, 0.01589454, 0.0096803, 0.004748912,
  0.007892986, 0.002996314, 0.004916007, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.254051e-10, -1.622565e-05, -3.246349e-09, 0, -3.239472e-05, 
    0.002528994, 0.002731313, -1.668811e-05, 0.004074759, -8.385134e-05, 
    4.659355e-07, 0.002073738, 0.002544587,
  -4.36516e-05, -6.331866e-07, 0.0003494785, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001662886, -1.356599e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.268963e-05, 
    -2.716468e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -2.089912e-06, 5.276859e-05, -6.969876e-05, 0.0002457432, 0, 0, 0, 0, 0, 0, 
    0, 0, -5.209758e-05, 0.0005702644, -2.092862e-05, 0, -1.938022e-10, 
    0.001685112, 0.005059344, 0.009246091, 0.01035306, 0.004674559, 
    -4.335523e-06, -4.196043e-05, 5.659865e-05, -1.10363e-06, 0, 0, 0,
  0.007321055, 0.007465732, 0.004017835, 0.005624877, 0.01187042, 
    0.008555539, 0.009089328, 0.003292742, 0.01167604, 0.01150233, 
    0.01184638, 0.01179692, 0.01621937, 0.007233963, 0.007930059, 
    0.008998577, 0.02356426, 0.03874781, 0.04590357, 0.04095853, 0.04924474, 
    0.0204808, 0.01261358, 0.007935292, 0.0001782802, 0.001749964, 
    0.007108527, 0.003092788, 0.003368517,
  0.1160587, 0.09752508, 0.08994441, 0.04254631, 0.07083394, 0.11234, 
    0.09904528, 0.09491083, 0.06118073, 0.05023497, 0.06741509, 0.06742775, 
    0.07066061, 0.07853692, 0.04836573, 0.06474444, 0.09323625, 0.09278614, 
    0.09537325, 0.09179775, 0.1402622, 0.1567574, 0.1168879, 0.03463557, 
    0.03192733, 0.0459625, 0.04319175, 0.06633288, 0.1032311,
  0.1066938, 0.1062748, 0.08643401, 0.1272498, 0.1631719, 0.1184211, 
    0.08217861, 0.1060092, 0.08468635, 0.1133043, 0.1525705, 0.1440168, 
    0.08257478, 0.06930241, 0.06753815, 0.09664552, 0.166959, 0.142804, 
    0.1059158, 0.1639368, 0.1856286, 0.1127409, 0.1032967, 0.08503953, 
    0.1606504, 0.1881308, 0.1187771, 0.1892176, 0.1830996,
  0.02561586, 0.01977428, 0.07248709, 0.05368274, 0.07399515, 0.09043422, 
    0.1414578, 0.08225751, 0.109348, 0.1475918, 0.1529176, 0.08253626, 
    0.06275491, 0.05000979, 0.05787668, 0.1289953, 0.1248458, 0.08707655, 
    0.1649698, 0.1636941, 0.1240966, 0.04037888, 0.04483876, 0.03522396, 
    0.02185034, 0.0958168, 0.1437976, 0.1036927, 0.0460128,
  5.439506e-07, 0.0005854313, 0.04322333, 0.02997371, 0.06310207, 0.0818271, 
    0.06731702, 0.03266414, 0.08918457, 0.06287135, 0.003397111, 0.006311276, 
    0.008579614, 0.04858151, 0.1236063, 0.09523468, 0.06389501, 0.06470231, 
    0.09971981, 0.03248656, 0.02451643, 0.0005660424, -0.0001933869, 
    0.05798642, 0.04654231, 0.04570452, 0.03739095, 0.04583427, 0.003446854,
  4.963148e-06, 0.13885, 0.1784718, 0.05414963, 0.04279927, 0.09177887, 
    0.09893315, 0.05797484, 0.1488255, 0.05607328, 0.09645282, 0.07697816, 
    0.0867635, 0.1003157, 0.1054464, 0.09758551, 0.04799152, 0.06337266, 
    0.01785096, 0.005605213, 0.006311823, 0.005906138, 1.179877e-05, 
    0.2214689, 0.107293, 0.01665914, 0.02125706, 0.04138187, 4.007104e-05,
  0.1030233, 0.249032, 0.2175561, 0.006638411, 0.02966068, 0.006921811, 
    0.005455078, 0.04865963, 0.1940741, 0.2421638, 0.07105495, 0.04862427, 
    0.1498962, 0.1266393, 0.07528549, 0.007076913, 0.01273214, 0.01929625, 
    0.01187854, 0.00702406, 0.01007625, 0.02131479, 0.06131198, 0.2715945, 
    0.1666576, 0.04095114, 0.06241543, 0.03476155, 0.05485511,
  0.06568101, 0.02314766, 0.009628667, 0.0488974, 0.04205263, 0.008928574, 
    0.04997337, 0.0161345, 0.02142925, 0.05599341, 0.01504822, 0.06107188, 
    0.108013, 0.1006729, 0.04300212, 0.1276937, 0.1042581, 0.03852623, 
    0.03179685, 0.04648466, 0.1089046, 0.03241624, 0.006272197, 0.03162246, 
    0.03713299, 0.01599552, 0.01548317, 0.001922793, 0.1772581,
  0.1065273, 0.06349202, 0.005623911, 0.02375704, 0.08286643, 0.03665335, 
    0.03160129, 0.009375555, 0.03324701, 0.01504379, 0.02996678, 0.02082258, 
    0.02630173, 0.00479121, 0.0290845, 0.002798256, 0.007698046, 0.04193917, 
    0.07659261, 0.09745535, 0.1168714, 0.05949428, 0.0187172, 0.03993861, 
    0.01502152, 0.09882797, 0.07050805, 0.03295956, 0.06094669,
  0.06838133, 0.04095956, 0.05781413, 0.04937019, 0.07410494, 0.07632634, 
    0.06639625, -7.029163e-05, 0.03222988, 0.1549951, 0.1776289, 0.1464526, 
    0.1352183, 0.1310197, 0.1064907, 0.08091584, 0.07022295, 0.06118133, 
    0.04867245, 0.04165976, 0.04831154, 0.1068541, 0.1563117, 0.1095113, 
    0.1043713, 0.1328782, 0.1234323, 0.04086044, 0.05909559,
  0.02587617, 0.02859672, 0.04702494, 0.02944505, 0.0603501, 0.08683458, 
    0.01062495, 0.01696327, 0.03602416, 0.02263181, 0.04685132, 0.08773126, 
    0.1196961, 0.1801305, 0.2154159, 0.1982272, 0.1773163, 0.1751241, 
    0.1300699, 0.008475398, 0.0021739, 0.03231637, 0.1098684, 0.1655061, 
    0.1312409, 0.1085099, 0.1190305, 0.04676129, 0.04196574,
  0.02967213, 0.01180873, 0.003587517, 0.002295988, 0.003860528, 
    0.0009733736, -4.892864e-06, 5.969887e-05, -2.411619e-07, -2.329695e-05, 
    0.0002233262, 0.001351418, 0.01133689, 0.03133732, 0.04500671, 
    0.03790561, 0.05986297, 0.08126128, 0.05525081, 0.003817312, 0.00778859, 
    0.01280618, 0.02234649, 0.07387535, 0.09920619, 0.1022314, 0.06789115, 
    0.03931241, 0.0301662,
  0.01204059, 0.003430475, 0.007428105, 0.0006415662, 0.0005819818, 
    0.001765962, 0, 0, 0, 0, 0, 0, -4.439041e-06, -2.428898e-06, 0, 0, 
    -3.970095e-07, 0.0002470826, -2.970333e-05, 9.257929e-06, -6.427596e-05, 
    0.003891114, 0.004042408, 0.001391577, 0.02209073, 0.007109417, 
    0.01235929, 0.003324511, 0.01047853,
  0.002840708, 9.276086e-05, 0.0003903786, 0.000229623, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.541966e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.002846744, 
    -2.997312e-06, 0, -4.064606e-06, 0.001187086,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.55601e-07, 
    -6.983746e-05, 0.0001772714, -3.383321e-07, -6.394798e-06, -4.397371e-06, 
    2.864971e-06, -2.224243e-05, -1.615757e-06, -4.030903e-07, -2.613932e-07, 
    0, 0,
  -2.807154e-05, 0.003078224, 0.004698055, 0.001722567, -1.952923e-05, 0, 
    4.607781e-09, 0, 0, 0, -5.803042e-09, 0, -0.0001353777, 0.005628765, 
    0.001376785, -3.214299e-05, -6.707547e-05, 0.01714939, 0.03151383, 
    0.04472505, 0.02922034, 0.01072074, 0.01025158, 0.003316847, 0.003721688, 
    0.0001754425, -1.194806e-06, 0, 2.457776e-05,
  0.04359763, 0.04967793, 0.03545789, 0.05242883, 0.04909326, 0.04180579, 
    0.03850292, 0.02302362, 0.03268769, 0.03661307, 0.05625499, 0.06484134, 
    0.05465946, 0.05613622, 0.08302743, 0.07346438, 0.1039957, 0.1089737, 
    0.1232219, 0.1030973, 0.1228966, 0.07493485, 0.07085337, 0.07130418, 
    0.04034952, 0.02096533, 0.01845455, 0.01285722, 0.03885472,
  0.1590528, 0.1447499, 0.1663278, 0.1342109, 0.1440608, 0.1956798, 
    0.1626806, 0.1744408, 0.1260097, 0.116931, 0.1541842, 0.1522576, 
    0.1490508, 0.1384516, 0.1087705, 0.14927, 0.1572502, 0.1507538, 
    0.1418388, 0.1203337, 0.1962755, 0.1954603, 0.1731012, 0.07482457, 
    0.083597, 0.1096663, 0.09934358, 0.156915, 0.1683277,
  0.09663566, 0.09696744, 0.09407666, 0.1203218, 0.1431675, 0.09146561, 
    0.07972954, 0.1117269, 0.09396582, 0.1317071, 0.1499471, 0.150024, 
    0.08148526, 0.07323889, 0.0965092, 0.09883735, 0.164174, 0.1607902, 
    0.1155211, 0.1613936, 0.1848701, 0.1116167, 0.1192675, 0.1032377, 
    0.1740298, 0.2008353, 0.1342335, 0.1844946, 0.1736959,
  0.01576219, 0.01512355, 0.06564046, 0.03914529, 0.06709114, 0.08602031, 
    0.1193791, 0.06672238, 0.092391, 0.1206345, 0.1488221, 0.07389956, 
    0.07187938, 0.0472045, 0.04693635, 0.1110135, 0.1079522, 0.0935449, 
    0.1294746, 0.1460999, 0.1001134, 0.03253446, 0.03999894, 0.02475191, 
    0.01917848, 0.07704189, 0.1236793, 0.09223235, 0.02694809,
  5.527033e-07, 0.004264313, 0.02123629, 0.02369233, 0.04479492, 0.08547407, 
    0.06064593, 0.02854064, 0.08403265, 0.05535256, 0.001344326, 0.00785269, 
    0.01221093, 0.04176098, 0.1240711, 0.08098738, 0.04941103, 0.05969428, 
    0.09543024, 0.02777587, 0.007121422, 8.037135e-05, -0.0002557678, 
    0.04952345, 0.03966268, 0.04040314, 0.01683567, 0.0246829, 0.0005536017,
  1.671046e-06, 0.1431528, 0.1500319, 0.04543335, 0.0435646, 0.06491867, 
    0.08380152, 0.04532218, 0.1309808, 0.04486221, 0.09500684, 0.06760743, 
    0.0840161, 0.08208664, 0.09383168, 0.08404973, 0.03836805, 0.04878312, 
    0.007164486, 0.002691884, 0.001299053, 0.0002675349, 2.117505e-05, 
    0.1712669, 0.09299993, 0.01201598, 0.0212198, 0.02174977, 3.352581e-05,
  0.07968825, 0.2206647, 0.1531315, 0.007520256, 0.02088757, 0.00613363, 
    0.006409639, 0.03010314, 0.1273066, 0.1979908, 0.05781629, 0.03668349, 
    0.1154007, 0.1205553, 0.06857327, 0.008253012, 0.007860757, 0.02018996, 
    0.006552801, 0.003346414, 0.008163905, 0.01510324, 0.07739346, 0.232594, 
    0.1395428, 0.04824401, 0.05267143, 0.02473426, 0.04091842,
  0.03762606, 0.01416695, 0.008320819, 0.03089651, 0.03252354, 0.005983421, 
    0.03261489, 0.01368914, 0.01390821, 0.05418485, 0.01512701, 0.05427821, 
    0.09353159, 0.09527251, 0.04423444, 0.1192293, 0.08445154, 0.0394301, 
    0.02008122, 0.03808467, 0.09590256, 0.0223433, 0.003576363, 0.03225555, 
    0.03204248, 0.01668278, 0.006308493, 0.0005431921, 0.1367932,
  0.09493749, 0.04798412, 0.008646284, 0.02563188, 0.05910042, 0.0268894, 
    0.0238174, 0.002713552, 0.03193703, 0.01644061, 0.01953421, 0.01925364, 
    0.02622671, 0.005846216, 0.01951957, 0.00207254, 0.006589944, 0.02925868, 
    0.04511791, 0.08751499, 0.108282, 0.05004155, 0.01228059, 0.03097492, 
    0.01095688, 0.07424645, 0.05062129, 0.03706779, 0.06022625,
  0.07204993, 0.06741298, 0.07380708, 0.08669965, 0.09141503, 0.07824072, 
    0.0584423, 0.001936191, 0.05508939, 0.152139, 0.161458, 0.1466664, 
    0.1352291, 0.1184286, 0.09538177, 0.07211033, 0.05743542, 0.04597313, 
    0.04003264, 0.04164258, 0.05252441, 0.08602566, 0.1290903, 0.1015033, 
    0.08408423, 0.1401049, 0.1072029, 0.0384448, 0.079802,
  0.08823673, 0.0963394, 0.1257529, 0.07106724, 0.1287588, 0.1085004, 
    0.02534837, 0.1294777, 0.1091773, 0.05170199, 0.080285, 0.1142822, 
    0.1415263, 0.1937783, 0.2245645, 0.2068566, 0.1742818, 0.1945681, 
    0.1568878, 0.0647919, 0.01491406, 0.07893769, 0.1339441, 0.1555359, 
    0.1666926, 0.1486794, 0.141249, 0.08001933, 0.06896842,
  0.1231009, 0.04644328, 0.05959158, 0.03501777, 0.1163791, 0.01789336, 
    0.0005379657, -9.270463e-07, -4.886939e-06, 5.191252e-05, 0.005435873, 
    0.009479076, 0.03420138, 0.0498995, 0.06971408, 0.04690725, 0.09579754, 
    0.1596759, 0.1675276, 0.02974526, 0.0520239, 0.07417186, 0.06036279, 
    0.115303, 0.1491268, 0.1507891, 0.1247445, 0.07900899, 0.07378037,
  0.0400684, 0.0278431, 0.04952485, 0.04528858, 0.01856471, 0.008927431, 
    0.006561346, -4.503984e-06, 0, 0, 0, 0, -5.469718e-05, 0.0006131654, 
    0.001350639, 0.00895671, 0.001754037, 0.02874756, 2.42068e-05, 
    0.002855382, 0.002919394, 0.0121335, 0.01323124, 0.04625167, 0.1191189, 
    0.04846741, 0.02174806, 0.01139103, 0.03847606,
  0.01685082, 0.02814256, 0.01595402, 0.02592974, 0.009081057, 0.01023983, 
    0.008186823, 0, 0, 0, 0, 0, 0, 0.003455459, 0.001355676, 0.0005108778, 
    4.96841e-06, 1.681597e-05, -4.366668e-06, 1.261012e-05, -1.954417e-05, 
    1.209516e-05, -0.0004120459, -0.0025882, 0.04717159, -7.263522e-05, 
    -8.252264e-09, 0.00125825, 0.01408235,
  -1.203804e-05, 0, -2.126991e-11, 0.0002808615, 0.001595026, 0, 0, 0, 0, 
    -7.273187e-08, 4.891191e-09, 1.160535e-09, 0, 0, 0, 0, -1.648885e-06, 
    0.000293443, -1.206152e-05, 0, -1.588855e-05, 0.0004823605, -3.06286e-05, 
    -0.0001576557, -0.0001273002, 0, 0, -4.399137e-05, 1.55383e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.031457e-05, 0.001975097, 
    0.006580822, 0.002127596, 0.00313708, 0.0002266886, -3.816013e-05, 
    -2.530556e-05, 0.0005899339, 0.003290294, 0.001583895, -0.001197856, 
    0.004221086, 0, 0,
  0.0006000942, 0.007550743, 0.006860271, 0.008439645, -0.0001585451, 
    -4.425179e-06, 0.0005706686, 0.0001074312, -4.144085e-08, 7.560808e-05, 
    0.0009167262, -4.546981e-06, -0.0002954624, 0.01096928, 0.01381052, 
    0.01647839, 0.02027979, 0.04819269, 0.08632414, 0.1122458, 0.08658772, 
    0.08329593, 0.05354311, 0.01827286, 0.03000432, 0.009884503, 0.005751153, 
    0.004406927, 0.003014821,
  0.08410709, 0.08844637, 0.0796079, 0.09961786, 0.1041738, 0.08800133, 
    0.09199165, 0.07963333, 0.08915442, 0.1050391, 0.1185661, 0.173523, 
    0.1559319, 0.1496315, 0.1771563, 0.1811751, 0.1877931, 0.1638607, 
    0.2089819, 0.1424912, 0.1765349, 0.1539747, 0.1500637, 0.1887597, 
    0.1008552, 0.0695193, 0.0784006, 0.06560069, 0.07800418,
  0.1841918, 0.1680168, 0.1753081, 0.151507, 0.1458896, 0.2048717, 0.1660786, 
    0.1789475, 0.1520653, 0.1614362, 0.1986131, 0.20048, 0.1601521, 
    0.1495834, 0.1258799, 0.1531222, 0.1595739, 0.1495874, 0.1522912, 
    0.130592, 0.2117048, 0.186136, 0.1627242, 0.1272206, 0.128337, 0.1452041, 
    0.1259007, 0.1683037, 0.1883259,
  0.08378778, 0.08031449, 0.07559784, 0.1037086, 0.1236274, 0.07985646, 
    0.07926917, 0.09856685, 0.08517234, 0.1215563, 0.1330023, 0.1316255, 
    0.06691207, 0.06385971, 0.09277345, 0.0920718, 0.1545254, 0.1503154, 
    0.1181034, 0.1601987, 0.1772046, 0.0928835, 0.1316437, 0.1104977, 
    0.1432863, 0.1723783, 0.1210665, 0.1667223, 0.1716167,
  0.005888662, 0.005243994, 0.04483888, 0.03047116, 0.06036109, 0.09151842, 
    0.1156311, 0.05933613, 0.08507309, 0.08806194, 0.1432603, 0.06534681, 
    0.04616746, 0.03421136, 0.04440945, 0.1028579, 0.104969, 0.08113476, 
    0.1165076, 0.1345906, 0.1027374, 0.02710668, 0.03021666, 0.01227249, 
    0.01578411, 0.07109826, 0.1069048, 0.08026822, 0.02325259,
  3.467048e-07, 0.001020304, 0.008907985, 0.01280973, 0.03547199, 0.08804534, 
    0.06158138, 0.02856481, 0.06771065, 0.04550958, 0.0007614199, 
    0.006484382, 0.01614892, 0.04081533, 0.1137849, 0.06691808, 0.04027582, 
    0.05134687, 0.08620629, 0.02251523, 0.001399251, 0.0009227977, 
    -3.417502e-05, 0.04028789, 0.03193187, 0.03553956, 0.01107391, 
    0.009280031, 1.656309e-05,
  2.718977e-06, 0.1410445, 0.1256548, 0.04157542, 0.04001307, 0.04253482, 
    0.07218741, 0.03941784, 0.1085605, 0.03410871, 0.09860907, 0.06483532, 
    0.07960902, 0.06107993, 0.08014201, 0.06970406, 0.02629266, 0.03059782, 
    0.005220187, 0.001825097, 0.001123554, -0.0001311111, 7.876277e-05, 
    0.1131419, 0.08209717, 0.01156106, 0.01865546, 0.006760942, 9.727334e-06,
  0.05513132, 0.1851955, 0.1090969, 0.008432943, 0.01701931, 0.005733955, 
    0.00839749, 0.01543235, 0.07945388, 0.1587847, 0.05333515, 0.02332988, 
    0.08127919, 0.1045072, 0.06174364, 0.006656627, 0.006359383, 0.02128835, 
    0.006650963, 0.001207727, 0.006878911, 0.009041865, 0.07793616, 
    0.2022179, 0.1226429, 0.06473725, 0.05370363, 0.01959886, 0.03353076,
  0.02420004, 0.008517528, 0.006634728, 0.02227317, 0.02656974, 0.004306927, 
    0.02009302, 0.009673122, 0.009208904, 0.04887587, 0.01329169, 0.05091086, 
    0.07091699, 0.08316213, 0.05340774, 0.1076863, 0.07118435, 0.04359204, 
    0.00977762, 0.02139945, 0.07917878, 0.01389401, 0.002429051, 0.02728843, 
    0.03171313, 0.01769166, 0.003609459, 0.00420813, 0.1025433,
  0.09173796, 0.03322391, 0.007656939, 0.02680787, 0.04659851, 0.02031522, 
    0.009750679, 0.001087946, 0.02422369, 0.01409481, 0.01586599, 0.01656632, 
    0.02601661, 0.002867787, 0.01117148, 0.001219529, 0.005732019, 
    0.01886985, 0.04934603, 0.06196466, 0.09188064, 0.04149242, 0.009292893, 
    0.02607644, 0.007946704, 0.04839442, 0.03845475, 0.03273964, 0.06123742,
  0.06160785, 0.07306901, 0.064961, 0.07382154, 0.09848268, 0.07361558, 
    0.0513666, 0.003799717, 0.08494617, 0.1471901, 0.1492752, 0.1562875, 
    0.1436894, 0.1032584, 0.08203222, 0.06622057, 0.04404857, 0.03272725, 
    0.0353193, 0.03095456, 0.04976337, 0.07198232, 0.112137, 0.09607334, 
    0.07456596, 0.1292622, 0.1073055, 0.03293613, 0.05776747,
  0.1031905, 0.1140085, 0.1585544, 0.123285, 0.1316891, 0.1006022, 
    0.05194939, 0.2035078, 0.1741436, 0.09751235, 0.08630612, 0.1218719, 
    0.1402623, 0.187531, 0.2338113, 0.2074298, 0.1700416, 0.1720717, 0.1341, 
    0.1214208, 0.05586351, 0.1086347, 0.1264556, 0.1459734, 0.1592337, 
    0.1424642, 0.1431043, 0.07273035, 0.06105126,
  0.1948511, 0.1424533, 0.1408973, 0.1292572, 0.1394076, 0.07925281, 
    0.03173466, 0.001461046, 0.0003431154, 0.01615273, 0.03611773, 0.0164435, 
    0.0645963, 0.06332964, 0.1077544, 0.0566156, 0.1149895, 0.1950726, 
    0.2334241, 0.1133923, 0.1149023, 0.1308193, 0.1357735, 0.1293965, 
    0.1804145, 0.1591695, 0.1402117, 0.09299251, 0.1065364,
  0.1808149, 0.09725062, 0.1476266, 0.1261518, 0.1191557, 0.0593409, 
    0.0261598, 0.01204888, 0.000726523, -1.218787e-05, -5.501731e-08, 0, 
    -0.0002654734, 0.02629003, 0.02830075, 0.03076058, 0.03148803, 0.0737765, 
    0.03704824, 0.04908387, 0.06597693, 0.05933439, 0.09408129, 0.08109836, 
    0.198063, 0.08542433, 0.03094743, 0.04860862, 0.1265965,
  0.1198045, 0.1037828, 0.06938604, 0.09093633, 0.09776892, 0.05776995, 
    0.01721812, 0.02200803, 0.008379092, -9.177405e-06, -2.500515e-06, 
    3.392248e-05, 0.0003591171, 0.02235979, 0.03520679, 0.02087643, 
    0.01491349, 0.02796031, 0.02321984, 0.01983169, 0.03215333, 0.01414034, 
    0.02321397, 0.02315034, 0.09351349, 0.001379675, -2.299401e-06, 
    0.02740821, 0.06882845,
  0.01419317, 0.0172008, 0.01821739, 0.01483868, 0.01742032, 0.01836895, 
    0.01644483, 0.01552041, 0.005821259, 0.01101137, 0.02283811, 0.01040917, 
    0.007412968, 0.001170453, 0.004489939, 0.005345218, 0.008133729, 
    0.00799918, 0.007174316, 0.01637606, 0.02756057, 0.02779675, 0.004522516, 
    0.002352176, 0.005697716, 0.0002316921, -0.001098868, 0.005713065, 
    0.007017251,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0010033, 0.01978792, 0.02122071, 
    0.01857098, 0.009896323, 0.009670869, 0.003673331, 0.002994946, 
    0.0002998868, 0.004942393, 0.03211165, 0.03046639, 0.01497618, 
    0.01546751, 0.001080645, 0,
  0.06264501, 0.0533522, 0.04171479, 0.0299146, 0.001044079, 0.001490151, 
    0.009934915, -6.678737e-05, -0.0003668903, 0.001170285, 0.001017013, 
    -0.0001484926, 0.002024692, 0.05723718, 0.07004614, 0.08962317, 
    0.0862804, 0.1333763, 0.178808, 0.1874584, 0.1926491, 0.2191246, 
    0.2012515, 0.1363055, 0.1159142, 0.04477817, 0.04203179, 0.03275643, 
    0.04657942,
  0.147361, 0.1172936, 0.1178501, 0.1945998, 0.1657613, 0.1341173, 0.1232733, 
    0.1656489, 0.1601983, 0.1759015, 0.1706179, 0.2154824, 0.2096363, 
    0.2038621, 0.2209036, 0.2303881, 0.1977276, 0.180648, 0.2317895, 
    0.1756231, 0.2135032, 0.1865748, 0.2283787, 0.227777, 0.1753392, 
    0.1691317, 0.1528371, 0.1171619, 0.1217809,
  0.1915427, 0.1941065, 0.183383, 0.1512086, 0.1497383, 0.1906848, 0.1551038, 
    0.1648898, 0.1558124, 0.1676433, 0.2003044, 0.1991932, 0.1588029, 
    0.1538804, 0.1137107, 0.1342587, 0.1404455, 0.1481557, 0.1400958, 
    0.1525279, 0.2170585, 0.1897678, 0.1563607, 0.1420485, 0.1406615, 
    0.1584337, 0.1544335, 0.1786631, 0.1907847,
  0.07392301, 0.06986196, 0.04745378, 0.08913673, 0.1054261, 0.07352061, 
    0.08521464, 0.08104865, 0.08020435, 0.1083763, 0.1302977, 0.1242702, 
    0.05665772, 0.06071676, 0.08625703, 0.0910739, 0.143126, 0.1394105, 
    0.1128194, 0.1567669, 0.1781682, 0.08642849, 0.1473666, 0.1163116, 
    0.1215098, 0.1434291, 0.125033, 0.1514136, 0.1738485,
  0.00604359, 0.006509861, 0.02893814, 0.02834137, 0.05605591, 0.08565486, 
    0.08453768, 0.05558564, 0.05694322, 0.07519434, 0.1347339, 0.05815463, 
    0.02660124, 0.03099381, 0.04286162, 0.1008832, 0.0888536, 0.06883398, 
    0.1007323, 0.1104169, 0.09601544, 0.02150603, 0.02559055, 0.004780301, 
    0.02125115, 0.06612302, 0.09132934, 0.0615916, 0.01992583,
  4.560307e-07, 0.0005118316, 0.00235123, 0.008257467, 0.03157962, 
    0.08401671, 0.0590074, 0.02006578, 0.05007198, 0.02984052, 0.0007133812, 
    0.005190938, 0.03244923, 0.0436708, 0.09473786, 0.05529093, 0.02555402, 
    0.0453197, 0.07017893, 0.02051804, 9.393822e-05, 0.0003717796, 
    1.095206e-06, 0.02627485, 0.02533991, 0.03438878, 0.007118704, 
    0.00168627, 2.258934e-06,
  1.015237e-06, 0.1427293, 0.1071722, 0.0517398, 0.03628505, 0.03441193, 
    0.05787724, 0.03811539, 0.09923919, 0.02377382, 0.09304416, 0.05622818, 
    0.08270863, 0.05108462, 0.07281131, 0.0567397, 0.02296424, 0.01984535, 
    0.004504278, 0.001263143, 0.0005787399, 0.000112362, 0.001794289, 
    0.07814564, 0.07814102, 0.01124257, 0.02121237, 0.001929344, 7.237001e-06,
  0.04991298, 0.1550516, 0.09035733, 0.006187302, 0.01609192, 0.004504597, 
    0.004906977, 0.01119859, 0.05331419, 0.1449642, 0.0469466, 0.01540944, 
    0.05686032, 0.09581847, 0.05463677, 0.006457481, 0.005311701, 0.01876083, 
    0.01379095, 0.0007249002, 0.009994456, 0.008227451, 0.0884825, 0.1811594, 
    0.1266077, 0.07746987, 0.0567314, 0.01903934, 0.02842703,
  0.01762753, 0.002187497, 0.004403378, 0.01954961, 0.01683377, 0.003172865, 
    0.01232899, 0.006024901, 0.006363265, 0.04447554, 0.01239278, 0.05883819, 
    0.05828132, 0.08845741, 0.0542773, 0.09570953, 0.05758395, 0.04036679, 
    0.009629056, 0.02002806, 0.06880246, 0.01161835, 0.001978421, 0.02442846, 
    0.02919203, 0.01848807, 0.000883884, 0.006147352, 0.08058494,
  0.09026122, 0.01880755, 0.005353899, 0.02271803, 0.03770985, 0.01366701, 
    0.00254253, 0.0006857743, 0.01182908, 0.01130513, 0.01444722, 0.01550712, 
    0.01509792, 0.003217464, 0.005168006, 0.001291217, 0.003155732, 
    0.01447356, 0.04059307, 0.03700523, 0.06864214, 0.03870966, 0.006480374, 
    0.02753627, 0.01443474, 0.03147641, 0.01839051, 0.02557305, 0.04924968,
  0.05462993, 0.07029371, 0.06052553, 0.06676614, 0.09471866, 0.06527039, 
    0.04763424, 0.008036551, 0.1192834, 0.1399367, 0.1364649, 0.147137, 
    0.1390503, 0.08336426, 0.06839354, 0.04641974, 0.02537177, 0.02659982, 
    0.0276732, 0.02389744, 0.04507356, 0.06524418, 0.08900806, 0.08616528, 
    0.066083, 0.1215757, 0.09747914, 0.03035351, 0.03674355,
  0.09630399, 0.1091135, 0.1436574, 0.1420737, 0.1209893, 0.0947703, 
    0.1222868, 0.1867099, 0.1557532, 0.09424677, 0.08978642, 0.1335088, 
    0.1422086, 0.1891195, 0.2371178, 0.2093754, 0.1597575, 0.1474288, 
    0.1077091, 0.1225748, 0.1146734, 0.1098919, 0.1186731, 0.1389685, 
    0.1464037, 0.1386976, 0.1460648, 0.06237854, 0.06922226,
  0.2055931, 0.1797287, 0.1444894, 0.1194623, 0.1301486, 0.1074644, 
    0.1012327, 0.01591312, 0.01232462, 0.04780301, 0.07426674, 0.08215318, 
    0.122716, 0.1214065, 0.141434, 0.1055565, 0.1665681, 0.233987, 0.2432147, 
    0.1703439, 0.1231882, 0.1373897, 0.1511374, 0.1747563, 0.1926205, 
    0.1613468, 0.1436741, 0.1014241, 0.1590371,
  0.2227105, 0.1714897, 0.1677062, 0.1343946, 0.1246499, 0.08961365, 
    0.08090229, 0.06925857, 0.05933177, 0.01631577, 0.01584076, 
    -6.915566e-05, 0.04589308, 0.05827471, 0.06950798, 0.07730086, 
    0.07005107, 0.1361289, 0.1039749, 0.10221, 0.1111712, 0.1272816, 
    0.1342229, 0.1338461, 0.2152639, 0.09799911, 0.06614934, 0.1132504, 
    0.1767893,
  0.1639358, 0.1653327, 0.1773642, 0.1300159, 0.1674785, 0.1413794, 
    0.06695141, 0.08493104, 0.06082547, 0.04300062, 0.01021939, 0.01035272, 
    0.03845161, 0.07212491, 0.08112942, 0.0606854, 0.07380569, 0.05561364, 
    0.04210924, 0.07011426, 0.08102567, 0.06105822, 0.0537723, 0.04015902, 
    0.1340569, 0.01574755, -7.328047e-05, 0.09713854, 0.13412,
  0.06248057, 0.07769383, 0.1082805, 0.0998805, 0.09649432, 0.09888108, 
    0.1184639, 0.1120967, 0.07052199, 0.06197049, 0.08431464, 0.06820899, 
    0.04389339, 0.02972196, 0.02547684, 0.01870726, 0.02043249, 0.02290116, 
    0.03905036, 0.05193119, 0.05234461, 0.05313953, 0.03019056, 0.02506134, 
    0.02904884, 0.00482311, -0.003205588, 0.01600334, 0.04341492,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01191304, 0.0259208, 0.02430086, 
    0.03768728, 0.0337596, 0.023138, 0.007443589, 0.00569238, 0.005331785, 
    0.02811147, 0.1381095, 0.1195234, 0.05110437, 0.04251039, 0.007950957, 
    0.0001562846,
  0.1794532, 0.1267202, 0.1433663, 0.08454606, 0.003868261, 0.00149479, 
    0.03583848, 0.0003503035, -0.0003700477, 0.01113058, 0.0008858676, 
    -0.0004508667, 0.02453183, 0.1483112, 0.1816982, 0.1737126, 0.1655278, 
    0.2043335, 0.2366275, 0.2402484, 0.2531022, 0.2902297, 0.3281568, 
    0.2057832, 0.1942889, 0.1161914, 0.1517503, 0.1462123, 0.09334894,
  0.2028355, 0.1761859, 0.1957912, 0.2551039, 0.2224767, 0.1900777, 0.178577, 
    0.2266521, 0.2113857, 0.220673, 0.1994037, 0.2528347, 0.2475036, 
    0.2270755, 0.2459572, 0.2267856, 0.203957, 0.1745675, 0.2326533, 
    0.197434, 0.2334378, 0.2222205, 0.265624, 0.245532, 0.2329603, 0.2227422, 
    0.2087625, 0.204095, 0.226363,
  0.1853929, 0.1913608, 0.190743, 0.1549421, 0.1538882, 0.1898672, 0.1613584, 
    0.1646726, 0.1597736, 0.1873634, 0.200609, 0.1803232, 0.1516731, 
    0.1585204, 0.1103717, 0.1164256, 0.1342998, 0.1523173, 0.1573637, 
    0.1620261, 0.2053477, 0.1790717, 0.1379123, 0.1508059, 0.1727419, 
    0.1921697, 0.172442, 0.1782356, 0.1852859,
  0.0753877, 0.07059842, 0.04773027, 0.08478278, 0.09731118, 0.06749141, 
    0.09454702, 0.08070512, 0.06490651, 0.1015537, 0.1144081, 0.1100832, 
    0.05465555, 0.0537043, 0.08227703, 0.1066625, 0.1323425, 0.1329862, 
    0.1085521, 0.1459383, 0.1795305, 0.08438626, 0.1420284, 0.1236993, 
    0.09081821, 0.1214425, 0.1166932, 0.1393757, 0.1733112,
  0.001412934, 0.007381712, 0.0214879, 0.02594772, 0.05223439, 0.07831232, 
    0.05959557, 0.0403199, 0.02818189, 0.06625742, 0.1288256, 0.053529, 
    0.01874709, 0.03053075, 0.03626361, 0.1016419, 0.08113272, 0.0620488, 
    0.09626447, 0.09271816, 0.09931746, 0.02036254, 0.01392473, 0.004255779, 
    0.02433618, 0.06190063, 0.07704747, 0.05065738, 0.01813832,
  8.820088e-08, 0.0005032018, 0.001400115, 0.006471158, 0.02614954, 
    0.08226674, 0.05891315, 0.01838907, 0.04050619, 0.01976077, 0.0005752592, 
    0.003784551, 0.04265108, 0.0393081, 0.07700066, 0.04779934, 0.01729081, 
    0.04794904, 0.06300861, 0.01455721, 3.106542e-05, 7.079753e-06, 
    2.452214e-07, 0.01342264, 0.0184337, 0.02790372, 0.004952532, 
    0.0001939562, 1.327486e-06,
  6.316259e-06, 0.1484035, 0.09689488, 0.05587273, 0.02682639, 0.03191535, 
    0.05646566, 0.03968893, 0.09554051, 0.01964713, 0.09806854, 0.05143955, 
    0.08902144, 0.04976829, 0.0664374, 0.04668009, 0.02399662, 0.01892903, 
    0.005870939, 0.0009316691, 0.0004210209, -5.394904e-06, 0.0003339573, 
    0.05511404, 0.07802915, 0.008208965, 0.02222705, 0.001252558, 5.493694e-06,
  0.05051984, 0.1358739, 0.06942337, 0.008746636, 0.01583161, 0.004454703, 
    0.005583511, 0.009382496, 0.04155534, 0.1481495, 0.05534722, 0.01127348, 
    0.05098535, 0.08535676, 0.05138487, 0.00936807, 0.005139321, 0.01073815, 
    0.01856885, 0.0008282835, 0.01915754, 0.0153883, 0.1070383, 0.1887693, 
    0.1337131, 0.0896834, 0.06473929, 0.02248257, 0.02153698,
  0.01760959, 0.003956771, 0.003716623, 0.02089347, 0.009829692, 0.002780032, 
    0.01004421, 0.003844508, 0.004659242, 0.04181068, 0.01102643, 0.05521714, 
    0.05098286, 0.0854294, 0.0621382, 0.07488362, 0.05644552, 0.03160151, 
    0.006405292, 0.02066652, 0.06312749, 0.007988526, 0.001968179, 
    0.02297053, 0.02580962, 0.01958475, -5.791515e-05, 0.02251494, 0.06524374,
  0.0884003, 0.01018638, 0.004536764, 0.01873518, 0.03138182, 0.006138747, 
    0.001006657, 0.0003974352, 0.006416757, 0.01080347, 0.01525581, 0.01633, 
    0.01187175, 0.003715277, 0.0007374624, 0.001205795, 0.0007131937, 
    0.01027091, 0.03370555, 0.02747745, 0.04108326, 0.03706156, 0.003298339, 
    0.02749512, 0.006026695, 0.01785681, 0.01227159, 0.01425519, 0.0257808,
  0.04729435, 0.0728384, 0.06255461, 0.05972448, 0.09046534, 0.05311921, 
    0.04587662, 0.02002887, 0.1434383, 0.1356495, 0.135824, 0.1344238, 
    0.1345662, 0.1024037, 0.05842719, 0.02667213, 0.01325537, 0.02944051, 
    0.01759158, 0.01803249, 0.03338715, 0.05730851, 0.07752035, 0.07013693, 
    0.05688075, 0.1074235, 0.07198876, 0.02324892, 0.0216941,
  0.08744211, 0.1120404, 0.1408466, 0.1328576, 0.1078215, 0.08919664, 
    0.1677871, 0.1566289, 0.1383158, 0.08552975, 0.08998784, 0.1357139, 
    0.1380514, 0.1797266, 0.2345376, 0.2008936, 0.1601785, 0.126511, 
    0.0909203, 0.1166967, 0.1457611, 0.1067331, 0.1195937, 0.1496289, 
    0.1352924, 0.1257562, 0.1321068, 0.05816123, 0.06630151,
  0.1942708, 0.1785276, 0.1389944, 0.1144541, 0.1216778, 0.1044272, 
    0.1281922, 0.05005801, 0.05040938, 0.1228335, 0.1459886, 0.1318815, 
    0.1615331, 0.1490315, 0.1629756, 0.1507705, 0.1957176, 0.2492124, 
    0.2356859, 0.1623803, 0.1221173, 0.1533664, 0.1587679, 0.186511, 
    0.2064682, 0.169986, 0.1363755, 0.1059868, 0.1618138,
  0.2442579, 0.1871634, 0.1772564, 0.2052319, 0.1517936, 0.1049039, 
    0.1083845, 0.1114481, 0.1369417, 0.08634447, 0.07046919, 0.01798973, 
    0.1229244, 0.1469582, 0.09200673, 0.1498706, 0.1309571, 0.1992339, 
    0.133487, 0.1047342, 0.1517415, 0.1748021, 0.1408252, 0.1460077, 
    0.2062775, 0.117355, 0.05731087, 0.1405781, 0.2115976,
  0.2251885, 0.2014603, 0.2251586, 0.1837582, 0.1741109, 0.1480675, 
    0.09282047, 0.1024718, 0.106075, 0.1853222, 0.07562106, 0.08302065, 
    0.1113666, 0.1239557, 0.1051731, 0.1076732, 0.1058803, 0.08606905, 
    0.07362488, 0.09874857, 0.126142, 0.1201049, 0.11286, 0.07615338, 
    0.1476969, 0.03106391, 0.002084729, 0.1510822, 0.1850708,
  0.1442125, 0.1512422, 0.1727231, 0.1790615, 0.1470163, 0.143863, 0.1656134, 
    0.1637618, 0.1035186, 0.1095928, 0.1159378, 0.1070548, 0.09434588, 
    0.09272063, 0.0930253, 0.06039176, 0.03827733, 0.068284, 0.08550915, 
    0.08515111, 0.08970115, 0.09765918, 0.06361265, 0.0313556, 0.04646282, 
    0.021076, 0.01331808, 0.03599501, 0.1331837,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.096444e-05, -1.096444e-05, 
    -1.096444e-05, -1.096444e-05, -1.096444e-05, -1.096444e-05, 
    -1.096444e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.0003346974, -3.783066e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002260213, 
    0.02809409, 0.06327744, 0.07825123, 0.1315994, 0.09803841, 0.07199374, 
    0.02978557, 0.01531196, 0.01235399, 0.07212055, 0.2240907, 0.2604515, 
    0.1757418, 0.1416722, 0.0198518, 0.002538941,
  0.2540408, 0.2380491, 0.2213365, 0.171546, 0.01780067, 0.01741861, 
    0.09783198, 0.0033896, 0.01152071, 0.02880967, 0.01232987, -9.9133e-05, 
    0.06393904, 0.2108725, 0.2740555, 0.2797185, 0.254946, 0.2852367, 
    0.3159663, 0.3076881, 0.284219, 0.3370115, 0.3671569, 0.2776074, 
    0.266436, 0.1467583, 0.1724245, 0.1793868, 0.2490333,
  0.2583839, 0.2485156, 0.2616828, 0.2946774, 0.2615011, 0.2606839, 
    0.2156838, 0.3094924, 0.2787368, 0.2668339, 0.2498346, 0.2853563, 
    0.2577545, 0.2441358, 0.2499224, 0.2481003, 0.2069389, 0.1765452, 
    0.2292463, 0.2147068, 0.239638, 0.2325093, 0.2484802, 0.2479949, 
    0.2420052, 0.2127974, 0.2251261, 0.2308069, 0.2674501,
  0.1845143, 0.1949356, 0.1953021, 0.1636267, 0.1570446, 0.1893413, 
    0.1668432, 0.171472, 0.1668349, 0.2094103, 0.1940948, 0.1745652, 
    0.1557895, 0.1494371, 0.1077133, 0.1048063, 0.1317091, 0.1408585, 
    0.1574032, 0.1495865, 0.2012853, 0.2013655, 0.1384066, 0.1646858, 
    0.1606283, 0.2026977, 0.1785316, 0.1805312, 0.1946375,
  0.08521652, 0.05831763, 0.04688007, 0.08329935, 0.1012665, 0.0561469, 
    0.09352137, 0.06940982, 0.0674584, 0.09234327, 0.09062137, 0.08061466, 
    0.05004204, 0.05495515, 0.07884431, 0.1049517, 0.1201213, 0.1216351, 
    0.1129525, 0.1395032, 0.1671143, 0.07853112, 0.1475399, 0.1124618, 
    0.06849164, 0.1150023, 0.109612, 0.1322472, 0.1611873,
  0.0006444023, 0.009023872, 0.02148727, 0.02643385, 0.04957653, 0.06912486, 
    0.04038102, 0.02904807, 0.02177895, 0.06198014, 0.1154013, 0.04751451, 
    0.01382008, 0.03204492, 0.03091238, 0.0950368, 0.08107002, 0.06488637, 
    0.08906648, 0.0773869, 0.1035932, 0.02336928, 0.009579288, 0.005053564, 
    0.02882151, 0.05788364, 0.08167349, 0.05182242, 0.0187814,
  1.183391e-07, 0.0004825148, 0.0006236453, 0.005627806, 0.02307231, 
    0.07577849, 0.05852725, 0.02535876, 0.04179136, 0.0119463, 0.0005799719, 
    0.002286726, 0.0342846, 0.03751555, 0.07223398, 0.04173963, 0.02094342, 
    0.04957236, 0.05998163, 0.008627094, 2.030605e-05, 1.593628e-06, 
    2.126105e-07, 0.005930494, 0.01594462, 0.0220452, 0.007023104, 
    9.498568e-05, 4.57498e-07,
  0.000185031, 0.1510306, 0.0968577, 0.05415532, 0.02827093, 0.03013316, 
    0.05948886, 0.03819413, 0.093715, 0.01880352, 0.09354715, 0.0639736, 
    0.09440211, 0.05062786, 0.06527077, 0.03459153, 0.02463581, 0.01924207, 
    0.00551175, 0.000815084, 0.0007276622, 0.00013837, 0.001518616, 
    0.0424388, 0.08293712, 0.006346278, 0.02753261, 0.0009896404, 5.36042e-06,
  0.0547093, 0.1276768, 0.06300341, 0.00942328, 0.01212113, 0.003819967, 
    0.004356735, 0.00872768, 0.0381292, 0.1470779, 0.06481138, 0.008932781, 
    0.05071465, 0.07826566, 0.04859421, 0.00786235, 0.003678339, 0.005124855, 
    0.01863083, 0.000501555, 0.02126159, 0.01528677, 0.1287322, 0.1875395, 
    0.1214241, 0.07983651, 0.05949653, 0.03098387, 0.02728432,
  0.01754134, 0.00420678, 0.002765466, 0.03802163, 0.005815728, 0.00291491, 
    0.009863924, 0.002942377, 0.003742598, 0.03992142, 0.009820726, 
    0.04565619, 0.04755306, 0.08789054, 0.06837154, 0.06613585, 0.05595759, 
    0.02897487, 0.003869331, 0.02392757, 0.05651794, 0.005567217, 
    0.001619606, 0.0190861, 0.02173081, 0.01113672, -0.0001413653, 
    0.03308176, 0.04410895,
  0.08313593, 0.008264306, 0.008895178, 0.01199021, 0.03129822, 0.003178521, 
    0.0007261435, 0.0003158655, 0.00468875, 0.009356857, 0.01591916, 
    0.01719073, 0.009245457, 0.002884207, 0.0005284009, 0.001241736, 
    0.0004689361, 0.008413762, 0.02571521, 0.01605592, 0.01371599, 
    0.03786987, 0.001461369, 0.02614868, 0.003780055, 0.01737173, 
    0.009942113, 0.006705661, 0.04499613,
  0.04143329, 0.07186038, 0.06546895, 0.06010019, 0.08636114, 0.04720809, 
    0.05902306, 0.02706833, 0.1476715, 0.1374771, 0.1373704, 0.1257467, 
    0.1240483, 0.1207651, 0.04338397, 0.02410132, 0.01134316, 0.03337998, 
    0.01413423, 0.01106783, 0.03071046, 0.05585998, 0.06292123, 0.05698982, 
    0.05140709, 0.09526485, 0.04864764, 0.01817194, 0.009979619,
  0.08008085, 0.1011661, 0.1465917, 0.1240505, 0.09622905, 0.07972929, 
    0.1890252, 0.1348411, 0.1215332, 0.06976325, 0.0922991, 0.1331867, 
    0.1293281, 0.1709252, 0.2272898, 0.1980015, 0.1544548, 0.1135581, 
    0.08731465, 0.1120838, 0.1342925, 0.1115955, 0.1218917, 0.1632055, 
    0.1277508, 0.1187845, 0.1136688, 0.05376449, 0.06281564,
  0.1954557, 0.1738084, 0.1403505, 0.1141711, 0.1153222, 0.1083302, 
    0.1528748, 0.1292902, 0.105382, 0.2133761, 0.1911142, 0.1539076, 
    0.1766144, 0.1741481, 0.1585991, 0.1598206, 0.1990005, 0.2428463, 
    0.2136784, 0.1562236, 0.1332973, 0.1623312, 0.1659666, 0.1969075, 
    0.2261064, 0.1683196, 0.133963, 0.1145174, 0.1616211,
  0.2682607, 0.2074453, 0.1725238, 0.215997, 0.1644355, 0.1175469, 0.1574244, 
    0.1443601, 0.2070163, 0.1227934, 0.09256095, 0.06619769, 0.1491783, 
    0.2277172, 0.1239612, 0.1998023, 0.2268696, 0.2607796, 0.1632559, 
    0.1094802, 0.168355, 0.2126571, 0.1539842, 0.1470128, 0.2232649, 
    0.137251, 0.05575629, 0.1539402, 0.2501236,
  0.2601913, 0.2125219, 0.2468197, 0.1944523, 0.1598106, 0.1285228, 
    0.09541175, 0.1111987, 0.1292606, 0.2129593, 0.1510885, 0.1548991, 
    0.1937892, 0.2005589, 0.159756, 0.1455653, 0.1263744, 0.1139227, 
    0.1293427, 0.1482235, 0.1788798, 0.1445988, 0.1515467, 0.1154282, 
    0.1754505, 0.04849176, 0.007079888, 0.2398523, 0.2240633,
  0.1954309, 0.1789135, 0.2077999, 0.2305996, 0.1624773, 0.1519415, 
    0.1698004, 0.1746125, 0.1238, 0.1262091, 0.1479474, 0.1414109, 0.1316346, 
    0.1369393, 0.1439735, 0.1156714, 0.09760914, 0.1043418, 0.08944105, 
    0.09449674, 0.115328, 0.138059, 0.1012343, 0.07004999, 0.0823832, 
    0.02678327, 0.01954934, 0.07026882, 0.2250776,
  2.192887e-05, 2.192887e-05, 2.192887e-05, 2.192887e-05, 2.192887e-05, 
    2.192887e-05, 2.192887e-05, -2.876495e-05, -1.158061e-05, 5.603743e-06, 
    2.278809e-05, 3.997244e-05, 5.715679e-05, 7.434114e-05, 0.0005197049, 
    0.0005368893, 0.0005540737, 0.000571258, 0.0005884424, 0.0006056267, 
    0.000622811, 0.000137064, 0.0001026953, 6.832662e-05, 3.395792e-05, 
    -4.107793e-07, -3.477948e-05, -6.914818e-05, 2.192887e-05,
  0.0002043859, -2.466005e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003447138, 
    0.07366336, 0.08133166, 0.1288966, 0.1989916, 0.2119056, 0.1623235, 
    0.1071496, 0.0625276, 0.04033706, 0.1560826, 0.2372879, 0.3058456, 
    0.3105704, 0.2850715, 0.07734647, 0.008106328,
  0.2460649, 0.2743218, 0.2556578, 0.277067, 0.05756614, 0.0488645, 0.146343, 
    0.03312634, 0.04427858, 0.0669299, 0.03206714, 0.006046943, 0.1170193, 
    0.2334532, 0.3331318, 0.3440423, 0.2972764, 0.3024658, 0.3557129, 
    0.329208, 0.3100041, 0.3530754, 0.3902583, 0.2898495, 0.2978574, 
    0.1744659, 0.2007923, 0.2216288, 0.2638292,
  0.2701944, 0.2597555, 0.2688015, 0.2919999, 0.2577023, 0.2738489, 
    0.2222667, 0.3154196, 0.3158779, 0.2863223, 0.2698482, 0.2884766, 
    0.2686422, 0.2577798, 0.2584707, 0.2540541, 0.2320626, 0.1845533, 
    0.2316589, 0.2175195, 0.2382848, 0.2365741, 0.249751, 0.2488115, 
    0.2525404, 0.2088698, 0.2194722, 0.2439668, 0.2721665,
  0.183818, 0.1995622, 0.2040845, 0.1652485, 0.1610961, 0.1954397, 0.1677115, 
    0.1746115, 0.1607777, 0.2025758, 0.1941311, 0.1761517, 0.1434447, 
    0.150136, 0.1182258, 0.0996284, 0.132026, 0.1443052, 0.1647205, 
    0.1602479, 0.1871337, 0.170093, 0.1406008, 0.151812, 0.1701116, 
    0.1834721, 0.1807536, 0.1771421, 0.1918097,
  0.08396593, 0.05649927, 0.04004416, 0.08209939, 0.08701484, 0.04804614, 
    0.08047035, 0.07855516, 0.0621876, 0.07777957, 0.08073828, 0.07246371, 
    0.05206279, 0.05821316, 0.07063093, 0.1079618, 0.1197544, 0.1180369, 
    0.1121416, 0.1427853, 0.1619366, 0.07339099, 0.1334976, 0.09649491, 
    0.04897686, 0.09398596, 0.1115301, 0.1242091, 0.1590616,
  7.16365e-05, 0.01130923, 0.02263312, 0.02515437, 0.05104425, 0.05823116, 
    0.03144495, 0.01993686, 0.02233511, 0.05876884, 0.1054542, 0.04170579, 
    0.01859128, 0.03057049, 0.0260212, 0.09435005, 0.08390208, 0.0652409, 
    0.08862324, 0.06700768, 0.0981689, 0.0215575, 0.009910946, 0.006009143, 
    0.02827678, 0.0551562, 0.07554123, 0.04723438, 0.01525822,
  1.355495e-07, 0.0006121445, 0.000710316, 0.005701544, 0.02090788, 
    0.06411944, 0.05760656, 0.02554017, 0.03892113, 0.007587296, 
    0.0005995082, 0.001128935, 0.02514393, 0.03266709, 0.07332585, 
    0.04578358, 0.02535631, 0.05341762, 0.04525992, 0.004564203, 
    7.367803e-05, 1.501607e-06, 5.789472e-08, 0.001515284, 0.01793489, 
    0.02020907, 0.01060207, 9.744073e-05, 4.043103e-07,
  -4.645863e-05, 0.1514244, 0.1024363, 0.05321861, 0.02934801, 0.03350552, 
    0.06312106, 0.04388947, 0.1023016, 0.02308549, 0.09538511, 0.07386501, 
    0.1013471, 0.05022455, 0.06071763, 0.03284062, 0.0286925, 0.02147007, 
    0.004494015, 0.001199294, 0.001081695, 0.001192727, 0.007832132, 
    0.04696532, 0.08953646, 0.004685021, 0.03146892, 0.0009598335, 
    1.759819e-06,
  0.06990576, 0.1263056, 0.07267793, 0.00695822, 0.008090561, 0.003835832, 
    0.004614649, 0.007084928, 0.03892899, 0.1516491, 0.05485408, 0.00867722, 
    0.05508872, 0.07832988, 0.0459446, 0.007626674, 0.004551466, 0.004345099, 
    0.01772663, 0.0006241308, 0.03043555, 0.01651247, 0.1434983, 0.1809809, 
    0.1265625, 0.07305236, 0.05418756, 0.03869911, 0.03999184,
  0.01359011, 0.01253137, 0.002518531, 0.06460941, 0.004007988, 0.004353402, 
    0.01280626, 0.002783803, 0.005127681, 0.04192148, 0.008847527, 
    0.04236897, 0.05010829, 0.1027999, 0.08564874, 0.06841879, 0.06571743, 
    0.02711478, 0.004430334, 0.03010146, 0.06673937, 0.005715915, 0.00298199, 
    0.01235754, 0.02087572, 0.005883973, -3.122601e-05, 0.03231198, 0.03758829,
  0.05928261, 0.007447827, 0.009665784, 0.006279644, 0.04354608, 0.001731369, 
    0.004597531, 0.0004188054, 0.004391592, 0.01050141, 0.01649242, 
    0.01862731, 0.01343743, 0.001427072, 0.0005832121, 0.001492211, 
    0.0007801372, 0.00952065, 0.01331769, 0.01222359, 0.005239033, 
    0.04006063, 0.001339577, 0.02600079, 0.001861142, 0.02419246, 
    0.003526056, 0.004681598, 0.05804715,
  0.03245427, 0.07107288, 0.05111217, 0.05854085, 0.08999948, 0.0438586, 
    0.08851482, 0.04686803, 0.1462035, 0.158177, 0.1428191, 0.1265616, 
    0.1242704, 0.1094001, 0.03996371, 0.01522301, 0.00917004, 0.03558106, 
    0.01026124, 0.006934992, 0.0242752, 0.04827382, 0.05038191, 0.05423829, 
    0.03947153, 0.08186503, 0.04546747, 0.01070361, 0.006295617,
  0.06874986, 0.09909964, 0.1418477, 0.1274025, 0.09171528, 0.07350355, 
    0.1953187, 0.1152605, 0.1064581, 0.06512916, 0.08943281, 0.1344552, 
    0.1285703, 0.1545228, 0.2144768, 0.1969178, 0.1510982, 0.1205336, 
    0.09278595, 0.1046965, 0.133542, 0.1170438, 0.1268812, 0.1538366, 
    0.1300764, 0.1047706, 0.09831758, 0.05116813, 0.06116753,
  0.1884331, 0.1696609, 0.1398483, 0.1117943, 0.1073261, 0.1174323, 
    0.1625584, 0.1660134, 0.1609892, 0.234753, 0.2038498, 0.1843017, 
    0.1929732, 0.1779583, 0.1601408, 0.1576092, 0.1966544, 0.2188746, 
    0.2022745, 0.1605877, 0.1418054, 0.1615002, 0.1697516, 0.2128494, 
    0.223879, 0.1686185, 0.1419897, 0.101231, 0.1485578,
  0.2656498, 0.2114825, 0.1678641, 0.2138272, 0.1625606, 0.1095191, 
    0.1689536, 0.1876382, 0.2493627, 0.2036809, 0.1139798, 0.1379108, 
    0.2124406, 0.2594819, 0.1227791, 0.2093598, 0.2365336, 0.2909404, 
    0.2093976, 0.1265514, 0.1726656, 0.2246279, 0.1801183, 0.1581806, 
    0.2252641, 0.1370715, 0.06029735, 0.1577768, 0.2589379,
  0.2623306, 0.2241749, 0.2368094, 0.18097, 0.1504656, 0.1061736, 0.09412422, 
    0.1100498, 0.1346731, 0.194764, 0.1764932, 0.197035, 0.2381753, 
    0.2348074, 0.1814899, 0.1475027, 0.1484106, 0.1347553, 0.1378044, 
    0.1729515, 0.2151125, 0.144231, 0.1449742, 0.1239127, 0.1736153, 
    0.06439683, 0.01530484, 0.285837, 0.2204624,
  0.2110286, 0.1969177, 0.2275402, 0.2305043, 0.1667879, 0.1521647, 
    0.1663861, 0.1791779, 0.1289806, 0.152114, 0.160068, 0.1521043, 0.154657, 
    0.1617772, 0.1810162, 0.1469155, 0.1160173, 0.1134018, 0.117832, 
    0.1086416, 0.1451661, 0.1723854, 0.1291625, 0.1064601, 0.1449854, 
    0.06416208, 0.03479393, 0.1508235, 0.2464748,
  9.921378e-05, 9.06216e-05, 8.202943e-05, 7.343725e-05, 6.484508e-05, 
    5.62529e-05, 4.766073e-05, 0.0002531708, 0.0004209437, 0.0005887166, 
    0.0007564895, 0.0009242624, 0.001092035, 0.001259808, -0.0006712595, 
    -0.0005750298, -0.0004788, -0.0003825703, -0.0002863406, -0.0001901108, 
    -9.388112e-05, 0.001034807, 0.0007793965, 0.0005239861, 0.0002685756, 
    1.31652e-05, -0.0002422452, -0.0004976557, 0.0001060875,
  0.006727635, -0.000117339, 0, 0, 0, -2.540824e-06, 0, 0, 0, 0, 0, 
    0.0001632059, 0.01042103, 0.1267566, 0.104087, 0.1473211, 0.2586132, 
    0.2570436, 0.248181, 0.1851567, 0.1536708, 0.118237, 0.2350541, 
    0.2418472, 0.2949623, 0.3439479, 0.3125547, 0.1911292, 0.02526144,
  0.2297846, 0.2830914, 0.2687707, 0.3162159, 0.1076629, 0.09593193, 
    0.1648603, 0.09111589, 0.0992077, 0.1221907, 0.06507688, 0.04092509, 
    0.1597013, 0.2313928, 0.339844, 0.3713329, 0.3094564, 0.3113105, 
    0.3796411, 0.3495128, 0.2959167, 0.3371464, 0.3761638, 0.2679521, 
    0.3182103, 0.1921387, 0.1897206, 0.2234311, 0.2728399,
  0.2808532, 0.2631096, 0.2801753, 0.3052995, 0.2604577, 0.2819159, 
    0.2351657, 0.3069566, 0.3283792, 0.2966009, 0.2686617, 0.2861325, 
    0.2616925, 0.2654343, 0.2604983, 0.2321209, 0.2507544, 0.2039324, 
    0.2397448, 0.2180005, 0.2272151, 0.226271, 0.2408473, 0.2372195, 
    0.2443419, 0.1967971, 0.2187627, 0.2398797, 0.2684063,
  0.1996152, 0.1960452, 0.206686, 0.1402461, 0.1546203, 0.1981183, 0.1664742, 
    0.1798586, 0.150261, 0.2104478, 0.1878212, 0.1723799, 0.1338294, 
    0.1456074, 0.12034, 0.08681969, 0.1269259, 0.1396306, 0.1789171, 
    0.1487364, 0.1888721, 0.1838278, 0.1570187, 0.1447924, 0.152046, 
    0.2185407, 0.1691732, 0.1709886, 0.1931774,
  0.0774501, 0.05934801, 0.04353728, 0.07668142, 0.08262444, 0.05410313, 
    0.07931954, 0.07089768, 0.06647127, 0.07720359, 0.06812117, 0.07279266, 
    0.04827734, 0.05725884, 0.06461421, 0.1075606, 0.1222856, 0.104823, 
    0.1169309, 0.1364148, 0.1611936, 0.06981608, 0.1151287, 0.09175052, 
    0.03708774, 0.08253309, 0.1030667, 0.1183401, 0.1495997,
  0.001576251, 0.01515474, 0.02754234, 0.02702105, 0.04904188, 0.05714357, 
    0.03096718, 0.01542582, 0.02277165, 0.05405692, 0.1039067, 0.03676419, 
    0.02280759, 0.03001383, 0.02477489, 0.08940643, 0.08392002, 0.06767218, 
    0.08720532, 0.06176332, 0.1032709, 0.02003936, 0.01104299, 0.00536739, 
    0.03070979, 0.05744098, 0.07853141, 0.04993427, 0.01333632,
  6.175727e-07, 0.0006990134, 0.0009250302, 0.007346516, 0.02474846, 
    0.06320844, 0.06545554, 0.04426544, 0.04249287, 0.01684596, 0.0007319259, 
    0.001201127, 0.02143171, 0.02661271, 0.07187086, 0.05082863, 0.03551246, 
    0.06583744, 0.04247664, 0.004407166, 4.464787e-05, 3.246382e-06, 
    1.3228e-07, 0.001524724, 0.02345029, 0.02829934, 0.01277403, 
    0.0001734603, 1.432886e-06,
  4.690228e-05, 0.1590868, 0.1083253, 0.06546889, 0.03467081, 0.05451209, 
    0.07898498, 0.06170987, 0.1184113, 0.02823713, 0.1003288, 0.09553145, 
    0.1184925, 0.06229146, 0.06924437, 0.03871447, 0.03738243, 0.02820475, 
    0.004465138, 0.001527019, 0.001701305, 0.003689824, 0.003454243, 
    0.06812783, 0.1083989, 0.006084238, 0.03984424, 0.001797836, 2.593543e-06,
  0.1003787, 0.1485693, 0.1002978, 0.006754423, 0.01157764, 0.004292886, 
    0.005250487, 0.008983038, 0.04560917, 0.157755, 0.0626149, 0.01066681, 
    0.0807744, 0.08944479, 0.05270219, 0.0077637, 0.006985914, 0.005806302, 
    0.01577465, 0.002284132, 0.03520939, 0.01969466, 0.1302898, 0.2082771, 
    0.147246, 0.07369231, 0.05998465, 0.05135459, 0.05409759,
  0.01694657, 0.04264613, 0.01157752, 0.1092942, 0.004096012, 0.006352468, 
    0.0211601, 0.004283464, 0.009724637, 0.04524115, 0.01252019, 0.05093543, 
    0.05945509, 0.1176306, 0.09691941, 0.0783367, 0.07652275, 0.02432553, 
    0.01090529, 0.03523917, 0.07830672, 0.006955805, 0.005787546, 0.01327154, 
    0.0206956, 0.003504584, 0.0001524936, 0.03887243, 0.05268923,
  0.01438101, 0.00580591, 0.01160317, 0.004115872, 0.07935126, 0.002788585, 
    0.009126715, 0.0009455996, 0.009262821, 0.01467456, 0.01587767, 
    0.02137177, 0.01838964, 0.0009652683, 0.0007906526, 0.001504336, 
    0.002117581, 0.01056712, 0.002969126, 0.01194331, 0.003813798, 
    0.03910881, 0.001945614, 0.02771002, 0.002514239, 0.0381271, 0.003205541, 
    0.0008836601, 0.06871658,
  0.01895533, 0.0561466, 0.02823836, 0.03999155, 0.09478937, 0.0424881, 
    0.09744526, 0.0509186, 0.1515263, 0.175783, 0.152624, 0.1167355, 
    0.1271753, 0.1017476, 0.04607622, 0.01522048, 0.006872488, 0.04314451, 
    0.01001292, 0.004696024, 0.02413154, 0.03727296, 0.03902793, 0.04422026, 
    0.03876562, 0.07096307, 0.04280065, 0.00943303, 0.004217623,
  0.06214939, 0.08270784, 0.1377935, 0.1252333, 0.09339556, 0.06379841, 
    0.1865521, 0.0956488, 0.08663264, 0.07012736, 0.08778021, 0.1300222, 
    0.124653, 0.1429902, 0.1918473, 0.1854266, 0.1454904, 0.1132188, 
    0.09380431, 0.09193991, 0.137471, 0.1142876, 0.1312262, 0.1591546, 
    0.1263295, 0.1043154, 0.08633927, 0.04657266, 0.07093016,
  0.1726877, 0.1778946, 0.1369674, 0.1083091, 0.1069747, 0.1277608, 
    0.1625555, 0.1795114, 0.2201058, 0.234784, 0.2107894, 0.2046517, 
    0.2066587, 0.1678569, 0.1697957, 0.1504532, 0.1943991, 0.1942043, 
    0.1879123, 0.1670711, 0.1463736, 0.1535211, 0.1685914, 0.2085385, 
    0.2268518, 0.1894678, 0.1246327, 0.1111729, 0.1478324,
  0.2467926, 0.2091174, 0.1588794, 0.2099865, 0.1506967, 0.1110791, 
    0.1547662, 0.1896478, 0.2637881, 0.2060051, 0.1525421, 0.1603172, 
    0.262864, 0.2583395, 0.1203924, 0.2108192, 0.2200091, 0.2993516, 
    0.2121009, 0.1231211, 0.164854, 0.2228623, 0.1811887, 0.1829178, 
    0.2384097, 0.1371712, 0.07166889, 0.1561071, 0.2480898,
  0.2443988, 0.2123123, 0.2322265, 0.1691248, 0.1526325, 0.09199128, 
    0.08190142, 0.1131332, 0.1310377, 0.1786043, 0.1874302, 0.1898398, 
    0.2303647, 0.2483903, 0.1746599, 0.147128, 0.1662759, 0.1343243, 
    0.1407901, 0.1491801, 0.2022479, 0.1436605, 0.1420587, 0.1277449, 
    0.161868, 0.1151755, 0.03593816, 0.299848, 0.2094643,
  0.2094988, 0.2007561, 0.2297158, 0.2264626, 0.1748111, 0.1487163, 
    0.1654935, 0.1888487, 0.1273224, 0.1519255, 0.1519962, 0.1373216, 
    0.1432184, 0.1491218, 0.1772418, 0.1523864, 0.1223177, 0.1044399, 
    0.1114478, 0.1515371, 0.2036356, 0.1955558, 0.1404632, 0.1392381, 
    0.1878095, 0.1062498, 0.1045005, 0.1544281, 0.2538508,
  0.006284607, 0.005720255, 0.005155902, 0.00459155, 0.004027198, 
    0.003462845, 0.002898493, 0.005027459, 0.006589411, 0.008151364, 
    0.009713315, 0.01127527, 0.01283722, 0.01439917, 0.01723035, 0.01766137, 
    0.01809239, 0.01852342, 0.01895444, 0.01938546, 0.01981648, 0.0185674, 
    0.01713878, 0.01571016, 0.01428154, 0.01285292, 0.01142429, 0.009995673, 
    0.006736089,
  0.01917782, 0.003672518, -3.979388e-05, 0, 0, -8.790036e-05, 1.992415e-05, 
    0, 0, 0, 0.0003070039, 0.01745338, 0.02368032, 0.1748005, 0.1085648, 
    0.1538337, 0.2719971, 0.292114, 0.2898681, 0.3185978, 0.2713538, 
    0.2607662, 0.313209, 0.2411192, 0.2943572, 0.3365193, 0.3216108, 
    0.2542859, 0.07849836,
  0.2324735, 0.2929329, 0.2773668, 0.3334781, 0.1805013, 0.1303448, 
    0.1989191, 0.165773, 0.1615093, 0.1802759, 0.1263233, 0.0724512, 
    0.1605769, 0.2302051, 0.3425795, 0.3885691, 0.3073368, 0.3246258, 
    0.3979982, 0.3696103, 0.354209, 0.3447829, 0.3861431, 0.2804987, 
    0.3173153, 0.2234527, 0.1907559, 0.2450311, 0.2773283,
  0.3033383, 0.2578235, 0.2624807, 0.3026198, 0.2476914, 0.2728564, 
    0.2334411, 0.3263401, 0.3351232, 0.3221265, 0.3059223, 0.2774131, 
    0.2494579, 0.270229, 0.2775643, 0.2486497, 0.2547979, 0.2044048, 
    0.2341532, 0.2030248, 0.2154514, 0.2088037, 0.2292784, 0.2541261, 
    0.2373404, 0.2379722, 0.2301628, 0.2433479, 0.2734104,
  0.1804079, 0.1933587, 0.2181508, 0.1410078, 0.1603535, 0.1878279, 
    0.1597239, 0.1660337, 0.1619532, 0.2051983, 0.1957588, 0.1804417, 
    0.1270933, 0.1518818, 0.1157864, 0.07840723, 0.1292406, 0.1538188, 
    0.1750753, 0.1508593, 0.1791328, 0.1637668, 0.1609581, 0.1294813, 
    0.1606718, 0.1948613, 0.1761669, 0.1718909, 0.1915836,
  0.07103414, 0.06356416, 0.04142244, 0.0836046, 0.08868091, 0.06226651, 
    0.08199122, 0.06982771, 0.06851238, 0.07821326, 0.0622751, 0.08972748, 
    0.05923304, 0.05683085, 0.06902294, 0.1097393, 0.1238257, 0.1015299, 
    0.1256527, 0.135199, 0.1685434, 0.07096312, 0.1034274, 0.09128875, 
    0.03756656, 0.06779718, 0.1029042, 0.1126996, 0.149699,
  0.003024023, 0.01950374, 0.03791222, 0.02512247, 0.06356474, 0.05744803, 
    0.03520054, 0.02030759, 0.02496242, 0.05037206, 0.1266665, 0.04003101, 
    0.02722433, 0.02904703, 0.02739315, 0.08540414, 0.0907896, 0.07051335, 
    0.07879676, 0.07554427, 0.1257238, 0.02286335, 0.01340777, 0.005103817, 
    0.04332046, 0.06082086, 0.08540145, 0.05639758, 0.01356124,
  9.990032e-07, 0.003449986, 0.0009902272, 0.01172025, 0.02904207, 
    0.06606544, 0.073142, 0.04341467, 0.05342397, 0.02377099, 0.001397353, 
    0.002195216, 0.0257456, 0.01995946, 0.07140721, 0.05766857, 0.04690973, 
    0.0860706, 0.04420126, 0.004490868, 0.0001192414, -1.606388e-06, 
    1.454803e-07, 0.001135943, 0.02318247, 0.01751815, 0.01237626, 
    0.0003785384, 2.126093e-06,
  5.944245e-05, 0.1582806, 0.1234737, 0.08596457, 0.04296947, 0.06281216, 
    0.09662598, 0.06564049, 0.129657, 0.03673616, 0.102995, 0.111206, 
    0.124167, 0.06595585, 0.0709203, 0.04745866, 0.03899073, 0.03507579, 
    0.005239401, 0.001189255, 0.001798465, 0.003692271, 0.00766877, 
    0.09666918, 0.1297077, 0.007807603, 0.04308006, 0.002174851, 6.387651e-05,
  0.1124916, 0.1908408, 0.124757, 0.01056144, 0.01252947, 0.003313827, 
    0.003758963, 0.009139054, 0.06068992, 0.1954879, 0.07562679, 0.01331465, 
    0.09293711, 0.100501, 0.05603648, 0.007315585, 0.007689543, 0.005964666, 
    0.01393368, 0.008555377, 0.02803868, 0.02657158, 0.1466346, 0.2375828, 
    0.1819625, 0.07546998, 0.07142062, 0.0582064, 0.0714341,
  0.03290749, 0.03180472, 0.02161933, 0.161313, 0.004824988, 0.007521727, 
    0.03003937, 0.005502551, 0.01088766, 0.04441431, 0.01510861, 0.05144829, 
    0.06271221, 0.1233237, 0.1063222, 0.0902083, 0.08641201, 0.0224315, 
    0.0152541, 0.04388159, 0.09294368, 0.007107044, 0.009708505, 0.01704327, 
    0.02046672, 0.001960801, 0.0009098965, 0.02686457, 0.0805895,
  0.00486264, 0.002286479, 0.008592417, 0.004633677, 0.09496842, 0.002631139, 
    0.01715078, 0.001072529, 0.03303741, 0.01268936, 0.0156677, 0.02150199, 
    0.01988323, 0.0012311, 0.001603112, 0.001331683, 0.005689697, 
    0.006180707, 0.0004964492, 0.005868134, 0.00137857, 0.03878603, 
    0.003613914, 0.03256893, 0.006786454, 0.04595076, 0.008713699, 
    0.002693088, 0.0450907,
  0.009404606, 0.03818416, 0.01970898, 0.02409263, 0.09468669, 0.03921153, 
    0.07234413, 0.05119465, 0.1489938, 0.1967577, 0.1575265, 0.1204144, 
    0.1425599, 0.0947405, 0.06037467, 0.01409674, 0.005608932, 0.04243428, 
    0.01219273, 0.007984535, 0.02586663, 0.03330327, 0.02981826, 0.03993848, 
    0.04278824, 0.06296089, 0.03493862, 0.01365458, 0.001897713,
  0.05656459, 0.06228646, 0.1291282, 0.1180654, 0.09892295, 0.06042905, 
    0.1745628, 0.07656061, 0.06196354, 0.07007489, 0.08486561, 0.1296593, 
    0.1221473, 0.1335567, 0.1786454, 0.1790207, 0.1476884, 0.1118104, 
    0.1064591, 0.0912827, 0.1398343, 0.10606, 0.1345701, 0.1651612, 
    0.1263537, 0.1064749, 0.09601969, 0.04525626, 0.06734417,
  0.171136, 0.168595, 0.135121, 0.1018756, 0.1071305, 0.1257342, 0.1556538, 
    0.2028755, 0.2323446, 0.2287253, 0.2169488, 0.2063684, 0.2119766, 
    0.1706746, 0.1892725, 0.1558132, 0.1840803, 0.1931224, 0.1934337, 
    0.1667345, 0.1437579, 0.1579426, 0.1614936, 0.2258947, 0.2312344, 
    0.1860769, 0.1211783, 0.1036538, 0.148676,
  0.2405097, 0.204911, 0.1408449, 0.1859718, 0.1399999, 0.1168634, 0.1566607, 
    0.1994648, 0.2713776, 0.1967818, 0.1663622, 0.1594895, 0.2689843, 
    0.2571193, 0.1207278, 0.2105383, 0.2190897, 0.3120646, 0.2137803, 
    0.1087957, 0.1553343, 0.2217962, 0.2093595, 0.1911846, 0.2532879, 
    0.1490013, 0.07836127, 0.1687007, 0.2494828,
  0.2358134, 0.2126149, 0.2356896, 0.1738291, 0.1507286, 0.08959562, 
    0.06962321, 0.1166687, 0.1295951, 0.1699873, 0.1839669, 0.1733753, 
    0.223774, 0.2456874, 0.1909486, 0.1460492, 0.1540906, 0.1345527, 
    0.1456487, 0.1318647, 0.1905632, 0.1312152, 0.1404134, 0.1251079, 
    0.1633743, 0.1928893, 0.08064206, 0.303361, 0.2173042,
  0.2188824, 0.2018915, 0.2402058, 0.2238295, 0.1761357, 0.1443947, 
    0.1633602, 0.1848077, 0.1226395, 0.1612302, 0.1522868, 0.1340365, 
    0.1378341, 0.1350711, 0.1688894, 0.1617167, 0.1225478, 0.09117518, 
    0.106058, 0.1824306, 0.2063088, 0.2052141, 0.1518742, 0.1623932, 
    0.2042652, 0.1451535, 0.1897256, 0.1464701, 0.2605345,
  0.01376628, 0.0127796, 0.01179292, 0.01080624, 0.009819556, 0.008832875, 
    0.007846192, 0.01342232, 0.01531012, 0.01719793, 0.01908573, 0.02097354, 
    0.02286134, 0.02474914, 0.02288338, 0.02318256, 0.02348174, 0.02378092, 
    0.0240801, 0.02437929, 0.02467847, 0.02638381, 0.0251835, 0.0239832, 
    0.0227829, 0.02158259, 0.02038229, 0.01918198, 0.01455563,
  0.0773934, 0.01769838, 0.01103279, 0.0005913008, -2.696734e-06, 
    -0.000663338, -0.000628295, -0.0006541255, 5.819374e-05, 1.282991e-05, 
    0.006922478, 0.0233007, 0.04065827, 0.2054963, 0.1588583, 0.2227035, 
    0.3127964, 0.343788, 0.3370081, 0.3847696, 0.4042505, 0.3558302, 
    0.343577, 0.2551608, 0.3101984, 0.3631437, 0.3430937, 0.2639049, 0.1748558,
  0.2485923, 0.3345769, 0.2967941, 0.3655946, 0.2552648, 0.1610665, 
    0.2154581, 0.2530704, 0.2090666, 0.2403131, 0.2268906, 0.101177, 
    0.1585391, 0.2402429, 0.3469629, 0.3761561, 0.3249983, 0.3442967, 
    0.3850178, 0.3761465, 0.3492553, 0.340881, 0.3647853, 0.279523, 0.341917, 
    0.2283431, 0.1931266, 0.2676955, 0.2474993,
  0.341346, 0.3191662, 0.312442, 0.3364866, 0.314786, 0.3058679, 0.2435867, 
    0.3345446, 0.3502123, 0.3341233, 0.2866304, 0.2816648, 0.2678016, 
    0.2897739, 0.2644301, 0.2275529, 0.251878, 0.2057936, 0.2247162, 
    0.2156642, 0.2318703, 0.2101054, 0.24652, 0.2161687, 0.2414894, 
    0.2446751, 0.2553422, 0.2495114, 0.296868,
  0.1922409, 0.1792462, 0.2114661, 0.1493099, 0.1660762, 0.2070071, 
    0.1738585, 0.1881186, 0.1867411, 0.2128654, 0.2014397, 0.1848795, 
    0.1316283, 0.1529055, 0.1067104, 0.07888417, 0.1339843, 0.1537418, 
    0.1714627, 0.1502992, 0.1686615, 0.1777492, 0.1609044, 0.1250496, 
    0.1646944, 0.1872446, 0.177165, 0.1710979, 0.1743596,
  0.07056825, 0.06707741, 0.04424734, 0.0975231, 0.09003472, 0.07288714, 
    0.07855374, 0.08324553, 0.07391586, 0.08004577, 0.0616782, 0.08609474, 
    0.05872472, 0.06166565, 0.07740691, 0.1131644, 0.1337456, 0.1091944, 
    0.1335824, 0.1341617, 0.1647917, 0.07217823, 0.09549587, 0.09270211, 
    0.05298571, 0.07128765, 0.1065839, 0.112632, 0.1490996,
  0.01117923, 0.02170896, 0.06186642, 0.02477593, 0.07310206, 0.06384354, 
    0.04107136, 0.02483498, 0.02725925, 0.04807427, 0.1180843, 0.03869328, 
    0.04616321, 0.03081573, 0.03647017, 0.08619142, 0.08537262, 0.06739476, 
    0.08005831, 0.07756606, 0.1419712, 0.03075932, 0.01731304, 0.004417103, 
    0.05830446, 0.07613859, 0.08692057, 0.07381295, 0.01928427,
  2.131332e-05, 0.01276647, 0.001826728, 0.01724637, 0.02703634, 0.06048196, 
    0.06442475, 0.04714521, 0.06577686, 0.0166427, 0.001478752, 0.00485891, 
    0.02547482, 0.02642896, 0.07409889, 0.05073509, 0.05194284, 0.08484869, 
    0.04720409, 0.005312133, 0.00235101, 3.714834e-06, 1.231668e-07, 
    0.0007615035, 0.02704476, 0.02188889, 0.01379329, 0.001136798, 
    1.147637e-06,
  0.001231627, 0.1420929, 0.1418238, 0.1032913, 0.03765111, 0.05208512, 
    0.08097867, 0.06701013, 0.1088338, 0.03344218, 0.1037226, 0.1015328, 
    0.1200279, 0.05525943, 0.06070261, 0.04516628, 0.034276, 0.03656583, 
    0.005644702, 0.001743245, 0.002607357, 0.005399508, 0.007888432, 
    0.09621745, 0.1336534, 0.01254605, 0.04679196, 0.001594037, 6.438218e-05,
  0.07805394, 0.1892067, 0.1264543, 0.01679925, 0.008761163, 0.003803171, 
    0.004578084, 0.009092439, 0.06855889, 0.2222981, 0.07481791, 0.01283079, 
    0.07913907, 0.07606696, 0.04226333, 0.007058564, 0.007652644, 0.00599304, 
    0.01184447, 0.004103779, 0.02249232, 0.02328248, 0.1254857, 0.2452445, 
    0.2036928, 0.06610721, 0.07518286, 0.04576654, 0.04919838,
  0.03368824, 0.01460844, 0.01921842, 0.1982801, 0.004231622, 0.005451884, 
    0.03303285, 0.006625126, 0.01201623, 0.03884072, 0.01297488, 0.04446039, 
    0.04630107, 0.1045443, 0.1019987, 0.08935627, 0.07354201, 0.02586683, 
    0.01878473, 0.04728395, 0.09717116, 0.007509936, 0.01316622, 0.02097941, 
    0.01541379, 0.003253464, 0.001022242, 0.01425197, 0.08149341,
  0.0008656689, 0.0007291093, 0.006599014, 0.004168886, 0.06300318, 
    0.001232461, 0.01924956, 0.0008957362, 0.05934662, 0.007581056, 
    0.01637861, 0.02155664, 0.01866156, 0.002627859, 0.002867449, 
    0.002498555, 0.01055086, 0.0007647782, 0.0002371309, 0.000741799, 
    0.0004113094, 0.03271998, 0.005823051, 0.03565641, 0.008577474, 
    0.04997443, 0.007420741, 8.948336e-05, 0.01217617,
  0.005056406, 0.02457822, 0.01015323, 0.01963386, 0.0975658, 0.03127918, 
    0.02729647, 0.04451577, 0.1441921, 0.2087585, 0.1728371, 0.1261758, 
    0.1461285, 0.08348073, 0.06814223, 0.01520409, 0.01003452, 0.04624563, 
    0.01519971, 0.008407511, 0.02051032, 0.03723907, 0.02767676, 0.05215838, 
    0.04991649, 0.06604993, 0.03004905, 0.01576344, 0.001261851,
  0.05399546, 0.04472816, 0.1344004, 0.1135226, 0.10569, 0.05551511, 
    0.1705082, 0.04845836, 0.03846059, 0.08276698, 0.08103755, 0.1225438, 
    0.1212181, 0.1363265, 0.1773809, 0.1775596, 0.1555509, 0.1082554, 
    0.09805636, 0.1011617, 0.1410214, 0.1024633, 0.1276555, 0.1612603, 
    0.128227, 0.1044904, 0.08706893, 0.04892458, 0.06738131,
  0.1619969, 0.1610539, 0.1428573, 0.1059946, 0.1053765, 0.122727, 0.1692086, 
    0.2173044, 0.217838, 0.2256156, 0.2172944, 0.1996042, 0.2182535, 
    0.184934, 0.2089098, 0.1640139, 0.1952816, 0.2011765, 0.1861486, 
    0.1781669, 0.1563729, 0.1677459, 0.1732265, 0.2196445, 0.2357066, 
    0.1968984, 0.1264482, 0.109031, 0.1390294,
  0.244601, 0.2156774, 0.151346, 0.197256, 0.14934, 0.1326291, 0.1658652, 
    0.2146006, 0.2749279, 0.2035794, 0.1605783, 0.1539425, 0.2587465, 
    0.2652591, 0.1167759, 0.2075431, 0.2294908, 0.3343494, 0.2254047, 
    0.09598254, 0.1702189, 0.2139233, 0.2128379, 0.1878847, 0.2436894, 
    0.1467366, 0.1268392, 0.1761051, 0.2682179,
  0.2390207, 0.1903045, 0.2269075, 0.1733131, 0.1371845, 0.08799304, 
    0.06157093, 0.1016439, 0.1310879, 0.1760621, 0.1915631, 0.1811315, 
    0.2102183, 0.235996, 0.2005512, 0.1336659, 0.1646004, 0.1429143, 
    0.1545215, 0.140892, 0.171523, 0.1230202, 0.1564656, 0.1312061, 
    0.1488382, 0.2415227, 0.1293274, 0.3107716, 0.2198718,
  0.2346064, 0.2326315, 0.2809169, 0.2251861, 0.1634118, 0.1347746, 
    0.1701567, 0.1840303, 0.1313, 0.1604936, 0.152336, 0.1288578, 0.1378609, 
    0.1307519, 0.1650144, 0.1562637, 0.1211234, 0.08635259, 0.1168905, 
    0.2135833, 0.2021894, 0.2090982, 0.1656279, 0.152592, 0.1953481, 
    0.1655298, 0.2120847, 0.1406516, 0.2678784,
  0.03935826, 0.0359525, 0.03254674, 0.02914099, 0.02573523, 0.02232947, 
    0.01892371, 0.0290094, 0.03116137, 0.03331334, 0.03546531, 0.03761728, 
    0.03976925, 0.04192123, 0.03925078, 0.04193962, 0.04462846, 0.0473173, 
    0.05000614, 0.05269498, 0.05538382, 0.06303114, 0.06159609, 0.06016104, 
    0.05872598, 0.05729093, 0.05585588, 0.05442083, 0.04208286,
  0.1750273, 0.03664485, 0.01924461, 0.004788102, 0.002300672, 0.01600462, 
    0.00812393, 0.01017272, 0.005845995, 0.0002851197, 0.01140563, 
    0.04237735, 0.06495433, 0.2120197, 0.1832365, 0.2892829, 0.3441054, 
    0.3846995, 0.3522466, 0.412148, 0.4774331, 0.4238766, 0.3439192, 
    0.2450008, 0.2864106, 0.3760816, 0.3442996, 0.2807474, 0.2252182,
  0.294926, 0.3746251, 0.3782639, 0.3754638, 0.2972576, 0.1664065, 0.2268993, 
    0.2979044, 0.262695, 0.2825474, 0.2863102, 0.1215266, 0.1521417, 
    0.255818, 0.3943954, 0.3982177, 0.3122715, 0.3823392, 0.3927598, 
    0.3269333, 0.3410767, 0.3637984, 0.3836223, 0.2841044, 0.3731784, 
    0.2346149, 0.1932822, 0.3301863, 0.2725653,
  0.3118739, 0.2930381, 0.2979766, 0.339605, 0.2975792, 0.3245742, 0.2616228, 
    0.3629188, 0.384609, 0.3515171, 0.3149063, 0.2882354, 0.2799672, 
    0.2786604, 0.2776007, 0.2339482, 0.2599735, 0.2198839, 0.2526664, 
    0.2128606, 0.2361071, 0.2207367, 0.2278721, 0.2286343, 0.2156599, 
    0.2581211, 0.2881783, 0.2463477, 0.2832898,
  0.2078662, 0.1739545, 0.2156518, 0.1592954, 0.1688186, 0.2094075, 0.179009, 
    0.1914888, 0.2002865, 0.2115062, 0.1930271, 0.1894711, 0.136125, 
    0.1577904, 0.1050839, 0.0804313, 0.1438285, 0.1679085, 0.1797285, 
    0.1453905, 0.1711336, 0.1779995, 0.1569411, 0.1255928, 0.1596726, 
    0.190286, 0.1844296, 0.1842928, 0.1677087,
  0.07778153, 0.07329495, 0.04562083, 0.09893645, 0.09336279, 0.08723882, 
    0.0800176, 0.08974618, 0.07987635, 0.09120276, 0.07132857, 0.0801596, 
    0.07685079, 0.0708281, 0.09305365, 0.1306199, 0.1459331, 0.1217147, 
    0.1435368, 0.1282756, 0.1667821, 0.06532817, 0.100897, 0.09715201, 
    0.06367706, 0.08003065, 0.1148988, 0.1121939, 0.160902,
  0.01239449, 0.01643416, 0.06940956, 0.02510745, 0.09101412, 0.05241798, 
    0.04486675, 0.01867618, 0.02894974, 0.04936666, 0.08662596, 0.03625942, 
    0.06461755, 0.03761777, 0.04327497, 0.08976816, 0.06899533, 0.0650551, 
    0.08579184, 0.07760075, 0.14509, 0.04304804, 0.02139934, 0.006340623, 
    0.06379604, 0.06593359, 0.07409962, 0.08725405, 0.01822766,
  -1.600585e-06, 0.04378019, 0.003523381, 0.01202618, 0.02368778, 0.05201826, 
    0.05191109, 0.04832571, 0.05852403, 0.005624953, 0.008000877, 0.02423177, 
    0.02800127, 0.02857346, 0.06682268, 0.0446864, 0.05156202, 0.08376441, 
    0.04421123, 0.01046473, 0.00202243, 0.0007212877, 9.279475e-08, 
    0.0001372997, 0.02485828, 0.02905632, 0.01766542, 0.004089593, 
    -1.183174e-06,
  0.0002774944, 0.1151089, 0.1488974, 0.1097119, 0.03045768, 0.04440365, 
    0.07195265, 0.06701551, 0.09553646, 0.03128159, 0.09425611, 0.09235626, 
    0.1247949, 0.05087041, 0.05098779, 0.04292032, 0.0307318, 0.03329819, 
    0.006476178, 0.00112731, 0.004766852, 0.003986365, 0.00640129, 0.0681521, 
    0.1146672, 0.01868575, 0.05395759, 0.001115393, 2.231681e-05,
  0.05095655, 0.1169302, 0.05207575, 0.02413502, 0.006693849, 0.004191121, 
    0.005556102, 0.008568315, 0.05878819, 0.1889012, 0.07081322, 0.0132213, 
    0.0710009, 0.06315433, 0.0355626, 0.008915267, 0.01186558, 0.008233973, 
    0.01339095, 0.004762697, 0.02236222, 0.01743004, 0.1085897, 0.180842, 
    0.1862759, 0.05842546, 0.07395882, 0.03888843, 0.03870409,
  0.01698278, 0.00595353, 0.009649241, 0.2298089, 0.003015436, 0.005213677, 
    0.02995984, 0.007738873, 0.01160063, 0.03188016, 0.01519153, 0.03999955, 
    0.04230258, 0.0972854, 0.08777843, 0.07887515, 0.05751829, 0.02389195, 
    0.02421657, 0.04812476, 0.0836232, 0.01050837, 0.01398883, 0.02380437, 
    0.01398703, 0.00246524, 0.0005993128, 0.004731488, 0.03011266,
  2.402886e-05, 7.248618e-05, 0.001082683, 0.001347719, 0.0165446, 
    0.0002202494, 0.02278238, 0.0002601416, 0.0349883, 0.002564584, 
    0.01563886, 0.02328669, 0.01923324, 0.007116233, 0.005533728, 
    0.007215395, 0.01310262, 0.00555333, -1.736204e-05, -0.0001949387, 
    0.002622492, 0.03043922, 0.009284347, 0.03817984, 0.01195336, 0.05287334, 
    0.006297658, 1.453495e-05, 0.0004886043,
  0.001211144, 0.01687259, 0.01126043, 0.01421427, 0.09860034, 0.02645576, 
    0.007102236, 0.03422001, 0.1355583, 0.2179946, 0.177617, 0.1269545, 
    0.1466671, 0.07616877, 0.07616787, 0.01360492, 0.01667549, 0.05236445, 
    0.01627781, 0.01078508, 0.01145061, 0.04530257, 0.03343769, 0.06746985, 
    0.05636013, 0.08006389, 0.02869913, 0.01704445, 0.0006853707,
  0.05296523, 0.03866705, 0.141189, 0.114745, 0.105054, 0.03977239, 
    0.1667111, 0.03864967, 0.02870774, 0.08358422, 0.08168654, 0.120345, 
    0.1272474, 0.1367995, 0.1696143, 0.1854779, 0.1566663, 0.1231199, 
    0.09052511, 0.1053914, 0.1498305, 0.1074608, 0.1416608, 0.1630946, 
    0.1432755, 0.1094475, 0.09060862, 0.05827958, 0.07759728,
  0.1587211, 0.1632826, 0.1302055, 0.1261353, 0.1009109, 0.1272458, 
    0.1882376, 0.2272718, 0.1926202, 0.2139751, 0.2267446, 0.201999, 
    0.2176335, 0.2129048, 0.2261354, 0.1853106, 0.2090699, 0.1905701, 
    0.1825214, 0.1837394, 0.1439973, 0.1668577, 0.1674934, 0.2357937, 
    0.2358057, 0.2002937, 0.1356244, 0.1311362, 0.1439032,
  0.2548264, 0.2018424, 0.1624253, 0.1976081, 0.1533534, 0.1364771, 
    0.1891357, 0.2322678, 0.281474, 0.2140168, 0.1482487, 0.147144, 0.258992, 
    0.2616798, 0.1171072, 0.215598, 0.2459718, 0.3501421, 0.2204464, 
    0.1038499, 0.1731705, 0.2098686, 0.1953498, 0.1763905, 0.2536585, 
    0.1513433, 0.1499953, 0.1672773, 0.2485983,
  0.2468041, 0.1852474, 0.2282675, 0.1794855, 0.1554104, 0.1123429, 
    0.06789555, 0.09632077, 0.1266124, 0.1672522, 0.2024827, 0.1836779, 
    0.1907969, 0.2437146, 0.2006751, 0.1356891, 0.194211, 0.1500136, 
    0.1731265, 0.1533712, 0.16424, 0.1375175, 0.1593794, 0.1342905, 
    0.1431208, 0.2544692, 0.1693035, 0.3222494, 0.2416883,
  0.2548131, 0.2525626, 0.3073382, 0.2589821, 0.1856884, 0.1414319, 
    0.1841408, 0.1867008, 0.139364, 0.1637937, 0.1582809, 0.1309692, 
    0.1392225, 0.1292672, 0.1691086, 0.1601108, 0.1273898, 0.08985595, 
    0.1346071, 0.216042, 0.1947866, 0.213369, 0.1826463, 0.1440828, 
    0.1926011, 0.1731167, 0.2136387, 0.1236375, 0.2793387,
  0.09950393, 0.09355982, 0.08761572, 0.08167162, 0.07572751, 0.0697834, 
    0.0638393, 0.07740065, 0.07980301, 0.08220538, 0.08460775, 0.08701012, 
    0.08941249, 0.09181485, 0.0712947, 0.07917061, 0.08704654, 0.09492247, 
    0.1027984, 0.1106743, 0.1185502, 0.1222727, 0.1179385, 0.1136044, 
    0.1092702, 0.104936, 0.1006018, 0.09626761, 0.1042592,
  0.2569093, 0.1310901, 0.01723669, 0.0178816, 0.01875071, 0.0446869, 
    0.03035036, 0.0328792, 0.01542767, 0.005390423, 0.02136033, 0.05324518, 
    0.1075026, 0.2140442, 0.1818199, 0.2456461, 0.3162446, 0.3692451, 
    0.3569196, 0.4378716, 0.5192595, 0.4511342, 0.3440912, 0.2507358, 
    0.2716821, 0.3602304, 0.3727483, 0.3036061, 0.2773899,
  0.3229248, 0.3713134, 0.3232666, 0.4035501, 0.3396472, 0.1577234, 0.249527, 
    0.2949731, 0.3137069, 0.3029005, 0.2844292, 0.1277679, 0.1662967, 
    0.2973315, 0.3774858, 0.4234013, 0.3364377, 0.3470122, 0.4214685, 
    0.3477703, 0.3243351, 0.3316703, 0.3759089, 0.2925596, 0.351261, 
    0.2441305, 0.1860579, 0.3107728, 0.2934399,
  0.3570126, 0.3562706, 0.3506255, 0.3624005, 0.292743, 0.3465729, 0.294481, 
    0.3821928, 0.3991075, 0.342918, 0.3019661, 0.3075576, 0.3046969, 
    0.3130508, 0.2824298, 0.2487223, 0.2686324, 0.224, 0.2210523, 0.2230498, 
    0.2324261, 0.2115915, 0.2510519, 0.2261111, 0.2418157, 0.2732432, 
    0.3056766, 0.2410048, 0.3106833,
  0.2123026, 0.1919857, 0.2214686, 0.1648501, 0.1687247, 0.2121372, 
    0.1823876, 0.1970438, 0.2062008, 0.2151663, 0.2019954, 0.1922075, 
    0.1403589, 0.1637761, 0.1014041, 0.1061883, 0.1651922, 0.1847576, 
    0.1960948, 0.1753026, 0.1969559, 0.2018964, 0.1776256, 0.1389939, 
    0.1713992, 0.1833119, 0.2031586, 0.1881262, 0.1819731,
  0.08526763, 0.0864591, 0.05543401, 0.1091433, 0.09888241, 0.09734423, 
    0.0926923, 0.09926614, 0.09375398, 0.1276313, 0.08294943, 0.07126792, 
    0.07224669, 0.08744937, 0.1253733, 0.1465334, 0.1614792, 0.1389447, 
    0.1498442, 0.1371473, 0.1598956, 0.08299814, 0.1053334, 0.1096538, 
    0.0750376, 0.09808704, 0.1435326, 0.1149523, 0.1685868,
  0.01257416, 0.01748371, 0.07096057, 0.02365091, 0.0779563, 0.03800549, 
    0.04438387, 0.01698899, 0.02820225, 0.0412126, 0.04668258, 0.01885611, 
    0.101654, 0.05052749, 0.04229021, 0.1013624, 0.06156904, 0.06967475, 
    0.08815376, 0.06675023, 0.1492911, 0.06621845, 0.02580773, 0.00629519, 
    0.07431515, 0.06994206, 0.07196203, 0.08328759, 0.03229748,
  1.494145e-07, 0.02794518, 0.05026341, 0.01892802, 0.03127857, 0.04754529, 
    0.05896625, 0.0542733, 0.05811186, 0.003845698, 0.01281338, 0.04257918, 
    0.03451948, 0.03144688, 0.06426329, 0.04749745, 0.05466871, 0.09742294, 
    0.04399873, 0.02138859, 0.008346021, 0.006928258, 1.040936e-07, 
    7.604333e-05, 0.02691304, 0.0496998, 0.03996813, 0.01584983, 1.594428e-05,
  5.104103e-05, 0.09727049, 0.1161005, 0.1171283, 0.03395438, 0.04124386, 
    0.06539506, 0.06782624, 0.08946054, 0.03024669, 0.1022466, 0.08799508, 
    0.1239674, 0.04476389, 0.04578561, 0.04324758, 0.03072777, 0.03136926, 
    0.009611368, 0.003348583, 0.007378153, 0.003794363, 0.003062856, 
    0.0679263, 0.1075255, 0.02520493, 0.0666283, 0.002173695, 4.291279e-06,
  0.03606261, 0.08514666, 0.03032813, 0.04357085, 0.006326664, 0.006022447, 
    0.00711607, 0.008476292, 0.05414843, 0.1761921, 0.06802782, 0.01669526, 
    0.05998679, 0.05232831, 0.03580046, 0.01328288, 0.01441465, 0.01073727, 
    0.01779878, 0.0071739, 0.02671187, 0.01734085, 0.09343864, 0.1578364, 
    0.1802975, 0.05377842, 0.07438426, 0.03481222, 0.03218769,
  0.005326645, 0.003271066, 0.0052859, 0.2326905, 0.003032257, 0.005597041, 
    0.02455543, 0.0111847, 0.01218529, 0.02958765, 0.0214072, 0.03751177, 
    0.04286048, 0.09619471, 0.08566995, 0.06797945, 0.05023191, 0.02765639, 
    0.03388782, 0.0554338, 0.07673638, 0.0123169, 0.01676361, 0.02907573, 
    0.01662243, 0.0009818882, 3.353012e-05, 0.001079712, 0.01282497,
  5.561231e-06, 7.724628e-06, 2.34815e-05, 0.0003374599, 0.004657858, 
    7.772345e-05, 0.0141516, 0.0001159604, 0.02576203, 0.0115851, 0.01520195, 
    0.02790225, 0.02485817, 0.01046249, 0.01577428, 0.01364655, 0.01785369, 
    0.0156309, 1.592357e-05, -9.788041e-05, 0.0003685471, 0.02837967, 
    0.01226584, 0.04686131, 0.01673607, 0.05896049, 0.01147234, 9.347174e-06, 
    1.692917e-05,
  0.004406706, 0.008296324, 0.01413509, 0.01427232, 0.09551503, 0.01659821, 
    -0.001760187, 0.02519555, 0.1096728, 0.2331003, 0.1909491, 0.1216167, 
    0.1339778, 0.07812969, 0.09440078, 0.01914256, 0.02448785, 0.06286348, 
    0.0308874, 0.01697113, 0.01046295, 0.05814179, 0.04496629, 0.07275152, 
    0.062938, 0.08572539, 0.03050676, 0.01574297, 0.000269202,
  0.04635126, 0.03768136, 0.1543123, 0.1275702, 0.09131066, 0.03245086, 
    0.1622743, 0.03260925, 0.02169586, 0.08104791, 0.0848631, 0.1232382, 
    0.1264497, 0.1342734, 0.1691623, 0.2103216, 0.1568326, 0.129599, 
    0.08808667, 0.1219899, 0.1618278, 0.1203101, 0.1576343, 0.169212, 
    0.1484896, 0.1227961, 0.09389191, 0.06980447, 0.09722774,
  0.1677377, 0.1695289, 0.1598116, 0.1445982, 0.1049324, 0.1437428, 0.208582, 
    0.2354862, 0.166846, 0.1836973, 0.2065314, 0.1959772, 0.2321424, 
    0.2359916, 0.2694869, 0.2301887, 0.2364913, 0.2253801, 0.1845563, 
    0.1879637, 0.1441274, 0.1934382, 0.2080499, 0.2634332, 0.2733387, 
    0.2101275, 0.1614422, 0.1659294, 0.1626542,
  0.2337966, 0.2136458, 0.1889529, 0.2163148, 0.1880119, 0.1596112, 
    0.2398829, 0.2451389, 0.3007359, 0.1997487, 0.1503168, 0.1586484, 
    0.2657955, 0.3063339, 0.1393068, 0.2486956, 0.2784273, 0.363376, 
    0.2588784, 0.129125, 0.1831453, 0.2238337, 0.2455336, 0.213971, 
    0.2624242, 0.167388, 0.1833572, 0.1941941, 0.2418565,
  0.2739885, 0.1848357, 0.2385544, 0.2139637, 0.2108895, 0.1095038, 
    0.08147632, 0.1101601, 0.1351251, 0.175008, 0.2504913, 0.2396401, 
    0.2185603, 0.2745862, 0.2351108, 0.1440364, 0.2115422, 0.1471989, 
    0.2067076, 0.1808169, 0.1722475, 0.1570687, 0.162659, 0.122165, 
    0.1463362, 0.2689949, 0.2074625, 0.3251772, 0.2835396,
  0.2596065, 0.2941493, 0.3337416, 0.2822452, 0.2196988, 0.1741644, 
    0.2171006, 0.2119963, 0.1578975, 0.1871674, 0.1728835, 0.1474293, 
    0.1608747, 0.150587, 0.1645647, 0.1602529, 0.1358212, 0.09210415, 
    0.1041809, 0.1976656, 0.2007025, 0.230556, 0.2046851, 0.1474841, 
    0.1922287, 0.1830796, 0.2150721, 0.1204446, 0.3026505,
  0.1866047, 0.1776485, 0.1686922, 0.1597359, 0.1507797, 0.1418234, 
    0.1328671, 0.1548714, 0.1592802, 0.163689, 0.1680978, 0.1725066, 
    0.1769154, 0.1813242, 0.1729005, 0.1841065, 0.1953126, 0.2065186, 
    0.2177246, 0.2289306, 0.2401366, 0.2420152, 0.2353566, 0.2286981, 
    0.2220395, 0.215381, 0.2087224, 0.2020638, 0.1937697,
  0.3389983, 0.2135645, 0.04883349, 0.02928096, 0.02326649, 0.06639002, 
    0.05780225, 0.05275622, 0.02834735, 0.01280962, 0.03052926, 0.08814628, 
    0.1479647, 0.2293739, 0.221619, 0.2532555, 0.2967793, 0.3363757, 
    0.3401413, 0.4463725, 0.5456406, 0.4628579, 0.3347701, 0.2495343, 
    0.2538538, 0.3605046, 0.3685773, 0.3243544, 0.2658195,
  0.2980976, 0.3714406, 0.3035029, 0.3824619, 0.3595135, 0.157193, 0.3043472, 
    0.3099949, 0.3369808, 0.3063745, 0.2727212, 0.1204699, 0.1689538, 
    0.3294603, 0.3644406, 0.3892354, 0.3158388, 0.3076059, 0.3662179, 
    0.3206417, 0.3172857, 0.3354587, 0.3479669, 0.3103524, 0.335135, 
    0.2224019, 0.159606, 0.2754725, 0.2947544,
  0.3595472, 0.3376858, 0.3638537, 0.3347239, 0.314599, 0.3595883, 0.3038447, 
    0.3953712, 0.3869621, 0.3659843, 0.3094331, 0.3182625, 0.3139435, 
    0.3055211, 0.2924198, 0.253824, 0.2873143, 0.2420655, 0.2183225, 
    0.2094107, 0.2338153, 0.2363715, 0.2916478, 0.2281942, 0.2379681, 
    0.2823078, 0.322459, 0.2641066, 0.2915101,
  0.2344273, 0.214955, 0.2381419, 0.1656261, 0.1689138, 0.2106768, 0.203727, 
    0.2140528, 0.2162436, 0.2204856, 0.2189915, 0.2201003, 0.1604758, 
    0.1825968, 0.09602658, 0.1288987, 0.1908423, 0.2030219, 0.2188174, 
    0.2004623, 0.2181832, 0.2118779, 0.1940598, 0.1397692, 0.1825949, 0.2047, 
    0.2029452, 0.2189713, 0.1973671,
  0.1030172, 0.09835555, 0.06201439, 0.1106861, 0.1034757, 0.1080109, 
    0.1013691, 0.1229134, 0.1144493, 0.1459822, 0.1171761, 0.07299721, 
    0.06733926, 0.09236697, 0.1433682, 0.1731389, 0.1811357, 0.1538873, 
    0.1559188, 0.1447526, 0.1658007, 0.09881845, 0.1184687, 0.1265356, 
    0.08574782, 0.114521, 0.1585165, 0.1166151, 0.1659455,
  0.01804652, 0.0184569, 0.07601571, 0.02761221, 0.07073438, 0.03914411, 
    0.04773369, 0.01764868, 0.03142322, 0.03744139, 0.01773949, 0.009691455, 
    0.09491809, 0.04712334, 0.04849702, 0.1142409, 0.07118119, 0.07890949, 
    0.09543528, 0.08244155, 0.1486037, 0.07617384, 0.03552407, 0.006022418, 
    0.07569405, 0.07783081, 0.08026897, 0.08553313, 0.04617724,
  2.547768e-05, 0.01133431, 0.05258825, 0.02733305, 0.03579973, 0.04776105, 
    0.06335251, 0.06979204, 0.06198427, 0.003093481, 0.003661101, 0.05196947, 
    0.04024344, 0.03942196, 0.120199, 0.05584103, 0.05414576, 0.1093773, 
    0.04446569, 0.0286686, 0.03108378, 0.01848061, -2.078127e-06, 
    3.946997e-05, 0.03011483, 0.04931622, 0.05431047, 0.03500032, 0.0008894537,
  -8.472498e-06, 0.08097397, 0.1070942, 0.1217032, 0.03676355, 0.04232228, 
    0.06244393, 0.07050793, 0.08520716, 0.03139555, 0.1110637, 0.08260346, 
    0.1246746, 0.04362469, 0.04201286, 0.03952058, 0.02883441, 0.03013001, 
    0.01557217, 0.008022142, 0.008696869, 0.003799751, 0.0008087236, 
    0.07006721, 0.102979, 0.04396008, 0.08630068, 0.004190542, 0.0001620169,
  0.0285752, 0.07043126, 0.023831, 0.1039506, 0.007010354, 0.007720318, 
    0.00985872, 0.01058809, 0.06569976, 0.1761283, 0.06961218, 0.01953294, 
    0.05446891, 0.04425272, 0.03427435, 0.01656657, 0.01926579, 0.01633788, 
    0.02123356, 0.01630632, 0.03180362, 0.0275082, 0.07686807, 0.1464171, 
    0.1740005, 0.04906119, 0.07507651, 0.03626041, 0.03460433,
  0.002238022, 0.001003171, 0.003944498, 0.1743943, 0.003917803, 0.006075076, 
    0.02088845, 0.01188335, 0.01311812, 0.02969001, 0.03270083, 0.04065499, 
    0.04276786, 0.09213512, 0.08488505, 0.0617379, 0.048928, 0.03506603, 
    0.04577049, 0.06156944, 0.07621466, 0.01492878, 0.02889345, 0.03370696, 
    0.02382841, 0.001111079, 1.693892e-05, 4.982878e-05, 0.007142023,
  3.309332e-06, 4.080283e-06, 3.381549e-06, 0.0001279142, 0.003515149, 
    9.421513e-05, 0.003889805, 0.0001268663, 0.0159162, 0.009056401, 
    0.0160574, 0.04177841, 0.03590253, 0.02973039, 0.02600672, 0.02006791, 
    0.02473648, 0.0217227, 3.184925e-05, 0.0007120363, 6.616367e-06, 
    0.03425998, 0.01805816, 0.04796626, 0.0209555, 0.06637107, 0.01577584, 
    4.881243e-06, 1.103246e-05,
  0.003424977, 0.001872581, 0.01173355, 0.01171904, 0.08838908, 0.009715815, 
    -0.003678481, 0.01876623, 0.08681151, 0.2486545, 0.1976736, 0.1279158, 
    0.1241708, 0.0754769, 0.09510472, 0.02298334, 0.03928576, 0.07927656, 
    0.036268, 0.01888725, 0.009417889, 0.06998278, 0.05539718, 0.08160499, 
    0.06490679, 0.08880858, 0.04462554, 0.0121608, 0.000520625,
  0.03591647, 0.03670153, 0.1583042, 0.1329634, 0.06089531, 0.01795672, 
    0.1640019, 0.0224429, 0.0183901, 0.06405622, 0.08610576, 0.1248885, 
    0.1366893, 0.1417209, 0.1676176, 0.2143433, 0.1714863, 0.1425627, 
    0.09568682, 0.1392426, 0.145596, 0.1154195, 0.1692669, 0.1857336, 
    0.1652591, 0.1343924, 0.1039667, 0.09087323, 0.1292,
  0.1930204, 0.209532, 0.1543469, 0.1381085, 0.1099331, 0.1538468, 0.2007135, 
    0.2390337, 0.1406822, 0.1351655, 0.182626, 0.1946888, 0.2374359, 
    0.2728658, 0.2751756, 0.2666446, 0.2467981, 0.2441387, 0.1800556, 
    0.1802463, 0.1257849, 0.1686036, 0.220082, 0.2803641, 0.2882007, 
    0.2219347, 0.1767948, 0.2007705, 0.1857254,
  0.2532797, 0.2387897, 0.2134204, 0.2064921, 0.1797261, 0.1728286, 
    0.2248419, 0.2280053, 0.3227741, 0.1774559, 0.1531448, 0.1731007, 
    0.2605506, 0.2883112, 0.1664739, 0.2435915, 0.2746828, 0.3579681, 
    0.243372, 0.1336649, 0.1802676, 0.2004513, 0.2059394, 0.2076574, 
    0.2394471, 0.1766618, 0.2145458, 0.213086, 0.2512233,
  0.2901484, 0.1882097, 0.2199715, 0.1847973, 0.1962429, 0.1247278, 
    0.1074235, 0.1027668, 0.1468729, 0.1984337, 0.2594022, 0.2164427, 
    0.1936386, 0.2183257, 0.2199967, 0.1238456, 0.1794957, 0.1193883, 
    0.1606846, 0.1396305, 0.1884335, 0.1361983, 0.1592975, 0.1037289, 
    0.1405541, 0.2942308, 0.2077458, 0.3061714, 0.3177553,
  0.2922792, 0.2866267, 0.3294472, 0.2785924, 0.2205498, 0.158029, 0.2193633, 
    0.2193363, 0.1683647, 0.1900196, 0.1769953, 0.1484285, 0.1501058, 
    0.1512372, 0.1612947, 0.1465433, 0.1136184, 0.1003499, 0.1097238, 
    0.1905931, 0.2170299, 0.2471711, 0.2123922, 0.1538782, 0.1866223, 
    0.1930378, 0.2171578, 0.1390039, 0.2858995,
  0.2604305, 0.2523368, 0.2442431, 0.2361493, 0.2280556, 0.2199619, 
    0.2118682, 0.2397867, 0.2476655, 0.2555444, 0.2634232, 0.2713021, 
    0.2791809, 0.2870597, 0.2869223, 0.2969728, 0.3070232, 0.3170737, 
    0.3271242, 0.3371746, 0.3472251, 0.3357796, 0.325944, 0.3161085, 
    0.3062729, 0.2964373, 0.2866017, 0.2767661, 0.2669055,
  0.3683235, 0.2778891, 0.1302605, 0.04114081, 0.04057662, 0.08194969, 
    0.0756909, 0.077512, 0.04605762, 0.02559761, 0.0515918, 0.1219252, 
    0.1849578, 0.2332949, 0.2405377, 0.2489473, 0.317525, 0.3117755, 
    0.3226305, 0.4236273, 0.5790104, 0.4835609, 0.3242009, 0.2396403, 
    0.2830411, 0.3251401, 0.3519225, 0.3363423, 0.2808355,
  0.2781923, 0.380942, 0.3121606, 0.3612978, 0.3583976, 0.1529121, 0.3477704, 
    0.3220096, 0.3581735, 0.3300115, 0.271394, 0.1238358, 0.1628753, 
    0.3369433, 0.4061928, 0.4030093, 0.3336605, 0.3057619, 0.3492274, 
    0.2949102, 0.3091463, 0.3555981, 0.3817736, 0.3195564, 0.3490283, 
    0.2181602, 0.1665131, 0.2824293, 0.2881953,
  0.3243476, 0.3139806, 0.3164913, 0.3098167, 0.3010821, 0.3625813, 
    0.2797937, 0.3986423, 0.37855, 0.3560474, 0.3110359, 0.3251401, 
    0.3229431, 0.3062189, 0.3089342, 0.2553152, 0.2687902, 0.2561104, 
    0.2361738, 0.2303872, 0.2424317, 0.2568765, 0.2988763, 0.2389659, 
    0.277703, 0.2538313, 0.2958382, 0.2724285, 0.2783224,
  0.2279913, 0.2186563, 0.2496715, 0.177665, 0.1882631, 0.2170461, 0.225914, 
    0.2264818, 0.2433989, 0.2294205, 0.2310702, 0.2216334, 0.1677656, 
    0.1922818, 0.1112734, 0.1649495, 0.2228204, 0.2294329, 0.262316, 
    0.1977952, 0.240502, 0.2127309, 0.1897964, 0.142864, 0.2126178, 
    0.2159806, 0.2098086, 0.2357812, 0.2059336,
  0.1100701, 0.1129739, 0.07894656, 0.1262238, 0.1023468, 0.1205597, 
    0.116308, 0.1466813, 0.1263726, 0.1527167, 0.1232029, 0.09480564, 
    0.06718766, 0.09941598, 0.1505874, 0.1734794, 0.1913704, 0.165217, 
    0.1597197, 0.1562882, 0.16966, 0.1209157, 0.1320903, 0.1441296, 
    0.07086865, 0.114687, 0.1703893, 0.1270658, 0.1670299,
  0.02183078, 0.01558727, 0.05649164, 0.03182469, 0.06615269, 0.05092768, 
    0.05677013, 0.02634838, 0.03788806, 0.03232111, 0.01469038, 0.002491328, 
    0.05050695, 0.07437971, 0.05963877, 0.1122306, 0.0895794, 0.09633787, 
    0.1075989, 0.08016001, 0.1381373, 0.08740342, 0.04989326, 0.005776393, 
    0.07003485, 0.08267484, 0.08901985, 0.08920197, 0.04730454,
  0.0003337379, 0.002704143, 0.0168051, 0.03282038, 0.034182, 0.04801276, 
    0.06591164, 0.06664447, 0.05488447, 0.002710176, 0.003766315, 
    0.008658775, 0.04553252, 0.04069075, 0.1165089, 0.05458016, 0.05233658, 
    0.1123574, 0.04244952, 0.04314122, 0.06714997, 0.05369002, 0.0001962529, 
    1.965449e-05, 0.04144165, 0.05221491, 0.05351252, 0.06429066, 0.0143526,
  0.0001406869, 0.06611148, 0.09888698, 0.1284505, 0.03521997, 0.03969356, 
    0.05745658, 0.06554034, 0.07932785, 0.02983141, 0.0939418, 0.06914365, 
    0.1326499, 0.04352694, 0.03794365, 0.03217715, 0.02558726, 0.02653277, 
    0.01694157, 0.01193422, 0.009417214, 0.005255369, 8.214994e-05, 
    0.07060663, 0.1033707, 0.0420096, 0.0945088, 0.008179335, 0.0008364609,
  0.02574706, 0.06224267, 0.02156179, 0.130341, 0.008330401, 0.009555725, 
    0.01241457, 0.01109968, 0.07518499, 0.1715749, 0.06988461, 0.02014345, 
    0.04982894, 0.0404367, 0.03189014, 0.01613846, 0.02165252, 0.02029537, 
    0.02077553, 0.01577155, 0.03972215, 0.03294666, 0.06387816, 0.1374073, 
    0.166381, 0.04237168, 0.0680501, 0.04509062, 0.03932785,
  0.001004267, 0.0002406639, 0.0009260591, 0.1096228, 0.005071325, 
    0.008184788, 0.01985312, 0.009687274, 0.01470757, 0.0352104, 0.04126983, 
    0.04152506, 0.04216432, 0.0823823, 0.07581767, 0.05246207, 0.05106733, 
    0.04592638, 0.05692902, 0.06804898, 0.07239383, 0.01721182, 0.04446406, 
    0.04521851, 0.03125266, 0.001785524, 7.321962e-06, 1.231086e-05, 
    0.00433585,
  2.693487e-06, 1.711447e-06, 8.734532e-07, 4.122582e-05, 0.002207005, 
    0.0001185125, 0.0002502417, 0.0001855594, 0.006552555, 0.007111672, 
    0.02334885, 0.05491587, 0.0447243, 0.03580096, 0.0418017, 0.03614487, 
    0.03227255, 0.02740781, 0.002073156, -0.0001260955, 4.490595e-06, 
    0.05015943, 0.02475239, 0.04715192, 0.02267223, 0.06637767, 0.02974675, 
    1.628375e-06, 5.415928e-06,
  0.001584768, 0.0003598921, 0.01064487, 0.007462932, 0.07721116, 
    0.006414072, -0.003172448, 0.01278999, 0.07646259, 0.2521816, 0.1824469, 
    0.1392892, 0.1326658, 0.07584094, 0.09272681, 0.03962656, 0.04728023, 
    0.0839899, 0.04098272, 0.02969826, 0.009575771, 0.07841186, 0.05533347, 
    0.08149526, 0.08051045, 0.08685031, 0.05761231, 0.02542072, 0.003915444,
  0.02056926, 0.03605711, 0.1472866, 0.1270455, 0.04500999, 0.008673119, 
    0.162916, 0.02052451, 0.01544996, 0.05766595, 0.08957041, 0.1176881, 
    0.1369272, 0.1424703, 0.181269, 0.2183348, 0.1891426, 0.1394011, 0.12908, 
    0.143356, 0.1142481, 0.1185286, 0.1828615, 0.1884519, 0.1784696, 
    0.1474135, 0.1113141, 0.1059533, 0.1289027,
  0.2151444, 0.2119846, 0.1631466, 0.1307988, 0.08337773, 0.1356799, 
    0.1713241, 0.2428316, 0.1163776, 0.1082579, 0.149118, 0.1914481, 
    0.2170883, 0.3031068, 0.2676263, 0.2757037, 0.2815654, 0.2478904, 
    0.179864, 0.1888481, 0.1160945, 0.1286615, 0.1700739, 0.2861232, 
    0.2866464, 0.2236817, 0.2047295, 0.2097798, 0.2034931,
  0.2690852, 0.2550476, 0.2413549, 0.1993774, 0.1826166, 0.1892352, 
    0.1737542, 0.1945425, 0.3008267, 0.1854234, 0.141858, 0.1885456, 
    0.2603392, 0.2827912, 0.1622641, 0.210882, 0.2494882, 0.3538695, 
    0.2053678, 0.1235516, 0.1849778, 0.1804376, 0.180385, 0.2130284, 
    0.2413811, 0.1839651, 0.246131, 0.2441912, 0.2662773,
  0.2967727, 0.2347012, 0.2158614, 0.1648281, 0.1611774, 0.1213623, 
    0.0770186, 0.1064766, 0.1429395, 0.2059655, 0.2211631, 0.2002541, 
    0.1641686, 0.2109827, 0.1964816, 0.1077956, 0.1448127, 0.112682, 
    0.1124973, 0.09792241, 0.1684233, 0.1119017, 0.1457867, 0.1046996, 
    0.1452844, 0.3119661, 0.1988258, 0.2682231, 0.2942353,
  0.2906277, 0.2709664, 0.3320976, 0.2503451, 0.1997143, 0.1461267, 
    0.1866831, 0.1860611, 0.1366643, 0.1750766, 0.1647819, 0.1547959, 
    0.1368087, 0.1294502, 0.1393334, 0.139889, 0.09409299, 0.07347767, 
    0.1339138, 0.2045724, 0.2111675, 0.2300333, 0.2196911, 0.1622492, 
    0.1869761, 0.2042809, 0.2230597, 0.1552794, 0.2548282,
  0.3095116, 0.3049006, 0.3002895, 0.2956784, 0.2910674, 0.2864563, 
    0.2818452, 0.3319516, 0.3433677, 0.3547838, 0.3661999, 0.377616, 
    0.3890321, 0.4004483, 0.387911, 0.3938026, 0.3996942, 0.4055858, 
    0.4114774, 0.4173691, 0.4232607, 0.4071594, 0.3944628, 0.3817661, 
    0.3690695, 0.3563728, 0.3436762, 0.3309796, 0.3132005,
  0.3598066, 0.3379216, 0.2207053, 0.06492186, 0.06299896, 0.1040219, 
    0.0944512, 0.09269685, 0.05391591, 0.03258417, 0.1030539, 0.1321791, 
    0.2153203, 0.21235, 0.2066207, 0.2542104, 0.3261109, 0.289603, 0.3003424, 
    0.4047875, 0.5980781, 0.5006961, 0.3257405, 0.2543569, 0.3141454, 
    0.314881, 0.3449634, 0.3126732, 0.3094462,
  0.3216433, 0.3436642, 0.3190182, 0.3399359, 0.3229984, 0.1409214, 
    0.3657102, 0.3406693, 0.3675535, 0.3299621, 0.2666458, 0.1129924, 
    0.1598982, 0.3664686, 0.4586174, 0.4067816, 0.3663384, 0.3238585, 
    0.3992659, 0.3309283, 0.3621157, 0.3695405, 0.4139751, 0.3397084, 
    0.3375835, 0.3095417, 0.184891, 0.3167892, 0.2855054,
  0.4017005, 0.3477, 0.3196611, 0.3232343, 0.3089262, 0.3609449, 0.3543276, 
    0.4329959, 0.4162633, 0.3795559, 0.3454396, 0.3474149, 0.361212, 
    0.3401274, 0.3419104, 0.2956716, 0.2968382, 0.2803061, 0.2832198, 
    0.2975983, 0.2944598, 0.341098, 0.3160415, 0.3169461, 0.3441746, 
    0.2801099, 0.3488485, 0.3033492, 0.3339677,
  0.2530142, 0.250177, 0.2951075, 0.2216069, 0.221613, 0.2465547, 0.2550637, 
    0.2777033, 0.2705658, 0.2672632, 0.2628478, 0.2642197, 0.2151161, 
    0.2410415, 0.1700576, 0.2336609, 0.2670089, 0.287426, 0.3055299, 
    0.246905, 0.2685352, 0.2243955, 0.2302048, 0.1473104, 0.2280456, 
    0.2365613, 0.2455392, 0.2836653, 0.2457733,
  0.1357787, 0.1414941, 0.1044898, 0.1567153, 0.1272499, 0.1601122, 
    0.1324067, 0.1788474, 0.1605047, 0.1984062, 0.1503628, 0.1097955, 
    0.09036179, 0.140623, 0.1737828, 0.184943, 0.2140797, 0.188015, 
    0.1814111, 0.1703373, 0.1928381, 0.1456652, 0.1717706, 0.1531924, 
    0.0697939, 0.1262853, 0.1629802, 0.1513054, 0.1899423,
  0.03428192, 0.02265679, 0.04233934, 0.05304891, 0.06287676, 0.07020454, 
    0.06883061, 0.0540401, 0.05404373, 0.0393641, 0.0180817, 9.696136e-05, 
    0.02409368, 0.1058258, 0.08812776, 0.1377372, 0.0898628, 0.104645, 
    0.1210528, 0.08105287, 0.1285054, 0.1159774, 0.07627986, 0.004902343, 
    0.06091423, 0.08898775, 0.1058506, 0.08283652, 0.06095641,
  0.0139625, 0.002467869, 0.01326639, 0.03371258, 0.03256693, 0.05653559, 
    0.07112893, 0.07667921, 0.06270554, 0.002260366, 0.00274928, 0.00239979, 
    0.03928508, 0.04332426, 0.08911501, 0.06389463, 0.06383481, 0.1046441, 
    0.03630216, 0.03723254, 0.05891817, 0.07346928, 0.01384721, 5.623563e-06, 
    0.0510743, 0.06648132, 0.04463545, 0.0737246, 0.06630442,
  0.004207256, 0.05076544, 0.0896749, 0.1265398, 0.03146547, 0.03494828, 
    0.05164815, 0.05867248, 0.06449618, 0.02625648, 0.07353861, 0.05866227, 
    0.1220986, 0.03911303, 0.03224497, 0.02682713, 0.02230772, 0.02318971, 
    0.0188359, 0.01615585, 0.01170357, 0.009519349, 8.840781e-05, 0.06542563, 
    0.09944989, 0.03510262, 0.08229285, 0.01681143, 0.00415197,
  0.02742081, 0.05382672, 0.01984533, 0.09249286, 0.01088223, 0.01203203, 
    0.01484919, 0.01192219, 0.08266655, 0.173801, 0.06437054, 0.01927979, 
    0.04442447, 0.03219852, 0.02790096, 0.01656904, 0.01883003, 0.01944011, 
    0.02001714, 0.01669838, 0.04155803, 0.0346706, 0.04799204, 0.1247674, 
    0.1553443, 0.03607649, 0.05966573, 0.04113816, 0.03807169,
  0.0004788842, 8.004487e-05, 9.423625e-05, 0.07147324, 0.007323471, 
    0.0157108, 0.02156843, 0.01212446, 0.01690587, 0.03646608, 0.04983445, 
    0.03714276, 0.04001467, 0.0712475, 0.07032979, 0.04892865, 0.05669191, 
    0.05855706, 0.06962433, 0.07293037, 0.06466383, 0.0178555, 0.05503561, 
    0.05218831, 0.03746677, 0.005550213, 0.0001864418, 9.863868e-07, 
    0.002726097,
  2.095061e-06, 7.980744e-07, 3.446968e-07, 6.916984e-05, 0.001320191, 
    0.0002044499, 0.0002081758, 0.0001781999, 0.00264314, 0.01782089, 
    0.02763833, 0.06643151, 0.04453491, 0.03087941, 0.03703445, 0.05245721, 
    0.04535723, 0.06933242, 0.01799285, 0.0001274558, 2.032417e-06, 
    0.0675729, 0.04043513, 0.04365867, 0.02815181, 0.05147436, 0.05534603, 
    3.950751e-06, 3.536093e-06,
  0.0003646851, 0.0002533168, 0.01366223, 0.005538923, 0.06485392, 
    0.005446607, -0.002609913, 0.01028398, 0.06643695, 0.252118, 0.1719022, 
    0.1957881, 0.1756052, 0.1213678, 0.09829251, 0.06172277, 0.06535283, 
    0.1146842, 0.05487713, 0.03814866, 0.007989052, 0.09172332, 0.05663326, 
    0.09298418, 0.09261785, 0.09109735, 0.07271007, 0.05830047, 0.007926,
  0.01082931, 0.0367182, 0.1242172, 0.1286568, 0.03246563, 0.004192145, 
    0.1568342, 0.01552477, 0.01320525, 0.04772468, 0.09526459, 0.1098415, 
    0.1455051, 0.1742452, 0.207333, 0.2541017, 0.225633, 0.1633769, 0.170774, 
    0.1480365, 0.1085237, 0.1196293, 0.2032735, 0.2169307, 0.2006521, 
    0.1648013, 0.1272833, 0.1288279, 0.1217498,
  0.2058717, 0.215024, 0.1610284, 0.1145393, 0.06600649, 0.1250294, 
    0.1536721, 0.2377173, 0.09319815, 0.07435501, 0.1162234, 0.1953109, 
    0.245967, 0.3338634, 0.3076265, 0.3091049, 0.2666741, 0.2707809, 
    0.1949434, 0.2372267, 0.0985691, 0.1227244, 0.1628734, 0.2904284, 
    0.3003455, 0.2521273, 0.2558596, 0.2499782, 0.2258708,
  0.2594388, 0.2919696, 0.2502829, 0.2394218, 0.1642371, 0.1546726, 
    0.1484972, 0.1864787, 0.269387, 0.2021835, 0.1219738, 0.1939641, 
    0.2558727, 0.3130579, 0.2227305, 0.2135843, 0.2878888, 0.350219, 
    0.2310009, 0.1131636, 0.1718294, 0.1860953, 0.1598632, 0.2331886, 
    0.2779492, 0.2034414, 0.2615408, 0.2895533, 0.2858689,
  0.3129386, 0.2505497, 0.240021, 0.1990221, 0.237849, 0.1484644, 0.09618134, 
    0.1422626, 0.1479148, 0.221998, 0.1955339, 0.1831093, 0.1753219, 
    0.1820155, 0.1993527, 0.1193736, 0.1318024, 0.1138098, 0.1064378, 
    0.09703988, 0.16634, 0.1027081, 0.1157562, 0.1211859, 0.1299857, 
    0.324792, 0.1709146, 0.2397472, 0.3558193,
  0.2637222, 0.2647066, 0.3424508, 0.2420547, 0.2004633, 0.1689014, 
    0.2077685, 0.1829161, 0.1376753, 0.1528553, 0.2119903, 0.1705857, 
    0.1398009, 0.1245309, 0.1317437, 0.1409316, 0.09188241, 0.08572783, 
    0.1147954, 0.1570786, 0.180792, 0.2042947, 0.2317598, 0.1789138, 
    0.1738651, 0.2138143, 0.228363, 0.1529644, 0.2787997,
  0.3526247, 0.3518659, 0.3511071, 0.3503483, 0.3495895, 0.3488307, 
    0.3480719, 0.3586443, 0.371695, 0.3847458, 0.3977965, 0.4108472, 
    0.423898, 0.4369487, 0.437179, 0.438966, 0.4407529, 0.4425399, 0.4443269, 
    0.4461139, 0.4479009, 0.4467133, 0.4326344, 0.4185554, 0.4044766, 
    0.3903976, 0.3763187, 0.3622398, 0.3532317,
  0.3526637, 0.3520482, 0.3003882, 0.09087397, 0.08974694, 0.1341968, 
    0.1245975, 0.1262526, 0.06451362, 0.03837232, 0.1448652, 0.1651738, 
    0.2284945, 0.1694578, 0.2122654, 0.2289682, 0.2998322, 0.3371653, 
    0.3154546, 0.3923247, 0.6145706, 0.5332125, 0.3305525, 0.2736996, 
    0.3162245, 0.3254994, 0.3520617, 0.2827084, 0.3321277,
  0.3866363, 0.3884625, 0.3168319, 0.309761, 0.3012879, 0.1508833, 0.3498788, 
    0.3982658, 0.3646813, 0.3323654, 0.2656792, 0.1032245, 0.1695758, 
    0.3682241, 0.5031306, 0.4152089, 0.4171626, 0.3981236, 0.4901319, 
    0.4341032, 0.4163138, 0.4110928, 0.4192725, 0.3695751, 0.3461991, 
    0.3166964, 0.2127825, 0.3868059, 0.2945051,
  0.4368776, 0.3694658, 0.3539293, 0.3483876, 0.3125384, 0.347336, 0.3661835, 
    0.4416049, 0.4647576, 0.4206963, 0.376363, 0.3634421, 0.4043396, 
    0.376406, 0.3452927, 0.3403785, 0.3644787, 0.2858341, 0.3341593, 
    0.3545771, 0.3491569, 0.4161578, 0.3627258, 0.3704624, 0.399464, 
    0.3911551, 0.3747631, 0.3811355, 0.3753143,
  0.2882549, 0.3125776, 0.3296248, 0.2523774, 0.2496326, 0.2807754, 
    0.2958984, 0.2909856, 0.2819133, 0.3008775, 0.2852258, 0.3137526, 
    0.2715484, 0.3016021, 0.2266102, 0.2642281, 0.2768681, 0.2999023, 
    0.3123912, 0.3131695, 0.320691, 0.3127285, 0.3318914, 0.1597424, 
    0.2489641, 0.2648447, 0.2385077, 0.3251858, 0.2815318,
  0.1675512, 0.1723652, 0.1554506, 0.1915123, 0.1722367, 0.1743596, 
    0.1673087, 0.2364351, 0.2274296, 0.27653, 0.1818414, 0.1657474, 
    0.08264537, 0.169341, 0.2043318, 0.1973223, 0.2320871, 0.2442315, 
    0.2009556, 0.2204627, 0.2281733, 0.1492817, 0.2077371, 0.1787352, 
    0.07760544, 0.1236376, 0.1481716, 0.1475187, 0.2165764,
  0.08214928, 0.03603544, 0.03619184, 0.08971845, 0.06476238, 0.08049646, 
    0.09916431, 0.1237112, 0.1241891, 0.07087537, 0.02160736, -1.12464e-05, 
    0.01368829, 0.1230462, 0.08178459, 0.1497424, 0.1141773, 0.1480712, 
    0.1747931, 0.1104505, 0.1403815, 0.1170985, 0.1197224, 0.004544249, 
    0.06327666, 0.1068203, 0.1318102, 0.08738212, 0.07524946,
  0.0548146, 0.002515, 0.002906936, 0.04285417, 0.03991017, 0.06637336, 
    0.06725633, 0.07849379, 0.08964694, 0.002085451, 0.0009436366, 
    0.001532572, 0.04999464, 0.05156673, 0.102386, 0.06374413, 0.09319892, 
    0.1027115, 0.0371034, 0.03457794, 0.04694964, 0.09918429, 0.07745794, 
    6.883082e-05, 0.05583156, 0.1048593, 0.04671277, 0.05029092, 0.1051806,
  0.007885923, 0.03704442, 0.08219597, 0.1213344, 0.03127554, 0.03482411, 
    0.04622229, 0.04896941, 0.05189382, 0.02488809, 0.06044429, 0.06037337, 
    0.1143145, 0.036113, 0.03160673, 0.02666566, 0.02256279, 0.02397887, 
    0.02479947, 0.02695893, 0.01837253, 0.02571312, 0.001254445, 0.05812912, 
    0.0990675, 0.02282031, 0.07412849, 0.0359696, 0.02698029,
  0.02997545, 0.04365108, 0.01834252, 0.05950499, 0.01820918, 0.01745725, 
    0.01862855, 0.01586464, 0.07953826, 0.175451, 0.05716508, 0.02140706, 
    0.04116348, 0.03055621, 0.02654365, 0.01902274, 0.01791948, 0.01977385, 
    0.02006487, 0.01678675, 0.03821241, 0.03172629, 0.03733442, 0.1115796, 
    0.1466017, 0.03536437, 0.05292984, 0.03849293, 0.03989331,
  0.0002299689, 2.999786e-05, 1.275016e-05, 0.0434835, 0.01358112, 
    0.03567558, 0.02755321, 0.01690711, 0.02102671, 0.04838355, 0.05057316, 
    0.03550313, 0.0379678, 0.0600976, 0.06749103, 0.04556644, 0.06544891, 
    0.08832505, 0.093493, 0.07433625, 0.06227259, 0.02253293, 0.06317195, 
    0.05871017, 0.04609821, 0.02219559, 0.003382117, 3.725729e-07, 0.001973988,
  1.487924e-06, 4.216409e-07, 1.273298e-07, 6.166389e-05, 0.0005754043, 
    0.0002772857, 0.0001258281, 5.117161e-05, 0.0007114615, 0.0405324, 
    0.04467961, 0.07111749, 0.04197773, 0.03040863, 0.03526529, 0.06281165, 
    0.07776456, 0.1109337, 0.06287181, 0.007443879, 9.325573e-07, 0.07450686, 
    0.08226997, 0.06295153, 0.04123106, 0.06035463, 0.07658917, 0.007397574, 
    2.119003e-06,
  4.683226e-05, 0.004135459, 0.01318253, 0.004930045, 0.05216599, 
    0.002421767, -0.002283345, 0.00578993, 0.06113692, 0.2594098, 0.1911878, 
    0.2159716, 0.2009602, 0.1577526, 0.1472877, 0.1324434, 0.1414451, 
    0.1540867, 0.1148475, 0.05267999, 0.007938665, 0.1091629, 0.07121034, 
    0.1379785, 0.114769, 0.1326556, 0.08174379, 0.07293437, 0.009081844,
  0.007158444, 0.02924381, 0.092879, 0.1355787, 0.02198033, 0.002828222, 
    0.1514294, 0.01142191, 0.01160441, 0.04472245, 0.09868288, 0.1093268, 
    0.1939964, 0.2178339, 0.2532762, 0.2869012, 0.2514786, 0.2435599, 
    0.2577749, 0.1596774, 0.08606987, 0.1267503, 0.2115769, 0.1961984, 
    0.2442213, 0.1622872, 0.166216, 0.1418027, 0.1280617,
  0.185878, 0.2727213, 0.1389766, 0.1204487, 0.05533073, 0.1239346, 
    0.1573578, 0.2314967, 0.07585102, 0.05140683, 0.09858814, 0.1997472, 
    0.2802891, 0.3756139, 0.4016292, 0.3275108, 0.2788656, 0.2930795, 
    0.2333104, 0.2464717, 0.08935925, 0.1199994, 0.1741481, 0.3037766, 
    0.3425633, 0.2747069, 0.3442555, 0.2846729, 0.2424935,
  0.2807942, 0.3291327, 0.2326571, 0.1973384, 0.2017536, 0.1687101, 
    0.1317301, 0.1462837, 0.2095278, 0.1276619, 0.1259005, 0.1830932, 
    0.2398146, 0.310093, 0.3164723, 0.2361512, 0.3139933, 0.3572295, 
    0.2428178, 0.06460497, 0.1450182, 0.1652723, 0.1723418, 0.2598899, 
    0.3314283, 0.2198514, 0.2584329, 0.3147821, 0.3079951,
  0.3308445, 0.2552689, 0.2313964, 0.2390464, 0.2825235, 0.115906, 0.1243924, 
    0.1530123, 0.1708421, 0.2413405, 0.1928683, 0.228312, 0.1653776, 
    0.1640983, 0.2011998, 0.1097591, 0.1328421, 0.1093397, 0.1124655, 
    0.104996, 0.1664053, 0.09101821, 0.1184893, 0.1264197, 0.1315566, 
    0.3352935, 0.1540769, 0.2253485, 0.4213766,
  0.333195, 0.3416661, 0.336031, 0.2641179, 0.2075603, 0.1845215, 0.1941587, 
    0.1502888, 0.1200393, 0.1806644, 0.1737835, 0.1724343, 0.1556996, 
    0.1452947, 0.1432576, 0.1483146, 0.1345382, 0.1015086, 0.1393981, 
    0.1754773, 0.1843079, 0.2123469, 0.2200774, 0.1911504, 0.1573224, 
    0.2136792, 0.2102834, 0.1673036, 0.300125,
  0.3740732, 0.375968, 0.3778628, 0.3797576, 0.3816524, 0.3835472, 0.385442, 
    0.4001679, 0.4140986, 0.4280292, 0.4419599, 0.4558907, 0.4698213, 
    0.483752, 0.4789675, 0.476529, 0.4740906, 0.4716522, 0.4692137, 
    0.4667753, 0.4643368, 0.4578617, 0.4444746, 0.4310876, 0.4177006, 
    0.4043135, 0.3909265, 0.3775395, 0.3725574,
  0.3499639, 0.365207, 0.3369541, 0.1552776, 0.1182794, 0.1616202, 0.1697578, 
    0.1718127, 0.08033745, 0.04774961, 0.1738818, 0.2128515, 0.2684239, 
    0.1101223, 0.2021115, 0.2592595, 0.2958004, 0.3802162, 0.3249844, 
    0.4096808, 0.6423074, 0.5706556, 0.3366025, 0.2821323, 0.3123339, 
    0.3889217, 0.3282481, 0.2717782, 0.3228755,
  0.3984735, 0.379743, 0.3045983, 0.2561063, 0.2710622, 0.1692121, 0.2943124, 
    0.407745, 0.3594647, 0.3298405, 0.2670585, 0.1043609, 0.1576545, 
    0.3715977, 0.513611, 0.4292927, 0.4211237, 0.4836662, 0.5488015, 
    0.4708822, 0.4933643, 0.4813826, 0.4105372, 0.3812639, 0.3692387, 
    0.2881256, 0.2516022, 0.4212762, 0.343037,
  0.4499693, 0.3707263, 0.3562399, 0.371183, 0.3273738, 0.3604867, 0.3661921, 
    0.4136148, 0.4687448, 0.3969309, 0.3525872, 0.3996899, 0.4581429, 
    0.4048828, 0.3202258, 0.348962, 0.3577608, 0.3592713, 0.3397609, 
    0.3576867, 0.3480803, 0.4480465, 0.4436604, 0.3406834, 0.4555145, 
    0.4612645, 0.445511, 0.39342, 0.4024249,
  0.3237845, 0.3345078, 0.3336122, 0.2748233, 0.2769839, 0.3014601, 
    0.3342349, 0.2925963, 0.2959705, 0.3044497, 0.2833825, 0.3025026, 
    0.2616861, 0.2818896, 0.2162327, 0.2753925, 0.300221, 0.2773213, 
    0.3085308, 0.3496746, 0.3823708, 0.3848715, 0.3326043, 0.1780848, 
    0.2187804, 0.2465897, 0.2839829, 0.3357807, 0.2887968,
  0.2171195, 0.2227193, 0.1917474, 0.2488894, 0.2323207, 0.2557142, 
    0.2478617, 0.2715955, 0.2434773, 0.298037, 0.1727715, 0.1441245, 
    0.07373968, 0.2124723, 0.2444201, 0.2178003, 0.2181801, 0.2532962, 
    0.2143889, 0.2392286, 0.2644852, 0.1855001, 0.2285235, 0.2269078, 
    0.05310803, 0.1076142, 0.12311, 0.1421989, 0.242876,
  0.1672995, 0.04462877, 0.03326363, 0.119866, 0.08038399, 0.1284887, 
    0.1359431, 0.1408083, 0.2125214, 0.07910655, 0.01976899, -1.339882e-05, 
    0.01304946, 0.1031539, 0.07902984, 0.1063685, 0.1252403, 0.1246888, 
    0.1743566, 0.09926058, 0.1714379, 0.1157465, 0.1161784, 0.005849413, 
    0.08864211, 0.1216474, 0.1432591, 0.1020085, 0.1096387,
  0.1604347, 0.0006319331, 0.001805961, 0.04492885, 0.07253965, 0.07104899, 
    0.07339564, 0.1058734, 0.1089499, 0.008334832, 0.000295548, 0.0008099749, 
    0.07225092, 0.0663747, 0.09640621, 0.06350846, 0.08690281, 0.1081979, 
    0.05885775, 0.04677608, 0.05583154, 0.1125243, 0.2152524, 0.0002126388, 
    0.05411559, 0.09135845, 0.0555379, 0.05247656, 0.1636795,
  0.02458386, 0.03353083, 0.04677944, 0.1400923, 0.04668191, 0.04335427, 
    0.04903056, 0.04774877, 0.04959871, 0.02882545, 0.06006119, 0.06686162, 
    0.1029502, 0.03729565, 0.0348554, 0.03095266, 0.03202254, 0.03288954, 
    0.04208332, 0.06173431, 0.05069508, 0.1048813, 0.02171856, 0.05197379, 
    0.08962137, 0.009354059, 0.08865198, 0.08642917, 0.1019114,
  0.03817864, 0.03194905, 0.01343593, 0.03511992, 0.03658969, 0.03769982, 
    0.03625146, 0.02214974, 0.07630612, 0.1672406, 0.05330807, 0.02637584, 
    0.04171895, 0.03357104, 0.03236234, 0.02651667, 0.02032569, 0.0229145, 
    0.02544772, 0.01869191, 0.03415204, 0.03375855, 0.02585922, 0.09653387, 
    0.1257506, 0.037884, 0.05275764, 0.03758574, 0.04463894,
  0.0001264375, 1.226375e-05, 1.916742e-06, 0.02522086, 0.01594046, 
    0.1564881, 0.03830062, 0.03443576, 0.02872811, 0.07839715, 0.06326133, 
    0.04074671, 0.0401265, 0.06106091, 0.06788538, 0.05285073, 0.08677871, 
    0.1234761, 0.1135044, 0.09085555, 0.07121042, 0.07766709, 0.0589003, 
    0.06215704, 0.06533411, 0.0919594, 0.03205543, 4.334562e-06, 0.00114263,
  9.300088e-07, 2.489123e-07, 6.42744e-08, 8.699411e-05, 0.00022022, 
    0.0006622325, 1.159916e-05, 6.558742e-06, 0.0002679671, 0.07840672, 
    0.06962042, 0.08181713, 0.05352955, 0.04346935, 0.0539391, 0.07908479, 
    0.05906128, 0.1254353, 0.1684931, 0.02987017, 1.922037e-06, 0.08653267, 
    0.0791299, 0.06844012, 0.09656478, 0.09335878, 0.09288655, 0.0597196, 
    1.404451e-06,
  -3.102502e-06, 0.01276571, 0.01241932, 0.004376204, 0.0445405, 0.001529977, 
    -0.001928123, 0.002051605, 0.05063118, 0.2604207, 0.2018957, 0.2482276, 
    0.2451919, 0.1644628, 0.1894396, 0.193529, 0.1936062, 0.1754903, 
    0.2407804, 0.1097325, 0.006879349, 0.1291469, 0.0615019, 0.1124212, 
    0.1343947, 0.127352, 0.1248821, 0.1416968, 0.01489305,
  0.006875582, 0.01457482, 0.06858093, 0.129878, 0.01579091, 0.001495792, 
    0.1424309, 0.009012029, 0.01058934, 0.0404746, 0.1002519, 0.104417, 
    0.1972349, 0.2012895, 0.2378956, 0.2657928, 0.237237, 0.2851106, 
    0.286767, 0.1569078, 0.07311457, 0.1374957, 0.195795, 0.1808513, 
    0.2447805, 0.1735119, 0.2055314, 0.1938505, 0.1239408,
  0.1843985, 0.2380622, 0.1225175, 0.09894824, 0.04169238, 0.1295491, 
    0.148817, 0.2353445, 0.06140031, 0.03617328, 0.09633526, 0.1890646, 
    0.2857849, 0.349537, 0.3390514, 0.2785901, 0.2898531, 0.3111802, 
    0.2937676, 0.2426138, 0.08008862, 0.1275243, 0.1923217, 0.3249267, 
    0.3873199, 0.4214956, 0.3586909, 0.2179989, 0.2372601,
  0.2714831, 0.3170627, 0.2224753, 0.1755796, 0.1567593, 0.1490275, 
    0.1496071, 0.1382712, 0.1332221, 0.07128197, 0.1128898, 0.1572092, 
    0.1919916, 0.2931021, 0.3766449, 0.254002, 0.3232693, 0.3759664, 
    0.2170634, 0.03904347, 0.134101, 0.1540963, 0.2082198, 0.2725047, 
    0.4661168, 0.1603357, 0.2157769, 0.3005646, 0.3026487,
  0.3225338, 0.2516657, 0.2361052, 0.2431114, 0.2390248, 0.132658, 0.1200282, 
    0.127837, 0.1947991, 0.2638621, 0.2019379, 0.2793771, 0.1848187, 
    0.2053365, 0.2008716, 0.1224764, 0.1420524, 0.1021423, 0.1120378, 
    0.1178925, 0.1394466, 0.08540495, 0.1348656, 0.1293115, 0.1042399, 
    0.346897, 0.1418615, 0.186618, 0.417982,
  0.3318319, 0.3909618, 0.3372917, 0.2791483, 0.2359861, 0.1884357, 
    0.2034738, 0.1523531, 0.1420619, 0.2027908, 0.1751838, 0.1732344, 
    0.2070666, 0.1747356, 0.1694127, 0.1834957, 0.1582225, 0.1439132, 
    0.1974845, 0.22001, 0.1974612, 0.2291274, 0.2039221, 0.2032916, 
    0.1571582, 0.1998052, 0.1841107, 0.1822244, 0.3325581,
  0.3990711, 0.4014917, 0.4039123, 0.4063329, 0.4087535, 0.4111741, 
    0.4135947, 0.4215821, 0.4349256, 0.4482691, 0.4616127, 0.4749562, 
    0.4882997, 0.5016432, 0.510042, 0.5060339, 0.5020258, 0.4980177, 
    0.4940096, 0.4900016, 0.4859935, 0.4666843, 0.4549283, 0.4431722, 
    0.4314162, 0.4196602, 0.4079041, 0.3961481, 0.3971346,
  0.3569662, 0.376563, 0.3705755, 0.2285956, 0.1509343, 0.1905745, 0.2002629, 
    0.2001858, 0.08450233, 0.08417305, 0.2137399, 0.2470809, 0.2986587, 
    0.071732, 0.1819022, 0.2542342, 0.269439, 0.3996474, 0.3375175, 
    0.3874764, 0.667703, 0.6198478, 0.3580586, 0.2582822, 0.3246315, 
    0.4264998, 0.3321165, 0.2598865, 0.3331924,
  0.3479479, 0.305603, 0.2862395, 0.2054628, 0.2533125, 0.1792471, 0.2068538, 
    0.4128825, 0.3487282, 0.3253369, 0.2587799, 0.1010639, 0.1591727, 
    0.3147077, 0.439962, 0.4472068, 0.4184392, 0.4949134, 0.5387602, 
    0.4970087, 0.5422134, 0.5026778, 0.4415226, 0.4155869, 0.3743548, 
    0.2755722, 0.3482938, 0.4365304, 0.3333328,
  0.4412338, 0.3647967, 0.33844, 0.3681699, 0.3204416, 0.3739117, 0.3699264, 
    0.3819509, 0.4190453, 0.3804809, 0.3386689, 0.4223555, 0.4823794, 
    0.3986948, 0.3372587, 0.3680197, 0.3946998, 0.4155186, 0.3879196, 
    0.3559777, 0.3704941, 0.4222795, 0.4322439, 0.3282256, 0.4190039, 
    0.4704092, 0.4698454, 0.3676672, 0.3769682,
  0.3622488, 0.3436231, 0.3598884, 0.3028947, 0.2863449, 0.328951, 0.344403, 
    0.3110736, 0.303479, 0.3189713, 0.2956098, 0.3025432, 0.2698099, 
    0.216957, 0.2262719, 0.2387522, 0.3116871, 0.2782035, 0.2976708, 
    0.3590733, 0.3834881, 0.3482471, 0.2851883, 0.1832645, 0.1592846, 
    0.2363903, 0.2640822, 0.3300539, 0.3417765,
  0.2956162, 0.291489, 0.2010621, 0.2245125, 0.2457773, 0.2098271, 0.2210746, 
    0.2471867, 0.2366044, 0.2487308, 0.1732274, 0.1564238, 0.03826841, 
    0.1609978, 0.2943873, 0.1776474, 0.2249969, 0.2506435, 0.20389, 
    0.2536398, 0.2388757, 0.2369348, 0.2356281, 0.2668058, 0.05109539, 
    0.08551762, 0.1239938, 0.1637769, 0.2680328,
  0.2087748, 0.1074125, 0.01692275, 0.0902667, 0.1149026, 0.118059, 
    0.1308399, 0.1887286, 0.2144916, 0.05499308, 0.03798738, -2.35234e-05, 
    0.008570503, 0.06718879, 0.073733, 0.1216771, 0.08821198, 0.09074407, 
    0.1311549, 0.1068159, 0.1623065, 0.1009933, 0.1159158, 0.01179237, 
    0.0969298, 0.1146058, 0.1439619, 0.1113413, 0.1555551,
  0.2975093, -0.0001337932, 0.0006160391, 0.0673928, 0.08081233, 0.07973064, 
    0.08179992, 0.09725673, 0.1129311, 0.01097528, 9.768872e-05, 
    0.0003193541, 0.02991771, 0.06171126, 0.08898586, 0.07814792, 0.07851522, 
    0.1064593, 0.05497704, 0.05726361, 0.06834595, 0.08453815, 0.3013484, 
    0.000312122, 0.0531076, 0.09077469, 0.09199518, 0.05980089, 0.1156402,
  0.2799596, 0.03163039, 0.02836494, 0.1022412, 0.0804684, 0.07123919, 
    0.08192397, 0.05591089, 0.06542975, 0.04236691, 0.05963482, 0.05857653, 
    0.1072827, 0.07066678, 0.04473443, 0.06967242, 0.09959449, 0.07327627, 
    0.09773842, 0.1219787, 0.1265645, 0.1347308, 0.2476768, 0.03398236, 
    0.05564262, 0.002367177, 0.09938173, 0.09705068, 0.2200136,
  0.0503206, 0.02040512, 0.006672535, 0.03083488, 0.154825, 0.1976548, 
    0.1556385, 0.1175361, 0.05381545, 0.1231988, 0.1039813, 0.09913197, 
    0.056438, 0.0515425, 0.0477032, 0.0657665, 0.04985026, 0.0554175, 
    0.05941122, 0.03187296, 0.03977629, 0.04872891, 0.02327782, 0.07541518, 
    0.08454823, 0.04868343, 0.06333989, 0.04319257, 0.07572933,
  9.860769e-05, 2.473182e-06, 6.821188e-07, 0.01554925, 0.02387059, 
    0.1395427, 0.09129986, 0.1787021, 0.04776886, 0.1957447, 0.08763399, 
    0.06670292, 0.06115585, 0.06697549, 0.06132408, 0.05208407, 0.08235788, 
    0.1466786, 0.1497104, 0.1801268, 0.08637446, 0.1063452, 0.1080464, 
    0.06445649, 0.07696763, 0.2019025, 0.3599238, 0.0003460436, 0.0003354709,
  5.994126e-07, 1.701886e-07, 3.584326e-08, 0.0001692564, 9.541126e-05, 
    0.00473189, -4.962192e-06, -0.0003214223, 0.0001711765, 0.1237268, 
    0.1070289, 0.0982331, 0.07508696, 0.04298854, 0.03635584, 0.05011869, 
    0.06091877, 0.0693349, 0.2466918, 0.2078092, 2.99041e-05, 0.08713613, 
    0.03718092, 0.04517674, 0.06044875, 0.09696594, 0.1437277, 0.103774, 
    8.123664e-07,
  -6.422405e-06, 0.01371226, 0.009731171, 0.005002355, 0.04022032, 
    0.001233467, -0.001631482, -9.680956e-05, 0.04953898, 0.252186, 
    0.2165499, 0.2319441, 0.2844381, 0.2181678, 0.2555727, 0.2088765, 
    0.244179, 0.2000151, 0.3083776, 0.1175826, 0.007280286, 0.1484188, 
    0.05815412, 0.1066871, 0.1055682, 0.1223954, 0.1480606, 0.1500756, 
    0.01465093,
  0.006360784, 0.01157382, 0.05468536, 0.1265838, 0.02063604, 0.001071772, 
    0.133974, 0.01033356, 0.01009248, 0.03637192, 0.1009372, 0.1036572, 
    0.1801944, 0.1885366, 0.2205473, 0.2812623, 0.2615111, 0.2438935, 
    0.3025809, 0.1521221, 0.06737125, 0.1278916, 0.1658387, 0.1806097, 
    0.2763316, 0.2285369, 0.243885, 0.2810187, 0.1260356,
  0.1815789, 0.2217197, 0.07790719, 0.08907371, 0.04645076, 0.1139168, 
    0.1415055, 0.2129276, 0.04770168, 0.03548578, 0.0872564, 0.1994105, 
    0.2878533, 0.3362477, 0.268654, 0.2331071, 0.2677473, 0.319089, 
    0.2798681, 0.2492823, 0.0839265, 0.1242328, 0.1854934, 0.3377702, 
    0.3941969, 0.4578049, 0.3355484, 0.1570581, 0.2155153,
  0.2369019, 0.2775627, 0.2259412, 0.1631527, 0.1632874, 0.1464122, 
    0.1505784, 0.1181411, 0.09708118, 0.0423224, 0.06580896, 0.1059005, 
    0.1637169, 0.2493689, 0.45939, 0.2974651, 0.3339912, 0.3552209, 
    0.2268333, 0.03551183, 0.1310228, 0.1684121, 0.215764, 0.242729, 
    0.5221764, 0.1305846, 0.1597244, 0.23807, 0.2643088,
  0.3394901, 0.1978754, 0.2263615, 0.2301475, 0.2031418, 0.1374941, 
    0.1130951, 0.1348666, 0.2147898, 0.2483591, 0.2235687, 0.2831653, 
    0.2155265, 0.2249828, 0.1924209, 0.131989, 0.15035, 0.1198163, 
    0.09528684, 0.1413858, 0.1417009, 0.09139422, 0.1387491, 0.1281073, 
    0.07785974, 0.3438036, 0.1444057, 0.1401719, 0.421261,
  0.3269736, 0.3925233, 0.3310816, 0.2479288, 0.2581201, 0.2133244, 
    0.2298039, 0.146935, 0.1645952, 0.1964436, 0.1865695, 0.2009033, 
    0.2020549, 0.2166726, 0.2330849, 0.229155, 0.1988569, 0.1768, 0.2261521, 
    0.2518233, 0.223726, 0.2363603, 0.2167822, 0.2209965, 0.1609109, 
    0.1913183, 0.1836264, 0.1764813, 0.3130268,
  0.42602, 0.4295217, 0.4330234, 0.4365251, 0.4400268, 0.4435285, 0.4470302, 
    0.4618979, 0.4732041, 0.4845103, 0.4958165, 0.5071226, 0.5184288, 
    0.529735, 0.5366639, 0.5300044, 0.5233448, 0.5166852, 0.5100256, 
    0.503366, 0.4967064, 0.4650612, 0.456913, 0.4487647, 0.4406164, 
    0.4324681, 0.4243198, 0.4161715, 0.4232187,
  0.3806198, 0.4188244, 0.4107327, 0.2576415, 0.1852866, 0.1998676, 
    0.2174184, 0.2202071, 0.09368055, 0.100671, 0.2504775, 0.3118434, 
    0.3623566, 0.04412885, 0.1587663, 0.2616018, 0.2780614, 0.371015, 
    0.3185276, 0.3791543, 0.7233375, 0.6414595, 0.365774, 0.2504418, 
    0.3074093, 0.4535531, 0.3347178, 0.2660987, 0.3921221,
  0.3039086, 0.234012, 0.2755128, 0.1626719, 0.2290391, 0.1910716, 0.1347385, 
    0.3932571, 0.3430167, 0.3331941, 0.2373884, 0.09066828, 0.1544788, 
    0.2432427, 0.3705477, 0.4994146, 0.3780131, 0.4516378, 0.4946374, 
    0.5196069, 0.528483, 0.5090833, 0.46474, 0.4295194, 0.386981, 0.2794701, 
    0.3172636, 0.3844522, 0.3448699,
  0.4090796, 0.3291945, 0.2918246, 0.3445708, 0.312117, 0.3642046, 0.362666, 
    0.3384131, 0.3620581, 0.3468043, 0.3366014, 0.4199899, 0.4976071, 
    0.3875186, 0.3460613, 0.3794551, 0.4114576, 0.4363243, 0.4262865, 
    0.3802112, 0.3723161, 0.4073597, 0.3936261, 0.2866708, 0.390479, 
    0.4219521, 0.4708586, 0.3591414, 0.3474296,
  0.3379498, 0.3474135, 0.3729547, 0.3002709, 0.3007089, 0.3459823, 
    0.3401023, 0.309137, 0.3061653, 0.3081263, 0.2923277, 0.3122467, 
    0.2262927, 0.2028232, 0.1998626, 0.2040682, 0.2761528, 0.256274, 
    0.3106586, 0.3342343, 0.3136476, 0.2860219, 0.2624654, 0.1941956, 
    0.1231701, 0.2099719, 0.2446654, 0.3261316, 0.3686216,
  0.2820195, 0.2571476, 0.147327, 0.1774457, 0.2105851, 0.1844187, 0.1872522, 
    0.1994302, 0.2401619, 0.1887911, 0.0961001, 0.08215186, 0.02096695, 
    0.0924083, 0.327977, 0.1427943, 0.2075195, 0.1929778, 0.1741467, 
    0.2154414, 0.2166872, 0.2132416, 0.1596447, 0.296334, 0.0422918, 
    0.09425553, 0.1123205, 0.19909, 0.3046841,
  0.1476929, 0.09890269, 0.01112597, 0.09430996, 0.08981889, 0.07772952, 
    0.09718001, 0.1086777, 0.1102231, 0.02515988, 0.0323517, -5.332742e-05, 
    0.007040679, 0.03365581, 0.04638162, 0.09532645, 0.08027342, 0.08821499, 
    0.1051059, 0.07879117, 0.09777405, 0.04928852, 0.06784324, 0.02048403, 
    0.08084787, 0.08785552, 0.08034183, 0.08026102, 0.123349,
  0.1659441, -0.0001699401, 0.0001621231, 0.07606339, 0.04255213, 0.06515735, 
    0.04172725, 0.06158319, 0.07488315, 0.004386053, 3.447827e-05, 
    0.0001280897, 0.0128255, 0.05622503, 0.05408712, 0.04125266, 0.05979972, 
    0.05227934, 0.02312649, 0.0511574, 0.01512637, 0.04400263, 0.1370497, 
    0.06204807, 0.05359027, 0.07783073, 0.03136228, 0.01456018, 0.04420238,
  0.4051879, 0.06202494, 0.0211516, 0.09672689, 0.09929225, 0.03711641, 
    0.05914357, 0.06150181, 0.05294607, 0.02238972, 0.0472799, 0.0293044, 
    0.09365349, 0.05861255, 0.04504474, 0.02615446, 0.02702528, 0.03666347, 
    0.03154576, 0.02900961, 0.03527937, 0.05447356, 0.3804358, 0.02147799, 
    0.03533471, 0.0004958837, 0.03543675, 0.02304413, 0.0915474,
  0.1331216, 0.01412618, 0.001924791, 0.02562968, 0.04950698, 0.03989279, 
    0.0516154, 0.03121214, 0.05247537, 0.07749173, 0.04454041, 0.0982917, 
    0.03320522, 0.03696757, 0.04046904, 0.1078253, 0.1210227, 0.1258213, 
    0.09438933, 0.119181, 0.06899272, 0.1927243, 0.03937409, 0.05363736, 
    0.0531222, 0.03999556, 0.08365769, 0.08978824, 0.1675924,
  7.821719e-05, -1.940677e-07, 4.772164e-07, 0.009252525, 0.0223373, 
    0.04701855, 0.05848699, 0.06519035, 0.01599423, 0.0760017, 0.04631278, 
    0.04941796, 0.04065752, 0.0402, 0.03067089, 0.02546166, 0.04247332, 
    0.07870346, 0.1092366, 0.1148189, 0.05369321, 0.01610119, 0.2392745, 
    0.07774019, 0.03003488, 0.05760439, 0.2599369, 0.05085641, 9.858027e-05,
  4.386604e-07, 1.346096e-07, 2.520092e-08, 0.0004105358, 4.214121e-05, 
    0.008206776, -4.108179e-05, 0.01744386, 0.0001066586, 0.2106767, 
    0.1566132, 0.0856297, 0.05204186, 0.02274716, 0.01136184, 0.01245268, 
    0.0197885, 0.03314503, 0.2039829, 0.2056928, 0.0001828043, 0.07897417, 
    0.01511395, 0.01850371, 0.01935389, 0.04623055, 0.09685129, 0.05722503, 
    5.097606e-07,
  2.111035e-06, 0.009796805, 0.0100252, 0.003525339, 0.03126789, 0.001295162, 
    -0.001419828, -0.0002471563, 0.05126411, 0.2262774, 0.2202001, 0.2048187, 
    0.2956305, 0.246999, 0.1723827, 0.2016766, 0.2548629, 0.1834626, 
    0.2287467, 0.131039, 0.006499656, 0.1582284, 0.04591383, 0.09639214, 
    0.08363916, 0.08215967, 0.08894179, 0.09234326, 0.01571048,
  0.004494162, 0.006181713, 0.04548043, 0.1304969, 0.01939483, 0.000530745, 
    0.1283974, 0.008484074, 0.008543446, 0.03291435, 0.09635665, 0.09150912, 
    0.1649401, 0.1729957, 0.2003551, 0.2411833, 0.2738533, 0.2028337, 
    0.3046006, 0.1440501, 0.06323809, 0.1254581, 0.1458623, 0.2015355, 
    0.2845555, 0.1955977, 0.2158066, 0.2252944, 0.1160792,
  0.1466025, 0.1969621, 0.05700508, 0.07419109, 0.03355627, 0.089913, 
    0.1118221, 0.1924067, 0.03670564, 0.03394552, 0.0809755, 0.2031432, 
    0.272118, 0.3410078, 0.2153772, 0.1962419, 0.2621573, 0.3108927, 
    0.2727019, 0.2341328, 0.07810923, 0.1091691, 0.1504432, 0.3257153, 
    0.3799621, 0.4319243, 0.2991195, 0.1360348, 0.1891465,
  0.1781923, 0.2679893, 0.207643, 0.1502206, 0.1716693, 0.1713645, 0.1426666, 
    0.1091296, 0.07079297, 0.02681668, 0.03344922, 0.06092694, 0.1289856, 
    0.1833165, 0.3775211, 0.3343058, 0.3328055, 0.3350835, 0.1983232, 
    0.04045998, 0.1288094, 0.1818026, 0.1901668, 0.2201279, 0.449054, 
    0.1241346, 0.1189721, 0.150922, 0.191145,
  0.295163, 0.1637584, 0.266799, 0.2139214, 0.1891476, 0.1327722, 0.1301938, 
    0.1181651, 0.1996059, 0.2147077, 0.2156648, 0.2675382, 0.2260283, 
    0.2241967, 0.2137724, 0.1580819, 0.1535434, 0.134626, 0.1226273, 
    0.1706118, 0.1827045, 0.09764023, 0.1511193, 0.1383379, 0.07731579, 
    0.3434545, 0.1639682, 0.0974886, 0.3720073,
  0.3655233, 0.3742798, 0.3339924, 0.2266517, 0.3035814, 0.2571774, 
    0.2685649, 0.1887518, 0.2121706, 0.220264, 0.228714, 0.228211, 0.1993512, 
    0.2517937, 0.2932345, 0.2910141, 0.2441453, 0.1930985, 0.2351716, 
    0.2797653, 0.2656194, 0.2500422, 0.2320402, 0.258167, 0.156016, 
    0.2056277, 0.180614, 0.1594284, 0.3022436,
  0.4311221, 0.430769, 0.430416, 0.4300629, 0.4297099, 0.4293568, 0.4290038, 
    0.4261177, 0.4370939, 0.4480701, 0.4590463, 0.4700225, 0.4809987, 
    0.4919749, 0.5066972, 0.5014029, 0.4961086, 0.4908142, 0.4855199, 
    0.4802256, 0.4749313, 0.4639023, 0.4585735, 0.4532447, 0.4479159, 
    0.442587, 0.4372582, 0.4319294, 0.4314045,
  0.4172053, 0.483137, 0.4205296, 0.2825645, 0.1963496, 0.1917425, 0.2166423, 
    0.246266, 0.1008686, 0.1040104, 0.2309796, 0.3329837, 0.454487, 
    0.0234566, 0.1625441, 0.2754191, 0.2954242, 0.3451946, 0.2966167, 
    0.3807386, 0.7454897, 0.6969956, 0.3421527, 0.2366564, 0.2845089, 
    0.4612003, 0.356696, 0.2433904, 0.4605375,
  0.2324661, 0.1635582, 0.2468398, 0.1124213, 0.1988129, 0.1994146, 
    0.07914379, 0.3607703, 0.3399532, 0.3231026, 0.2060038, 0.09654059, 
    0.1477585, 0.1833125, 0.3327416, 0.4605579, 0.3659547, 0.3870494, 
    0.4363386, 0.4926021, 0.4771604, 0.5293442, 0.4627731, 0.4374421, 
    0.3708993, 0.3023205, 0.294367, 0.3049065, 0.3338313,
  0.351156, 0.2935, 0.2595654, 0.3038985, 0.3072258, 0.3350752, 0.3214995, 
    0.3024226, 0.3146667, 0.2975689, 0.3112232, 0.3730279, 0.4761544, 
    0.3579277, 0.324057, 0.3740982, 0.3887547, 0.415587, 0.4355289, 
    0.3888095, 0.374345, 0.3751436, 0.3420446, 0.2579322, 0.3391269, 
    0.3919375, 0.416716, 0.3255217, 0.3119833,
  0.3224472, 0.3620134, 0.3754706, 0.2958187, 0.3182448, 0.3527796, 
    0.3281159, 0.2773649, 0.2976734, 0.2894881, 0.2627532, 0.2795892, 
    0.2016446, 0.203289, 0.1573073, 0.1756276, 0.2407242, 0.2772181, 
    0.2946458, 0.2907021, 0.2611064, 0.2664817, 0.2456913, 0.1769982, 
    0.1031998, 0.1815627, 0.2237266, 0.3162336, 0.3398934,
  0.2585474, 0.1755628, 0.11494, 0.1420341, 0.1809038, 0.1710416, 0.1327014, 
    0.1647271, 0.1804948, 0.1476679, 0.05997753, 0.04323341, 0.01053141, 
    0.05112345, 0.3206156, 0.1382716, 0.1788602, 0.160706, 0.1278805, 
    0.178728, 0.2081977, 0.1469141, 0.1044337, 0.3047457, 0.03092764, 
    0.07927701, 0.09719604, 0.1723848, 0.2662659,
  0.06081219, 0.08119964, 0.007971096, 0.03756732, 0.05678898, 0.04813028, 
    0.06697579, 0.04995583, 0.04725821, 0.01535445, 0.01670937, 
    -2.300478e-05, 0.008422145, 0.01927729, 0.03115793, 0.06908546, 
    0.04941558, 0.06623565, 0.1089217, 0.05710798, 0.06106801, 0.02493348, 
    0.02875837, 0.04709832, 0.06186718, 0.05303774, 0.05660437, 0.04080768, 
    0.05010857,
  0.1091706, -0.0004496141, -2.24835e-06, 0.01274186, 0.004885789, 0.0262768, 
    0.01860939, 0.03207885, 0.03130819, 0.0004850477, 9.307891e-06, 
    3.543531e-05, 0.009861179, 0.02900788, 0.02177136, 0.02089307, 0.0176923, 
    0.02168458, 0.004094174, 0.008353858, 0.002004085, 0.009137076, 
    0.03863185, 0.1531048, 0.04480346, 0.06539419, 0.007932094, 0.001488075, 
    0.009899662,
  0.1519623, 0.06732085, 0.0142827, 0.09901232, 0.01695479, 0.01206035, 
    0.01745936, 0.01458246, 0.02046642, 0.003327269, 0.03431415, 0.01132151, 
    0.06133984, 0.01251523, 0.01718942, 0.008078246, 0.006053992, 
    0.006036332, 0.006112282, 0.006289535, 0.008734668, 0.01102686, 
    0.1190854, 0.009468034, 0.02928311, 0.0001734759, 0.01196535, 
    0.005061957, 0.02695983,
  0.03074317, 0.01010961, 0.0009513185, 0.02172745, 0.007357015, 0.007672617, 
    0.008055221, 0.005033616, 0.04655543, 0.05116318, 0.0180661, 0.01427318, 
    0.02024631, 0.02025866, 0.008347935, 0.01352593, 0.04888291, 0.05553333, 
    0.08139957, 0.1897415, 0.09263194, 0.1158714, 0.2557994, 0.04678451, 
    0.04009713, 0.01914177, 0.04509183, 0.02247356, 0.03490616,
  4.400546e-05, -4.213684e-07, 1.135062e-07, 0.008449148, 0.02057051, 
    0.01174197, 0.02250261, 0.01276319, 0.002445485, 0.01709479, 0.01321239, 
    0.009600487, 0.02111581, 0.01805039, 0.01194651, 0.009665742, 0.0201108, 
    0.02488455, 0.05061114, 0.04109585, 0.02014186, 0.003022508, 0.2803181, 
    0.08425608, 0.007572377, 0.01484971, 0.08411886, 0.1531186, 0.0001338618,
  3.673009e-07, 1.189233e-07, 1.931567e-08, 0.0007804697, 4.414619e-05, 
    0.005558377, -2.182192e-05, 0.004228805, 5.96227e-05, 0.2314492, 
    0.09520256, 0.03227218, 0.01470238, 0.003064503, 0.001202253, 
    0.001913329, 0.008200716, 0.01815488, 0.09342265, 0.0830396, 0.004043587, 
    0.06644616, 0.004851645, 0.006605499, 0.007388005, 0.02242266, 
    0.05953956, 0.04318337, 3.611214e-07,
  -8.496406e-08, 0.007314907, 0.01149793, 0.003037245, 0.02376632, 
    0.00173188, -0.001278059, -0.0003837256, 0.04897299, 0.2086657, 0.220265, 
    0.1960283, 0.2812367, 0.240235, 0.120506, 0.1649936, 0.1773164, 
    0.09708792, 0.1036032, 0.09058665, 0.004785377, 0.1611154, 0.03915139, 
    0.06206884, 0.05309553, 0.06241673, 0.04139951, 0.05397739, 0.01940386,
  0.001908102, 0.002795629, 0.03476119, 0.1480153, 0.01737213, 4.18666e-05, 
    0.1208287, 0.005915508, 0.006948082, 0.03293517, 0.09098082, 0.08156839, 
    0.1497932, 0.1697848, 0.1843197, 0.2207405, 0.2657802, 0.1870911, 
    0.2233468, 0.1431335, 0.05368384, 0.1224142, 0.1284823, 0.1969245, 
    0.2396009, 0.1415422, 0.139527, 0.1457068, 0.1000281,
  0.1198411, 0.1679056, 0.05039269, 0.05953036, 0.05497173, 0.06086172, 
    0.08827382, 0.1587538, 0.0291898, 0.03141734, 0.07338464, 0.1904707, 
    0.2282103, 0.3012114, 0.166463, 0.1631011, 0.2405989, 0.300505, 
    0.2513778, 0.2239157, 0.0711768, 0.1044814, 0.1265717, 0.2973974, 
    0.3505893, 0.3876724, 0.2802619, 0.1234236, 0.1697803,
  0.150684, 0.2688206, 0.187332, 0.1380741, 0.1877683, 0.1457579, 0.1405424, 
    0.08015367, 0.0506085, 0.01838342, 0.02029965, 0.03590029, 0.0958847, 
    0.1248591, 0.282952, 0.3445304, 0.3050246, 0.3127789, 0.1447815, 
    0.04720596, 0.1189454, 0.1584028, 0.1733047, 0.2175668, 0.3563234, 
    0.1229143, 0.0910553, 0.1006889, 0.1469411,
  0.2675382, 0.1359305, 0.2598886, 0.2007082, 0.2137205, 0.1551808, 
    0.1309452, 0.1041607, 0.168702, 0.2082386, 0.1984434, 0.2673187, 
    0.2260978, 0.2384642, 0.2575333, 0.2029575, 0.2034744, 0.1501679, 
    0.1222018, 0.229278, 0.2127925, 0.1189821, 0.1406856, 0.1574918, 
    0.09028955, 0.3532934, 0.1769495, 0.05822442, 0.3107067,
  0.4259995, 0.4019032, 0.3514798, 0.2911786, 0.3461184, 0.3009193, 0.303515, 
    0.2201779, 0.2213047, 0.2638881, 0.2656232, 0.2639876, 0.2298517, 
    0.2975754, 0.3274876, 0.3642626, 0.3029499, 0.2409941, 0.2676482, 
    0.32515, 0.2860847, 0.2450907, 0.2473371, 0.2860911, 0.1381406, 
    0.2247773, 0.1828812, 0.1372762, 0.314396,
  0.2510103, 0.2432043, 0.2353983, 0.2275922, 0.2197862, 0.2119802, 
    0.2041742, 0.2052775, 0.2222821, 0.2392868, 0.2562914, 0.273296, 
    0.2903006, 0.3073052, 0.3521826, 0.3543286, 0.3564747, 0.3586207, 
    0.3607668, 0.3629128, 0.3650589, 0.3997136, 0.3883689, 0.3770243, 
    0.3656797, 0.354335, 0.3429904, 0.3316457, 0.2572551,
  0.419997, 0.4692469, 0.3524196, 0.24401, 0.1766679, 0.1677214, 0.1905968, 
    0.216959, 0.1111716, 0.07695076, 0.1584847, 0.2931671, 0.4975619, 
    0.008579236, 0.1987243, 0.306878, 0.3549394, 0.3296958, 0.2716714, 
    0.3977748, 0.7682034, 0.7340505, 0.3005137, 0.2153527, 0.3088074, 
    0.4724182, 0.3553112, 0.2129578, 0.4348154,
  0.1760458, 0.1104022, 0.2333329, 0.07192162, 0.1663939, 0.1940171, 
    0.03843296, 0.325814, 0.3213792, 0.2945192, 0.1767139, 0.1024852, 
    0.1332081, 0.1463601, 0.2927935, 0.4078521, 0.3076524, 0.3229086, 
    0.3817138, 0.4420127, 0.436136, 0.5160264, 0.4361565, 0.4260372, 
    0.357671, 0.3197607, 0.3176194, 0.2484786, 0.3177279,
  0.2825145, 0.2442631, 0.2180429, 0.2651742, 0.2680793, 0.2811105, 
    0.2661871, 0.2544791, 0.2649307, 0.2438118, 0.266976, 0.3299937, 
    0.4383765, 0.3258889, 0.2865566, 0.3413289, 0.3556201, 0.4173263, 
    0.4075048, 0.346127, 0.3359801, 0.3454988, 0.2887971, 0.2280589, 
    0.3025263, 0.3642319, 0.3582716, 0.2884531, 0.281146,
  0.300801, 0.3465225, 0.3489554, 0.2736284, 0.3081039, 0.3300384, 0.3027283, 
    0.2359271, 0.2520058, 0.2549692, 0.2194193, 0.2326205, 0.1617685, 
    0.1693127, 0.1269775, 0.1429506, 0.2049095, 0.2685996, 0.2647766, 
    0.2491984, 0.2335925, 0.2351816, 0.2077288, 0.1490028, 0.07708895, 
    0.1389296, 0.2104701, 0.287068, 0.3205873,
  0.2127288, 0.1146265, 0.0741099, 0.1119865, 0.1445324, 0.1338058, 
    0.09495923, 0.1352789, 0.1217132, 0.1218152, 0.04293429, 0.02448765, 
    0.006648493, 0.03486096, 0.2818741, 0.1100325, 0.1624729, 0.1294142, 
    0.09010623, 0.1548269, 0.1769465, 0.1007952, 0.06326523, 0.307168, 
    0.0222726, 0.05740322, 0.07516895, 0.1291654, 0.2203567,
  0.02541028, 0.04803766, 0.006404067, 0.01440854, 0.0234783, 0.0206668, 
    0.04032061, 0.02083972, 0.02537393, 0.01107197, 0.008327129, 
    -4.190292e-06, 0.009643277, 0.01018984, 0.04167179, 0.03405284, 
    0.03664733, 0.0391406, 0.0779546, 0.03023349, 0.03382438, 0.01406461, 
    0.01087199, 0.03682479, 0.05204346, 0.02953323, 0.04039414, 0.01460358, 
    0.02135316,
  0.05856838, 8.703992e-07, -4.26551e-05, 0.004301635, -0.001473721, 
    0.009930953, 0.006811651, 0.01425047, 0.01032587, 6.583791e-05, 
    2.609874e-06, 1.12228e-05, 0.003137301, 0.008809838, 0.009483845, 
    0.006747563, 0.00351788, 0.0104677, 0.000673337, 0.002701933, 
    0.0006944342, 0.003363982, 0.01414941, 0.08528534, 0.03006721, 
    0.05400056, 0.002506565, 0.0002122364, 0.003357286,
  0.05988241, 0.04166301, 0.01585264, 0.08351378, 0.006853402, 0.002895605, 
    0.005551141, 0.003274008, 0.007450253, -0.0006849705, 0.02547014, 
    0.004420836, 0.04208537, 0.00313581, 0.005987629, 0.003894853, 
    0.001059538, 0.001954378, 0.002370767, 0.002110336, 0.00299017, 
    0.003618872, 0.04435125, 0.01054277, 0.02695778, 5.903597e-05, 
    0.003965585, 0.00208227, 0.01013786,
  0.008651514, 0.01635598, 0.0008326391, 0.01778708, 0.002278192, 
    0.002932392, 0.002818796, 0.00158535, 0.03819632, 0.03757887, 
    0.005853828, 0.003628736, 0.01001779, 0.0123678, 0.001388024, 
    0.003111267, 0.008291272, 0.009184066, 0.0158136, 0.03388777, 0.03315523, 
    0.0315897, 0.2299917, 0.04433741, 0.0340132, 0.01123133, 0.01598565, 
    0.005999126, 0.007040107,
  3.29514e-05, -2.339612e-07, -6.836387e-08, 0.006381553, 0.02214161, 
    0.005045637, 0.005332485, 0.005337517, 0.000375692, 0.006908668, 
    0.003723094, 0.002118837, 0.005382601, 0.006764824, 0.004257486, 
    0.006808314, 0.009282889, 0.006168506, 0.01739101, 0.01172058, 
    0.008476078, 0.001009442, 0.2094329, 0.07537218, 0.004028413, 
    0.005745702, 0.03276197, 0.05910565, 0.0001499895,
  3.36261e-07, 1.110024e-07, 1.909498e-08, 0.000422626, -1.790056e-06, 
    0.00103233, -1.93104e-05, 0.00117223, 3.22457e-05, 0.09672461, 
    0.02651918, 0.01111298, 0.003599267, 0.0004797936, 0.0002339233, 
    0.0004741858, 0.003137042, 0.006127996, 0.03458469, 0.04257396, 
    0.01228652, 0.05648031, 0.0008169169, 0.004330717, 0.002032107, 
    0.01478576, 0.03256669, 0.01581857, 3.00438e-07,
  -2.860755e-06, 0.005428073, 0.008987911, 0.002897523, 0.01780971, 
    0.001173087, -0.001234233, -0.0004173605, 0.04198768, 0.1778822, 
    0.2022023, 0.1839545, 0.2712745, 0.1816135, 0.08758286, 0.1115881, 
    0.09229695, 0.04474592, 0.04974077, 0.07718098, 0.003132064, 0.1553701, 
    0.03024063, 0.04870263, 0.03917304, 0.04499533, 0.01520994, 0.02908288, 
    0.02351553,
  0.001106236, 0.0007150723, 0.02293145, 0.1562445, 0.01672603, 1.712939e-05, 
    0.1066105, 0.004189353, 0.005737312, 0.03184759, 0.0874918, 0.07739912, 
    0.1253709, 0.1626726, 0.1683348, 0.1998232, 0.2522796, 0.1730657, 
    0.1617703, 0.1339401, 0.04818468, 0.113863, 0.1028503, 0.1850687, 
    0.1806167, 0.0932514, 0.08499867, 0.08773698, 0.07813585,
  0.09037825, 0.1395596, 0.03625014, 0.04687552, 0.06692924, 0.04674412, 
    0.06678064, 0.1287906, 0.02075347, 0.02472981, 0.06756552, 0.1725166, 
    0.1900025, 0.2478218, 0.1299954, 0.133495, 0.2245267, 0.2662207, 
    0.2098863, 0.2164702, 0.05847768, 0.09000632, 0.1083646, 0.2744249, 
    0.3172521, 0.3498727, 0.2410734, 0.1011454, 0.1417783,
  0.1134503, 0.2618799, 0.1646453, 0.1289393, 0.1778003, 0.1255976, 0.117842, 
    0.06057049, 0.04031904, 0.01491209, 0.01381982, 0.02100768, 0.08219041, 
    0.08732003, 0.2275899, 0.3520011, 0.2731855, 0.2842491, 0.09203674, 
    0.04652692, 0.1000378, 0.1381201, 0.1559697, 0.2121576, 0.3130074, 
    0.09857519, 0.0741751, 0.07304794, 0.1162578,
  0.2247676, 0.1108956, 0.2403296, 0.1733502, 0.2048687, 0.1653633, 
    0.1092242, 0.09364508, 0.1331434, 0.1855643, 0.1842723, 0.2337664, 
    0.2312118, 0.2756444, 0.2856373, 0.2700566, 0.2656955, 0.1518417, 
    0.1581521, 0.2373305, 0.2177639, 0.1414294, 0.1273717, 0.1888302, 
    0.1022732, 0.3413363, 0.1797034, 0.03333361, 0.2752131,
  0.4824502, 0.3991459, 0.3749534, 0.354167, 0.346635, 0.3404182, 0.3385538, 
    0.2745787, 0.2221382, 0.300707, 0.2965395, 0.3117231, 0.290206, 
    0.3432369, 0.3650013, 0.4342574, 0.3710236, 0.2988875, 0.3109736, 
    0.3463404, 0.3293417, 0.2224093, 0.2502542, 0.311103, 0.1294426, 
    0.2146553, 0.1615922, 0.1368357, 0.3257086,
  0.1602143, 0.1569353, 0.1536563, 0.1503773, 0.1470983, 0.1438194, 
    0.1405404, 0.1321622, 0.1429152, 0.1536682, 0.1644211, 0.175174, 
    0.185927, 0.1966799, 0.2301065, 0.2344088, 0.2387112, 0.2430135, 
    0.2473158, 0.2516182, 0.2559205, 0.2355768, 0.2238005, 0.2120242, 
    0.2002479, 0.1884716, 0.1766953, 0.164919, 0.1628375,
  0.4020688, 0.3819865, 0.2631294, 0.1470344, 0.1342824, 0.1347411, 
    0.1221008, 0.1604665, 0.09204195, 0.06284178, 0.07034846, 0.2702767, 
    0.4645431, 0.003758878, 0.2682856, 0.395977, 0.389266, 0.3300713, 
    0.2385638, 0.3845276, 0.7657965, 0.7672221, 0.2516176, 0.1952418, 
    0.359272, 0.5025379, 0.3348243, 0.1844152, 0.3815597,
  0.135211, 0.07413548, 0.1889892, 0.04300567, 0.1360349, 0.1828163, 
    0.02583959, 0.2680585, 0.3000803, 0.2533171, 0.1571884, 0.102608, 
    0.1042711, 0.1163942, 0.2446301, 0.3465632, 0.2309368, 0.2554581, 
    0.3187642, 0.3794886, 0.3780836, 0.4630201, 0.402383, 0.4138427, 
    0.3292924, 0.3228937, 0.3430592, 0.19188, 0.277487,
  0.2224734, 0.1952223, 0.1682909, 0.2112204, 0.2008412, 0.2175298, 
    0.2162051, 0.199764, 0.2157807, 0.1959037, 0.2238882, 0.2787946, 
    0.374332, 0.2746467, 0.2232532, 0.2798689, 0.3022759, 0.3767905, 
    0.3495411, 0.2813809, 0.2920257, 0.294481, 0.2459169, 0.1764114, 
    0.2699632, 0.3186918, 0.2945123, 0.2315349, 0.2255663,
  0.2527198, 0.2903419, 0.2937635, 0.2233356, 0.2599832, 0.2664016, 
    0.2573472, 0.1816327, 0.1954361, 0.1993536, 0.1665772, 0.1797734, 
    0.1181303, 0.1281543, 0.101356, 0.1063565, 0.1651026, 0.2119296, 
    0.2121887, 0.208793, 0.1869487, 0.1844966, 0.1690468, 0.1245646, 
    0.058077, 0.105137, 0.1813629, 0.2541895, 0.2734629,
  0.1584884, 0.06719137, 0.04643456, 0.08121146, 0.1038198, 0.08407302, 
    0.06679861, 0.1036158, 0.082435, 0.09426218, 0.0296598, 0.01652412, 
    0.004899718, 0.02320824, 0.2458701, 0.08001122, 0.1187237, 0.1033378, 
    0.0605543, 0.1262342, 0.1432497, 0.08372989, 0.03932521, 0.2922089, 
    0.01443556, 0.04118014, 0.05270278, 0.08886634, 0.1780385,
  0.01116976, 0.02388318, 0.006448695, 0.005575862, 0.01115386, 0.009666731, 
    0.02208717, 0.01340048, 0.01410671, 0.00716552, 0.006471632, 
    -1.399419e-06, 0.01070332, 0.006209012, 0.03213198, 0.01669678, 
    0.02406112, 0.02144277, 0.04072345, 0.01372143, 0.01839414, 0.00738377, 
    0.005580256, 0.02369196, 0.04691358, 0.01500633, 0.02211181, 0.00507684, 
    0.009349711,
  0.02960228, -3.773011e-05, 2.322896e-05, 0.002052264, -0.001811069, 
    0.00377033, 0.001764177, 0.006571602, 0.00342067, 3.255063e-05, 
    9.969575e-07, 5.02758e-06, 0.00133161, 0.004619825, 0.004576907, 
    0.001733036, 0.0008680511, 0.004621081, 0.0001586922, 0.001610471, 
    0.0003624248, 0.001917989, 0.00753452, 0.04149291, 0.01920731, 
    0.04389349, 0.0009813223, 9.231014e-05, 0.001661805,
  0.02989558, 0.02777079, 0.02253829, 0.06310068, 0.004336524, 0.001279694, 
    0.001846761, 0.001080258, 0.002634829, -0.0006308024, 0.01725363, 
    0.001537362, 0.02266238, 0.001335074, 0.002611588, 0.001826287, 
    0.000479564, 0.0008081696, 0.001327325, 0.001138404, 0.001597631, 
    0.00175379, 0.02301103, 0.00792975, 0.02791161, 3.584131e-05, 
    0.0006197494, 0.001121668, 0.00530494,
  0.004426429, 0.02653345, 0.0004777471, 0.01149076, 0.001167364, 0.00162356, 
    0.001524112, 0.0008634783, 0.03282601, 0.03334102, 0.003701421, 
    0.001716261, 0.005641847, 0.006158321, 0.0004747295, 0.001371127, 
    0.003287519, 0.003414939, 0.00658651, 0.0128852, 0.006943448, 
    0.008414309, 0.1048749, 0.04975782, 0.03245659, 0.004861769, 0.009237093, 
    0.002918886, 0.002643532,
  2.141321e-05, -8.064471e-08, -7.055227e-09, 0.007719037, 0.01725222, 
    0.002926077, 0.001407246, 0.003097842, 0.0001456556, 0.003434164, 
    0.0008022732, 0.0008639758, 0.0009426869, 0.002009089, 0.001404554, 
    0.003235778, 0.003477187, 0.002067671, 0.004477006, 0.004256484, 
    0.003629882, 0.0006064887, 0.137443, 0.06325015, 0.001956472, 
    0.003080126, 0.01675973, 0.02941767, 6.615488e-05,
  3.177264e-07, 1.056534e-07, 1.882883e-08, 4.104469e-05, 4.784994e-05, 
    0.000376943, -3.122359e-05, 0.0004240733, 1.826243e-05, 0.03731334, 
    0.01048389, 0.003600887, 0.001061256, 0.0001827858, 0.0001259564, 
    0.0002583664, 0.001167152, 0.00245347, 0.01847409, 0.02598515, 0.0103897, 
    0.04392061, 0.0002802123, 0.002637815, 0.0008524061, 0.008154311, 
    0.01852045, 0.008886199, 2.806253e-07,
  -2.108902e-06, 0.003740355, 0.004907716, 0.00181048, 0.01220471, 
    0.0008602947, -0.001213836, -0.0004114595, 0.034527, 0.1341434, 0.173149, 
    0.1476171, 0.2029251, 0.1250824, 0.06581332, 0.05659266, 0.05985222, 
    0.02279096, 0.02888519, 0.06234239, 0.002557022, 0.1365493, 0.02373846, 
    0.03338657, 0.02960381, 0.02689233, 0.007730256, 0.01499485, 0.01700734,
  0.0007553568, 0.0001035532, 0.01204279, 0.1482446, 0.03397691, 
    2.158818e-05, 0.08939413, 0.003302304, 0.004374186, 0.03018511, 
    0.0825518, 0.07549913, 0.1053865, 0.1336834, 0.1370616, 0.1639878, 
    0.2079321, 0.1468634, 0.1089514, 0.1191373, 0.04119595, 0.1049011, 
    0.0803262, 0.172367, 0.1274436, 0.0585041, 0.04399154, 0.05385027, 
    0.05452483,
  0.07007079, 0.1136694, 0.02360194, 0.03299285, 0.06404162, 0.03279681, 
    0.05188078, 0.1039063, 0.0160037, 0.01896222, 0.06019348, 0.1515197, 
    0.156249, 0.1899591, 0.09841531, 0.1136963, 0.1980341, 0.2106012, 
    0.1644192, 0.2032807, 0.04804521, 0.06830862, 0.08859907, 0.2540768, 
    0.2829665, 0.3596593, 0.1908465, 0.07768664, 0.09685734,
  0.09019273, 0.2400455, 0.1414662, 0.1173082, 0.1626092, 0.1105125, 
    0.09756899, 0.04837389, 0.03013587, 0.01235534, 0.01049526, 0.01554866, 
    0.08362526, 0.05645882, 0.1883066, 0.3279382, 0.2405707, 0.2454745, 
    0.05801035, 0.04243669, 0.0863214, 0.1344637, 0.1563741, 0.1999322, 
    0.2698027, 0.07767896, 0.05230503, 0.05363832, 0.09474149,
  0.1758279, 0.08411095, 0.2239865, 0.1422995, 0.1910216, 0.1554922, 
    0.09499243, 0.07810768, 0.1009922, 0.1455943, 0.1620887, 0.2007407, 
    0.22232, 0.296805, 0.2597229, 0.3190668, 0.2459618, 0.1673744, 0.1908097, 
    0.2393497, 0.2543165, 0.1469394, 0.1166471, 0.2018766, 0.1312036, 
    0.3148829, 0.1907331, 0.01513097, 0.2473761,
  0.5304244, 0.409942, 0.3922286, 0.3712891, 0.3507617, 0.3512916, 0.3857351, 
    0.3170854, 0.2354861, 0.311619, 0.3084844, 0.327581, 0.3553904, 
    0.3970079, 0.4288966, 0.4766568, 0.4263802, 0.3654374, 0.3096262, 
    0.3526044, 0.3755664, 0.210378, 0.2325898, 0.3383305, 0.1289551, 
    0.1914968, 0.1321271, 0.126171, 0.3002582,
  0.1208695, 0.1163119, 0.1117542, 0.1071966, 0.1026389, 0.09808125, 
    0.09352359, 0.08261435, 0.08919197, 0.09576958, 0.1023472, 0.1089248, 
    0.1155024, 0.12208, 0.1419175, 0.149038, 0.1561585, 0.163279, 0.1703995, 
    0.17752, 0.1846405, 0.180618, 0.1714776, 0.1623371, 0.1531966, 0.1440562, 
    0.1349157, 0.1257752, 0.1245156,
  0.4181328, 0.3334733, 0.1719195, 0.1124668, 0.1012778, 0.08288434, 
    0.08437779, 0.07346115, 0.05894122, 0.07700115, 0.0690958, 0.2037583, 
    0.3410468, 0.000309784, 0.3416625, 0.4642295, 0.4173457, 0.3253541, 
    0.2005742, 0.365175, 0.7656491, 0.8066629, 0.217218, 0.1692366, 
    0.3879674, 0.5332624, 0.3201013, 0.1672291, 0.3467269,
  0.1114745, 0.05501617, 0.1482808, 0.02321974, 0.1020598, 0.165875, 
    0.02192741, 0.2096149, 0.2558143, 0.2001727, 0.1330059, 0.09649037, 
    0.07066305, 0.1013693, 0.2023263, 0.2885679, 0.1745632, 0.1988591, 
    0.2461256, 0.3020461, 0.3071657, 0.3906241, 0.3469737, 0.3930065, 
    0.2985145, 0.3169482, 0.3033549, 0.1419032, 0.2592258,
  0.1655624, 0.1475577, 0.126227, 0.1573421, 0.1445411, 0.1631273, 0.1558858, 
    0.145323, 0.1675192, 0.1470415, 0.1784944, 0.2211339, 0.2966139, 
    0.2077029, 0.1554773, 0.2147688, 0.2315892, 0.3041156, 0.278466, 
    0.2214069, 0.2298785, 0.2209013, 0.1849492, 0.1239119, 0.2260889, 
    0.2663687, 0.2364158, 0.1782624, 0.1707103,
  0.1926038, 0.2321877, 0.2252056, 0.1717033, 0.2011286, 0.2090598, 0.210437, 
    0.1361743, 0.1388489, 0.1409192, 0.1163431, 0.1227244, 0.07598606, 
    0.08496971, 0.07434675, 0.07562564, 0.1184365, 0.1526022, 0.1485074, 
    0.153527, 0.1461045, 0.1313619, 0.1252715, 0.1016672, 0.03795354, 
    0.07283577, 0.1396171, 0.2096864, 0.2201578,
  0.1095109, 0.03782213, 0.03034939, 0.05223399, 0.06516598, 0.05110089, 
    0.04624332, 0.07240787, 0.04746851, 0.06347383, 0.01754039, 0.009708636, 
    0.003427057, 0.01341401, 0.2096274, 0.05378208, 0.06771043, 0.07241448, 
    0.03730209, 0.09066558, 0.1013065, 0.06439772, 0.02355817, 0.2632991, 
    0.00901513, 0.02645402, 0.03470902, 0.05266379, 0.1207106,
  0.007002776, 0.01419226, 0.007623171, 0.002973804, 0.006055797, 
    0.004614209, 0.009206755, 0.007312493, 0.008002255, 0.003905087, 
    0.006690452, -6.085675e-07, 0.01287484, 0.003602022, 0.01919432, 
    0.007057578, 0.01397392, 0.01240793, 0.02275427, 0.006963331, 
    0.008576644, 0.003792579, 0.003577088, 0.01637422, 0.038096, 0.006523275, 
    0.01053917, 0.002314433, 0.004757741,
  0.01814099, -0.0001289568, -2.997825e-05, 0.001226587, -0.00134387, 
    0.0008521396, 0.0005921488, 0.002745121, 0.001456485, 2.300135e-05, 
    1.280352e-07, 2.148563e-06, 0.0007597921, 0.003048567, 0.002532679, 
    0.0006394591, 0.0004268119, 0.001938527, 8.345024e-05, 0.001025761, 
    0.0002303519, 0.001304232, 0.004961343, 0.02638668, 0.01218988, 
    0.03554853, 0.0005413679, 5.584825e-05, 0.001029675,
  0.01838315, 0.01557174, 0.0209315, 0.05372835, 0.002467479, 0.0006735823, 
    0.0007477065, 0.000520873, 0.001016403, -0.0003051322, 0.01034433, 
    0.0004601606, 0.009238675, 0.0006689795, 0.0009915542, 0.0006968546, 
    0.0003053647, 0.0003646908, 0.0008767855, 0.0007559945, 0.001039745, 
    0.001065025, 0.01467524, 0.007149739, 0.02930495, 2.036972e-05, 
    -0.0001907102, 0.0007213749, 0.003396618,
  0.002372502, 0.02716044, 0.0003368384, 0.006974936, 0.0007282334, 
    0.001061866, 0.0009951864, 0.0005601925, 0.02351835, 0.03538079, 
    0.002187929, 0.001056248, 0.002698819, 0.002820181, 0.000214048, 
    0.0008021175, 0.001927056, 0.001916238, 0.003946329, 0.007462445, 
    0.002592613, 0.004586052, 0.05034949, 0.05444839, 0.03286283, 0.00200859, 
    0.004619984, 0.001617273, 0.001480769,
  1.47049e-05, 7.909375e-08, 2.186441e-08, 0.01130118, 0.0101332, 
    0.001987304, -7.847091e-06, 0.002107792, 9.919591e-05, 0.001748591, 
    0.0004740728, 0.0004812234, 0.000427124, 0.0006329922, 0.0004618404, 
    0.001564035, 0.001168473, 0.001022414, 0.001964053, 0.00222292, 
    0.001528011, 0.0004394596, 0.09796892, 0.05179524, 0.0008839692, 
    0.001991877, 0.01058869, 0.01784891, -4.012929e-06,
  3.083929e-07, 1.028616e-07, 1.796669e-08, 1.065289e-05, -1.322995e-07, 
    0.000204124, -1.941969e-05, 0.0001687558, 2.00883e-05, 0.01224759, 
    0.005118, 0.001672314, 0.0005794001, 0.0001182862, 8.221631e-05, 
    0.0001692418, 0.0005766712, 0.001195018, 0.01217551, 0.01827029, 
    0.005021183, 0.03543608, 0.0001801607, 0.0008578936, 0.0005456597, 
    0.004225432, 0.01202727, 0.005969111, 2.723351e-07,
  -7.230701e-07, 0.002584628, 0.002689466, 0.001207118, 0.008511405, 
    0.0004773563, -0.001142422, -0.000486875, 0.03062799, 0.0886042, 
    0.1402614, 0.09527475, 0.1269018, 0.07608364, 0.04305789, 0.03785541, 
    0.04021376, 0.01364419, 0.01847966, 0.04776147, 0.002241987, 0.1126205, 
    0.01796398, 0.01785612, 0.02041705, 0.01656524, 0.004284273, 0.00935025, 
    0.01303516,
  0.0006205711, 3.532018e-05, 0.005912471, 0.1334271, 0.03334485, 
    2.882696e-05, 0.07580965, 0.00273219, 0.003081669, 0.02664335, 
    0.07426791, 0.06535769, 0.08350471, 0.1075548, 0.1013458, 0.1222829, 
    0.1588282, 0.1087199, 0.06733229, 0.1008175, 0.0356176, 0.09176247, 
    0.06140997, 0.1595225, 0.08734489, 0.03314259, 0.02449844, 0.03266491, 
    0.03851776,
  0.04959752, 0.08879352, 0.01636748, 0.02222168, 0.06009623, 0.02400425, 
    0.04069559, 0.08564562, 0.01219292, 0.01436665, 0.05060256, 0.1246598, 
    0.1298929, 0.1440046, 0.07490918, 0.08532003, 0.1525546, 0.1483307, 
    0.1096474, 0.1894443, 0.03774437, 0.05390472, 0.07374787, 0.2283531, 
    0.2546336, 0.3566773, 0.1472875, 0.05109123, 0.05788642,
  0.05937427, 0.2091237, 0.1212732, 0.1030017, 0.1477586, 0.09411378, 
    0.08080612, 0.03490822, 0.02077168, 0.009612797, 0.008173863, 0.01844834, 
    0.08812615, 0.03860547, 0.1490099, 0.2931981, 0.2140054, 0.2071118, 
    0.0446766, 0.03631039, 0.07463585, 0.1314251, 0.1515885, 0.2005927, 
    0.2238936, 0.05997058, 0.03263926, 0.03911192, 0.07638933,
  0.1370815, 0.06078403, 0.2113976, 0.1101665, 0.1759112, 0.1476897, 
    0.1185511, 0.08069416, 0.09302753, 0.147693, 0.1468915, 0.1595428, 
    0.2003036, 0.2493478, 0.2042553, 0.2838293, 0.2184282, 0.164527, 
    0.2364959, 0.22751, 0.2520812, 0.1583722, 0.1131988, 0.2275735, 
    0.1520924, 0.2726716, 0.1903463, 0.004899499, 0.2051886,
  0.5238638, 0.3608993, 0.358197, 0.3382096, 0.331497, 0.3579178, 0.3600182, 
    0.2924073, 0.2609932, 0.2888501, 0.3172331, 0.3035948, 0.3441971, 
    0.4105259, 0.4062007, 0.4409037, 0.3680153, 0.3391596, 0.3162115, 
    0.3414332, 0.3550504, 0.1722513, 0.2209242, 0.3404874, 0.1074292, 
    0.1673722, 0.1048485, 0.1085444, 0.2610266,
  0.1059829, 0.1047484, 0.1035138, 0.1022792, 0.1010447, 0.09981009, 
    0.09857552, 0.09775895, 0.1017718, 0.1057846, 0.1097975, 0.1138103, 
    0.1178232, 0.121836, 0.1215862, 0.1258921, 0.1301981, 0.134504, 
    0.1388099, 0.1431159, 0.1474218, 0.1493327, 0.1422485, 0.1351643, 
    0.1280801, 0.1209959, 0.1139117, 0.1068275, 0.1069706,
  0.3799014, 0.2447051, 0.09331179, 0.03296395, 0.03962377, 0.06019806, 
    0.04238541, 0.03126459, 0.02384824, 0.07113112, 0.06552026, 0.1530973, 
    0.2925013, -0.002379873, 0.3818809, 0.4503408, 0.4194722, 0.324532, 
    0.1638376, 0.3829153, 0.759545, 0.8241966, 0.2026491, 0.1532074, 
    0.3718065, 0.544347, 0.2963898, 0.1506444, 0.3638448,
  0.1005808, 0.04579761, 0.1230746, 0.01605003, 0.08150895, 0.144602, 
    0.0187382, 0.1804745, 0.2288176, 0.1601982, 0.1153596, 0.08970256, 
    0.05320177, 0.08776347, 0.1770612, 0.2462233, 0.1432892, 0.1662372, 
    0.1964223, 0.2457508, 0.2601356, 0.3260782, 0.3138445, 0.3727949, 
    0.2543176, 0.2897998, 0.2731079, 0.1105994, 0.2457638,
  0.1301322, 0.1180067, 0.09943819, 0.1248936, 0.1105378, 0.1314116, 
    0.1236279, 0.1119969, 0.1330051, 0.1178637, 0.1483631, 0.17761, 
    0.2454781, 0.1648352, 0.1150076, 0.1706372, 0.1878621, 0.2478222, 
    0.2293819, 0.1824385, 0.1789114, 0.1628632, 0.1381742, 0.09121315, 
    0.1878347, 0.2219429, 0.1895225, 0.146035, 0.1358353,
  0.1570239, 0.1912788, 0.179276, 0.1353124, 0.1602407, 0.1709447, 0.1765969, 
    0.1066009, 0.1067318, 0.1023873, 0.08331195, 0.08601086, 0.05186042, 
    0.05766922, 0.05561423, 0.05464758, 0.08533163, 0.1055407, 0.1025446, 
    0.1138206, 0.1130519, 0.09206934, 0.09001642, 0.0897468, 0.02352178, 
    0.05059195, 0.1093742, 0.1657293, 0.1883644,
  0.07825215, 0.02421428, 0.02048411, 0.03198308, 0.03989176, 0.03088804, 
    0.03303305, 0.04592029, 0.02899179, 0.04096069, 0.008620461, 0.007107448, 
    0.002491797, 0.007882286, 0.1858295, 0.03494171, 0.04035711, 0.04626974, 
    0.02380697, 0.06050889, 0.06599799, 0.04513442, 0.01414762, 0.2373564, 
    0.006061597, 0.01676491, 0.0226325, 0.03214915, 0.08418396,
  0.005198351, 0.01015333, 0.008479672, 0.002034204, 0.003357688, 
    0.002386286, 0.004402606, 0.004635008, 0.005261513, 0.002385661, 
    0.003914912, -3.984615e-07, 0.0112534, 0.002052038, 0.01426845, 
    0.003884796, 0.007967584, 0.007130741, 0.01297797, 0.003883814, 
    0.004219264, 0.002089963, 0.00264572, 0.01233933, 0.02949088, 
    0.003314487, 0.005041377, 0.001334461, 0.00326138,
  0.01318775, -0.0001505249, -5.401935e-05, 0.0008707019, -0.000868315, 
    0.0004103286, 0.0003174451, 0.001338228, 0.0009343622, 1.719015e-05, 
    3.850446e-08, -2.348914e-07, 0.0005259857, 0.001812881, 0.001239436, 
    0.0003434171, 0.0003132451, 0.001027307, 6.573502e-05, 0.0007087205, 
    0.0001665096, 0.0009900599, 0.003715817, 0.01946509, 0.01077589, 
    0.03344656, 0.0003846349, 3.977153e-05, 0.0007394615,
  0.01310332, 0.008329336, 0.02029514, 0.05035031, 0.001406548, 0.0004403999, 
    0.0004217945, 0.0002502709, 0.000488728, -0.0002570528, 0.006969145, 
    0.0002038424, 0.004456033, 0.0004137992, 0.0004382859, 0.0003077575, 
    0.0002261033, 0.0002355103, 0.0006532278, 0.0005678597, 0.0007654461, 
    0.0007560173, 0.01069488, 0.007790543, 0.02461705, 7.0795e-05, 
    -0.0002892162, 0.0005280528, 0.002487051,
  0.001370994, 0.02063447, 0.0005557016, 0.00471311, 0.0005194397, 
    0.0007738844, 0.0007307413, 0.0003914005, 0.01772628, 0.03978732, 
    0.001084691, 0.0007553284, 0.001259268, 0.001239301, 0.0001418293, 
    0.0005528237, 0.001339324, 0.00130534, 0.002750679, 0.005200819, 
    0.001480791, 0.003184277, 0.03111919, 0.04169195, 0.02660077, 
    0.0009268652, 0.002259906, 0.0009461234, 0.001030416,
  1.136267e-05, 1.195983e-07, 2.687655e-08, 0.01035105, 0.006284263, 
    0.001513862, -0.0009393668, 0.001595116, 4.474045e-05, 0.001093547, 
    0.0003676763, 0.0003404873, 0.0002586917, 0.0002578958, 0.000217832, 
    0.0007485227, 0.0004979564, 0.0006884555, 0.001270822, 0.001453773, 
    0.0007386204, 0.0003358815, 0.0646958, 0.03725246, 0.0003678064, 
    0.001460022, 0.007691284, 0.01271353, 0.0006271083,
  3.038987e-07, 9.89944e-08, 1.682386e-08, 8.157755e-06, 6.405405e-07, 
    0.0001351297, -1.579654e-05, 0.0001043939, 0.0001240683, 0.006546015, 
    0.003081047, 0.001028823, 0.0004074488, 8.796901e-05, 6.122096e-05, 
    0.0001269586, 0.0003464319, 0.0007303372, 0.009114822, 0.01422491, 
    0.00279753, 0.03052732, 0.0001422688, -0.0001315349, 0.0004154388, 
    0.002078264, 0.008953012, 0.004504073, 2.671391e-07,
  -2.545991e-08, 0.001681795, 0.001896185, 0.0007832405, 0.007197037, 
    0.0004353744, -0.001106151, -0.0008841486, 0.03090789, 0.05836866, 
    0.1047056, 0.05806595, 0.07904053, 0.04830841, 0.02811737, 0.02648311, 
    0.02666495, 0.009531948, 0.01248134, 0.03173859, 0.002090919, 0.09474114, 
    0.01535147, 0.007939085, 0.01210617, 0.01015311, 0.002923349, 
    0.006136422, 0.01002884,
  0.0004005638, 3.646484e-05, 0.003279648, 0.1274379, 0.02913819, 
    3.523238e-05, 0.06736168, 0.002412594, 0.002152282, 0.02225646, 
    0.06653006, 0.05021725, 0.06695498, 0.08800597, 0.07789894, 0.09199287, 
    0.1195964, 0.07350506, 0.04420493, 0.08566572, 0.03182524, 0.08051098, 
    0.04654285, 0.1488746, 0.06272571, 0.01908299, 0.01580312, 0.02075264, 
    0.02806327,
  0.03451766, 0.07153884, 0.01245961, 0.01469713, 0.05477059, 0.01913006, 
    0.03358559, 0.07494662, 0.01031755, 0.0121291, 0.04574725, 0.1049111, 
    0.1050327, 0.1132544, 0.06093878, 0.06552806, 0.1161365, 0.1095013, 
    0.07179992, 0.1781544, 0.03190111, 0.04575419, 0.06891874, 0.20541, 
    0.234619, 0.3416836, 0.111053, 0.03639204, 0.03665221,
  0.03484471, 0.1889253, 0.1107713, 0.105827, 0.1408798, 0.08639319, 
    0.07280861, 0.03051012, 0.01697781, 0.00876826, 0.006570519, 0.04889008, 
    0.1167573, 0.03291149, 0.126403, 0.2495942, 0.2010527, 0.1794423, 
    0.05113763, 0.03192969, 0.06617165, 0.1279057, 0.1296873, 0.2166161, 
    0.1892979, 0.04708347, 0.02307006, 0.02974518, 0.06396919,
  0.1069938, 0.04608147, 0.2057851, 0.08489861, 0.1784153, 0.1427595, 
    0.1707012, 0.1176943, 0.1206088, 0.1700308, 0.1510108, 0.1387849, 
    0.2221841, 0.1961888, 0.1650733, 0.2212494, 0.203329, 0.1502756, 
    0.2508984, 0.194998, 0.2378435, 0.1593456, 0.1643257, 0.2415969, 
    0.1731173, 0.2384388, 0.1859856, 0.004259925, 0.1710213,
  0.4933484, 0.3244442, 0.298907, 0.2978674, 0.3047106, 0.3124895, 0.2976617, 
    0.2340062, 0.2160085, 0.1913732, 0.233057, 0.2347765, 0.2436413, 
    0.300189, 0.3057169, 0.3103071, 0.2573028, 0.2492108, 0.2301489, 
    0.2577502, 0.273004, 0.1406252, 0.2028655, 0.3617401, 0.09752692, 
    0.1294024, 0.08964597, 0.09154323, 0.2103257,
  0.1007678, 0.09941874, 0.0980697, 0.09672066, 0.09537162, 0.09402258, 
    0.09267354, 0.0770104, 0.08021492, 0.08341943, 0.08662395, 0.08982847, 
    0.09303299, 0.0962375, 0.1031563, 0.1074838, 0.1118114, 0.1161389, 
    0.1204664, 0.124794, 0.1291215, 0.1326955, 0.1265125, 0.1203295, 
    0.1141465, 0.1079635, 0.1017805, 0.09559745, 0.101847,
  0.2902082, 0.1730684, 0.03476106, 0.02589571, 0.01196291, 0.04293023, 
    0.01885831, 0.007285872, 0.01536353, 0.06357899, 0.05730775, 0.1340585, 
    0.2786989, -0.00106286, 0.3782467, 0.4096398, 0.405888, 0.3385249, 
    0.1547559, 0.3889696, 0.7622882, 0.8129612, 0.2091628, 0.151241, 
    0.3111113, 0.5274608, 0.2979581, 0.1552819, 0.3391421,
  0.1040673, 0.04131776, 0.1107324, 0.01394904, 0.06305451, 0.1304484, 
    0.01681913, 0.1692458, 0.2125832, 0.1488516, 0.1081331, 0.0852083, 
    0.04690703, 0.08036548, 0.1665148, 0.2220196, 0.1284533, 0.1491843, 
    0.1689093, 0.2163293, 0.2335477, 0.2914086, 0.2865236, 0.3471212, 
    0.2269078, 0.2664123, 0.2573, 0.09729107, 0.2233614,
  0.1109, 0.1025867, 0.08457984, 0.1078162, 0.09376888, 0.1148565, 0.1074391, 
    0.09436105, 0.114442, 0.1017457, 0.1290053, 0.1505675, 0.2114785, 
    0.1389805, 0.09557514, 0.1436706, 0.158682, 0.213349, 0.1933615, 
    0.1552319, 0.1494401, 0.1315028, 0.1122759, 0.07638476, 0.1566681, 
    0.1919597, 0.1613665, 0.1280465, 0.1187703,
  0.1353994, 0.1588778, 0.1520068, 0.1130759, 0.1354963, 0.1423739, 0.148922, 
    0.09025612, 0.08903582, 0.08526912, 0.06556613, 0.0677898, 0.03950131, 
    0.04478747, 0.04496835, 0.04314282, 0.06725232, 0.0785322, 0.07609851, 
    0.08972194, 0.0905167, 0.0709205, 0.06937475, 0.1054276, 0.01710208, 
    0.03920018, 0.08921021, 0.1372342, 0.1587975,
  0.05754675, 0.01847368, 0.01489813, 0.02083695, 0.02710317, 0.02146073, 
    0.02419833, 0.03067686, 0.02033218, 0.02848647, 0.005794506, 0.005902533, 
    0.001808311, 0.005168199, 0.1909412, 0.02289578, 0.02753658, 0.03271539, 
    0.01662863, 0.04169093, 0.04566362, 0.03178217, 0.009796877, 0.2374557, 
    0.004004228, 0.01153393, 0.01491751, 0.02273428, 0.06243332,
  0.00428688, 0.008210672, 0.0152511, 0.001656718, 0.002486777, 0.001731021, 
    0.002829937, 0.003478517, 0.00403649, 0.001849395, 0.002284156, 
    -3.012548e-07, 0.01432131, 0.001428181, 0.008337971, 0.002887723, 
    0.005039511, 0.003999958, 0.008405478, 0.002435968, 0.002399304, 
    0.001446401, 0.002185174, 0.009601532, 0.03955533, 0.002241543, 
    0.003179277, 0.001008976, 0.002649756,
  0.01063805, -8.056345e-05, -5.2257e-05, 0.000699734, -0.000860545, 
    0.0002885834, 0.0002289289, 0.0009475206, 0.0007365664, 1.430849e-05, 
    2.900869e-08, -2.50199e-05, 0.0004170961, 0.001113808, 0.0007697442, 
    0.0002554894, 0.000261037, 0.0007013684, 5.61471e-05, 0.0005469009, 
    0.0001348307, 0.0008248324, 0.003084253, 0.01585451, 0.03098946, 
    0.05770158, 0.0003119114, 3.225559e-05, 0.0006053433,
  0.01060786, 0.006153525, 0.01931377, 0.07769553, 0.0009628284, 
    0.0003435213, 0.0003186085, 0.0001690384, 0.0003249429, -0.0004003296, 
    0.005518299, 0.0001434151, 0.003099918, 0.0003165741, 0.0002780056, 
    0.000200732, 0.0001850067, 0.0001818359, 0.0005429453, 0.0004742155, 
    0.0006315792, 0.0006153703, 0.008758762, 0.03524104, 0.05206616, 
    0.005466482, -0.0002295152, 0.0004244756, 0.002053408,
  0.0009994364, 0.02283137, 0.003845043, 0.004874927, 0.0004150118, 
    0.0006278452, 0.000580661, 0.0003176256, 0.02290291, 0.06946665, 
    0.0007603852, 0.0006113401, 0.0007675803, 0.0007648568, 9.36928e-05, 
    0.0004350983, 0.001048392, 0.001014308, 0.002192019, 0.004075861, 
    0.001083931, 0.002502971, 0.02273527, 0.04219206, 0.07954903, 
    0.000558854, 0.001327651, 0.0006903832, 0.0008199326,
  0.0004830933, -9.5498e-07, 2.710437e-08, 0.01563211, 0.004329332, 
    0.001264665, -0.0001550062, 0.001291696, -9.97168e-05, 0.0008219058, 
    0.0002546907, 0.0002758572, 0.0001997795, 0.0001700991, 0.0001526502, 
    0.0004764872, 0.0003267513, 0.000549249, 0.001005914, 0.001146945, 
    0.0005031189, 0.000284603, 0.07820795, 0.03384476, 0.0002171254, 
    0.001213633, 0.00630934, 0.01022627, 0.01476506,
  3.035673e-07, 9.81679e-08, 1.620829e-08, 6.768371e-06, -2.908538e-06, 
    0.0001021964, -1.105353e-05, 8.823178e-05, 0.001564293, 0.00346719, 
    0.002289711, 0.0007505876, 0.0003305623, 6.772111e-05, 5.201305e-05, 
    0.0001088998, 0.0002750263, 0.0005475241, 0.007606189, 0.01208589, 
    0.001770227, 0.02950495, 0.0001228999, -0.0004907912, 0.0003530711, 
    0.001407996, 0.007403351, 0.003773163, 2.665458e-07,
  2.307532e-07, 0.001313081, 0.001806824, 0.0005192485, 0.007992103, 
    0.0003663139, -0.001168494, -0.001406383, 0.03929188, 0.04684834, 
    0.07195677, 0.03786057, 0.05440538, 0.03428537, 0.01961066, 0.01953338, 
    0.01909057, 0.007258441, 0.009702834, 0.0227346, 0.001720074, 0.09787617, 
    0.04099105, 0.00431912, 0.007859788, 0.006742591, 0.002245026, 
    0.004330479, 0.007586733,
  0.0004155636, -0.0001488925, 0.002189321, 0.1237878, 0.02596659, 
    3.164363e-05, 0.06141855, 0.002178677, 0.001694149, 0.01899796, 
    0.06836142, 0.03832223, 0.05779056, 0.06909671, 0.06287398, 0.07320394, 
    0.09116066, 0.05479881, 0.03255295, 0.07886793, 0.02931677, 0.0743423, 
    0.04048368, 0.1325857, 0.05078328, 0.01279894, 0.01192188, 0.01595508, 
    0.02262298,
  0.02734055, 0.06472202, 0.01157989, 0.01106693, 0.05080113, 0.01657098, 
    0.03078263, 0.08758923, 0.01028023, 0.01475583, 0.05045824, 0.1063556, 
    0.08998513, 0.09649524, 0.0522762, 0.05454925, 0.09713241, 0.08851145, 
    0.05340726, 0.1914806, 0.03054141, 0.04403134, 0.07292645, 0.2090429, 
    0.2291613, 0.2980043, 0.0858121, 0.0278226, 0.02713128,
  0.02216247, 0.2005025, 0.1181715, 0.1300569, 0.186998, 0.09796473, 
    0.07353418, 0.03690167, 0.0204483, 0.01326921, 0.009494391, 0.1810413, 
    0.19339, 0.03672451, 0.1135403, 0.2325695, 0.2294779, 0.1655067, 
    0.08415791, 0.0359972, 0.07025177, 0.1506289, 0.1131976, 0.2593058, 
    0.1668512, 0.04097638, 0.01839561, 0.02508309, 0.05639062,
  0.08791055, 0.03944527, 0.2318883, 0.06722077, 0.1941462, 0.1384125, 
    0.2638465, 0.2189335, 0.2178092, 0.2298532, 0.2100258, 0.1635319, 
    0.2998068, 0.1770474, 0.1608007, 0.1883611, 0.2418245, 0.1597312, 
    0.2789573, 0.1833004, 0.2453934, 0.1717395, 0.2511945, 0.2642806, 
    0.1737473, 0.2123905, 0.2156325, 0.01026024, 0.1458172,
  0.4524424, 0.3003705, 0.2606999, 0.2700784, 0.2815727, 0.2770325, 
    0.2592614, 0.1955801, 0.1753634, 0.1415376, 0.1736689, 0.1741069, 
    0.1747921, 0.2240742, 0.2154257, 0.2357837, 0.1946664, 0.2022599, 
    0.1827142, 0.2005518, 0.2083176, 0.1324219, 0.2055629, 0.3863648, 
    0.09010232, 0.1075913, 0.08617607, 0.08727498, 0.1888603 ;

 average_DT = 730 ;

 average_T1 = 106 ;

 average_T2 = 836 ;

 climatology_bounds =
  106, 836 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
