netcdf reduced_ocean_monthly_1x1deg.199301-199712.sos {
dimensions:
	lat = 2 ;
	bnds = 2 ;
	lon = 2 ;
	time = UNLIMITED ; // (2 currently)
variables:
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	float sos(time, lat, lon) ;
		sos:_FillValue = 1.e+20f ;
		sos:missing_value = 1.e+20f ;
		sos:units = "psu" ;
		sos:long_name = "Sea Surface Salinity" ;
		sos:cell_methods = "area:mean yh:mean xh:mean time: mean" ;
		sos:cell_measures = "area: areacello" ;
		sos:standard_name = "sea_surface_salinity" ;
		sos:interp_method = "conserve_order1" ;
	double time(time) ;
		time:units = "days since 1958-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 1958-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "om5_b05_noHiLatHenyey_55" ;
		:associated_files = "areacello: 19930101.ocean_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Mon Jun 17 18:57:22 2024" ;
		:hostname = "pp337" ;
		:history = "Tue Oct 22 11:05:33 2024: ncks --dmn lat,0,1 --dmn lon,0,1 --dmn time,0,1 ocean_monthly_1x1deg.199301-199712.sos.nc -o reduced_ocean_monthly_1x1deg.199301-199712.sos.nc\n",
			"fregrid --standard_dimension --input_mosaic ocean_mosaic.nc --input_file all --interp_method conserve_order1 --remap_file .fregrid_remap_file_360_by_180.nc --nlon 360 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file out.nc" ;
		:external_variables = "areacello" ;
		:NCO = "netCDF Operators version 5.1.5 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
}
