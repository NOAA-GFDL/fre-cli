netcdf tracer_level.0002-0002.radon {
dimensions:
	bnds = 2 ;
	lat = 2 ;
	lon = 2 ;
	pfull = 65 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	float radon(time, pfull, lat, lon) ;
		radon:_FillValue = -1.e+10f ;
		radon:missing_value = -1.e+10f ;
		radon:units = "vmr*1e21" ;
		radon:long_name = "radon-222" ;
		radon:interp_method = "conserve_order1" ;
		radon:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 17:15:31 2024" ;
		:hostname = "pp329" ;
		:history = "Tue Sep 23 14:27:36 2025: ncks -d lon,0,1 tracer_level.0002-0002.radon.nc_lat01 tracer_level.0002-0002.radon.nc_lat01_lon01\n",
			"Tue Sep 23 14:26:18 2025: ncks -d lat,0,1 tracer_level.0002-0002.radon.nc tracer_level.0002-0002.radon.nc_lat01\n",
			"Tue Aug 12 16:31:13 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0002-0002.radon.nc reduced/tracer_level.0002-0002.radon.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00020101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.3.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5 ;

 lat_bnds =
  -90, -89,
  -80, -79 ;

 lon = 0.625, 13.125 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 radon =
  5.84339e-21, 5.84339e-21,
  1.198741e-20, 1.299412e-20,
  1.185919e-20, 1.185919e-20,
  2.707962e-20, 2.905326e-20,
  3.511195e-20, 3.511195e-20,
  6.797557e-20, 7.752918e-20,
  1.002282e-19, 1.002282e-19,
  1.787181e-19, 1.90655e-19,
  2.568689e-19, 2.568689e-19,
  3.396632e-19, 4.168067e-19,
  6.702528e-19, 6.702528e-19,
  5.990152e-19, 7.488989e-19,
  2.00547e-18, 2.00547e-18,
  1.299381e-18, 1.545818e-18,
  5.258524e-18, 5.258524e-18,
  3.388956e-18, 3.675393e-18,
  1.187743e-17, 1.187743e-17,
  1.118741e-17, 1.088408e-17,
  2.72789e-17, 2.72789e-17,
  3.127639e-17, 3.732474e-17,
  6.386993e-17, 6.386993e-17,
  5.399635e-17, 6.145649e-17,
  2.272603e-16, 2.272603e-16,
  1.596789e-16, 1.650774e-16,
  9.672524e-16, 9.672524e-16,
  8.529583e-16, 7.466007e-16,
  4.591861e-15, 4.591861e-15,
  6.189363e-15, 4.978484e-15,
  1.61205e-14, 1.61205e-14,
  2.657154e-14, 2.419917e-14,
  5.170192e-14, 5.170192e-14,
  9.461897e-14, 9.876561e-14,
  8.748715e-14, 8.748715e-14,
  2.660231e-13, 2.979323e-13,
  1.323306e-13, 1.323306e-13,
  5.338106e-13, 6.930059e-13,
  3.53954e-13, 3.53954e-13,
  1.325008e-12, 1.546789e-12,
  1.563455e-12, 1.563455e-12,
  5.538631e-12, 5.603272e-12,
  8.223117e-12, 8.223117e-12,
  1.895778e-11, 2.092674e-11,
  5.810028e-11, 5.810028e-11,
  7.823552e-11, 9.149771e-11,
  3.209372e-10, 3.209372e-10,
  4.049505e-10, 4.375319e-10,
  1.591832e-09, 1.591832e-09,
  2.469798e-09, 2.333356e-09,
  8.500012e-09, 8.500012e-09,
  1.236298e-08, 1.171917e-08,
  5.857941e-08, 5.857941e-08,
  6.779644e-08, 6.766712e-08,
  3.12504e-07, 3.12504e-07,
  3.301741e-07, 3.471152e-07,
  1.958516e-06, 1.958516e-06,
  1.62583e-06, 1.74109e-06,
  8.129346e-06, 8.129346e-06,
  7.850933e-06, 8.773354e-06,
  3.785294e-05, 3.785294e-05,
  3.667513e-05, 3.924871e-05,
  0.00016837, 0.00016837,
  0.000165512, 0.0001391753,
  0.001031774, 0.001031774,
  0.001068673, 0.001042599,
  0.007043442, 0.007043442,
  0.006093835, 0.00683558,
  0.02378623, 0.02378623,
  0.01572161, 0.01846066,
  0.04555744, 0.04555744,
  0.03094472, 0.03610782,
  0.07273281, 0.07273281,
  0.05700063, 0.06288863,
  0.1068113, 0.1068113,
  0.1022332, 0.1058445,
  0.154615, 0.154615,
  0.1742871, 0.1678025,
  0.2110141, 0.2110141,
  0.2683745, 0.242781,
  0.2746139, 0.2746139,
  0.3727483, 0.3279251,
  0.3400338, 0.3400338,
  0.461947, 0.4135256,
  0.3937578, 0.3937578,
  0.5203037, 0.4807975,
  0.4325204, 0.4325204,
  0.5530845, 0.5221275,
  0.4566895, 0.4566895,
  0.5711287, 0.5427616,
  0.4699539, 0.4699539,
  0.5839799, 0.5554429,
  0.4766698, 0.4766698,
  0.5926505, 0.5604157,
  0.4749982, 0.4749982,
  0.5966731, 0.5570363,
  0.4701429, 0.4701429,
  0.5956888, 0.5484015,
  0.4624002, 0.4624002,
  0.5916227, 0.5404015,
  0.451346, 0.451346,
  0.5824398, 0.5350035,
  0.4358947, 0.4358947,
  0.5679162, 0.5242132,
  0.4166179, 0.4166179,
  0.5459655, 0.50828,
  0.3984487, 0.3984487,
  0.5189677, 0.4884913,
  0.3832363, 0.3832363,
  0.4899096, 0.4624029,
  0.3667257, 0.3667257,
  0.4574514, 0.4291912,
  0.3462757, 0.3462757,
  0.4236823, 0.3943839,
  0.3244964, 0.3244964,
  0.391773, 0.3641616,
  0.3042182, 0.3042182,
  0.3598081, 0.3389662,
  0.2848201, 0.2848201,
  0.328214, 0.3159839,
  0.2643491, 0.2643491,
  0.3016985, 0.293511,
  0.2442631, 0.2442631,
  0.2845521, 0.2755138,
  0.2307505, 0.2307505,
  0.2721483, 0.2620395,
  0.2229644, 0.2229644,
  0.2615055, 0.252426,
  0.2186493, 0.2186493,
  0.2546053, 0.2472809,
  0.216563, 0.216563,
  0.2524069, 0.2451792 ;

 time = 547.5 ;

 time_bnds =
  365, 730 ;
}
