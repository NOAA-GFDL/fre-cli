netcdf \00010101.ps.atmos_daily.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float hfls(time, grid_yt, grid_xt) ;
		hfls:_FillValue = 1.e+20f ;
		hfls:missing_value = 1.e+20f ;
		hfls:units = "W m-2" ;
		hfls:long_name = "Surface Upward Latent Heat Flux" ;
		hfls:cell_methods = "time: mean" ;
		hfls:cell_measures = "area: area" ;
		hfls:comment = "Lv*evap" ;
		hfls:time_avg_info = "average_T1,average_T2,average_DT" ;
		hfls:standard_name = "surface_upward_latent_heat_flux" ;
	float huss(time, grid_yt, grid_xt) ;
		huss:_FillValue = 1.e+20f ;
		huss:missing_value = 1.e+20f ;
		huss:units = "1.0" ;
		huss:long_name = "Near-Surface Specific Humidity" ;
		huss:cell_methods = "time: mean" ;
		huss:cell_measures = "area: area" ;
		huss:coordinates = "height2m" ;
		huss:time_avg_info = "average_T1,average_T2,average_DT" ;
		huss:standard_name = "specific_humidity" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:_FillValue = NaN ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float prw(time, grid_yt, grid_xt) ;
		prw:_FillValue = 1.e+20f ;
		prw:missing_value = 1.e+20f ;
		prw:units = "kg m-2" ;
		prw:long_name = "Water Vapor Path" ;
		prw:cell_methods = "time: mean" ;
		prw:cell_measures = "area: area" ;
		prw:time_avg_info = "average_T1,average_T2,average_DT" ;
		prw:standard_name = "atmosphere_water_vapor_content" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float rlut(time, grid_yt, grid_xt) ;
		rlut:_FillValue = 1.e+20f ;
		rlut:missing_value = 1.e+20f ;
		rlut:units = "W m-2" ;
		rlut:long_name = "TOA Outgoing Longwave Radiation" ;
		rlut:cell_methods = "time: mean" ;
		rlut:cell_measures = "area: area" ;
		rlut:time_avg_info = "average_T1,average_T2,average_DT" ;
		rlut:standard_name = "toa_outgoing_longwave_flux" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float sfcWind(time, grid_yt, grid_xt) ;
		sfcWind:_FillValue = 1.e+20f ;
		sfcWind:missing_value = 1.e+20f ;
		sfcWind:units = "m s-1" ;
		sfcWind:long_name = "Near-Surface Wind Speed" ;
		sfcWind:cell_methods = "time: mean" ;
		sfcWind:cell_measures = "area: area" ;
		sfcWind:coordinates = "height10m" ;
		sfcWind:time_avg_info = "average_T1,average_T2,average_DT" ;
		sfcWind:standard_name = "wind_speed" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float ts(time, grid_yt, grid_xt) ;
		ts:_FillValue = 1.e+20f ;
		ts:missing_value = 1.e+20f ;
		ts:units = "K" ;
		ts:long_name = "Surface Temperature" ;
		ts:cell_methods = "time: mean" ;
		ts:cell_measures = "area: area" ;
		ts:time_avg_info = "average_T1,average_T2,average_DT" ;
		ts:standard_name = "surface_temperature" ;
	float zg500(time, grid_yt, grid_xt) ;
		zg500:_FillValue = 1.e+20f ;
		zg500:missing_value = 1.e+20f ;
		zg500:units = "m" ;
		zg500:long_name = "Geopotential Height at 500 hPa" ;
		zg500:cell_methods = "time: mean" ;
		zg500:cell_measures = "area: area" ;
		zg500:time_avg_info = "average_T1,average_T2,average_DT" ;
		zg500:standard_name = "geopotential_height" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 hfls =
  29.90368, 49.35181, 49.9096, 95.12691, 71.87212, 35.03489, 47.63442, 
    50.20385, 53.5752, 11.16579, 14.51125, 27.03942, 11.70793, 14.27759, 
    -0.3786513,
  85.97427, 75.98698, 57.91388, 77.04918, 35.42171, 26.09041, 44.20863, 
    40.81323, 50.58518, 40.09371, 21.50808, 49.16239, 49.14007, 5.695109, 
    -0.3838496,
  77.86563, 86.58753, 82.07342, 79.01974, 63.59566, 5.253563, 42.06587, 
    43.8668, 50.82354, 48.50815, 47.83553, 52.98396, 56.59428, 50.79833, 
    23.60787,
  90.28301, 79.84243, 84.45894, 86.84377, 96.03311, 70.30258, 5.590069, 
    37.44505, 66.14964, 48.09973, 42.62407, 47.77813, 53.16575, 54.2935, 
    40.27913,
  108.1024, 96.88148, 87.83829, 87.85508, 89.05102, 96.91717, 82.45899, 
    7.665728, 23.434, 30.05699, 38.93267, 44.75055, 51.67457, 57.85662, 
    60.49834,
  111.5299, 111.7298, 101.9088, 96.64767, 93.89856, 92.98494, 86.36525, 
    85.89212, 63.87637, 54.17691, 35.88317, 47.81981, 51.35664, 57.47815, 
    59.41167,
  142.48, 126.0268, 119.2533, 111.6749, 106.4043, 106.0936, 105.7216, 
    104.1531, 96.93313, 94.34602, 76.10916, 52.9972, 54.02652, 56.78365, 
    56.2613,
  160.5278, 143.6519, 129.296, 121.3241, 115.8553, 113.2635, 111.5116, 
    110.4745, 105.2159, 105.8064, 92.3639, 59.81791, 54.64816, 56.76723, 
    56.20507,
  150.6531, 140.6597, 129.5796, 121.8886, 115.4403, 112.5857, 109.8309, 
    111.2056, 112.5377, 108.7657, 99.57213, 64.77615, 57.7329, 57.47926, 
    52.13752,
  130.8871, 124.7921, 120.3337, 114.0291, 108.5477, 105.3859, 107.403, 
    107.7126, 95.67406, 57.05529, 68.44485, 65.23853, 54.89882, 53.54874, 
    48.85418,
  19.94387, 68.18848, 35.11386, 77.19118, 53.91861, 27.53799, 39.91742, 
    39.15331, 30.5566, 8.709927, 6.694763, 16.43366, 8.347309, 7.020243, 
    -1.035404,
  94.01846, 63.43055, 68.16828, 77.42448, 37.32515, 15.14052, 46.80177, 
    45.37751, 38.44511, 26.12229, 12.31758, 26.77488, 30.09464, 3.41725, 
    -1.226893,
  136.9446, 119.7449, 95.17655, 95.66568, 65.04585, 2.645418, 37.6474, 
    49.59634, 51.96608, 34.23428, 30.95558, 31.09142, 29.64791, 30.73212, 
    12.87078,
  145.8134, 144.2041, 137.166, 121.9089, 106.4885, 69.11348, 2.082128, 
    35.04427, 61.74097, 39.09015, 32.89597, 32.47304, 30.65792, 26.59863, 
    21.80292,
  140.8575, 139.7991, 135.6308, 130.8493, 119.6519, 108.6756, 80.07188, 
    4.914348, 10.67877, 20.84244, 32.31161, 32.82687, 32.6984, 30.39337, 
    29.32289,
  136.3033, 136.7004, 131.5711, 129.3912, 126.5813, 120.7381, 109.4274, 
    104.0917, 68.36091, 65.57024, 27.8831, 33.6718, 33.63538, 33.11654, 
    30.79506,
  134.0072, 133.4505, 128.346, 124.3258, 121.1189, 119.2733, 115.7979, 
    110.9834, 103.5854, 110.1534, 65.93564, 35.3195, 34.24898, 35.51768, 
    34.48705,
  132.0383, 130.3293, 126.3854, 122.4379, 116.0227, 110.2302, 104.9459, 
    103.797, 107.2649, 115.0891, 82.69083, 37.3639, 35.0563, 36.77258, 
    35.45859,
  121.8291, 121.4803, 118.6989, 116.8132, 114.5379, 112.4398, 110.5155, 
    110.9144, 113.3944, 110.972, 87.62427, 38.8427, 35.22116, 36.03963, 
    32.42701,
  104.0649, 105.2761, 106.6556, 105.4754, 104.2499, 106.519, 111.2164, 
    111.2786, 96.00427, 57.59768, 61.20727, 38.20073, 33.92863, 33.76033, 
    30.82523,
  29.49665, 79.39426, 36.22445, 66.26254, 38.2092, 15.41371, 24.21033, 
    24.48758, 14.63505, 2.524331, 4.54463, 10.4499, 3.422899, 3.775796, 
    -1.475031,
  99.55483, 107.1141, 100.3814, 83.37931, 22.29678, 7.595412, 29.30658, 
    26.37353, 16.6594, 17.80875, 8.695395, 17.84048, 24.64693, 0.227561, 
    -1.737749,
  103.4131, 108.9124, 111.5458, 104.6378, 61.59361, 2.802226, 23.29206, 
    25.85521, 24.45564, 25.46906, 22.63697, 21.23371, 20.75711, 31.25564, 
    7.687753,
  107.2414, 108.6677, 114.9735, 118.6814, 115.5807, 58.64091, 2.099117, 
    19.09479, 31.21553, 24.77027, 22.57123, 22.27404, 20.89271, 18.62674, 
    19.85809,
  112.411, 112.5591, 115.7835, 123.7976, 127.4977, 104.6736, 57.6132, 
    4.565296, 4.721332, 12.36031, 22.25357, 24.86841, 23.59048, 22.24597, 
    20.97233,
  117.1093, 118.8862, 118.9836, 123.8579, 130.4616, 120.5527, 96.96727, 
    89.75337, 58.5301, 62.34965, 23.91878, 25.80862, 24.56903, 23.34992, 
    20.58767,
  125.197, 127.1145, 125.566, 126.8255, 129.7521, 124.0255, 112.465, 
    107.3583, 105.8252, 115.1535, 53.1879, 29.93278, 25.48637, 25.08777, 
    24.93339,
  129.218, 132.7282, 132.9009, 133.1095, 130.4518, 125.4616, 119.5993, 
    120.1405, 120.1186, 124.772, 67.88586, 32.96475, 27.17938, 27.13265, 
    25.45874,
  124.2681, 129.776, 132.8704, 134.642, 131.5636, 124.6623, 120.7146, 
    124.0693, 126.605, 123.8061, 79.37349, 35.25262, 30.18461, 28.38721, 
    25.50344,
  112.2394, 118.5169, 125.1055, 128.377, 128.4959, 124.6787, 121.5553, 
    118.413, 105.4979, 67.91891, 61.62674, 35.53001, 34.50707, 30.05908, 
    29.44142,
  30.186, 69.28781, 31.06088, 58.54395, 15.96561, 4.620884, 14.55353, 
    13.90488, 12.6291, 2.516629, 0.08817343, 6.27221, 2.267228, 1.925579, 
    -0.5842738,
  76.43607, 74.09801, 64.90688, 53.85924, 11.82014, 4.326458, 13.74294, 
    17.06936, 17.14952, 13.72735, 3.454065, 11.49145, 17.80231, 0.1519339, 
    -0.6532018,
  73.31511, 61.42937, 62.24793, 60.46941, 32.29095, 1.437121, 10.94933, 
    19.07415, 24.72638, 20.27587, 16.40111, 12.39819, 12.49832, 17.63468, 
    5.994524,
  64.27818, 56.91526, 64.82674, 67.00723, 61.38698, 29.21724, -0.9560582, 
    8.484658, 19.52128, 17.59842, 13.38289, 12.58552, 12.94139, 11.7723, 
    12.58611,
  56.88434, 59.40531, 66.11562, 66.77129, 60.15685, 59.47005, 60.73809, 
    1.913983, 1.959728, 6.339938, 11.84248, 14.41221, 14.31263, 14.03899, 
    13.24203,
  59.13514, 65.76833, 68.94794, 63.59967, 53.0408, 62.47777, 101.1762, 
    104.3756, 59.04048, 63.25182, 21.98762, 16.94074, 14.82189, 13.24846, 
    13.05468,
  66.43985, 72.16913, 71.20568, 58.61789, 47.93162, 69.23689, 102.617, 
    114.6154, 122.7928, 131.7735, 53.16456, 20.55632, 16.28527, 14.81254, 
    16.99631,
  79.22583, 78.72034, 75.36917, 57.70323, 59.79492, 86.53474, 116.2762, 
    126.0243, 133.4176, 134.9903, 52.05973, 22.9968, 16.82232, 18.68106, 
    18.8256,
  86.39959, 84.33742, 76.67826, 65.11486, 76.66173, 101.989, 121.4774, 
    122.6847, 127.7903, 127.3481, 59.16478, 25.83772, 18.96892, 22.60896, 
    17.56969,
  82.10811, 79.4471, 74.3224, 79.92526, 90.79325, 106.555, 119.7112, 
    119.0771, 104.7615, 64.15684, 44.37476, 26.20104, 26.78516, 22.69279, 
    21.8245,
  36.72674, 81.28628, 42.7725, 62.04868, 12.70072, 3.76093, 16.40561, 
    14.87112, 15.64011, 5.036236, 0.4752112, 5.133053, 1.451237, 1.659036, 
    -0.07729162,
  88.24762, 90.31697, 76.54839, 58.91077, 5.428793, 8.784087, 20.42345, 
    17.18258, 14.91925, 14.53654, 3.636008, 9.195682, 13.24052, 1.155654, 
    -0.03052879,
  88.41698, 79.50895, 65.36109, 62.22869, 44.06359, 2.832501, 18.19785, 
    20.30075, 18.67632, 14.73027, 14.26157, 10.05181, 8.753593, 9.843642, 
    4.233417,
  92.827, 76.27119, 64.16093, 74.79767, 95.81362, 61.10793, 0.7413305, 
    12.99763, 15.36454, 12.65689, 10.6776, 8.94291, 7.449193, 6.694005, 
    7.335553,
  95.04328, 78.2803, 68.45449, 77.66142, 92.79767, 103.6608, 88.86219, 
    1.818138, -0.8169997, 2.180555, 8.341966, 9.496581, 7.581588, 6.61267, 
    6.959939,
  97.1233, 83.79354, 73.23766, 77.5854, 85.7849, 96.5926, 115.8155, 103.431, 
    46.08648, 45.8288, 16.7435, 11.03699, 8.031536, 6.566501, 7.002732,
  103.468, 93.03603, 79.83617, 78.98044, 81.47308, 89.50407, 104.6459, 
    106.0877, 107.396, 114.6892, 45.79217, 14.09298, 8.311985, 6.690997, 
    7.770307,
  113.2272, 100.9135, 83.53759, 78.87901, 81.04982, 91.24094, 110.6284, 
    117.9091, 122.1383, 116.7452, 36.88425, 15.36965, 8.722073, 7.851161, 
    7.529326,
  114.955, 104.7511, 86.78647, 78.46326, 79.75532, 96.0891, 117.7008, 
    117.1062, 117.1589, 111.1448, 41.56239, 15.84196, 9.023249, 9.529157, 
    9.556837,
  106.1012, 91.87922, 78.07041, 76.89349, 82.38218, 96.99767, 118.4921, 
    113.6096, 96.60474, 51.79499, 31.48509, 14.90121, 11.94797, 13.33376, 
    13.79647,
  38.42847, 86.24054, 50.74516, 77.28505, 25.98875, 11.07192, 17.71925, 
    16.68664, 14.39678, 3.697607, 0.7760437, 2.277699, 0.2863366, 1.192304, 
    -0.3061956,
  94.83387, 101.8266, 99.5528, 89.31242, 18.1683, 8.21797, 20.72439, 
    15.52581, 10.16745, 8.871483, 2.075456, 6.024156, 8.96297, 0.6530478, 
    -0.07454053,
  98.64342, 100.9419, 102.7324, 100.4351, 63.25273, 1.982138, 16.34619, 
    15.96945, 10.27515, 9.143429, 6.998737, 5.765967, 7.795322, 9.332646, 
    2.92713,
  106.617, 103.0239, 101.8157, 104.8686, 115.3563, 69.49582, 2.71488, 
    7.231191, 8.275229, 6.174344, 4.700841, 4.115173, 4.105628, 6.653508, 
    5.375134,
  113.7324, 106.4996, 100.6247, 98.5798, 109.3904, 115.075, 88.72878, 
    2.340438, -0.6090736, 0.931077, 3.71731, 4.049097, 3.372426, 5.169108, 
    6.129706,
  121.4625, 108.6822, 98.70801, 92.25932, 101.9606, 109.7147, 112.195, 
    94.00412, 35.01019, 30.77778, 9.600596, 4.315543, 3.819422, 6.572888, 
    7.634212,
  132.5433, 113.4959, 98.57487, 89.82738, 96.96941, 102.0061, 100.4616, 
    95.8113, 84.82072, 81.96284, 29.51884, 5.482117, 3.663484, 6.211717, 
    8.228372,
  136.9637, 114.5358, 96.54081, 90.36079, 95.60961, 98.44691, 100.3844, 
    107.9918, 107.6623, 93.50208, 22.51789, 6.29215, 3.26133, 7.204817, 
    8.026834,
  130.8438, 110.3816, 94.72894, 89.33306, 93.2246, 95.40867, 99.18629, 
    103.9554, 103.4363, 88.22191, 23.56927, 6.958236, 4.935464, 7.890628, 
    10.04526,
  111.6337, 91.8197, 84.34911, 82.35535, 86.10698, 88.0366, 98.55688, 
    102.4768, 83.2356, 38.64003, 23.44515, 7.703847, 5.622465, 7.255063, 
    12.02281,
  32.50927, 81.45358, 43.80713, 71.60387, 12.81567, 6.982353, 9.667059, 
    7.020205, 7.605055, 0.5317229, -0.9479934, 1.495114, 0.8275149, 2.068601, 
    -0.3387798,
  91.1184, 97.6827, 103.4084, 94.75546, 16.56893, 6.65987, 11.51831, 
    7.545704, 6.14158, 6.75714, -0.07978026, 6.261873, 8.234672, 0.8442042, 
    -0.3063043,
  100.7904, 100.0999, 109.7211, 109.7658, 67.59688, 2.290895, 8.849565, 
    7.151902, 5.533168, 7.292179, 7.216505, 7.172476, 9.167984, 9.623001, 
    4.323376,
  110.2588, 106.229, 111.7948, 117.355, 115.0207, 66.79968, 3.239507, 
    2.227865, 3.637924, 4.219467, 4.993548, 4.54461, 6.620676, 7.630599, 
    6.571214,
  122.7285, 115.1463, 116.1139, 117.7818, 111.7654, 99.51218, 66.73161, 
    4.002596, 0.6218349, 1.272291, 3.841454, 5.166663, 5.290385, 9.149816, 
    6.353565,
  137.1347, 123.4726, 120.4826, 118.7013, 110.7266, 94.22355, 81.31451, 
    51.53695, 16.9724, 12.23622, 3.594113, 5.170259, 10.22675, 12.17357, 
    9.564744,
  149.1279, 133.3751, 127.4895, 121.1564, 111.2926, 94.67313, 79.86821, 
    58.64264, 45.60876, 39.25768, 13.85659, 5.801545, 10.11314, 12.16992, 
    12.24926,
  151.9458, 138.549, 130.919, 125.2543, 112.8746, 95.80505, 77.1086, 
    65.81042, 64.69772, 54.3854, 9.961553, 4.563283, 9.22791, 12.68642, 
    12.35505,
  137.3895, 135.6548, 132.2379, 127.1491, 113.7518, 94.57756, 73.16664, 
    59.55267, 62.97247, 53.91339, 9.757659, 3.515329, 7.934896, 13.90606, 
    15.25981,
  114.8731, 113.884, 118.5555, 116.9369, 104.844, 86.97745, 64.56825, 
    51.59933, 50.42272, 20.0403, 15.59557, 3.957745, 6.366655, 11.54648, 
    15.59239,
  30.18808, 84.62022, 43.47585, 63.60222, 9.003234, 2.140717, 6.241577, 
    6.751247, 9.361827, 1.787945, 0.5546011, 3.325044, 1.050202, 1.336251, 
    -0.3785072,
  89.2901, 107.056, 112.5555, 97.24577, 9.210705, 1.825709, 6.087929, 
    7.500794, 7.729077, 8.685429, 1.684649, 7.172385, 9.063536, 0.6593789, 
    -0.3660343,
  96.14007, 107.9689, 122.341, 111.2797, 57.71985, 0.8191461, 2.804862, 
    6.527435, 6.606506, 8.496464, 7.978731, 7.953539, 7.795706, 9.637957, 
    3.809421,
  97.4012, 109.3972, 120.3036, 116.0186, 100.9226, 51.7659, 2.197204, 
    1.652244, 5.18921, 5.277846, 5.755652, 5.979486, 6.740044, 6.920969, 
    6.015733,
  93.2859, 109.5849, 119.8859, 115.7827, 96.33742, 75.78777, 47.55151, 
    3.103341, 0.3949554, 0.6734973, 3.511671, 6.431262, 5.271238, 6.232954, 
    7.017113,
  89.23018, 109.4818, 117.9915, 111.6573, 95.82558, 76.7115, 59.08517, 
    33.2608, 14.47476, 13.9872, 3.431054, 6.833865, 6.161099, 7.151192, 
    5.899425,
  98.00774, 110.4625, 115.2062, 107.4661, 95.04036, 76.5915, 62.00294, 
    41.10871, 35.69903, 37.89821, 17.13119, 8.840962, 7.948787, 7.917403, 
    5.938035,
  105.9171, 107.6985, 109.5422, 104.3143, 95.82286, 77.88793, 62.95683, 
    48.22698, 46.18477, 48.10065, 13.29519, 10.88321, 10.55753, 10.07931, 
    7.368233,
  97.09384, 101.3303, 106.2748, 100.9473, 94.26534, 79.95941, 67.11412, 
    53.08924, 47.90296, 44.94852, 10.68196, 10.87008, 12.11396, 12.03743, 
    10.61857,
  88.62538, 88.4072, 91.07698, 90.8297, 86.56057, 75.29155, 68.15191, 
    58.31402, 44.30017, 20.33135, 18.17934, 10.54808, 12.98565, 13.729, 
    14.36697,
  24.57923, 87.54375, 45.5293, 68.36984, 10.51135, 3.388565, 8.643313, 
    7.343522, 8.642472, 1.565436, 0.1354226, 1.037474, 0.1093328, 0.3236986, 
    -0.7445637,
  66.03447, 107.1877, 130.8473, 120.37, 8.502699, 2.100133, 10.46188, 
    8.150336, 6.572431, 6.325274, 1.254235, 3.032681, 4.606669, 0.2559429, 
    -0.7981956,
  61.08755, 99.68035, 135.1019, 132.9292, 64.70701, -0.8013177, 7.425273, 
    8.847104, 7.398215, 5.81604, 5.07602, 3.267292, 3.568213, 5.569273, 
    1.46137,
  65.62801, 97.86332, 129.3069, 131.4884, 125.4186, 64.50034, 0.6746535, 
    2.226521, 4.782799, 4.206266, 3.163759, 2.478707, 2.421834, 3.53519, 
    2.52588,
  67.70213, 97.5533, 125.668, 124.2423, 112.4326, 105.0493, 67.44787, 
    1.951169, -0.355635, 0.6797235, 3.732384, 3.542207, 2.870119, 2.811302, 
    3.617533,
  68.72215, 99.01833, 120.6139, 114.9863, 103.4812, 93.47498, 90.98562, 
    66.36252, 21.0097, 14.88989, 5.896696, 5.54091, 3.250336, 2.695906, 
    3.472968,
  77.41035, 102.5833, 116.5281, 106.8948, 93.52341, 81.57275, 76.43265, 
    64.22813, 47.40879, 37.97075, 17.2997, 6.924463, 3.255536, 2.801549, 
    2.726642,
  76.54099, 101.5757, 110.2919, 100.1256, 87.11421, 74.26595, 66.52436, 
    60.61691, 64.39285, 57.56174, 11.91743, 7.315583, 3.450686, 2.664583, 
    2.325415,
  70.31889, 93.75163, 104.1219, 92.75918, 79.21854, 68.23678, 59.23326, 
    49.88986, 52.16423, 49.24265, 8.475417, 7.523419, 5.309663, 3.84711, 4.059,
  67.93323, 73.58688, 85.36782, 82.24178, 70.97454, 59.83671, 55.28371, 
    46.8718, 38.73386, 14.93961, 19.63724, 12.15921, 7.461158, 7.223077, 
    6.809978,
  26.47719, 85.46861, 31.56744, 40.74089, 7.722154, 2.261551, 5.036795, 
    4.349507, 7.859059, 0.5124635, -1.049118, -0.4210033, -0.5028114, 
    0.356695, -0.7079582,
  105.5777, 117.1837, 116.1522, 92.40034, 6.315258, 1.103365, 5.304066, 
    5.153759, 4.660228, 4.870198, -0.4541016, 1.545104, 4.368216, -0.3715715, 
    -1.419207,
  109.9012, 111.473, 120.6357, 108.7367, 51.29454, 0.3283034, 2.710755, 
    3.947121, 3.45694, 4.184247, 3.185236, 2.239609, 4.351305, 7.880531, 
    1.335079,
  109.5466, 110.2223, 113.0833, 104.9857, 98.38891, 51.20784, 1.804374, 
    1.058605, 1.724231, 1.663301, 1.35853, 0.8497254, 2.154696, 4.192729, 
    2.590097,
  108.4224, 107.4779, 107.7327, 98.52992, 88.61711, 76.47887, 46.60236, 
    2.728671, 0.5688186, 0.6144986, 0.6512331, 1.064924, 1.841826, 3.136277, 
    5.737541,
  106.1909, 104.7672, 102.5325, 91.69552, 85.74497, 73.91805, 61.00898, 
    39.89679, 9.986721, 6.454754, 2.626477, 1.669256, 1.443214, 3.198856, 
    5.099245,
  100.0508, 101.554, 100.0589, 89.2617, 81.37468, 70.13655, 61.33883, 
    47.35518, 30.81644, 20.66212, 8.993962, 2.462138, 1.733932, 3.318035, 
    6.65327,
  89.29751, 94.89266, 96.01482, 86.53867, 79.63798, 70.52106, 61.46402, 
    52.88126, 43.17549, 34.13777, 6.48778, 3.152555, 2.043488, 3.7796, 
    6.266811,
  75.13184, 84.42372, 92.91314, 83.94262, 74.71026, 65.95347, 58.05433, 
    51.62436, 46.49327, 33.88717, 4.542201, 4.52388, 1.71512, 3.46715, 
    5.833891,
  70.85905, 67.70951, 75.36549, 73.44813, 67.69289, 59.36004, 54.16603, 
    49.34906, 37.14367, 9.934594, 18.45495, 6.934974, 2.587228, 2.019352, 
    4.524894,
  18.78163, 52.77678, 14.90022, 14.59516, 5.93289, 0.9605854, 3.03368, 
    2.898131, 5.360455, -0.7691152, -1.395314, -0.5525165, 0.08213606, 
    0.6453346, -0.2734925,
  82.27737, 73.54359, 57.80042, 39.78855, 4.272964, 0.6006019, 2.471731, 
    3.74517, 3.173373, 2.207945, -1.644575, 1.952385, 4.281771, 0.05585356, 
    -1.083858,
  86.27838, 68.86145, 58.49443, 47.59401, 21.96551, 0.4693513, 1.189526, 
    2.880363, 3.071236, 2.178289, 0.5825414, 2.390519, 5.917029, 9.506378, 
    2.369711,
  87.53782, 68.60797, 57.92356, 45.58937, 40.29551, 24.07293, 1.390242, 
    0.5794807, 3.438195, 2.258563, 0.8166333, 1.460459, 3.351725, 5.83935, 
    3.906226,
  87.6755, 73.34155, 63.54002, 51.13981, 38.86657, 36.26987, 22.59074, 
    1.842122, 1.340012, 1.826331, 2.456657, 1.968187, 3.239811, 2.014405, 
    6.575009,
  97.17207, 84.75861, 74.2229, 61.23966, 47.24783, 32.87975, 32.20639, 
    31.69081, 7.027502, 5.677295, 2.993354, 3.910709, 3.601695, 2.348301, 
    5.274329,
  112.6707, 100.8946, 88.19744, 75.48951, 61.24736, 41.68485, 29.67625, 
    32.5138, 29.98355, 20.04575, 7.942853, 9.602835, 11.69892, 5.334942, 
    7.946824,
  118.1627, 111.0942, 99.89064, 86.17458, 70.8885, 55.67154, 41.00448, 
    34.87667, 40.8327, 30.91412, 6.064475, 8.9467, 11.96924, 10.02819, 
    12.53911,
  92.75445, 95.06287, 93.87996, 87.25611, 74.63335, 59.32275, 42.71797, 
    34.45713, 42.58983, 30.40879, 3.159762, 6.107217, 8.336852, 13.0379, 
    12.56552,
  39.55753, 45.69468, 57.62575, 64.87571, 66.90756, 58.24409, 46.98421, 
    38.7984, 34.37933, 18.54759, 14.1199, 6.09305, 5.813642, 10.29587, 
    17.05504,
  13.30149, 32.53336, 8.355282, 7.407232, 4.22814, 1.048014, 0.7153053, 
    0.5866193, 1.625545, -1.428348, -1.940767, -0.9561903, -1.127535, 
    -0.09182524, -1.584681,
  68.3721, 56.88147, 40.11684, 26.03813, 4.508847, 0.5273022, 0.9635403, 
    0.3278145, -0.0009985565, 0.6875437, -2.445827, 2.52393, 6.510187, 
    -1.549051, -2.793425,
  81.39851, 65.60841, 47.99545, 39.95062, 14.0932, 0.810169, 0.7681339, 
    0.7338738, 0.5268404, 0.6401086, 0.1434827, 2.424726, 7.236571, 10.65053, 
    3.623119,
  88.70378, 73.79662, 60.76027, 51.87826, 39.78304, 19.37771, 1.885115, 
    0.5253685, 1.039932, -0.08564169, 0.03022117, 0.8721144, 4.214062, 
    8.791627, 7.751519,
  101.6248, 84.05923, 72.09203, 58.90822, 42.36943, 30.58704, 29.08043, 
    2.308074, 0.9087524, 0.1503799, -0.453934, 0.01041596, 2.467347, 
    4.409618, 10.49641,
  124.374, 100.4672, 82.80069, 65.71591, 50.5032, 35.18113, 39.07077, 
    32.55652, 4.37772, 3.244015, 1.955873, -0.1146376, 0.9613274, 2.619037, 
    8.54131,
  145.0918, 121.5093, 95.17712, 72.43375, 54.97179, 43.27481, 46.91421, 
    47.55139, 21.87001, 12.02665, 0.9822231, 0.4269893, 0.7771398, 1.805971, 
    5.175327,
  84.00933, 95.23468, 92.83062, 82.95136, 67.74385, 53.99934, 52.55643, 
    55.76779, 48.22968, 20.26272, 1.448886, 0.6188775, 0.9310435, 1.857559, 
    5.942267,
  29.90461, 28.22689, 39.70499, 47.87196, 56.61988, 56.90285, 52.57628, 
    50.88248, 49.68959, 25.42119, 0.7054198, 0.6385462, 0.4554259, 2.111306, 
    9.812976,
  47.57483, 30.0147, 18.88925, 16.17144, 22.56445, 34.83792, 45.58129, 
    45.74036, 33.89213, 10.32452, 9.544725, 1.571931, 0.5819535, 1.788452, 
    11.1174,
  13.57814, 34.1977, 12.2607, 9.249291, 0.5059137, 0.7741088, 3.914135, 
    1.709165, 0.8641163, -2.033188, -1.920604, -1.175854, -2.425058, 
    -1.072011, -2.287942,
  74.78226, 60.23242, 41.62208, 24.98189, 1.29598, 0.8391411, 1.800985, 
    5.049444, 0.5213516, 0.4465938, -1.461738, 2.136908, 6.219481, -2.815194, 
    -3.692159,
  104.0417, 75.02303, 54.88061, 47.97498, 9.977523, 0.9378572, 1.874602, 
    0.6005602, 0.1346452, 0.2656295, 0.5669618, 3.213577, 9.15824, 6.46928, 
    1.046759,
  111.0852, 91.2922, 68.40704, 57.97689, 34.92154, 19.50797, 1.576279, 
    0.3586957, 0.9098591, -0.1441196, 0.6145869, 1.436572, 6.872272, 
    9.558455, 3.188888,
  112.609, 96.64046, 80.47746, 64.25097, 49.81643, 27.98478, 25.65077, 
    2.555064, 1.333963, 0.8687795, 1.896384, 0.2914441, 2.005431, 4.037496, 
    5.690548,
  127.1416, 105.1932, 87.03973, 69.5534, 54.22186, 31.27092, 33.49612, 
    20.94199, 5.129068, 1.758508, 1.192667, 0.2278414, 1.043189, 2.727348, 
    5.636965,
  143.252, 115.2759, 92.98357, 75.30956, 59.79359, 40.08524, 36.57541, 
    33.77793, 23.47128, 9.547459, 1.881151, 1.342453, 0.9182288, 1.058129, 
    4.482892,
  129.3354, 114.8389, 97.59138, 82.43187, 69.3362, 52.93929, 42.8776, 
    44.81554, 40.03536, 20.41593, 3.822012, 2.024852, 1.172462, 0.8066443, 
    5.054892,
  83.22093, 87.92197, 84.60986, 74.09715, 66.51075, 57.17056, 45.71261, 
    42.73257, 43.8128, 19.65173, 5.719695, 2.500978, 1.216195, 0.8742379, 
    8.876205,
  49.56099, 50.45634, 54.73209, 51.43567, 46.83803, 39.51837, 35.63923, 
    30.77153, 20.21692, 11.56435, 13.89837, 6.384721, 2.708577, 1.359933, 
    2.586909,
  23.41496, 49.97394, 21.3794, 17.12297, 9.025062, 4.073584, 5.569523, 
    3.969945, 0.1256429, 0.1748729, 0.1838249, -1.81349, -2.532548, 
    -1.070713, -1.295746,
  102.8972, 113.078, 101.1623, 63.43551, 4.357746, 2.141901, 5.054039, 
    5.89582, 1.016136, 0.123897, -0.3247503, 0.1553202, 0.9931154, -2.406762, 
    -2.305177,
  131.1096, 107.578, 105.7801, 91.31606, 32.81245, 0.49412, 1.669903, 
    4.069776, 0.966688, 0.4910338, 0.8994322, 3.041832, 4.777748, 2.005229, 
    -0.1447813,
  124.8587, 100.9399, 92.42648, 84.71326, 68.12788, 25.80164, 1.089392, 
    0.9511096, 0.551167, 0.2553824, 0.4369473, 4.464934, 4.321387, 3.827909, 
    0.8551162,
  120.2555, 98.7739, 83.09498, 68.2732, 53.19942, 38.30709, 23.57843, 
    0.7229719, -0.1056403, 1.294129, 0.910893, 5.231286, 3.469577, 1.549408, 
    1.553757,
  117.8531, 102.2303, 83.61473, 65.45231, 50.02188, 37.28321, 31.27781, 
    13.15704, 4.682369, 2.492971, 1.844992, 5.442476, 2.79801, 0.3859285, 
    1.249109,
  122.7208, 106.3293, 88.25124, 71.63872, 59.36905, 49.06512, 45.49749, 
    34.44044, 10.49614, 7.618894, 4.471473, 3.554519, 2.136803, 0.257809, 
    0.5811884,
  126.7441, 107.3773, 92.54943, 79.67731, 70.74802, 61.4152, 54.72653, 
    48.96899, 36.64364, 10.6842, 5.784152, 3.475363, 1.692901, 0.2138115, 
    1.19219,
  120.0001, 106.3708, 97.67731, 84.4561, 74.64599, 67.32226, 57.91807, 
    50.4833, 42.52057, 8.942161, 3.080378, 1.727621, 2.347973, 0.7866868, 
    1.549434,
  105.3979, 91.47171, 85.90102, 78.07801, 68.15745, 59.60543, 53.51885, 
    43.82676, 19.27892, 4.433223, 15.33205, 12.64189, 6.926015, 3.822307, 
    1.624696,
  22.22833, 41.37538, 26.72543, 18.32915, 7.438858, 1.596839, 5.425286, 
    2.449892, 1.986639, 0.7831967, 0.08850629, 0.001944832, -2.485955, 
    -1.065739, -1.748997,
  91.24485, 115.6091, 113.8874, 65.07887, 4.520698, 0.2312146, 5.564359, 
    4.209386, 3.166172, 2.751459, -0.1489739, 0.9640814, 2.42536, -1.007937, 
    -1.325,
  123.2562, 130.4299, 142.3843, 126.6546, 48.81153, -1.261877, 1.284333, 
    5.18229, 5.850114, 1.7462, 1.701533, 3.880837, 3.872205, 4.79714, 1.124696,
  124.9263, 130.1762, 135.0383, 130.4988, 115.7138, 46.80382, 1.172284, 
    1.626661, 0.8985941, 1.27995, 2.013076, 5.829338, 3.696787, 3.810457, 
    3.563014,
  127.5713, 129.1324, 128.0264, 119.7102, 104.8124, 86.13882, 40.59246, 
    1.370446, 0.6574772, 0.8781065, 2.284708, 4.543116, 2.786208, 0.4796868, 
    3.941795,
  130.1723, 129.5411, 123.8853, 111.4149, 97.59155, 80.6694, 63.58323, 
    25.23462, 6.342264, 3.1422, 1.922023, 4.164571, 3.01382, 0.03829878, 
    3.104929,
  136.105, 130.1023, 117.1698, 101.8401, 87.08183, 71.64167, 60.77864, 
    44.38995, 20.78153, 8.88689, 5.473445, 4.665816, 3.763793, 0.2467589, 
    1.909569,
  134.9875, 121.0809, 106.4883, 91.64308, 79.61833, 65.30515, 56.09495, 
    49.81306, 36.52143, 5.017908, 1.399805, 3.910501, 5.261173, 2.439451, 
    0.2336047,
  118.4609, 109.0607, 99.55521, 82.19293, 69.74351, 62.12638, 55.14629, 
    48.93284, 42.53249, 8.116418, 3.57538, 7.980077, 7.450477, 4.076424, 
    0.8442473,
  96.87086, 82.99832, 76.27638, 68.51903, 61.49507, 56.25101, 53.88441, 
    48.39561, 22.9142, 6.003797, 12.9489, 9.511526, 5.841746, 3.440416, 
    1.272064,
  22.6576, 32.4407, 18.17668, 11.54107, 3.767122, 0.6167119, 2.206626, 
    1.242267, 1.02083, -0.7703428, -1.128839, 0.30199, 0.2912996, 1.08073, 
    -0.7883871,
  104.5952, 102.4739, 90.40776, 36.42833, 2.40574, -0.2851488, 1.943156, 
    1.327826, 1.461751, 1.114768, -1.799542, 0.1077398, 4.438672, -0.2801046, 
    -1.316779,
  134.59, 124.3738, 125.5938, 102.6243, 39.6147, -1.008629, 0.4807245, 
    0.8904589, 2.473561, 2.526087, 2.62651, 2.219491, 3.614229, 5.362515, 
    0.9192011,
  127.8646, 118.3296, 114.8677, 114.6179, 105.9822, 42.28569, 1.23608, 
    1.014671, 0.5810108, 1.670663, 3.58618, 5.066324, 2.401541, 6.277529, 
    2.598217,
  116.82, 110.0764, 105.7363, 104.7175, 101.714, 89.84661, 47.13345, 
    1.814595, 1.092597, 0.9263912, 3.462831, 5.695686, 4.510716, 6.316182, 
    4.13028,
  109.3323, 106.2468, 100.7064, 98.01514, 95.51157, 88.2784, 73.84159, 
    28.1215, 4.637388, 3.252171, 2.072342, 5.487834, 6.244354, 1.758876, 
    4.931785,
  107.6027, 105.5856, 98.34628, 92.20093, 90.53793, 83.53003, 75.43031, 
    58.51278, 32.12598, 7.967865, 4.807187, 4.652191, 7.83581, 2.331764, 
    4.884169,
  102.7907, 98.10677, 93.18297, 87.43872, 86.05378, 81.12525, 72.84167, 
    67.84283, 53.13207, 6.824866, 3.561195, 6.098897, 6.900964, 5.395291, 
    3.982335,
  87.96717, 88.31148, 88.83035, 78.97267, 72.97, 72.61009, 68.49818, 61.1498, 
    53.6131, 16.7996, 0.8701842, -0.4665387, 3.903913, 2.39498, 2.630861,
  65.93203, 63.70838, 64.57483, 61.38929, 58.09587, 56.21888, 56.8648, 
    54.0829, 34.17706, 6.281018, 9.603544, 0.8643194, 0.07140119, 2.834181, 
    1.59824,
  17.08274, 22.79878, 12.19366, 6.518814, 0.9467631, 0.6370949, 2.524407, 
    2.412424, 3.345431, 1.178244, 0.5990047, 1.947864, -3.061199, -0.3629045, 
    -2.075095,
  89.72498, 78.88132, 70.80174, 19.49694, 0.8558829, 0.2982442, 0.5296374, 
    4.013184, 5.226988, 5.396495, 2.585808, 5.731801, 4.715858, -1.312606, 
    -1.986089,
  125.9799, 109.1019, 105.8027, 77.85902, 28.76685, 0.3009539, 0.7404091, 
    1.241367, 3.300524, 3.742934, 6.396356, 8.760115, 9.395368, 7.533149, 
    2.697002,
  126.5396, 111.0333, 101.0616, 95.2252, 86.14955, 32.39393, 1.476258, 
    1.1478, 1.847766, 3.035673, 4.693535, 9.132061, 10.54852, 10.21661, 
    4.947008,
  123.994, 110.3615, 99.37972, 90.56306, 84.56766, 75.50903, 39.64746, 
    1.908824, -0.1341741, 1.216959, 3.030031, 4.887264, 9.314935, 9.321968, 
    8.712398,
  118.4656, 110.6659, 97.24171, 86.96208, 80.12447, 74.22636, 66.38262, 
    29.21091, 4.293637, 1.129684, 0.6290677, 2.606295, 7.735639, 8.159175, 
    10.53386,
  114.1842, 108.3779, 94.47625, 83.08455, 76.17387, 68.49342, 65.19955, 
    53.25021, 27.70503, 4.474119, 0.8748928, 1.706829, 6.735674, 7.688566, 
    9.97698,
  108.1836, 99.39413, 89.15707, 79.99306, 73.23821, 64.03442, 57.10177, 
    52.6415, 38.28222, 7.933767, 0.7634932, 1.308966, 3.388895, 4.429898, 
    9.216691,
  87.18431, 86.3454, 84.96982, 73.35369, 64.98226, 59.65019, 52.29439, 
    44.0552, 39.48341, 15.87989, 2.627708, 1.461246, 0.444689, -0.5053429, 
    6.303177,
  47.43485, 47.05842, 48.2165, 46.88092, 43.49154, 37.90566, 35.46536, 
    32.77933, 20.92215, 7.014334, 13.57057, 4.201021, -0.2979303, -0.3725488, 
    3.212216,
  10.53724, 16.54176, 7.117758, 2.504647, 1.682591, 0.4128057, 0.2766299, 
    0.09710203, 0.6932734, -0.9842138, -0.5500378, 2.870814, 1.543371, 
    0.6008071, -0.3279994,
  74.27631, 63.69739, 51.66106, 10.81565, 0.7135787, -0.0780296, 0.7539436, 
    0.5714356, 1.062332, 0.9171147, 0.0526816, 5.926825, 6.276806, 0.4043359, 
    -0.1970292,
  102.1033, 82.89684, 68.58689, 42.45002, 15.7169, -0.04038233, 0.9750904, 
    1.097207, 0.6391953, 1.610436, 1.511192, 6.331003, 5.515947, 5.363008, 
    1.909152,
  94.2893, 73.99242, 59.22892, 53.97691, 53.13985, 25.88139, -0.5031691, 
    0.4601661, 0.6478425, 2.041674, 0.4924111, 4.852791, 6.516751, 4.714964, 
    4.085649,
  91.00934, 73.39039, 63.3561, 60.73801, 63.66508, 58.23418, 34.45382, 
    -0.2865628, -0.4529567, 0.6246152, 0.4340631, 2.115819, 6.811916, 
    5.050382, 3.940291,
  91.50684, 80.97996, 72.70546, 69.38122, 66.99736, 61.93395, 49.38157, 
    19.98278, 1.467786, 0.8163297, 0.4999828, 1.111216, 6.37607, 5.176373, 
    3.410509,
  102.2583, 93.00263, 81.38353, 73.52991, 67.73954, 55.82565, 44.06916, 
    28.2466, 8.091382, 1.590002, 3.603325, 0.4251748, 8.575987, 7.192189, 
    4.129333,
  117.3091, 98.69096, 84.92051, 74.10898, 63.5275, 47.44484, 32.31718, 
    23.53262, 11.17871, 1.414122, 2.255944, 0.8335972, 5.082013, 8.726713, 
    5.790557,
  116.3438, 98.79052, 86.3037, 64.16962, 46.22614, 35.11141, 26.80191, 
    19.49836, 19.52842, 2.802256, 0.3982889, 1.860684, -0.3052516, 9.17203, 
    7.959656,
  85.03412, 60.63144, 43.46054, 30.9631, 23.43472, 17.54529, 13.05361, 
    11.47727, 5.306835, 1.182497, 6.138447, 4.773204, -0.1487855, 0.1926806, 
    6.418915,
  7.246726, 7.722124, 2.542367, 1.151054, -0.07612758, -0.8464163, 0.5221314, 
    1.700409, 3.198539, 0.3243846, 0.08580402, 0.6634401, -0.1916987, 
    -0.2634647, -0.6662365,
  58.2199, 37.29919, 22.75604, 4.520345, -1.917446, -2.903551, 0.4648795, 
    0.8115535, 2.708542, 2.76171, 0.7949862, 2.166757, 1.796563, -0.5174991, 
    -1.155372,
  79.22413, 50.22612, 38.10333, 37.55997, 9.458339, -4.661607, -0.5554881, 
    0.6033998, 3.045292, 2.915061, 3.225939, 1.227774, 0.9243242, 1.7286, 
    0.5306609,
  77.64022, 52.14898, 45.12033, 57.78852, 63.11992, 21.69567, -4.955317, 
    -0.8598396, 0.1724278, 3.034958, 1.172018, 1.126351, 0.8137801, 1.893374, 
    1.500754,
  76.92761, 59.07192, 56.1985, 64.07368, 69.28941, 57.11776, 18.87615, 
    -0.393273, -0.392643, 0.05242146, 0.9163216, 0.9349968, 0.889462, 
    1.348927, 2.945161,
  80.68804, 72.46483, 65.87189, 63.92653, 64.63512, 53.8386, 32.24916, 
    6.037809, 0.4705498, 1.151992, 2.375057, 2.528286, 0.6164359, 0.7661468, 
    2.62862,
  87.63432, 79.33015, 67.46415, 62.40193, 60.74817, 44.32622, 29.77818, 
    16.20581, 3.666794, 2.050765, 4.515259, 1.164024, 1.153472, 0.6023744, 
    1.416373,
  107.0292, 88.11824, 74.2562, 66.67204, 58.00711, 37.96879, 23.13296, 
    16.79456, 7.003991, 4.458494, 3.97069, 2.632654, 1.545469, 1.077764, 
    1.10984,
  120.0127, 100.9114, 87.51768, 66.10465, 44.65312, 29.81259, 21.70095, 
    12.85546, 20.47687, 7.983472, 5.416316, 4.646871, 3.401493, 3.171158, 
    0.6614599,
  116.0796, 90.63185, 68.54478, 51.21669, 34.01461, 25.30859, 15.53687, 
    18.15434, 10.32999, 2.254669, 7.632349, 6.066761, 6.463171, 3.882585, 
    1.426278,
  11.09611, 10.35876, 4.550984, 3.553478, -0.3129986, -1.001043, -0.3654585, 
    -1.909333, -1.253081, -1.521389, -2.075215, -0.9933099, -1.139876, 
    -0.4398958, -0.5344399,
  61.02659, 48.06143, 38.10545, 7.428717, -3.03936, -3.080598, 0.07463632, 
    -2.917236, -2.01302, -0.3237132, -1.566895, 0.343835, -0.2687302, 
    -0.8874721, -0.7694766,
  102.2306, 80.73547, 72.74444, 59.77872, 11.72549, -6.219584, -0.9898472, 
    -1.439836, -0.8284131, -0.4333771, 0.7292968, -0.4291794, -0.009113139, 
    0.7599922, 0.5420966,
  107.7566, 90.48556, 79.81256, 78.41113, 76.17835, 21.98814, -6.907546, 
    -1.613366, -0.7476686, -1.373742, -1.124215, -0.07554233, -0.02159486, 
    1.448426, 0.8455588,
  100.816, 91.61137, 83.3195, 80.33856, 77.1692, 62.42758, 22.78151, 
    2.472059, 1.319631, -3.535224, -1.603065, -0.6341151, 0.5534724, 1.07504, 
    2.444677,
  97.00207, 90.35598, 83.10506, 77.17623, 70.48801, 61.35701, 46.10346, 
    12.26883, -1.569687, -1.045488, -0.7801447, 0.4420822, 0.5284873, 
    0.7073554, 2.70805,
  117.2422, 102.9123, 87.42103, 76.73817, 69.58231, 60.27348, 53.95155, 
    40.01564, 10.7631, 0.563759, 0.2021647, -0.01071768, 0.4107583, 
    0.2465282, 2.026705,
  134.3343, 114.3648, 98.56543, 85.10333, 75.54594, 65.06734, 53.71107, 
    44.37587, 15.56352, 3.592594, 0.1145135, 0.08604349, 0.8994926, 
    0.6351922, 1.927069,
  125.7478, 115.8997, 107.6107, 85.74478, 72.18227, 64.81384, 54.3349, 
    26.85908, 27.24333, 7.301414, 0.920945, 0.6371266, 0.7114252, 2.835636, 
    1.795042,
  102.4674, 92.4741, 83.31606, 76.30054, 70.70908, 51.52143, 25.69902, 
    25.90574, 13.18707, 3.061278, 10.52678, 3.170315, 0.8643384, 5.493074, 
    1.271303,
  14.58924, 16.78651, 10.6947, 8.427719, 1.065692, 1.286234, 2.688967, 
    0.5406233, -1.103798, -4.557888, -5.559404, -4.7809, -3.58154, 
    -0.3985161, 0.08429023,
  63.89902, 64.33423, 68.15115, 23.23631, -1.381936, 0.4095814, 4.436946, 
    1.387655, -0.4176323, -2.481973, -4.805069, -3.039433, -2.310397, 
    -0.902095, 0.2273798,
  100.4755, 102.544, 105.2819, 89.39794, 22.39526, -3.385552, 6.246519, 
    2.007766, 0.2501453, -1.418857, -1.83044, -2.676917, -1.890622, 
    0.3202477, 3.138744,
  94.44328, 96.11738, 96.97085, 101.8043, 99.63952, 37.9515, -5.252584, 
    1.93853, 2.157538, 0.9811754, -0.5571719, -1.343664, -0.8591319, 
    1.149935, 6.47956,
  88.68691, 87.99039, 90.73826, 96.89995, 99.25885, 91.00958, 47.88388, 
    -3.710571, 5.539172, 0.7220715, 0.985905, -1.424792, -1.023717, 
    0.8506967, 7.915033,
  90.99182, 90.4763, 91.69444, 93.82588, 93.943, 89.95068, 78.79163, 
    39.35892, 2.719269, -1.518754, -2.093357, -1.078406, -0.8990402, 
    1.104421, 7.991939,
  105.8016, 104.9553, 96.90771, 90.13425, 86.89614, 78.24458, 72.35986, 
    58.15146, 31.03196, 4.111075, -0.2803243, -1.075849, -0.4818511, 
    1.675105, 9.507362,
  107.1344, 99.29503, 89.72141, 78.418, 72.18621, 62.51011, 52.66475, 
    48.25158, 28.13189, 3.673615, -1.328251, -1.215957, -0.06426112, 
    4.294222, 8.811193,
  90.27811, 85.33817, 83.36359, 61.23458, 48.87893, 43.47573, 40.93189, 
    28.91154, 27.32003, 5.934484, -0.6122813, -0.8283917, -0.1801715, 
    7.123547, 8.089182,
  76.29438, 59.90445, 50.89516, 42.09608, 36.43325, 25.21506, 18.30215, 
    24.93946, 20.5172, 9.006474, 11.31887, 2.105595, 1.458268, 11.84436, 
    10.06992,
  15.72382, 19.07047, 10.70595, 7.113619, -0.6367933, 1.363595, 3.806137, 
    -0.2206943, -1.613441, -1.564519, -1.055347, -0.4605925, -1.327691, 
    -0.4374749, -1.302706,
  62.23787, 67.84962, 74.99915, 28.27457, -3.28436, 3.188649, 7.877884, 
    0.60919, -0.6572022, -1.339212, 0.8426532, 3.191484, -1.094352, 
    -2.434501, -1.815938,
  125.7949, 124.0461, 126.0558, 106.2739, 18.06061, 4.509028, 12.26436, 
    3.356738, 0.8128174, 1.42373, 4.641937, 1.424961, -1.052207, -0.3982835, 
    2.00405,
  135.1759, 131.3084, 125.604, 121.8303, 114.664, 47.97168, -2.910938, 
    6.12469, 8.305097, 7.596898, 4.87257, 0.9738377, 0.9320605, 2.058074, 
    7.833517,
  138.3601, 134.2627, 126.9165, 121.4669, 116.163, 103.3968, 54.09521, 
    3.516146, 4.112544, 6.704878, 5.296577, 0.3917941, 1.435472, 2.512043, 
    9.978131,
  129.419, 131.443, 128.7714, 119.5501, 110.619, 96.38457, 76.9692, 43.10973, 
    7.056839, 2.640622, 0.4069771, 0.9048219, 2.178325, 3.39434, 8.868921,
  117.5053, 124.1768, 118.0266, 110.1082, 97.46327, 79.39495, 61.92112, 
    39.97672, 19.38669, 6.607297, 1.081368, 0.8099793, 2.017826, 7.226653, 
    11.05634,
  104.5738, 100.1254, 96.15104, 89.78866, 80.24786, 65.37197, 44.86188, 
    30.39183, 17.83506, 2.98122, -0.962851, 4.089853, 3.27943, 11.71073, 
    9.343472,
  91.6655, 87.76267, 86.63747, 67.34834, 58.8918, 52.90306, 36.70835, 
    21.57247, 15.76316, 4.457379, -0.02230215, 4.856136, 6.428777, 15.64835, 
    7.751491,
  68.79224, 56.1526, 48.44509, 41.20295, 38.58993, 29.03275, 16.46228, 
    13.00393, 9.805787, 2.6528, 11.01609, 9.077023, 13.82538, 19.40878, 
    12.06738,
  20.60157, 30.32688, 19.89192, 15.88396, 2.453444, 6.697354, 12.18001, 
    2.74144, 0.6514192, -1.074935, -0.3154721, 0.6796522, -0.1562666, 
    1.455447, -1.414905,
  68.29458, 82.65501, 82.98494, 42.02277, -0.6128617, 14.4743, 22.7748, 
    5.11364, 2.850668, 0.9826097, 0.5877157, 5.08845, 4.513945, -0.6439924, 
    -1.483436,
  123.899, 145.898, 155.5166, 133.6622, 29.59651, 0.4474408, 31.42752, 
    10.40829, 2.882557, 1.965476, 3.908322, 4.813197, 5.317468, 2.042396, 
    2.154827,
  87.04647, 112.8011, 130.3719, 144.513, 150.7506, 67.82391, 1.031154, 
    14.67446, 13.43662, 4.940795, 5.153761, 6.765351, 4.549097, 4.390751, 
    8.450621,
  52.67962, 61.86754, 77.87392, 101.2584, 125.0484, 137.7057, 90.30102, 
    2.356297, 3.353236, 10.72205, 12.78035, 6.095914, 4.626577, 5.371455, 
    10.88862,
  38.24305, 38.59344, 40.7076, 52.74179, 71.71147, 94.86112, 118.6036, 
    94.47249, 16.92625, 7.052399, 6.424479, 5.805183, 5.191628, 9.314658, 
    7.60779,
  41.93066, 37.36334, 26.95583, 26.85499, 32.28986, 45.95699, 62.85778, 
    82.65483, 67.14292, 17.50184, 9.85369, 5.877537, 5.700848, 12.14485, 
    8.841957,
  47.59095, 35.06035, 23.88915, 18.40948, 18.12976, 25.71507, 29.21385, 
    41.80032, 36.72779, 16.42183, 11.18068, 6.265831, 10.91283, 12.15478, 
    4.963975,
  63.56519, 57.4529, 44.70818, 23.2788, 14.65771, 16.59018, 25.2606, 
    26.94181, 23.28276, 19.42702, 12.92336, 10.4985, 13.11523, 11.61774, 
    4.606426,
  65.46201, 56.60966, 41.9995, 26.29555, 15.37045, 6.685363, 7.679442, 
    13.22472, 15.76409, 11.76514, 22.25762, 15.66688, 18.20195, 14.46988, 
    9.143884,
  22.31285, 41.82386, 23.81147, 19.84408, 1.913201, 7.394906, 15.21095, 
    2.941142, 1.371723, -0.745594, -0.5474017, 0.8977721, -0.05770789, 
    0.340385, -0.4151376,
  60.24287, 76.22002, 67.01897, 33.8489, 0.08519208, 17.09135, 24.19915, 
    4.906903, 2.703791, 1.536101, 1.021081, 3.028128, 1.920331, -0.2932227, 
    -0.1344599,
  129.073, 139.5308, 151.3822, 128.5015, 30.57735, -0.766568, 28.06095, 
    9.183539, 4.207488, 2.278802, 4.007248, 2.195721, 1.527375, 1.34636, 
    -0.6190421,
  71.36657, 130.7758, 146.0695, 160.6456, 158.6333, 62.49929, -1.411533, 
    12.44693, 11.30653, 5.460469, 4.152697, 3.486592, 2.78645, 3.450991, 
    3.013888,
  19.32068, 76.99693, 117.6985, 135.3599, 155.0155, 142.1637, 91.00884, 
    -1.471523, 0.3412119, 7.764553, 12.71935, 5.746925, 3.715983, 6.524325, 
    5.59503,
  49.47943, 41.90141, 83.13833, 101.7558, 121.6066, 126.553, 126.9997, 
    90.95529, 19.34705, 7.405837, 7.564253, 9.83874, 5.752183, 5.678336, 
    3.028652,
  86.1485, 58.89543, 58.26816, 74.37655, 93.902, 102.0984, 104.5146, 
    96.96236, 72.1911, 22.33753, 12.01586, 7.443448, 6.58411, 4.833464, 
    2.50026,
  113.4389, 74.77645, 47.49895, 43.21021, 56.47236, 67.45911, 70.78571, 
    75.81577, 64.91847, 16.34413, 12.06474, 10.6332, 7.060524, 1.812683, 
    1.59411,
  134.8289, 116.9446, 89.39108, 52.38294, 33.32264, 28.78196, 35.29733, 
    41.1111, 34.26794, 15.21102, 9.442139, 14.66119, 5.44729, 3.259635, 
    2.266409,
  117.2437, 108.7467, 97.17236, 78.41349, 62.59727, 40.71472, 15.35693, 
    17.45927, 14.42144, 12.34039, 17.30555, 18.46424, 11.18237, 6.489121, 
    8.142972,
  19.89256, 38.32197, 23.92707, 16.20843, 0.1235649, 4.226707, 9.525249, 
    0.9393094, 3.09822, 0.01007217, -0.5800887, 0.8250026, 0.1331111, 
    -0.1268196, -0.2605721,
  55.4377, 66.36122, 55.91887, 24.03334, -1.471316, 11.40703, 10.69614, 
    1.457098, 0.8986131, 1.900687, 0.5258155, 1.554246, 2.064913, 0.0321008, 
    -0.2022071,
  139.9185, 118.7841, 127.4246, 90.10793, 23.28973, -3.109636, 8.88983, 
    2.146485, 0.6237631, 0.620444, 3.061792, 0.2374202, -0.08518, 1.155644, 
    0.09802637,
  138.7178, 138.8376, 148.6567, 161.5416, 138.7313, 47.10777, -3.120254, 
    2.008982, 1.993137, 0.709151, 0.6035123, 0.3502293, -0.0004253625, 
    0.8147698, 2.333973,
  120.8029, 126.7297, 137.3749, 149.0183, 153.7443, 132.3467, 81.57898, 
    -2.065093, -2.273005, 1.589857, 4.034198, 2.718947, 0.9015378, 1.882506, 
    3.78464,
  105.729, 116.7153, 124.7765, 131.653, 140.1079, 134.7871, 129.0983, 
    83.74647, 20.76351, 8.892305, 9.277593, 6.082729, 1.574183, 1.358453, 
    0.7865368,
  99.74789, 108.0068, 111.3518, 115.5965, 120.994, 119.4792, 116.5507, 
    104.6818, 79.20172, 29.50753, 12.8985, 3.873017, 1.844878, 1.403048, 
    0.2956401,
  106.0831, 95.43082, 96.10548, 99.86343, 104.737, 104.9484, 99.24001, 
    99.0429, 79.9278, 18.85373, 6.013254, 2.924318, 1.924449, 0.2722466, 
    -0.5743543,
  109.3908, 92.57372, 89.33399, 81.73631, 83.99887, 86.65121, 87.77892, 
    84.01328, 62.5155, 9.605803, 2.018128, 3.640275, 1.184665, 0.02972057, 
    -0.6723465,
  118.5799, 93.41724, 74.78822, 61.09295, 59.93667, 55.70576, 47.02143, 
    44.05295, 27.64898, 4.355146, 20.8393, 11.43981, 4.431174, 1.808198, 
    2.046512,
  20.99783, 34.96086, 19.54382, 11.34887, 1.211518, 1.701319, 9.63632, 
    3.670358, 6.784611, 1.711643, -0.2112006, 1.409892, 0.05721566, 
    -0.1645085, -0.5037336,
  63.27058, 69.04553, 59.93394, 17.27278, -0.539054, 3.159139, 4.322719, 
    2.373714, 2.456975, 5.384324, 0.2043052, 2.294691, 4.096256, 0.002093374, 
    -0.3678253,
  146.8741, 118.4246, 114.6226, 59.11048, 20.66039, -2.599115, 1.537438, 
    1.069307, 0.9125943, 1.108115, 3.738207, 1.476287, 0.9181105, 2.023468, 
    0.1710481,
  166.4726, 159.787, 154.1886, 140.2215, 109.0107, 36.95096, -1.684811, 
    -0.510194, 0.4456949, 0.3688377, 0.2544344, 0.4800326, 0.341624, 
    0.837231, 0.8030855,
  160.7214, 153.2652, 148.9286, 144.3466, 132.2302, 111.0273, 72.36047, 
    -0.6806368, -1.104578, 0.5506509, 1.100345, 1.599476, 0.3967465, 
    0.9456145, 1.53078,
  161.1817, 148.8614, 141.5025, 134.8767, 129.4132, 121.2184, 105.1389, 
    60.90562, 17.07412, 10.03014, 3.388005, 2.480997, 0.5734553, 0.3286156, 
    0.5311942,
  160.6834, 156.5592, 139.9457, 127.0052, 121.4512, 113.5024, 103.786, 
    86.42385, 63.31908, 23.57274, 6.351859, 0.8659413, 0.6260529, 0.2638762, 
    0.02923573,
  157.9491, 144.1775, 132.8425, 122.1266, 113.5636, 106.471, 93.27217, 
    86.82108, 67.68479, 13.71044, 0.9636956, 0.1246292, 0.4871922, 
    -0.07826704, -0.1344487,
  141.8503, 136.0471, 134.2692, 114.6693, 101.83, 94.73858, 85.71942, 
    78.26839, 59.29343, 3.759375, -0.3686389, 0.5323474, 0.2991954, 
    -0.151412, 0.08454645,
  112.7322, 107.3674, 102.1606, 91.31337, 87.60993, 76.61287, 60.09325, 
    51.21246, 11.30759, 1.20857, 11.84962, 2.734981, 0.7090364, 0.474739, 
    0.6024845,
  22.23557, 31.86886, 16.60464, 12.37874, 4.077756, 1.152878, 5.734324, 
    2.26664, 7.314206, 1.098366, -0.9157621, -0.01312651, -0.2673116, 
    -0.001310782, -0.521365,
  78.35322, 64.58408, 60.62361, 20.76217, 4.31933, 0.05428689, 2.273893, 
    1.229744, 1.269176, 5.978805, -0.6641939, 0.9222888, 4.413029, 
    -0.2352125, -0.5051381,
  146.9324, 109.49, 106.9174, 43.38867, 30.00633, -1.562005, 0.3198791, 
    0.9749001, 0.9638099, 1.392915, 2.60321, 0.7150165, 1.256325, 2.322798, 
    0.3247022,
  182.0668, 167.938, 152.2977, 116.7198, 89.17094, 39.09883, -0.196683, 
    0.2328766, 1.116352, 0.2832803, -0.001485779, -0.3052641, -0.2137082, 
    0.2538901, 0.3330145,
  181.2013, 164.3027, 145.9015, 134.4036, 114.7405, 90.38945, 61.93287, 
    1.18782, -0.2507572, -0.30248, -0.2397035, 0.07863513, -0.2816444, 
    0.028429, 1.020561,
  187.3037, 163.5353, 141.3132, 125.2299, 115.9747, 101.7845, 80.3368, 
    46.59472, 16.14249, 9.915348, 1.265805, 0.8271359, -0.2130556, 
    -0.1396713, 0.5810201,
  192.9508, 173.0439, 142.7937, 122.384, 109.3453, 101.1221, 90.67538, 
    76.4241, 53.09095, 19.24258, 3.534718, 0.314263, -0.1946273, -0.2789749, 
    -0.5259003,
  191.6284, 163.6473, 138.6517, 119.4478, 105.75, 97.9306, 88.52231, 
    84.07422, 50.8004, 8.81254, 1.037233, 0.5060514, 0.06616116, -0.6467129, 
    -0.6022408,
  177.6573, 157.3645, 141.5645, 113.9118, 97.00634, 85.96732, 79.54613, 
    71.48424, 45.66077, 2.469692, 0.9841859, 1.492721, 0.9228254, -0.447767, 
    0.2154918,
  152.5922, 134.033, 115.3111, 95.84639, 85.08085, 71.62435, 56.33461, 
    46.95739, 5.874403, 3.73544, 8.057158, 1.174014, 0.7223753, 0.7775673, 
    -0.1122638,
  15.87134, 18.76693, 8.131706, 8.242081, 3.347142, 0.6719509, 2.564712, 
    1.420087, 7.469917, 2.131357, 0.1379902, 1.462156, 0.6622924, 0.407781, 
    0.01095961,
  61.58652, 40.36055, 36.06594, 13.7854, 3.197062, -1.009471, 0.242777, 
    0.3142565, 0.8181628, 6.600163, 0.4639015, 2.737119, 5.284531, 0.388549, 
    -0.1621939,
  114.4022, 71.91082, 66.90151, 27.19086, 22.72086, -0.8458874, -0.7628998, 
    0.245169, 1.534502, 2.81328, 2.833883, 2.183099, 3.269195, 3.670285, 
    0.5326001,
  144.7977, 125.3666, 107.7047, 70.9413, 54.74907, 26.07757, 0.8888339, 
    -1.084572, 0.9244533, 1.857922, 1.553599, 1.339986, 1.626328, 1.804221, 
    0.5858628,
  150.7523, 132.5568, 112.3114, 97.93046, 79.83254, 58.59063, 36.56096, 
    0.7614123, -1.642516, -0.1647211, 1.161354, 1.977741, 1.037422, 
    0.7029938, 1.329924,
  161.7714, 139.1353, 114.0029, 98.62347, 91.32633, 82.46001, 67.61968, 
    40.37791, 13.98211, 9.887424, 0.6553971, 2.058656, 2.246067, 0.9230723, 
    2.053214,
  177.8549, 153.09, 121.7386, 101.3309, 91.36643, 87.53484, 85.46003, 
    74.94579, 50.33876, 19.64761, 5.294463, 3.060111, 2.522828, 1.587924, 
    0.8527647,
  189.5227, 155.9552, 124.6182, 103.8313, 91.05861, 85.92097, 80.11664, 
    79.29354, 39.04864, 10.95281, 4.532603, 2.362721, 2.75802, 1.687791, 
    2.593197,
  184.7265, 157.3777, 137.3161, 106.1584, 88.28087, 79.49378, 74.92304, 
    66.16909, 35.10575, 3.628879, 3.096787, 4.341189, 2.096451, 1.533079, 
    4.770424,
  164.3042, 139.0993, 116.9511, 94.88786, 80.84007, 68.55215, 52.82988, 
    42.53783, 4.156323, 2.425681, 8.466454, 2.578623, 1.914096, 0.9313082, 
    4.20955,
  6.918462, 11.30589, 4.783022, 8.69015, 4.768448, 1.038756, 2.790328, 
    2.589309, 5.931563, 1.362358, 0.01560024, 0.5925379, 0.2112717, 
    0.7091407, -0.5106096,
  33.27906, 24.22874, 23.6187, 12.52046, 3.160642, -0.2595853, 1.336006, 
    1.877489, 2.086587, 5.29507, 1.073556, 2.557749, 4.674639, 0.211956, 
    -0.3366299,
  66.98876, 44.38277, 48.4646, 23.19744, 20.2512, -0.08458579, 0.0195942, 
    1.80874, 2.512485, 3.583096, 3.728193, 2.05739, 2.469242, 2.492198, 
    0.5137846,
  81.02215, 71.12636, 64.85213, 49.43845, 42.07266, 23.68692, 0.9287721, 
    -0.03818915, 1.402941, 1.427831, 0.9624852, 0.3414597, 0.6625904, 
    1.626881, 1.63386,
  80.31509, 66.34386, 56.23251, 55.61992, 53.63073, 43.01221, 36.50462, 
    1.089334, -0.3449547, 0.0481331, 0.1600429, -0.02580942, 0.07104061, 
    2.055907, 1.797926,
  84.46951, 68.27753, 58.98163, 57.04462, 58.12016, 58.02185, 46.09645, 
    27.17335, 11.92252, 6.886523, 1.102544, 0.9043821, 2.054952, 1.63114, 
    1.199638,
  97.10349, 83.99274, 72.23737, 66.48504, 65.54422, 64.80518, 63.54066, 
    56.14337, 36.10329, 16.47599, 7.805425, 2.817779, 3.149524, 1.727736, 
    0.4304023,
  111.714, 94.03904, 83.57626, 77.36305, 72.64751, 72.5695, 69.74502, 
    70.58344, 31.25874, 12.88601, 7.05876, 6.251244, 3.722001, 2.951324, 
    3.671376,
  118.7129, 105.0685, 101.132, 86.33358, 77.4146, 74.11215, 73.00768, 
    63.03328, 36.00825, 12.99251, 9.210077, 8.12495, 4.353728, 1.092728, 
    3.167009,
  116.1531, 102.1497, 95.80022, 82.74215, 78.20937, 64.57455, 51.88446, 
    43.58713, 16.92286, 8.909548, 14.94246, 4.641979, 3.18861, 1.091094, 
    5.082088,
  6.866405, 12.11227, 7.440466, 7.557224, 4.192243, 1.041064, 2.527581, 
    3.49837, 9.989483, 4.059295, 0.7319483, 1.412251, 0.00743485, 0.5891928, 
    -0.5462293,
  33.39428, 25.84284, 23.35131, 12.64, 3.152363, 0.03681581, 1.838713, 
    2.42672, 2.962511, 9.301719, 1.132095, 4.568504, 8.271872, 0.6829286, 
    -0.6231328,
  74.53683, 49.05962, 54.76242, 26.08775, 20.35403, -0.4757505, 0.609773, 
    2.37357, 3.543193, 4.735531, 5.736291, 3.236716, 5.324316, 6.268993, 
    1.075771,
  86.70895, 83.66671, 84.12639, 61.58627, 51.69527, 24.59933, 0.464794, 
    -0.2430109, 1.850308, 1.817282, 0.9601849, 0.8730577, 2.616858, 4.156607, 
    2.992189,
  80.39858, 77.28609, 79.4409, 82.1995, 72.66193, 55.49557, 42.76293, 
    1.217695, -0.2517184, 0.1942339, 0.9318044, 1.030453, 1.55189, 3.018736, 
    2.421076,
  74.72267, 70.36242, 69.028, 70.83138, 71.21909, 67.92098, 48.08621, 
    24.21361, 12.97038, 12.0619, 1.496627, 2.336644, 3.127031, 1.366861, 
    1.327822,
  70.14317, 70.26904, 65.92292, 64.57822, 63.61613, 65.46491, 59.46345, 
    44.84966, 30.92755, 14.32806, 8.216029, 4.576352, 3.724916, 0.2453773, 
    0.4877162,
  68.01521, 69.17648, 65.38541, 63.42719, 59.53327, 61.70404, 57.48721, 
    58.38144, 26.24035, 11.09135, 7.315159, 5.867043, 3.843086, 1.832813, 
    2.370294,
  72.47325, 72.38429, 73.85424, 65.43279, 59.07335, 57.65696, 55.32922, 
    48.44593, 25.63393, 9.270832, 6.72471, 6.658771, 4.758523, 1.899341, 
    4.302763,
  76.81453, 69.99756, 66.92525, 59.07172, 55.8156, 45.4808, 41.87849, 
    41.00342, 18.69978, 11.42786, 13.04423, 5.782802, 1.541925, 0.8644131, 
    3.986528,
  6.388035, 8.90411, 4.962897, 4.139628, 1.943253, 1.350938, 3.135601, 
    4.140835, 7.17861, 2.240658, 0.709874, 2.173063, 0.8170034, 0.09931247, 
    -0.5647999,
  25.75513, 19.19607, 14.94981, 6.481943, 1.980212, 0.2751198, 2.613648, 
    4.42171, 3.64321, 5.947108, 1.086976, 4.270164, 7.530069, -0.02620844, 
    -1.133828,
  68.41074, 40.94712, 39.49126, 17.41117, 16.62776, -0.0742311, 1.041465, 
    4.233152, 4.297518, 3.995972, 5.500649, 4.027871, 5.123505, 8.494543, 
    1.807762,
  84.04762, 68.12806, 60.70402, 45.54222, 46.05194, 24.82908, -0.3182441, 
    0.3090553, 0.4179733, 0.8659896, 1.156277, 1.057529, 2.291552, 3.354586, 
    5.267365,
  79.82899, 62.36317, 55.444, 60.55046, 70.627, 62.06534, 49.56425, 
    0.7589381, -0.6031016, -0.1922876, 0.5572335, 0.8089683, 1.144537, 
    2.498991, 3.236842,
  82.05742, 60.95105, 50.19255, 53.02166, 69.75645, 74.07005, 55.64823, 
    29.89597, 15.72624, 17.33043, 3.082911, 2.042516, 0.9659197, 0.7868986, 
    1.45302,
  90.76971, 68.03381, 51.27436, 51.53168, 60.48287, 71.09749, 68.1192, 
    48.22852, 29.40718, 16.00048, 9.578324, 3.637832, 1.315687, 0.1304238, 
    0.3802457,
  94.19666, 70.73887, 55.31953, 51.98014, 54.12405, 60.81882, 60.51667, 
    61.67469, 25.23521, 10.39421, 6.610447, 3.282655, 1.285171, 0.1427898, 
    0.3759757,
  88.18517, 76.79643, 67.95038, 55.78798, 50.40701, 50.52664, 51.24622, 
    46.14695, 18.48466, 6.013133, 4.631451, 3.451361, 1.142103, 0.4416799, 
    2.017945,
  68.82475, 65.08752, 58.61722, 49.71735, 44.45569, 35.97164, 37.32862, 
    37.18366, 11.6181, 11.69871, 12.59933, 3.654423, 1.814511, 1.480222, 
    2.239727,
  4.388189, 5.709753, 3.275817, 4.545206, 4.005537, 1.692399, 1.695522, 
    1.977994, 7.584723, 3.321341, 1.320626, 2.62773, 0.5780239, -0.2434583, 
    -0.6588875,
  19.54116, 15.21366, 9.333258, 4.051891, 1.564445, 0.3647751, 2.50382, 
    2.529792, 5.16563, 10.08803, 3.865289, 5.933836, 8.623833, 0.0781113, 
    -0.882863,
  63.86889, 43.11731, 35.07822, 13.29846, 9.447755, 0.3447632, 0.4391579, 
    2.552718, 5.004588, 8.020439, 8.178792, 4.06084, 4.826558, 9.230638, 
    2.609009,
  91.56107, 79.43638, 66.25795, 42.07096, 34.76308, 17.58269, 1.161399, 
    0.8782402, 2.99053, 3.620505, 2.558389, 0.2890934, 1.1295, 3.316309, 
    6.546983,
  96.24668, 84.19604, 75.2868, 65.51451, 57.80898, 46.41997, 43.7305, 
    2.139687, -0.2280078, 0.4420246, 0.60956, 0.1849463, 0.5101025, 2.600175, 
    4.471726,
  101.8371, 87.89344, 80.18446, 69.64695, 62.5693, 57.87349, 47.34915, 
    27.69484, 16.69691, 19.65109, 4.726748, 1.25349, 0.4518113, 0.5157449, 
    0.7601919,
  108.7448, 93.66865, 79.57963, 67.82495, 62.03089, 62.24409, 60.34958, 
    42.26848, 30.03499, 15.57199, 9.226762, 2.728594, 0.8791099, -0.1059055, 
    -0.03699078,
  105.755, 82.97324, 69.71866, 61.26823, 58.04163, 62.13078, 63.22522, 
    65.12022, 27.13642, 7.506483, 3.423671, 2.166056, 0.8241341, -0.2111501, 
    -0.3894435,
  91.98398, 70.78197, 59.30465, 50.15725, 49.13982, 53.82518, 58.84792, 
    48.13334, 10.7264, 2.146027, 0.9437912, 1.831651, 0.7519641, 0.1378007, 
    0.7936348,
  70.52986, 51.20567, 36.87776, 31.63184, 34.71836, 36.86619, 39.20161, 
    29.62205, 4.867118, 6.938465, 13.6, 3.359471, 1.96418, 1.880352, 1.297778,
  4.044114, 6.816444, 2.591328, 3.341135, 2.977991, 1.061741, 1.683389, 
    2.072923, 5.544252, 1.414718, 0.1695678, 2.416718, 1.508582, 0.03083469, 
    -0.2535711,
  20.78418, 17.72585, 9.642958, 3.396045, 1.480908, 0.2798037, 0.3274716, 
    1.322605, 2.812196, 4.997379, 1.637199, 5.17753, 7.512562, 0.1208669, 
    -0.326828,
  80.41451, 58.03146, 42.65614, 14.10658, 8.784615, -0.1013111, 0.2998252, 
    0.1962056, 1.633297, 3.477793, 4.650483, 4.02741, 4.53861, 5.023382, 
    1.809947,
  129.2487, 109.3778, 91.0023, 57.75541, 37.91636, 15.55416, 0.5197056, 
    0.3381503, 2.200316, 1.086949, 0.6325354, 0.5314354, 0.844766, 3.603487, 
    4.797509,
  142.2511, 117.7249, 100.3143, 85.74317, 71.43305, 41.65548, 43.24298, 
    1.176609, -1.221175, 0.3158872, 0.4032465, 0.4754507, 0.4596883, 
    2.188372, 4.132111,
  154.6587, 127.9421, 108.6336, 89.15532, 73.53083, 50.48246, 48.82312, 
    34.62307, 17.03575, 17.83146, 7.612364, 2.495625, 0.617137, 0.4563054, 
    0.8530292,
  168.7473, 146.8099, 117.9049, 91.71568, 74.40262, 52.22624, 48.55627, 
    38.5601, 29.69434, 16.53453, 10.13646, 2.450294, 1.074703, 0.204908, 
    0.3505172,
  174.245, 144.4797, 116.1113, 92.47206, 73.87418, 58.18258, 43.51696, 
    48.29106, 25.47779, 5.600669, 2.412003, 1.579889, 0.6247523, -0.1213053, 
    -0.2287036,
  161.0893, 135.01, 117.8717, 89.03242, 69.99001, 52.90858, 41.89174, 
    30.9488, 3.421309, -0.4220638, 1.124134, 2.172003, 0.5699536, 0.04365128, 
    0.1990537,
  128.4202, 106.845, 87.41223, 65.43203, 52.7134, 31.5861, 18.62258, 
    12.98102, 0.8293166, 4.063568, 14.12666, 5.07519, 1.920794, 2.749535, 
    0.9467462,
  14.55886, 16.60509, 10.59774, 8.299086, 3.463044, 1.173187, 3.684113, 
    2.849663, 4.408836, 0.8552094, 0.439912, 1.152976, 0.3831888, 0.1364698, 
    -0.1279447,
  26.49326, 28.49026, 22.98479, 13.21264, 2.421565, -0.03705001, 1.410222, 
    1.184445, 2.380005, 3.463023, 0.9818017, 3.768773, 4.403581, 0.08725008, 
    -0.1738581,
  78.56872, 81.49058, 61.45955, 31.7697, 13.58117, -1.288976, 0.1987442, 
    0.4304881, 1.365633, 2.810546, 3.299643, 2.245838, 2.784974, 3.399297, 
    1.216147,
  135.2973, 143.6265, 144.2414, 105.165, 70.1602, 22.22945, -0.2664168, 
    0.1321648, 0.4227335, 0.7584792, 0.7588061, 0.5889272, 1.575834, 
    2.631922, 3.176378,
  134.873, 144.8641, 152.7446, 153.5213, 136.9306, 87.12828, 55.70242, 
    0.7168612, -1.026034, -0.02191875, 1.047182, 1.299143, 0.5948645, 
    2.10823, 3.098607,
  137.0857, 146.1478, 153.0368, 149.6087, 140.7331, 119.0614, 87.04352, 
    39.554, 13.56976, 14.00337, 10.31241, 3.716467, 0.5048596, 0.1646888, 
    0.1363548,
  141.2507, 158.7949, 156.6927, 146.0507, 135.9337, 117.5361, 96.63229, 
    50.94432, 28.03129, 13.27633, 10.55942, 2.286835, 0.8982582, -0.03143292, 
    -0.247006,
  134.7119, 148.5623, 154.1508, 146.1526, 131.8513, 115.1963, 88.50205, 
    70.79274, 27.83645, 8.05227, 2.678135, 1.586658, 0.5943199, -0.5030316, 
    -0.5328822,
  120.2707, 139.0359, 157.8953, 145.3652, 126.6838, 102.7665, 81.90085, 
    47.70535, 2.819022, 1.151671, 4.035663, 5.124688, 1.126728, -0.3183497, 
    -0.6377057,
  92.88868, 108.1187, 125.096, 117.2876, 105.6353, 72.67341, 49.33298, 
    17.38741, -1.125652, 0.996522, 12.10302, 9.217152, 6.228098, 3.211774, 
    0.1747036,
  9.359711, 11.05099, 14.00344, 10.5895, 3.771117, 1.77404, 5.003469, 
    2.803015, 4.071799, 0.619143, 0.2035917, 1.676034, 0.3604806, 0.133038, 
    -0.2233906,
  10.08576, 15.52411, 20.85332, 11.63595, 1.791251, 0.366443, 1.063257, 
    0.8512682, 2.032284, 3.295501, 0.9763303, 4.263405, 4.514638, 
    -0.02770502, -0.2838835,
  27.45222, 33.79779, 36.80569, 26.45945, 18.28937, -1.29635, -0.1167192, 
    0.5073723, 1.142544, 3.044527, 3.05782, 3.302544, 4.033011, 3.136504, 
    1.280124,
  54.04808, 63.13784, 96.67687, 94.26723, 63.16162, 27.40109, -0.2738751, 
    -0.2678546, 0.2802677, 1.444661, 0.8855215, 1.124036, 1.943436, 2.809242, 
    2.706087,
  54.14397, 58.71478, 101.7011, 149.0736, 146.1932, 94.85861, 65.01464, 
    0.7948853, -1.268608, -0.003814073, 1.295211, 1.52725, 0.7339991, 
    2.02069, 2.959548,
  59.96632, 59.48887, 91.94228, 137.4881, 156.2213, 147.4291, 104.8511, 
    44.02245, 13.96584, 16.0402, 10.10425, 4.404938, 0.6095792, 0.625601, 
    1.09404,
  68.47215, 67.17393, 87.24362, 126.3329, 141.8921, 142.9786, 130.2811, 
    62.18128, 27.39512, 15.2422, 11.70349, 2.592869, 0.9247746, 0.1183376, 
    0.3746546,
  70.18999, 62.10947, 80.71021, 116.2985, 132.4234, 132.093, 122.0757, 
    105.5466, 43.6262, 4.821988, 2.290868, 1.479908, 0.8221701, -0.3191255, 
    -0.04507909,
  61.83972, 56.03202, 81.89761, 111.8281, 122.4777, 116.9855, 109.4424, 
    86.3607, 11.37132, 0.471317, 0.8673828, 2.235812, 0.7680944, -0.2824779, 
    -0.4952983,
  44.54456, 41.33125, 61.87999, 88.78664, 100.3192, 89.33984, 73.04132, 
    33.68549, 2.164055, 3.817274, 16.62353, 7.678683, 4.073222, 1.24646, 
    -0.0002392718,
  5.404897, 8.487907, 5.315319, 3.563461, 1.646193, 1.098958, 5.541072, 
    3.471275, 4.955183, 1.044714, 0.4324035, 2.138086, 0.780611, 0.283708, 
    -0.2702653,
  2.165627, 5.983566, 5.533259, 5.268647, 1.904035, 0.2359195, 0.9517161, 
    0.904033, 3.216601, 4.088559, 2.021407, 4.880505, 5.170397, 0.03081079, 
    -0.2668653,
  28.74813, 12.01199, 9.783665, 15.8192, 16.8573, -0.8991542, -0.09182227, 
    0.6437547, 2.458055, 3.561493, 4.113936, 3.946652, 3.973447, 3.729563, 
    1.245814,
  57.22603, 34.88296, 35.326, 53.30899, 55.37593, 28.28452, -0.4980192, 
    -0.2021589, 0.7558404, 1.751584, 1.730412, 2.146008, 2.379544, 3.019785, 
    3.068314,
  61.75705, 36.32748, 37.17508, 91.89911, 102.0839, 75.94101, 63.94812, 
    0.8292408, -1.112996, -0.07514083, 1.141065, 2.542381, 2.134119, 
    3.033406, 3.448534,
  61.31998, 42.05828, 34.56693, 79.24259, 124.8896, 121.8721, 94.26723, 
    43.29134, 15.02395, 20.31949, 10.61833, 4.887038, 2.670412, 1.887479, 
    1.664036,
  53.62528, 46.00749, 33.22266, 66.66516, 111.9665, 120.4312, 113.5221, 
    51.59859, 24.31259, 20.89156, 14.1416, 4.166949, 2.818989, 1.22363, 
    1.358363,
  47.03439, 42.46827, 30.6738, 62.27616, 106.1074, 116.4902, 115.2927, 
    97.83349, 38.53641, 8.164229, 4.771861, 2.842199, 1.926087, 0.6547892, 
    0.8034915,
  43.93756, 46.09156, 33.86147, 63.88824, 102.002, 105.5986, 110.8208, 
    91.49403, 15.72137, 1.342314, 1.455084, 2.57056, 1.628764, 0.3454459, 
    0.2870009,
  41.35513, 33.95655, 25.20681, 60.30651, 88.57633, 87.41327, 75.60003, 
    34.6511, 1.738208, 3.908272, 16.47932, 5.951554, 3.472338, 2.074309, 
    0.9644018,
  12.34895, 23.72948, 16.95962, 9.878695, 0.6679932, -1.05396, 2.872085, 
    3.445674, 6.585554, 1.205214, 0.07100741, 2.049047, 0.6086206, 0.2973502, 
    -0.1855525,
  20.05295, 23.57977, 18.97778, 8.325895, -0.8929101, -1.323132, 0.3703938, 
    0.8752767, 3.970492, 4.943547, 1.950812, 4.722537, 4.736569, 0.188696, 
    -0.09056067,
  59.01222, 46.62051, 28.9908, 13.2154, 9.575144, 0.7798293, 0.1197056, 
    0.5853129, 2.342686, 3.842464, 4.182871, 3.663407, 3.381278, 2.997191, 
    1.115695,
  77.25736, 73.01712, 67.31779, 43.44421, 38.577, 28.41826, 1.600067, 
    -0.198049, 0.6989279, 1.589285, 1.73758, 1.994432, 2.084929, 2.555553, 
    2.66598,
  68.50197, 62.60684, 63.49672, 68.01614, 58.40202, 60.09602, 55.62456, 
    1.763298, -1.260073, -0.1724547, 1.051453, 2.424623, 2.254079, 2.611152, 
    2.619644,
  47.61856, 49.89893, 54.11147, 61.52852, 86.07258, 92.47985, 70.46204, 
    34.0975, 15.2597, 24.30936, 11.69364, 5.142875, 3.357468, 1.819349, 
    1.370107,
  33.54693, 38.50911, 45.90456, 53.47615, 80.75874, 95.82201, 77.83356, 
    33.64388, 19.63742, 28.40892, 16.5892, 5.519827, 3.795207, 1.556324, 
    1.043219,
  47.08414, 37.4615, 43.01911, 54.21694, 81.76984, 96.63639, 92.35482, 
    80.64072, 30.20992, 7.724949, 5.027131, 3.886546, 2.997612, 1.176997, 
    0.6731918,
  62.57632, 51.70843, 56.54266, 67.57208, 88.67961, 88.04257, 93.71989, 
    87.59763, 13.80927, 1.830784, 1.726526, 3.143086, 2.285978, 0.9743386, 
    0.314999,
  55.88556, 48.05275, 56.46151, 67.78201, 82.72865, 83.65289, 75.49938, 
    33.98481, 2.896862, 4.038934, 15.02788, 5.033606, 4.224604, 2.806138, 
    1.725357,
  11.38116, 24.2413, 15.36138, 11.34831, 4.402399, 1.915132, 4.670912, 
    -0.1791007, 2.046124, 0.4612974, 0.4832015, 2.467858, 0.6645582, 
    0.2374889, -0.2195697,
  18.89774, 13.70928, 11.51379, 6.917161, 0.4816031, -0.4234578, -0.9065337, 
    -1.571236, 0.4073871, 4.412258, 2.658629, 5.448883, 4.732843, -0.0682177, 
    -0.3144331,
  43.90399, 31.6975, 21.27318, 5.178652, 2.873506, -3.031407, -1.370559, 
    -0.06736714, 0.136452, 3.523693, 5.180663, 3.91813, 3.101057, 1.931496, 
    0.5061494,
  53.45724, 54.36798, 55.24842, 41.37078, 29.14405, 18.07778, 0.2433975, 
    -0.8256311, 0.348949, 1.490141, 1.860195, 0.939934, 1.002515, 1.17886, 
    0.6895242,
  48.56254, 42.59452, 50.04825, 66.57832, 49.18287, 46.43287, 41.32749, 
    -0.07078708, -1.023355, -0.02950838, 0.7139902, 0.9331197, 0.7702572, 
    0.9060776, 0.7420447,
  44.89578, 34.49855, 40.97416, 63.76461, 88.18393, 77.77001, 53.47974, 
    28.28688, 15.70396, 24.32817, 13.61855, 4.163005, 1.936447, 0.5139781, 
    0.3514528,
  42.09401, 31.71765, 39.11277, 64.08595, 86.96937, 86.42196, 69.01888, 
    28.08468, 19.93396, 32.91476, 20.97504, 5.107639, 2.478744, 0.4627276, 
    0.1288947,
  47.49926, 35.60483, 48.46841, 74.52361, 82.31356, 85.63415, 76.26558, 
    60.30485, 22.56143, 6.502588, 3.668226, 3.434296, 1.907518, 0.4140908, 
    0.1137049,
  93.53347, 76.49297, 82.31866, 83.79047, 81.98648, 73.93304, 70.71094, 
    64.18654, 6.811677, 1.257604, 0.5246304, 2.696961, 1.779478, 0.7065251, 
    0.3333307,
  126.4319, 102.3365, 92.29211, 81.84277, 74.89867, 72.86861, 61.74554, 
    34.00574, 3.976048, 3.192465, 12.78266, 4.624208, 3.494203, 2.15305, 
    1.460148,
  13.83617, 25.94479, 19.25668, 16.78261, 7.600307, 6.853483, 11.80828, 
    5.844065, 3.142127, -2.357169, -0.9584278, 1.924985, 0.5590072, 
    0.3432139, -0.6671764,
  20.67979, 10.02046, 10.1259, 6.128447, -1.134687, 0.3003163, 1.557444, 
    -0.5843254, -0.7728994, -0.1459848, 0.1090207, 5.840993, 6.294119, 
    -0.6658747, -0.6942703,
  38.06145, 27.02188, 17.53258, 4.754651, 2.821937, -3.121923, -0.5931786, 
    -1.08818, -1.89172, -1.090536, 1.589399, 2.762485, 3.219573, 4.384929, 
    1.535175,
  43.91561, 38.84271, 34.69165, 19.15962, 14.24852, 14.366, -2.349682, 
    -0.8828033, -0.6170915, -0.8806016, -0.5449321, 0.7699458, 2.292385, 
    2.923526, 2.905548,
  57.08944, 35.02924, 26.62428, 25.58481, 18.04945, 28.24698, 25.68878, 
    1.846705, -1.411829, -0.3384869, -0.02351947, 1.657039, 2.643474, 
    3.316209, 3.050165,
  73.70503, 43.84743, 25.02929, 16.33171, 25.57077, 41.20292, 34.36587, 
    20.12507, 10.9604, 17.85535, 10.21513, 4.181758, 3.402912, 1.695614, 
    0.7198355,
  100.7815, 87.64117, 44.47017, 30.37009, 48.13451, 63.54127, 53.92683, 
    21.61746, 13.77804, 27.35834, 19.08873, 6.432719, 3.403971, 1.154366, 
    0.3013713,
  105.9972, 108.571, 97.47346, 84.28847, 82.19557, 79.1996, 71.38497, 
    54.7188, 15.30219, 4.022578, 5.030489, 4.147271, 2.313595, 0.5010047, 
    0.2007132,
  101.7465, 98.67638, 97.25077, 89.6267, 80.46864, 70.81818, 71.21621, 
    57.75574, 5.631276, 0.5062013, 1.697488, 2.280216, 1.280911, 0.2912831, 
    0.4232097,
  99.90714, 92.38465, 88.55293, 80.25062, 71.60961, 66.25438, 58.67944, 
    30.72969, 3.482317, 2.098287, 9.653114, 2.874056, 2.191787, 0.7981873, 
    1.071755,
  5.183647, 12.72801, 8.686093, 10.1685, 3.876512, 6.888312, 12.94714, 
    4.864653, 1.492113, -1.173732, -0.2964106, 2.256327, 0.2866695, 
    -0.06687397, -0.8869894,
  10.38618, 9.655508, 7.722704, 5.324511, 0.1497669, 5.126477, 5.931157, 
    1.15372, -0.2251447, 0.2862049, 2.173511, 6.889573, 5.426901, -1.171602, 
    -0.8501444,
  34.01496, 21.46774, 13.81747, 8.756476, 3.708832, -1.433366, 2.281929, 
    1.506517, -0.01103867, 0.5946547, 3.762893, 4.186195, 3.61023, 2.919265, 
    0.7757559,
  59.25295, 57.30571, 47.73619, 24.98057, 10.69937, 11.73436, -1.497935, 
    -0.4029495, -0.3808522, -0.005865283, 0.56893, 1.124302, 0.8598834, 
    1.255444, 3.409332,
  67.47971, 63.59373, 57.71818, 38.94672, 20.31402, 22.34825, 24.44481, 
    1.744249, -1.487697, 0.1535186, 1.098534, 1.144915, 0.7355295, 0.9820973, 
    4.21455,
  72.46187, 77.00417, 71.57227, 59.30402, 40.34632, 29.67512, 26.67362, 
    15.71203, 9.735662, 14.79052, 11.2427, 3.990831, 1.73896, 0.2594633, 
    0.7509582,
  69.20894, 90.30524, 87.58894, 81.16476, 76.23361, 63.34146, 45.4051, 
    13.42008, 6.573867, 17.60049, 16.52743, 5.058398, 2.899371, 1.092824, 
    1.744892,
  62.21234, 79.46809, 83.87737, 82.89995, 82.15086, 78.98485, 68.93133, 
    44.04487, 5.798854, 0.8609774, 2.676554, 2.592448, 3.143722, 1.448665, 
    1.256547,
  65.25019, 72.8667, 82.04556, 81.97169, 79.0891, 71.77863, 71.31044, 
    45.6724, 3.593518, -0.1287052, 0.7006037, 2.481032, 3.360813, 2.274962, 
    1.153378,
  67.74423, 65.95383, 71.81374, 74.01299, 69.66163, 63.60931, 54.18094, 
    26.35069, 3.064302, 1.391166, 7.916646, 4.329821, 5.401638, 4.175929, 
    2.736255,
  3.899038, 9.17772, 5.761263, 10.69158, 5.396436, 2.727552, 6.928013, 
    4.602211, 2.988006, -0.466958, 0.7963279, 3.504035, 0.6924875, 0.6660094, 
    -0.7557452,
  6.648255, 4.342385, 3.847083, 8.34293, 2.646766, 2.873374, 3.380169, 
    2.613879, 2.168083, 2.553164, 4.972426, 8.102619, 5.963445, -0.5647514, 
    -0.5868906,
  21.8222, 29.47264, 13.2507, 6.05553, 5.407341, -0.8542578, 1.344201, 
    2.160426, 1.303005, 1.840725, 6.362077, 6.336686, 3.803827, 3.366808, 
    0.938206,
  28.06132, 48.28136, 62.04911, 47.35456, 13.3193, 5.798284, -0.5296165, 
    0.47923, 1.74609, 0.423499, 1.432031, 2.501482, 2.476824, 3.858428, 
    4.148554,
  30.17177, 41.24666, 59.73441, 69.56509, 50.51907, 36.43223, 15.33461, 
    0.9014785, -0.1413856, -0.576661, 1.749107, 3.965732, 3.099115, 4.694294, 
    5.985976,
  39.98779, 40.19173, 58.15473, 67.97734, 70.54916, 63.42082, 37.28935, 
    17.73143, 7.190026, 8.761929, 7.479939, 5.152677, 5.589265, 2.816618, 
    3.101128,
  55.38453, 47.78082, 59.24928, 63.34394, 66.35192, 65.34595, 56.4798, 
    24.27891, 11.88127, 9.442648, 9.255536, 5.569592, 5.259742, 2.562783, 
    2.776191,
  60.92366, 53.31963, 59.89239, 59.1121, 61.85505, 61.14209, 54.43132, 
    35.17119, 7.457906, 0.8870412, 2.513535, 4.53313, 4.983537, 1.494376, 
    1.680545,
  57.949, 61.08184, 66.79913, 58.33969, 57.82745, 50.78621, 46.76939, 
    29.76441, 3.134448, 0.5116138, 0.888831, 3.313326, 2.363811, 2.065266, 
    2.766559,
  55.48414, 62.52527, 59.02903, 51.84928, 48.92208, 43.27856, 29.23684, 
    15.44535, 2.867059, 1.467955, 3.276219, 3.920672, 5.080344, 5.743951, 
    5.568815,
  2.435209, 1.499518, 1.040914, 0.1595782, -0.6345119, -0.1744883, 4.714468, 
    2.097344, -0.5553514, -3.053376, -0.8289124, 0.7122684, -0.2814075, 
    0.1930377, -0.3476243,
  7.351909, 0.7018722, -0.3369588, -1.406151, -3.136816, 0.3074705, 1.527739, 
    0.7096329, -0.3100904, -1.927197, -0.3944449, 3.159023, 2.988323, 
    -1.052958, -0.7505062,
  38.8214, 28.67903, 11.87147, 0.3597491, -3.368663, -5.513414, -0.8082934, 
    0.4221407, 0.01756535, -0.7601136, 0.7804992, 2.291548, 1.213281, 
    1.151809, 0.2293782,
  46.81808, 49.40308, 59.82494, 46.18501, 14.11111, 3.17097, -3.300416, 
    -2.180513, -0.291216, 0.05891332, -0.1590987, 1.193045, 1.355539, 
    1.600671, 2.564805,
  50.18024, 51.86064, 59.28167, 64.73302, 46.61271, 30.5472, 11.04847, 
    -2.364887, -1.482873, -0.0430776, 0.6779694, 1.624109, 0.8505027, 
    1.967148, 3.485492,
  67.96906, 66.32769, 66.3128, 62.36168, 57.80955, 42.6006, 20.14351, 
    6.021194, 2.219466, 7.117272, 3.906554, 1.720248, 1.953739, 1.337427, 
    1.296786,
  81.14077, 78.29267, 70.48584, 59.35223, 49.11701, 43.47285, 41.67857, 
    6.770081, 2.684553, 10.10499, 3.368714, 1.492151, 1.985837, 1.747409, 
    1.830149,
  74.66233, 77.99712, 66.54198, 59.14003, 44.80952, 46.12711, 48.17435, 
    18.71973, 3.146075, 3.153499, 1.324597, 1.025485, 2.157059, 0.9869643, 
    1.029231,
  70.4637, 71.6287, 70.24158, 64.60006, 42.98298, 40.32517, 50.24158, 
    16.34215, 1.929987, 2.138925, 0.9733394, 1.156568, 0.9525593, 1.544628, 
    2.055114,
  50.54245, 43.58863, 50.13107, 55.59089, 37.90025, 37.1836, 35.79466, 
    5.233744, 2.345862, 2.293691, 2.437469, 1.531, 2.962146, 4.640205, 
    5.039995,
  1.75976, 3.15207, 1.780996, 1.254351, -0.3531309, 2.040078, 5.921021, 
    2.892453, 2.817059, -0.08675341, 2.39088, 2.067647, -1.31549, -1.379833, 
    -2.514129,
  6.828779, 2.569663, -0.01877049, -0.2749247, -0.9954996, 4.956987, 
    4.286738, 1.911723, 2.084765, 1.845596, 1.472567, 4.168598, 2.925955, 
    -1.801167, -2.370799,
  22.09287, 26.90104, 16.68692, 4.62763, 0.3800509, -0.481227, 5.099034, 
    4.145948, 4.785136, 1.539754, 2.123123, 7.245882, 6.949527, 7.09549, 
    2.427346,
  36.52017, 40.43914, 41.96263, 40.81761, 14.52163, 2.005637, -1.341529, 
    0.4519238, 3.674053, 4.459483, 3.742679, 4.563221, 7.430385, 7.506978, 
    5.315083,
  46.24939, 30.52752, 36.21714, 50.60452, 49.1669, 44.41604, 7.026293, 
    -2.319753, 1.972545, 1.429634, 3.485823, 3.486864, 4.50065, 6.087221, 
    4.820377,
  43.73701, 26.2527, 33.95047, 49.89194, 55.91448, 57.43909, 37.75434, 
    13.5756, 7.994363, 10.57634, 2.664799, 5.344742, 4.739399, 3.622988, 
    2.468236,
  42.55763, 34.03909, 35.60477, 41.23074, 48.81012, 53.76504, 53.67685, 
    15.30097, 8.972592, 11.696, 4.10859, 2.533807, 4.381945, 1.819244, 
    2.087968,
  41.18981, 38.41803, 37.69562, 37.32046, 45.18844, 49.59167, 45.26008, 
    24.16005, 7.220518, 5.642119, 1.815897, 1.421811, 1.076081, 0.2475117, 
    -0.1472333,
  38.96841, 38.51645, 43.5158, 37.28323, 38.00712, 35.44163, 37.24181, 
    18.58155, 3.342819, 2.119658, 1.351051, 0.67397, 0.7215001, 0.1337224, 
    1.071651,
  27.09497, 19.93931, 26.69957, 26.28618, 27.98245, 26.2296, 21.74064, 
    7.966285, 2.512035, 2.541886, 2.717835, 1.352167, 1.186508, 1.822415, 
    2.276566,
  1.813704, 3.233923, 1.42038, 0.8710449, 0.9309641, 1.522079, 3.369287, 
    -0.3714291, 1.860776, -0.7279969, 0.3405536, 2.48272, -0.5630535, 
    -0.4231899, -0.9576259,
  12.94027, 3.282207, 0.8623229, 0.7945129, -0.2858466, 1.443991, 1.016557, 
    -0.903657, 1.595984, 0.8944393, 1.426157, 3.540465, 4.153048, -1.071944, 
    -0.8471001,
  51.39279, 25.97791, 9.906734, 2.649966, -0.01392651, -2.902716, 3.534369, 
    1.847623, 1.56935, 1.697822, 2.918848, 3.82763, 3.629143, 6.112501, 
    1.769353,
  58.07429, 33.68622, 19.87171, 16.4403, 5.761203, -0.7022638, -2.301128, 
    -1.253146, 1.001728, 1.573573, 2.107579, 4.471217, 3.237418, 3.663099, 
    4.316433,
  56.22093, 23.22289, 16.17121, 21.1525, 23.08997, 13.3852, 4.555724, 
    -2.329021, -1.595542, 0.3280798, 3.322966, 3.84945, 3.262823, 3.145422, 
    7.21811,
  40.84507, 14.47975, 13.82396, 21.88189, 28.8143, 23.5573, 13.53786, 
    5.613025, 3.350636, 1.539751, 3.724298, 3.770087, 1.963499, 2.115255, 
    1.297411,
  40.07626, 25.51195, 17.00105, 12.30455, 29.22553, 26.36129, 27.28509, 
    8.98771, 7.761366, 3.230379, 3.863431, 2.082626, 1.547749, 0.207461, 
    0.07938775,
  38.482, 25.70419, 21.38906, 18.47438, 30.68266, 29.23041, 23.47178, 
    13.91358, 7.671986, 2.767738, 1.346714, 1.806335, 1.637243, 0.5773134, 
    -0.2078891,
  33.09498, 23.80731, 29.43639, 25.79855, 27.27843, 14.7153, 23.428, 
    15.06896, 9.159411, 2.517804, 1.701407, 1.588092, 0.5893769, -0.09988259, 
    0.1385928,
  23.09861, 17.68579, 22.22136, 22.43556, 17.1166, 12.4227, 13.56156, 
    13.12247, 11.40312, 0.9617061, 2.115476, 3.493823, 1.164714, 1.269663, 
    0.7063378,
  6.575338, 6.432883, 5.418181, 4.692688, 1.660913, 0.1987141, 1.532393, 
    0.04169042, 2.956045, 0.6849058, -0.5398725, 1.856838, 0.8340239, 
    -0.441386, -0.8446481,
  16.07882, 8.331029, 6.300362, 3.24943, 0.930096, 2.774775, 3.984691, 
    -2.340515, 0.9000363, 1.61772, -0.03579338, 2.956389, 3.783712, 
    0.07773563, -0.3962367,
  52.99281, 26.65591, 13.87701, 3.79846, 1.563375, 0.3269563, 5.923834, 
    1.454613, -0.3102602, 1.521006, 1.768864, 1.741721, 3.514367, 5.881544, 
    2.999811,
  62.69874, 38.33881, 28.03369, 20.46, 6.055729, 2.429345, -0.4092607, 
    -3.160959, 1.71267, -0.5792942, 1.319132, 2.702005, 1.929079, 3.351481, 
    4.347421,
  60.48857, 30.62448, 22.34435, 20.19608, 15.93394, 15.7582, 3.846551, 
    -0.2937633, 1.235642, -0.6556017, 0.8781714, 1.436438, 1.310595, 
    0.7952416, 1.153039,
  53.34589, 28.20593, 20.6624, 16.92747, 19.54651, 22.50174, 15.35082, 
    4.752454, 2.856608, 2.951216, -1.135097, 0.6584123, 0.617467, 0.1742976, 
    0.2268053,
  49.9691, 30.33211, 22.62495, 17.2753, 24.50376, 26.32432, 27.03874, 
    10.28474, 7.575606, 3.716303, 1.17684, -1.600904, 0.05190624, -0.7273785, 
    -0.7341955,
  48.85194, 35.97629, 29.43616, 25.78283, 29.75191, 28.82881, 20.80861, 
    14.98266, 8.090235, 2.726654, 2.455, -1.458659, -0.3237881, -1.362072, 
    -1.479417,
  51.41874, 42.77354, 35.73101, 24.88937, 19.81708, 20.10754, 16.78421, 
    11.25112, 8.539948, 5.734523, 3.952251, -1.621395, -0.8462371, -1.847281, 
    -1.887854,
  49.38015, 35.07935, 17.52637, 22.75365, 22.56615, 19.73224, 10.14246, 
    3.488858, 9.247434, 2.383208, 3.712861, -0.1987698, -1.064581, -1.870129, 
    -1.166813,
  12.22508, 14.01371, 10.55903, 5.251404, 1.961942, 0.7817435, 1.760427, 
    0.5178299, 3.481184, -1.150722, -1.287246, 0.03928632, -0.5484998, 
    -0.1726217, -0.5957912,
  22.8591, 18.86709, 8.781142, 2.060932, 0.8685549, 1.817579, 2.003814, 
    2.583795, 0.6694894, -0.04367967, -2.227202, 0.3560876, 1.417251, 
    -0.8509544, -1.083931,
  56.15536, 33.5559, 21.87171, 5.928852, 2.422089, -0.2192911, 3.648763, 
    3.257291, 2.126432, -0.1197812, 0.6363172, 1.320962, 1.424607, 1.043934, 
    -0.5362309,
  73.09976, 60.7655, 50.5693, 33.72653, 13.15106, 4.014913, 1.088654, 
    1.484929, 1.56562, -0.4281753, -0.4162622, -0.4136262, 1.540546, 
    1.637417, 0.8682584,
  70.62804, 50.89082, 46.21961, 47.12318, 47.41882, 43.09353, 15.34427, 
    -0.05361024, 3.126911, 0.9477517, 2.840892, 1.602696, -0.2599959, 
    -0.8831921, -0.04135275,
  62.68394, 52.8858, 52.08575, 53.29713, 56.65408, 51.76535, 38.50487, 
    13.44943, 12.30747, 4.600828, 3.165449, 0.143951, -0.7430436, -2.650143, 
    -2.427988,
  64.46273, 63.24615, 60.34185, 51.11412, 52.03843, 49.09736, 43.97701, 
    21.91533, 11.40303, 7.068031, 3.206474, 0.2635052, -0.9757362, -2.471223, 
    -3.879834,
  73.00603, 72.39917, 65.66953, 49.31604, 48.79176, 44.44981, 28.86527, 
    19.41625, 10.63785, 5.86399, 4.034077, -1.551673, -2.871127, -3.733658, 
    -5.410429,
  88.75619, 82.76125, 68.7824, 45.41068, 30.93999, 23.98317, 21.73852, 
    14.20187, 9.373736, 4.282205, 2.621496, 0.001373522, -1.954821, 
    -5.103332, -5.800098,
  81.30153, 61.73955, 45.77644, 23.83769, 16.5107, 10.55713, 13.35587, 
    4.853877, 11.26841, 3.636683, 4.39241, 2.029356, -0.3994178, -2.688092, 
    -3.973614,
  7.850387, 11.39418, 7.551475, 3.677087, -0.2523759, 1.001588, 3.711318, 
    1.513677, 0.3686389, -2.381731, -1.086272, -0.3081718, -3.447302, 
    -2.371452, -3.397798,
  17.96573, 11.11967, 7.434206, 1.170885, -0.1163275, 1.230591, 2.912275, 
    1.821283, 1.013014, -2.29414, -1.237043, 1.198811, -0.7908339, -4.008371, 
    -4.470683,
  41.93896, 24.28555, 19.80186, 5.747272, 2.178439, -1.57813, 4.557709, 
    1.797949, 2.98475, 0.9967035, -1.125303, -0.2281228, 0.4758794, 1.263509, 
    1.400398,
  62.80862, 60.41133, 58.02987, 40.0605, 14.74758, -0.5184395, -3.893912, 
    0.4526912, 4.902908, 4.967141, 2.874815, 3.936849, 4.62953, 4.909822, 
    2.959107,
  72.46993, 57.56159, 53.64738, 53.38183, 52.60046, 44.63266, 16.06561, 
    4.292862, 12.58871, 4.26583, 9.261398, 7.193728, 4.788824, 3.680939, 
    3.898804,
  79.40703, 64.70467, 57.67032, 53.49766, 55.41567, 52.44248, 41.4352, 
    14.55321, 13.82872, 4.393772, 4.877415, 6.192197, 5.312916, 6.176622, 
    5.313393,
  85.20586, 75.07565, 63.12983, 53.10936, 47.90722, 44.51086, 35.27472, 
    17.78139, 8.943485, 4.180688, 7.248631, 7.716616, 7.346115, 7.045784, 
    4.796766,
  78.31598, 72.3533, 61.35637, 47.32912, 40.73555, 34.32608, 16.58623, 
    5.481494, 6.779449, 8.993547, 9.077344, 7.792743, 8.803036, 6.226724, 
    6.893404,
  76.13242, 69.62039, 62.26483, 44.15334, 30.46054, 14.1625, 5.400001, 
    2.342519, 10.14131, 18.0301, 16.22876, 5.938043, 3.734259, 3.13833, 
    4.194368,
  62.9539, 50.96459, 43.68787, 25.42104, 10.20332, 1.009764, -1.208714, 
    1.08524, 12.84785, 5.857971, 25.2241, 13.68259, 5.97333, 3.538811, 
    3.091584,
  9.018078, 10.77715, 11.04554, 7.453901, 1.108978, 2.762038, 7.002882, 
    -0.6503437, -1.536595, -3.019669, -1.575047, 0.2672043, -2.239011, 
    -1.794592, -1.659637,
  16.01173, 14.22042, 9.239686, 4.077148, 0.1600491, 3.734255, 6.592985, 
    -0.3411807, -1.047285, -2.178634, -1.410621, 1.458638, 0.7391939, 
    -1.470661, -1.696468,
  38.19559, 25.00936, 19.6281, 9.585414, 5.089429, 0.593056, 8.044885, 
    3.772893, 0.4452186, -1.372459, -0.3847176, 0.04525021, 1.332554, 
    0.7441847, -1.613763,
  65.522, 60.83107, 59.59883, 43.81694, 22.15567, 7.638948, 1.780224, 
    4.471048, 1.596539, -1.519086, -0.02040853, 0.1594061, 0.3389495, 
    -0.283601, -1.503618,
  80.58009, 63.46978, 59.13079, 57.62725, 54.66072, 45.52105, 21.43842, 
    3.21863, 2.25485, 7.74108, 10.44473, 0.3508781, 0.1155617, 0.6057773, 
    1.741912,
  93.06045, 75.54879, 64.05084, 54.76829, 54.36369, 53.78077, 51.91803, 
    19.56646, 6.483203, 9.267973, 7.886806, 4.487195, 3.643326, 2.014488, 
    0.8005832,
  100.8877, 84.89015, 69.5838, 56.36555, 55.87269, 54.48233, 53.1521, 
    38.5017, 14.98616, 10.22228, 8.225001, 5.512803, 3.412123, 2.139031, 
    0.4484325,
  92.80727, 79.3015, 67.14082, 56.68347, 54.06336, 54.41021, 46.20864, 
    34.42593, 15.0808, 8.200409, 9.315218, 5.654869, 5.737627, 2.600223, 
    1.21774,
  82.32118, 72.36709, 63.74429, 49.27013, 43.56567, 35.58694, 35.3182, 
    25.17199, 13.5621, 16.52664, 19.60349, 9.255196, 3.973143, 1.419564, 
    1.556426,
  61.91172, 48.70434, 42.09173, 31.61938, 23.44073, 21.34387, 23.15768, 
    13.63381, 16.97772, 11.278, 20.98499, 9.986096, 3.764356, 2.033145, 
    0.8272324,
  7.643978, 9.235319, 10.15579, 7.827963, 1.970072, 1.41857, 2.889863, 
    -1.526411, -1.339511, -1.975543, -0.5376485, 1.643853, 0.2351148, 
    -0.4128199, -1.490507,
  10.96478, 9.150533, 8.35072, 4.428903, 0.2530223, 1.844547, 4.181346, 
    -0.9527066, -0.5089256, -0.5451484, 0.5212233, 2.908957, 1.662556, 
    -1.301691, -1.94733,
  43.6748, 25.53168, 14.25606, 6.142734, 1.767628, -2.687583, 4.996476, 
    3.255873, -0.2244196, -0.8003115, 1.232925, 1.437861, 1.547228, 2.7576, 
    0.2869851,
  63.57059, 56.72898, 47.04182, 30.00669, 8.073073, 0.2412503, -1.832915, 
    2.904889, 2.092639, 0.4461304, 0.8298481, 0.5038842, 0.4132968, 
    -0.4811483, 0.1547062,
  65.80724, 47.72176, 38.19818, 29.61188, 22.96041, 13.40199, 5.845812, 
    -0.4594698, 2.019348, 3.454977, 3.365364, -0.4398556, 0.09699421, 
    -0.07197373, 2.092665,
  60.39717, 46.66221, 31.78154, 23.48742, 23.05187, 21.80632, 17.85914, 
    12.8472, 1.897609, -0.3777013, 1.477907, 1.05799, 2.736135, 3.077568, 
    3.471955,
  58.04517, 45.27096, 30.00443, 20.5348, 20.60451, 21.09889, 23.02508, 
    14.44758, -0.9386146, 0.184706, 1.180655, 2.289254, 3.612411, 4.175875, 
    3.650101,
  50.88394, 35.25235, 24.06096, 20.80255, 17.85658, 24.50613, 18.81511, 
    12.82308, 1.956903, 2.434424, 2.15794, 2.362243, 4.532862, 3.73765, 
    3.379681,
  38.24327, 33.11184, 24.81027, 15.46826, 14.33457, 13.03548, 15.89174, 
    8.751036, 8.471144, 13.14837, 19.73645, 5.454602, 2.930194, 2.651608, 
    4.429123,
  26.68371, 16.25958, 13.14424, 9.515829, 8.223699, 11.89366, 8.537031, 
    8.322426, 14.26101, 8.943339, 22.4901, 5.013624, 1.833764, 1.884833, 
    2.46417,
  1.626505, -0.157152, -2.587794, 0.1977393, -2.365137, 0.6808322, 0.4363789, 
    -2.863973, -4.626109, -5.282138, -3.834164, -1.679859, -1.299588, 
    -0.4116406, -0.7168422,
  1.076251, -1.923954, -0.1793424, 0.9558343, -3.036156, -0.07858675, 
    -0.1941225, -2.7723, -4.351609, -4.693684, -2.592196, -0.9884319, 
    -0.5648823, -2.447341, -1.792405,
  16.39749, 2.73616, 0.9160926, 2.822285, -0.9227214, -2.640282, -1.75264, 
    -2.135846, -3.386327, -3.058849, -0.7416697, -1.146829, -0.9414723, 
    -0.04988914, -1.335372,
  27.39722, 13.35059, 10.48034, 2.954791, -0.1037834, -2.043643, -1.175703, 
    -3.315588, -2.735032, -0.9743633, -1.099424, -1.045072, -0.3118467, 
    -0.7934534, -1.089383,
  20.92707, 7.451521, 4.440421, -0.7851969, -3.821951, -3.826364, -2.053238, 
    0.6282496, 0.5919082, 0.3871288, 3.020656, 2.231344, 1.466076, 
    -0.6892903, -0.8279525,
  20.76311, 10.70467, 1.058484, -3.491356, -2.977879, -1.710162, 1.182781, 
    2.355821, 2.656244, 3.048964, 2.505289, 3.349787, 1.885191, 0.8210471, 
    0.4431589,
  18.47518, 9.144469, -0.08488012, -4.226247, -2.746601, 2.834538, 8.149645, 
    7.596794, -0.7854706, -0.382321, -0.6938693, 1.271089, -1.095223, 
    -0.1410411, 0.7036033,
  20.66465, 7.81869, -0.4774307, -2.30922, 0.1645658, 8.649256, 10.12191, 
    10.9256, 4.010998, 2.419244, 3.492096, 0.1299944, 2.375196, 2.091136, 
    0.4706825,
  12.58478, 5.260535, 2.639871, 0.5342295, 3.8884, 3.989344, 9.206285, 
    9.60856, 7.718661, 7.036959, 7.635525, 4.665065, 4.233239, 0.8802065, 
    2.819674,
  5.816957, 1.155093, 2.222514, 0.2008693, 1.214052, 3.420396, 4.750662, 
    3.530115, 6.790024, 3.34013, 12.44898, 9.182978, 2.870599, 1.482044, 
    0.8482374,
  4.903165, 5.998007, 2.363876, 1.31142, -2.964505, -3.071554, -1.406302, 
    -3.188286, -5.689812, -3.990845, -6.924283, -6.275736, -7.003881, 
    -2.95203, -4.030611,
  8.34295, 3.937001, -0.944772, -3.43071, -3.988939, 1.946086, -1.239746, 
    -6.919049, -7.849659, -9.855776, -8.785881, -5.706223, -4.858743, 
    -4.229399, -3.474815,
  54.69243, 26.38986, 10.33014, 0.4711803, 2.71939, 1.541544, 7.298374, 
    -6.981695, -9.06566, -9.048694, -6.840137, -5.548235, 1.161948, 
    0.1550977, -0.2225691,
  79.30001, 64.38274, 49.18232, 25.06607, 6.00966, 6.002729, 4.784188, 
    -1.999281, -4.810891, -4.941515, -1.905724, 2.713062, 1.391408, 
    -0.4060074, -0.4945868,
  89.54347, 60.63388, 44.14243, 32.37734, 22.9546, 15.85623, 6.69173, 
    5.792382, 8.14572, 9.316611, 11.20369, 5.925487, 1.960713, -0.2761218, 
    3.27299,
  94.1323, 65.93013, 41.3963, 26.18207, 20.46601, 14.97147, 9.615466, 
    4.81168, 3.637586, 10.06447, 5.095219, 2.340595, 1.157685, 2.743717, 
    2.648859,
  79.38768, 60.19711, 36.95291, 18.63198, 17.28156, 12.24056, 11.19394, 
    9.02281, 3.532353, -1.071153, -1.086932, 0.1216355, 2.069445, 3.479093, 
    2.129116,
  67.82021, 51.83459, 32.06626, 17.28247, 11.58634, 12.32793, 8.676758, 
    7.292012, 2.030042, -1.771412, -2.314343, 1.769676, 1.274908, 3.115482, 
    2.789776,
  61.09227, 45.57125, 29.80877, 9.221329, 5.424506, 2.000367, 3.412956, 
    1.408714, -1.213799, 1.277075, 5.54247, 2.450085, 2.222856, 2.72857, 
    3.894973,
  40.4322, 24.36454, 14.43414, 2.893696, -1.733174, -1.591292, -1.712387, 
    -3.527731, -1.195574, -2.415206, 4.664673, 1.306085, 3.955405, 2.297874, 
    2.073648,
  6.984534, 11.73732, 7.719885, 4.877561, -0.9635597, 0.1371802, 4.981512, 
    1.675785, 3.214798, 1.287914, 2.105367, 2.052469, -0.793635, -0.3916246, 
    -1.75676,
  17.75848, 12.36057, 1.015459, -1.773596, -2.614132, 6.411448, 10.12586, 
    4.237305, 3.795216, 2.013545, 1.438633, 2.439005, -0.006047727, 
    -1.187926, -2.466514,
  84.88357, 59.7076, 27.93799, 4.791508, 10.7142, 7.497671, 20.89803, 
    12.18564, 6.753211, 3.78937, 0.3964724, -0.4618669, 0.7860574, 1.075681, 
    -0.4312948,
  113.05, 101.3821, 85.42408, 66.6934, 32.58694, 13.76767, 7.967448, 
    21.40243, 6.238531, -3.061912, 0.01065032, 1.358978, 1.62467, 1.198058, 
    -1.137567,
  129.1444, 99.1372, 81.96249, 70.76983, 59.17099, 37.82913, 20.99562, 
    5.420468, 11.88976, 6.883071, 7.891559, 1.822116, 2.115934, 0.4189573, 
    -1.154777,
  133.5298, 103.4775, 80.77534, 65.08003, 54.67845, 39.56319, 29.84733, 
    16.59066, 6.164475, 7.086111, 5.471366, 2.276669, 1.224151, 0.3255824, 
    -1.607568,
  114.7221, 94.48264, 71.42841, 48.08504, 38.77205, 30.50669, 24.4695, 
    14.96484, 7.809525, 3.549786, 2.410255, 1.426457, 0.5204886, -1.132837, 
    -1.390476,
  97.51422, 80.02534, 59.228, 37.19104, 26.02057, 23.20504, 11.61088, 
    6.50558, 3.126206, 0.44941, -0.1026707, 0.2764811, -0.4220562, -1.982721, 
    -0.219417,
  95.81113, 78.58762, 56.51763, 29.53951, 18.73184, 8.28157, 7.706101, 
    4.033734, 1.785909, 1.037547, 1.502794, -0.5257959, -2.314677, -2.608016, 
    -0.2297243,
  66.95355, 48.36655, 34.10338, 13.61543, 6.924318, 4.879791, 3.702683, 
    1.704093, 1.562057, 3.953677, 2.587463, -0.318615, -3.039964, -2.601941, 
    -0.5939938,
  8.433226, 14.76523, 9.931136, 13.84939, 4.595325, 5.056677, 7.54457, 
    1.39725, 2.25457, 0.6846545, 3.832284, 2.816854, 2.043978, 3.68303, 
    2.986075,
  24.44161, 18.62675, 5.091505, 3.243083, -0.5083394, 14.59779, 27.93085, 
    9.404482, 4.3372, 3.525371, 3.986953, 4.879425, 3.903668, 1.29563, 
    2.376209,
  107.2721, 79.11096, 37.98656, 10.92586, 2.102499, 7.763313, 42.86227, 
    16.10644, 5.082078, 3.76889, 3.270571, 3.974495, 4.171533, 4.664287, 
    3.733107,
  132.5238, 128.6175, 114.4006, 96.44434, 43.50419, 6.728018, 6.458217, 
    30.19988, 19.00261, 7.087803, 3.773136, 0.9930974, 3.510649, 4.491348, 
    2.234997,
  139.4191, 118.0734, 105.6508, 92.3395, 83.74704, 52.93619, 28.30206, 
    5.478143, 14.02979, 8.537084, 15.64136, 2.040949, 2.349695, 4.030582, 
    -0.3074164,
  135.8859, 115.8104, 98.78111, 86.68181, 79.96814, 68.80487, 56.00101, 
    31.59575, 8.528331, 9.463281, 8.118515, 1.201321, 0.8904682, 2.844539, 
    2.586166,
  111.5596, 100.524, 82.75582, 67.03834, 64.02609, 59.57596, 54.06664, 
    41.33876, 23.05293, 3.993142, 2.612886, 1.539085, 3.628761, 3.029142, 
    1.975479,
  103.0773, 91.11559, 77.61054, 60.93111, 52.483, 52.75173, 41.73192, 
    36.06158, 22.31095, 5.603849, 2.370614, 0.7347124, 0.5392958, 0.4027804, 
    1.363778,
  98.90613, 91.86177, 80.16806, 54.50221, 38.59829, 28.08579, 29.14231, 
    26.17961, 15.26084, 9.441341, 12.11848, 2.734362, 2.836132, 2.760169, 
    0.2164001,
  85.65278, 80.22507, 72.57728, 48.7252, 29.75609, 18.96057, 10.87392, 
    6.343828, 5.785064, 8.761722, 11.60802, 8.302004, 3.263608, 0.3915396, 
    -1.428494,
  8.598839, 12.60285, 8.82789, 11.8054, -0.9651868, 4.090631, 7.466276, 
    0.3335201, -0.4603038, 0.07416751, 2.354001, 2.625161, 0.5373743, 
    -0.418413, -1.01712,
  29.32501, 13.98756, 5.366831, 0.783029, -2.003118, 11.70432, 23.2676, 
    2.438988, -0.3588927, 0.08873336, 1.647132, 2.810888, 0.4834746, 
    -1.997543, -1.109092,
  91.24198, 78.95042, 48.42895, 14.76437, -0.7778364, -0.8827861, 48.57378, 
    14.71005, 0.9907182, -0.6955885, 2.540988, 2.158676, -0.4018443, 
    -0.137693, 0.507758,
  83.14867, 96.427, 101.1141, 97.14822, 41.56054, 5.385226, 2.954977, 
    36.75001, 15.08702, -0.1767632, -0.7799471, 2.699054, 3.02222, 3.564715, 
    3.805798,
  60.61082, 52.12328, 59.497, 67.70856, 75.59782, 51.81737, 29.24124, 
    6.640471, 11.07547, 9.862411, 17.02239, 7.116921, 3.518059, 1.926052, 
    0.9759572,
  60.95817, 42.01963, 32.60752, 29.2443, 33.56203, 38.56037, 44.5044, 
    38.26422, 2.80108, 4.473489, 6.353438, 8.48274, 6.365528, 4.364683, 
    2.705247,
  81.9411, 66.12932, 54.50425, 46.17118, 47.45642, 46.97384, 50.46146, 
    48.68244, 33.77202, 6.305119, 7.954051, 7.499958, 5.026536, 3.608469, 
    3.010875,
  111.0779, 94.99518, 81.97506, 73.77521, 72.33942, 70.8806, 56.93114, 
    46.06016, 32.08177, 2.213649, 3.860754, 2.472544, 2.746574, 2.035348, 
    1.45874,
  126.5454, 117.5681, 104.887, 87.31127, 76.97518, 63.9777, 52.74137, 
    42.48478, 22.34432, 10.44001, 25.98902, 7.59622, 4.623483, 0.763741, 
    -0.1560046,
  118.8097, 112.3504, 104.8298, 85.87143, 66.84686, 48.52433, 28.16592, 
    12.35269, 13.51187, 9.724479, 18.21206, 8.850883, 2.020109, -0.09405952, 
    -0.4601309,
  10.9514, 17.58259, 16.61627, 17.5868, 1.232492, 4.033365, 9.206289, 
    -1.286613, -2.451065, -2.726454, -1.794955, 0.2845971, -1.449125, 
    -1.339469, -1.850559,
  34.29975, 20.2452, 11.20235, 4.602374, -2.014219, 14.69912, 25.53616, 
    3.694875, -1.895076, -1.703998, 1.30982, 3.324961, -0.2005305, -2.894871, 
    -2.151715,
  56.15651, 50.448, 45.13408, 14.90881, 1.101234, 0.5788496, 43.56945, 
    15.66062, 1.187028, -1.581149, 4.356527, 1.401173, -0.2896102, 
    -0.5815083, -1.215201,
  52.28486, 48.0868, 48.91588, 53.3501, 33.96002, 4.929929, 2.039088, 
    32.76545, 19.79228, 1.851014, 1.338186, 1.794279, -1.658955, -0.9735625, 
    -1.174687,
  54.59466, 41.54119, 36.90854, 37.00881, 37.66311, 36.54256, 26.87868, 
    3.29043, 6.708549, 11.92383, 13.44654, 1.799009, -0.8448159, -1.66616, 
    -1.597265,
  74.56741, 56.91481, 49.56064, 43.00965, 43.2901, 32.9485, 43.11827, 
    36.91218, 5.484413, 0.5770407, 4.935421, 3.607596, 2.978589, 2.917304, 
    3.166155,
  90.80222, 76.6973, 59.31364, 50.23574, 50.90833, 52.14195, 40.76438, 
    36.55199, 25.30531, 8.33453, 4.522566, 6.017321, 3.504299, 1.967942, 
    1.443788,
  96.09171, 88.43172, 73.59711, 60.69981, 55.12657, 53.49904, 46.72903, 
    40.81102, 27.64492, 2.219496, 0.4371805, -0.3080081, -0.9157287, 
    -0.9954056, 0.02645,
  87.93005, 89.29797, 82.89723, 70.26093, 66.24009, 61.88292, 57.78361, 
    51.12474, 30.14552, 20.37409, 41.73618, 4.638021, -0.572404, -1.508417, 
    -1.910929,
  70.74546, 77.08968, 77.84695, 64.21171, 59.19159, 47.59967, 26.08377, 
    12.56047, 14.8853, 10.61998, 24.60779, 7.121814, 3.054089, 1.985719, 
    0.9971849,
  9.324906, 16.69868, 13.96491, 18.25063, 2.554796, 7.021338, 13.65743, 
    4.146435, 0.666465, -0.1922874, 2.558734, 4.268527, 1.931365, 1.03482, 
    0.4309795,
  27.9847, 22.50804, 13.02631, 7.807407, -0.5744366, 19.58294, 29.89682, 
    8.427144, 1.569432, 0.3690257, 6.816765, 10.23121, 4.520355, -1.478583, 
    -0.5634794,
  50.08276, 39.31733, 36.52443, 10.5202, 1.875208, 1.754473, 40.14448, 
    20.86116, 7.937434, 1.966771, 8.588349, 7.148789, 2.999469, 2.745234, 
    0.9317961,
  50.65396, 47.67327, 50.34447, 51.17544, 23.10808, 3.730291, -0.1435679, 
    26.49561, 19.16544, 3.591655, 6.266503, 7.332445, 4.088881, 3.869726, 
    1.895801,
  51.45573, 39.89571, 38.78256, 41.43379, 43.51101, 30.07928, 17.55989, 
    3.952733, 10.6856, 8.255809, 14.0484, 5.624501, 2.744027, 1.535325, 
    1.58158,
  64.03122, 49.73091, 40.56884, 35.82761, 36.48739, 39.37555, 44.66961, 
    28.41446, 3.072989, -0.5219243, 0.5885051, -0.7488438, -1.293101, 
    -0.2444824, 0.5021273,
  80.51273, 67.6141, 53.40797, 48.50321, 48.08891, 46.84576, 48.0011, 
    45.57572, 27.60418, 5.552867, 1.549825, 0.7469596, 0.8511103, -0.2434367, 
    -1.117394,
  103.3358, 91.40045, 78.73042, 75.26903, 75.06483, 74.74384, 64.58522, 
    58.82447, 32.13204, 4.540134, 1.59696, 1.30769, 0.7852826, 0.1789705, 
    -0.3937433,
  119.3757, 111.757, 102.4609, 94.42988, 89.09182, 79.57234, 71.73164, 
    53.74294, 25.49446, 15.4818, 25.44591, 1.990078, 0.3691415, 0.1209832, 
    0.0864189,
  103.3761, 100.6836, 97.04888, 82.71478, 69.85825, 51.04074, 27.31229, 
    17.91287, 17.44399, 9.443393, 14.98931, 0.8871168, 0.7284331, 0.6647623, 
    1.410578,
  9.636248, 18.53181, 17.8991, 18.41269, 2.594181, 2.961803, 12.41312, 
    2.187389, 0.1507019, -0.924073, 1.30465, 4.661441, 0.813588, -0.6463923, 
    -1.070585,
  21.51109, 18.40498, 13.91358, 7.288987, 4.452792, 25.26661, 29.81849, 
    5.436512, -0.6340856, -1.150665, 3.617606, 9.327283, 5.141623, -1.077569, 
    -0.351234,
  49.65343, 37.99233, 34.35171, 10.2187, 4.844835, 3.965756, 37.15806, 
    16.57026, 4.826535, -0.998875, 6.811653, 5.403562, 0.9898329, 2.039024, 
    0.6420643,
  54.57508, 48.39342, 47.95551, 37.6662, 23.13886, 9.837066, 3.559628, 
    22.81029, 11.83185, 1.345773, 3.304636, 2.645577, -0.08900806, 2.066498, 
    2.10437,
  65.90444, 58.81204, 57.28429, 56.86474, 36.14133, 29.69939, 18.81632, 
    3.902354, 7.702297, 7.125417, 14.61763, 7.792048, 1.524594, 0.9575947, 
    0.246574,
  77.91571, 74.75957, 70.1835, 70.80016, 77.02394, 51.37048, 36.07191, 
    23.85742, 3.759778, 1.449831, 2.980891, 2.360238, 1.555035, 0.4058156, 
    -0.7616412,
  81.25413, 82.06901, 73.17374, 73.63916, 83.69462, 92.18371, 84.09587, 
    55.91685, 23.42458, 4.133821, 1.923625, 0.4650187, 0.42904, -0.9166317, 
    -0.480867,
  82.7374, 73.09833, 61.98402, 62.68536, 68.73109, 78.54485, 76.56322, 
    74.28017, 31.29856, 8.672359, 1.719594, 1.053408, 1.064021, -0.2022473, 
    -0.9776288,
  87.29636, 70.22615, 60.01299, 56.52241, 58.66514, 57.60682, 52.40772, 
    36.06271, 18.96962, 14.36251, 16.09633, 2.265358, 0.1053375, 0.06190119, 
    0.07955436,
  92.00948, 70.17563, 60.08638, 44.70596, 38.26158, 29.69507, 17.95294, 
    13.97866, 12.60489, 7.763633, 8.167176, 0.7049639, 0.9859377, 0.5439801, 
    1.330531,
  9.532152, 15.07024, 10.17675, 14.09601, -1.466819, 3.016914, 10.19523, 
    1.000336, 0.7237169, -0.8104279, 1.421367, 3.575162, -0.006445527, 
    -0.5851552, -0.922075,
  32.29867, 22.71077, 7.98823, 4.667947, -1.391326, 16.49268, 20.73861, 
    2.364363, -0.04056245, 0.623805, 4.56824, 9.345811, 4.955382, -0.6983109, 
    -0.6778686,
  57.09753, 52.84748, 34.59722, 3.547364, 2.375182, 2.777515, 27.00433, 
    8.734971, 1.227926, -0.5066484, 11.03157, 8.698533, 1.506434, 1.772234, 
    0.2450126,
  50.75285, 56.55313, 47.77981, 35.20155, 16.08528, 3.439861, 0.9009537, 
    12.76919, 7.25918, 0.6244166, 3.671712, 4.822048, 2.155133, 2.450563, 
    3.334762,
  74.57838, 70.32983, 55.79291, 46.83341, 36.07377, 19.45507, 8.349995, 
    0.4790759, 5.121462, 4.929121, 10.85987, 3.953933, 3.07485, 3.300693, 
    2.635084,
  112.6278, 97.93974, 70.9129, 48.26275, 53.52996, 47.91853, 37.86052, 
    18.16743, 2.805291, 1.741678, 4.164302, 4.869164, 1.177387, 1.182161, 
    1.311607,
  136.8904, 112.3687, 76.60861, 47.47672, 51.96491, 70.8413, 81.6526, 
    66.77481, 25.67349, 8.96559, 5.909829, 1.689631, 1.47276, 0.4335572, 
    1.262715,
  135.598, 102.187, 59.79013, 54.45629, 57.41259, 65.62025, 63.59294, 
    51.82744, 16.50178, 6.667192, 3.505495, 3.144705, 3.014321, 0.5775229, 
    0.9144019,
  146.5731, 123.1042, 97.23866, 74.51564, 61.48671, 47.87324, 42.43169, 
    26.8125, 12.80769, 11.57434, 12.33461, 3.750223, 0.9901108, 0.7279097, 
    0.2506637,
  161.111, 131.0173, 112.7525, 79.2656, 59.40571, 33.23883, 18.69444, 
    11.43204, 7.779245, 6.483746, 6.177783, 1.014662, 0.4925878, 0.2088311, 
    1.002726,
  9.919583, 17.30066, 13.33459, 13.46007, 2.021158, 6.802731, 15.07888, 
    0.1479663, 2.973409, 1.73219, 3.186131, 5.873537, 2.262995, 0.6032555, 
    -0.3786741,
  24.7067, 13.68934, 6.596042, 3.371925, -0.5432887, 19.86605, 23.23781, 
    3.361459, 1.969206, 4.285196, 7.62679, 11.62411, 7.950454, 0.9147947, 
    -0.2572634,
  52.51332, 46.78766, 30.74556, 5.9697, 3.520129, 0.7515644, 25.26168, 
    12.10259, 2.339298, 0.03238342, 14.84769, 11.22279, 4.573127, 4.009881, 
    1.437504,
  56.53345, 62.41013, 69.09586, 56.95918, 26.83195, 6.569636, -0.6496505, 
    9.960818, 6.519596, 2.170712, 2.61076, 2.729575, 2.843359, 3.107018, 
    3.641677,
  68.08393, 73.92796, 75.47882, 69.65369, 61.86928, 37.134, 8.600003, 
    -0.05769422, 2.204556, 1.938686, 4.506897, 0.6559052, 0.2765961, 
    2.994403, 2.678076,
  118.9202, 105.9989, 88.89292, 69.44013, 52.24389, 45.43345, 47.53197, 
    18.27439, 2.168753, 1.065404, 0.4851954, 1.299094, -0.8249782, -1.667298, 
    -1.443798,
  147.0782, 128.5827, 102.7159, 73.27668, 55.07247, 50.03984, 54.90751, 
    50.07997, 13.63427, 5.466974, 1.850582, -0.6116993, -0.7319043, 
    -1.462537, -2.096854,
  173.2031, 148.1383, 122.6028, 99.81889, 92.83425, 90.36578, 79.34074, 
    68.27064, 20.41072, 6.043579, 2.552256, 1.535738, 0.4711268, -0.382011, 
    -1.052914,
  203.5812, 175.6058, 155.0753, 126.31, 103.1597, 79.64197, 50.98777, 
    37.31024, 19.60047, 11.44101, 5.159283, 1.655578, 0.8168426, 0.1090562, 
    -0.3112368,
  179.1599, 152.1294, 130.8291, 75.67622, 47.0814, 28.08339, 22.19984, 
    20.5327, 11.40032, 6.42815, 2.575958, 0.6490391, 0.3062659, 0.2124477, 
    0.2630271,
  3.043342, 8.365808, 5.369421, 9.215887, 1.966169, 5.611006, 11.43017, 
    4.556148, 4.304733, 1.715453, 1.145565, 2.67446, 0.3744179, -0.1641784, 
    -0.3257529,
  17.54303, 7.558211, 5.650983, 4.139949, -0.004418987, 9.244152, 12.23877, 
    4.201063, 3.849452, 4.863791, 4.308456, 7.194433, 3.962681, -0.2330336, 
    -0.4167754,
  50.90778, 38.47618, 17.40399, 3.772252, 3.804351, 1.491036, 10.87245, 
    6.746195, 4.619035, 6.398775, 14.11361, 8.660316, 0.6244587, 1.351249, 
    0.1347473,
  38.13242, 37.74413, 51.46238, 38.57705, 15.71435, 4.829234, -0.3523106, 
    6.344265, 6.979866, 5.856353, 6.800614, 6.469513, 0.93029, 0.8285818, 
    1.844436,
  80.40564, 76.0312, 68.30048, 60.88083, 47.34915, 24.37303, 8.356426, 
    0.222752, 1.713577, 3.350927, 4.852377, 3.40659, 1.425452, 1.403393, 
    1.331456,
  125.7306, 108.1225, 94.80416, 81.04377, 72.10369, 57.38212, 39.74213, 
    19.89432, 7.552169, 6.879227, 4.095043, 2.802652, 2.094643, 1.052696, 
    0.1091699,
  143.397, 131.5803, 113.9259, 100.4089, 93.43165, 81.93346, 61.1445, 
    35.74632, 11.61308, 9.740399, 4.916357, 1.017124, 0.008159536, 0.8099894, 
    0.8727504,
  156.709, 147.9612, 131.81, 121.6289, 112.4514, 105.3272, 79.9861, 62.3393, 
    13.18185, 1.543528, 3.235308, 1.842857, -0.07243426, -0.3327206, 0.1456727,
  150.1356, 142.3047, 135.2259, 118.7727, 84.22401, 60.89654, 50.22097, 
    33.9062, 11.11467, 3.16426, 4.912498, 2.115764, -0.3344897, -0.8898684, 
    -0.7113947,
  125.951, 116.6237, 105.5057, 57.44862, 31.01858, 16.82476, 14.81504, 
    19.35372, 9.990909, 1.6057, 2.145909, 0.4759702, -0.1684238, -0.05160339, 
    1.022957,
  3.703366, 5.328925, 2.409638, 5.203924, 3.516695, 6.945303, 10.52868, 
    2.919256, 1.092333, 3.061877, 2.841709, 5.492331, 3.245187, 2.272308, 
    1.115501,
  20.0192, 13.02908, 2.694352, -0.2348914, 1.077765, 10.69617, 9.990748, 
    4.132512, 1.939239, 4.15437, 6.028474, 14.4713, 12.5657, -0.701148, 
    -0.2512487,
  40.53384, 40.49393, 22.05552, 1.244189, -0.07679018, -0.8206546, 9.389323, 
    6.139486, 4.717746, 4.205225, 13.26749, 8.180907, 4.643218, 6.03524, 
    1.733894,
  50.30874, 33.35743, 41.96211, 43.28929, 11.14722, 3.954144, -0.5897752, 
    3.793497, 3.745774, 2.17082, 2.821061, 4.318365, 2.319355, 3.622356, 
    3.664846,
  119.4392, 95.3829, 65.39652, 33.85017, 43.61244, 25.07795, 9.049622, 
    1.005051, 0.8478833, -0.1652538, 2.64957, 1.710611, 1.073408, 1.686107, 
    1.306363,
  133.7411, 130.9825, 121.6312, 89.47735, 60.07737, 46.35794, 37.62235, 
    15.39829, 6.866483, 6.932343, 4.723991, 4.127508, 2.260173, 0.5512128, 
    0.2708068,
  129.875, 130.7195, 130.8659, 126.2543, 120.4123, 96.29472, 59.5789, 
    35.27776, 12.69217, 13.12875, 7.091452, 1.964399, 1.148754, -0.09505803, 
    0.2529273,
  126.2949, 120.6446, 116.8556, 117.1977, 122.7118, 120.6154, 90.62038, 
    55.10666, 10.41197, 2.326861, 1.847398, 2.208391, 2.110735, 0.3502366, 
    0.2155268,
  122.3575, 119.4451, 121.6735, 113.8707, 76.31185, 61.00161, 50.04784, 
    29.99663, 11.46244, 3.637101, 1.695829, 2.365681, 1.06745, 1.664598, 
    0.6937389,
  117.2753, 103.5383, 97.72542, 52.43141, 24.28182, 13.8316, 12.37644, 
    18.36254, 10.92406, 0.8243782, 0.6450568, 1.536807, 2.16355, 2.038485, 
    2.132248,
  5.404662, 5.548995, 3.48376, 4.579548, 2.449775, 4.55773, 10.63186, 
    6.497167, 8.299306, 2.032952, 0.2111214, 8.194454, 5.147171, 3.70605, 
    1.61638,
  15.37467, 4.978432, 3.500475, 1.197817, 0.8857738, 8.226168, 12.17997, 
    6.550169, 2.867821, 10.00323, 4.864781, 13.55169, 14.97183, 1.108641, 
    0.0625532,
  71.00584, 24.69325, 13.41101, 1.072333, 3.071448, 0.1189457, 9.238224, 
    8.41756, 4.390395, 7.350257, 13.64221, 7.055607, 4.363616, 9.204147, 
    4.212916,
  125.3304, 68.39661, 41.69936, 42.84666, 8.470553, 5.404868, -0.3771086, 
    4.43244, 4.89044, 3.0748, 4.135899, 4.909578, 2.24617, 5.130326, 8.702857,
  138.0486, 124.1039, 61.27312, 43.60243, 55.47449, 19.68179, 12.21521, 
    -1.646871, -1.164386, 0.7872146, 3.490983, 3.789318, 2.544544, 3.844365, 
    6.536257,
  120.3097, 132.8836, 121.6302, 60.59538, 55.89475, 65.39383, 43.72617, 
    19.4368, 11.33265, 12.25248, 10.52455, 8.709432, 4.435757, 0.7043632, 
    0.639948,
  120.4004, 127.0722, 136.3846, 109.3294, 70.86607, 64.02545, 54.99581, 
    45.26957, 18.48922, 18.65232, 13.46588, 6.391707, 1.803993, 0.9900978, 
    1.588242,
  126.3867, 123.0048, 126.7984, 122.0542, 105.6477, 80.1215, 54.47491, 
    32.6825, 9.806539, 3.821202, 1.111728, 5.182357, 2.857636, 0.2141911, 
    1.534527,
  146.8946, 135.0059, 131.907, 118.6689, 68.66545, 48.27018, 32.4186, 
    15.55002, 3.88831, 0.8870779, -0.4581871, 3.042228, 2.160665, 0.6764488, 
    1.609753,
  133.8706, 120.3392, 103.957, 50.53819, 19.19444, 11.57842, 9.344169, 
    13.72622, 4.995981, -1.097878, -0.7836344, 2.981674, 2.463599, 3.92635, 
    4.051002,
  3.061623, 9.935167, 3.182284, 8.601567, 6.007753, 4.955175, 15.09131, 
    8.362559, 9.421849, 2.450495, 0.9297222, 3.726008, -0.7765248, -2.501439, 
    -3.580653,
  32.34975, 8.585974, 5.917196, 4.335653, 1.687588, 5.683316, 8.645703, 
    4.663864, 1.762085, 11.05885, 2.186305, 10.32763, 11.07622, -2.637249, 
    -3.309569,
  115.3409, 58.21879, 17.58278, 4.596961, 3.868526, 0.3529231, 6.256145, 
    4.09295, 1.996274, 7.655152, 10.63347, 2.201042, 1.757927, 8.052748, 
    1.832955,
  133.1365, 114.108, 80.22078, 48.4216, 12.92784, 9.483373, -1.017406, 
    0.1537119, 2.152223, 0.9898846, 0.1820195, -0.05799042, -0.6312618, 
    3.685024, 9.085467,
  136.9311, 115.3339, 93.33306, 71.13115, 56.38411, 24.7161, 17.75023, 
    -1.685235, -1.481161, -1.312224, -1.598098, -0.556206, -0.06713495, 
    3.253809, 7.969224,
  144.8104, 131.5429, 110.8139, 81.15955, 72.75014, 69.00186, 38.98925, 
    20.18613, 14.19769, 16.12295, 5.927698, 2.41379, 1.645448, -0.04448749, 
    -0.1920199,
  152.2795, 151.5925, 127.71, 99.46967, 82.73849, 77.40237, 71.90533, 
    46.79424, 23.50245, 28.55996, 15.57052, 4.829176, 2.825353, 0.851712, 
    -0.7309126,
  161.8659, 159.3571, 138.894, 115.6721, 96.04369, 77.58031, 67.60442, 
    51.06643, 13.2613, 6.335359, 4.27108, 4.83948, 4.602006, 0.9942273, 
    -0.1390413,
  168.4556, 165.7915, 156.2322, 117.0866, 53.92212, 43.05979, 35.72849, 
    21.42727, 8.254116, 3.462464, 3.241389, 5.26355, 2.281567, 0.5472095, 
    1.277106,
  138.9886, 128.0429, 112.0602, 49.29536, 18.8522, 12.57961, 12.70736, 
    22.94083, 9.206445, 2.536146, 4.685773, 3.822316, 3.40547, 0.7706236, 
    2.715749,
  2.988695, 10.68878, 4.812542, 6.796207, 2.280535, 5.098886, 16.68489, 
    8.260121, 10.27993, 4.400008, 5.09793, 7.662319, 2.211668, -0.09167443, 
    -1.926595,
  37.46715, 13.90726, 7.546229, 5.844191, 1.429928, 3.145568, 13.70928, 
    9.739537, 5.340526, 13.55306, 5.888784, 13.04649, 13.52344, 0.4975284, 
    -0.9580925,
  88.60468, 48.38886, 19.96867, 6.03303, 3.545408, -1.249829, 7.379891, 
    6.943944, 6.046851, 11.14251, 9.492773, 6.377231, 6.187712, 8.322006, 
    2.338556,
  112.5458, 95.98917, 86.3651, 61.1755, 15.44929, 15.90929, -0.5142096, 
    2.197108, 4.318505, 2.131122, 2.398215, 2.325512, 2.530718, 8.058232, 
    9.427196,
  128.1574, 105.4604, 97.60448, 98.17224, 70.93217, 36.48241, 33.04419, 
    -1.50028, -1.278496, -1.270542, 0.2614288, 1.802472, 3.602487, 5.525944, 
    9.650279,
  144.7057, 122.4088, 108.2948, 100.9612, 109.0533, 94.14673, 41.19624, 
    22.74452, 15.41737, 15.12023, 5.861205, 4.854538, 4.353373, 2.635706, 
    2.20961,
  158.7811, 140.6536, 119.0758, 104.409, 109.1863, 109.3083, 92.82559, 
    45.05149, 20.67967, 28.96074, 15.5394, 4.929102, 2.452058, 0.2838337, 
    -0.3332829,
  170.078, 147.98, 123.8432, 105.5147, 102.7632, 94.57954, 83.68662, 
    54.83899, 6.588829, 2.68788, 2.909161, 1.33106, 0.01399682, -0.3491144, 
    -0.01370925,
  166.5055, 149.9943, 133.5864, 88.99371, 48.89985, 45.23363, 37.0808, 
    15.12213, 3.046529, -0.5109892, -0.9228903, 0.3754868, 1.293017, 
    0.7489223, 2.526384,
  127.6838, 106.2238, 83.8574, 30.72374, 6.731597, 3.061593, 4.394678, 
    15.48422, 3.902503, -0.09801307, -0.570269, 0.4017186, 2.465174, 
    0.3002842, 3.156206,
  0.7899338, 4.575413, 1.780321, 5.360276, 1.025493, 3.587324, 7.667677, 
    5.006925, 6.74924, 1.292111, 0.7698832, 7.357461, 3.953676, 2.383729, 
    -0.4447821,
  38.23088, 9.719289, 3.309002, 2.5491, 1.13868, 3.488976, 7.348588, 
    2.782895, 0.8213834, 6.603689, 2.220237, 12.19481, 17.03778, 2.558912, 
    -0.6425495,
  108.0762, 64.33129, 26.8918, 11.13461, 15.45371, 0.1665143, 2.096756, 
    -0.08141546, -0.158044, 6.523411, 8.539541, 7.653617, 11.93951, 14.39084, 
    4.4688,
  138.1736, 130.3413, 118.7677, 69.25672, 26.63862, 24.5829, -0.8386088, 
    -2.161829, -0.3704646, 0.2515953, 2.192067, 3.490644, 4.836611, 9.658442, 
    10.59946,
  133.9267, 119.9264, 115.9913, 108.0926, 53.9598, 31.53693, 28.33328, 
    0.2080507, -0.1494615, 0.8308439, 0.8337133, 1.921846, 1.52099, 7.626162, 
    11.28213,
  120.7359, 111.4906, 102.274, 93.83176, 90.09401, 61.95076, 24.65998, 
    19.47858, 13.57546, 19.35438, 5.971211, 4.189891, 2.696282, 2.84146, 
    1.403776,
  106.4425, 102.5116, 91.75366, 81.12626, 83.55528, 80.82541, 65.38277, 
    29.15407, 21.4608, 25.80549, 10.48247, 4.477657, 3.262295, 2.038724, 
    0.2330539,
  100.4746, 98.03016, 87.24811, 77.2887, 77.79671, 70.28101, 62.41821, 
    41.50972, 10.89768, 5.37367, 2.688962, 2.328418, 0.8185675, 0.8990702, 
    -0.103413,
  89.6946, 91.30871, 89.60931, 67.12952, 40.25208, 34.95858, 30.44538, 
    10.47873, 2.356475, 0.3722575, -0.03275099, -0.05601056, -0.07182936, 
    -0.06304086, 1.509454,
  61.32689, 57.39396, 52.57165, 20.24905, 9.354373, 4.387329, 5.3309, 
    6.569396, 1.205815, 0.3604477, 0.08012602, 0.0727319, 0.3872516, 
    0.1607266, 2.395898,
  5.673601, 11.63837, 5.664033, 5.573139, 3.822894, 2.787962, 7.303291, 
    7.701485, 11.80382, 6.082405, 2.69853, 5.997936, 1.970697, -0.1624503, 
    -2.681576,
  38.48741, 17.37552, 10.62248, 7.681941, 3.693772, 0.11239, 2.303665, 
    3.239144, 7.409675, 15.70318, 5.586512, 12.26287, 10.76519, -0.234419, 
    -2.169636,
  77.47474, 45.52302, 20.75062, 9.451737, 11.06845, -1.183607, 1.727966, 
    3.84601, 4.444406, 8.408164, 9.418921, 7.104014, 9.337223, 8.116943, 
    2.604858,
  94.35476, 88.63383, 80.42104, 43.06142, 16.93812, 14.70293, 0.7821622, 
    -0.7375525, -0.03014299, 2.701111, 5.13627, 5.328602, 6.038811, 5.884924, 
    6.46787,
  92.60941, 82.7131, 80.08508, 72.59095, 33.41475, 24.08871, 22.41379, 
    1.334594, -0.0444024, 1.004017, 3.27095, 1.794034, 4.048741, 3.749029, 
    5.200914,
  69.48475, 65.59474, 61.87865, 58.13654, 58.67712, 45.90973, 18.86834, 
    22.47316, 11.31627, 14.42587, 1.461923, 2.964928, 2.088866, 2.022695, 
    0.8196942,
  50.45742, 50.1705, 44.23718, 41.48241, 51.10054, 57.35799, 51.75927, 
    25.53228, 17.36204, 15.39815, 3.836805, 2.624846, 1.30087, 0.6709396, 
    0.4697837,
  48.55468, 49.06136, 43.15909, 40.67619, 48.96564, 49.32332, 43.54312, 
    27.32493, 5.916618, 3.714964, 1.599302, 1.960805, 1.889458, 1.398737, 
    0.3001082,
  55.53613, 59.86457, 56.08726, 42.69505, 24.66681, 20.08923, 18.05309, 
    6.001796, 2.751878, 2.335023, 0.8628984, 0.04528611, 0.9368213, 
    0.6135628, 2.667342,
  44.83483, 39.60159, 32.79221, 9.988139, 4.614219, 2.069551, 2.172424, 
    2.129323, 1.701478, 1.378016, 0.1449208, 0.07738672, 0.4564783, 
    0.3463978, 2.882521,
  3.807262, 10.65962, 6.088942, 9.247755, 8.424295, 4.150636, 6.576757, 
    5.122167, 12.20291, 6.662595, 3.037291, 5.810923, 4.128937, 0.6036286, 
    -1.600672,
  15.91818, 7.365229, 7.17765, 6.170622, 3.915471, 0.2004982, 6.294865, 
    4.912925, 8.752883, 14.45077, 2.677036, 10.91493, 18.72832, -2.355054, 
    -3.429125,
  47.72126, 22.38335, 10.94606, 5.620122, 6.231019, -0.7638651, 4.423758, 
    4.910983, 5.703192, 9.159429, 5.191825, 8.835026, 16.13761, 13.89504, 
    1.649734,
  59.8266, 51.5264, 45.08557, 28.85809, 13.00891, 14.49243, 0.7770862, 
    1.578783, 9.688672, 6.999934, 5.620124, 5.908081, 9.612594, 8.01161, 
    7.551116,
  70.09881, 53.83348, 44.58155, 41.46489, 22.83873, 25.42594, 22.72285, 
    -0.5970554, 4.955249, 7.493343, 4.02878, 1.886892, 4.392962, 4.381302, 
    9.17795,
  87.26139, 71.92995, 58.87762, 45.70492, 38.35206, 38.37043, 20.47924, 
    20.98756, 14.01325, 12.25667, 2.629669, 2.12003, 0.6345705, -0.4071553, 
    0.8689408,
  88.14307, 77.65264, 65.81824, 50.17055, 41.18291, 36.61623, 52.41901, 
    29.28051, 19.69386, 10.65981, 4.290544, 2.090034, -0.2635911, -1.335444, 
    -1.84508,
  74.47139, 61.19081, 49.08209, 40.09215, 42.75396, 41.92321, 41.56329, 
    28.39035, 10.86794, 8.486175, 5.037026, 2.633173, 0.8711451, -0.2336554, 
    -0.8818481,
  66.9439, 50.50374, 44.43298, 36.81223, 23.12269, 18.45275, 16.18618, 
    5.99614, 5.859745, 7.246586, 4.458266, 1.662878, 1.379327, -0.2693075, 
    2.107361,
  53.4633, 37.71749, 33.76222, 6.370066, 2.90202, 1.002344, 1.311635, 
    2.582903, 2.598416, 2.623667, 0.3239742, 0.7589166, 0.5902497, 
    -0.3580109, 1.490278,
  5.970777, 12.04284, 9.969385, 8.883695, 8.090846, 1.760396, 4.24878, 
    1.55993, 4.548876, 1.349956, 1.452004, 2.979613, 0.2985502, -1.268135, 
    -0.113153,
  29.40181, 11.96063, 8.90564, 7.589459, 3.243542, -0.1222754, 3.627908, 
    2.752867, 4.288167, 7.647427, 5.618585, 8.054809, 8.180506, -0.8063442, 
    -0.4872782,
  80.99802, 36.5196, 13.85992, 4.031024, 5.341089, -1.11948, 3.168245, 
    3.679539, 3.535969, 8.298427, 9.973845, 7.579525, 5.886652, 8.909203, 
    6.487288,
  86.5119, 78.79455, 74.15643, 43.35979, 10.4289, 5.082088, -0.3415588, 
    3.29023, 5.778468, 3.742826, 9.726416, 7.090722, 4.539525, 3.537922, 
    12.02358,
  83.78008, 57.22052, 62.35383, 57.60373, 18.07155, 13.50328, 14.2921, 
    0.1776404, 2.19602, 1.455992, 2.105608, 1.961362, 2.338878, 2.538415, 
    9.701479,
  83.56735, 58.39245, 62.93098, 60.12107, 52.81957, 42.1082, 16.01365, 
    12.65804, 7.631045, 5.894701, 1.084252, 0.5687811, -0.1582994, 4.464565, 
    5.143251,
  93.81342, 77.49091, 75.93842, 65.90534, 75.50696, 80.09862, 68.09823, 
    27.04657, 10.45184, 4.573747, 2.349161, -0.3277874, -0.2066951, 3.759228, 
    4.299592,
  102.9003, 88.0678, 83.36039, 85.03275, 102.7213, 97.94154, 80.05118, 
    30.77123, 8.126666, 2.257672, -0.4272868, -1.439368, 2.686309, 3.568018, 
    2.095468,
  105.5293, 95.5341, 105.2243, 94.94392, 58.51999, 48.03277, 34.73695, 
    11.92268, 6.457448, 1.477303, -0.4142101, 0.6201785, 2.082223, 3.032688, 
    4.289776,
  94.96902, 89.17733, 90.43118, 22.2816, 11.32724, 7.387245, 6.709749, 
    11.56002, 4.963806, 0.8278776, -1.019371, -0.2752171, 0.9143337, 
    1.012303, 1.923231,
  10.8473, 18.16075, 16.59517, 10.46447, 3.204747, 4.739457, 8.835649, 
    2.442744, 2.887864, 0.6173652, 1.053265, 3.324991, 1.062063, 0.8838992, 
    -0.7328515,
  21.29783, 15.93943, 16.44745, 8.000452, 2.989288, 6.943119, 8.307812, 
    2.762227, 3.068642, 5.11371, 3.577806, 6.110896, 7.106818, -0.3100891, 
    -1.032779,
  54.82008, 35.23146, 27.30505, 12.47789, 8.971059, 2.482983, 8.068266, 
    3.397163, 1.320232, 5.432103, 3.98285, 1.654284, 4.170973, 7.739233, 
    2.805328,
  55.71623, 71.17043, 87.46861, 64.81257, 15.3501, 8.065226, -0.06081075, 
    0.5850395, 1.381314, 1.256742, 1.282837, 1.424591, 3.295589, 5.167778, 
    5.247733,
  50.95375, 47.22168, 60.9451, 67.82958, 31.9623, 15.90691, 14.30326, 
    1.654236, 0.9137887, -0.02624129, -0.4257951, 0.6080714, 2.593694, 
    4.269022, 5.625473,
  99.0628, 86.59691, 82.52103, 79.42303, 69.30188, 40.58114, 13.96982, 
    19.29168, 10.01495, 8.228806, 0.9657458, 0.9109624, 1.761126, 3.407151, 
    3.826215,
  141.8063, 129.9046, 111.7458, 94.77632, 94.68422, 94.54005, 67.88239, 
    21.79366, 7.441621, 4.155895, 4.35167, 2.19973, 1.990655, 0.6810285, 
    0.2449064,
  173.7704, 164.7486, 145.819, 126.6018, 127.4205, 117.6832, 87.8119, 
    29.09389, 5.507992, 2.444004, 1.671912, 1.497142, 0.271037, 0.08805656, 
    -0.00937655,
  196.6922, 189.5668, 174.1656, 125.065, 81.12553, 62.63584, 37.53814, 
    12.89812, 2.476467, 1.373136, 0.3917704, 1.146111, 0.8633564, 0.8570692, 
    2.186048,
  167.6246, 154.3451, 118.1628, 25.85355, 14.3624, 6.27533, 5.45688, 
    14.38298, 3.3496, 2.276276, 0.3936279, 0.8438295, 1.234116, 0.4296832, 
    1.894847,
  6.717868, 14.90379, 17.14935, 13.941, 1.994292, 4.404149, 7.665853, 
    1.166133, 1.295968, -0.1485356, 0.5828787, 1.494596, 0.2919521, 
    0.8382845, -0.004525182,
  15.7201, 15.94295, 16.23755, 9.69235, 3.009358, 7.261256, 5.398427, 
    1.065801, 0.5411004, 1.451902, 1.002917, 3.737195, 4.133713, -0.1292174, 
    -0.1905923,
  45.57643, 30.42903, 20.37746, 11.90903, 11.49738, -0.395142, 1.686651, 
    0.3560112, 0.1053782, 1.873847, 2.677229, 2.576149, 4.858668, 8.568286, 
    2.793417,
  56.73268, 69.4944, 85.09476, 62.25507, 22.78151, 17.29721, -1.40381, 
    -0.06827955, 0.5209522, -0.05564907, 0.8634862, 0.9394608, 3.965825, 
    5.446682, 3.83549,
  97.27412, 90.56219, 104.0787, 107.5739, 35.63, 18.52357, 18.25853, 
    -0.2944423, 0.1548417, 0.2628221, 0.468281, 0.5465664, 3.446313, 
    4.586314, 4.689394,
  137.5724, 128.2232, 119.4812, 111.1593, 85.62065, 41.68147, 8.847628, 
    10.93466, 4.230277, 4.358967, 0.8688876, 1.248802, 2.677544, 3.275026, 
    4.016756,
  151.036, 145.9497, 125.9809, 104.9364, 99.03716, 82.59054, 39.32248, 
    11.01635, 4.372634, 3.721895, 1.929913, 1.419456, 1.276283, 0.8721017, 
    1.543148,
  153.2684, 145.1635, 124.6664, 104.5877, 99.86815, 85.78118, 58.66644, 
    18.11948, 5.11406, 2.13169, 0.4457825, 0.4439321, 0.1632933, 0.07973691, 
    1.35773,
  160.6536, 150.8909, 131.5316, 97.21337, 70.25398, 51.61681, 25.20997, 
    8.094605, 2.392662, 0.843794, 0.06382936, -0.1905777, -0.2162997, 
    0.2735058, 1.737774,
  133.0045, 119.6874, 81.69778, 15.82498, 6.351663, 5.499237, 2.951801, 
    6.4422, 1.911971, 0.4387189, -0.1613601, -0.2964325, -0.2403323, 
    -0.04749517, 0.777725,
  3.656258, 7.167528, 7.540684, 6.446011, 1.642161, 3.612134, 7.435907, 
    3.122318, 3.38802, 0.02068568, 0.09810527, 0.6005309, -0.09561584, 
    -0.07191042, -0.7605262,
  9.288404, 7.027572, 6.80075, 4.344369, 2.072933, 2.838658, 3.727733, 
    1.913186, 0.2935774, 1.429502, 0.6956308, 1.771896, 1.140498, -0.8472306, 
    -1.066647,
  47.14822, 24.84071, 13.25029, 9.203364, 12.95606, -2.453154, 2.50193, 
    1.348795, -0.2246843, 1.124301, 1.444334, 0.8036211, 2.283727, 4.171575, 
    1.090504,
  62.57385, 73.37763, 72.2149, 44.55949, 21.87885, 18.81751, -1.351005, 
    -0.4842702, 0.3821291, 0.3600661, 0.8547824, 1.645294, 3.36919, 5.996624, 
    3.942664,
  86.64374, 79.28466, 90.00928, 91.0856, 24.9072, 16.67237, 20.10452, 
    -0.3761629, 0.3669469, 0.4834587, 0.9901174, 0.8748327, 4.101905, 
    4.184525, 5.247979,
  109.7096, 98.999, 96.70618, 92.29388, 62.55156, 28.13688, 8.667454, 
    10.54852, 2.642658, 1.400823, 0.7575825, 0.884762, 2.68405, 3.637408, 
    3.587086,
  126.9679, 119.5393, 104.5848, 89.07006, 81.88863, 65.84589, 26.13843, 
    2.886411, 1.456634, 1.286935, 1.188196, 1.136019, 1.351161, 0.9505464, 
    1.936031,
  131.7411, 119.748, 97.63679, 81.40974, 77.37193, 65.70816, 45.67576, 
    13.90806, 2.560983, 1.198634, 0.5230988, 0.3552896, 0.1789786, 0.1609935, 
    1.828872,
  131.3989, 117.7366, 98.90179, 73.7401, 55.97231, 39.2348, 19.11161, 
    4.267552, 1.884445, 0.7582474, 0.1009862, 0.02927023, -0.08787226, 
    0.3520556, 1.618823,
  107.5871, 94.96961, 58.3739, 8.617567, 2.826733, 2.324134, 3.193919, 
    2.216947, 1.066565, 0.2896398, 0.09608596, -0.1108482, -0.2029659, 
    0.02361427, 0.6186045,
  5.19751, 8.486818, 4.814653, 2.940401, 0.5431216, 0.3018713, 2.738617, 
    3.486621, 7.241432, 3.48326, 1.129009, 2.709696, 0.4705891, -0.1446217, 
    -0.8162465,
  10.55801, 3.2642, 2.194049, 1.353446, 0.06791573, 0.2297352, 5.253278, 
    5.046925, 6.136176, 8.078125, 1.104558, 2.632577, 2.401822, -0.3592823, 
    -0.4176695,
  31.97244, 15.17405, 5.653316, 2.2239, 8.328739, -0.7099618, 2.230315, 
    2.619374, 2.159065, 3.93473, 2.380321, 0.4067617, 0.9667298, 1.65126, 
    1.572274,
  53.24646, 59.46415, 55.30265, 28.98717, 15.00034, 20.11322, -0.4503989, 
    -0.6714479, -0.2784406, -0.4618838, 0.1025366, 0.5695838, 1.574734, 
    2.995717, 3.04537,
  78.65922, 70.41429, 75.19558, 70.95703, 14.50677, 17.2427, 21.6966, 
    -0.09512186, -0.1235256, 0.3450509, 0.7004942, 0.6768405, 1.831092, 
    2.6988, 4.456103,
  88.00204, 84.00136, 82.79287, 78.66214, 51.31026, 21.94109, 8.438101, 
    12.66038, 3.2736, 2.812805, 0.544319, 0.4020651, 1.187011, 1.929428, 
    3.70929,
  88.92047, 93.62904, 88.1881, 79.784, 81.28005, 69.34258, 26.11041, 4.43259, 
    1.387761, 0.8789319, 0.4081855, 0.2506776, 0.2754418, 0.2538801, 1.076859,
  83.86174, 90.6964, 82.13145, 74.67203, 79.40794, 74.64634, 51.57473, 
    13.2099, 2.817374, 0.8985233, -0.06597362, -0.2152603, -0.3174117, 
    -0.2154959, 1.574007,
  79.37604, 84.79029, 81.25388, 71.72398, 62.9432, 47.5089, 22.63457, 
    6.021813, 2.542269, 0.7049531, -0.1362174, -0.283403, -0.3833803, 
    0.1072144, 2.447974,
  80.21519, 78.61595, 55.27074, 11.44846, 3.528527, 2.752672, 6.921828, 
    3.80952, 0.993763, -0.04957977, -0.3746369, -0.3040196, -0.02427871, 
    0.0263174, 1.09318,
  5.67055, 9.725774, 7.669638, 5.136595, 2.579179, 0.2979728, 2.457583, 
    2.368788, 4.80913, 1.530809, -0.02524396, 1.072637, 1.319449, 0.3467499, 
    -0.4481342,
  14.39752, 5.83843, 6.260094, 4.475141, 1.979375, -0.1946894, 2.631612, 
    2.859612, 5.27788, 9.096496, 0.2910242, 1.653879, 3.426524, 0.1933549, 
    -0.09262436,
  52.0363, 21.5927, 8.741211, 5.180288, 8.092701, -0.8470914, -0.4659574, 
    0.09124587, 0.576705, 3.267192, 2.531073, 0.4695855, 1.4314, 1.90883, 
    1.502699,
  67.14145, 64.9388, 56.43419, 25.40125, 9.227283, 11.43916, 0.2541684, 
    -1.065523, -0.06995848, 0.5073367, 1.686889, 2.303581, 4.479073, 
    4.604462, 2.459281,
  77.92933, 64.82967, 65.71933, 52.29609, 8.873663, 9.297225, 13.30322, 
    0.7865784, -0.7780553, -0.198835, 0.3903871, 0.9232666, 3.475113, 
    4.263199, 5.319134,
  90.11845, 76.10561, 69.75836, 55.43331, 35.52626, 16.11519, 8.671752, 
    12.90069, 5.985867, 4.021914, 0.3338702, 0.574201, 1.66519, 1.918205, 
    4.327782,
  101.5985, 93.17658, 79.86345, 62.96686, 65.33945, 61.5106, 24.24233, 
    8.836763, 5.064083, 3.005413, 1.417763, 0.7030746, 0.3472625, -0.3294203, 
    0.9399443,
  114.1845, 104.2142, 84.27591, 70.32843, 76.27316, 71.62971, 50.23944, 
    12.41875, 4.566344, 1.605396, 0.3840801, 0.1312973, -0.1670596, 0.108404, 
    2.34409,
  121.1992, 108.3613, 97.4715, 82.50688, 69.10529, 48.73384, 18.7709, 
    6.883577, 3.867786, 0.8506292, -0.1220345, -0.2182516, 0.02834091, 
    0.7004718, 4.196331,
  115.8486, 108.2527, 72.02443, 24.8007, 8.179914, 6.056065, 4.423459, 
    6.072254, 1.984586, 0.01090452, -0.5587403, -0.2808461, -0.001063216, 
    0.204336, 1.826964,
  11.54867, 17.37876, 8.063355, 7.860371, 3.999559, 0.3109089, 0.5689675, 
    0.2822036, 3.052584, 0.9097395, -0.1150491, -0.1321779, 0.1177961, 
    0.7095652, 0.1228292,
  21.1428, 12.34083, 9.747813, 6.026583, 2.644008, -0.6791436, -0.1852928, 
    0.03401369, 1.883022, 4.316, -0.1882009, 0.4122207, 2.102487, 0.1905383, 
    -0.1160363,
  71.3574, 25.35953, 7.462311, 4.770664, 4.795106, 0.1118171, -0.1075549, 
    -0.07416849, 0.646031, 2.158161, 1.5458, 1.259321, 3.272127, 3.578202, 
    1.541879,
  84.11239, 72.84257, 49.10973, 18.35873, 6.259519, 6.961913, 0.8495733, 
    -0.1540351, 0.1256157, 0.3361664, 1.033255, 1.365934, 4.148954, 4.606797, 
    2.681902,
  82.7017, 61.35749, 55.96498, 43.39519, 7.56679, 10.26333, 10.21464, 
    1.259433, -0.0954951, 0.3436172, 0.3889436, 0.3328735, 2.681817, 
    3.837993, 5.1575,
  90.34059, 66.30574, 56.15143, 46.72179, 31.81917, 16.57863, 10.32136, 
    10.37988, 4.12169, 3.327969, 0.5509236, 0.3129369, 0.6347235, 2.240233, 
    4.307891,
  100.3274, 76.20246, 61.37107, 52.08746, 56.41391, 48.37729, 17.26945, 
    8.281069, 4.854741, 2.854274, 1.615025, 0.3979927, -0.2194347, 
    -0.2684039, 0.848268,
  107.6398, 77.49471, 65.5695, 58.96395, 62.00769, 53.18819, 32.05578, 
    7.687101, 3.744697, 2.092644, 0.8045279, 0.2660027, -0.3313507, 
    -0.2421832, 0.8665036,
  105.6097, 85.97968, 84.54659, 68.85693, 54.97475, 35.92559, 11.58811, 
    4.857293, 3.143354, 1.124414, 0.2541626, 0.01306429, 0.02686094, 
    0.8197756, 1.880534,
  100.419, 90.60516, 64.21002, 20.74092, 7.431217, 4.880765, 3.753916, 
    3.956063, 1.449094, 0.2595717, 0.02604047, 0.05242974, 0.1345348, 
    0.4503486, 0.8572792,
  11.83619, 22.99591, 12.36693, 14.84892, 13.10919, 3.693322, 4.173384, 
    4.25271, 8.515423, 1.532866, -0.2435024, 0.07870225, 0.004271477, 
    0.2770025, -0.1017341,
  19.50448, 16.19491, 16.21157, 14.78753, 8.915738, -0.4193445, 0.421266, 
    0.2212876, 2.062337, 3.771689, -0.1256625, 0.1706998, 0.9723972, 
    -0.007753437, -0.3007939,
  67.19077, 22.1488, 14.92296, 14.19353, 11.95963, -0.9090081, -0.5610941, 
    -0.4232486, 0.175795, 1.256115, 0.8851469, 0.667051, 1.818213, 2.209314, 
    0.9972326,
  79.15439, 81.35339, 64.94257, 24.69242, 12.27971, 13.16549, 0.1849137, 
    -0.435004, -0.1639811, 0.6681167, 0.6434435, 0.8942712, 2.51711, 
    2.588857, 1.88757,
  72.07687, 67.84425, 71.39023, 52.29934, 8.027168, 11.02086, 13.63384, 
    1.083637, 0.2285142, 0.5551902, 0.5845169, 0.5672135, 2.099679, 2.765115, 
    3.857199,
  73.97555, 67.15411, 61.75819, 47.82977, 28.65155, 10.30993, 8.473467, 
    9.164921, 2.873649, 1.310981, 0.5352521, 0.2718397, 0.6062523, 1.744136, 
    2.773165,
  78.49584, 70.20548, 61.58579, 48.2364, 49.62294, 44.58906, 15.66588, 
    6.133017, 2.242143, 1.085201, 0.6055212, 0.1849464, 0.08927092, 
    0.4724765, 1.083649,
  78.94669, 62.76155, 56.73933, 43.33948, 48.02684, 54.00951, 34.44335, 
    6.227245, 2.001958, 0.6992696, 0.07335107, -0.0701769, -0.2028826, 
    0.3515594, 1.651679,
  63.07409, 48.41979, 55.33009, 46.68198, 41.67961, 32.44452, 11.10764, 
    3.536266, 1.268302, 0.5148509, -0.01234477, -0.1591747, -0.1405032, 
    0.5044838, 0.9399914,
  65.28851, 65.236, 45.36783, 12.87227, 4.832604, 2.77896, 2.479931, 
    1.783077, 0.4284729, -0.01031226, -0.104773, -0.04862448, -0.01024742, 
    0.2709261, 0.890308,
  10.8392, 23.21521, 12.56945, 17.47039, 25.44368, 8.186007, 6.53209, 
    8.798946, 22.01563, 9.200668, 2.004982, 4.127731, 1.77433, 1.399245, 
    -0.2551858,
  15.50376, 18.90195, 17.34176, 28.74774, 25.67242, 3.863486, 5.702753, 
    6.390363, 12.54282, 17.29476, 3.101218, 4.8781, 7.460557, 0.7814217, 
    -0.4133363,
  53.22631, 22.10369, 20.62799, 27.91838, 26.59956, 2.081108, 2.181812, 
    3.501578, 5.276311, 7.835544, 6.057002, 3.451842, 4.735728, 5.949153, 
    1.719577,
  82.15392, 96.11846, 73.99022, 32.01351, 22.43459, 21.38559, -0.1357147, 
    0.2669183, 0.5456308, 0.6203493, 0.4724799, 0.6771669, 2.428495, 
    3.277301, 1.578358,
  82.02149, 79.20547, 89.00423, 62.72267, 14.10935, 13.43366, 15.40137, 
    0.5202878, -0.2200069, 0.1832183, 0.2684982, 0.7977595, 1.317373, 
    2.021243, 2.239004,
  80.1842, 72.31213, 72.96432, 57.06808, 34.49603, 11.17569, 10.3083, 
    10.25164, 3.117356, 1.318091, 0.7348217, 0.6641459, 0.7924606, 1.249391, 
    1.840172,
  93.46763, 77.99214, 62.35846, 49.86139, 54.42788, 43.26928, 13.13167, 
    4.02714, 1.805032, 1.212473, 0.6631275, 0.2012716, 0.137136, 0.7355942, 
    1.200694,
  106.0354, 105.9277, 79.63313, 52.22376, 45.51665, 45.14109, 21.37033, 
    3.047945, 1.055532, 0.1171535, -0.5078809, -0.5689842, -0.6346155, 
    -0.1452589, 0.6766188,
  78.66259, 90.46304, 61.49598, 41.68807, 39.43059, 24.65677, 5.984545, 
    1.965793, 0.8886191, 1.249473, 0.7979415, 0.3172632, 0.2400873, 1.074226, 
    0.3525315,
  51.87991, 56.40879, 39.53695, 11.04988, 3.61424, 2.947459, 3.757467, 
    3.586523, 2.168127, -0.1207415, 2.588243, 3.743545, 0.856315, 1.740583, 
    1.422594,
  4.861222, 15.72794, 8.713657, 13.87104, 28.10395, 8.412468, 3.401807, 
    5.312284, 12.45551, 5.430481, -0.3722726, 1.841876, 3.440318, 3.334133, 
    0.5342036,
  5.774328, 12.7903, 12.84588, 33.15369, 28.07406, 7.556361, 5.44016, 
    5.456695, 9.284754, 13.81939, 0.9448144, 4.85483, 12.3669, 2.732349, 
    0.1659373,
  37.72918, 19.8348, 19.14215, 36.63178, 30.1344, 3.363928, 5.483388, 5.731, 
    7.249324, 8.090333, 5.738497, 5.021003, 8.674994, 14.26111, 6.517949,
  73.50238, 85.81784, 65.58782, 31.68972, 31.66522, 24.45702, 0.6530718, 
    2.892592, 2.925189, 3.932106, 3.41364, 4.25672, 7.62671, 9.091498, 
    8.308447,
  71.13004, 65.51322, 72.9939, 40.91003, 16.80278, 18.53588, 17.55744, 
    -0.1641239, -1.557237, -0.5303828, 0.4029958, 0.9742602, 4.191885, 
    6.414646, 6.76476,
  74.98309, 53.65291, 46.3551, 30.98924, 17.93388, 8.669602, 9.815477, 
    10.69413, 2.878281, 0.9714341, -0.1267242, -0.4928004, 0.6096256, 
    1.877695, 3.726814,
  86.84468, 63.65748, 42.98892, 28.22618, 31.22551, 21.67572, 4.559857, 
    2.212714, 1.6271, 1.227969, 0.7491938, -0.06552706, -0.2772889, 
    -0.3335385, 0.8545909,
  76.75304, 56.19761, 47.66187, 35.12498, 37.88404, 39.89046, 18.84997, 
    1.343487, 2.461893, 0.6637682, -0.4372057, -0.5894601, -0.6160679, 
    -0.6372433, 0.1305282,
  71.32171, 64.25014, 46.22392, 34.89961, 30.77222, 24.76188, 6.841307, 
    3.661548, 1.81673, 1.136982, 0.8942366, 1.183867, -0.1093379, -0.3874333, 
    -0.6871905,
  76.6328, 69.32568, 44.71354, 14.40037, 6.881322, 5.364603, 3.974302, 
    4.010021, 1.722203, 0.123343, 2.164967, 2.935886, 1.216502, 1.592733, 
    0.1165873,
  -0.4273238, 3.276105, 0.03714529, 7.815932, 22.56041, 8.368209, 2.229458, 
    -0.2223839, 2.402169, 1.407232, 0.5042242, 1.851164, -0.4084104, 
    -0.2439892, -1.987758,
  0.8666633, 2.445336, -0.05024532, 17.47935, 18.34064, 4.691138, 4.701615, 
    3.912, 2.774121, 3.363321, 0.6883966, 0.8212711, 4.624248, -0.2235038, 
    -1.426507,
  21.96124, 8.570964, 0.9271173, 13.6664, 15.92388, 2.285938, 3.932944, 
    5.683958, 6.296341, 5.112996, 0.4483516, 0.6825258, 2.532755, 4.929281, 
    1.41396,
  70.73785, 61.11496, 19.70867, 5.593863, 14.19547, 11.39392, 0.502667, 
    2.616303, 4.110201, 4.609333, 4.581661, 3.259047, 3.052796, 3.512667, 
    2.781576,
  83.0798, 53.03295, 31.71466, 7.657673, 4.27426, 7.55847, 8.891111, 
    0.5593026, -0.6344045, -0.1175535, 1.130353, 2.003499, 4.986237, 
    5.095906, 4.598041,
  88.2558, 53.68273, 19.18872, 9.671991, 7.041349, 5.102061, 5.994498, 
    6.053902, 1.773229, 0.9824852, -0.2370408, -0.1562546, 0.6675343, 
    3.864242, 6.073554,
  82.28978, 46.82551, 28.08831, 19.98647, 21.08026, 17.62513, 5.865068, 
    2.353285, 2.198824, 1.509286, 0.6788749, 0.1268783, -0.05238351, 
    -0.1083458, 2.810174,
  63.82428, 46.81022, 43.69988, 31.15797, 27.85072, 28.36303, 12.84109, 
    3.661087, 2.947954, 2.551395, 1.125887, 0.3208056, -0.05918572, 
    -0.2778388, 0.396659,
  58.48931, 53.84549, 49.07985, 27.82285, 19.38963, 12.41728, 3.331457, 
    1.673977, 2.304894, 2.01459, 0.5831644, 1.657123, 0.6305035, 0.06151982, 
    0.2031639,
  54.33384, 47.43537, 27.93066, 6.326366, 2.756556, 2.605112, 2.145129, 
    1.223187, 1.154724, 0.7802762, 0.6078269, 0.9487783, 1.209023, 0.2221872, 
    0.3256447,
  3.684631, 4.08075, 0.2859094, 0.8814225, 3.670865, 1.482001, 0.06676659, 
    0.4260716, 3.098648, 3.423337, 1.571887, 2.57142, 1.200672, -0.3889331, 
    -1.156935,
  8.090662, 4.995725, 1.237493, 3.172431, 3.413388, 0.1351701, 0.7175878, 
    0.9980589, 4.476013, 5.141616, 2.422787, 4.043149, 4.86408, 1.703099, 
    0.649738,
  28.14509, 11.06774, 4.303152, 4.353348, 3.84983, -0.05945795, 0.4164984, 
    0.8683228, 1.853719, 2.922011, 1.690247, 2.106673, 4.567719, 4.659844, 
    2.916863,
  76.15073, 78.01968, 47.31974, 7.551461, 3.509595, 3.027906, 0.3226441, 
    0.5768516, 0.6866046, 1.00811, 2.055053, 2.561825, 2.849086, 1.399809, 
    1.482209,
  89.46608, 74.28904, 70.88906, 23.9317, 2.239194, 2.048493, 4.06191, 
    0.6275893, 0.140651, 0.2652193, 0.4978381, 1.270947, 3.132858, 3.093828, 
    2.558681,
  98.51198, 82.23742, 60.99824, 31.44277, 7.151089, 2.523163, 3.451585, 
    4.578448, 2.423858, 1.198637, 0.335195, 0.3899222, 1.247271, 2.423773, 
    4.988541,
  100.6584, 92.73135, 74.49662, 43.98015, 33.49788, 15.67307, 5.273983, 
    3.104388, 2.937211, 2.847014, 1.049616, 0.5768713, 0.4482953, 0.66857, 
    2.445466,
  98.1997, 90.89803, 76.41012, 50.41419, 36.13034, 27.51586, 11.66159, 
    3.276643, 2.460793, 2.818633, 1.43196, 0.2702031, -0.01547746, 0.2239985, 
    1.392993,
  90.26559, 85.62133, 72.52638, 42.96567, 24.17389, 8.20799, 3.419057, 
    2.925812, 3.483984, 1.735618, 1.228108, 0.2986873, -0.0743221, 
    0.08416065, 1.16037,
  75.9727, 69.05685, 43.4494, 6.573717, 1.028726, 0.3326435, 3.746036, 
    4.241874, 2.156991, 1.42913, 1.467996, 0.556071, 0.124756, -0.0443415, 
    0.8406942,
  2.351553, 4.009615, 2.252579, 2.773167, 3.418243, 0.7811267, 0.3033568, 
    0.7897016, 4.51555, 3.922743, 1.947094, 2.780937, 2.385322, 0.5208082, 
    -0.2309592,
  7.033609, 4.907873, 3.99912, 5.865242, 5.584814, 0.2020098, 0.3694468, 
    0.5192615, 2.066455, 4.119112, 2.518719, 6.638576, 5.903725, 2.023, 
    0.06259236,
  14.65076, 11.42974, 7.06249, 12.19302, 11.7059, 0.2011797, 0.3500323, 
    0.5695592, 0.926734, 0.9757853, 1.233881, 3.961579, 5.72313, 8.545634, 
    4.072796,
  52.2044, 54.09664, 47.34865, 21.73653, 16.98277, 11.42955, 0.4346025, 
    0.2204999, 0.3791922, 0.5076889, 0.5198283, 1.650355, 3.076025, 3.758928, 
    2.228349,
  62.53919, 51.51494, 62.72518, 45.48926, 14.68581, 10.9688, 10.12974, 
    1.36328, 0.2758661, 0.2082997, 0.3471243, 0.8529164, 2.091373, 2.453037, 
    2.797,
  73.36969, 59.65648, 49.83633, 47.68164, 26.11435, 8.893585, 5.215225, 
    3.406776, 0.9360161, 1.153316, 0.2727052, 0.5604218, 1.179755, 1.867801, 
    2.812186,
  73.85642, 69.85751, 59.67293, 49.28366, 57.87881, 36.09228, 2.929753, 
    0.5257015, 1.314473, 2.111635, 1.029456, 0.4297367, 0.6258087, 0.750742, 
    1.669497,
  65.48328, 65.07365, 59.5294, 50.8446, 61.0148, 52.30626, 7.315322, 
    0.9297743, 2.25244, 1.496498, 0.447577, 0.8896948, 0.2274915, 0.2583407, 
    1.781682,
  52.554, 56.53284, 52.99469, 41.20096, 40.08561, 17.01281, 0.8471344, 
    1.373711, 1.865311, 1.322642, 0.1417222, 0.9669469, -0.006519757, 
    0.08748209, 1.892817,
  45.02328, 42.18379, 29.76134, 8.988804, 4.740166, 2.59306, 0.3842889, 
    2.5689, 0.5976768, 0.08462161, 0.8771222, 0.396146, -0.02472048, 
    -0.06328566, 1.138373,
  2.300995, 2.361568, 2.426171, 2.753386, 3.254011, 1.419723, 0.3907295, 
    1.480547, 6.723227, 2.931984, 2.458729, 4.384097, 3.375063, 2.510935, 
    0.3267907,
  3.477895, 2.291207, 2.419004, 5.856915, 5.035282, 0.738941, 0.3723212, 
    0.6994641, 2.767679, 5.497154, 2.627797, 7.957488, 8.407701, 0.2391775, 
    0.5286603,
  8.39947, 6.221568, 8.420113, 12.41463, 13.57286, 1.054223, 0.8038583, 
    0.3653117, 0.5799308, 0.7570009, 1.852075, 4.971475, 5.331409, 5.89567, 
    1.715951,
  23.42164, 32.53154, 37.64045, 18.74732, 14.3918, 13.952, 1.054239, 
    -0.03430216, 0.07490564, 0.4031581, 1.061761, 2.234338, 2.754371, 
    2.228328, 1.192048,
  29.22384, 32.09546, 52.83768, 34.63951, 11.39, 10.87491, 16.20868, 
    0.3930405, -0.3128931, -0.04455961, 0.04794206, 0.5209416, 1.378732, 
    1.50446, 1.38361,
  33.18467, 39.53269, 48.71627, 40.64257, 21.31288, 9.947336, 10.56124, 
    9.979589, 4.886375, 4.122796, 0.1381256, -0.05657944, 0.50638, 1.328853, 
    1.624983,
  31.35317, 51.01718, 57.55498, 46.51522, 44.36878, 31.41408, 6.657743, 
    1.979375, 3.734653, 4.597652, 1.683388, 0.1253376, 0.443267, 1.001837, 
    1.754642,
  34.6623, 55.59682, 60.47985, 49.39672, 53.44055, 46.13645, 12.62778, 
    2.198033, 3.163447, 2.047927, 0.444139, 0.505592, 0.1049719, 0.451748, 
    2.535789,
  35.42574, 56.28335, 61.58158, 46.97224, 45.6629, 29.00507, 5.040436, 
    2.841676, 2.768405, 0.8075979, 0.3009181, -0.003995119, 0.002969628, 
    0.3315992, 2.392484,
  28.99605, 37.72072, 36.60376, 9.796973, 2.215836, 4.19385, 3.002904, 
    4.589749, 1.887634, 0.1943022, 0.1585017, -0.03325316, -0.004004086, 
    0.03311896, 1.416927,
  4.883693, 4.102324, 2.75677, 3.156696, 1.764416, 0.9792817, 0.6125085, 
    0.4776635, 3.001575, 2.534261, 3.342364, 5.290596, 2.974765, 1.283951, 
    -0.6221771,
  8.595101, 4.666385, 3.254221, 5.106872, 2.499079, 0.4799702, -0.3225281, 
    0.04333827, 2.159887, 4.401349, 3.655995, 8.066654, 10.38057, 0.1424071, 
    -0.6209782,
  16.4099, 3.804045, 5.426168, 9.423949, 8.677708, -0.09701408, 0.3049491, 
    -0.01387185, 1.294527, 2.577166, 5.258713, 6.871713, 8.670003, 8.689172, 
    2.520248,
  37.11533, 34.73862, 30.98181, 19.57974, 10.09529, 7.470888, 0.6704596, 
    -0.09582085, 0.204854, 1.528606, 3.874446, 6.405844, 7.001568, 6.043038, 
    3.018545,
  43.14322, 40.28235, 58.90965, 41.12901, 5.278722, 4.867928, 12.01766, 
    1.32122, 0.4448565, 0.9084683, 2.130006, 4.247341, 4.700891, 4.641981, 
    3.063535,
  57.99453, 58.21171, 59.69763, 44.87881, 11.50875, 4.056562, 5.896285, 
    11.05785, 9.159115, 8.26519, 2.153447, 1.914432, 2.184474, 2.585407, 
    1.674746,
  77.95793, 83.74498, 78.25047, 47.58453, 29.50572, 22.99711, 9.364751, 
    8.816206, 7.301561, 7.467116, 4.714387, 2.329598, 0.4463904, 0.8447622, 
    1.690895,
  96.53639, 92.40634, 79.69035, 48.04139, 43.52765, 48.53591, 17.44327, 
    8.275489, 5.465236, 3.684618, 2.09626, 1.249537, -0.2039489, 0.5911705, 
    2.086097,
  101.4362, 96.08561, 76.37713, 50.45122, 52.06279, 35.97363, 12.98441, 
    6.783604, 3.196595, 1.024756, 0.5562966, 0.151096, -0.2694436, 0.5284119, 
    1.919554,
  92.11091, 81.27283, 60.18583, 14.59058, 2.935287, 7.479004, 8.520308, 
    5.169296, 1.781313, 0.2967876, 0.1051744, 0.09877828, -0.08473895, 
    -0.007272923, 1.223932,
  4.668708, 6.849855, 6.42121, 4.674072, 1.564188, -0.4880522, 1.817666, 
    2.882821, 4.445787, 1.952995, 1.410568, 2.08726, 1.137238, 1.258354, 
    -1.472813,
  5.830475, 5.749892, 6.120476, 4.86586, 1.267497, 1.021889, 2.18447, 
    2.672678, 4.02611, 2.684999, 1.278315, 4.809789, 7.477136, -0.2392289, 
    -0.9640595,
  12.61083, 7.921938, 7.337439, 7.754283, 11.44298, 2.194594, 2.004274, 
    2.018594, 1.302177, 0.416637, 1.478555, 3.886358, 6.639899, 8.897132, 
    3.867942,
  45.0276, 45.25999, 36.8357, 20.71714, 19.51031, 14.38188, 1.345029, 
    0.5466756, -0.3194268, 0.2642373, 1.390062, 3.589552, 6.200471, 7.13942, 
    5.556482,
  66.96138, 59.03704, 72.73389, 46.94592, 19.1413, 15.72889, 15.72932, 
    1.909995, 0.05380915, 0.4565151, 1.845281, 3.449103, 6.069872, 7.640751, 
    8.031403,
  92.7716, 84.33831, 75.89066, 59.0121, 31.71758, 13.84073, 13.14981, 
    10.5321, 5.652829, 5.240585, 2.508447, 3.575984, 4.628502, 6.024165, 
    7.255136,
  108.2574, 102.4792, 90.29147, 67.28561, 60.00935, 43.19684, 12.60972, 
    9.185802, 6.617886, 6.565799, 5.173086, 4.316753, 3.711812, 4.717747, 
    6.422554,
  113.3079, 105.3056, 94.24276, 79.52562, 79.60015, 68.40063, 16.88849, 
    8.494495, 6.281794, 4.512864, 3.977029, 3.2905, 1.600385, 3.010233, 
    4.502589,
  101.4707, 101.2459, 94.47416, 80.59113, 76.22179, 46.33571, 13.42437, 
    8.170601, 4.79352, 2.746018, 1.702099, 1.517549, 0.1362019, 1.77257, 
    2.112885,
  77.76922, 77.12516, 65.1589, 26.04194, 6.098595, 9.766381, 8.691834, 
    6.603673, 3.535313, 1.08321, 0.1616936, 0.5088454, -0.08313687, 
    -0.08930721, 1.293219,
  3.100008, 4.099173, 6.133759, 9.541554, 11.57551, 3.299335, 2.485725, 
    4.432418, 5.736284, 3.638894, 3.029941, 5.889144, 3.796546, 3.29522, 
    0.6332447,
  3.844487, 3.429998, 3.371543, 13.66193, 10.21906, 2.997845, -0.01868136, 
    0.5383117, 0.9276854, 1.661077, 0.5970407, 4.462331, 6.04478, 1.800521, 
    -0.12504,
  18.28401, 3.608126, 3.580051, 11.68506, 14.95634, 0.971024, 0.6138013, 
    0.6070004, 0.6556183, 0.3046237, 2.065961, 4.49679, 6.315914, 8.341487, 
    4.436844,
  55.13063, 65.32529, 52.32653, 20.45237, 23.38254, 17.97648, -0.3967291, 
    0.05149603, 1.182914, 0.5454715, 1.085775, 3.531743, 6.041306, 8.475038, 
    6.699168,
  65.88514, 68.60415, 83.06216, 43.74836, 17.27627, 24.22329, 20.22432, 
    0.6013698, -0.9046689, 0.2042826, 1.848462, 1.869702, 5.392762, 8.379976, 
    8.711992,
  72.3456, 73.88579, 77.43362, 59.28424, 28.77593, 20.93573, 23.71957, 
    18.85182, 8.196144, 3.396592, 0.7246168, 1.143585, 3.290339, 5.237389, 
    5.163613,
  71.78493, 80.18375, 86.14674, 77.00641, 73.81576, 45.456, 18.44542, 
    14.23652, 8.536168, 4.510201, 2.040801, 1.824845, 2.559567, 3.656407, 
    5.05996,
  69.10917, 74.71553, 80.36491, 85.32169, 95.73299, 73.33387, 15.44874, 
    10.08299, 7.975521, 4.980104, 2.257447, 2.261472, 1.797465, 3.897358, 
    5.665244,
  66.03913, 69.08877, 68.91737, 68.62911, 70.60031, 35.88372, 10.60319, 
    8.452637, 7.003137, 4.869344, 2.687916, 3.006421, 2.758023, 4.521598, 
    4.214575,
  59.67851, 55.26898, 42.98279, 16.29581, 4.988076, 5.49485, 6.567346, 
    7.42759, 5.244138, 1.516068, 0.5355871, 1.759651, 2.141913, 2.268962, 
    2.770617,
  3.786617, 0.8278634, 0.7791872, 0.9905252, 3.362811, 1.338477, 0.3684489, 
    0.471951, 1.658003, 0.2158145, 1.808434, 2.153279, 1.414801, 0.9828026, 
    1.637991,
  5.184176, 0.4311159, 1.231067, 2.838351, 4.474618, 0.7996763, 1.079712, 
    0.1315162, 0.7755572, 1.087053, 0.5803766, 3.663506, 3.790093, 0.1825817, 
    1.220953,
  9.171069, 1.749374, 2.905763, 4.618219, 8.355799, -0.2220231, 1.362524, 
    2.495358, 1.674017, 1.714796, 2.648196, 5.009607, 4.799857, 3.159851, 
    4.934968,
  28.12668, 38.21116, 38.48243, 8.401937, 15.37255, 10.99036, -0.4236094, 
    1.446497, 2.675229, 2.81153, 5.121954, 6.299585, 6.207986, 5.184294, 
    6.591967,
  29.68461, 30.5533, 50.15492, 29.95018, 10.91608, 15.40176, 13.51394, 
    -0.4063004, -0.4143673, 1.774595, 4.856896, 5.330851, 6.795208, 5.870798, 
    8.145043,
  31.01435, 25.59237, 35.26314, 37.00967, 21.02713, 14.27472, 15.00632, 
    8.829243, 3.436631, 3.264296, 0.9343172, 3.404771, 5.817935, 6.173594, 
    6.362609,
  28.70747, 24.5754, 29.88685, 40.75003, 50.58478, 29.75536, 10.84933, 
    6.25296, 3.084437, 2.133439, 1.010957, 1.56967, 3.181698, 3.250814, 
    4.603945,
  28.22808, 20.76215, 21.60999, 38.2442, 57.41748, 43.34024, 7.951873, 
    4.681819, 3.239569, 1.142235, 0.1608018, 0.595297, 1.031427, 1.630651, 
    2.585516,
  24.29605, 18.38501, 15.90413, 24.03548, 42.64967, 17.14012, 5.46073, 
    3.30488, 2.804355, 1.236741, -0.1602671, -0.01561482, 0.2735596, 
    1.143487, 1.990149,
  15.26146, 9.212502, 5.018726, 3.109477, 7.247283, 2.925599, 2.814787, 
    3.641155, 2.274778, -0.02461991, -0.5624911, -0.4997331, -0.1748355, 
    -0.1148544, 1.005016,
  -0.6028699, 1.517733, 7.588304, 5.87142, 2.129146, 0.9563702, 0.3062836, 
    0.4904389, 2.333215, 1.108399, 2.381243, 3.288762, 2.498851, 2.230231, 
    0.06299105,
  -1.633554, 3.61223, 9.695563, 6.872405, 2.585436, 0.8588639, 0.2582201, 
    -0.1892339, 0.5751101, 1.710769, 1.402354, 3.244408, 5.698324, 0.3604001, 
    -0.3354633,
  -5.067599, 6.494913, 12.54507, 8.85272, 7.89408, 0.5430618, -0.05197317, 
    -0.775255, -0.09861023, 0.4866236, 1.725611, 3.204885, 3.079217, 4.05607, 
    2.925479,
  0.2354597, 25.60706, 41.09566, 15.04557, 11.56073, 8.328782, 0.5339527, 
    -0.3435651, 0.3658124, 0.8942069, 2.10204, 2.900415, 3.808108, 3.998188, 
    6.072144,
  10.87835, 26.81026, 61.75676, 38.87823, 14.54752, 13.37702, 10.27526, 
    -0.04838913, -0.5429714, 0.141965, 0.8197838, 2.219501, 6.228166, 
    7.604512, 9.522365,
  27.37496, 32.56651, 51.29385, 59.10408, 31.22532, 17.42676, 15.9252, 
    8.637461, 1.942776, 2.421789, -0.4220669, 1.989762, 6.720506, 7.898459, 
    9.875306,
  40.61568, 49.72939, 64.57462, 78.43969, 76.80183, 39.7756, 15.07228, 
    5.673485, 2.109687, 1.838778, -0.004289802, 0.9692703, 2.682272, 
    4.077904, 6.794394,
  54.3243, 62.11516, 70.81566, 91.73597, 96.19634, 61.8841, 12.95025, 
    6.172598, 2.469671, 0.6730853, -0.2067067, 0.0808302, 0.3139282, 
    2.205702, 3.876223,
  61.07602, 67.85934, 74.40559, 92.56882, 90.46246, 35.54125, 10.48653, 
    5.437595, 2.387531, 0.1851862, -0.6221381, -0.5429806, -0.4323131, 
    0.7340401, 3.911272,
  57.4537, 58.22273, 57.0379, 45.99911, 20.0841, 9.128695, 5.91441, 5.456153, 
    1.472142, -0.9368068, -1.497058, -1.383981, -0.6783106, 0.1359821, 
    2.997884,
  7.318686, 10.84064, 6.729604, 5.433356, 5.80046, 3.105603, 1.86235, 
    0.072451, 0.6814735, 1.068785, 2.127643, 3.146497, 1.831392, 1.042432, 
    -0.3510335,
  18.1126, 10.11779, 8.081397, 6.218411, 4.937365, 2.155654, 2.136831, 
    -0.4588808, 0.0185537, 0.1728484, 0.7100097, 2.375489, 3.881108, 
    -0.3877048, -0.7312545,
  64.48603, 16.19795, 10.12402, 10.46791, 9.678364, 0.2211054, 0.4764669, 
    -0.1013228, 0.8620815, 0.1454703, 1.038417, 2.287936, 2.375898, 3.954909, 
    1.932591,
  93.79971, 83.24054, 54.83145, 18.02868, 22.30338, 15.98337, -0.0486377, 
    1.502033, 3.638739, 3.675715, 2.940939, 2.746523, 3.206758, 4.52855, 
    3.150389,
  106.0666, 91.95938, 94.41954, 42.57404, 23.60519, 23.54159, 20.41924, 
    -0.7922622, -0.6994917, 2.887318, 4.340294, 4.982509, 6.37614, 7.749938, 
    9.141271,
  115.828, 100.4216, 88.0771, 56.97961, 32.03094, 23.11051, 22.86636, 
    17.5422, 5.99636, 4.603033, 1.922287, 3.856361, 5.139132, 5.94202, 
    8.060028,
  118.88, 113.1295, 100.4654, 75.4794, 74.52648, 33.86583, 19.03415, 
    12.30143, 7.055051, 4.925736, 3.489358, 3.458104, 4.065313, 4.14416, 
    5.842474,
  122.9565, 116.7438, 106.7367, 94.69292, 99.78172, 54.39201, 16.28388, 
    10.58971, 6.386002, 3.379349, 2.402856, 3.509658, 2.634903, 4.090534, 
    4.960438,
  122.568, 119.7371, 114.6406, 102.5154, 89.97865, 33.33917, 13.96584, 
    8.226449, 6.879876, 6.010885, 2.381555, 2.111883, 3.20966, 4.418206, 
    8.385304,
  117.5825, 113.7722, 102.4789, 55.98895, 21.13209, 12.99303, 6.482527, 
    13.99813, 7.651762, 2.25122, 0.9960874, 1.873787, 2.331853, 3.847841, 
    9.104542,
  4.824709, 7.36099, 10.97393, 10.15679, 1.943771, 1.522736, 0.2311996, 
    0.5992182, 0.5546879, 0.09974568, 0.5680224, 1.426171, 1.729578, 
    1.943739, -0.1633599,
  5.767891, 2.044913, 9.106802, 10.18109, 5.229106, 0.9267544, 1.111531, 
    0.339122, 1.044386, 0.4706256, 0.6310326, 1.97287, 4.237631, 0.9372703, 
    -0.01042539,
  35.19564, 6.163779, 6.621233, 17.05257, 15.35847, 0.1039428, 1.426925, 
    1.547173, 2.107789, 1.497252, 2.012168, 1.956168, 2.414199, 4.803495, 
    2.814204,
  66.6483, 65.5153, 45.71462, 22.25013, 27.92909, 18.39972, 0.8234559, 
    1.891659, 2.946154, 1.995354, 4.080049, 3.492318, 2.680469, 4.24701, 
    3.700963,
  81.49687, 75.99548, 79.7112, 34.34558, 24.68509, 24.79478, 20.86877, 
    0.06591882, 0.3148839, 0.869074, 2.434841, 3.937008, 3.945552, 4.077097, 
    5.046245,
  91.9594, 84.89751, 76.25156, 50.50771, 34.74559, 23.33096, 19.48069, 
    11.09611, 4.907143, 1.503306, 0.7292252, 1.179138, 5.109678, 4.153013, 
    4.187423,
  99.46354, 101.3562, 94.25571, 76.53255, 79.43056, 32.03046, 17.75087, 
    8.227773, 6.509311, 5.017823, 1.107644, 1.162715, 0.9593285, 2.175733, 
    3.289807,
  105.6655, 109.2395, 108.6018, 103.0275, 106.7792, 48.14185, 16.12048, 
    6.45777, 4.02384, 6.04216, 3.744202, 1.045004, 0.7574002, 1.467597, 
    1.573552,
  107.5763, 113.3946, 117.3164, 112.7635, 79.12921, 28.47614, 17.83411, 
    8.119097, 7.792799, 9.897443, 5.312364, 2.048369, 0.8791103, 1.654514, 
    2.20784,
  102.2295, 106.6313, 95.88714, 41.98183, 15.0934, 15.34169, 12.47494, 
    26.59154, 17.86773, 6.380649, 1.609595, 2.004822, 1.487556, 2.149907, 
    3.25196,
  5.285139, 3.748814, 4.532318, 5.670751, 1.951017, 1.567717, 0.9676319, 
    1.942033, 1.736056, 0.5214776, 1.034697, 1.493221, 0.5350586, 0.8531367, 
    -0.07032847,
  3.874789, 1.433203, 7.987153, 9.625844, 4.591314, 1.996761, 0.9818811, 
    0.806678, 0.9000989, 1.67931, 1.389567, 2.066661, 2.353095, -0.346195, 
    -0.3980517,
  23.67856, 3.11483, 3.092916, 12.88925, 13.72591, 1.472495, 1.136783, 
    0.782811, 1.031044, 0.6069379, 1.105001, 1.425665, 1.550608, 3.219422, 
    1.553978,
  60.72243, 52.48366, 35.67108, 12.34489, 21.27707, 11.33092, 0.4966468, 
    1.433536, 2.455431, 2.05977, 2.28374, 2.009116, 2.139485, 4.279339, 
    2.59477,
  81.73034, 74.71846, 74.13635, 28.47614, 19.03768, 20.13288, 13.91847, 
    0.05407612, 0.15927, 2.811097, 2.334413, 2.023052, 2.065185, 4.141603, 
    5.171132,
  97.16325, 88.22865, 77.59306, 45.52495, 31.71294, 22.08353, 16.25514, 
    5.504369, 3.679429, 2.93278, 1.042741, 2.377719, 1.638199, 3.896314, 
    6.079379,
  106.9651, 105.9587, 100.0325, 76.57029, 79.0815, 28.05847, 15.78863, 
    6.787226, 6.179605, 4.536752, 1.482008, 1.909627, 1.272145, 2.031934, 
    5.441141,
  113.7856, 114.5183, 112.5392, 107.7332, 103.8542, 36.42612, 16.13631, 
    8.977583, 7.422339, 5.15835, 3.166581, 1.516614, 2.199187, 2.147871, 
    4.257576,
  113.491, 115.8434, 116.8499, 104.2326, 55.63613, 18.63796, 13.937, 
    12.13492, 12.72903, 11.72709, 3.98648, 1.05267, 1.265082, 2.042032, 
    4.113522,
  103.6393, 102.1735, 80.69353, 28.0724, 10.85872, 11.35567, 11.11989, 
    37.05957, 25.48475, 10.38622, 1.54705, 1.041537, 1.19467, 1.949237, 
    2.82735,
  7.528659, 6.394569, 4.231641, 3.536368, 4.196097, 2.061661, 0.9271627, 
    1.0963, 1.600368, 1.960997, 3.58461, 4.664391, 3.01344, 2.846281, 
    0.4142387,
  7.993546, 3.666073, 4.593429, 4.009929, 3.723494, 1.097299, 0.591141, 
    1.209564, 1.371129, 2.217343, 3.748157, 6.196518, 6.563229, 2.144306, 
    0.167623,
  29.98208, 4.065713, 5.905755, 6.937643, 7.304817, 0.837226, 0.8524007, 
    0.9684073, 0.9398182, 0.571797, 1.720054, 2.86982, 3.215818, 3.794856, 
    1.58367,
  56.16795, 47.80771, 29.25559, 8.83627, 17.85647, 8.510339, 0.3268602, 
    1.34399, 1.264472, 2.031605, 2.137275, 2.569014, 2.943532, 3.652306, 
    2.143026,
  69.84217, 63.45285, 62.67034, 18.3849, 12.9831, 13.86917, 8.647532, 
    0.2810959, 0.1868224, 3.371208, 4.076894, 2.588528, 1.982133, 2.301776, 
    3.350608,
  68.85592, 63.88346, 55.77436, 31.57676, 22.3257, 14.38694, 10.97648, 
    6.086995, 3.374323, 1.854836, 0.7273425, 1.529891, 1.4074, 2.367737, 
    2.930608,
  65.2249, 67.88283, 66.16308, 51.42847, 56.32231, 17.32176, 9.317806, 
    6.18602, 5.212429, 2.859483, 0.8890572, 0.951853, 1.217256, 1.678709, 
    3.695765,
  63.20224, 68.47717, 71.18243, 71.16914, 67.00467, 19.17788, 8.466969, 
    5.748768, 4.655041, 3.196281, 1.465516, 0.9458634, 1.172117, 1.42414, 
    3.645888,
  56.90355, 62.30481, 68.29637, 60.77003, 28.74366, 9.709247, 6.660195, 
    6.322032, 7.76182, 6.782423, 2.428527, 0.6934484, 0.7310641, 1.998205, 
    3.383957,
  53.20149, 54.14106, 47.03406, 17.78683, 6.719689, 6.276511, 6.546012, 
    29.55685, 18.97895, 5.082357, 0.6260036, 0.4148763, 0.4207712, 1.81785, 
    2.755612,
  4.850502, 3.715029, 3.484643, 3.544889, 2.215552, 1.942088, 0.9461548, 
    0.7573617, 0.8786879, 0.4369748, 1.966389, 3.350972, 1.90194, 1.686576, 
    0.7870319,
  4.418643, 2.230198, 2.574523, 2.493595, 1.313597, 0.8688964, 0.5062152, 
    0.7215922, 1.169587, 0.9094969, 0.8174405, 2.346475, 3.431905, 1.553638, 
    0.589952,
  19.17283, 2.467386, 2.21903, 4.696699, 4.107194, -0.3587637, 0.8172749, 
    0.379269, 0.5776908, 0.3294183, 1.081334, 2.806901, 3.660981, 3.595542, 
    2.56513,
  48.5038, 41.94487, 22.30172, 3.726253, 9.04313, 4.919139, -0.6156572, 
    2.194817, 1.642743, 2.166386, 2.698266, 2.499055, 1.961941, 1.940864, 
    1.495513,
  68.53171, 64.14784, 63.00041, 11.59189, 9.036364, 7.442227, 6.424255, 
    -3.036725, -0.6791197, 3.707416, 8.093385, 5.591036, 3.11158, 3.352319, 
    3.765277,
  93.50875, 76.48975, 53.05798, 22.17395, 18.95177, 12.30842, 10.55849, 
    5.068061, 2.744432, 2.57493, 3.15262, 5.967537, 4.107214, 3.610545, 
    3.426885,
  103.3982, 83.55264, 65.51006, 45.33494, 55.7642, 19.60227, 9.303172, 
    7.491072, 4.532809, 4.384219, 3.814455, 4.630567, 5.097586, 3.406405, 
    3.417827,
  96.2045, 78.97001, 75.01481, 71.02224, 69.97356, 22.80568, 9.395497, 
    7.174377, 5.494128, 4.570037, 3.893882, 3.307354, 3.462529, 3.60433, 
    3.027348,
  81.61256, 79.76242, 84.40027, 69.63884, 32.68226, 13.52172, 10.93357, 
    10.91395, 9.858034, 7.531061, 4.426867, 2.670925, 2.95838, 3.463207, 
    1.479509,
  67.24663, 68.06326, 57.68629, 23.46097, 14.07249, 11.6113, 11.69521, 
    34.65848, 23.66191, 4.731172, 3.336362, 3.559617, 0.9704375, 2.307102, 
    0.9573624,
  0.9883307, 1.080438, 2.087926, 1.615033, 0.9280567, 1.632521, 1.492245, 
    1.016651, 0.9453088, 0.2364622, 0.8729611, 1.32013, 0.4410416, 0.6848392, 
    0.1128265,
  1.147584, -0.4424507, 0.08025589, -0.9951419, -3.003913, 0.1115374, 
    1.604519, 3.298189, 2.180052, 2.305278, 3.106663, 3.923657, 2.331158, 
    -0.3035396, -0.1532522,
  26.84565, 3.562199, 2.241441, 1.216942, -2.826556, -0.5721899, 2.126301, 
    2.373783, 3.18741, 2.602002, 2.426391, 3.298259, 2.470993, 2.180933, 
    1.154505,
  82.90778, 70.49482, 31.53517, 4.000267, -1.025565, -1.420977, -0.4311159, 
    3.820894, 4.620136, 4.683168, 5.768, 3.864054, 3.646432, 4.883905, 3.25469,
  98.5244, 68.93769, 48.5838, 4.014882, 3.235893, 4.230677, 4.589463, 
    -1.161544, 0.9521347, 7.511703, 11.84921, 7.181654, 5.390148, 4.681074, 
    5.515906,
  97.33441, 58.8721, 20.67627, 9.07215, 12.44233, 6.264477, 5.698705, 
    1.713189, -0.1906358, -0.5806182, 2.695682, 7.127763, 6.511882, 6.715789, 
    6.102044,
  89.65833, 54.90863, 33.67859, 33.15928, 46.21794, 11.00114, 3.586214, 
    2.934413, 2.826959, 2.597646, 1.84384, 3.082066, 5.12649, 5.17448, 
    5.056757,
  73.41934, 57.16958, 54.84872, 60.17173, 55.21128, 15.4347, 5.661821, 
    4.381782, 3.741886, 1.890396, 2.127206, 2.873435, 4.616548, 4.212647, 
    3.812542,
  72.06872, 70.02728, 70.35423, 56.86324, 24.97804, 10.44588, 7.571742, 
    9.896577, 11.67283, 16.28549, 8.163043, 3.960906, 4.352692, 4.895405, 
    2.413567,
  70.60476, 66.49147, 50.85108, 18.93768, 10.39917, 9.610326, 10.46256, 
    30.51844, 26.10915, 8.601774, 8.991468, 4.343666, 1.400139, 3.755486, 
    2.476792,
  0.9731301, 0.3718249, 0.5944481, -0.0008970905, 4.73108, -0.2146392, 
    4.833642, 1.365021, 1.886499, -0.6463867, 1.896559, 2.260355, 0.7840748, 
    0.9176442, 0.5169712,
  2.345938, 0.05703383, 0.7144285, 1.329552, -2.375367, -2.578068, 3.094835, 
    2.896504, 3.344388, 3.103351, 5.807034, 7.961399, 6.286482, 2.575931, 
    1.85043,
  50.01178, 9.521712, 6.234345, 4.426964, 0.9193082, 3.002578, 4.479799, 
    5.79635, 3.722157, 3.069706, 2.914883, 5.19529, 5.042544, 4.66607, 
    2.114428,
  90.86244, 87.73253, 53.80875, 5.580637, 1.935054, 6.171917, 2.952215, 
    4.04834, 5.808293, 5.749458, 6.154044, 4.3865, 4.195712, 4.608287, 
    5.199652,
  98.54713, 66.85395, 40.33101, 9.81486, 11.81558, 7.988523, 5.842246, 
    0.9098969, 2.323466, 6.765242, 11.78488, 6.516198, 4.345763, 4.244966, 
    5.628799,
  79.59863, 36.91941, 15.63009, 28.59671, 16.84852, 4.927894, 3.219029, 
    2.435232, 0.8780584, -0.3604071, 2.516979, 5.950199, 5.048316, 4.812806, 
    5.061022,
  50.60142, 25.48916, 47.49709, 30.928, 41.10728, 7.211793, 2.554702, 
    1.62325, 0.5524995, 0.3890103, 0.7336062, 1.855902, 2.628482, 2.395838, 
    1.984065,
  36.35589, 58.81057, 44.98701, 48.31343, 48.42033, 10.02787, 4.772476, 
    2.968031, 2.192621, 1.375933, 1.122221, 2.104425, 2.541085, 1.585461, 
    1.806059,
  70.59795, 63.74699, 58.08544, 46.96217, 19.11234, 9.159964, 6.928482, 
    8.698941, 11.05844, 13.19687, 4.38787, 1.555785, 3.204401, 3.071176, 
    0.3806412,
  82.49471, 67.52493, 46.25892, 15.56119, 8.745009, 9.295753, 7.887672, 
    23.33418, 22.44018, 6.956616, 7.362689, 1.682884, 0.2022299, 2.53904, 
    -0.007378838,
  5.937538, 6.305572, 4.322502, 1.37244, 0.4938816, 2.232822, 6.728917, 
    3.513563, 2.310299, -0.1696083, 0.5774165, 0.8316671, 0.7628711, 
    2.716136, 3.166397,
  10.15029, 6.882953, 3.916265, 2.202524, -0.3775803, 2.123917, 1.172223, 
    0.1699456, 0.1096677, 0.4884017, 0.2179096, 0.5167186, 0.5133069, 
    0.9974283, 2.193728,
  32.30763, 8.938284, 4.997713, 3.744852, 2.790122, 2.523584, 0.8112922, 
    0.4831456, 0.7020801, 0.6576236, 0.6626107, 0.6423431, 1.031002, 
    0.7739263, 1.23676,
  61.75907, 62.84497, 57.62858, 16.16411, 4.974273, 3.053246, -1.258246, 
    1.622446, 2.007194, 1.833875, 2.215497, 1.755143, 1.460495, 1.364617, 
    0.2636522,
  75.89421, 64.36103, 63.16822, 13.20879, 3.478745, 3.635364, 1.148712, 
    -0.5745736, 0.1228955, 4.144567, 8.117682, 3.797458, 1.883925, 2.058336, 
    2.464998,
  86.72151, 65.62926, 41.11961, 14.62837, 6.465036, 0.06917249, 0.6121171, 
    -0.4347376, -0.7761884, -0.4424909, 1.169821, 3.514153, 3.192312, 
    3.01385, 2.162414,
  86.30855, 67.12823, 44.52944, 22.28353, 22.30773, 1.601747, 0.6238034, 
    1.403731, 1.563106, 1.124226, 1.707807, 2.929781, 3.860103, 3.299892, 
    2.565926,
  73.81803, 57.89239, 47.14967, 33.546, 27.23651, 4.136489, 2.854042, 
    2.883674, 3.079797, 2.047841, 1.743688, 3.00709, 2.941306, 2.300826, 
    2.7495,
  41.11039, 50.84583, 51.38219, 32.77885, 11.30726, 4.892712, 4.407865, 
    6.478714, 10.13997, 9.852685, 2.731486, 2.267623, 2.943807, 2.964318, 
    1.881067,
  43.9267, 43.85178, 33.46407, 13.50219, 6.12682, 4.515655, 5.150437, 
    17.63333, 20.0165, 5.965184, 3.730931, 0.5237694, 0.5839024, 2.784193, 
    1.476701,
  4.716744, 5.15873, 5.023942, 3.104895, 0.8585042, 1.295869, 1.875245, 
    0.1399084, 0.7526517, -0.8215626, 1.085841, 1.784386, -0.1293641, 
    -0.3273894, -1.772853,
  7.652506, 4.632188, 4.495714, 2.033956, 0.1771537, 2.586056, 2.002676, 
    0.438918, 0.3748494, 0.1798149, 0.239587, 1.287245, 0.4279779, -1.470806, 
    -1.374268,
  24.22955, 7.904748, 3.989346, 4.262218, 4.585125, -0.4632673, 2.7005, 
    2.266011, 0.3769006, 1.114024, 1.930316, 2.288854, 1.470774, 0.7912278, 
    0.9378165,
  46.94034, 50.07157, 49.91345, 22.43657, 7.497532, 9.0791, -0.6240214, 
    2.261029, 1.873767, 1.978017, 2.959969, 2.696462, 1.85055, 1.157654, 
    1.458593,
  62.23387, 50.99144, 59.05331, 28.79849, 6.445056, 9.406315, 6.402256, 
    -1.937499, -0.1424298, 2.633765, 6.570449, 3.040801, 1.246931, 1.897202, 
    2.38096,
  73.37996, 54.73251, 45.51503, 26.72418, 12.63119, 4.181505, 5.687135, 
    4.26251, 4.134654, 0.6237935, 0.7576794, 1.810121, 1.116924, 1.523118, 
    1.754822,
  75.60751, 63.11632, 50.83038, 31.43295, 32.04863, 3.669123, 1.02432, 
    2.205846, 1.615041, 1.394648, 0.8756307, 0.6465906, 2.20112, 2.300049, 
    1.341564,
  69.10398, 58.81414, 48.24575, 38.92723, 38.5776, 3.467721, 1.056533, 
    1.180803, 1.374444, 1.430549, 1.287225, 2.959297, 2.857121, 1.89502, 
    2.679203,
  53.11034, 50.70695, 49.35711, 33.62244, 7.25505, 3.367058, 3.898704, 
    4.408228, 5.396223, 4.584219, 2.288461, 2.147559, 2.836077, 2.42025, 
    2.14142,
  44.85237, 25.95175, 12.12912, 4.15855, 3.569469, 5.166556, 6.632286, 
    12.37117, 13.51073, 3.3563, 2.059081, 1.16374, 0.6117242, 2.053012, 
    2.510128,
  6.97179, 8.473328, 8.260953, 5.159526, 1.460864, 0.6100988, 0.8795227, 
    1.771169, 2.005049, 1.585453, 2.990865, 6.755682, 4.187778, 4.967916, 
    3.692251,
  8.316617, 6.118778, 5.469402, 2.414379, 0.6564699, 1.927669, -0.005417849, 
    0.3062019, 1.475075, 3.128104, 4.676201, 7.802202, 6.978359, 2.775382, 
    1.695737,
  22.8042, 3.610071, 3.28747, 4.549757, 4.110651, 1.535806, 1.409869, 
    0.4414407, 1.460404, 1.504868, 2.043373, 1.789398, 2.789864, 3.577061, 
    1.901496,
  35.06679, 34.22791, 28.98119, 11.14366, 7.434839, 6.978791, 0.7153062, 
    2.297671, 2.45806, 1.975387, 1.675732, 0.898307, 1.349121, 0.9254077, 
    1.78077,
  41.42165, 36.4784, 31.88983, 16.23014, 5.469238, 7.300159, 7.673354, 
    -1.930296, 0.2869052, 1.649423, 4.871013, 2.460362, 0.5047768, 0.4857584, 
    0.951097,
  45.69893, 37.05814, 27.4302, 20.39886, 11.64172, 4.725463, 4.656454, 
    2.833184, 0.4889927, -0.317599, -0.2745006, 0.2992582, -0.2118175, 
    0.2882505, 0.002054538,
  57.77436, 46.85925, 40.49239, 30.85232, 32.06718, 8.104975, 2.837595, 
    1.354684, 0.1502484, 0.3110676, 0.1542378, -0.3374955, 0.0561825, 
    0.1999422, 0.5067286,
  78.8204, 68.29929, 58.79893, 52.65309, 53.32987, 10.42849, 4.308452, 
    3.116583, 0.6559739, 0.01720612, -0.4419246, 0.4286579, 1.429446, 
    1.589608, 1.515105,
  98.53683, 89.17432, 79.13008, 58.35683, 22.4869, 10.74093, 8.84655, 
    8.79024, 7.067042, 5.513819, 1.862811, 1.502138, 2.039402, 1.027941, 
    0.6656837,
  110.308, 91.95644, 61.11036, 19.84615, 12.55558, 11.50317, 9.01223, 
    18.86876, 11.08036, 1.67197, 0.4682118, 0.1905358, 0.3666477, 0.6135273, 
    0.6356544,
  4.160027, 4.586697, 9.274728, 6.514206, 2.463774, 2.553691, 7.729863, 
    8.158063, 8.617881, 6.990738, 5.269188, 7.040046, 3.040633, 2.628419, 
    2.057083,
  5.9206, 7.300184, 7.599895, 1.958245, 0.1929478, 4.213069, 3.194656, 
    0.5248065, 5.277707, 6.823534, 8.679059, 8.500693, 7.858272, 1.363165, 
    0.6219943,
  34.10173, 12.72907, 8.381871, 6.48763, 4.394839, 2.839454, 4.089733, 
    3.230683, 0.9589726, 2.077628, 2.419225, 0.2166737, 0.780066, 0.7741818, 
    1.293822,
  67.16784, 68.35654, 60.66537, 25.75596, 9.567767, 4.60991, 0.568832, 
    2.690186, 1.635064, 1.279318, 0.1596563, 1.001941, 1.102104, 2.173998, 
    2.032252,
  87.58175, 78.82859, 84.49123, 35.95831, 13.20619, 10.95598, 6.161593, 
    0.5783809, 0.919099, 1.735943, 3.440017, 2.176421, 1.561654, 1.761667, 
    2.764574,
  105.3115, 91.21653, 80.16167, 43.32114, 20.22636, 12.52642, 9.941882, 
    6.54377, 4.744534, 3.474154, 1.999701, 2.883343, 3.101236, 3.236555, 
    2.882727,
  117.1913, 109.4801, 96.55862, 59.02219, 48.62256, 13.11574, 10.5133, 
    10.27842, 9.769902, 8.219139, 6.374357, 5.451779, 5.492411, 4.931026, 
    5.349729,
  120.2549, 114.2906, 102.5718, 93.68229, 77.98672, 14.50444, 11.30259, 
    9.434158, 9.124426, 6.689562, 5.285571, 6.235288, 6.103418, 6.042924, 
    5.719238,
  115.2013, 108.8004, 98.85052, 71.91947, 24.57799, 10.55879, 8.438096, 
    8.537345, 6.769842, 3.087331, 0.5262995, 0.9149148, 1.40213, 1.214355, 
    1.253802,
  95.14699, 86.03129, 53.80653, 12.32921, 6.228151, 5.001123, 4.649474, 
    13.61299, 6.894752, 0.6524461, -0.01138695, -0.3360703, -0.239038, 
    0.02891872, 0.3933912,
  1.087937, 0.5502371, 2.494855, 2.709439, 2.88655, 7.075269, 10.79565, 
    6.303271, 4.697691, 7.727278, 7.229247, 8.51133, 5.3558, 4.655726, 
    4.367366,
  1.186525, 0.7194525, 0.1631539, 0.4477427, 0.7069143, 8.748765, 9.388798, 
    4.212044, 1.042505, 1.353114, 4.371141, 6.715565, 5.072834, 2.170435, 
    1.075122,
  38.68798, 6.668305, 0.7481418, 0.4266492, 0.9455038, 3.376653, 9.760843, 
    5.682912, 3.906456, 3.023446, 3.736398, 4.975507, 2.466371, 1.833511, 
    0.4495694,
  77.21099, 70.94633, 52.10038, 13.55392, 2.98498, 4.146758, 0.8062451, 
    5.267113, 8.747134, 6.261388, 5.449243, 4.593559, 3.762469, 2.788573, 
    1.105057,
  93.76833, 73.91801, 67.0296, 18.49985, 6.222656, 8.15122, 7.78415, 
    0.3124375, 2.524092, 6.572063, 9.203359, 6.60309, 4.984631, 4.334185, 
    3.385242,
  93.72858, 74.17405, 53.06562, 21.11496, 9.845778, 6.875267, 7.535035, 
    6.788743, 5.722797, 5.614832, 4.187018, 6.670662, 6.715157, 7.412227, 
    6.69558,
  88.13131, 76.49547, 56.48246, 24.27653, 30.01388, 6.949121, 5.279763, 
    6.847844, 6.216441, 5.898899, 4.434446, 4.433773, 5.739051, 6.188897, 
    7.376545,
  74.07816, 58.66056, 42.25734, 66.39984, 57.41656, 6.07821, 4.263055, 
    4.46616, 3.709394, 2.858965, 2.047588, 2.513915, 2.471574, 3.620574, 
    5.566427,
  67.51485, 65.70714, 84.43806, 81.95083, 20.57637, 4.356122, 2.942687, 
    3.10084, 3.847634, 3.172922, 1.464911, 1.603256, 1.19395, 1.342769, 
    3.461938,
  82.10021, 78.16814, 65.34999, 21.83143, 5.399924, 3.125486, 3.221883, 
    9.057036, 6.59949, 1.109305, 0.6091262, 0.334787, 0.008506588, 0.3605321, 
    1.632255,
  1.322678, 2.123792, 4.164842, 1.45896, 0.1275659, 1.275448, 3.170033, 
    0.2886815, 0.3526458, -0.5833734, -0.02441043, 1.19933, 0.6495506, 
    2.139575, 4.482076,
  2.004382, 1.065488, 0.82715, 1.055127, 0.1638094, 3.297366, 2.101003, 
    1.19283, 1.016736, -0.8883684, -0.2899148, 2.267725, 1.556001, 1.672394, 
    2.486608,
  20.76229, 6.926438, 1.915214, 0.9570093, -0.9160673, -0.5248804, 2.632175, 
    2.391387, 0.7001362, 0.7465469, 2.368631, 2.968931, 2.688945, 1.759952, 
    1.281275,
  52.56932, 46.48169, 35.14451, 10.84596, 0.008860965, 1.114074, 1.039699, 
    1.745105, 4.272821, 4.754217, 4.791212, 3.457026, 2.749883, 1.821966, 
    0.2042372,
  57.83919, 50.79058, 55.99577, 19.45569, 3.152509, 5.920071, 5.189651, 
    1.926142, 2.1653, 3.2871, 5.228909, 3.670093, 3.08927, 2.001475, 1.291043,
  61.54322, 58.44996, 56.14491, 29.19585, 14.9017, 10.02247, 9.925682, 
    7.393608, 3.434526, 2.151645, 2.227674, 3.555789, 3.3797, 3.006686, 
    2.56038,
  113.4034, 115.3435, 112.5219, 55.87261, 40.82108, 16.86116, 9.284957, 
    5.330311, 2.749285, 2.105038, 2.292758, 2.582649, 2.464363, 2.92193, 
    3.576437,
  156.6646, 149.8633, 134.1249, 116.2657, 61.83635, 11.46171, 6.065669, 
    3.593014, 2.851645, 2.393826, 1.940459, 2.080788, 1.718402, 2.610148, 
    4.372986,
  163.4815, 149.9184, 129.3388, 80.72134, 20.38715, 6.987159, 4.35626, 
    3.694618, 3.95719, 2.878648, 1.718822, 1.66307, 1.781418, 2.466476, 
    4.158681,
  125.4008, 112.473, 69.33456, 14.86604, 5.665285, 3.968363, 3.669911, 
    11.19304, 7.143874, 1.125681, 1.848114, 1.51351, 0.8254482, 1.380596, 
    2.654655,
  5.184154, 10.4012, 10.77939, 9.504035, 7.414597, 2.779443, 2.981009, 
    2.123757, 4.128672, 3.467206, 5.337275, 10.59754, 4.972414, 3.905413, 
    1.762937,
  7.894533, 8.907721, 10.39915, 13.3287, 14.8465, 6.441638, 3.543865, 
    2.539921, 3.764867, 6.645877, 4.420756, 7.599854, 6.510765, 2.572308, 
    1.181229,
  37.23787, 15.28241, 11.211, 11.98707, 13.49964, 3.548388, 5.228603, 
    3.852262, 2.266169, 4.876801, 5.858673, 3.640619, 3.482469, 4.444963, 
    2.321303,
  57.7307, 65.20927, 61.71103, 23.10632, 9.518402, 10.15612, 4.798563, 
    7.395302, 6.540289, 5.315745, 3.676048, 1.688911, 1.328981, 0.9034364, 
    -0.45923,
  68.54419, 64.70197, 74.61343, 29.72099, 6.875449, 9.50428, 15.07704, 
    3.985679, 2.78906, 2.125562, 3.616982, 2.045898, 0.8453902, 0.618242, 
    0.06585244,
  89.91651, 84.39545, 78.36874, 33.69728, 16.89509, 8.43806, 5.777116, 
    8.467237, 3.862755, 1.954482, 1.080285, 1.574874, 1.091559, 0.857919, 
    0.5204855,
  87.26546, 85.96262, 74.09392, 28.8024, 18.84216, 9.258579, 6.515335, 
    3.654363, 1.977989, 1.90059, 1.248518, 1.052168, 1.68168, 1.940245, 
    1.727611,
  71.01513, 66.08773, 56.71876, 44.078, 20.69141, 4.428043, 2.994734, 
    2.452662, 2.055293, 1.857108, 1.264445, 1.397522, 2.086542, 3.055534, 
    3.587206,
  75.5746, 69.63298, 63.84282, 42.48516, 8.238497, 3.532988, 2.650404, 
    2.459729, 2.599751, 3.948255, 3.874433, 1.754641, 1.297025, 2.39574, 
    2.31244,
  79.90501, 73.75326, 51.54237, 7.170615, 2.753691, 2.272519, 1.244608, 
    3.555784, 3.171737, 1.601562, 5.797743, 1.697822, 0.2161006, 1.504457, 
    1.338078,
  5.851404, 13.20418, 16.44506, 15.28454, 14.6142, 3.842422, 4.016097, 
    5.644266, 6.84875, 6.248717, 7.576801, 12.18638, 8.225635, 2.43858, 
    3.033328,
  9.915243, 13.24953, 14.95967, 30.32431, 22.57847, 4.938068, 1.045076, 
    2.117066, 4.871033, 7.795453, 6.738258, 9.12789, 6.512569, 2.008884, 
    1.710109,
  53.41221, 28.18104, 23.4825, 33.03344, 23.83605, 3.751148, 1.007419, 
    1.261094, 5.000661, 8.00227, 7.346055, 4.552041, 4.584992, 8.037123, 
    7.970729,
  71.89898, 88.29851, 91.24792, 39.72113, 28.10325, 16.43694, 2.760245, 
    1.764783, 2.888948, 3.06766, 4.569711, 1.738808, 2.891261, 3.211987, 
    7.824443,
  70.21291, 72.31601, 89.29205, 32.82484, 23.36751, 24.63191, 17.59468, 
    3.179342, -0.2781606, 0.7787404, 2.686516, 0.860285, 1.071338, 1.739503, 
    4.169616,
  65.64422, 57.68931, 52.61151, 18.61243, 18.2989, 20.36704, 20.97094, 
    14.21741, 5.968769, 2.898597, 1.31937, 0.880502, 1.426054, 0.9842529, 
    1.865098,
  76.19357, 59.34848, 40.23378, 11.54833, 13.58963, 14.43704, 13.95962, 
    12.59019, 8.639886, 6.38184, 2.492861, 1.307615, 0.6327702, 1.427597, 
    1.457496,
  92.66783, 80.41936, 60.19171, 32.58891, 17.2213, 5.543457, 5.75283, 
    7.59988, 6.143927, 5.305562, 3.598323, 2.052817, 1.00524, 1.800457, 
    2.500075,
  101.7919, 96.35878, 82.41, 46.24577, 13.48097, 6.551675, 3.274623, 
    3.040076, 4.224718, 3.941929, 3.068573, 2.313309, 2.020118, 2.091336, 
    2.545387,
  43.8055, 32.34571, 21.28072, 10.35725, 6.668612, 8.396729, 3.748792, 
    1.919505, 1.570578, 0.6406033, 3.366325, 2.187899, 1.864318, 2.50037, 
    2.031224,
  1.531133, 1.078259, 2.166166, 5.020624, 24.80695, 10.7894, 1.730217, 2.646, 
    3.578845, 8.81739, 12.06463, 11.94094, 9.388659, 5.345649, 3.855946,
  4.27143, 1.388392, 0.7295358, 10.44947, 16.83053, 6.329895, 2.575503, 
    3.221339, 2.417585, 9.235346, 11.00083, 12.76283, 6.618962, 3.8243, 
    1.709981,
  26.33061, 7.19471, 3.86634, 10.91765, 10.74065, 4.377716, 2.980933, 
    2.326699, 4.81414, 6.522428, 8.287464, 6.203538, 6.112091, 6.437729, 
    5.59505,
  43.12186, 38.46487, 39.32754, 10.57838, 12.69277, 7.998024, 4.695981, 
    5.230376, 3.96837, 4.190134, 3.597017, 1.417874, 3.909355, 6.143681, 
    5.734393,
  59.8429, 37.107, 36.77884, 5.175008, 9.876561, 12.51432, 3.893995, 
    4.322541, 2.673418, 0.5866979, 1.57855, -0.3351623, 2.769705, 3.489688, 
    6.016744,
  78.05318, 51.55544, 26.15628, 2.517675, 7.235917, 10.72631, 4.998803, 
    2.171864, 1.87915, -0.5414635, -0.8197181, 2.417581, 3.076067, 2.113792, 
    4.155154,
  94.60332, 74.64199, 43.17618, 7.033528, 3.389569, 8.188538, 6.419537, 
    1.097793, -0.4420864, -0.1226995, -1.412983, 2.751209, 3.276476, 
    4.453021, 5.794816,
  111.61, 94.80289, 64.3786, 27.8003, 5.338083, 4.460488, 4.417305, 1.829085, 
    -2.195684, -1.939556, -1.044423, 3.510343, 3.380529, 5.304296, 7.525681,
  127.5346, 107.7408, 79.80571, 30.31748, 7.05999, 8.330577, 2.790274, 
    2.4511, 0.5983832, -2.34073, -0.169365, 3.622088, 3.47604, 5.041762, 
    6.43079,
  129.3702, 115.8463, 69.93726, 18.05674, 3.920355, 6.157795, 4.409606, 
    1.657547, 1.06208, -1.023567, -0.6063229, 3.086423, 2.970793, 5.792549, 
    8.417458,
  5.392992, 7.10312, 3.074578, 6.214971, 2.285697, 0.7410472, 1.285361, 
    2.60697, 4.831236, 8.151539, 3.879118, 4.88413, 3.487341, 2.410195, 
    -0.5805813,
  16.40239, 14.25385, 9.361386, 3.60464, 2.660492, 1.492021, 0.7564152, 
    2.965994, 6.046965, 1.662202, 5.078314, 6.192488, 10.1504, 8.287816, 
    -1.121171,
  75.39969, 38.81816, 16.89114, 9.479999, 1.251772, 0.05498458, 0.7237055, 
    0.7998354, 3.286242, 3.496372, 7.28543, 8.154481, 8.127668, 7.254055, 
    5.121826,
  109.8681, 109.6727, 86.02099, 22.42844, 2.689581, 0.5020962, 1.36329, 
    0.7382814, 3.995782, 4.450266, 4.393402, 5.498856, 8.504573, 10.00264, 
    11.47569,
  128.6496, 123.0953, 105.4701, 20.2325, 5.288925, 1.298015, 3.098219, 
    2.579057, 1.46534, 0.6694022, 4.930083, 8.026071, 10.80359, 11.30696, 
    10.86942,
  142.7725, 139.6605, 103.2128, 24.29509, 11.86294, 2.435861, 1.693551, 
    2.382753, 1.892304, 4.232513, -0.2543254, 9.596797, 8.925919, 5.861864, 
    5.736435,
  157.9521, 160.6952, 126.0356, 42.38845, 19.77561, 2.359786, 4.907101, 
    0.7287047, 0.6247162, 6.913689, 3.392831, 5.928944, 5.185967, 6.135111, 
    6.657076,
  169.3437, 174.4378, 143.0173, 100.4274, 33.80375, 1.967181, 1.524508, 
    2.982308, 1.696904, 5.742179, 3.20001, 4.504247, 4.467327, 7.426926, 
    6.019959,
  171.3329, 178.3788, 156.0607, 103.286, 23.03964, 2.740684, 0.8060032, 
    1.635835, 3.783175, 3.993806, 3.11034, 5.055525, 5.987531, 6.888416, 
    5.986832,
  133.298, 124.805, 84.78484, 29.07913, 12.26606, 3.796831, 1.616182, 
    4.667257, 3.680499, 2.796976, 4.250107, 4.159015, 7.561662, 5.71216, 
    7.567675,
  1.544467, 2.087695, 1.32849, 1.990486, 11.02511, 6.896401, 4.661807, 
    8.029529, 12.41466, 10.12422, 9.766298, 7.847055, 9.061702, 11.53012, 
    6.224305,
  7.253767, 3.106004, 1.629433, 3.310472, 11.33531, 4.397444, 3.294017, 
    7.283557, 7.588115, 8.85457, 8.42948, 12.55433, 18.22574, 8.529901, 
    6.996657,
  73.92358, 34.90188, 9.547541, 3.981495, 3.716835, 4.643897, 2.063211, 
    3.504686, -0.1008381, 0.592003, 9.494267, 14.68769, 15.74755, 18.84682, 
    13.68632,
  97.96046, 92.98058, 76.07868, 14.85817, 2.838658, 3.0083, 3.339872, 
    0.4116389, 1.597472, 3.046897, 5.888569, 12.80221, 14.54755, 16.01468, 
    19.0575,
  109.6934, 94.53535, 81.31237, 11.15026, 1.824545, 1.924889, 3.845844, 
    -0.06600938, 1.267144, -0.1293221, 6.003521, 11.82702, 13.16989, 14.8366, 
    16.44559,
  117.7986, 101.7622, 69.66949, 15.64401, 8.895355, 2.968563, 3.800458, 
    6.664581, 3.526735, 8.460585, 2.337968, 12.6455, 12.127, 11.62063, 10.1331,
  119.2155, 112.9171, 87.46294, 35.36578, 13.49704, 2.915179, 2.969805, 
    2.592125, 3.43943, 5.837554, 10.77615, 13.05644, 11.37345, 7.166646, 
    5.22565,
  116.6421, 112.8864, 97.47898, 71.5264, 28.89347, 3.374111, 0.8891766, 
    3.347916, 1.117153, 9.091572, 8.846946, 7.513453, 6.523007, 4.105535, 
    3.021631,
  114.4991, 114.5759, 107.3089, 61.78621, 16.22955, 4.262167, 0.2021916, 
    -0.1026734, 9.336631, 7.213042, 4.49162, 5.055476, 3.388853, 2.729587, 
    3.655685,
  82.12142, 75.05859, 47.63642, 18.78416, 7.271586, 1.327584, 0.2344884, 
    1.018197, 8.299723, 6.774635, 4.337028, 2.243717, 2.545465, 1.809838, 
    4.428433,
  1.07215, 2.990634, 1.643653, 7.7667, 8.169886, 6.258756, 3.197139, 
    9.110783, 9.626805, 6.879174, 6.76707, 11.39769, 8.728559, 8.742643, 
    4.955742,
  4.110196, 1.247227, 1.961161, 8.804523, 9.093617, 2.198006, 2.013281, 
    9.116291, 5.915938, 10.05828, 5.349485, 16.21955, 22.26495, 9.341016, 
    5.438158,
  36.02866, 18.79485, 12.02032, 14.75469, 6.502272, 5.919912, 0.9768114, 
    7.935176, 6.313883, 8.667553, 9.72227, 14.64304, 21.83322, 26.66927, 
    17.70331,
  45.14111, 49.39048, 55.53159, 23.70643, 12.93986, 6.588696, 2.840415, 
    3.640269, 6.120068, 6.319683, 5.342984, 6.809323, 10.93035, 15.52055, 
    23.76548,
  47.79293, 46.02852, 48.23108, 15.38804, 13.18086, 13.74103, 8.534646, 
    1.856274, 1.773016, 3.120964, 4.861354, 3.730255, 6.069005, 7.737846, 
    14.33922,
  50.56912, 45.96446, 36.19939, 16.73396, 15.80511, 15.12319, 16.65932, 
    14.95581, 8.730628, 11.68512, 4.08628, 3.679972, 2.718155, 2.787049, 
    6.132087,
  49.64563, 52.65963, 44.10058, 23.52427, 14.17659, 11.95562, 8.036961, 
    7.536204, 9.145402, 7.958412, 4.912844, 3.292777, 2.619113, 1.997356, 
    2.741044,
  48.1285, 52.27493, 51.41608, 39.34318, 21.06142, 8.852675, 4.766313, 
    4.077987, 3.093341, 3.345087, 2.499325, 2.119914, 1.821534, 1.52589, 
    1.657996,
  47.48716, 50.92958, 52.9671, 30.95028, 15.0258, 7.29037, 3.143961, 
    2.106585, 1.534937, 1.016678, 0.8408984, 1.342133, 1.25219, 1.09655, 
    2.609094,
  33.85039, 29.9387, 20.98465, 11.25379, 10.6791, 8.723095, 2.780656, 
    1.73596, 0.6826808, 0.255316, 0.9457123, 1.00047, 0.9248466, 0.7307764, 
    3.887084,
  5.430496, 2.656425, 2.934492, 2.695522, 3.112795, 2.109907, 1.685515, 
    1.715166, 2.946063, 4.160662, 4.238678, 10.7377, 8.029756, 7.926235, 
    4.019492,
  3.208178, 3.268411, 2.484337, 3.205456, 7.636982, 2.74253, 2.698115, 
    2.278799, 2.954989, 5.987885, 4.638035, 7.836297, 13.70111, 7.139671, 
    4.706598,
  4.990718, 4.701018, 3.815387, 6.47988, 5.666598, 3.025068, 5.159425, 
    3.706108, 3.554162, 3.260877, 3.712324, 6.990311, 12.40148, 13.75058, 
    10.27984,
  7.863513, 18.18764, 25.5132, 9.857221, 7.511977, 6.22355, 3.293742, 
    3.660969, 4.378118, 3.701264, 2.775709, 3.053614, 5.902493, 8.524112, 
    11.24262,
  13.30505, 18.37437, 31.0695, 8.039486, 10.20428, 11.68548, 12.25267, 
    2.740296, 1.357745, 3.55765, 4.567912, 2.160627, 2.568948, 3.682211, 
    9.063853,
  22.20489, 24.66743, 27.89694, 12.48334, 19.25469, 17.38879, 18.50911, 
    18.88975, 11.50199, 9.19774, 4.670687, 3.467453, 1.32446, 1.967883, 
    4.040304,
  31.58784, 39.56049, 46.98375, 37.04245, 26.27177, 15.67152, 15.39475, 
    13.25814, 10.20726, 9.1445, 4.841232, 3.749395, 1.388519, 0.9392329, 
    2.819039,
  46.5642, 55.68031, 61.67252, 64.57757, 47.12326, 13.92815, 11.61231, 
    11.82545, 7.803073, 5.54513, 4.493846, 3.639294, 1.547931, 0.4637979, 
    1.151181,
  58.32315, 67.52096, 76.63924, 42.01188, 23.76044, 13.07598, 9.76196, 
    10.96766, 7.270822, 3.862808, 3.336233, 4.453131, 1.988994, 0.6188375, 
    1.721694,
  48.21098, 49.0313, 39.4785, 18.44148, 15.84967, 11.45533, 9.458151, 
    12.76051, 9.34308, 2.334214, 5.389732, 5.117229, 1.328113, 0.7526156, 
    2.008554,
  4.862671, 8.197927, 8.58928, 8.632913, 12.08425, 14.31383, 14.57296, 
    12.23147, 9.503485, 5.573126, 10.31037, 8.531377, 4.575723, 5.82917, 
    5.33141,
  11.38033, 10.68192, 9.115034, 11.9404, 16.68057, 12.49888, 15.31023, 
    15.16156, 7.696202, 6.596527, 7.246071, 8.8599, 10.04253, 5.111023, 
    5.021148,
  41.60959, 40.50496, 29.06922, 17.08721, 9.410078, 10.21932, 19.55936, 
    17.0442, 7.745421, 3.63822, 6.611332, 8.17079, 10.99574, 13.88164, 
    10.50342,
  58.53876, 72.51099, 89.79483, 36.72615, 12.03507, 10.16941, 5.069192, 
    18.241, 17.22429, 4.563772, 4.84123, 7.222148, 8.264648, 11.50543, 
    15.26337,
  67.08158, 69.72504, 88.20722, 27.65404, 20.45389, 16.30889, 10.45448, 
    2.649469, 11.67313, 11.11186, 3.917963, 4.208713, 7.509652, 11.57795, 
    15.65003,
  70.6562, 75.0041, 74.28895, 28.76848, 35.98701, 32.62075, 20.47143, 
    16.14425, 12.99373, 9.667359, 3.2873, 3.781112, 7.363853, 7.988725, 
    10.21926,
  68.70419, 82.03535, 85.90082, 65.95271, 39.69341, 20.98352, 22.25481, 
    17.77547, 11.06721, 6.039762, 4.676897, 4.187486, 5.133415, 4.950686, 
    4.3149,
  59.83649, 79.86295, 84.36034, 83.53894, 51.52629, 13.90021, 13.1248, 
    15.09265, 14.37841, 12.19771, 2.138852, 5.362439, 4.3734, 1.87194, 
    2.764188,
  48.5408, 67.2935, 73.29723, 35.15401, 18.22858, 9.227415, 9.812243, 
    11.63841, 15.65965, 12.82213, 7.385444, 5.095074, 2.496601, 0.9676537, 
    0.9942026,
  29.4277, 35.61985, 26.37409, 11.10352, 9.293483, 6.310747, 6.168753, 
    19.26593, 19.78505, 9.46373, 4.966846, 3.329596, 1.149862, 0.9561023, 
    1.940352,
  2.185654, 3.295396, 3.503964, 3.447723, 8.101805, 4.47787, 3.723436, 
    3.954555, 7.305046, 7.497001, 6.922509, 6.250088, 3.586005, 2.328387, 
    5.321836,
  2.535334, 4.690339, 2.062159, 4.701542, 9.383555, 3.859227, 5.933184, 
    7.64292, 9.889399, 9.015483, 2.448064, 6.291701, 3.657611, 2.823868, 
    0.7772301,
  16.21359, 15.59737, 10.4349, 4.798595, 2.941506, 2.35494, 11.35046, 
    9.898454, 10.92611, 8.492952, 7.42719, 5.097867, 6.785001, 9.631906, 
    3.802249,
  16.79363, 23.31626, 26.81675, 7.907197, 3.12273, 1.463861, 1.91976, 
    11.26478, 15.83474, 9.535234, 7.461492, 9.086025, 10.63216, 7.373973, 
    8.455014,
  16.04245, 13.17811, 17.91264, 2.595324, 2.914947, 3.576977, 3.357837, 
    -0.3103769, 6.462055, 10.98003, 7.07399, 4.837254, 8.406094, 9.962164, 
    11.3741,
  13.94076, 6.475413, 3.167701, 1.127657, 6.835409, 6.701187, 4.128849, 
    4.526775, 5.044464, 5.089999, 2.231476, 2.95228, 3.548718, 5.330081, 
    8.890325,
  11.70381, 6.611411, 3.073562, 1.799109, 4.011123, 3.124867, 3.117274, 
    3.200021, 3.287116, 3.974345, 4.042793, 4.008316, 3.17822, 3.697816, 
    5.091951,
  15.43057, 8.739462, 2.030895, 0.4710679, 4.360097, 2.315045, 1.774252, 
    2.601051, 2.788431, 3.340801, 3.454815, 2.963329, 2.495057, 1.896265, 
    2.028047,
  23.19872, 16.53645, 5.410735, 0.1140938, 3.086895, 2.917728, 2.303107, 
    3.000983, 3.760577, 3.600348, 2.684103, 2.853504, 1.971998, 1.785691, 
    1.902284,
  15.21884, 6.000307, 0.3392942, 0.3713567, 1.592116, 1.747717, 2.476525, 
    5.436633, 6.106544, 2.042729, 2.198955, 2.966434, 1.117558, 1.100083, 
    3.008123,
  4.507793, 6.86301, 5.147821, 2.755777, 2.012081, 2.085034, 2.11511, 
    1.05248, 1.35888, 0.5587899, 6.969561, 9.258104, 6.281995, 4.162966, 
    1.451036,
  6.183812, 9.754218, 4.660101, 1.411546, 1.346591, 1.002577, 0.7455794, 
    0.4631866, 0.7071003, 1.759782, 4.82418, 10.00292, 11.3067, 6.558167, 
    1.329319,
  9.002967, 9.986646, 7.057298, 3.002881, 1.117365, 3.979897, 1.080436, 
    1.18328, 0.373367, 1.495904, 3.998015, 6.983577, 10.54894, 15.09812, 
    12.20202,
  21.52468, 22.09698, 20.94165, 5.747143, 2.593776, 1.423217, 3.549464, 
    0.8651205, 1.338251, 1.622158, 1.708515, 4.704922, 8.80357, 12.14365, 
    12.63282,
  34.2441, 25.74604, 28.86388, 7.169082, 4.877475, 3.767886, 2.364406, 
    3.569916, 4.280862, 5.741333, 4.442442, 4.020899, 6.24017, 10.1717, 
    14.48308,
  46.60497, 35.63313, 24.53602, 9.387211, 10.76296, 6.795468, 4.529414, 
    3.77472, 3.826755, 3.277727, 1.628566, 1.571759, 2.386353, 7.233619, 
    11.85766,
  56.17752, 50.00061, 35.81004, 23.36695, 16.18975, 8.607845, 6.211532, 
    8.005191, 6.855396, 5.419368, 2.831987, 0.3003073, 2.171335, 5.573012, 
    8.835835,
  62.77597, 56.59643, 42.14393, 30.86049, 20.77591, 11.84206, 8.121896, 
    10.44164, 8.439621, 8.648725, 5.109609, 1.987559, 4.647085, 6.757268, 
    5.511618,
  61.25751, 55.19579, 44.65454, 20.03787, 13.46713, 10.47675, 9.943113, 
    10.45841, 11.98672, 11.83254, 6.711522, 6.034197, 6.319945, 5.124641, 
    2.979795,
  38.60883, 28.02277, 20.69193, 15.30311, 12.83812, 11.47574, 10.09606, 
    13.26868, 14.06204, 8.659932, 6.74556, 4.889194, 3.87467, 1.431709, 
    0.9504742,
  2.881394, 8.736198, 13.43569, 12.6596, 12.33491, 13.23385, 10.20724, 
    4.236462, 6.183592, 5.874156, 7.115574, 6.72578, 6.245918, 7.923496, 
    6.274902,
  0.8198931, 6.426811, 9.886168, 10.39687, 10.20473, 12.32701, 9.75843, 
    5.682397, 5.044305, 5.479272, 5.069458, 7.0643, 8.350929, 6.646269, 
    6.182791,
  -2.507138, 4.088897, 8.592834, 7.73794, 10.32536, 10.64919, 13.75608, 
    9.057183, 9.695284, 9.566417, 10.27078, 7.361718, 6.189159, 10.23969, 
    9.087637,
  -2.75457, 4.646664, 11.53543, 6.039237, 5.519374, 7.121274, 8.064709, 
    8.061245, 10.79648, 15.2914, 13.39247, 9.33596, 6.662205, 5.99086, 
    7.513615,
  -2.929192, -2.343942, 6.967244, 0.9934083, 4.533331, 6.634311, 5.525456, 
    3.982596, 9.795732, 16.60034, 16.47005, 12.16336, 8.337921, 7.250272, 
    8.35574,
  -2.674703, -4.619043, -1.920466, 0.5999869, 9.052237, 6.794258, 5.051827, 
    5.625656, 4.655973, 7.187147, 7.980967, 12.13842, 7.5142, 3.750374, 
    1.771577,
  -3.061074, -1.633921, -2.18662, 0.2911763, 5.815282, 5.542179, 4.532947, 
    5.206798, 4.623103, 6.654486, 11.03862, 10.55909, 10.10905, 4.123791, 
    4.929831,
  0.5909364, 1.360021, -2.063891, -0.9612098, 4.517266, 4.073059, 4.429997, 
    4.882267, 2.24817, 2.862254, 8.471854, 8.299404, 7.926065, 6.675158, 
    6.77227,
  2.667364, 3.077454, 0.6873364, -0.1018106, 2.107971, 3.532266, 4.412507, 
    4.522281, 4.14853, 2.698275, 2.340304, 3.827747, 4.251781, 2.496605, 
    3.103616,
  -3.747858, -3.367479, 0.351918, 5.691972, 5.256416, 4.494318, 4.856214, 
    6.826885, 7.932067, 3.406953, 1.241649, 1.352838, 0.9961576, 1.379219, 
    2.007988,
  -3.062284, 3.353079, 5.820369, 2.249537, 1.7512, 1.697058, 1.234061, 
    1.640337, 5.629883, 11.45099, 9.014266, 10.28798, 9.379801, 3.767337, 
    5.794563,
  -6.996556, 5.169112, 6.317901, 3.405718, 2.094221, 2.586413, 2.136274, 
    1.240597, 1.489426, 2.05731, 8.004048, 9.890061, 9.742509, 5.322901, 
    3.077203,
  -12.67662, 4.059248, 7.69, 6.23035, 2.564513, 4.095087, 1.526637, 1.506197, 
    1.656975, 1.688932, 6.641018, 10.26173, 9.034347, 8.164462, 4.693578,
  -7.615162, 9.710073, 18.90732, 9.88353, 3.875032, 2.061631, 3.018545, 
    2.55638, 3.490787, 5.451431, 6.933038, 5.974592, 7.394292, 7.607588, 
    5.950253,
  0.843915, 6.092087, 22.52425, 11.74532, 7.263287, 2.854669, 2.32328, 
    1.297651, 2.068781, 7.229664, 5.792607, 5.448836, 7.770357, 8.760791, 
    9.24736,
  10.2957, 7.489223, 17.5736, 15.85173, 13.22528, 6.197799, 2.980661, 
    2.775271, 2.047493, 1.933439, 3.072391, 4.21726, 6.752596, 6.585618, 
    7.795026,
  18.32187, 18.67555, 25.89332, 23.99622, 19.82565, 9.215453, 5.70759, 
    3.467103, 2.282207, 2.575821, 3.456251, 3.742357, 5.346025, 6.509552, 
    3.404184,
  25.07792, 27.68949, 31.06569, 26.19583, 23.35193, 11.23616, 7.515803, 
    6.586007, 4.008044, 3.600106, 4.156508, 4.69917, 4.614934, 4.569488, 
    4.157092,
  28.01575, 30.21822, 30.84817, 16.01024, 13.31253, 12.51225, 10.8592, 
    9.520554, 5.801706, 5.421232, 5.152856, 5.044979, 5.223949, 4.642862, 
    4.350308,
  10.54393, 13.52696, 15.72836, 13.51063, 13.98276, 14.80164, 12.34835, 
    11.75001, 10.47546, 5.174981, 6.349761, 7.258062, 4.472754, 4.705554, 
    3.795896,
  2.841259, 7.988783, 12.61235, 11.91574, 11.43779, 11.23471, 3.954237, 
    3.355638, 3.496151, 6.277546, 5.296018, 7.638427, 9.433766, 8.090599, 
    6.492411,
  -0.5011747, 4.787261, 7.07553, 13.34137, 14.58493, 11.48901, 5.382614, 
    2.185736, 2.93866, 3.967714, 7.305147, 9.568355, 8.786737, 6.231173, 
    5.591025,
  1.001657, 4.31248, 14.44714, 13.79311, 16.56147, 15.02635, 10.31158, 
    5.327566, 5.566949, 5.718362, 6.022138, 8.426184, 11.97222, 5.643385, 
    5.481119,
  14.25533, 17.56484, 28.98732, 18.2644, 15.42615, 14.90514, 11.49095, 
    6.39663, 7.996686, 9.378657, 6.857357, 7.421883, 7.754342, 11.8116, 
    12.07361,
  28.28499, 20.11082, 32.27657, 16.94417, 17.78864, 14.6152, 11.56737, 
    8.980584, 11.17022, 13.62265, 10.90449, 7.712538, 6.344635, 7.432448, 
    10.42294,
  44.15793, 30.13121, 30.89543, 26.356, 38.55605, 13.18669, 11.89317, 
    10.36036, 8.170752, 9.547725, 7.279684, 6.589468, 6.535543, 7.441706, 
    6.811846,
  51.08417, 47.21262, 42.67922, 49.30761, 43.31556, 15.62627, 11.1335, 
    8.743901, 8.399725, 7.662001, 7.593393, 9.251077, 7.019889, 6.717224, 
    5.740667,
  59.90534, 59.65398, 54.9374, 51.68674, 35.17572, 14.02525, 9.565447, 
    8.586807, 7.819817, 7.586133, 8.178695, 9.454895, 9.716278, 7.132096, 
    7.328769,
  63.36945, 62.48767, 56.38887, 27.99783, 13.44679, 14.58315, 10.22829, 
    7.818739, 5.936183, 9.027888, 7.385133, 6.929204, 8.446905, 8.763441, 
    7.906971,
  46.8642, 32.94846, 29.3222, 19.26842, 14.41926, 11.5478, 7.701475, 
    14.13682, 13.04054, 5.166982, 3.431246, 4.492945, 5.804305, 7.169309, 
    8.65891,
  7.561979, 10.5785, 13.28607, 11.64753, 10.46158, 11.52289, 9.134056, 
    9.952115, 12.59728, 11.25796, 8.60621, 9.65609, 6.906155, 6.555454, 
    9.266559,
  31.70922, 21.2114, 12.70707, 10.33565, 10.85297, 7.402137, 7.850227, 
    10.77799, 13.5136, 13.84005, 10.01937, 12.13943, 9.417019, 5.420595, 
    9.180529,
  58.03568, 63.27522, 59.16276, 17.20509, 9.74855, 7.767203, 9.950963, 
    7.718219, 9.766683, 10.85283, 10.86824, 12.03679, 10.71041, 12.27326, 
    9.200017,
  70.13158, 76.88829, 79.14274, 20.68784, 7.598713, 6.37426, 3.715374, 
    8.096236, 11.76392, 12.3782, 10.11965, 11.81794, 13.01873, 11.67558, 
    10.76891,
  78.27828, 73.89172, 75.84969, 19.36727, 11.62658, 5.957719, 4.26986, 
    0.6353078, 6.614648, 15.44417, 13.1053, 8.859039, 9.612075, 11.34647, 
    12.31619,
  91.64589, 79.86754, 70.33263, 35.29053, 36.37516, 5.975729, 3.241467, 
    2.433869, 1.491402, 0.9844564, 2.1818, 4.131538, 6.811574, 10.20574, 
    11.19817,
  102.5043, 95.06926, 80.0368, 61.58727, 38.79556, 8.160635, 3.733692, 
    2.576974, 2.051522, 1.160601, 1.800364, 3.122813, 5.982359, 6.933913, 
    11.39157,
  114.1472, 106.0601, 90.61613, 58.39238, 34.54935, 10.16875, 5.524529, 
    4.379939, 3.899431, 2.427327, 2.323598, 2.971032, 4.24797, 5.293612, 
    9.727464,
  118.0147, 108.3176, 83.57051, 24.74678, 13.55949, 13.12133, 7.615272, 
    7.49595, 7.194677, 7.253037, 3.059306, 2.738317, 3.197109, 4.341107, 
    9.875411,
  88.63766, 59.51375, 43.83028, 15.87599, 10.78613, 13.62701, 10.02984, 
    18.07822, 16.19599, 4.789424, 1.72684, 1.453826, 1.82144, 2.932528, 
    6.300864,
  5.499453, 8.726829, 11.54674, 6.127238, 3.928906, 4.506772, 5.66159, 
    1.990898, 2.296442, 4.441831, 3.684679, 3.467187, 8.881363, 9.685594, 
    7.818371,
  33.29337, 21.55747, 13.07979, 4.755254, 3.246158, 5.414366, 4.099549, 
    2.256679, 2.337595, 3.713462, 2.648931, 3.046508, 4.39339, 5.006205, 
    4.254564,
  73.52367, 69.5163, 52.02278, 8.174847, 4.396859, 5.46748, 6.473722, 
    3.562288, 3.978452, 2.499206, 2.927315, 3.366009, 4.760866, 7.460059, 
    7.616699,
  99.685, 93.60006, 78.23587, 15.73284, 4.317244, 4.150824, 4.9333, 6.062065, 
    5.400423, 4.005831, 3.150311, 3.066239, 4.414666, 5.036112, 7.827782,
  115.029, 96.04568, 80.35657, 11.24857, 5.606457, 4.875593, 3.792017, 
    2.112912, 3.996059, 6.946276, 5.684484, 2.411227, 2.601687, 3.46628, 
    5.5599,
  134.9387, 110.9101, 81.49118, 30.22821, 20.05102, 3.630234, 2.809151, 
    2.608998, 0.4755908, 0.05084966, 0.5149128, 1.406747, 1.875683, 2.69133, 
    4.520948,
  150.5311, 136.2547, 104.032, 59.00658, 27.34947, 3.947368, 2.35365, 
    3.066171, 2.422667, 0.7885829, 1.147089, 1.609577, 2.526404, 2.292016, 
    4.158794,
  163.8034, 155.2028, 126.0463, 64.17219, 28.94842, 7.735057, 5.647287, 
    4.924236, 4.472781, 2.783131, 0.9578558, 1.727751, 2.483281, 1.986893, 
    5.185342,
  164.5967, 158.1429, 111.8428, 34.26023, 15.99206, 9.695072, 7.936027, 
    7.678981, 5.782933, 3.809203, 0.7145897, 1.470772, 1.424672, 2.141333, 
    5.50455,
  119.8574, 81.21732, 62.75498, 29.99428, 15.64822, 11.81383, 8.434342, 
    10.96685, 8.972972, 3.335684, 0.4152024, 1.459174, 0.8876746, 1.762581, 
    4.070777,
  8.60025, 9.002213, 13.26919, 7.844097, 4.755306, 7.166138, 5.566926, 
    6.057733, 6.661591, 6.452715, 3.238002, 1.720872, 4.053388, 4.844605, 
    5.891252,
  67.86707, 38.19833, 16.56716, 9.71252, 6.589056, 6.004233, 4.706165, 
    5.328254, 7.033742, 8.069564, 2.326668, 1.741121, 4.040216, 3.863026, 
    3.176942,
  117.2004, 109.6122, 88.79044, 15.40432, 6.766704, 4.388942, 7.168262, 
    7.70879, 6.758944, 3.870188, 2.985892, 2.676258, 4.945501, 4.484684, 
    1.873682,
  142.3132, 133.6788, 114.1426, 22.56004, 10.41792, 8.70954, 7.255595, 
    8.33451, 5.597026, 4.702219, 3.294883, 2.684442, 4.450986, 3.708818, 
    1.872725,
  155.6479, 134.3035, 112.0644, 17.49621, 9.571495, 7.979961, 14.27761, 
    4.984465, 1.866744, 5.489538, 5.14563, 2.257222, 3.052085, 2.665544, 
    2.399437,
  172.1685, 147.0112, 114.355, 42.49898, 20.09212, 4.370454, 8.686808, 
    16.76372, 7.561567, 4.420062, 3.286273, 2.313531, 1.665398, 2.446575, 
    3.266085,
  181.7325, 171.2238, 138.2692, 69.76372, 26.83731, 4.804699, 5.898106, 
    8.533187, 5.9883, 4.65952, 6.295118, 4.062171, 1.996971, 2.205065, 
    3.264904,
  185.7123, 184.4846, 153.0569, 73.63882, 29.76643, 9.905721, 8.914259, 
    6.536284, 3.115416, 5.380068, 4.569646, 4.113071, 2.161377, 1.420222, 
    3.414776,
  168.1904, 170.7769, 108.3673, 40.01251, 21.79222, 11.69569, 8.725744, 
    4.077286, 1.606377, 2.88329, 2.466753, 2.807827, 1.429603, 1.310026, 
    3.721398,
  95.47284, 72.94338, 51.47762, 29.4625, 15.85362, 11.35995, 7.02543, 
    8.756062, 4.134668, 2.445299, 2.084527, 2.182917, 0.914324, 1.33028, 
    3.925075,
  7.328326, 6.121211, 6.258678, 4.14569, 8.44083, 7.36287, 6.388352, 
    4.957801, 5.8873, 10.02741, 10.7013, 11.65089, 6.978548, 5.871327, 
    2.195255,
  64.51016, 35.17912, 11.72988, 6.508191, 11.84584, 8.846544, 5.81873, 
    5.918783, 6.920636, 10.40532, 9.508422, 8.168675, 8.36772, 2.48082, 
    3.718155,
  92.19244, 85.49278, 74.31934, 13.71828, 13.1618, 8.381676, 5.594738, 
    5.640454, 6.5861, 7.1848, 5.800246, 6.677136, 5.944429, 4.83776, 4.323193,
  99.15993, 95.38464, 98.67122, 26.07488, 16.42313, 19.56247, 7.670455, 
    5.49078, 5.886168, 5.574191, 2.383614, 2.71489, 4.90526, 4.436031, 
    5.691648,
  96.84238, 84.1896, 87.08839, 19.29139, 17.05101, 18.92898, 22.55672, 
    4.145845, 1.698282, 6.00892, 3.743587, 0.2683751, 2.016763, 5.477644, 
    5.67562,
  104.3193, 83.16039, 77.58901, 40.57868, 28.05355, 13.09999, 12.46807, 
    14.36148, 5.294984, 3.660906, 1.280656, 1.364026, 3.379137, 6.695633, 
    5.605469,
  114.1502, 101.2488, 85.30779, 50.98479, 28.01057, 9.940554, 6.856648, 
    5.597165, 4.950172, 2.779768, 1.812234, 1.918743, 5.220222, 7.787095, 
    6.66967,
  117.3997, 112.5516, 86.30108, 47.51235, 26.19162, 10.90839, 5.942521, 
    4.129916, 2.712693, 1.784938, 1.690211, 1.968385, 3.622254, 5.19559, 
    9.082059,
  111.0101, 109.837, 59.70457, 26.80517, 15.31613, 11.09599, 5.852375, 
    3.46231, 2.644133, 3.167474, 1.901918, 2.408542, 2.48878, 3.193586, 
    6.821055,
  66.73417, 49.95588, 31.04224, 19.43809, 11.3269, 10.06573, 6.898151, 
    9.338926, 5.978864, 2.332226, 1.531443, 2.036895, 2.016988, 5.651986, 
    6.952555,
  3.849754, 3.053372, 3.368417, 4.43496, 12.77251, 9.358564, 9.222911, 
    7.890825, 7.486408, 9.266343, 9.691402, 8.267819, 8.458175, 18.87391, 
    18.59392,
  20.76486, 13.82237, 7.019867, 8.434639, 12.82601, 8.635664, 12.22927, 
    9.466063, 11.65254, 15.71316, 10.07443, 10.92097, 19.16342, 11.36895, 
    8.91898,
  42.65711, 50.04939, 52.33981, 13.53567, 9.586612, 4.667419, 12.68806, 
    10.74374, 9.145519, 10.9456, 10.65289, 10.94341, 11.10764, 13.95003, 
    10.32329,
  61.00829, 67.3985, 77.85639, 20.30095, 14.20687, 14.12382, 9.452978, 
    14.46397, 10.40348, 8.085188, 6.527815, 6.964655, 8.749253, 8.321346, 
    6.213634,
  76.78813, 68.89873, 70.39104, 15.27809, 15.06819, 16.9043, 16.25434, 
    5.120355, 3.247671, 8.482716, 6.101467, 2.536915, 3.287513, 5.05205, 
    4.917218,
  97.41567, 79.33905, 72.19421, 33.57134, 24.05188, 11.90638, 11.05343, 
    11.82318, 4.403016, 5.136017, 3.808249, 3.614318, 3.306119, 1.941941, 
    2.607238,
  107.6972, 100.8022, 87.21191, 48.68129, 24.21466, 11.52771, 6.003272, 
    5.977537, 5.228048, 3.320371, 3.331703, 3.901328, 4.801236, 1.231315, 
    4.099072,
  107.0322, 108.9426, 87.50924, 47.18524, 23.46497, 11.29878, 2.702665, 
    5.169593, 4.905815, 3.886457, 4.371002, 3.66636, 3.914898, 6.221284, 
    8.866199,
  98.62885, 100.9306, 54.26655, 26.34493, 14.96682, 7.465344, 4.245193, 
    1.408821, 5.934634, 6.291594, 5.967872, 6.099745, 6.711753, 6.920098, 
    10.19396,
  57.42607, 43.86367, 25.98228, 16.53937, 15.30319, 16.23314, 11.49034, 
    14.93497, 3.802915, 2.946954, 4.160329, 6.494595, 5.915293, 7.522305, 
    7.94818,
  3.566761, 3.87427, 6.728243, 5.884182, 11.05245, 6.228174, 4.078508, 
    4.754014, 10.99527, 14.93788, 15.14072, 9.84854, 9.935251, 8.126615, 
    5.342975,
  28.03857, 11.65374, 7.796602, 10.0162, 13.47486, 5.52739, 4.115419, 
    4.810824, 8.38905, 17.09109, 13.58242, 10.86041, 15.56294, 9.154056, 
    6.338931,
  58.5332, 55.39669, 42.85614, 13.6325, 7.230445, 3.736089, 5.74914, 
    4.312372, 5.545632, 7.618773, 11.12658, 12.63801, 11.15867, 16.77543, 
    12.71747,
  66.18395, 67.20757, 63.98086, 16.53939, 8.699865, 10.124, 4.891482, 
    4.73035, 5.824681, 5.090775, 10.11007, 14.25765, 10.18703, 16.50342, 
    13.99039,
  67.53646, 62.51812, 60.76432, 12.10354, 14.55731, 16.21155, 15.30424, 
    7.061203, 6.036041, 8.266672, 11.65677, 10.26785, 11.80804, 10.85785, 
    13.93024,
  69.55882, 63.89245, 57.57579, 31.86823, 25.61656, 17.44722, 15.2696, 
    16.04265, 9.419142, 7.125101, 7.474017, 8.31655, 9.063935, 8.446479, 
    12.84437,
  70.65202, 72.66086, 62.84706, 37.26368, 21.43703, 16.65172, 14.8164, 
    16.35596, 9.769937, 7.572482, 6.423601, 8.021536, 8.709203, 10.51668, 
    11.52664,
  74.16582, 74.19184, 52.44307, 26.60149, 17.67955, 13.44885, 12.60528, 
    17.53622, 11.57605, 9.172241, 6.974484, 7.661826, 8.279538, 10.03051, 
    10.73678,
  68.01365, 56.15356, 25.49244, 12.46337, 9.510063, 9.442392, 11.46624, 
    15.99475, 13.86963, 8.913006, 6.230647, 7.286419, 8.215082, 8.639404, 
    9.499717,
  32.20455, 15.61025, 8.682547, 5.573016, 4.497946, 9.186203, 11.05717, 
    23.65603, 15.7443, 7.12312, 5.087882, 5.407416, 7.064843, 8.747198, 
    8.840172,
  9.970611, 15.97986, 17.51085, 4.385594, 0.9970059, 4.325548, 3.107603, 
    2.032347, 5.267882, 9.965943, 13.97323, 8.908046, 9.19235, 6.557547, 
    7.066316,
  29.11652, 13.36007, 4.3255, 1.665688, 6.041646, 5.357241, 3.498793, 
    4.282879, 6.795442, 10.35239, 13.49434, 8.33042, 9.176368, 4.135893, 
    4.697537,
  37.30932, 23.22827, 12.4392, 1.585815, 2.135628, 4.641763, 5.221207, 
    7.08053, 8.442834, 9.808507, 11.78244, 10.43777, 4.370228, 8.813113, 
    6.874298,
  29.56773, 24.87879, 23.40627, 5.986911, 6.689305, 4.49867, 4.198097, 
    5.364468, 9.201216, 11.71253, 13.96566, 11.31124, 7.269896, 8.264771, 
    5.405505,
  22.67543, 15.00978, 22.58265, 7.902592, 7.89247, 2.474913, 5.510178, 
    2.717117, 6.745743, 10.27929, 14.13393, 12.68571, 9.546244, 5.622525, 
    6.044777,
  30.09735, 18.16458, 17.38119, 11.59653, 9.681346, 3.625762, 2.920346, 
    5.105989, 4.690075, 7.534822, 8.52477, 10.72006, 9.39475, 6.524132, 
    9.207852,
  35.67212, 27.95454, 20.84762, 11.45211, 8.737482, 6.922668, 2.856996, 
    5.575809, 7.813278, 9.525449, 11.11857, 10.30254, 9.661806, 10.24084, 
    9.97448,
  34.08242, 27.4998, 17.38562, 12.96506, 11.44707, 4.363573, 4.713223, 
    8.24171, 9.95227, 8.083672, 10.6563, 9.57123, 10.01743, 10.12555, 10.50456,
  26.2407, 21.23063, 10.38297, 10.04777, 6.707352, 3.454801, 7.498309, 
    8.925797, 13.01645, 10.27294, 10.10005, 9.627208, 9.024674, 7.508452, 
    8.535956,
  7.12417, 7.123618, 8.301513, 4.376601, 3.423824, 3.579875, 8.930795, 
    19.89916, 15.14746, 7.845837, 7.957963, 8.344316, 11.17095, 6.485116, 
    9.805947,
  4.890178, 8.36952, 12.25101, 4.404466, 4.805227, 6.757946, 3.615366, 
    4.885802, 4.071138, 4.657548, 4.659622, 8.102696, 6.025641, 3.018242, 
    4.286691,
  6.10418, 5.779694, 4.876995, 5.828803, 10.09137, 10.53902, 6.186901, 
    5.312587, 5.227722, 1.810453, 6.090585, 9.928888, 7.540864, 4.354355, 
    1.728018,
  8.058874, 12.18339, 16.50448, 7.853742, 10.86388, 12.63111, 7.486751, 
    7.017419, 1.773554, 1.341855, 7.576833, 10.17557, 9.298622, 12.2966, 
    6.234345,
  11.47497, 22.45592, 30.65296, 11.52489, 7.917209, 8.839954, 7.727059, 
    6.405945, 3.160053, 2.72777, 3.93838, 10.39328, 15.20809, 12.90866, 
    5.018439,
  16.35203, 20.68826, 31.11222, 10.96729, 8.962104, 6.490561, 7.811536, 
    2.143283, 1.190117, 4.329862, 13.3513, 11.6089, 16.27911, 9.995098, 
    8.596031,
  19.4981, 24.52841, 27.02635, 14.26941, 12.28788, 8.073498, 10.1888, 9.255, 
    6.516285, 3.382238, 11.08532, 5.065669, 12.74009, 9.552246, 5.617711,
  17.44376, 24.77666, 21.69642, 14.75412, 11.12673, 8.804317, 10.05119, 
    12.51957, 8.832857, 10.50788, 12.29448, 4.123833, 12.41881, 8.346192, 
    6.887335,
  13.66321, 22.36371, 15.51296, 10.27464, 9.232313, 5.676457, 11.11839, 
    13.55585, 11.28449, 11.85298, 11.72149, 4.245555, 8.233635, 7.572932, 
    7.787826,
  14.42036, 15.9506, 6.721179, 6.200553, 6.503844, 5.70474, 11.16311, 
    15.98806, 11.84591, 13.14684, 10.79438, 4.944166, 9.273602, 9.808477, 
    10.86709,
  3.276735, 1.300131, 4.04726, 4.088091, 6.14043, 5.985323, 11.47903, 
    26.80778, 17.93631, 9.876597, 8.484647, 9.605101, 13.4257, 14.77127, 
    5.850417,
  3.263049, 4.62766, 8.557801, 5.322009, 4.136843, 6.231505, 6.069133, 
    10.79311, 10.12722, 10.99804, 9.190219, 11.06909, 11.58208, 9.46937, 
    9.9856,
  10.7122, 6.94889, 6.631312, 4.659211, 4.93432, 5.118151, 4.079061, 
    3.729159, 8.09825, 9.252338, 9.260014, 11.63809, 10.74586, 8.566541, 
    10.70943,
  13.89577, 18.67985, 14.79441, 3.616826, 3.971192, 6.275032, 4.463066, 
    5.598712, 6.700251, 3.622124, 3.580835, 11.57271, 13.76377, 15.4212, 
    14.49975,
  11.65898, 15.28403, 17.03556, 4.571686, 6.506822, 8.073175, 6.038073, 
    4.706618, 7.430376, 7.902549, 8.769999, 11.77095, 14.37641, 16.36399, 
    13.08145,
  7.422705, 6.425015, 17.53628, 2.67354, 7.512209, 7.086072, 8.964714, 
    4.770696, 8.204809, 13.09609, 16.12298, 12.07735, 15.61726, 13.99909, 
    17.24846,
  4.267732, 4.141009, 13.62621, 6.382339, 8.841192, 5.329917, 7.329643, 
    9.655697, 7.466586, 8.459816, 10.4587, 9.630569, 15.48537, 15.95939, 
    17.73623,
  4.495773, 12.96701, 22.84259, 7.106149, 8.272775, 4.578414, 6.147465, 
    9.207762, 7.960179, 10.39544, 10.69793, 10.3051, 15.37848, 16.88128, 
    17.05769,
  7.116405, 19.92949, 28.24549, 9.618274, 8.002812, 5.688048, 6.476102, 
    9.385939, 8.694263, 13.11047, 11.88796, 16.73848, 18.7516, 17.94102, 
    13.8805,
  9.697922, 19.73104, 16.93647, 10.94364, 7.46316, 3.962421, 6.586277, 
    11.74572, 12.28942, 13.4284, 15.47745, 19.90262, 18.50677, 19.85263, 
    21.14141,
  1.341851, 6.854074, 10.13166, 11.05689, 6.71936, 5.485516, 6.659157, 
    20.04692, 17.23549, 12.56781, 12.94208, 16.06218, 20.23822, 19.05944, 
    24.94065,
  2.428061, 4.767389, 10.6884, 7.906828, 6.333433, 9.117081, 3.95745, 
    5.036367, 8.614313, 13.40126, 12.27934, 10.37899, 12.2328, 9.225894, 
    9.569738,
  3.034466, 5.313538, 10.20881, 9.030788, 15.48862, 10.68589, 5.767509, 
    1.793309, 1.38562, 3.815394, 8.264238, 11.54216, 11.43268, 11.39549, 
    10.41501,
  7.19802, 11.41099, 18.34055, 11.09625, 11.83496, 11.17417, 3.551114, 
    7.140288, 3.010844, 8.282678, 10.48815, 12.37123, 11.08025, 10.22067, 
    9.801101,
  7.515399, 16.82648, 27.56869, 13.50066, 9.374884, 8.506158, 5.108508, 
    6.464664, 9.559613, 11.43905, 12.64779, 12.54269, 11.74279, 12.11889, 
    15.72336,
  10.70897, 17.14866, 24.86811, 11.44863, 7.294089, 8.236723, 8.61191, 
    6.096262, 7.111052, 18.036, 19.72378, 9.27916, 9.596687, 8.932878, 
    11.07216,
  10.72721, 22.80102, 21.84391, 14.35432, 11.15508, 6.775081, 3.147584, 
    6.424003, 0.3839175, 3.3041, 7.908071, 12.64959, 13.06633, 8.092402, 
    9.405892,
  12.40565, 31.64401, 27.88708, 15.43688, 9.030682, 6.668097, 1.675905, 
    3.049578, 1.546535, 3.5642, 7.118373, 13.35764, 15.94882, 12.60602, 
    8.478079,
  16.99381, 39.33361, 29.44738, 15.49414, 6.824984, 5.639039, 0.9580542, 
    1.648452, 3.185537, 5.076983, 8.267848, 16.27735, 19.99493, 20.6433, 
    15.90463,
  16.31865, 38.12187, 18.61556, 7.728917, 8.345243, 2.666736, 0.6795259, 
    3.690876, 6.122715, 11.1991, 11.568, 12.88359, 20.67296, 21.19988, 
    29.27293,
  1.389845, 14.78848, 16.08811, 6.963767, 7.603142, 7.506783, 1.032212, 
    18.33889, 16.7644, 7.825875, 4.03207, 8.795056, 18.89489, 19.47961, 
    30.18831,
  3.102998, 4.357877, 12.7644, 2.107681, 1.859948, 3.242443, 1.459903, 
    1.226448, 1.420359, 6.588012, 5.943287, 1.519664, 10.12604, 12.94362, 
    11.00387,
  11.74495, 6.067078, 5.093845, 1.203454, 4.058632, 3.415967, 0.8944877, 
    1.19951, 1.259244, 1.497597, 0.5027329, 4.343766, 2.018905, 8.339373, 
    8.11013,
  20.09376, 22.0161, 18.33811, 3.022542, 2.493734, 3.009749, 1.724377, 
    1.316962, 0.9138656, 1.778133, 1.077303, 4.196865, 9.828581, 10.6759, 
    8.706294,
  16.73915, 21.23059, 22.33049, 9.91891, 2.853702, 1.993553, 1.981688, 
    3.271491, 3.797257, 4.654199, 3.55047, 8.383936, 11.04272, 13.99707, 
    10.62233,
  16.61185, 11.06449, 16.27404, 10.19516, 5.269343, 4.818093, 6.619477, 
    2.653608, 2.061328, 12.56912, 9.858357, 8.17476, 11.47461, 12.21679, 
    10.58492,
  13.4547, 8.536606, 8.668521, 10.30678, 11.96041, 9.126333, 7.777462, 
    4.99474, 2.3651, 3.441282, 5.186492, 8.457027, 15.39989, 12.07217, 
    11.39566,
  6.234204, 5.246871, 8.085712, 6.463365, 7.473558, 7.029294, 6.547052, 
    7.601271, 8.096537, 5.699979, 6.822537, 8.309536, 11.10545, 16.3121, 
    17.76647,
  5.763628, 6.172034, 6.663489, 5.686531, 7.903007, 7.871511, 8.995727, 
    8.099094, 6.505847, 6.726331, 7.77212, 6.68263, 9.05361, 21.17251, 
    26.46635,
  7.533319, 5.893977, 0.05037434, 1.250563, 3.722174, 5.708616, 7.461498, 
    7.255921, 6.767971, 9.023995, 7.535404, 8.391029, 11.13181, 18.99672, 
    37.7818,
  3.675863, -0.2037102, -1.195224, 1.214914, 2.370047, 5.148553, 5.35533, 
    10.53659, 12.72378, 8.372473, 4.431711, 6.134954, 5.296117, 15.70193, 
    29.29008,
  3.698663, 6.993743, 11.22246, 5.059876, 6.039533, 5.256106, 3.707842, 
    2.519738, 2.197643, 2.641068, 3.920362, 1.488369, 3.674355, 7.518199, 
    6.079666,
  4.928657, 4.673802, 4.462546, 4.170086, 5.288352, 6.272125, 1.57329, 
    5.051361, 3.770569, 0.5615773, 3.224133, 1.653801, 1.12792, 6.381642, 
    5.657463,
  4.168359, 3.374981, 6.108449, 5.047543, 6.721209, 9.914344, 8.024018, 
    6.000731, 4.738085, 2.966486, 2.792916, 2.185208, 3.241462, 7.88799, 
    7.455299,
  2.015721, 1.51993, 3.812742, 4.260083, 6.889945, 7.066133, 5.277748, 
    7.029979, 3.378168, 3.554039, 2.20457, 1.923734, 5.151281, 7.698529, 
    8.494789,
  1.814235, -0.2683868, 2.052361, 2.605045, 4.040477, 4.655022, 4.05384, 
    4.51477, 3.61763, 6.908442, 7.712345, 7.275168, 7.059041, 5.996127, 
    6.396163,
  3.236475, 0.7731532, -0.7810687, 1.438325, 3.636889, 4.261291, 3.504158, 
    3.166973, 5.435647, 7.116991, 6.517343, 6.249733, 7.280231, 5.491056, 
    5.008281,
  4.970069, 3.156476, 0.7418267, 1.336848, 4.044131, 5.131059, 3.386864, 
    3.655378, 4.486467, 4.921389, 4.197061, 3.642584, 4.948885, 5.263684, 
    7.513462,
  3.742634, 3.345432, 2.2659, 1.076696, 4.447221, 4.326276, 4.693994, 
    7.26801, 5.567674, 5.480121, 3.610262, 5.463867, 7.001881, 10.88335, 
    13.49804,
  2.666843, 3.705126, -0.7410621, 2.211224, 4.008677, 4.509508, 7.502392, 
    8.910254, 8.633676, 11.76557, 7.418527, 12.5914, 13.40681, 15.31748, 
    20.49517,
  -0.7159987, -0.900821, 0.1479765, 4.663583, 6.833539, 8.665475, 6.637954, 
    13.67203, 23.58749, 18.34795, 13.72489, 12.54233, 10.7812, 12.32434, 
    15.58037,
  0.1656243, 2.319293, 4.6616, 1.436163, 4.413756, 5.193686, 3.875297, 
    3.08334, 3.790123, 6.220513, 11.80471, 7.808686, 4.174501, 4.850694, 
    5.425972,
  -0.4810048, 0.2339258, -0.02573851, 2.509351, 6.494301, 6.170464, 3.517258, 
    5.724344, 7.29845, 8.398755, 10.49284, 7.870717, 5.806197, 3.527175, 
    3.013306,
  0.09525087, 0.3990347, 1.858006, 2.22869, 6.503281, 8.070031, 7.072868, 
    4.689245, 3.853079, 8.676162, 8.168503, 7.399605, 6.051108, 4.345552, 
    2.510798,
  3.396074, 7.430838, 13.4986, 6.545696, 5.845045, 5.822472, 11.16948, 
    3.665502, 3.3828, 7.581913, 5.995976, 5.7439, 4.811232, 5.000166, 3.107364,
  10.17889, 12.47121, 23.20735, 10.1699, 7.651584, 8.696817, 8.330287, 
    11.31826, 10.79297, 7.29486, 6.683514, 6.315381, 7.486825, 8.274854, 
    8.976293,
  16.10909, 22.72724, 25.21763, 18.95819, 10.98941, 8.652195, 9.420591, 
    10.30316, 9.119826, 7.338478, 6.434547, 4.645281, 4.534564, 4.585266, 
    9.946978,
  20.19512, 32.14788, 35.74609, 28.61042, 12.35305, 8.066519, 7.349457, 
    9.284249, 8.533371, 5.791759, 3.048462, 2.371394, 4.780166, 5.814444, 
    7.43925,
  27.16446, 40.23287, 42.4046, 25.55957, 14.24874, 7.569474, 3.72982, 
    4.817757, 9.813375, 11.83221, 10.62672, 11.34424, 13.22398, 18.93765, 
    21.57236,
  32.93812, 44.02299, 30.73703, 14.96282, 11.03172, 5.874668, 5.194036, 
    11.69511, 16.318, 24.25999, 13.91115, 11.207, 14.61318, 18.87906, 23.68738,
  27.59323, 26.8289, 20.92009, 9.799467, 6.554521, 4.963527, 9.056844, 
    19.48471, 34.27755, 23.0826, 13.31792, 10.44015, 11.54986, 16.24663, 
    20.19979,
  8.268119, 11.67398, 18.74247, 12.7673, 12.9837, 17.57036, 10.88553, 
    12.05954, 13.36845, 18.68342, 15.56008, 10.2344, 8.75268, 9.570903, 
    7.913126,
  26.15542, 24.93779, 12.69706, 12.46959, 20.62157, 15.4435, 9.594753, 
    10.6057, 11.12382, 14.0141, 13.59103, 13.55854, 9.372939, 8.184203, 
    11.64852,
  37.36398, 43.51627, 42.88236, 12.18546, 11.57405, 10.77279, 9.059589, 
    6.976532, 10.91507, 7.467656, 6.236696, 11.50407, 11.88964, 9.252571, 
    9.870075,
  39.7684, 46.66708, 53.53392, 21.16324, 12.2002, 6.876094, 6.595149, 6.5914, 
    8.886246, 12.30085, 5.577707, 5.414877, 5.393193, 11.92928, 11.99424,
  39.80787, 38.48735, 45.46465, 20.0787, 12.90341, 13.6537, 8.95077, 
    4.666912, 9.642086, 14.0267, 8.75152, 5.201325, 2.424131, 2.616125, 
    4.107554,
  38.45251, 35.44275, 31.99342, 24.01562, 17.19767, 6.201495, 11.3804, 
    13.1754, 12.40476, 8.992059, 3.43156, 4.952149, 6.949904, 1.707857, 
    1.664704,
  34.54494, 33.33323, 29.78918, 23.67758, 14.4497, 3.394742, 8.771663, 
    12.66904, 9.694573, 10.88727, 6.231199, 5.818328, 11.128, 7.076066, 
    2.797444,
  30.90437, 29.24553, 25.74581, 16.72448, 15.54472, 3.523092, 8.052455, 
    12.39412, 9.710041, 9.292461, 8.251925, 9.968689, 10.55197, 11.12713, 
    11.81029,
  25.08175, 21.168, 12.85898, 4.783157, 13.03908, 3.411011, 8.908837, 
    15.63343, 17.34891, 25.21638, 13.48447, 14.0674, 7.947894, 8.845376, 
    10.8716,
  10.07691, 5.60551, 8.211735, 5.117954, 9.635515, 5.058187, 6.865208, 
    18.52609, 29.62942, 19.77876, 14.60102, 12.70707, 4.821976, 6.654059, 
    7.499269,
  7.543873, 10.51484, 14.20067, 7.171754, 6.699269, 8.377863, 4.206725, 
    2.394727, 2.795386, 6.337041, 9.179949, 4.039693, 3.841182, 11.18928, 
    10.74164,
  11.73453, 12.52928, 10.37848, 8.139856, 7.306808, 5.350225, 3.813114, 
    4.150894, 4.011644, 3.325429, 3.954359, 0.7292451, 1.090856, 7.928382, 
    11.31894,
  14.78505, 17.74044, 14.30644, 6.697569, 3.440502, 5.833285, 4.681493, 
    5.217937, 6.499227, 4.936364, 4.616441, 3.304236, 2.452352, 3.897513, 
    6.944229,
  13.709, 15.87573, 13.12525, 3.603558, 2.919828, 3.348198, 3.718325, 
    5.692192, 7.882963, 6.16053, 6.965611, 3.71078, 3.016286, 5.401289, 
    2.860288,
  14.66679, 6.053901, 5.749027, -0.05362627, 1.248169, 4.315604, 6.11221, 
    5.330626, 6.118578, 11.84135, 6.776822, 3.11616, 3.564464, 6.132977, 
    3.392307,
  13.03205, 5.668536, -3.658348, -4.098618, 0.9486298, 2.407065, 4.780694, 
    6.226083, 8.185602, 9.498763, 8.484384, 2.307686, 2.589551, 2.807807, 
    5.887866,
  9.460395, 2.07667, -4.722362, -5.377267, -0.4242864, 1.420611, 4.49164, 
    4.560507, 7.180746, 5.702461, 7.745849, 3.331405, 2.250814, 5.359306, 
    6.682524,
  8.01103, 4.0963, -3.91676, -4.208228, -0.4284883, 2.553318, 2.252498, 
    4.625714, 7.778192, 7.171224, 8.339314, 3.29683, 2.012242, 7.983048, 
    9.616318,
  4.524299, 1.639648, -3.750426, -2.004682, 0.4665222, 2.483672, 3.958586, 
    7.521948, 10.57378, 12.42112, 2.698123, 2.674531, 2.093055, 4.164421, 
    13.8059,
  1.427397, -3.107951, -3.241139, 0.5419702, 4.125966, 3.75535, 6.157871, 
    13.05962, 17.3628, 7.08253, 3.706746, 3.277603, 2.664988, 2.965195, 
    12.00215,
  1.244221, 4.470081, 8.300922, 5.190804, 7.324387, 9.419172, 8.741382, 
    9.548864, 7.038557, 5.859206, 6.970069, 6.755681, 7.615614, 7.493334, 
    7.415357,
  -1.313506, -0.1845954, 1.592807, 4.184769, 5.12642, 6.040272, 6.514388, 
    8.883796, 5.558699, 4.43585, 4.098222, 6.121568, 6.930393, 8.837068, 
    7.264675,
  -1.803123, -0.9045669, 1.381377, 1.927863, 4.163505, 10.22108, 10.10711, 
    5.654576, 3.963351, 2.724377, 3.858508, 5.621318, 6.710712, 9.49201, 
    7.064321,
  -0.05637009, 4.524695, 8.331161, 4.668943, 6.262191, 7.389825, 11.22047, 
    6.893852, 8.558782, 11.76393, 7.156417, 7.449942, 7.672348, 9.447997, 
    6.828112,
  5.047029, 7.419824, 15.96922, 9.360303, 9.561107, 9.319517, 6.684943, 
    13.33366, 11.69252, 12.66022, 8.891078, 9.412317, 10.12041, 8.160169, 
    8.319633,
  10.86459, 17.83925, 18.65407, 18.27371, 16.60394, 14.45272, 13.31799, 
    11.30295, 10.76948, 13.07184, 8.713123, 8.759282, 7.298552, 5.90432, 
    4.475357,
  15.82459, 28.2417, 28.98735, 22.13422, 16.42811, 17.25995, 11.79275, 
    13.30018, 12.18856, 3.132445, 5.752433, 5.926584, 5.324461, 6.023223, 
    4.867625,
  22.68285, 37.18311, 33.57843, 19.27213, 15.53847, 14.67737, 15.12586, 
    15.19487, 9.304438, 3.199432, 1.985801, 2.436435, 4.060706, 5.906721, 
    8.795792,
  31.68187, 40.97467, 28.45724, 18.03641, 14.65133, 14.4525, 16.87537, 
    16.79188, 12.8919, 8.601127, 2.196365, 1.462218, 1.900501, 3.878307, 
    13.03079,
  33.15828, 30.58878, 28.26091, 17.14489, 12.48145, 10.31359, 10.59077, 
    16.92417, 17.40353, 5.857203, 1.601991, 1.371948, 2.267248, 4.277776, 
    10.2835,
  10.36752, 21.75031, 25.73421, 17.20876, 17.48476, 16.22233, 11.38585, 
    13.13427, 14.80223, 19.1037, 14.03898, 7.493299, 8.440176, 11.28384, 
    9.476693,
  30.07917, 32.63542, 22.80719, 23.10202, 18.97793, 15.52418, 9.128589, 
    11.60377, 15.10942, 20.87526, 18.15072, 8.791713, 5.885915, 7.293345, 
    5.905128,
  42.03172, 56.66647, 54.79564, 23.52861, 13.06026, 11.92237, 7.930973, 
    8.5783, 14.15322, 18.13033, 19.50916, 11.76527, 3.475718, 7.496347, 
    8.154464,
  48.37279, 62.29063, 72.91969, 29.35015, 11.40493, 9.118362, 5.748271, 
    8.050293, 11.45825, 16.9885, 16.28882, 10.15163, 5.952173, 7.129281, 
    9.657153,
  59.05313, 60.36237, 71.4994, 32.49512, 21.02246, 19.35811, 14.60057, 
    5.638838, 10.52401, 15.62673, 16.61417, 13.46664, 10.60736, 9.966841, 
    13.35141,
  63.83967, 67.36143, 63.88878, 45.61504, 26.36804, 17.22353, 18.31539, 
    16.27094, 12.06798, 6.424187, 6.273992, 9.291859, 11.27382, 10.8861, 
    9.443326,
  67.51764, 74.16679, 69.61843, 41.79775, 18.72739, 17.61614, 14.37636, 
    15.9981, 14.30499, 4.512282, 4.625561, 9.185205, 8.955407, 8.993142, 
    8.254757,
  76.13284, 80.37405, 65.20152, 28.17505, 16.42254, 16.44341, 14.66336, 
    13.38991, 14.28893, 4.634561, 2.759951, 4.873106, 8.139421, 8.476818, 
    13.41592,
  79.91587, 77.21473, 43.22423, 18.31657, 15.24963, 14.53213, 15.08874, 
    16.84451, 15.46071, 12.83811, 3.652556, 2.330044, 3.317807, 3.902057, 
    6.937844,
  69.69057, 51.12549, 31.45366, 17.96336, 14.73926, 12.05872, 14.28434, 
    21.96461, 20.41109, 5.576531, 1.311583, 0.6749693, 3.141037, 3.085479, 
    3.707304,
  7.788261, 12.54239, 16.29298, 12.37994, 13.37633, 8.263979, 4.486209, 
    0.5305662, 2.58313, 13.93897, 17.18447, 16.00582, 17.26668, 19.62749, 
    20.2491,
  36.01708, 25.0232, 13.11654, 15.124, 10.72167, 7.831036, 4.713512, 
    4.261922, 2.708591, 3.142119, 15.56493, 16.76794, 14.96099, 16.40793, 
    15.73848,
  56.91779, 54.91385, 42.45166, 14.26261, 8.575786, 8.147855, 7.611736, 
    8.081338, 6.868736, 7.911653, 15.29162, 17.59083, 15.07671, 11.18607, 
    14.81212,
  67.33114, 66.99439, 65.41519, 21.25418, 8.463194, 7.102389, 7.405868, 
    8.381824, 11.09642, 13.05888, 15.98343, 19.38771, 11.22813, 6.655738, 
    11.99982,
  78.08723, 64.76997, 71.46594, 29.46219, 14.41237, 8.252255, 7.524677, 
    4.0428, 6.997653, 14.96054, 13.72963, 17.13467, 12.55678, 7.158261, 
    8.70034,
  83.4107, 77.31784, 65.58454, 42.91259, 16.0757, 12.15718, 8.771298, 
    5.27845, 4.362533, 6.372791, 7.599556, 11.6662, 15.23296, 11.9879, 
    10.58494,
  83.98241, 84.18285, 73.89082, 38.57868, 15.36672, 14.57227, 8.363623, 
    7.878942, 4.032967, 3.841871, 6.733795, 9.450808, 12.76837, 15.61678, 
    14.27713,
  86.18893, 86.77129, 66.18061, 27.22847, 17.00579, 15.47513, 8.880021, 
    7.805938, 5.676408, 7.026134, 4.924709, 7.126463, 11.73489, 14.9915, 
    18.31984,
  77.02799, 78.5263, 39.79071, 19.74931, 13.04404, 11.04362, 12.43337, 
    15.65325, 12.01128, 11.07171, 12.68935, 10.76204, 9.801614, 14.97896, 
    19.22178,
  54.63742, 42.42622, 26.01818, 18.25164, 14.51734, 13.5083, 10.59087, 
    24.26449, 21.04493, 8.34916, 6.017454, 9.395905, 13.40465, 14.04948, 
    18.35579,
  5.497958, 10.63298, 13.82455, 16.51604, 12.90255, 11.80268, 2.36095, 
    2.277098, 2.138938, 10.44565, 10.33544, 7.026186, 14.18582, 16.45301, 
    5.868669,
  10.71849, 17.43632, 11.9308, 16.23636, 16.41888, 12.29827, 3.037429, 
    3.22322, 3.430655, 2.752931, 5.497829, 15.05231, 13.43055, 16.11197, 
    9.76103,
  22.41759, 37.58424, 35.7631, 13.12041, 10.33181, 11.72251, 4.499533, 
    6.61417, 7.742911, 3.926147, 2.705962, 15.22593, 14.85149, 13.13087, 
    14.87948,
  34.0408, 47.35454, 51.02075, 22.81458, 9.652601, 5.027293, 5.781477, 
    9.741521, 13.92972, 13.79483, 6.712567, 12.88325, 12.73281, 8.176485, 
    11.64019,
  47.12363, 48.00031, 52.5615, 25.76431, 14.79293, 10.45373, 3.724363, 
    3.962574, 6.650102, 16.91203, 14.44213, 11.83243, 13.28423, 10.92467, 
    11.56099,
  53.12973, 55.53384, 48.42036, 32.89751, 20.94374, 16.80771, 8.463005, 
    7.216911, 6.816639, 7.978067, 9.006588, 10.95632, 10.873, 8.043322, 
    8.784369,
  54.55634, 61.28771, 51.69132, 28.44593, 18.32267, 17.67397, 14.18941, 
    15.01316, 10.18778, 8.288295, 11.28289, 11.89467, 10.6828, 10.60747, 
    11.61609,
  57.32635, 64.93594, 45.03381, 18.859, 16.27518, 16.75013, 14.37232, 
    16.08939, 15.1443, 10.64509, 12.33777, 13.38376, 10.95795, 11.80349, 
    14.7345,
  56.4032, 62.90526, 30.1568, 14.65042, 13.00666, 15.48983, 16.30471, 
    23.55122, 20.99109, 20.38221, 16.42139, 14.34084, 12.96846, 8.285271, 
    14.86078,
  46.6337, 39.83, 17.94389, 15.77668, 14.15324, 15.26583, 18.20901, 34.83502, 
    32.35036, 19.39153, 13.72505, 14.23088, 14.92675, 10.97943, 7.511686,
  7.723525, 12.89664, 17.17033, 4.528055, 7.528371, 5.674405, 5.455461, 
    5.31775, 3.553384, 9.766903, 12.82416, 12.36608, 12.15658, 14.22201, 
    11.6998,
  30.84887, 33.69226, 12.21353, 4.679984, 8.104187, 5.859103, 7.765375, 
    7.345448, 4.841114, 0.09290411, 7.439428, 13.63951, 6.703254, 11.26171, 
    9.067771,
  70.85416, 76.17008, 43.22066, 10.80556, 8.686883, 5.884037, 9.981493, 
    12.62571, 12.71708, 6.017685, 0.611897, 11.28273, 7.125917, 11.50421, 
    10.85069,
  82.12918, 77.50759, 61.08959, 22.19265, 14.80148, 4.954791, 9.995506, 
    18.53751, 22.11407, 16.35036, 2.141635, 10.9724, 8.646955, 4.122733, 
    12.11562,
  85.11153, 66.66723, 57.60413, 25.27261, 16.59992, 15.47751, 10.95483, 
    8.555141, 14.91551, 20.46667, 9.455559, 9.620892, 7.833592, 4.523813, 
    9.525325,
  78.74191, 65.92197, 51.36137, 31.90904, 20.56328, 16.42865, 15.18082, 
    11.59523, 9.825571, 9.503582, 7.685043, 11.46527, 9.598631, 9.939899, 
    5.458674,
  70.1334, 65.2062, 52.82906, 26.65571, 18.6771, 17.30482, 15.67264, 
    12.43676, 10.83189, 10.2872, 8.466265, 12.35121, 9.816046, 12.13595, 
    3.590798,
  68.08203, 64.40808, 42.90957, 19.70082, 18.41584, 19.60584, 16.56686, 
    11.14411, 10.70178, 12.22532, 11.24105, 7.326735, 11.21783, 11.56732, 
    10.7167,
  62.66553, 60.48977, 25.83979, 13.57955, 16.9887, 13.03612, 13.33406, 
    20.06588, 18.18107, 20.41701, 12.56583, 8.852895, 4.777715, 6.885974, 
    14.54075,
  52.07021, 40.38333, 14.16873, 12.77323, 14.83105, 7.116243, 12.74642, 
    38.95681, 34.23039, 15.04469, 7.978414, 6.551807, 7.439723, 6.425334, 
    9.298005,
  11.35785, 17.93757, 16.75392, 3.589066, 3.279122, 4.821199, 3.538975, 
    3.398077, 5.227629, 13.14487, 15.37409, 13.1763, 10.78499, 13.91124, 
    17.28684,
  39.93188, 23.90604, 10.35822, 5.181627, 6.911847, 6.170638, 5.357174, 
    8.079648, 7.226909, -0.2031514, 13.47705, 12.0284, 10.31809, 12.31236, 
    16.7494,
  66.87605, 60.62223, 37.50784, 11.07022, 8.753541, 7.014472, 9.745265, 
    10.7747, 9.713295, 6.983955, 5.455486, 11.07452, 10.37136, 10.78256, 
    12.75255,
  63.23594, 62.197, 59.59195, 17.32729, 10.67617, 8.56212, 7.493298, 
    13.58891, 17.57162, 13.37139, 8.413488, 12.78106, 13.2591, 9.4663, 
    8.030831,
  59.28547, 53.8509, 61.5587, 23.90729, 16.07461, 11.61527, 5.848393, 
    8.176632, 16.85364, 19.41058, 9.543209, 14.50158, 12.96873, 11.97238, 
    8.440109,
  50.04458, 49.82516, 52.86028, 33.60735, 18.29867, 12.28313, 5.431341, 
    6.799468, 9.465259, 10.58261, 8.789017, 13.97831, 14.30961, 14.23154, 
    11.22473,
  46.43584, 42.42823, 45.2118, 24.56499, 16.84744, 13.92831, 10.8602, 
    6.379042, 8.344514, 11.31656, 8.001163, 10.01378, 14.01595, 15.85071, 
    13.01869,
  48.01973, 38.51752, 26.46797, 12.71989, 13.71717, 15.65554, 14.86861, 
    8.280451, 7.686664, 10.83334, 9.798966, 8.255592, 10.20977, 17.39069, 
    17.45062,
  48.0521, 39.10248, 14.32099, 8.298391, 7.458748, 11.04567, 16.42772, 
    24.64387, 23.64751, 23.58349, 12.23726, 8.161564, 9.572968, 14.65996, 
    16.15636,
  42.28028, 27.13686, 10.96229, 9.885885, 4.44673, 7.261267, 13.46045, 
    37.08798, 36.02269, 20.10816, 5.568185, 5.290951, 9.539105, 11.17949, 
    13.50675,
  6.877773, 9.037984, 9.104986, 7.109881, 5.704978, 6.094941, 3.25515, 
    9.411878, 11.94612, 13.64448, 16.42357, 10.98765, 10.34775, 11.42545, 
    12.44482,
  13.14207, 8.028597, 9.863694, 13.09799, 12.37592, 7.171238, 3.202533, 
    12.42135, 13.31201, 10.44944, 11.98978, 8.869003, 9.314709, 15.50725, 
    17.07323,
  30.80671, 32.14265, 25.34835, 18.28952, 12.34094, 10.14124, 4.86982, 
    5.71305, 10.02265, 10.50925, 10.67626, 8.402069, 7.492185, 12.41626, 
    15.85843,
  36.15508, 34.08738, 39.98062, 18.81739, 12.13618, 6.230558, 8.854513, 
    8.919893, 14.5953, 13.8439, 10.22269, 9.29283, 10.34161, 10.36787, 
    11.73156,
  46.07389, 30.57623, 39.37285, 23.54445, 15.00002, 13.82146, 12.66904, 
    11.38496, 16.11139, 19.59479, 10.46683, 9.945402, 10.55811, 10.2803, 
    11.31176,
  57.44955, 34.30546, 31.95851, 24.24259, 15.58712, 14.15919, 14.79177, 
    12.65418, 12.4473, 8.837792, 8.112703, 8.700965, 11.32683, 9.630307, 
    10.86571,
  65.69898, 40.15903, 26.43834, 11.46893, 14.18733, 13.99947, 15.89493, 
    17.62473, 15.77666, 11.8176, 10.25569, 10.30039, 11.04058, 10.86047, 
    8.496489,
  73.38629, 46.17716, 18.57071, 4.205355, 13.4908, 12.89226, 16.48267, 
    18.79839, 19.05816, 15.53961, 13.08444, 11.23819, 11.55291, 12.87622, 
    8.456088,
  67.27866, 40.19442, 13.19443, 3.579009, 5.335648, 12.28688, 16.15636, 
    25.9921, 29.07544, 27.04084, 16.81115, 12.65586, 11.56562, 12.19334, 
    11.37902,
  49.91341, 18.26696, 7.585292, 4.710471, 6.341158, 10.14496, 9.891314, 
    37.44408, 37.28421, 21.88426, 14.4512, 11.87831, 10.68866, 10.9725, 
    11.58968,
  6.715446, 12.32842, 15.40867, 13.5513, 11.59027, 11.82118, 10.94069, 
    12.2537, 12.28413, 17.73377, 16.90086, 15.43751, 17.44181, 12.21171, 
    17.78164,
  17.70734, 10.93483, 15.17389, 16.35677, 15.65972, 15.57414, 10.76095, 
    6.667201, 3.705227, 13.39162, 16.44334, 12.08938, 13.7738, 13.42055, 
    15.81255,
  35.43459, 25.01751, 21.38885, 18.77332, 15.44243, 15.40972, 7.542663, 
    5.690144, 8.874345, 14.487, 14.39789, 14.15691, 12.36062, 11.84439, 
    11.17253,
  48.96354, 32.76634, 36.03181, 20.20765, 14.65326, 12.49079, 14.93885, 
    6.875226, 9.13181, 16.90089, 16.40772, 14.27134, 14.52286, 10.31567, 
    10.18725,
  59.98302, 36.29417, 35.81968, 22.06321, 14.08583, 16.25264, 15.05528, 
    11.55524, 14.58602, 22.22334, 19.07607, 15.88473, 14.19593, 8.40904, 
    8.042676,
  62.94639, 41.53881, 31.816, 21.91334, 12.04593, 14.38371, 16.40047, 
    14.97195, 12.50569, 14.32856, 16.41163, 14.70934, 11.76592, 8.495184, 
    8.116351,
  58.74076, 42.3931, 28.86825, 12.40123, 12.77734, 14.38322, 18.00116, 
    18.13213, 17.18326, 17.54985, 17.13127, 14.40718, 12.7266, 11.28407, 
    5.468468,
  54.3919, 42.33194, 19.76437, 9.572264, 12.12735, 11.40301, 17.64375, 
    19.55089, 17.48983, 19.41254, 16.01506, 16.23544, 12.23507, 7.434124, 
    5.984286,
  45.92741, 32.06921, 7.809226, 9.44243, 10.58931, 9.54985, 13.95936, 
    25.2734, 29.087, 29.45703, 21.58056, 16.37145, 13.38892, 5.385533, 
    6.756722,
  32.37474, 14.16473, 7.048883, 9.296768, 9.717568, 4.097017, 10.80062, 
    34.12718, 36.08545, 20.31762, 17.90829, 13.71879, 11.6866, 3.71448, 
    8.768255,
  8.032938, 13.40899, 17.46134, 14.55382, 13.8927, 12.60248, 14.06647, 
    11.57778, 6.212943, 16.84036, 20.15572, 18.08376, 18.59307, 17.50483, 
    20.34146,
  14.15094, 15.83059, 16.80738, 15.31092, 17.03792, 14.64316, 12.82467, 
    3.282656, 2.676466, 10.93109, 16.07293, 13.44213, 10.77262, 11.60975, 
    20.65064,
  29.04327, 33.709, 24.82872, 18.05468, 10.74806, 17.03085, 8.667212, 
    6.448468, 3.290141, 13.33934, 12.1704, 15.54228, 12.62144, 12.23847, 
    13.95635,
  37.4792, 42.73972, 34.58543, 19.54142, 11.91254, 12.80322, 14.46933, 
    8.775954, 5.992656, 7.6039, 12.89282, 14.39744, 14.33007, 15.11819, 
    15.15899,
  50.61591, 42.19562, 31.38528, 17.47073, 9.34383, 8.746971, 9.051016, 
    9.576797, 11.56098, 16.10034, 16.2179, 13.13513, 15.83627, 11.39718, 
    7.911573,
  57.47873, 50.81962, 24.05222, 12.77381, 8.277163, 7.34896, 10.71494, 
    10.21269, 11.75575, 13.64055, 14.86159, 13.71863, 14.44407, 6.721284, 
    7.668416,
  61.46396, 56.14077, 30.6185, 12.49082, 11.37968, 8.764655, 9.78797, 
    11.54253, 12.21446, 11.31664, 8.989518, 11.02408, 16.12036, 8.084015, 
    9.628716,
  67.51611, 64.33193, 28.68892, 12.97747, 12.03119, 9.368281, 7.895267, 
    10.13105, 11.55603, 11.355, 11.10521, 13.39695, 16.42082, 13.65259, 
    14.91258,
  72.66519, 61.98514, 18.9039, 12.65535, 15.56976, 13.16374, 8.6936, 
    10.42161, 13.59324, 17.77401, 11.82845, 12.96494, 13.08655, 12.36268, 
    13.97696,
  61.59923, 36.33981, 19.61254, 21.14592, 17.80334, 12.85232, 10.34087, 
    14.54907, 16.15623, 13.56748, 13.05512, 15.82899, 7.782891, 13.37257, 
    16.93018,
  6.988168, 14.58731, 21.36469, 15.87329, 16.55819, 18.98514, 6.48487, 
    5.748143, 10.17361, 16.85793, 20.13411, 17.75896, 17.18468, 16.31911, 
    18.27447,
  13.14603, 14.73461, 19.53094, 18.19739, 22.31904, 21.99365, 8.283031, 
    5.871309, 3.533367, 5.052707, 7.642642, 10.68006, 9.154794, 14.33224, 
    17.89424,
  32.20904, 33.30395, 22.87098, 15.086, 14.7598, 13.67892, 13.41511, 
    8.261147, 5.752046, 3.779579, 4.820117, 6.423785, 8.890957, 12.05176, 
    13.87286,
  43.2401, 41.81089, 36.675, 18.37753, 10.34746, 11.7197, 12.03605, 13.41238, 
    8.015157, 6.624731, 9.026718, 7.559973, 9.274303, 14.49922, 13.0188,
  59.85962, 46.15721, 50.43934, 27.95314, 14.75616, 12.56081, 11.66955, 
    8.400148, 7.338661, 6.740156, 6.414222, 8.708827, 10.33078, 13.62807, 
    10.64329,
  70.78371, 66.94212, 58.70377, 28.18425, 14.54559, 14.30024, 13.28745, 
    12.534, 11.27554, 8.380885, 6.996848, 10.10637, 12.05523, 10.53325, 
    12.13315,
  80.68179, 82.66698, 67.88811, 15.67459, 11.52004, 8.546787, 8.493925, 
    7.819068, 7.813515, 4.67627, 12.11533, 11.08967, 10.03197, 9.201376, 
    13.22907,
  90.65591, 89.14076, 50.79412, 14.08298, 11.98691, 10.73949, 6.574195, 
    10.51063, 11.50758, 3.085277, 9.857298, 7.959059, 10.18751, 17.09851, 
    23.21509,
  91.80629, 82.54716, 35.17587, 14.06592, 14.89615, 13.17996, 10.21679, 
    13.03515, 12.18792, 4.601978, 7.524978, 5.916307, 8.924169, 22.22228, 
    21.27428,
  76.30461, 60.19405, 29.62939, 21.20521, 17.41319, 12.77367, 8.705235, 
    13.34109, 21.14364, 17.75307, 6.946431, 12.79927, 14.67774, 22.60614, 
    22.09202,
  5.758521, 4.144353, 15.40836, 7.154235, 8.318884, 10.00456, 6.684937, 
    8.629564, 8.519511, 13.71324, 17.23175, 16.61023, 15.32006, 16.20073, 
    17.88052,
  17.97244, 6.165878, 10.25692, 8.78434, 15.91778, 16.85887, 11.03248, 
    8.31284, 9.212755, 11.96214, 14.97437, 12.41554, 11.1913, 14.96146, 
    15.82956,
  27.89193, 25.78156, 15.33184, 5.338192, 9.385045, 17.36632, 13.61965, 
    7.306216, 11.88844, 12.18046, 10.44772, 11.70048, 6.824229, 14.85359, 
    14.33676,
  39.82492, 36.1503, 28.85627, 10.21252, 6.616817, 13.24106, 15.91691, 
    10.94572, 4.839775, 12.42847, 9.137789, 11.4031, 10.59546, 15.14121, 
    11.95374,
  52.76485, 37.26874, 32.64409, 11.17803, 6.369572, 8.626211, 11.58239, 
    10.01306, 9.633202, 8.413174, 14.12192, 10.60822, 9.783205, 17.21995, 
    5.587873,
  61.12614, 50.61601, 27.63655, 16.08952, 12.1036, 9.042233, 9.617579, 
    8.030116, 8.922023, 4.935393, 11.73426, 13.60527, 10.4189, 7.651951, 
    5.035066,
  70.51151, 59.91182, 35.5963, 15.06801, 11.05229, 8.103308, 6.864552, 
    9.055945, 8.437325, 3.462355, 6.688447, 13.19036, 13.73597, 7.310639, 
    10.22237,
  79.30586, 69.73057, 32.66395, 13.81376, 16.25866, 9.875713, 10.17919, 
    12.12691, 8.070483, 14.09785, 9.442122, 8.119615, 14.42429, 10.8417, 
    18.06678,
  83.64369, 68.21067, 22.79014, 13.05622, 10.89057, 6.844739, 9.962316, 
    12.59793, 13.95575, 19.05423, 7.614426, 10.33541, 13.91198, 13.62971, 
    20.87919,
  70.19955, 48.85879, 18.75615, 14.90191, 9.480453, 7.694837, 9.683227, 
    18.28109, 23.41896, 17.13432, 10.26805, 13.40421, 10.24373, 15.69835, 
    17.24927,
  3.41916, 6.399547, 18.82784, 15.36017, 14.27095, 10.07725, 8.130836, 
    6.48456, 7.512996, 17.87113, 17.43375, 12.82426, 16.01165, 11.66127, 
    19.28174,
  5.51868, 5.364141, 8.640143, 10.97676, 20.33237, 17.72381, 6.507685, 
    8.911247, 7.405794, 12.67116, 13.49379, 9.097746, 8.511516, 12.47788, 
    16.3798,
  10.5684, 8.535389, 5.734289, 9.134773, 12.80533, 18.47189, 8.1623, 
    8.924248, 8.796438, 11.067, 8.351424, 7.109838, 8.812653, 8.957376, 
    15.21499,
  24.53983, 19.74155, 15.78221, 3.312295, 3.153027, 9.728602, 15.019, 
    11.14214, 7.279611, 11.29912, 8.347478, 5.233195, 11.348, 6.71005, 
    13.55889,
  43.03109, 27.51895, 21.33971, 4.99752, 4.897422, 4.526624, 6.639979, 
    9.573494, 8.768583, 7.433813, 12.49356, 6.500053, 7.392779, 10.59538, 
    4.798046,
  56.19929, 37.51949, 16.37327, 10.72934, 7.332155, 3.402068, 5.102149, 
    8.082973, 10.55772, 9.216221, 17.21273, 11.5663, 14.17847, 5.702229, 
    8.225226,
  62.46968, 44.52326, 22.8886, 6.648243, 10.00295, 1.573771, 3.914957, 
    6.099509, 10.11058, 8.476004, 15.01202, 11.41865, 12.74573, 5.297674, 
    10.84335,
  70.60891, 55.17264, 22.48785, 7.664191, 10.72282, 4.231557, 3.434581, 
    9.633255, 7.798875, 12.0011, 15.59923, 12.59197, 7.172909, 8.505163, 
    13.81146,
  77.33337, 59.60653, 16.78634, 12.37951, 7.364282, 9.732648, 11.63833, 
    15.45365, 13.27501, 14.49084, 7.570954, 8.280279, 4.959667, 17.00337, 
    12.59407,
  64.3293, 41.51203, 11.46606, 15.39434, 11.10596, 11.36327, 14.73824, 
    23.50173, 14.48728, 16.6015, 7.786547, 12.56713, 5.096466, 12.38565, 
    10.60094,
  3.470348, 1.598784, 4.286116, 2.00978, 4.953644, 5.755564, 4.761757, 
    6.976323, 4.407186, 15.94563, 12.42478, 8.111403, 12.87918, 15.64314, 
    24.05506,
  1.931205, 1.620348, 1.138003, 2.754, 8.181417, 7.480316, 5.592053, 
    7.792187, 5.140991, 11.22696, 17.23702, 5.645305, 6.772675, 14.96106, 
    20.00131,
  6.918729, 6.226316, 3.567798, 6.211318, 8.167244, 10.20765, 6.94675, 
    8.520072, 6.10383, 8.497935, 7.714614, 7.207084, 6.707394, 6.506366, 
    16.57839,
  32.41836, 29.76659, 24.94728, 8.978434, 5.023924, 6.507331, 7.904821, 
    11.04634, 5.869526, 8.261843, 9.68153, 8.361945, 4.680731, 4.542126, 
    11.71207,
  50.73875, 37.22104, 28.47091, 7.916408, 5.340957, 4.057829, 6.047693, 
    9.448908, 10.40038, 8.844907, 11.149, 13.91133, 6.269876, 3.461936, 
    4.675937,
  65.80371, 47.85772, 26.43733, 8.402964, 8.092356, 5.977933, 6.912254, 
    7.496046, 11.67754, 7.759419, 17.37096, 16.59704, 10.5872, 2.700231, 
    4.812826,
  70.47691, 45.01426, 24.39629, 9.575099, 8.485152, 6.672758, 9.777321, 
    4.701339, 8.570476, 6.121338, 19.71607, 16.78115, 15.09296, 7.233111, 
    12.84766,
  73.842, 50.8105, 18.43439, 4.838503, 7.411382, 6.732572, 5.453052, 
    6.679747, 7.18866, 4.50483, 14.86724, 17.95739, 7.101927, 9.65196, 
    18.54373,
  77.81596, 56.04181, 9.562604, 7.403165, 6.917504, 5.547619, 5.945759, 
    9.780274, 12.12716, 6.198795, 19.65711, 16.99339, 5.172892, 14.00076, 
    20.04161,
  66.02103, 42.57501, 13.39648, 13.25265, 6.786126, 7.434832, 9.834175, 
    17.59281, 14.81393, 12.62055, 22.31433, 18.86478, 6.055626, 17.35842, 
    16.52699,
  4.440773, 0.935373, 1.836842, 5.136169, 4.805624, 12.32139, 12.42274, 
    11.13585, 10.00546, 14.8221, 15.35668, 10.60103, 17.1867, 18.0545, 
    24.94994,
  1.335128, 0.4035858, 1.225007, 1.461839, 14.43114, 21.05404, 15.1633, 
    10.74721, 7.030887, 4.979886, 17.15174, 8.44484, 8.978731, 18.4598, 
    17.50628,
  5.732718, 5.54884, 3.289299, 2.031373, 12.7457, 21.05577, 11.96608, 
    3.418024, 8.012986, 3.716095, 11.89727, 10.11971, 8.672002, 7.580273, 
    11.71469,
  29.66675, 32.18366, 26.26745, 12.37096, 6.644321, 12.12986, 20.47025, 
    7.247484, 4.814388, 3.125429, 1.89548, 2.071212, 7.695697, 5.756413, 
    12.17127,
  52.99577, 40.11333, 32.91888, 9.231688, 11.56434, 11.46352, 9.987489, 
    11.40099, 5.459105, 8.754288, 4.195682, 4.817511, 7.159888, 6.330563, 
    7.506321,
  59.96083, 43.57471, 22.52403, 6.040102, 9.66155, 6.105524, 6.197764, 
    5.165223, 9.979511, 9.40985, 11.1813, 5.463935, 6.741442, 9.117826, 
    15.16746,
  58.01385, 40.16736, 21.15391, 5.669014, 7.738391, 8.493499, 6.197567, 
    5.401595, 8.03669, 6.363265, 8.122191, 7.36571, 9.031854, 13.11964, 
    16.15543,
  53.65418, 42.31271, 18.71255, 3.544302, 9.441879, 5.055749, 8.689484, 
    11.50783, 8.766451, 5.689193, 11.74093, 13.06111, 14.80841, 17.97929, 
    18.60157,
  56.9262, 40.20219, 11.14954, 13.12771, 11.85514, 8.119285, 11.90206, 
    14.77882, 11.65609, 6.389435, 12.8622, 14.37332, 15.31828, 17.69933, 
    16.24724,
  49.78788, 29.56965, 7.989432, 10.98966, 8.315238, 9.673043, 14.62434, 
    21.16737, 14.78967, 14.89439, 14.99697, 15.1513, 15.85429, 14.2468, 
    14.5211,
  1.052689, 0.7501506, 2.304278, 6.520503, 9.03481, 10.45967, 9.76571, 
    11.68762, 13.10699, 22.29563, 21.91487, 19.61813, 21.82584, 21.25393, 
    23.95694,
  5.347018, 2.48928, 1.567117, 8.379306, 11.05763, 12.55954, 11.41524, 
    11.97271, 11.9905, 16.91637, 18.32184, 17.37962, 15.50281, 24.7383, 
    24.90141,
  11.82696, 9.254821, 3.571768, 3.671124, 8.77551, 25.10318, 10.18189, 
    8.902757, 11.50325, 8.047616, 11.18657, 13.59886, 9.461036, 8.53809, 
    16.05809,
  19.97728, 23.08619, 20.62702, 3.566925, 1.721893, 7.676376, 22.00702, 
    6.438002, 12.17006, 13.12591, 11.26496, 6.91775, 2.312179, 4.580326, 
    12.12995,
  34.00259, 28.56869, 24.14772, 7.25853, 2.584663, 16.26124, 15.26428, 
    17.72865, 10.89865, 10.07385, 4.452502, 2.635291, 3.263027, 6.193014, 
    13.91254,
  40.67054, 35.08469, 26.02567, 9.967152, 11.24074, 13.09078, 12.05595, 
    8.71802, 9.849376, 5.435528, 5.86449, 3.433906, 8.025795, 10.10168, 
    14.84558,
  43.42514, 36.2203, 33.22927, 10.11053, 10.36821, 9.834541, 8.866509, 
    1.948306, 8.311742, 11.90319, 11.15211, 11.1599, 10.04215, 13.69344, 
    14.88597,
  44.08069, 47.11649, 25.80785, 7.070641, 7.454569, 3.390037, 3.663836, 
    4.851125, 3.612683, 9.46818, 8.89183, 10.30584, 13.2621, 16.57192, 
    18.10151,
  50.11969, 42.54392, 12.30128, 13.18132, 10.55694, 9.530314, 8.521116, 
    7.470567, 6.007597, 10.76812, 11.48088, 11.41694, 15.06773, 16.67263, 
    17.39165,
  43.7768, 30.97469, 11.94502, 14.8698, 11.80369, 10.0062, 8.449228, 
    7.469568, 11.11986, 14.74647, 17.2108, 14.0577, 16.36047, 15.42101, 
    16.7048,
  2.144505, 6.080233, 11.77136, 10.63235, 10.84712, 8.777886, 5.925197, 
    6.006824, 6.056172, 14.97975, 17.06913, 10.86444, 15.12529, 19.03837, 
    26.41262,
  4.324714, 3.248855, 4.269198, 11.75312, 14.89522, 16.16823, 7.092555, 
    6.821553, 6.993706, 10.46843, 15.31244, 10.75604, 9.87288, 22.95229, 
    23.72966,
  14.44616, 15.47274, 12.28631, 4.3065, 11.48192, 16.73623, 8.197906, 
    8.827467, 6.828997, 6.53932, 4.903303, 7.693083, 6.531944, 9.864511, 
    17.83292,
  27.76869, 29.33716, 22.60102, 7.551906, 4.186845, 14.31643, 20.86104, 
    9.005829, 4.254632, 14.79586, 13.02174, 7.047089, 6.689968, 8.532854, 
    12.9825,
  43.70464, 27.53937, 23.58735, 11.00887, 2.926831, 10.04625, 11.55812, 
    11.93144, 11.33844, 12.61861, 12.73752, 8.089684, 8.910219, 6.922346, 
    8.107888,
  44.6056, 36.81124, 28.27929, 10.91459, 5.142582, 10.31083, 10.61095, 
    6.773502, 9.353306, 8.319029, 6.476787, 6.17582, 5.690903, 9.746386, 
    13.07007,
  50.15731, 45.59332, 26.10708, 11.27542, 10.68097, 10.55702, 8.129569, 
    7.231575, 9.371279, 7.022415, 9.401423, 9.522603, 9.287497, 10.68174, 
    15.37757,
  57.92001, 49.67648, 18.65388, 8.40789, 12.57255, 8.703609, 6.032892, 
    5.045874, 1.99284, 8.495312, 7.718342, 8.015544, 11.53883, 13.41586, 
    14.53105,
  51.43838, 44.08336, 12.96223, 14.38689, 13.09901, 6.788805, 2.507638, 
    2.512784, 9.483463, 11.1537, 7.875422, 7.440582, 10.07455, 13.05326, 
    14.95724,
  38.07165, 32.0876, 15.74259, 13.26029, 7.405261, 5.007724, 4.403766, 
    6.736693, 11.77304, 14.58883, 8.139724, 12.23351, 13.05124, 13.96414, 
    14.79467,
  -6.264443, -26.91908, -15.76665, -14.22732, -9.858509, -8.358551, 
    -5.107698, -4.201129, -2.115158, 5.386226, 12.57308, 12.59485, 20.80372, 
    15.4069, 24.27922,
  -18.38193, -18.65717, -13.39192, -10.53487, -14.00443, -3.708397, 
    -3.870043, -0.6874745, 1.677173, 4.733657, 14.41184, 10.46583, 6.928644, 
    21.46854, 20.85795,
  -11.42867, -12.64906, -15.055, -11.10361, -3.624645, 4.983511, 2.076541, 
    2.070671, 5.002807, 6.448273, 7.043623, 6.686728, 4.527479, 2.530141, 
    10.42522,
  -3.110432, -7.104531, -4.042145, 0.365202, 1.057706, 6.749112, 11.30297, 
    4.323905, 5.341418, 5.156525, 4.829545, 3.334956, 14.51175, 14.17705, 
    7.060547,
  8.241092, 6.544611, 16.37358, 11.58074, 5.05667, 8.749697, 15.82717, 
    18.77068, 12.63701, 9.120246, 6.616762, 12.17869, 15.13031, 13.18904, 
    11.14101,
  60.11948, 60.38732, 47.54123, 20.83272, 14.67541, 10.84366, 7.214947, 
    7.644832, 10.11096, 4.429972, 6.977515, 1.881778, 14.95483, 13.03328, 
    9.512226,
  94.09591, 95.78027, 50.21995, 14.34904, 9.104912, 5.580969, 3.991683, 
    5.047433, 14.06457, 16.1166, 12.34384, 7.208489, 8.774491, 10.36505, 
    8.386978,
  102.5459, 95.9594, 30.68114, 8.209728, 7.019981, 17.36933, 11.21885, 
    16.42733, 13.11646, 13.97365, 5.993882, 4.680654, 5.620656, 11.02952, 
    11.60903,
  83.43255, 67.17517, 14.00094, 12.93116, 18.39815, 13.02088, 12.63881, 
    17.56543, 17.72518, 16.12977, 6.029284, 10.73522, 11.40555, 13.88137, 
    11.8197,
  55.26129, 37.79902, 18.34386, 15.96182, 16.33379, 19.56311, 18.5231, 
    17.8549, 15.714, 17.65476, 10.78538, 13.64742, 12.78928, 10.38169, 
    12.59964,
  11.70683, 18.3653, 22.05735, 21.35564, 17.823, 11.51751, 4.735464, 
    1.644286, 0.6695574, 1.7284, 0.05061525, -0.4486395, -1.308524, 
    0.7032454, 1.888583,
  18.97146, 27.81887, 29.98421, 19.7122, 13.44842, 7.678746, 0.9938695, 
    -0.2975031, -0.7553866, -0.8598412, -1.186297, -1.802809, -1.537413, 
    5.004765, 4.362836,
  43.34818, 48.19139, 28.62408, 9.719898, 6.125013, 10.12792, 1.395843, 
    3.173033, 2.980876, 2.706105, 1.875983, 2.172699, 2.459804, 4.02887, 
    8.577732,
  63.40197, 50.46941, 31.787, 13.47458, 2.789614, 4.253912, 15.40375, 
    10.02647, 11.71651, 9.065326, 9.387792, 7.628645, 6.484832, 6.159632, 
    10.56827,
  64.80869, 44.49906, 43.2963, 20.05289, 11.14091, 10.49652, 19.38328, 
    15.83837, 10.018, 13.70175, 10.7021, 9.349363, 9.265002, 11.87735, 
    16.37517,
  60.02435, 63.00847, 55.74553, 24.50939, 17.19982, 14.48721, 11.64689, 
    15.61131, 15.34928, 13.88967, 13.69555, 12.09923, 14.02626, 15.73234, 
    17.01669,
  59.84966, 68.89664, 51.08505, 20.02444, 14.9987, 12.00825, 9.590569, 
    8.552321, 9.06249, 14.59465, 15.66996, 16.18767, 16.59928, 16.53682, 
    16.47891,
  63.06342, 71.44791, 35.47479, 21.75402, 18.09976, 13.70917, 8.010562, 
    6.203384, 5.150041, 8.54986, 8.944345, 12.02746, 13.36598, 15.92315, 
    15.14301,
  63.22895, 56.7981, 25.15486, 24.76536, 23.66552, 23.07464, 14.9363, 
    13.58038, 10.05381, 5.923649, 6.326432, 6.706583, 10.55296, 11.04525, 
    16.36906,
  52.81639, 37.13614, 22.14342, 21.82749, 19.80278, 19.42467, 20.10823, 
    11.49558, 12.55115, 11.77539, 10.3223, 10.45848, 13.3746, 13.66767, 
    11.12703,
  8.61282, 13.19019, 20.99467, 16.19617, 20.3016, 15.36298, 14.3207, 
    13.00137, 14.2318, 19.47133, 20.27602, 16.66297, 21.82516, 18.87853, 
    19.57307,
  8.931422, 15.11815, 20.62332, 15.87441, 19.08537, 23.65466, 16.63254, 
    13.53898, 15.80025, 15.24474, 19.83048, 18.36449, 11.24722, 17.9357, 
    14.3031,
  19.25789, 27.46902, 30.80114, 15.90826, 13.28791, 29.64966, 20.60552, 
    9.186102, 14.88309, 14.16381, 16.24588, 17.43419, 16.31824, 8.04283, 
    7.489881,
  33.37011, 39.16499, 42.05682, 23.48958, 5.646733, 14.72783, 23.27662, 
    13.37562, 12.19009, 16.19726, 16.47249, 17.39671, 15.90833, 5.475546, 
    2.692462,
  60.91443, 50.03797, 50.10135, 13.38111, 3.266021, 3.95399, 18.40044, 
    12.40837, 15.43968, 22.1876, 22.15912, 15.78539, 14.36921, 3.224076, 
    1.365597,
  77.59283, 62.79076, 42.37325, 6.189962, 2.23694, 3.470289, 14.16137, 
    13.99688, 16.2916, 15.16584, 17.86453, 19.82048, 11.02004, 4.586681, 
    3.112336,
  70.79397, 61.76108, 35.25137, 10.60156, 3.9342, 4.566758, 3.913487, 
    10.88775, 9.471572, 5.648141, 7.957106, 15.45097, 7.279519, 5.201444, 
    6.92552,
  60.00951, 51.22642, 21.07968, 13.89341, 13.54323, 13.45732, 5.23887, 
    2.781708, 7.240596, 2.539653, 11.83644, 11.86721, 5.666739, 7.145016, 
    10.83524,
  48.17029, 33.7452, 13.10373, 14.78285, 16.53254, 17.34003, 7.411523, 
    3.329941, 2.412639, 2.471824, 7.20998, 10.91452, 5.743856, 6.59342, 
    13.47913,
  39.17635, 22.23773, 13.06163, 17.83344, 17.48438, 12.3527, 11.97118, 
    5.203453, 4.915187, 8.222867, 9.967899, 8.556453, 7.747008, 7.040644, 
    14.66173,
  20.03617, 28.47845, 22.9596, 19.43888, 12.35705, 7.552725, 7.951385, 
    8.204475, 10.36616, 22.38078, 27.66355, 19.66032, 24.73537, 27.36381, 
    31.12869,
  36.33786, 32.88894, 24.07356, 17.29417, 11.96215, 10.47375, 6.214447, 
    4.58973, 6.385615, 14.19298, 24.66607, 12.97644, 8.538712, 20.45544, 
    24.3003,
  53.00218, 53.16099, 39.07163, 16.74723, 12.08408, 18.64069, 7.005366, 
    5.478376, 8.785187, 8.421756, 7.851758, 10.3525, 13.16957, 16.82614, 
    18.87516,
  70.74493, 70.52991, 58.09069, 30.03556, 12.2431, 20.63652, 16.11272, 
    10.27007, 10.24782, 6.869072, 4.841591, 6.570316, 14.98638, 19.75104, 
    11.69125,
  81.48768, 75.42994, 75.38001, 30.59463, 15.67185, 14.75722, 25.4605, 
    20.36999, 15.87502, 9.386223, 4.801088, 7.147267, 16.55444, 12.89338, 
    3.84858,
  67.9754, 74.98195, 64.1483, 28.48201, 17.92754, 16.86305, 16.5106, 
    19.93697, 17.25578, 17.30004, 13.91673, 10.50238, 14.71941, 4.784759, 
    0.9057176,
  54.70329, 68.24432, 50.05915, 19.93969, 22.77242, 23.77393, 15.28859, 
    13.2588, 15.61072, 14.75333, 4.612092, 13.49261, 12.33383, 3.117588, 
    1.396059,
  45.45616, 55.45109, 30.67289, 20.75136, 19.70855, 17.69798, 10.56267, 
    3.61329, 11.69045, 3.661052, 5.698514, 13.33938, 7.72693, 4.184271, 
    3.755773,
  40.57389, 36.65299, 16.23867, 15.14881, 13.25589, 10.88988, 11.23814, 
    2.641629, 2.408215, 4.397508, 11.70621, 7.958366, 4.879762, 5.678761, 
    8.886791,
  32.68651, 22.5894, 17.56008, 12.96997, 11.41831, 2.084443, 1.97507, 
    2.42297, 3.481315, 11.63773, 8.83126, 8.441237, 7.505974, 12.64687, 
    17.22169,
  12.3696, 11.43908, 16.33296, 27.32851, 29.44186, 26.45038, 18.19617, 
    14.5107, 11.6636, 12.78257, 12.2052, 14.1265, 17.96175, 20.27814, 37.82316,
  6.6684, 8.054525, 15.83793, 25.06632, 33.00315, 32.24537, 18.96839, 
    14.11455, 12.90941, 11.63466, 15.8978, 12.28305, 15.34391, 23.97062, 
    27.87721,
  4.965343, 11.8887, 27.70721, 22.52083, 22.62855, 29.97397, 21.65795, 
    13.96914, 11.10402, 9.861292, 10.0142, 10.54698, 10.48139, 8.413127, 
    16.50465,
  6.393619, 13.01903, 33.59111, 30.12408, 19.66498, 21.61675, 26.6084, 
    21.21212, 14.59842, 9.730254, 10.81234, 9.766061, 6.658182, 5.31481, 
    17.05374,
  6.100163, 11.4166, 31.31106, 19.88482, 17.46712, 23.29917, 25.78482, 
    16.13692, 12.89693, 12.20192, 8.947715, 8.696534, 8.267585, 5.919476, 
    2.787603,
  9.317011, 14.01189, 22.48755, 18.73844, 18.6737, 19.22013, 17.70699, 
    19.72077, 16.17925, 14.77545, 12.40693, 9.768432, 8.042312, 2.154536, 
    0.6904411,
  20.35775, 20.86621, 17.46413, 15.11347, 17.96159, 17.43948, 16.81113, 
    17.61609, 19.20505, 14.48639, 10.64581, 11.40744, 6.702174, 1.546048, 
    1.205845,
  33.50116, 27.61531, 10.99356, 13.38119, 14.7474, 14.79862, 15.79077, 
    16.2347, 16.48611, 11.5688, 12.98801, 11.10876, 6.545703, 2.791526, 
    2.983909,
  45.79203, 27.04623, 6.097048, 9.613022, 13.90335, 14.38704, 13.8635, 
    4.090816, 11.15982, 15.4584, 11.72145, 9.545033, 6.839579, 5.133961, 
    5.931625,
  37.89606, 19.62281, 11.10623, 7.032169, 10.89777, 11.18698, 5.749728, 
    3.454597, 15.48616, 17.56014, 10.52631, 10.93269, 10.71568, 10.4501, 
    13.09787,
  11.53955, 4.584304, 4.004596, 6.578456, 10.80242, 8.202847, 5.775881, 
    6.588036, 19.79609, 25.82554, 21.78052, 20.73399, 26.07714, 25.55074, 
    31.75487,
  2.56271, 1.916862, 3.355546, 11.77007, 16.01582, 10.97761, 5.641521, 
    6.829933, 15.49628, 14.55171, 15.7789, 10.77978, 7.997125, 21.44116, 
    24.06103,
  4.893883, 7.992308, 15.02233, 12.03758, 10.56381, 17.79942, 9.184389, 
    7.480519, 13.57949, 12.81813, 10.62761, 7.043021, 7.40087, 8.3178, 
    11.75899,
  5.914086, 9.519802, 20.79112, 21.24557, 5.641688, 12.31047, 23.06036, 
    12.16288, 13.7459, 15.1533, 12.0651, 6.243584, 5.965768, 7.41121, 9.280957,
  13.50502, 6.534273, 12.67628, 12.8139, 8.969102, 8.822799, 17.46134, 
    14.95861, 14.30583, 19.43762, 13.20758, 5.973072, 6.169975, 7.93812, 
    9.929553,
  27.25586, 10.96496, 3.45327, 7.58877, 13.01471, 14.15108, 12.51193, 
    15.73993, 17.46627, 18.12475, 14.70452, 8.165968, 6.391984, 8.470404, 
    11.57528,
  34.92734, 27.95017, 10.65139, 6.149621, 5.730191, 7.988264, 8.714106, 
    13.12014, 14.2493, 18.06724, 11.9866, 9.625648, 7.901898, 11.50998, 
    12.4963,
  41.62952, 33.36133, 11.67766, 10.24133, 6.294, 5.970921, 6.498485, 
    10.67491, 19.09879, 16.62603, 11.88993, 11.10848, 11.00591, 11.5806, 
    11.11769,
  50.97833, 39.90852, 10.63669, 7.109428, 8.186041, 6.260462, 11.02906, 
    4.084928, 16.882, 17.67501, 10.76051, 12.14578, 11.99203, 11.33028, 
    10.74888,
  38.0696, 31.41508, 15.99712, 8.613798, 4.974508, 8.807147, 12.19332, 
    6.282895, 18.51908, 20.70601, 13.57399, 11.98083, 11.72364, 11.57351, 
    10.61001,
  7.832784, 15.51733, 20.36206, 15.81406, 11.82652, 13.03029, 3.353928, 
    3.476107, 9.31391, 25.0873, 24.85071, 19.58102, 23.80264, 23.02835, 
    24.99666,
  18.63339, 24.91558, 25.88132, 15.16949, 21.17362, 14.92909, 3.293533, 
    5.060398, 4.38993, 21.21821, 20.02078, 14.6996, 16.61095, 22.44303, 
    23.11859,
  32.46791, 37.34135, 33.59319, 13.05697, 14.40037, 16.22461, 6.586367, 
    12.30525, 5.353866, 16.71501, 14.67529, 13.88341, 13.20163, 12.08605, 
    18.23815,
  48.22322, 47.82127, 37.6501, 18.5605, 4.24967, 9.665717, 17.65432, 
    12.36127, 8.119591, 18.18344, 15.31989, 11.97963, 11.03445, 10.65961, 
    13.55728,
  59.10706, 44.28194, 32.73224, 10.14074, 3.267872, 9.099473, 15.18804, 
    20.18185, 14.28772, 19.80173, 12.791, 11.30857, 10.91973, 8.573812, 
    8.353578,
  61.69434, 38.69693, 22.01244, 8.525206, 7.001395, 9.737794, 7.471753, 
    13.61797, 12.09812, 16.54107, 15.31004, 11.38784, 10.17301, 5.7992, 
    4.280759,
  70.92319, 55.34903, 30.35342, 11.14319, 9.207504, 13.70141, 15.1849, 
    17.76607, 9.497787, 14.41115, 11.77877, 10.13908, 8.086697, 4.005731, 
    2.899902,
  77.15557, 62.08293, 25.91095, 16.24067, 19.4165, 17.3907, 15.85449, 
    9.582596, 14.80202, 13.79603, 14.59609, 10.30972, 6.186405, 4.677367, 
    4.301747,
  74.45507, 50.45792, 19.07707, 16.43457, 18.4827, 18.74096, 11.53669, 
    12.19673, 15.20178, 15.90902, 14.19071, 8.074122, 4.971472, 6.439032, 
    3.90723,
  58.00768, 37.44032, 20.68603, 18.49792, 18.08877, 12.81313, 13.0739, 
    16.53733, 17.7355, 18.28947, 16.0418, 8.177767, 4.728948, 5.468945, 
    4.602667,
  20.67292, 26.56934, 23.47156, 7.825364, 9.216705, 11.70887, 6.522962, 
    6.608855, 11.71482, 25.25801, 23.74709, 20.79641, 16.18163, 15.19668, 
    16.94449,
  37.87484, 29.20663, 20.33151, 9.75684, 19.78157, 21.49301, 11.19969, 
    15.26942, 10.14338, 19.44829, 23.08555, 12.90732, 9.230033, 18.12941, 
    17.62198,
  44.79375, 35.39701, 29.74194, 17.28862, 18.40137, 23.56784, 21.528, 
    15.69101, 12.26848, 15.52848, 16.692, 11.41351, 10.13598, 6.100878, 
    9.381322,
  50.43176, 35.28436, 29.80159, 25.44327, 16.85144, 20.45393, 18.07369, 
    14.47473, 12.17739, 17.38238, 14.10551, 12.19654, 7.631859, 6.890477, 
    9.226314,
  51.28371, 32.61539, 30.50114, 17.97676, 15.38342, 17.7725, 18.80578, 
    12.11542, 10.13604, 22.32904, 13.51435, 11.2659, 8.259786, 9.657365, 
    8.75991,
  54.15301, 37.31388, 30.04454, 18.48675, 18.57289, 17.55347, 15.82106, 
    11.66006, 12.9175, 15.62854, 18.17707, 10.88723, 8.956675, 9.8673, 
    9.064577,
  58.7838, 45.51759, 28.29448, 17.20693, 19.59076, 18.28929, 17.01397, 
    15.92901, 12.30023, 13.85371, 14.23008, 12.43202, 9.744147, 10.75056, 
    7.833069,
  65.92616, 49.49175, 22.30115, 19.82412, 20.136, 18.26906, 18.30077, 
    17.79747, 13.94866, 13.12813, 14.78594, 11.93674, 10.24946, 9.705562, 
    6.696263,
  65.51857, 40.58012, 15.52067, 19.59216, 18.99566, 18.72129, 18.05757, 
    19.56, 16.56663, 16.17914, 12.83287, 11.98842, 10.56473, 7.074993, 
    3.998869,
  52.58772, 28.8831, 19.05426, 20.81444, 19.4239, 19.23461, 22.09691, 
    23.84362, 18.58982, 18.17477, 14.23201, 11.86255, 9.178358, 6.593968, 
    3.302645,
  13.30849, 21.23796, 24.67132, 15.3088, 18.35317, 19.88028, 15.53869, 
    14.23194, 14.17015, 19.9379, 21.18303, 19.68615, 25.08701, 24.61969, 
    23.32995,
  25.82377, 26.11526, 24.64007, 20.30181, 27.11903, 27.02014, 16.5522, 
    13.41188, 14.98052, 15.70827, 19.66776, 15.35845, 11.26658, 17.49016, 
    21.91789,
  33.23355, 31.54807, 31.22598, 24.42302, 20.28308, 23.47053, 22.38128, 
    14.69296, 10.37217, 11.12518, 13.53461, 9.407236, 8.566299, 7.120051, 
    10.81052,
  36.86235, 31.09943, 32.91282, 26.91268, 15.52146, 21.70727, 20.20762, 
    17.44453, 12.05737, 13.51574, 10.47309, 8.924372, 8.737784, 7.275603, 
    5.98844,
  35.9502, 29.2996, 35.50156, 21.71711, 18.94692, 16.87445, 18.99889, 
    11.15111, 9.965952, 17.23323, 10.87008, 7.404287, 7.618285, 6.613521, 
    3.796123,
  34.68417, 32.40396, 34.8422, 19.57869, 20.65826, 19.53238, 13.73627, 
    9.605035, 9.175706, 11.32212, 12.3243, 5.563505, 9.083276, 9.363367, 
    5.918387,
  34.07454, 36.35489, 30.04441, 16.78554, 21.34293, 22.45398, 15.47357, 
    10.09307, 9.242736, 7.870856, 7.475092, 4.55808, 6.775396, 11.27333, 
    9.387296,
  35.93103, 41.21257, 23.27297, 20.68091, 22.67832, 22.55381, 15.69433, 
    10.23979, 9.947652, 7.719276, 5.569939, 3.437488, 5.100147, 6.968444, 
    8.893247,
  38.32018, 35.99499, 17.95364, 20.43704, 22.16354, 22.1634, 16.62886, 
    10.7896, 8.216588, 5.688432, 3.743183, 3.451274, 4.23865, 4.790259, 
    6.495662,
  32.68859, 27.81971, 18.2824, 22.40644, 21.84753, 22.9868, 15.19622, 
    11.73853, 7.382404, 7.080549, 5.292193, 3.97531, 4.079859, 4.254381, 
    4.468119,
  12.65716, 19.09266, 20.42741, 18.08443, 17.49421, 23.57756, 14.20006, 
    15.07064, 13.9286, 18.381, 17.49862, 12.85396, 16.64833, 14.47728, 10.4122,
  21.38442, 14.22497, 19.57705, 20.17506, 28.21524, 30.47487, 15.38035, 
    14.08881, 10.45937, 15.36286, 17.39279, 13.39614, 11.76848, 16.8594, 
    12.75409,
  23.42347, 19.51081, 25.46827, 21.6217, 21.57245, 22.7147, 21.81214, 
    13.91344, 9.990849, 12.11442, 14.51061, 14.39674, 13.48238, 12.35741, 
    11.27421,
  23.96582, 27.09156, 32.99677, 26.34299, 16.50054, 16.36147, 16.93416, 
    19.34787, 13.18003, 11.21695, 12.42649, 13.68014, 12.3999, 11.70058, 
    9.590538,
  25.53042, 30.97597, 36.75995, 19.32753, 16.04509, 12.38972, 11.19022, 
    15.20962, 12.97391, 18.75768, 12.54016, 11.37887, 9.487269, 9.299488, 
    8.538425,
  29.48817, 36.75145, 29.6939, 16.32043, 18.08001, 12.13124, 9.284995, 
    8.157001, 12.18583, 11.75763, 11.66641, 11.1839, 8.900006, 8.312118, 
    9.749546,
  34.7758, 42.00829, 22.87277, 15.81701, 16.90415, 13.03114, 10.56665, 
    9.834696, 8.142509, 8.789031, 9.513555, 9.465465, 8.859795, 11.95677, 
    12.30939,
  39.1841, 42.68778, 18.21285, 16.27877, 14.29444, 12.23458, 9.763014, 
    8.693445, 6.974805, 7.533439, 8.496694, 7.560774, 6.406343, 9.254333, 
    8.491739,
  42.62754, 33.8363, 11.78592, 17.74451, 13.31945, 10.67335, 8.193717, 
    6.917278, 4.746682, 4.174281, 5.987788, 5.212744, 3.411124, 2.03503, 
    4.665701,
  35.34274, 21.28841, 12.82498, 12.73258, 9.706232, 9.897425, 7.9382, 
    5.57759, 5.027272, 6.562498, 6.732523, 4.949568, 4.570282, 3.297996, 
    4.968776,
  11.45366, 16.12818, 14.75826, 16.1904, 14.7556, 17.37564, 12.17195, 
    11.26358, 9.68688, 17.66843, 18.08853, 13.98657, 19.48891, 19.3997, 
    11.21605,
  20.99311, 13.71218, 15.04628, 10.45013, 17.66277, 16.71913, 10.87524, 
    10.31149, 7.954154, 9.381289, 15.92948, 13.24141, 12.05661, 19.75101, 
    14.34794,
  24.23281, 17.50524, 18.37535, 10.00453, 12.92319, 13.07283, 10.22563, 
    7.903003, 6.985473, 4.412628, 6.144569, 10.358, 14.00849, 11.37719, 
    14.97447,
  20.95485, 24.17999, 22.44075, 11.66926, 8.830606, 9.311252, 16.02546, 
    9.210466, 6.478034, 3.977426, 4.594916, 8.794719, 14.02353, 11.45328, 
    12.56751,
  21.18426, 20.98461, 24.36827, 10.13003, 9.071306, 6.336375, 7.501396, 
    16.09417, 8.870616, 5.534025, 3.455068, 5.809086, 11.5406, 11.23295, 
    9.376825,
  22.28147, 21.45984, 18.72859, 9.86979, 10.25688, 9.547702, 8.954923, 
    8.030606, 9.873892, 6.030709, 4.646739, 3.701274, 10.25914, 12.31763, 
    10.52681,
  23.69108, 25.22548, 16.37276, 10.5962, 10.04527, 9.059516, 9.092169, 
    7.391588, 6.600261, 5.06871, 3.252232, 2.692637, 9.81918, 12.52461, 
    11.3858,
  29.38786, 30.31938, 17.2303, 9.926304, 8.241608, 7.111389, 6.332052, 
    6.183444, 6.816782, 6.196041, 2.522084, 3.221595, 6.683255, 11.66881, 
    13.16361,
  30.90928, 22.9507, 13.73618, 10.10708, 8.513638, 7.491898, 4.591991, 
    3.204163, 4.091784, 3.576189, 2.249206, 1.76595, 7.914572, 12.22017, 
    16.71458,
  23.78051, 14.21439, 12.61454, 10.78679, 10.54564, 9.223216, 5.897304, 
    1.81244, 3.141726, 8.139982, 5.73622, 2.78832, 7.180003, 11.98434, 16.8078,
  12.59793, 16.16844, 16.95613, 10.37744, 9.640266, 12.65704, 9.316386, 
    7.648838, 6.018374, 9.917238, 11.74652, 11.52074, 21.05432, 12.74947, 
    12.03827,
  15.26968, 13.57114, 12.39008, 6.410087, 13.5642, 14.03222, 8.920505, 
    7.153737, 6.530887, 6.066822, 4.759065, 5.921249, 15.96259, 22.59629, 
    17.09501,
  17.16685, 16.93486, 17.228, 8.496033, 10.65351, 13.49787, 6.730052, 
    4.243608, 4.7362, 6.129112, 1.393678, 6.958644, 15.37743, 13.06019, 
    10.92783,
  18.59482, 24.24876, 22.19997, 9.311351, 6.807811, 7.972583, 9.773348, 
    4.527816, 3.60752, 4.649704, 2.253338, 6.364528, 13.20576, 10.67047, 
    6.796807,
  21.32894, 23.10221, 24.59882, 7.378776, 6.806607, 4.438812, 3.845809, 
    8.023428, 12.22868, 3.933055, 5.405038, 6.670119, 13.31397, 9.23491, 
    3.77979,
  24.11618, 25.44602, 18.16949, 6.039575, 6.07342, 4.34751, 2.055287, 
    3.773426, 7.676521, 6.883921, 7.023417, 6.204734, 10.28231, 7.74362, 
    3.757477,
  27.43529, 31.00689, 13.84078, 6.950288, 6.481699, 4.622325, 3.287326, 
    0.8166238, 3.86471, 6.400523, 4.453972, 6.201047, 9.759119, 8.785497, 
    3.788746,
  33.69465, 35.52215, 8.722841, 7.374172, 7.418831, 6.322882, 8.04504, 
    10.12555, 6.60309, 5.731563, 5.19681, 7.041472, 7.71761, 7.067934, 
    4.493373,
  37.76385, 26.87361, 5.932891, 8.455732, 7.83878, 5.963837, 6.089672, 
    5.945134, 4.643686, 2.931392, 4.923823, 7.317121, 6.949379, 5.574504, 
    5.618864,
  30.17533, 17.09498, 5.863369, 7.637957, 7.495755, 6.270376, 4.814365, 
    2.220619, 2.637145, 6.539342, 7.469469, 9.126403, 6.593007, 6.286835, 
    6.899699,
  8.567593, 8.54374, 11.60991, 8.809821, 6.463219, 4.694684, 3.118199, 
    4.554829, 4.938961, 13.16981, 20.76913, 17.68925, 11.21518, 6.963334, 
    18.65711,
  9.073732, 6.858302, 7.323031, 7.452482, 11.34568, 4.649961, 1.624207, 
    2.348645, 4.920642, 8.321856, 14.84152, 15.43055, 6.318294, 19.4824, 
    16.77904,
  17.23026, 12.32372, 11.82439, 9.421904, 5.940925, 12.0605, 0.9701228, 
    1.952663, 5.671446, 7.056015, 8.492096, 12.62367, 6.932196, 6.931204, 
    7.654322,
  21.03031, 17.18739, 15.47495, 9.122602, 2.462201, 1.334932, 9.274655, 
    6.079445, 6.518226, 8.740311, 10.29388, 12.41125, 10.70413, 7.750091, 
    5.19054,
  28.0431, 20.94212, 18.54416, 5.084989, 2.044286, 0.5183562, 2.76561, 
    16.14866, 11.95251, 12.49708, 10.71152, 10.09588, 4.802048, 4.573822, 
    3.3424,
  36.17215, 27.50083, 13.52403, 4.101087, 4.797705, 2.90161, 3.52921, 
    6.683604, 11.57076, 16.27847, 11.72391, 8.664233, 6.396163, 3.219908, 
    3.064304,
  43.53293, 35.93544, 12.05655, 5.407646, 9.240858, 12.76199, 8.693397, 
    7.724588, 12.74688, 11.68139, 9.741421, 7.975317, 6.907883, 4.416088, 
    4.241112,
  52.62262, 39.28727, 6.079081, 2.578453, 4.460957, 6.926306, 9.585596, 
    9.893123, 9.467938, 9.347692, 8.702761, 7.664449, 7.112482, 4.400968, 
    4.323438,
  53.3215, 25.04185, 1.701516, 2.553516, 4.256514, 5.598606, 5.230043, 
    5.810997, 7.383848, 8.333507, 8.098393, 7.48136, 7.368634, 6.481071, 
    4.161956,
  41.98786, 14.8224, 1.798173, 2.500151, 4.154589, 5.880167, 6.549618, 
    4.3556, 7.930732, 13.4674, 12.55373, 8.42775, 7.963671, 7.071848, 5.182355,
  8.43847, 7.665533, 19.88071, 9.763407, 10.03752, 14.71269, 10.40222, 
    5.305618, 3.518566, 3.665474, 10.76032, 13.36056, 13.35131, 11.49664, 
    22.79476,
  8.117264, 12.77052, 11.61935, 9.89972, 16.01373, 10.88831, 5.95015, 
    5.641889, 2.807858, 3.583671, 7.206583, 10.35769, 2.890402, 22.80975, 
    22.85273,
  25.01507, 24.54656, 19.42073, 10.72633, 12.14735, 14.23838, 1.60958, 
    1.069041, 2.324171, 6.153235, 7.152952, 8.237816, 2.862723, 5.197846, 
    12.03398,
  36.9651, 32.49099, 21.64933, 11.55575, 8.089209, 5.092065, 7.131207, 
    4.928314, 2.744088, 3.617429, 7.554918, 8.423433, 6.413783, 8.309758, 
    5.517326,
  49.56208, 34.19906, 20.4476, 7.032544, 5.251742, 2.332401, 1.401342, 
    16.55868, 14.35192, 5.109431, 8.35854, 7.839812, 6.082312, 3.829111, 
    1.024641,
  55.02913, 36.55446, 17.24504, 6.333887, 3.169244, 1.533851, 1.521407, 
    2.353135, 6.679894, 5.632481, 5.220919, 3.739607, 1.686807, 0.9042706, 
    0.1304474,
  56.03024, 40.75604, 15.68888, 8.435202, 7.486131, 6.761258, 5.075723, 
    5.890526, 3.451956, 2.805005, 7.477798, 6.840862, 1.95156, 0.324746, 
    0.1799474,
  56.14755, 38.93675, 7.823962, 5.055108, 6.762186, 6.302385, 5.413774, 
    4.075044, 3.129173, 4.802251, 3.689919, 2.447497, 0.5464733, 0.262604, 
    0.4411125,
  53.36199, 26.4929, 5.292786, 6.850948, 7.485744, 6.0667, 4.003783, 
    2.604974, 2.843986, 3.304838, 2.694281, 1.298547, 0.7589821, 0.3146514, 
    -0.4831513,
  42.62313, 22.25065, 6.053689, 6.281606, 9.234455, 8.198108, 5.054195, 
    3.270765, 3.753474, 4.240134, 3.295431, 2.387506, 1.245857, 1.191107, 
    0.4111509,
  0.27092, -6.511103, 12.57977, 3.142401, 7.620152, 11.35999, 9.535837, 
    8.258607, 7.638741, 17.2842, 20.19435, 20.10801, 11.55763, 22.70936, 
    27.23103,
  -6.559516, -3.844723, 0.9507602, 6.41038, 16.30573, 19.68503, 17.22047, 
    15.19635, 9.673306, 3.559365, 4.944147, 7.176188, 5.409062, 30.75132, 
    26.75849,
  3.789136, 9.56834, 11.5234, 10.89032, 17.99051, 23.17799, 16.17131, 
    13.9669, 9.551299, 9.324139, 7.544462, 5.833868, 9.058233, 10.26601, 
    14.2354,
  17.11131, 22.32162, 21.01638, 16.87139, 15.81982, 21.6705, 20.27513, 
    13.19993, 7.213296, 9.078578, 4.28314, 6.457832, 12.3142, 14.01498, 
    6.161561,
  38.06559, 30.03217, 26.80264, 16.93306, 15.14508, 15.64734, 14.16045, 
    21.88955, 11.85648, 8.061538, 12.20512, 13.64844, 13.25573, 9.246065, 
    2.079079,
  57.27669, 42.0735, 24.36302, 13.3057, 12.13509, 11.90827, 10.20605, 
    4.799886, 4.04516, 3.102105, 8.799254, 12.26587, 9.616983, 2.949789, 
    0.4056179,
  62.46306, 48.39338, 21.13881, 6.9421, 8.755397, 7.789361, 4.512269, 
    2.639557, 1.381663, 5.187835, 10.08951, 12.85209, 4.131297, 0.5724345, 
    0.2625961,
  50.91619, 38.01831, 6.057644, 6.655156, 5.888712, 6.328432, 6.99123, 
    4.113466, 11.07001, 8.820556, 12.46994, 5.824893, 0.6865296, 0.2165973, 
    -0.4525371,
  35.79502, 19.91251, 6.470825, 5.133379, 6.386581, 4.140378, 3.729975, 
    4.309793, 10.8088, 11.54966, 9.473263, 0.9354373, 0.3009413, 0.03633662, 
    -1.588324,
  25.22402, 13.55481, 5.664901, 7.885609, 6.487161, 4.715539, 7.400829, 
    6.608604, 6.513666, 6.266469, 1.130152, 0.3888564, 0.5788435, 0.2078911, 
    -1.290158,
  2.176733, -11.94272, -2.064931, -12.85594, -5.631726, -0.6703945, 3.36689, 
    7.764378, 7.405427, 21.56738, 32.53291, 21.48896, 18.76091, 17.52499, 
    19.58994,
  -11.76149, -19.53, -15.8799, -6.59666, -0.319781, 10.76974, 14.79476, 
    11.09446, 10.61356, 13.95864, 19.41393, 12.08405, 12.42151, 20.49573, 
    23.16228,
  -8.026366, -8.574936, -3.970496, -2.069314, 6.063198, 28.08202, 21.73236, 
    23.87115, 23.37977, 20.32949, 15.37259, 9.916632, 12.43165, 13.97595, 
    13.72614,
  -4.191896, -1.005988, 6.073674, 8.771507, 10.04778, 24.47206, 31.13068, 
    19.9914, 15.77109, 13.78772, 2.038789, 12.82538, 15.43475, 12.48019, 
    5.185595,
  4.15344, 5.329939, 12.05852, 10.34981, 15.48382, 19.07309, 21.47959, 
    25.93233, 14.82098, 4.654637, 4.924001, 15.09024, 9.293985, 3.350936, 
    0.4738207,
  14.22799, 16.50046, 11.43952, 10.15372, 16.98698, 14.14508, 11.67806, 
    10.38635, 6.599316, 3.963387, 13.6973, 9.349893, 2.988021, 0.3156215, 
    -0.06770415,
  29.50883, 32.5881, 13.77268, 12.02836, 15.33421, 15.8526, 11.82961, 
    11.98067, 7.254375, 9.445777, 12.0851, 3.813476, 0.4536389, -0.1702673, 
    -0.5165606,
  49.28839, 46.41393, 14.78599, 11.66315, 14.96009, 15.3588, 11.31803, 
    5.373975, 10.06064, 9.497027, 9.828887, 1.727405, 0.04080589, -0.4771863, 
    -1.148224,
  57.22205, 42.11052, 16.47914, 11.9228, 14.40946, 13.52595, 11.00788, 
    3.171258, 6.686672, 3.765622, 4.927526, 0.5580705, 0.04558711, 
    -0.3610503, -1.627018,
  46.07793, 34.28185, 19.59406, 13.2283, 13.46993, 13.88681, 12.32219, 
    3.953157, 3.2871, 8.18723, 2.476811, 0.1647802, 0.03880776, -0.1975633, 
    -1.219713,
  -4.147393, -16.43505, -8.412409, -22.57549, -20.28947, -20.83917, 
    -13.64951, -5.669203, -1.935385, 4.423413, 18.93797, 17.0504, 17.90084, 
    17.84129, 11.14418,
  -6.728379, -11.63503, -17.20167, -15.73976, -27.43173, -5.931147, 
    -3.980245, 0.3760605, 1.611362, 6.130231, 16.07107, 16.62704, 9.753775, 
    14.98515, 10.60901,
  -3.810333, -6.579579, -10.28077, -24.11864, -8.458549, 1.507776, 2.756049, 
    4.939929, 9.044388, 11.78728, 15.89195, 11.27222, 5.847999, 6.995395, 
    12.29089,
  -2.612548, -3.545375, -4.686307, -6.395066, -3.17565, 3.680776, 21.97365, 
    14.40767, 11.9733, 14.57472, 5.233856, 7.527257, 9.961079, 11.23799, 
    9.86907,
  -0.450873, -1.960051, -1.965988, -1.905984, 1.490436, 8.43507, 13.87844, 
    22.77344, 13.56278, 9.822192, 13.54012, 11.4395, 8.462229, 4.129997, 
    3.154752,
  1.40567, 1.87845, -1.675985, 0.6708002, 6.346532, 12.48333, 10.65854, 
    13.01593, 14.55803, 9.284698, 8.571388, 5.191796, 3.236097, 0.7122454, 
    0.168148,
  5.922332, 11.13159, 3.842421, 8.187355, 14.27789, 11.87077, 10.78079, 
    9.683919, 13.40759, 4.488038, 2.851832, 0.7511089, 0.009642864, 
    -0.04174066, 0.1857365,
  15.60959, 25.8763, 11.78597, 12.10393, 11.79495, 9.581464, 10.65352, 
    8.785681, 4.647746, 1.632388, 0.2516644, 0.02740831, -0.1512069, 
    -0.1471377, -0.1193526,
  33.96501, 34.75739, 16.51312, 14.10535, 14.2007, 12.41427, 7.451115, 
    5.228532, 3.13677, 0.7795125, 0.01119609, -0.08235431, -0.1590146, 
    -0.2159959, -0.6341516,
  39.84189, 40.30688, 28.80433, 13.10294, 11.09651, 8.883783, 3.653308, 
    4.147968, 3.442711, 1.072461, 0.5396932, 0.2718238, 0.03567366, 
    -0.1975774, -0.9022255,
  3.287091, -0.881871, 27.51654, -2.183754, -3.959461, -4.702731, -2.920518, 
    -3.616134, -8.624144, -9.706544, 7.091648, 8.903819, 9.983317, 3.681126, 
    0.577556,
  -13.81182, -4.384143, -5.04021, -2.563686, -3.14909, -3.952543, -1.672399, 
    -3.870835, -5.318893, -6.208678, 1.221637, 5.337231, 7.378316, 8.961232, 
    12.50447,
  -5.90799, -2.441995, -2.460402, -5.380542, -3.758126, -3.802741, -3.048175, 
    -2.185001, -3.525801, -4.839705, 1.316428, 6.466814, 7.080966, 3.94649, 
    12.57194,
  -1.243535, -2.196008, -2.334274, -2.454709, -3.257234, -3.248444, 
    -0.1002093, -1.241514, -2.487925, -0.2205251, 1.162407, 6.480269, 
    10.18091, 11.35482, 11.31944,
  3.40031, -1.290029, -1.912532, -2.69984, -3.134463, -4.013269, -3.584856, 
    3.769518, 6.325662, 3.296987, 3.480759, 5.219017, 9.113793, 12.00906, 
    11.28361,
  9.241507, 2.085858, -3.336339, -3.144201, -2.049419, -2.337677, -1.283809, 
    0.8323193, 4.39463, 4.805566, 6.125978, 7.371345, 11.6118, 11.06558, 
    7.069271,
  19.89216, 14.33745, 1.753858, 0.4094881, 1.201629, 1.897059, 3.730765, 
    4.741585, 4.223503, 6.698957, 10.0749, 8.997593, 6.110569, 2.920519, 
    3.21504,
  37.50039, 32.27234, 9.147055, 3.879104, 6.862293, 10.44909, 9.355798, 
    9.595165, 11.82243, 7.657557, 5.381583, 2.009965, 1.72818, 0.7947215, 
    0.8476912,
  50.80897, 37.15, 12.64318, 10.17547, 11.09916, 10.60829, 6.028713, 
    2.810813, 2.109066, 1.695677, -0.3852556, -0.08907128, 0.2018689, 
    0.1852647, 0.2244263,
  42.36637, 31.95621, 16.81948, 8.841791, 5.345426, 3.162478, -0.04323757, 
    -1.640614, -0.3480567, 0.3283378, 0.5309427, 0.7568015, 1.968741, 
    3.753271, 1.90594,
  1.618134, -1.517236, 12.90997, -2.480444, -4.166011, 2.074095, -5.584915, 
    -7.204406, -7.341968, -4.908231, 2.212737, 1.152159, -2.175275, 
    -7.254247, -7.004055,
  -3.4014, -1.047895, -0.5992566, -1.637504, -2.692073, -3.202607, -3.239207, 
    -5.743041, -6.805853, -5.357291, -0.6643443, -0.1504623, -3.279357, 
    -5.785015, -5.231091,
  -0.900268, 0.2019615, -0.9166107, -3.050785, -1.867096, 3.625702, 
    -2.231955, -3.990796, -5.200041, -4.115524, -0.2654918, -0.5696293, 
    -3.236187, -5.513299, -3.307013,
  1.461131, 0.8013729, -0.3709798, -1.38018, -2.712719, -2.423266, 1.744738, 
    -3.40626, -2.7525, -1.335583, 0.1915875, 0.8611104, -2.562902, -2.391075, 
    0.02924897,
  3.501828, 2.151463, 2.171224, 0.2129844, -1.212618, -3.228298, -3.460879, 
    1.146727, 4.053803, -1.177502, -0.3773208, -0.4197448, 1.194105, 
    0.7467458, 1.526878,
  5.512121, 4.387985, 1.682631, -0.4211909, -0.1271574, -1.196981, -2.35782, 
    -2.286447, -1.73646, -2.727347, -2.126389, 0.3950771, 2.099711, 2.584181, 
    3.126847,
  9.057566, 9.423124, 1.998252, -0.24812, -0.1746752, -0.2175261, -0.7720022, 
    -1.208753, -2.250012, -2.773932, -2.464443, 0.4393823, 2.233094, 
    2.445789, 3.892203,
  20.03704, 20.09097, 3.242338, 1.351097, 2.324919, 1.190645, 0.1569107, 
    -0.1916415, -0.1668031, -0.1539022, 0.5984135, 2.292394, 2.673942, 
    3.229424, 3.912124,
  31.84216, 18.44663, 2.727938, 3.663011, 5.152979, 5.169881, 5.079674, 
    3.87425, 4.15778, 4.960778, 3.778647, 4.002702, 3.438644, 2.961719, 
    2.943242,
  24.80987, 13.02645, 4.876582, 3.379474, 4.157284, 4.22691, 3.494306, 
    2.320263, 4.12432, 5.032837, 4.904339, 3.50572, 2.828811, 1.462783, 
    1.140365,
  2.568382, -2.596121, 8.570573, -5.118668, -4.721945, 0.6607445, -4.977848, 
    -4.663084, -8.345125, -1.705098, 0.9574661, -0.7383643, -6.538862, 
    -6.436327, -5.187077,
  -2.902987, -2.935104, -1.957354, -2.889476, -2.114466, -4.273256, 
    -4.901767, -3.316114, -4.807358, -1.078782, 0.07309422, -1.199392, 
    -5.147185, -7.051937, -5.69028,
  1.996934, 1.559474, -2.799943, -4.307089, -2.517916, 0.5357499, -3.586151, 
    -2.782742, -2.713039, -1.328678, -0.1220631, -0.997658, -3.10932, 
    -5.611347, -5.405341,
  14.25713, 9.599308, 1.71308, -1.954603, -3.804884, -3.965322, -0.4372431, 
    -1.119108, 0.1713382, -0.681069, 0.1047586, -0.8081093, -1.433064, 
    -4.52937, -3.968328,
  28.94054, 13.15469, 7.095647, -0.2457267, -0.6125674, -4.601802, -6.801643, 
    4.550839, 6.383392, -0.01305341, -0.1312148, -0.9366425, -1.22694, 
    -4.208678, -7.865159,
  38.1482, 18.91143, 4.587734, -0.448559, 0.5188038, -1.295475, -5.596124, 
    -3.946429, -1.569041, -0.9812122, -0.763137, -1.18053, -1.075576, 
    -4.057195, -5.118319,
  49.42927, 32.6926, 4.256866, -0.4377215, -0.1494677, -1.223195, -4.104236, 
    -2.516088, -1.823276, -2.613024, -1.697653, -2.070595, -1.338282, 
    -4.276621, -3.37804,
  62.1712, 44.80917, 5.470869, -0.187463, -0.2733428, -2.341252, -3.282762, 
    -2.42122, -1.503193, -2.516959, -1.532793, -1.220779, -1.51572, -3.41594, 
    -2.365286,
  65.83267, 42.83955, 6.482137, 1.375661, -0.3469162, -1.993552, -1.379088, 
    -1.732409, -2.350254, -1.473097, -0.09053844, 0.4488867, -0.6901276, 
    -1.429336, -0.3757206,
  53.48554, 45.80099, 18.06269, 4.552822, 1.247448, -0.3894298, -1.437979, 
    -2.167591, -0.7926521, 1.0949, 1.706068, 1.662898, 0.4684212, -0.3854696, 
    0.1347782,
  4.370932, -0.2933652, 15.5562, -1.687296, 1.555266, 8.639315, -0.620842, 
    -0.2518605, 0.3433947, -0.489108, 0.741977, -0.3047384, -2.731645, 
    -3.476835, -5.390506,
  0.5272417, 0.210528, 1.153733, -1.019843, 1.896788, 0.6059975, -0.3812947, 
    0.7386543, -0.1611501, -0.1405117, -0.1138449, -0.9939874, -3.176179, 
    -4.712854, -5.935759,
  9.996258, 11.28969, 3.945705, -2.339272, 0.4261184, 10.60312, 0.3518514, 
    -0.2829768, -0.6964426, -0.2461863, -0.02652877, -0.7551466, -3.123709, 
    -5.315659, -10.53403,
  16.17906, 10.87252, 2.680624, -1.08809, -2.214868, -0.516091, 7.380663, 
    -0.2553811, -0.7116102, -0.07407353, -0.2741981, -0.9006311, -3.036454, 
    -5.203269, -5.640512,
  20.93183, 7.236433, 2.780237, -2.737993, -1.865126, -2.094421, -1.671003, 
    5.687954, 0.665873, -0.1076209, -0.1618982, -0.9482761, -3.373237, 
    -5.821029, -10.65476,
  21.53263, 8.054493, -1.399553, -3.865861, -1.40637, -0.1199916, -1.198132, 
    -1.902223, -1.476877, -0.5008059, -0.2910959, -1.299072, -3.834513, 
    -5.113991, -4.951426,
  25.12779, 11.91291, -1.499601, -1.647411, -0.110359, 0.570036, -0.2249326, 
    -1.199457, -1.773692, -0.9520845, -0.6332188, -2.059633, -3.713712, 
    -4.51399, -3.364656,
  28.01296, 17.51425, 0.5690218, 0.3050317, 0.7706268, 0.8185801, -0.4677839, 
    -2.468702, -1.879398, -0.3395211, -0.6064557, -1.926551, -3.214951, 
    -3.538361, -2.385666,
  31.30964, 12.94045, -0.4800107, 0.9254051, 1.604352, 0.3346806, 0.1028297, 
    -1.364894, -0.9897463, -0.2549985, -0.5015321, -1.315123, -2.610837, 
    -2.467548, -1.351764,
  21.75926, 7.274612, 0.5833266, 0.6735986, 0.3994799, -0.3661033, -1.151212, 
    -1.617765, -0.7001847, 0.6856741, 1.029491, -0.5390769, -2.586189, 
    -2.567561, -1.143576,
  4.961019, -3.741922, 12.15192, -5.577336, -0.06927869, 10.2788, -2.494992, 
    -0.8770299, 3.133606, 6.66333, 14.64061, 9.800074, 2.721885, -0.9378346, 
    -5.696407,
  -1.388751, -1.752248, -2.675271, -3.609149, 0.2859588, 4.498477, -2.857816, 
    -0.8653633, 1.52646, 2.614123, 7.56446, 3.470303, 0.9466785, 2.277756, 
    -0.5204603,
  0.06245596, 0.8188241, -0.1726032, -1.99117, -0.1175397, 7.581586, 
    0.3096229, 0.3469546, 0.6365851, -0.008953806, 0.03940203, 0.7013723, 
    0.6766622, -0.2329917, -1.014353,
  6.785868, 5.597761, 0.6490819, -2.670347, -4.531491, -0.986557, 10.99856, 
    0.7463551, -0.4358957, -0.2834357, -0.2190783, -0.2648683, -0.446121, 
    -0.6802471, -1.434088,
  12.90467, 0.271493, -2.719458, -7.430377, -5.629338, -4.899491, -3.081442, 
    18.11914, 11.70194, 0.8121837, -0.1773949, -0.3862971, -0.5559577, 
    -0.9414378, -3.094242,
  6.098626, -2.163714, -7.101274, -8.2833, -3.734939, -2.398386, -2.59791, 
    -0.07981317, 2.189752, 0.3245837, 0.07819828, 0.5158659, 0.7062638, 
    -0.627423, -2.547356,
  5.265429, 2.555361, -2.890774, -3.141018, -0.7165102, 0.0165503, 
    -0.4281736, -0.4056712, 0.5321437, 1.515287, 1.861769, 1.533441, 
    0.03066877, -1.371265, -2.219371,
  11.04347, 16.88262, 0.08062627, -0.4689171, 0.4057806, 0.288435, 
    -0.02625695, 0.5484281, 1.161216, 1.438485, 1.327363, -0.1327724, 
    -0.8722254, -1.675361, -1.784606,
  19.71962, 8.440375, -0.1637067, 0.3618952, 0.6211592, 0.6524211, 0.9764083, 
    1.593054, 1.256098, 0.8284692, -0.08311597, -0.5290591, -0.7124225, 
    -0.1771235, 1.849451,
  11.64792, 5.99645, 0.7120039, 1.153446, 1.169413, 1.113409, 0.6578507, 
    0.970546, 0.3637429, -0.01730341, -0.4277106, 0.6841739, -0.2640811, 
    0.8092532, 3.407258,
  -6.510394, -15.31701, 1.961054, -13.0244, -6.378893, 1.214491, -7.847484, 
    -4.901417, -3.003342, 5.241614, 6.315066, 9.135105, -1.720091, 18.85284, 
    21.34775,
  -18.02115, -15.48446, -13.34642, -11.04692, -7.602328, 0.4856575, 
    -4.489831, -2.095825, -2.846231, 0.1213824, 0.3022175, -0.2988414, 
    1.849848, 12.51901, 13.87056,
  -7.46283, -8.11691, -6.669977, -7.854461, -10.67729, -6.875374, -2.499522, 
    -1.220233, -1.596684, -1.3816, 0.506507, 0.236023, 5.134251, 7.003892, 
    6.946075,
  4.480688, 0.9771051, -1.540044, -3.043377, -5.79477, -3.46904, 2.251105, 
    -0.06112325, -0.3379204, 0.08192348, 0.2369982, 0.2001999, 4.135747, 
    5.913376, 0.8909553,
  8.170977, 1.957807, -0.1829218, -3.552298, -3.224415, -3.591611, -2.301879, 
    11.20892, 9.153218, 0.4872573, 0.1716891, 0.1476424, 2.041971, 4.075759, 
    -0.9368622,
  3.883029, -0.6500434, -2.662431, -4.463251, -3.053229, -2.155818, 
    -3.162465, -2.057711, 0.8227919, 0.2456718, 0.1047777, 2.66573, 4.755736, 
    3.40956, 0.3994907,
  3.926039, 0.04416157, -4.160913, -4.806431, -2.670872, -0.3599988, 
    -0.4415034, -1.028124, -1.052249, -0.6456597, 0.7216188, 1.982564, 
    3.586776, 2.472512, 3.344979,
  5.359735, 3.328457, -4.001319, -3.48671, -1.295168, 0.1255034, 0.508114, 
    -0.1113415, -0.6757913, -0.1140023, 1.011501, 2.836309, 2.500785, 
    2.036186, 5.503997,
  8.942272, 0.482573, -4.118088, -2.009914, -0.9761952, -0.175398, 0.569286, 
    0.8816673, 0.4711385, 0.4948948, 2.528375, 3.749323, 1.597677, 1.274678, 
    9.258679,
  6.728158, 1.394776, -2.484859, -0.6612574, -0.1254686, 0.3334582, 
    0.4261035, 0.1094898, 1.148506, 1.611909, 3.614851, 4.7851, 0.6104379, 
    2.59492, 14.57372,
  0.7196451, -7.975822, 1.788806, -13.52189, -12.06292, -1.540429, -22.77229, 
    -20.27337, -24.04303, 16.21311, 27.46848, 35.91137, 18.73455, 26.42367, 
    28.38704,
  -2.808883, -6.730259, -9.289168, -16.8807, -3.391762, 3.390886, -15.21173, 
    -16.48242, -19.36222, -11.22038, 33.80491, 9.679727, 9.573145, 12.47537, 
    4.370908,
  2.39621, -2.761476, -7.002375, -15.27559, -18.6696, -8.115306, -9.732765, 
    -6.531509, -6.99083, 0.006729853, 4.095418, 6.661496, 8.220447, 3.899725, 
    1.242082,
  11.97808, 1.591869, -5.064059, -9.731519, -13.97282, -11.43167, -3.447256, 
    -2.808286, -0.09184116, 2.112268, 3.035111, 5.410489, 7.55987, 4.760764, 
    1.916755,
  20.35929, 1.680554, -2.522014, -9.650543, -10.15965, -10.2313, -9.224944, 
    1.483384, 8.324732, 1.424763, 2.403156, 4.311026, 7.475469, 4.958546, 
    3.091241,
  18.63408, 6.053243, -1.194522, -7.935789, -7.643531, -6.912182, -6.297842, 
    -3.692837, 1.55383, 1.424369, 5.593338, 7.16558, 7.856499, 6.732728, 
    4.248428,
  17.77586, 11.9261, -1.252705, -5.975002, -7.085229, -6.109332, -5.124907, 
    -1.572039, 0.4850074, 2.50162, 4.578179, 8.634604, 10.86388, 14.15976, 
    13.3607,
  9.408153, 11.9932, -1.577832, -3.974321, -4.550255, -4.256197, -4.034045, 
    -0.6024281, 0.4266132, 3.204192, 3.454881, 6.07896, 11.80489, 13.37578, 
    15.84409,
  5.484, 3.335207, -1.387841, -1.830346, -2.467685, -2.953318, -2.483973, 
    0.3707921, 2.12701, 3.073712, 3.285091, 10.10884, 12.1788, 13.36993, 
    15.38445,
  3.715487, 1.451608, -1.004882, -1.105026, -1.464176, -1.623545, -2.123924, 
    -0.5715244, 1.963288, 2.942073, 4.585232, 11.75314, 11.76991, 14.79094, 
    24.38748,
  8.913525, -4.832813, 7.379843, -7.861134, -6.450587, 5.39198, -8.418597, 
    -17.21495, -20.97104, -9.750216, 16.8848, 26.63933, 22.99306, 29.21691, 
    36.22585,
  4.433646, -3.537243, -4.559417, -8.405585, 1.188743, 3.248339, -8.11386, 
    -9.711308, -13.01089, -8.97878, 30.93805, 8.774287, 7.2017, 5.060055, 
    -2.822627,
  8.268579, 4.825289, -2.927293, -6.185205, -2.951226, -0.09429117, 
    -2.603833, -1.289596, -0.8430613, 1.75815, 8.418125, 6.46937, 3.816463, 
    1.27514, -0.5825682,
  10.62424, 9.361568, -0.564144, -1.647886, -4.880064, 0.5290795, 16.51892, 
    10.81944, 8.585541, 8.155952, 7.854924, 6.322414, 6.034249, 3.29258, 
    4.157983,
  9.342201, 5.206222, 0.7219942, -2.889077, -3.503483, -2.12873, 1.307153, 
    17.98591, 18.0468, 10.66394, 8.708093, 11.50746, 13.58808, 9.910909, 
    10.89845,
  7.802233, 4.798426, 0.3174669, -3.437843, -3.530456, -1.083366, 0.131695, 
    2.492949, 11.90897, 11.87201, 12.27939, 15.73624, 17.07198, 19.5732, 
    16.31425,
  9.932139, 7.244789, -0.1146751, -3.85762, -5.230115, -1.940581, 1.429135, 
    5.997375, 7.809036, 8.115857, 12.20801, 16.91963, 20.32936, 14.99215, 
    18.37665,
  13.48166, 8.334335, 0.6415507, -3.28511, -5.784317, -2.139428, 3.663082, 
    8.294794, 11.62337, 14.74791, 13.92714, 20.23915, 19.16507, 18.83818, 
    17.89914,
  7.398991, 2.388106, -0.9869002, -1.224225, -3.458616, -1.617141, 5.654819, 
    9.226244, 15.89609, 15.6636, 18.69997, 19.45505, 17.56504, 16.98893, 
    17.09458,
  1.955861, 1.421483, -0.5255864, -0.9233766, -2.11635, -0.6794155, 6.324466, 
    9.360941, 12.85096, 22.66145, 21.26464, 17.99607, 18.66988, 18.3579, 
    22.52423,
  1.823607, -7.424862, -0.5306619, -6.066421, -0.5010303, 6.832705, 
    -4.547318, -7.856984, -9.682257, 28.35961, 46.64796, 28.80054, 33.81112, 
    32.31298, 37.7214,
  -10.52345, -7.700259, -6.541845, -5.997666, 9.180605, 8.197957, -3.380248, 
    -4.969745, -6.704763, 2.871866, 34.66692, 7.026197, 4.22334, 1.490578, 
    24.86356,
  -8.573708, -3.408177, -4.62172, -6.580183, 1.438239, 2.733453, 2.345028, 
    0.1894218, -0.7344291, -0.6137437, 4.401941, 1.693473, 0.9741892, 
    3.318598, 7.211857,
  -2.789741, -0.1277146, -2.459475, -3.248973, -8.749462, -0.4514731, 
    12.1228, 3.943524, 2.371354, 1.178627, 1.719349, 5.246585, 6.156436, 
    8.758434, 11.66353,
  3.006144, -1.29037, -1.455726, -5.262969, -5.157847, -4.398675, 1.343606, 
    18.52932, 15.69339, 3.422828, 6.073114, 13.5303, 17.62062, 14.75958, 
    12.11916,
  10.74896, 1.516598, -2.619925, -5.864933, -3.948495, -1.815875, -0.4663392, 
    2.949514, 6.68213, 8.296587, 14.04507, 17.93691, 16.65638, 14.72441, 
    10.93813,
  18.88148, 11.34503, -2.939336, -6.129443, -5.736492, -2.664325, 1.07237, 
    6.437846, 8.173758, 13.42679, 16.53749, 16.63471, 12.99604, 10.62657, 
    10.67417,
  28.83554, 17.98674, 0.3963219, -4.058008, -4.695744, -1.562267, 6.762086, 
    8.354485, 12.48024, 19.83974, 21.76213, 16.23775, 13.99885, 11.14631, 
    8.991014,
  28.6098, 10.82287, -0.6754897, -1.58873, -2.538727, 0.9826137, 8.302863, 
    11.47318, 20.01523, 21.6957, 17.86072, 16.72904, 13.05962, 10.00964, 
    5.610795,
  10.91281, 7.539503, 0.3002036, 0.4381634, 0.5533805, 2.938266, 9.908482, 
    13.93829, 18.36466, 25.2371, 22.59456, 16.34921, 12.99226, 8.942054, 
    6.165766,
  0.7848945, -3.969067, 14.22741, -3.792446, -2.123493, 3.669206, -2.904385, 
    -2.620071, -2.836656, 14.80673, 22.91328, 20.06245, 25.65721, 25.55735, 
    38.41447,
  -0.06865742, 0.9734083, 2.214914, -1.154622, 15.30181, 15.40137, -2.966721, 
    -3.103048, -3.871713, -2.18565, 12.75625, 1.263929, 5.124371, 8.320986, 
    21.35743,
  7.763336, 7.728192, 5.26395, 1.170235, 9.881612, 4.311645, 2.328798, 
    -2.572324, -4.050494, -5.585428, -4.353901, -3.165191, 1.064748, 
    8.503724, 10.89388,
  12.23656, 9.172229, 5.54982, 4.196282, -1.213095, 3.422523, 5.798754, 
    1.745097, -2.295562, -2.691494, -4.339436, -0.7063295, 7.112795, 
    10.22341, 10.5215,
  13.4437, 8.952654, 8.825218, 2.953887, -0.9274853, -0.2582878, -0.6440387, 
    10.34611, 7.735928, -0.3244685, -0.3217371, 3.201384, 10.45978, 12.31378, 
    9.99943,
  21.8742, 15.22506, 7.161778, 0.4756709, -1.029266, 1.740473, -0.7809207, 
    -0.8335601, 3.344539, 1.035892, 2.862604, 8.211963, 12.15566, 13.72397, 
    6.381405,
  20.87677, 15.34555, 0.145182, -4.401241, -4.091627, -2.695747, 2.026048, 
    1.629185, 0.2587465, -0.09453507, 4.581776, 10.61447, 13.73082, 13.51032, 
    8.799782,
  26.34293, 19.61622, 0.2769983, -4.807573, -2.098816, -0.7529991, 3.270832, 
    1.324707, 1.422388, 4.459772, 11.1174, 14.27191, 17.6881, 14.06471, 
    7.875827,
  31.15336, 17.28388, -1.128138, 2.786368, 1.728991, 1.89824, 3.587909, 
    4.004873, 6.889225, 10.89959, 15.30687, 16.91752, 18.88024, 11.35239, 
    7.71986,
  17.32312, 10.85014, 5.331714, 4.0477, 3.220314, 2.584853, 2.285998, 
    6.068783, 12.29908, 21.19501, 23.4604, 21.53663, 10.65138, 4.472248, 
    3.273166,
  -8.33881, -26.73639, -7.368721, -17.25685, -9.783465, -3.308181, -6.853177, 
    -3.936876, -4.026717, 0.3659101, 3.289272, 0.3261576, 7.543603, 14.4277, 
    25.26306,
  -6.806745, -9.613958, -6.615369, -7.330701, 1.619755, 5.556858, 0.1866812, 
    -1.575225, -2.280411, -0.2513773, 8.268064, -2.512388, -5.256567, 
    2.164334, 20.80977,
  8.64445, 9.656073, 6.954939, 0.9523409, 14.06634, 10.94572, 7.997824, 
    4.587051, 0.2383371, 0.5554094, 5.314187, -0.6472102, -5.103109, 
    -4.246277, 7.286836,
  28.18335, 28.10563, 18.50261, 14.97068, 5.126372, 14.95205, 11.76986, 
    7.916452, 1.2917, 3.681133, 1.647254, 0.1138393, -2.321034, -3.10411, 
    -1.496851,
  30.29918, 19.09172, 13.66768, 7.418185, 2.963469, 4.164293, 9.972059, 
    19.05574, 17.18122, 11.05422, 5.389474, 2.885062, -0.3420689, 
    -0.04159615, 1.632408,
  16.99599, 10.32342, 4.663301, 1.310465, -0.2762043, 1.697331, 3.338262, 
    5.826775, 10.81302, 9.584039, 9.209884, 4.706831, 1.599326, 2.045308, 
    4.340075,
  14.72655, 10.35101, 0.7494168, -1.298427, -1.334536, -1.574034, 3.192336, 
    3.72525, 2.378798, 2.898558, 4.039817, 3.588994, 1.456439, 3.973973, 
    6.022289,
  15.30067, 17.55772, 0.7894796, -2.622365, -1.313092, -1.064893, 2.962818, 
    1.638352, 1.141721, 3.043295, 4.053462, 2.112511, 1.761644, 4.880716, 
    8.602533,
  29.34163, 8.492267, -1.835323, -0.6670473, 2.76162, -0.1499191, 2.660597, 
    3.105668, 3.722282, 4.642664, 4.159206, 2.222528, 3.404658, 7.478527, 
    11.55794,
  22.12076, 6.258693, -0.8654261, 3.618958, 4.111524, 1.738101, 2.601567, 
    3.140573, 3.77144, 5.254741, 3.464926, 2.9617, 7.056148, 9.90075, 14.37307,
  9.238822, -1.977131, 33.46371, -12.92393, -0.8452339, 15.64939, -13.9908, 
    -14.97009, -11.31151, 11.91844, 11.72806, -0.6240765, -3.833571, 
    -8.83894, -7.04667,
  6.539925, 4.817078, 5.291521, -0.2668762, 20.3019, 18.09372, -7.642107, 
    -9.77089, -10.78351, -7.152123, 15.13324, -4.373903, -9.255125, 
    -4.006677, -4.840841,
  13.89649, 15.36682, 11.90282, 3.50977, 12.00502, 3.631448, 1.885945, 
    -2.660469, -4.068412, -5.997673, 2.140496, -1.349802, -7.028554, 
    -6.012941, -5.322127,
  31.19027, 36.21841, 26.85789, 21.69637, 3.735967, 11.69305, 15.8055, 
    5.653892, 2.699015, 2.73543, 1.604863, 1.522021, -1.748002, -4.065564, 
    -8.17404,
  30.88286, 26.63219, 32.46252, 20.15965, 7.247006, 4.640059, 8.490844, 
    23.69977, 23.04271, 11.44888, 7.720527, 7.825537, 3.31733, -2.00496, 
    -4.81187,
  24.72655, 24.26026, 17.61006, 8.327372, 3.749499, 5.131712, 4.794313, 
    5.097372, 14.43544, 10.17342, 12.13079, 10.23781, 5.62372, -0.3780084, 
    -2.105638,
  25.06071, 25.52196, 6.527069, 2.516051, 2.239561, 1.206952, 3.804794, 
    5.973567, 5.024543, 7.014791, 8.177003, 7.507563, 3.713946, 0.5982996, 
    -1.412515,
  24.12355, 19.31301, 3.476383, 0.9271459, 1.979526, 0.5643875, 3.189697, 
    5.093317, 3.416073, 6.683426, 7.160124, 4.991545, 1.558648, -0.1091269, 
    -0.792808,
  24.96962, 8.480358, 1.095487, 1.212712, 2.570132, 1.37865, 1.843094, 
    1.792259, 1.929499, 2.708786, 3.345494, 3.150211, 1.799049, 2.617472, 
    5.518963,
  17.32657, 7.041561, 2.161425, 2.891604, 2.389544, 2.976708, 4.420714, 
    6.605948, 4.795909, 4.523962, 4.444817, 3.351276, 3.433466, 5.395309, 
    12.67421,
  8.176683, 4.39013, 24.44608, 3.649145, 9.109997, 23.75352, 5.936916, 
    5.431261, 6.643263, 47.60961, 64.00889, 43.54144, 41.92301, 54.65121, 
    68.27501,
  9.239959, 8.74648, 10.11596, 5.701909, 26.27587, 38.90144, 7.449889, 
    6.725286, 4.137291, 13.5461, 43.39012, 24.61184, 8.170327, 25.87747, 
    51.59131,
  11.08691, 14.3196, 13.2223, 9.062407, 24.04435, 24.67077, 19.60567, 
    5.634683, 4.068923, 3.133593, 7.022612, 4.897765, -1.590685, 0.7008803, 
    10.77965,
  7.385082, 11.06819, 8.646822, 15.90706, 7.163321, 25.90882, 27.5735, 
    9.732686, 10.01906, 7.607781, 3.009487, -2.095328, -2.109119, -1.44371, 
    -0.810066,
  5.352914, 3.905856, 10.14491, 10.99335, 5.014756, 5.325069, 14.37302, 
    20.48741, 20.69181, 25.94593, 0.9143617, -2.511562, -1.809568, -1.842431, 
    -4.16129,
  5.724074, 2.362977, 6.90307, 3.847674, 0.937763, 2.018652, 3.757603, 
    10.0189, 19.77493, 8.69044, 0.09365802, -2.098971, -2.250294, -4.620791, 
    -7.34976,
  8.251154, 5.822141, 1.678624, 0.6925921, 0.8616877, 0.663379, 1.742486, 
    6.980169, 7.22506, 1.045989, -1.044374, -0.9718026, -0.8049871, 
    -1.957145, -2.314036,
  8.969744, 9.617889, 2.958584, 0.3556725, 0.4008829, 0.4375352, 0.8221993, 
    3.376147, 2.672026, 2.176263, 0.3598864, -0.03429336, 1.076823, 1.413269, 
    2.143791,
  13.96972, 7.198673, 0.9808953, 0.7446783, 0.8219213, 0.05076753, 1.132325, 
    2.390825, 2.103014, 1.843581, 0.8458765, 0.7351642, 2.33972, 4.013792, 
    6.778584,
  13.45646, 7.547286, 1.443544, 1.865457, 2.58852, 2.262874, 2.055548, 
    1.926793, 4.46871, 2.576873, 1.833029, 1.732889, 2.93581, 6.044458, 
    9.873237,
  4.506999, -10.22814, 8.067893, -15.98898, -4.356371, 6.498027, -20.7647, 
    -16.6489, -11.91706, 14.51108, 39.19768, 28.58261, 30.40942, 36.1525, 
    40.45944,
  3.950778, -1.754772, -6.828906, -9.795281, 2.997719, 8.147234, -4.437273, 
    -7.836836, -7.2558, -2.590218, 31.45256, 15.48053, 6.947873, 25.48116, 
    31.66662,
  27.09618, 16.16483, 8.138242, -1.299516, 1.109827, 5.832611, 1.856849, 
    -0.6438173, -0.4476835, -1.426932, 3.673469, 1.357575, 1.879599, 5.35536, 
    16.11265,
  48.70646, 41.21472, 21.07233, 13.37549, 0.5159354, 8.865669, 14.33796, 
    4.187973, 3.463931, 2.285736, 1.179491, 0.503481, 4.201794, 2.254535, 
    4.432119,
  46.65388, 38.27852, 33.64263, 15.64253, 1.279682, 0.1819286, 10.45427, 
    21.21609, 16.51129, 12.40848, 0.436837, 1.518301, 4.691846, 0.6819993, 
    -0.6461402,
  42.67638, 35.75754, 24.11729, 9.936125, 3.324455, 2.435499, 2.591563, 
    6.678504, 13.65107, 2.64626, 1.50353, 1.289132, 3.95758, -0.2118194, 
    -0.0372581,
  39.21024, 35.15302, 13.06336, 5.142559, 4.495366, 3.246495, 2.497615, 
    3.756133, 1.955531, 0.7134006, 1.263049, 0.3553453, 0.8198212, 0.5087093, 
    2.1718,
  35.23779, 29.88943, 9.119534, 4.796242, 5.318569, 6.209036, 5.376902, 
    5.53428, 1.971709, 1.797473, 0.1412912, 1.130476, 0.6166385, 0.9243749, 
    2.118587,
  27.49733, 12.24176, 2.699387, 1.237874, 2.217479, 3.428419, 5.67979, 
    4.684037, 1.818129, 1.362694, 2.765263, 2.894587, 1.455687, 1.318004, 
    2.465881,
  14.18764, 6.343552, 1.54003, 0.8972808, 2.361634, 2.854987, 5.049872, 
    4.298646, 1.129951, 3.944123, 2.896188, 2.275786, 3.717991, 2.561419, 
    7.692593,
  8.783351, 1.126383, 23.01756, -1.937707, 1.775887, 19.35512, -16.20685, 
    -27.37823, -25.9231, 34.60514, 34.45422, 8.397607, 36.4497, 19.314, 
    23.42551,
  7.771636, 1.04784, -0.2747752, -2.083687, 19.26577, 23.31323, -5.776835, 
    -14.02988, -19.94863, -12.80137, 12.3482, -16.20202, -13.56606, 12.47261, 
    19.43627,
  20.65558, 13.81419, 2.3646, -1.813711, 8.062943, -7.389494, 4.030321, 
    -3.779794, -11.49664, -23.53679, -22.56152, -18.06847, -16.26453, 
    -4.884269, 9.375942,
  40.72685, 28.93652, 9.179901, 2.350774, -3.917563, 4.352758, -4.956683, 
    -2.558573, -2.972108, -7.650071, -11.63551, -9.892001, -6.422813, 
    -2.534236, 2.864623,
  47.7527, 35.34045, 20.7017, 4.370521, -1.762146, -6.23547, -8.841539, 
    -10.87386, -4.834126, 4.667333, -5.208932, -5.794597, -1.624799, 
    -2.075354, -2.877484,
  53.49956, 37.75536, 26.16868, 4.352927, -2.246194, -2.640651, -7.497859, 
    -11.30659, -1.633203, -4.593372, -2.170239, 0.3766364, 1.522682, 
    0.5809437, 1.541065,
  53.97865, 43.54718, 20.50882, 4.484638, 0.3834527, -1.512302, -2.594483, 
    -4.540064, -5.703581, -3.473988, -1.233123, 1.456524, 2.438689, 2.892722, 
    4.568296,
  46.09804, 41.54121, 21.10943, 6.824957, 4.014452, 0.9298733, -1.665851, 
    -1.330899, -0.3133865, 1.545753, 2.803083, 4.778214, 2.929793, 4.237814, 
    4.728462,
  28.83927, 24.12976, 14.74424, 7.134625, 4.56677, 0.9901208, 1.099582, 
    2.276677, 3.520186, 5.597912, 6.815044, 6.678042, 5.453163, 4.580159, 
    3.750945,
  10.30487, 10.90309, 12.81136, 9.480818, 10.27766, 6.7303, 4.113461, 
    4.08599, 6.768725, 10.22543, 10.97741, 9.166041, 7.741628, 5.715598, 
    5.558072,
  10.52706, 2.78742, 18.97212, -4.223643, -5.380854, 17.00726, -12.74882, 
    -19.61555, -18.60858, 43.26891, 42.82094, 21.05235, 32.08455, 22.11112, 
    28.02687,
  12.80201, 9.069369, 8.587251, -2.064568, 11.56094, 29.68324, -3.115581, 
    -6.792934, -8.531089, -2.33428, 23.08773, -17.63704, -18.41823, 19.38135, 
    19.3291,
  25.15624, 24.52324, 15.54976, 6.429242, 18.95042, -0.7031863, 2.099121, 
    -2.067811, -4.792751, -7.86342, -10.24642, -12.43825, -20.9724, 
    -21.75792, 4.59729,
  35.33384, 33.39656, 21.61065, 15.80776, 7.909419, 12.84857, 0.4394726, 
    -0.7197385, -3.179365, -2.126742, -5.53533, -9.155457, -9.762171, 
    -14.34985, -8.394619,
  29.31226, 29.4223, 26.77158, 12.55313, 5.077404, 4.618428, 5.009659, 
    1.025894, -2.15787, 7.827966, -1.437406, -5.000208, -7.457767, -12.14753, 
    -19.65412,
  23.01346, 22.85874, 22.4522, 7.543766, 4.824805, 3.819819, 3.130197, 
    2.440917, 6.160995, -1.053297, 1.450272, -3.108169, -4.296419, -7.330915, 
    -12.1799,
  23.33409, 20.96055, 14.28001, 3.243609, 5.476511, 4.435947, 2.740995, 
    2.799923, -0.03112328, -2.535302, -3.601331, -3.414121, -3.824174, 
    -4.765811, -7.510549,
  28.73964, 18.50184, 14.25554, 4.093978, 5.992056, 4.921709, 1.897567, 
    2.736612, 0.5687385, -1.080007, -2.278389, -3.424779, -4.216028, 
    -4.162303, -4.982609,
  21.01072, 12.20263, 11.06686, 3.953772, 4.415639, 3.538579, 5.104635, 
    3.650499, 1.090185, -0.4151069, -1.687569, -2.836921, -3.354527, 
    -3.699563, -3.996943,
  9.195654, 8.592856, 9.753042, 6.241288, 7.470234, 6.23734, 6.351833, 
    4.16122, 2.035437, 0.8293924, -0.5853801, -1.547162, -2.484562, -3.03952, 
    -1.405348,
  9.283569, -3.410382, 5.615557, -23.464, -21.67934, -3.122368, -34.43726, 
    -35.27478, -41.5448, 43.06903, 49.29275, 24.70841, 45.43052, 33.4975, 
    56.06009,
  17.22889, 5.883337, -3.667138, -20.82168, 8.323461, 10.87991, -19.19934, 
    -22.59401, -24.50782, -7.405065, 21.79525, -10.71526, -10.63696, 
    26.31244, 27.89314,
  30.59347, 31.56714, 16.15322, -4.68488, -0.6044971, -13.58458, -4.158158, 
    -14.16053, -23.97878, -21.81699, -15.63609, -10.55757, -12.30042, 
    -8.815045, 8.108763,
  45.94678, 42.88017, 29.51938, 18.23229, -3.893125, 2.882535, -7.892148, 
    -6.703981, -11.10495, -9.52961, -11.68421, -6.687077, -4.465934, 
    -3.365241, -6.540054,
  37.05422, 34.66357, 33.69257, 23.39899, 5.250989, -3.590583, -3.652255, 
    -11.59809, -0.1682653, 5.976543, -4.405666, -4.979277, -3.15614, 
    -2.588243, -10.09259,
  25.54669, 20.98624, 25.94023, 17.49182, 9.50454, 3.424869, 0.6869732, 
    1.029232, 6.89183, 3.416284, 8.653063, -1.583371, -2.19488, -1.622304, 
    -3.698783,
  21.57989, 8.574471, 8.679533, 10.20708, 13.5749, 11.7569, 6.29473, 
    5.949222, 4.871881, 2.677306, 2.553352, 0.02258587, -0.6158526, 
    -1.000627, -1.511764,
  22.92344, 5.135534, 2.257733, 7.150038, 10.27864, 10.80469, 7.731019, 
    8.088209, 7.866637, 5.67842, 4.86866, 1.736959, 0.3791873, -0.0527039, 
    -0.6186883,
  23.04024, 7.549012, 1.496955, 2.093375, 7.095438, 9.22483, 9.348203, 
    11.99685, 11.93049, 9.053237, 5.710979, 2.184231, 2.226788, 1.432367, 
    -0.1648342,
  8.95603, 1.92344, 0.2441549, 3.142718, 6.988429, 8.424383, 9.81767, 
    11.55296, 12.96915, 12.5936, 10.40464, 7.082684, 5.002551, 2.743082, 
    2.725956,
  2.410712, -1.942522, 34.81259, -1.026032, 4.479422, 8.826697, -25.92081, 
    -45.13406, -45.81044, 56.50392, 65.20866, 26.17739, 58.23304, 49.07625, 
    88.76222,
  1.012921, -3.085735, -2.081845, -1.831633, 49.20998, 14.17959, -14.89217, 
    -33.58331, -44.38448, -15.13541, 31.40061, -21.07058, -32.1925, 46.53978, 
    66.72239,
  17.87432, 5.234182, -1.080926, -3.288618, 17.43454, -12.34384, -3.049399, 
    -17.00998, -36.7803, -41.60369, -33.01459, -37.75272, -39.97875, 
    -25.42138, 12.82028,
  42.01719, 30.13895, 3.615799, -1.955472, -7.306231, 3.914696, -20.13835, 
    -4.906138, -13.41107, -18.59382, -30.23593, -33.26091, -25.67199, 
    -17.05147, -3.5565,
  57.28447, 39.15798, 21.80513, 2.129856, -2.835824, -14.59327, -14.67744, 
    -37.20589, -16.06759, 6.725023, -16.3041, -24.49639, -21.44041, 
    -14.42536, -17.04887,
  42.9108, 44.45652, 31.52642, 7.272937, -2.395375, -5.53306, -22.36517, 
    -24.69203, -8.065418, -7.273682, -1.704108, -18.32451, -16.8744, 
    -12.01433, -8.097999,
  44.73549, 48.08462, 23.39513, 11.76415, 1.937233, -1.918497, -6.015941, 
    -11.1264, -15.15309, -14.55598, -15.39582, -13.69446, -12.71925, 
    -11.42002, -8.506005,
  47.59138, 41.08615, 22.90215, 16.27361, 11.82917, 1.719893, -2.415322, 
    -6.070196, -9.575216, -9.562228, -9.917851, -8.155359, -7.878132, 
    -7.339599, -8.602995,
  39.75224, 17.15945, 10.61546, 10.40156, 11.87544, 7.054586, 0.3559759, 
    0.02567648, -1.740079, -2.486393, -3.184426, -2.594942, -2.509681, 
    -2.529807, -4.602253,
  17.2882, 6.963691, 4.373751, 6.11458, 13.06264, 10.11943, 5.796793, 
    4.038726, 2.831785, 3.058843, 2.845948, 2.245825, 1.537632, 1.087546, 
    2.153493,
  3.163681, -0.1148655, 16.6295, 1.171271, 7.523092, 28.04642, -0.6350574, 
    -6.44892, -1.986472, 61.31538, 67.60756, 28.82223, 71.03835, 60.8048, 
    117.3155,
  0.4266997, -1.239901, -0.7607331, 0.03691828, 45.90921, 44.75702, 
    -1.886162, -5.39238, -5.337804, 0.06183699, 35.64378, -23.01021, 
    -24.13087, 74.26709, 99.9277,
  11.38618, 6.223752, 0.07030962, -0.3423976, 25.90446, -2.157321, 6.360395, 
    -3.516978, -4.483541, -27.4613, -43.82153, -30.78769, -35.24909, 
    -16.18486, 25.83948,
  35.51102, 22.57857, 1.222785, 0.1991669, -1.926375, 21.04213, -2.757545, 
    3.64329, -5.087921, -15.85838, -37.54645, -35.80604, -30.18942, 
    -18.39124, -1.523378,
  47.31236, 27.80067, 12.70558, 0.3353549, -3.449059, -5.18259, 2.70359, 
    -8.581849, -7.744313, 8.406247, -21.22906, -26.85977, -26.70205, 
    -18.2919, -11.28847,
  32.04221, 35.67815, 18.69378, 2.596593, -1.679235, -4.249856, -9.39783, 
    -9.045596, 2.213144, -2.193112, -0.5193694, -24.27601, -21.40582, 
    -17.11897, -8.174153,
  47.4451, 46.19199, 13.86836, 2.355797, -0.5490658, -2.472077, -7.45305, 
    -8.834955, -11.89811, -12.45212, -17.61066, -22.10048, -19.10714, 
    -17.152, -10.82546,
  54.53809, 48.273, 17.82028, 7.294885, 3.240343, -0.1966553, -5.993449, 
    -9.500063, -12.88028, -13.2091, -12.92623, -17.27656, -17.22673, 
    -16.83039, -12.44643,
  39.80802, 30.93507, 14.84368, 9.561326, 4.210364, -0.5315881, -2.31308, 
    -5.476195, -9.662354, -10.68531, -10.56624, -12.48429, -15.01889, 
    -14.73772, -11.78287,
  19.04305, 20.01595, 10.29216, 12.6389, 12.96039, 3.330249, -1.163898, 
    -3.864909, -5.749431, -8.424107, -9.353343, -10.97929, -11.48853, 
    -11.4431, -10.56309,
  3.540786, 2.598935, 20.33898, 4.58819, 9.477996, 22.32166, -0.2980984, 
    -1.740566, -0.6259034, 44.81991, 71.325, 35.96699, 73.62505, 61.02653, 
    89.08531,
  -2.196887, 0.5748385, 6.423485, 6.067542, 27.71469, 32.77969, -0.2430129, 
    -2.374896, -3.34435, 6.964757, 54.98528, 3.930795, 2.536107, 71.66277, 
    83.79198,
  2.173014, 6.676159, 7.49361, 3.836789, 18.02339, 2.747216, 8.55291, 
    -4.103326, -3.547363, -7.251332, -10.31044, -0.1210544, -8.277349, 
    -7.599751, 29.61217,
  12.94779, 16.46464, 9.489152, 7.212506, 1.552138, 25.67267, 2.630281, 
    7.645096, -3.275418, -8.030193, -17.39736, -13.72806, -9.516129, 
    -10.58768, 7.164935,
  16.03372, 18.81012, 12.37054, 3.755628, -0.4116108, 0.3860964, 7.930712, 
    3.334033, -2.888928, 9.125685, -9.398604, -12.60598, -7.704383, 
    -9.378465, -12.77787,
  13.11731, 24.13904, 13.20375, 1.512056, -0.7079181, -0.6129923, -1.397547, 
    0.09489345, 6.022583, -2.712105, 7.291915, -11.49469, -7.417047, 
    -7.003356, -9.408215,
  19.98664, 34.66796, 9.789346, 0.663168, -0.0707467, -0.4841461, -0.8618392, 
    -1.736901, -5.254347, -14.89423, -13.26754, -10.3067, -8.892595, 
    -7.82117, -8.769135,
  26.58099, 38.34003, 13.43721, 2.702815, 0.6052585, 0.1962099, -0.645403, 
    -1.080709, -4.268177, -11.40062, -10.67041, -11.62847, -10.324, 
    -7.253909, -5.166348,
  21.11982, 27.81017, 12.85135, 4.696507, 0.4065037, -0.07641088, -0.1499249, 
    0.3359508, -2.341281, -6.727863, -7.326422, -10.14646, -9.608006, 
    -8.69521, -4.022734,
  13.95255, 20.6263, 13.53811, 11.23819, 4.998913, -0.1916883, 0.07556101, 
    -0.006485153, -1.726797, -4.27911, -5.636862, -8.301988, -7.717674, 
    -8.02482, -6.884194,
  8.505408, 1.166176, 16.31195, 3.944232, 9.397185, 20.27451, 6.197559, 
    7.199944, 4.202302, 63.24072, 58.96786, 27.24309, 35.79866, 46.43909, 
    101.4929,
  0.3098592, 0.1414336, 0.7613322, 3.546805, 30.74776, 31.30085, 6.439806, 
    5.847007, 1.075507, 15.122, 64.08773, 11.33199, -0.9736633, 45.02871, 
    93.32632,
  0.7079218, 0.3743495, 0.6271619, 3.503035, 22.84511, 19.48786, 14.54798, 
    4.167799, 0.7227295, -0.03574219, 19.52776, 12.37372, -3.98758, 
    -15.22787, 32.63584,
  2.256089, 0.5555296, 0.616933, 6.51719, 7.430949, 31.6597, 17.16877, 
    20.982, 1.510894, -2.899461, -2.079111, -0.3726342, -8.49329, -19.04408, 
    3.120905,
  1.144431, -0.7262238, 5.233365, 10.71468, 9.034482, 11.84904, 26.50241, 
    19.15721, 11.74655, 14.44099, -1.459586, -0.7497969, -6.451662, 
    -19.39128, -23.50856,
  2.549067, 1.955222, 8.933493, 8.542169, 8.64341, 9.599121, 6.412053, 
    15.22744, 19.93791, 14.46657, 9.833583, -0.3961217, -4.544941, -16.20538, 
    -20.33986,
  9.765165, 10.16125, 1.985384, 0.988703, 2.90216, 5.056383, 5.066834, 
    4.703452, 6.190238, 3.241025, 0.8515327, -0.1425847, -4.647602, 
    -13.85817, -17.24264,
  22.03675, 11.8261, 1.423945, -0.6912557, 1.301231, 4.363756, 2.021703, 
    1.714607, 6.796333, 4.380194, 1.7318, -0.3977358, -5.504348, -13.01643, 
    -13.88054,
  21.81513, 4.899354, 0.9547924, 1.943287, 0.359844, 3.254478, 3.635701, 
    4.16113, 6.328898, 4.138492, 1.742875, -0.9455946, -5.746451, -13.07666, 
    -11.81589,
  14.30136, 4.022938, 3.644439, 5.65098, 3.611544, 2.926721, 4.551373, 
    6.517334, 7.575497, 3.993905, 2.940333, -1.151662, -4.724422, -10.92478, 
    -12.09309,
  10.88333, 6.89333, 30.96664, 9.157907, 13.89038, 27.03804, 13.10994, 
    7.15241, 0.6930008, 20.6331, 30.57813, 28.976, 48.32071, 40.42844, 
    78.79162,
  2.301409, 2.080948, 3.263663, 5.422714, 33.87572, 38.09546, 7.688189, 
    10.0197, 1.285419, 4.929044, 33.32828, 9.196508, -1.386133, 43.92007, 
    70.78606,
  1.062887, 2.906348, 2.647925, 1.032501, 22.82162, 18.83229, 14.94208, 
    6.694458, 4.247019, 1.431376, 34.41257, 26.55839, 2.73777, -7.371563, 
    24.29827,
  1.730494, 2.4648, 2.507087, 2.413806, 0.9766299, 20.728, 17.03017, 
    19.64763, 6.472195, 5.219203, 4.886965, 4.176173, -3.976362, -8.193698, 
    7.090415,
  1.860116, 0.6143277, 2.028711, 2.264664, 2.236318, 3.907608, 17.50616, 
    17.85267, 16.97728, 22.0835, 5.834577, -0.5829059, -3.685256, -6.774089, 
    -10.03998,
  3.841636, -0.5401679, -2.494952, -3.160645, -1.005944, 2.722351, 4.574387, 
    11.08345, 19.22344, 23.03929, 25.51372, 2.938745, -2.210304, -6.128382, 
    -9.183692,
  14.11183, 1.813288, -4.664318, -5.208842, -4.192281, -3.129141, -0.1475298, 
    2.142887, 4.990086, 7.66396, 9.485415, 6.09054, -0.9041244, -4.713547, 
    -7.532806,
  26.96924, 8.116384, -0.7147879, -2.624593, -2.045427, -1.958331, -3.891532, 
    -3.574209, 1.590985, 8.16889, 9.527815, 7.722002, 0.7398774, -2.990683, 
    -6.139617,
  32.80539, 14.70591, 1.940143, 1.230729, 0.5720527, -0.07222234, -2.137377, 
    -0.5339401, 2.18285, 7.709863, 10.18138, 6.817613, 1.579942, -2.351955, 
    -3.897361,
  31.49116, 21.23027, 6.259309, 4.348137, 3.749676, 1.076126, 3.012861, 
    4.741405, 5.852178, 16.61294, 13.89794, 7.886201, 0.9961908, -1.809693, 
    -4.685159 ;

 huss =
  0.0007530822, 0.0008768799, 0.0009092166, 0.0009961284, 0.0008377059, 
    0.0006539731, 0.0006554869, 0.0006321146, 0.0006374769, 0.0003675956, 
    0.0003955099, 0.0004174119, 0.0002630356, 0.0002883163, 0.0001339794,
  0.0009561618, 0.0009128363, 0.0008647798, 0.0009378794, 0.0007641964, 
    0.000571433, 0.0005947688, 0.0005371174, 0.0005777993, 0.0005743248, 
    0.000425976, 0.0005255786, 0.0005168005, 0.0002419239, 0.0001384041,
  0.0009307395, 0.0008935601, 0.0008646884, 0.0008629375, 0.0007758569, 
    0.000447036, 0.0005087287, 0.0005155887, 0.0005337982, 0.0005408757, 
    0.0005119591, 0.0005206638, 0.0005404028, 0.0005288417, 0.0003520976,
  0.00113384, 0.0008631091, 0.0007961398, 0.000777832, 0.0007899554, 
    0.0006982922, 0.0002854749, 0.0004015622, 0.0005369425, 0.0004798827, 
    0.0004437493, 0.0004648793, 0.0004996103, 0.0005274226, 0.0004602039,
  0.001308236, 0.0009967769, 0.0007881733, 0.0007331111, 0.0007056717, 
    0.0007090645, 0.0006824931, 0.0002410056, 0.0002850571, 0.000307249, 
    0.0003930083, 0.0004322271, 0.0004758358, 0.0005212312, 0.0005475282,
  0.001277564, 0.001101121, 0.0008742156, 0.0007632893, 0.0007157979, 
    0.0006666422, 0.0006203346, 0.000634043, 0.0004587235, 0.0003683333, 
    0.0003368547, 0.0004292976, 0.000463269, 0.0005085627, 0.0005444105,
  0.001292239, 0.001102979, 0.0009468182, 0.0008127367, 0.0007604, 
    0.000716044, 0.0006858966, 0.0006329794, 0.0005738842, 0.0005391051, 
    0.0005011102, 0.0004579447, 0.0004766339, 0.0004995739, 0.0005359706,
  0.001269325, 0.001140613, 0.0009690849, 0.0008696977, 0.0007979057, 
    0.0007449095, 0.0007039802, 0.0006580271, 0.0006178524, 0.000594656, 
    0.0005557326, 0.000506365, 0.000502655, 0.0005263335, 0.0005416659,
  0.001244844, 0.001108353, 0.0009590478, 0.00087578, 0.0008185451, 
    0.0007577097, 0.0007120819, 0.0006731761, 0.0006527828, 0.0006173366, 
    0.0005922007, 0.0005354744, 0.0005365719, 0.0005552122, 0.0005691127,
  0.00120875, 0.001076314, 0.0009777534, 0.0009040253, 0.0008143926, 
    0.0007660507, 0.000730239, 0.0006923698, 0.0006145052, 0.0004795597, 
    0.0005147595, 0.0005403934, 0.0005401413, 0.000535469, 0.0005393531,
  0.0008980546, 0.001073442, 0.0007530436, 0.0007996496, 0.0007115795, 
    0.0006337609, 0.0006757569, 0.000664669, 0.0005938851, 0.000487438, 
    0.0006053591, 0.0006448331, 0.0005523701, 0.0005115941, 0.0003655333,
  0.0009984722, 0.0009372503, 0.0009599963, 0.0008575451, 0.0006437195, 
    0.0006573037, 0.000687752, 0.0006974107, 0.0006615157, 0.0005874933, 
    0.0006035316, 0.0006897251, 0.0006359905, 0.0004011344, 0.0003123115,
  0.001074921, 0.0009965914, 0.000949616, 0.0009052905, 0.0007076812, 
    0.0004398235, 0.0006716397, 0.0006833635, 0.0007061739, 0.000649713, 
    0.0006716747, 0.0006925944, 0.000664248, 0.0006261519, 0.0004388681,
  0.001036437, 0.0009981121, 0.0009270424, 0.0008431557, 0.0007757313, 
    0.0006916833, 0.0003898216, 0.0005880829, 0.0006791412, 0.0006300923, 
    0.0006466847, 0.0006645711, 0.000654576, 0.0006103413, 0.0004900293,
  0.0009850053, 0.0009462467, 0.0008758054, 0.0008179686, 0.0007526397, 
    0.0007389758, 0.0007264304, 0.0004323155, 0.0004583884, 0.0005554088, 
    0.0005839331, 0.0006172941, 0.0006310287, 0.0006179803, 0.0005850727,
  0.00100065, 0.0009398441, 0.0008752222, 0.0008142266, 0.0007571048, 
    0.0007260385, 0.0007007107, 0.0006955507, 0.0005986123, 0.0005738524, 
    0.0005592173, 0.0005869356, 0.0006149106, 0.0006228877, 0.0006070727,
  0.001049451, 0.0009741975, 0.0008805915, 0.0008200234, 0.000767327, 
    0.0007287167, 0.0007060217, 0.0006818941, 0.0006670841, 0.0007052703, 
    0.0006286543, 0.0005583372, 0.0005866491, 0.0006084851, 0.000592471,
  0.001070552, 0.001012136, 0.0009234792, 0.0008583146, 0.0008035842, 
    0.000737306, 0.0006885672, 0.0006683614, 0.0006711602, 0.000704921, 
    0.0006311021, 0.0005381237, 0.0005557536, 0.0005766152, 0.0005672105,
  0.001083633, 0.001032597, 0.0009645977, 0.0009015722, 0.0008255244, 
    0.0007754309, 0.000734996, 0.0007179205, 0.0007071889, 0.0006815303, 
    0.0006291486, 0.0005264693, 0.0005363925, 0.0005512457, 0.0005467192,
  0.001096405, 0.001044034, 0.0009823715, 0.0009309803, 0.0008686552, 
    0.000819184, 0.0007656894, 0.0007355547, 0.0006617467, 0.0005681547, 
    0.0005667752, 0.0005314429, 0.0005299909, 0.0005417115, 0.0005458943,
  0.00135655, 0.000957029, 0.0009171431, 0.0007683452, 0.0007847981, 
    0.0008719563, 0.0008990131, 0.0008399659, 0.0007519785, 0.0005911266, 
    0.0005688903, 0.0005197859, 0.0004917724, 0.0005261312, 0.000397647,
  0.00105266, 0.0009244414, 0.0008820223, 0.0008166908, 0.0008227486, 
    0.0008938395, 0.0008435775, 0.0007689197, 0.0007478251, 0.0007469565, 
    0.0006169259, 0.0006135405, 0.0006456155, 0.0004667959, 0.0003591249,
  0.001022252, 0.0009121695, 0.0008965994, 0.0008758614, 0.0007884059, 
    0.0005282015, 0.0008091156, 0.0007307418, 0.0008211561, 0.0007840539, 
    0.0007080858, 0.000688506, 0.0007019042, 0.0007336077, 0.0005690817,
  0.001037595, 0.000917552, 0.0009029151, 0.0009244372, 0.0009551837, 
    0.0008529504, 0.0004783327, 0.0007189242, 0.000844559, 0.0007809772, 
    0.0007529865, 0.000746544, 0.0007570798, 0.0007377694, 0.0006500371,
  0.001061363, 0.0009329103, 0.0009097412, 0.0009228921, 0.000979447, 
    0.0009935297, 0.0009780178, 0.0005340397, 0.0005798342, 0.0007495183, 
    0.000801663, 0.0008105797, 0.0007985095, 0.0007743195, 0.0007421008,
  0.001092793, 0.000962796, 0.0009194835, 0.0009393317, 0.000981658, 
    0.001031706, 0.001059151, 0.001062984, 0.0009285291, 0.000889072, 
    0.0008250752, 0.0008427274, 0.0008258965, 0.0008209722, 0.0007943487,
  0.001142343, 0.001037194, 0.0009523911, 0.0009400369, 0.0009724433, 
    0.001024681, 0.001104523, 0.001156345, 0.00117752, 0.001154777, 
    0.0009591159, 0.0008804561, 0.0008590887, 0.0008834685, 0.0008635087,
  0.001166665, 0.001084921, 0.001017527, 0.0009777739, 0.00098604, 
    0.00101646, 0.001080766, 0.001176205, 0.00124537, 0.001251715, 
    0.001027212, 0.0009111268, 0.0009123381, 0.0009668338, 0.0008624067,
  0.00117681, 0.001115904, 0.001056893, 0.001002287, 0.0009845035, 
    0.001015987, 0.00106609, 0.001157736, 0.001246354, 0.001265802, 
    0.001057588, 0.0009349418, 0.0009632639, 0.0009499122, 0.0007702274,
  0.001193253, 0.001137045, 0.001062313, 0.001022832, 0.001004515, 
    0.001004244, 0.001034052, 0.001115969, 0.001112094, 0.001008649, 
    0.0009774503, 0.0009476212, 0.0009797541, 0.0008969891, 0.0008073791,
  0.001627185, 0.001509548, 0.001357412, 0.001181064, 0.001317018, 
    0.001360065, 0.001155056, 0.0008835946, 0.0007219403, 0.0003829865, 
    0.0004272309, 0.0003292248, 0.0002595325, 0.0003015403, 0.0001728117,
  0.001619205, 0.00134769, 0.001134195, 0.001035277, 0.000908931, 
    0.001100016, 0.001314754, 0.001084897, 0.0008672302, 0.0006225342, 
    0.0004528249, 0.0004215558, 0.0004344355, 0.0002632265, 0.0001726813,
  0.001543007, 0.001241649, 0.001038922, 0.00100364, 0.001034016, 
    0.0006833803, 0.00130439, 0.001133973, 0.000982509, 0.0007315299, 
    0.0005624832, 0.0004503138, 0.0004284699, 0.000503736, 0.0003884511,
  0.001403165, 0.001116892, 0.001022387, 0.001012057, 0.00102764, 
    0.001341936, 0.0007136638, 0.001069162, 0.0009523394, 0.0006865243, 
    0.0005382542, 0.0004492979, 0.0004391255, 0.0004859319, 0.0004871878,
  0.001259651, 0.001033163, 0.001014809, 0.001016426, 0.001020862, 
    0.001243402, 0.001435786, 0.0006782218, 0.0005928428, 0.0005330672, 
    0.0005076898, 0.0004604468, 0.000481087, 0.0005415746, 0.0005476545,
  0.001170587, 0.001023674, 0.001020593, 0.001016725, 0.001017304, 
    0.001225119, 0.001474348, 0.001267614, 0.0008449564, 0.000723758, 
    0.000517319, 0.0005026202, 0.0005421782, 0.0005924528, 0.0005231393,
  0.001108071, 0.001009802, 0.001025058, 0.001023635, 0.001069359, 
    0.001267876, 0.001416581, 0.001269477, 0.001146613, 0.001043686, 
    0.000680681, 0.0005857383, 0.0006191225, 0.0006142892, 0.0005862893,
  0.001047952, 0.001011261, 0.001055091, 0.001086339, 0.001177726, 
    0.001345669, 0.001377834, 0.001321993, 0.001225931, 0.001125887, 
    0.0007595569, 0.0006781573, 0.0006688548, 0.0006475661, 0.0006368958,
  0.001017296, 0.001026587, 0.001121003, 0.001198748, 0.001313804, 
    0.001407519, 0.001367448, 0.001349563, 0.001296851, 0.001184901, 
    0.0008603281, 0.0007526244, 0.0007148192, 0.0007080482, 0.0006962098,
  0.0009922312, 0.001070923, 0.001206234, 0.001319489, 0.001392032, 
    0.001417328, 0.001398169, 0.001380107, 0.001271977, 0.0009811533, 
    0.0008374979, 0.0007975359, 0.0007816156, 0.000742277, 0.0007940147,
  0.001244931, 0.001500216, 0.001518027, 0.001651438, 0.001625377, 
    0.001482349, 0.001083796, 0.0005888687, 0.0004478158, 0.0002904466, 
    0.0002569427, 0.0002614844, 0.0002300165, 0.0002828164, 9.693115e-05,
  0.001584934, 0.001652695, 0.001691091, 0.001635522, 0.001549146, 
    0.001266933, 0.0008635756, 0.0006096173, 0.0004933051, 0.0003930131, 
    0.0002985082, 0.0003892836, 0.0004560337, 0.0002105278, 8.913482e-05,
  0.001648976, 0.001702621, 0.001676034, 0.001637538, 0.001684307, 
    0.0007899839, 0.000874568, 0.0006835842, 0.0005567619, 0.0004712873, 
    0.0004627351, 0.0004345903, 0.0004524546, 0.0005335872, 0.000291738,
  0.001720609, 0.001707252, 0.001646413, 0.001639671, 0.001775707, 
    0.00139257, 0.0006251337, 0.0006531405, 0.0005855231, 0.0005366409, 
    0.0004771214, 0.0004510333, 0.0004884864, 0.000519788, 0.0003997945,
  0.001762109, 0.001710972, 0.00161092, 0.001591451, 0.001693794, 
    0.001697783, 0.001229759, 0.0005217785, 0.0004206049, 0.0004834959, 
    0.0004714851, 0.000477387, 0.0005233486, 0.0005751593, 0.0006096233,
  0.001765804, 0.001701539, 0.001576418, 0.001536617, 0.001578487, 
    0.001684929, 0.001532269, 0.001232063, 0.0007983778, 0.00065925, 
    0.000499821, 0.0005090066, 0.0005520935, 0.0006098123, 0.0006266892,
  0.001803496, 0.001676399, 0.001534792, 0.001493325, 0.001488797, 
    0.001624539, 0.001570885, 0.001323628, 0.001168588, 0.001017788, 
    0.0006608014, 0.0005387455, 0.0005938174, 0.0006497502, 0.0006695391,
  0.001819151, 0.001646176, 0.0014741, 0.001451923, 0.001467006, 0.001626738, 
    0.001548359, 0.001329417, 0.001240335, 0.001076151, 0.0006604787, 
    0.0005730179, 0.0006407145, 0.0006896465, 0.0007292586,
  0.001788189, 0.001579517, 0.001432194, 0.001430467, 0.001530756, 
    0.001678904, 0.00149353, 0.001309232, 0.001239069, 0.001096383, 
    0.0007117121, 0.0006164405, 0.0006933659, 0.0007289145, 0.0007595762,
  0.001690051, 0.001488864, 0.001415162, 0.001478484, 0.001611821, 
    0.001688063, 0.001448498, 0.001311227, 0.001169003, 0.0008710331, 
    0.0006851083, 0.0006731757, 0.0007302076, 0.0007467864, 0.0009168799,
  0.00088528, 0.001201036, 0.001079171, 0.00125862, 0.001014239, 0.001034869, 
    0.0009659665, 0.0006281153, 0.0004475539, 0.0002527351, 0.0002212355, 
    0.000376318, 0.000362545, 0.0003735471, 0.0001366704,
  0.001296363, 0.001383019, 0.001416203, 0.00146578, 0.001206658, 
    0.001146873, 0.000894357, 0.0005875426, 0.0004556496, 0.0003573807, 
    0.0002785535, 0.000474667, 0.000610749, 0.0003192766, 0.000151656,
  0.001364552, 0.001452958, 0.001496675, 0.001574523, 0.001456165, 
    0.0009470491, 0.0008003141, 0.0005728637, 0.0004803931, 0.0004580799, 
    0.0004601229, 0.000506894, 0.0006509511, 0.0006714613, 0.000356046,
  0.001441461, 0.001504462, 0.001556391, 0.001672607, 0.001727208, 
    0.001317889, 0.000594279, 0.0005274338, 0.0004936859, 0.0004924979, 
    0.0004695536, 0.00052552, 0.0006918043, 0.0006787174, 0.0004769487,
  0.001558232, 0.00156873, 0.001619871, 0.001735362, 0.001832251, 
    0.001683983, 0.001125137, 0.0004301983, 0.0003278341, 0.0004281811, 
    0.0004725989, 0.0005441894, 0.0007414487, 0.0007703389, 0.0007549651,
  0.001662471, 0.001665466, 0.001681468, 0.001796095, 0.001886602, 
    0.00177396, 0.001537758, 0.001216602, 0.0008166729, 0.0006324744, 
    0.0005109624, 0.0006097996, 0.0007381557, 0.0007931156, 0.0008247024,
  0.001735576, 0.001728542, 0.001744724, 0.001861559, 0.001903245, 
    0.00177547, 0.001584364, 0.001368414, 0.001118225, 0.0009636085, 
    0.0007170626, 0.0006543247, 0.000766579, 0.0008115225, 0.0008470005,
  0.001842155, 0.001794712, 0.001820874, 0.001917504, 0.001934704, 
    0.001770031, 0.001569013, 0.001341478, 0.001213365, 0.001072069, 
    0.0007431243, 0.0006946061, 0.0008016748, 0.0008381997, 0.0009229468,
  0.001903303, 0.001878514, 0.001899447, 0.001982551, 0.001950409, 
    0.001769725, 0.001554188, 0.001342279, 0.001222701, 0.00110814, 
    0.0007905091, 0.0007411053, 0.0007933188, 0.0008469958, 0.0009073482,
  0.001927466, 0.001914913, 0.001925961, 0.002005461, 0.001962456, 
    0.001789356, 0.001523918, 0.001323816, 0.001178437, 0.0009667049, 
    0.0007902536, 0.0007792472, 0.0008167436, 0.0008544762, 0.0009759422,
  0.000772438, 0.001163808, 0.0010059, 0.001219889, 0.0006638478, 
    0.0005627173, 0.0006315805, 0.0005536226, 0.0005698404, 0.0004648798, 
    0.0004917078, 0.0006475924, 0.000390827, 0.0002845594, 0.0001847626,
  0.00133039, 0.001358878, 0.001353296, 0.001324019, 0.0007065058, 
    0.0006569041, 0.0006965324, 0.0005668725, 0.0005829588, 0.0006339918, 
    0.0006075518, 0.0007922468, 0.0007004802, 0.0002596571, 0.0001687422,
  0.001467045, 0.001414186, 0.001396409, 0.001387421, 0.0009642097, 
    0.0006303654, 0.0006942466, 0.000579554, 0.0005710205, 0.0006404648, 
    0.0007308832, 0.0008222234, 0.0007878378, 0.0006394278, 0.0003634478,
  0.001588381, 0.001502888, 0.001453981, 0.001459778, 0.00140206, 
    0.001051989, 0.0006071811, 0.0005456786, 0.000593778, 0.0006425751, 
    0.0007123311, 0.0008540399, 0.0008345716, 0.0006993202, 0.000474708,
  0.001676755, 0.001584322, 0.001518958, 0.00153641, 0.001477903, 
    0.001331103, 0.001025055, 0.0003863266, 0.0003047553, 0.0004963411, 
    0.0006873384, 0.0008411941, 0.0008748884, 0.00080411, 0.0007477585,
  0.00174588, 0.001662803, 0.001574419, 0.001575332, 0.001535129, 0.00145588, 
    0.001288368, 0.001224113, 0.0008843751, 0.0008195325, 0.0006759848, 
    0.0008405477, 0.0008459722, 0.0008404177, 0.0007752199,
  0.001857922, 0.001750271, 0.001636379, 0.001625334, 0.001595527, 
    0.001502593, 0.001352495, 0.001204588, 0.001052843, 0.001021997, 
    0.0008472624, 0.0008264109, 0.0008687042, 0.0008616764, 0.0008023459,
  0.001958499, 0.001826381, 0.001703547, 0.001656095, 0.001649977, 
    0.001531689, 0.001452415, 0.001382723, 0.001226002, 0.001084211, 
    0.0008751647, 0.0008399083, 0.0008875154, 0.0009009796, 0.000876707,
  0.002021183, 0.001890926, 0.00178963, 0.001697908, 0.00167827, 0.001593973, 
    0.001539589, 0.001564428, 0.001370621, 0.00113467, 0.0009251445, 
    0.0008383736, 0.0008766534, 0.00092754, 0.0009199308,
  0.002033893, 0.001893284, 0.001803636, 0.001733431, 0.001705684, 
    0.001635366, 0.001647215, 0.001738247, 0.001509409, 0.001231084, 
    0.0009567636, 0.0008677692, 0.000840957, 0.0009351274, 0.0009560644,
  0.0008458176, 0.001190368, 0.0008845752, 0.001084112, 0.0006570603, 
    0.0005646124, 0.0006926673, 0.0007068245, 0.0006670813, 0.0004240672, 
    0.0003271729, 0.0003047152, 0.0002451753, 0.000259932, 0.0001568898,
  0.001496093, 0.001510897, 0.001399384, 0.001277391, 0.0006873483, 
    0.0005112923, 0.000702277, 0.0007348695, 0.0007319978, 0.0006415503, 
    0.0004539293, 0.0004806627, 0.000463364, 0.0002150851, 0.0001551139,
  0.001680422, 0.001684084, 0.001515253, 0.001398753, 0.0009546456, 
    0.0004645502, 0.000714039, 0.0007344856, 0.0007861954, 0.000744412, 
    0.0006692006, 0.0006173963, 0.000581963, 0.0005312226, 0.0003779555,
  0.001756507, 0.001748445, 0.001622341, 0.00150387, 0.001328078, 
    0.001041593, 0.0003740854, 0.0007271524, 0.0008317417, 0.0008160004, 
    0.000748889, 0.0006856118, 0.0006400816, 0.0005952384, 0.0004971575,
  0.001724403, 0.001799866, 0.001673218, 0.001536297, 0.001412271, 
    0.001253327, 0.001062977, 0.0003586949, 0.0004535542, 0.0007161964, 
    0.0008431548, 0.0007507892, 0.0007203926, 0.0006607264, 0.0006330814,
  0.001756601, 0.001826778, 0.001701048, 0.001573465, 0.001473585, 
    0.001294467, 0.001117284, 0.00111505, 0.0009746728, 0.0008537669, 
    0.0008141619, 0.0007889356, 0.000736739, 0.0007158141, 0.0006783006,
  0.001839038, 0.001846468, 0.001727474, 0.00162604, 0.001505711, 
    0.001366977, 0.001152952, 0.001121571, 0.001153011, 0.001043601, 
    0.0008733693, 0.0008198628, 0.0007661768, 0.0007316038, 0.0007075011,
  0.001937845, 0.001903498, 0.001797273, 0.00168416, 0.001550114, 
    0.001467586, 0.00123796, 0.001159139, 0.001213907, 0.001135179, 
    0.0008790755, 0.0008391079, 0.0008001305, 0.0007523518, 0.0007066864,
  0.002128603, 0.001998359, 0.001866944, 0.001771548, 0.00163725, 
    0.001559009, 0.001366663, 0.001207929, 0.001248538, 0.001188893, 
    0.0008963486, 0.0008594687, 0.0008102524, 0.0007735668, 0.0007376147,
  0.00240006, 0.002104545, 0.001973284, 0.00186841, 0.001720868, 0.001640318, 
    0.001467237, 0.001302073, 0.001296729, 0.001149365, 0.0008986455, 
    0.0008806097, 0.0008392516, 0.0008358302, 0.0008460688,
  0.0009499397, 0.001149502, 0.0007682691, 0.0009003985, 0.0005971981, 
    0.000568375, 0.00050288, 0.0004347326, 0.0004046461, 0.0002776233, 
    0.0002694313, 0.0003518319, 0.0002644564, 0.0002780122, 0.0001469581,
  0.001342832, 0.001474158, 0.001364417, 0.00119469, 0.0006357197, 
    0.0005701555, 0.0005671176, 0.0004952668, 0.0004546067, 0.0004283974, 
    0.0003414695, 0.0004923914, 0.0005315549, 0.0002249122, 0.0001758391,
  0.001423813, 0.001612327, 0.001540148, 0.001368562, 0.0008749946, 
    0.0004309369, 0.0006135506, 0.0005655137, 0.0005074158, 0.0004902874, 
    0.0004987904, 0.000530626, 0.000566921, 0.0005664405, 0.0004686276,
  0.001488455, 0.001662728, 0.001623156, 0.001500361, 0.001250613, 
    0.0009569713, 0.0004500638, 0.0006042387, 0.000532969, 0.0004999242, 
    0.0004968515, 0.0005274737, 0.000598839, 0.0006075615, 0.0005892752,
  0.00159126, 0.001716183, 0.001638218, 0.001518766, 0.00137599, 0.001248318, 
    0.001010921, 0.0004574817, 0.0003843172, 0.0004663018, 0.0005309322, 
    0.0005534811, 0.0006127105, 0.0006598222, 0.0006762806,
  0.001679538, 0.001758969, 0.001666014, 0.001550281, 0.001415143, 
    0.001316036, 0.001245789, 0.001186371, 0.0008895199, 0.0007372125, 
    0.0006253528, 0.000607106, 0.0006345148, 0.0006927265, 0.0007001914,
  0.001762336, 0.001824967, 0.001684023, 0.001551474, 0.001418927, 
    0.001337155, 0.001294001, 0.001299163, 0.001194505, 0.0009966001, 
    0.0007740417, 0.0006804593, 0.0006741179, 0.0007082425, 0.0007342691,
  0.001853498, 0.001842372, 0.001702707, 0.001551111, 0.001408467, 
    0.001363692, 0.001323492, 0.001366799, 0.00132725, 0.00120011, 
    0.0008475368, 0.0007592109, 0.0007294266, 0.0007415477, 0.0007675747,
  0.001802848, 0.001869602, 0.001728557, 0.001585005, 0.001447891, 
    0.001399313, 0.00134403, 0.001365151, 0.001402971, 0.001252707, 
    0.0009403671, 0.0008329428, 0.0007623697, 0.0007690038, 0.0007539341,
  0.001868906, 0.001863841, 0.001764924, 0.001634837, 0.001485711, 
    0.001445699, 0.001384234, 0.001382799, 0.001437627, 0.001259611, 
    0.0009653283, 0.0008624629, 0.0007916858, 0.0007723793, 0.0007599458,
  0.0006798884, 0.0009273534, 0.0005796482, 0.0006608103, 0.0004814486, 
    0.0004714799, 0.0005278075, 0.0005502158, 0.0005886609, 0.00045812, 
    0.0004042562, 0.0005589795, 0.0004087429, 0.0003560864, 0.0001946153,
  0.001176487, 0.001217431, 0.001106654, 0.00098748, 0.0004817574, 
    0.0004257961, 0.000531052, 0.0005457469, 0.0005764399, 0.0006147923, 
    0.0004663036, 0.0007179814, 0.0007537344, 0.0003987499, 0.0003305572,
  0.00138231, 0.001364927, 0.001269183, 0.001169216, 0.0007256914, 
    0.000329046, 0.000513851, 0.0005435139, 0.000555283, 0.0005686608, 
    0.0006163557, 0.0007253342, 0.0008122339, 0.0008388328, 0.0006753516,
  0.001476959, 0.001448341, 0.001373286, 0.001281204, 0.001096852, 
    0.0008199436, 0.0003577206, 0.0004773551, 0.0005557741, 0.000553521, 
    0.0005882949, 0.0006964356, 0.0008280664, 0.0009100551, 0.0008928301,
  0.001586157, 0.001521092, 0.001416144, 0.001337198, 0.001202348, 
    0.00111714, 0.0009070458, 0.0002796284, 0.0003022251, 0.0004461132, 
    0.0006012633, 0.0006826049, 0.0008393758, 0.0009476088, 0.001038018,
  0.0016845, 0.001584252, 0.001488847, 0.001426884, 0.001287733, 0.001214396, 
    0.001114098, 0.001043793, 0.0008507161, 0.0007033524, 0.0005808385, 
    0.000685019, 0.0008334256, 0.0009559054, 0.001054576,
  0.001782312, 0.001677385, 0.001535428, 0.001463733, 0.001377879, 
    0.001301077, 0.001213597, 0.001089582, 0.0009625062, 0.0008288816, 
    0.0006907607, 0.0007047806, 0.000842174, 0.000958983, 0.001076277,
  0.001884768, 0.001778794, 0.001622893, 0.001542567, 0.001431314, 
    0.001381897, 0.001327644, 0.001175244, 0.001110879, 0.001021823, 
    0.0007425516, 0.0007307242, 0.0008326205, 0.0009313844, 0.001029254,
  0.001969611, 0.001953857, 0.001751087, 0.001625228, 0.001518527, 
    0.001469287, 0.001410406, 0.001342807, 0.001226469, 0.001122528, 
    0.0008596066, 0.0007590873, 0.0008196975, 0.000912409, 0.0009862127,
  0.002047504, 0.00199633, 0.001895577, 0.001766649, 0.001590899, 
    0.001525608, 0.001485578, 0.001443221, 0.001365813, 0.001296134, 
    0.0009303325, 0.0007913189, 0.0008148858, 0.0009087075, 0.0009863926,
  0.0005373147, 0.0007805214, 0.0005494839, 0.000688454, 0.0006035151, 
    0.0005343809, 0.000637004, 0.0006768154, 0.000782443, 0.0006551942, 
    0.0006120364, 0.0007427997, 0.0004999139, 0.0004425556, 0.0002340348,
  0.001027295, 0.001005504, 0.0009166581, 0.0008526498, 0.0005107899, 
    0.0004301495, 0.0006526909, 0.0006751962, 0.0007709893, 0.0009061305, 
    0.0007893663, 0.0009951666, 0.000932599, 0.0004062481, 0.0003589842,
  0.001194022, 0.001099992, 0.001016954, 0.0009169065, 0.000756191, 
    0.0003515301, 0.0005720931, 0.0006900679, 0.0007957664, 0.0009209301, 
    0.0010626, 0.001146029, 0.001105798, 0.001030551, 0.0008822888,
  0.001263715, 0.001164421, 0.001088056, 0.001011363, 0.0009564605, 
    0.0008251561, 0.0003314013, 0.0005498652, 0.0007373804, 0.0008821575, 
    0.001074097, 0.001199308, 0.001253918, 0.001227383, 0.001170399,
  0.001384472, 0.00128414, 0.001205278, 0.0011191, 0.00106159, 0.0009778483, 
    0.00100376, 0.0003562877, 0.0004935193, 0.0007496522, 0.00105561, 
    0.001203255, 0.001278205, 0.001284672, 0.001289382,
  0.001573931, 0.00149022, 0.001390371, 0.001291875, 0.001173697, 
    0.001082886, 0.001017811, 0.001078487, 0.0008554214, 0.0008177335, 
    0.0009578709, 0.00114646, 0.001208172, 0.001255337, 0.001285275,
  0.001847709, 0.001745894, 0.001634079, 0.001521914, 0.001432419, 
    0.001259308, 0.001100925, 0.001113743, 0.0009630601, 0.0008648491, 
    0.0009729539, 0.001030203, 0.001079856, 0.001157657, 0.001176759,
  0.002167573, 0.002016585, 0.001866266, 0.001725203, 0.001628359, 
    0.001502276, 0.001414135, 0.001286658, 0.001152089, 0.0009404718, 
    0.0009455087, 0.0009860464, 0.001018292, 0.00106275, 0.001061653,
  0.002766941, 0.002561068, 0.002344088, 0.002050011, 0.001799255, 
    0.001653079, 0.001551699, 0.001477036, 0.001362495, 0.001017129, 
    0.0009170455, 0.000954263, 0.001006527, 0.001003009, 0.001081152,
  0.003370462, 0.003073762, 0.002814954, 0.002461525, 0.002052115, 
    0.001787674, 0.00163222, 0.001580021, 0.001502705, 0.001090751, 
    0.0009016439, 0.0009133887, 0.0009744045, 0.0009527082, 0.000928279,
  0.0005341409, 0.0008826249, 0.0009600315, 0.001047156, 0.0007562609, 
    0.000584148, 0.0008892031, 0.001049999, 0.001167649, 0.0008060374, 
    0.0007696306, 0.0009845537, 0.0008126931, 0.0007442924, 0.0005443592,
  0.001040602, 0.001075951, 0.0009898562, 0.0009579254, 0.0006458763, 
    0.0004938116, 0.0008551904, 0.001015583, 0.001103399, 0.001110524, 
    0.0009045989, 0.00116826, 0.001149286, 0.0006721864, 0.0006703583,
  0.00121307, 0.001147719, 0.001091314, 0.001044464, 0.00117624, 
    0.0004658278, 0.0006519388, 0.001005674, 0.001107991, 0.001102994, 
    0.001084485, 0.001137539, 0.001129116, 0.001069996, 0.001038198,
  0.001355185, 0.001272149, 0.001253757, 0.001222565, 0.001185567, 
    0.001282745, 0.000334508, 0.0006546882, 0.0009608683, 0.001023664, 
    0.001028946, 0.001054963, 0.001086033, 0.001063013, 0.001050826,
  0.001524473, 0.001497808, 0.001458212, 0.001387928, 0.001265825, 
    0.001212428, 0.001366718, 0.000367339, 0.0006267116, 0.0007608711, 
    0.0009521634, 0.0009843967, 0.001014404, 0.001011328, 0.0009952179,
  0.001735846, 0.001725, 0.001662737, 0.001593734, 0.001512472, 0.001266592, 
    0.001425831, 0.001206863, 0.0008933156, 0.0008955363, 0.0009561845, 
    0.0009532101, 0.0009628076, 0.0009675283, 0.0009682935,
  0.002045075, 0.001932436, 0.001862278, 0.001777547, 0.001738863, 
    0.001592762, 0.001503929, 0.00119044, 0.0009233949, 0.0008149219, 
    0.001059868, 0.000981533, 0.0009577794, 0.0009486928, 0.0009455047,
  0.002888527, 0.002589704, 0.002339725, 0.002073884, 0.001902553, 
    0.00176095, 0.001644253, 0.00154557, 0.001174547, 0.0008917419, 
    0.0009982439, 0.0009940504, 0.0009661579, 0.0009524039, 0.0009235491,
  0.002989678, 0.002987709, 0.002969476, 0.002798998, 0.002446956, 
    0.002086795, 0.001808255, 0.001745381, 0.00160857, 0.001083056, 
    0.001033956, 0.0009709422, 0.0009494151, 0.0009543331, 0.0009152948,
  0.002413466, 0.002476096, 0.002556591, 0.002960916, 0.00289151, 0.00256091, 
    0.00209713, 0.001861234, 0.001759731, 0.001230514, 0.001099309, 
    0.0009974861, 0.0009327075, 0.0009302826, 0.0008835403,
  0.000552893, 0.0008929609, 0.0009882366, 0.001260897, 0.001088799, 
    0.0006892661, 0.0008799786, 0.0009201678, 0.000943662, 0.0006675241, 
    0.000623949, 0.0008122245, 0.0007855237, 0.000775423, 0.0005889317,
  0.001104261, 0.001247855, 0.001326396, 0.00132429, 0.0009368055, 
    0.0005478994, 0.0007878274, 0.0008937292, 0.0008923783, 0.0008558935, 
    0.0007508846, 0.0008794786, 0.0009293854, 0.000703922, 0.0006539749,
  0.00128977, 0.001258296, 0.001239815, 0.001366237, 0.00152618, 
    0.0005731707, 0.0006570735, 0.0008422083, 0.0008530967, 0.0008403381, 
    0.000812908, 0.0008768275, 0.0009082113, 0.001000202, 0.0009943329,
  0.001365829, 0.001331817, 0.001278924, 0.001369915, 0.00145947, 
    0.001603981, 0.0005563722, 0.00061446, 0.0007305252, 0.0008060838, 
    0.0007800685, 0.0008539949, 0.0008914869, 0.0009640569, 0.001054368,
  0.00150186, 0.001454037, 0.001417143, 0.001442067, 0.001486795, 
    0.001723685, 0.00165601, 0.000374269, 0.0004001498, 0.0007283142, 
    0.0008174353, 0.0008468534, 0.0008667379, 0.0009219896, 0.001056243,
  0.001631551, 0.001597764, 0.0015486, 0.001528376, 0.001584384, 0.001627145, 
    0.001767067, 0.001675269, 0.00107615, 0.0009142941, 0.0008415225, 
    0.0009039906, 0.0008648193, 0.000872373, 0.0009711111,
  0.001846651, 0.001746741, 0.001689313, 0.001628597, 0.001652272, 
    0.001671363, 0.001750827, 0.001635544, 0.001357218, 0.001064977, 
    0.001070352, 0.001038734, 0.0009333307, 0.0008568658, 0.0009155434,
  0.002201915, 0.001986342, 0.001871417, 0.001804298, 0.001773144, 
    0.001768922, 0.001833677, 0.001769201, 0.001685568, 0.001431528, 
    0.001293811, 0.001198343, 0.001039515, 0.0009004368, 0.0008854038,
  0.002394401, 0.00226598, 0.002208276, 0.002136066, 0.0020488, 0.001976997, 
    0.001990201, 0.001976351, 0.001903861, 0.001815302, 0.001586839, 
    0.001381361, 0.001176397, 0.0009948596, 0.0009237388,
  0.002370987, 0.002291222, 0.002254694, 0.00230897, 0.002306225, 
    0.002317201, 0.002299361, 0.002301476, 0.002202974, 0.002048776, 
    0.001860846, 0.001585289, 0.001319788, 0.001102283, 0.0009940605,
  0.0006755121, 0.0008474457, 0.0007146689, 0.0007368508, 0.0007282908, 
    0.0006791523, 0.0007444739, 0.000720392, 0.0007642721, 0.0005719279, 
    0.000597754, 0.0007150251, 0.0007185221, 0.0007549985, 0.0005324639,
  0.001217584, 0.00133114, 0.001353839, 0.00122484, 0.0007395571, 
    0.0005881015, 0.0007312061, 0.0007829908, 0.0007713556, 0.0007045662, 
    0.000622788, 0.0008922705, 0.001015559, 0.0006633607, 0.0006205223,
  0.001406589, 0.001410181, 0.001433711, 0.001394995, 0.001291472, 
    0.0004760293, 0.0009073554, 0.0007851818, 0.0007767596, 0.0007278598, 
    0.0007847825, 0.001002138, 0.001101404, 0.001108407, 0.001020487,
  0.001421558, 0.001400608, 0.001430688, 0.001473772, 0.001503381, 
    0.001603098, 0.0008177204, 0.000769066, 0.0008854743, 0.0007979902, 
    0.0008216473, 0.001067279, 0.001138487, 0.001173758, 0.001087694,
  0.001408303, 0.00139127, 0.001350541, 0.001391966, 0.001502815, 0.00165702, 
    0.001787057, 0.001076275, 0.0008854249, 0.0009459851, 0.0009442134, 
    0.00119766, 0.001256358, 0.001258711, 0.001157919,
  0.001430536, 0.001409882, 0.001378882, 0.001382363, 0.001447495, 
    0.001482901, 0.001665601, 0.001998274, 0.001661808, 0.001411274, 
    0.001191822, 0.001383294, 0.00148565, 0.001424069, 0.001313887,
  0.001480456, 0.001453133, 0.001419892, 0.0014122, 0.001440885, 0.001491514, 
    0.001549642, 0.001680142, 0.002047418, 0.002005052, 0.001753208, 
    0.001749158, 0.001767343, 0.001652846, 0.001449171,
  0.001571106, 0.001532083, 0.001499469, 0.001484787, 0.00151539, 
    0.001577635, 0.00166841, 0.001745716, 0.001855526, 0.002109743, 
    0.002073617, 0.00202966, 0.001987494, 0.001834719, 0.001657312,
  0.001699813, 0.00167232, 0.001652212, 0.001652831, 0.00169244, 0.001748815, 
    0.00181815, 0.001890395, 0.001991543, 0.002105271, 0.002076475, 
    0.00207196, 0.002090856, 0.001962824, 0.001834271,
  0.001893193, 0.001808029, 0.001801415, 0.001833273, 0.001892647, 
    0.001963301, 0.002027125, 0.002119849, 0.002241175, 0.002143055, 
    0.002193006, 0.002110961, 0.002078997, 0.002020758, 0.001927831,
  0.0007152242, 0.0008318364, 0.0007638162, 0.000768077, 0.0006625067, 
    0.0005937974, 0.0006507834, 0.0006394563, 0.0006145029, 0.0005030361, 
    0.0005064808, 0.0006863811, 0.0007530211, 0.000934726, 0.0005782566,
  0.001162282, 0.001304111, 0.001308041, 0.001043943, 0.0006541855, 
    0.0005863697, 0.0006901795, 0.0006818559, 0.0006953478, 0.0007521355, 
    0.0006846727, 0.0009078538, 0.00123332, 0.001182003, 0.0006318286,
  0.001452836, 0.001534318, 0.001554312, 0.001393188, 0.0009059472, 
    0.0004818485, 0.0007574465, 0.0007563143, 0.0008719402, 0.0009974671, 
    0.00106104, 0.001312933, 0.001499479, 0.001589967, 0.000926148,
  0.001567465, 0.001638812, 0.00163147, 0.001535972, 0.001372576, 
    0.001092238, 0.0005287361, 0.000713298, 0.001277442, 0.001381364, 
    0.001348761, 0.001560515, 0.001753439, 0.001708115, 0.001072198,
  0.001603156, 0.001650623, 0.001642448, 0.00156528, 0.00146826, 0.001394933, 
    0.001367623, 0.000795011, 0.001049342, 0.001560173, 0.001673619, 
    0.001752669, 0.001880362, 0.001918858, 0.001279709,
  0.001640499, 0.001643406, 0.001599604, 0.00153851, 0.001483597, 
    0.001462336, 0.001448104, 0.001540226, 0.001508851, 0.001811892, 
    0.001760342, 0.001868297, 0.001952122, 0.002015541, 0.001586202,
  0.0016725, 0.001653704, 0.001604979, 0.001545453, 0.001521908, 0.001507511, 
    0.001514627, 0.001533778, 0.001724925, 0.002049942, 0.002002914, 
    0.001970698, 0.001978321, 0.002027512, 0.00176195,
  0.001669067, 0.001641816, 0.001597452, 0.001556685, 0.0015306, 0.001538252, 
    0.001547033, 0.001594135, 0.001704924, 0.001891246, 0.001866029, 
    0.001897239, 0.001969662, 0.002071979, 0.001978893,
  0.0016385, 0.001613835, 0.001578916, 0.00154789, 0.001527505, 0.001538938, 
    0.001579936, 0.001669915, 0.001755652, 0.001968544, 0.001931839, 
    0.001993196, 0.002019028, 0.002111709, 0.002200688,
  0.001577043, 0.001546877, 0.001538685, 0.001554168, 0.001572407, 
    0.001609553, 0.001671082, 0.001746873, 0.001944382, 0.0019266, 
    0.002081373, 0.002223962, 0.002272513, 0.002332616, 0.00238812,
  0.0006399217, 0.0007436967, 0.0006720006, 0.0007074457, 0.0006096797, 
    0.0005158479, 0.0005751852, 0.0006405133, 0.0008366935, 0.0009964192, 
    0.0009304913, 0.000911308, 0.000577361, 0.0003797749, 0.0002072982,
  0.001212562, 0.001250322, 0.001212675, 0.0008779019, 0.0005933613, 
    0.0004913741, 0.0006522388, 0.0006690617, 0.0009278533, 0.001243974, 
    0.00131382, 0.001371565, 0.001120669, 0.0005583861, 0.0003896057,
  0.001550528, 0.001509903, 0.001452224, 0.001303954, 0.0008521124, 
    0.0003978443, 0.000665337, 0.0007179885, 0.00103521, 0.001465134, 
    0.001696442, 0.001825414, 0.001609524, 0.0012815, 0.0008210012,
  0.001694216, 0.001629946, 0.001562512, 0.001503406, 0.001360213, 
    0.001063915, 0.0004733276, 0.0006757177, 0.001136875, 0.001697748, 
    0.001699669, 0.001802116, 0.001926178, 0.001642767, 0.001176294,
  0.001728136, 0.001661641, 0.001615873, 0.001592689, 0.001493573, 
    0.001398712, 0.001245145, 0.000520603, 0.0007356763, 0.001518421, 
    0.001733886, 0.001761356, 0.001873448, 0.001794476, 0.001499333,
  0.001747927, 0.001700606, 0.001665378, 0.001631599, 0.001583634, 
    0.001487135, 0.001402169, 0.001510815, 0.001242288, 0.001534973, 
    0.001713628, 0.001786427, 0.001799054, 0.001708836, 0.001791314,
  0.001785782, 0.001766114, 0.001728073, 0.001671967, 0.001590073, 
    0.001495953, 0.001460526, 0.001398789, 0.001346234, 0.001541825, 
    0.001839971, 0.001883263, 0.001745622, 0.001796509, 0.00195506,
  0.001793228, 0.001810102, 0.001814131, 0.001764478, 0.001661437, 
    0.001551032, 0.001510049, 0.001462653, 0.001389684, 0.001605127, 
    0.001763706, 0.001813625, 0.001869358, 0.001976732, 0.002115096,
  0.00179936, 0.001839361, 0.001862653, 0.00181951, 0.001746863, 0.001644525, 
    0.001546473, 0.001501706, 0.001479853, 0.001645314, 0.001588511, 
    0.001616553, 0.00195056, 0.002013252, 0.00216947,
  0.001804967, 0.001830861, 0.001829621, 0.001810204, 0.001771326, 
    0.001708287, 0.001631921, 0.001554876, 0.001569871, 0.001531968, 
    0.001772571, 0.001790676, 0.001791875, 0.002029203, 0.002202246,
  0.0005546997, 0.0006438819, 0.0005687734, 0.0006905457, 0.0006276005, 
    0.0005129021, 0.0007762783, 0.001018135, 0.001252765, 0.001243826, 
    0.00125186, 0.001450251, 0.00140048, 0.001222659, 0.0006667318,
  0.001077508, 0.001087011, 0.00108648, 0.0008024375, 0.0004941471, 
    0.0003988909, 0.0006993039, 0.000849886, 0.001128399, 0.001354674, 
    0.001327486, 0.001553943, 0.001682579, 0.00134884, 0.0008224295,
  0.001359686, 0.001340087, 0.001318234, 0.001223641, 0.000842914, 
    0.0002809544, 0.000627997, 0.0007396014, 0.00101136, 0.001333233, 
    0.001394806, 0.001542983, 0.001696993, 0.00154061, 0.001029769,
  0.001518312, 0.00146591, 0.001446389, 0.001408556, 0.001365549, 
    0.001190589, 0.0004497012, 0.0006766762, 0.0008755163, 0.001263477, 
    0.001350476, 0.001479164, 0.001658964, 0.001567368, 0.001132106,
  0.001596008, 0.0015498, 0.001499734, 0.001476685, 0.00145451, 0.001421796, 
    0.001418607, 0.0005866642, 0.0005048659, 0.0009783038, 0.00132427, 
    0.001408002, 0.00162087, 0.001605785, 0.001304505,
  0.001662869, 0.001644569, 0.001593091, 0.001559491, 0.001551103, 
    0.001517796, 0.001491101, 0.001577457, 0.00134732, 0.0012027, 
    0.001195421, 0.001430198, 0.001561503, 0.001617254, 0.00137821,
  0.001760017, 0.001744019, 0.001660342, 0.001606949, 0.001589101, 
    0.001580857, 0.001556474, 0.001564142, 0.001609548, 0.001534907, 
    0.001401651, 0.001428962, 0.00154877, 0.001656213, 0.001514172,
  0.001833746, 0.001758732, 0.001715945, 0.001690237, 0.001673387, 
    0.001666671, 0.00166148, 0.001636303, 0.001630707, 0.001677382, 
    0.001461319, 0.001418725, 0.00147637, 0.001606505, 0.00162753,
  0.001893629, 0.001875348, 0.001867759, 0.001857447, 0.001862801, 
    0.001864135, 0.001841903, 0.001818325, 0.001756637, 0.001740225, 
    0.001538153, 0.001433396, 0.0013849, 0.001397194, 0.001767821,
  0.00189059, 0.001956306, 0.002013876, 0.00205155, 0.002083672, 0.002117622, 
    0.002107689, 0.002072674, 0.002003253, 0.001772325, 0.001753278, 
    0.001581199, 0.001366842, 0.00132212, 0.001744313,
  0.0007241182, 0.0009032185, 0.000885118, 0.0009491201, 0.0007176324, 
    0.0005786545, 0.0007864104, 0.0008492902, 0.0008903458, 0.0005727883, 
    0.0005645187, 0.0005719436, 0.000259701, 0.0001440574, 8.19065e-05,
  0.001215434, 0.00118177, 0.00119123, 0.001013099, 0.0005383793, 
    0.0004769819, 0.0008191947, 0.0009546555, 0.0009949026, 0.0007990211, 
    0.000608502, 0.0006609882, 0.0003760233, 0.0001216634, 8.008149e-05,
  0.001327455, 0.001251052, 0.001190657, 0.001122814, 0.00096764, 
    0.0004069997, 0.0008184594, 0.00104674, 0.001142321, 0.0009812211, 
    0.0008674367, 0.0006841945, 0.0004265632, 0.0002747808, 0.0001684489,
  0.001405973, 0.0013454, 0.001305404, 0.001295012, 0.001313527, 0.001295781, 
    0.0008498309, 0.001120001, 0.001260284, 0.001075744, 0.0009242778, 
    0.0007748912, 0.0004679832, 0.0002964043, 0.0002333029,
  0.001480902, 0.001384801, 0.001327737, 0.001354692, 0.001428958, 
    0.001539308, 0.001575427, 0.001046569, 0.001124756, 0.001074435, 
    0.0009886094, 0.000830099, 0.0005806389, 0.0003588048, 0.0003164147,
  0.001500556, 0.001502338, 0.001495241, 0.001531269, 0.001619591, 
    0.00167521, 0.001721934, 0.001916439, 0.001747145, 0.001488174, 
    0.001012802, 0.0009333655, 0.0007152631, 0.0004361532, 0.0003739221,
  0.001585115, 0.001632098, 0.001662944, 0.001707396, 0.00176867, 
    0.001826991, 0.001861096, 0.001877925, 0.002009093, 0.001870518, 
    0.001353983, 0.001082057, 0.0009234918, 0.0005546029, 0.0004393814,
  0.001683079, 0.001685944, 0.001723017, 0.001775006, 0.001843165, 
    0.001893738, 0.001919581, 0.001894396, 0.001995322, 0.001996093, 
    0.001509255, 0.001237752, 0.001160859, 0.0007596762, 0.0005350077,
  0.00176689, 0.001757296, 0.001798232, 0.001848219, 0.00195022, 0.001973364, 
    0.002002429, 0.002096235, 0.002027673, 0.002069849, 0.00162487, 
    0.00138307, 0.001191263, 0.001068881, 0.0006670808,
  0.001888414, 0.001894016, 0.001959585, 0.00205647, 0.002093467, 
    0.002137283, 0.002273837, 0.002335529, 0.002370083, 0.001991491, 
    0.001911539, 0.001530083, 0.001273909, 0.001111755, 0.001158145,
  0.001011945, 0.001070649, 0.000900061, 0.001097145, 0.000978273, 
    0.0008341064, 0.001062182, 0.000929612, 0.0005320949, 0.000215528, 
    0.0001686452, 0.000196181, 0.0001625248, 0.0001944151, 0.0001696597,
  0.001118703, 0.001040105, 0.001119513, 0.001246139, 0.0009754961, 
    0.0008650382, 0.001250837, 0.00128711, 0.0007884277, 0.0004153641, 
    0.000258016, 0.0003062661, 0.000330714, 0.000183368, 0.0001826304,
  0.001184081, 0.001079991, 0.001055778, 0.001246713, 0.001468002, 
    0.0008529571, 0.001348443, 0.001518704, 0.001161882, 0.0006689625, 
    0.0004543115, 0.0003825845, 0.0003567094, 0.0003711366, 0.0003498574,
  0.001275005, 0.00117553, 0.001188951, 0.00138506, 0.001647404, 0.001863416, 
    0.001400426, 0.001549657, 0.00131492, 0.0008610422, 0.0005577827, 
    0.0004335799, 0.0003901842, 0.0003883474, 0.0004105546,
  0.001370085, 0.001309964, 0.001336675, 0.001532742, 0.001762114, 
    0.001972416, 0.002198869, 0.001540276, 0.001289247, 0.0009402534, 
    0.0006789364, 0.000523798, 0.0004232656, 0.0004274448, 0.0004520239,
  0.001483923, 0.001474753, 0.001495246, 0.00168535, 0.001845235, 0.00201331, 
    0.002106791, 0.002286825, 0.001686163, 0.001228366, 0.0007581012, 
    0.000608984, 0.0004962829, 0.000455825, 0.0004795869,
  0.001578284, 0.001586504, 0.001654015, 0.001738999, 0.001859031, 
    0.002035678, 0.002112809, 0.002069438, 0.002082617, 0.001568908, 
    0.001070801, 0.000765688, 0.0005828826, 0.0005112399, 0.0005214442,
  0.001681235, 0.001666268, 0.001696638, 0.001743512, 0.001891154, 
    0.002048455, 0.002090076, 0.002044824, 0.002148803, 0.001801384, 
    0.001206083, 0.0009024697, 0.0007288269, 0.00056999, 0.0005611127,
  0.001733423, 0.0017363, 0.001750985, 0.001798249, 0.001965513, 0.002032434, 
    0.002068631, 0.002153226, 0.001981073, 0.001985841, 0.00161863, 
    0.001285802, 0.0009926077, 0.0007077972, 0.0005921789,
  0.001783836, 0.001763607, 0.001779322, 0.001851615, 0.001964916, 
    0.001974782, 0.002094628, 0.002018015, 0.002007436, 0.001783119, 
    0.001840524, 0.001569021, 0.001245699, 0.0009175009, 0.0006752075,
  0.0006891138, 0.0009053152, 0.0009228467, 0.001148973, 0.001127763, 
    0.00115084, 0.001438358, 0.001423014, 0.001045001, 0.000871529, 
    0.0006844496, 0.0005937198, 0.000340051, 0.0003368688, 0.0002758084,
  0.001167, 0.001198509, 0.001297872, 0.001403518, 0.001098799, 0.001144961, 
    0.001524102, 0.001474195, 0.001231443, 0.001210722, 0.0008774535, 
    0.0008145621, 0.0005669123, 0.0003110611, 0.0002946844,
  0.001283128, 0.001259918, 0.001289319, 0.001348023, 0.001557069, 
    0.001194655, 0.001548743, 0.001518868, 0.001367108, 0.001217326, 
    0.001175581, 0.0009446606, 0.0006095088, 0.0005738156, 0.0005165777,
  0.001388078, 0.00136364, 0.001368269, 0.001438028, 0.001642602, 
    0.001916641, 0.001252117, 0.001415641, 0.001403864, 0.001323674, 
    0.001225082, 0.0009907987, 0.0006596657, 0.0006051211, 0.0005786285,
  0.001414535, 0.001426133, 0.001449454, 0.00153648, 0.001729385, 
    0.001853705, 0.002119693, 0.001551975, 0.001540363, 0.001302743, 
    0.001248281, 0.001010937, 0.0007269967, 0.0006369418, 0.0006451333,
  0.001419205, 0.001445715, 0.001496307, 0.001606587, 0.001751732, 
    0.001848792, 0.001946479, 0.002195363, 0.00185003, 0.001790744, 
    0.001399592, 0.001158239, 0.0008108285, 0.0006622463, 0.0006483495,
  0.001525165, 0.001537761, 0.001581834, 0.001662928, 0.001754125, 
    0.001827131, 0.001914349, 0.001979847, 0.002194604, 0.002003897, 
    0.001750783, 0.001296222, 0.0009588992, 0.0006782047, 0.0006592525,
  0.001622043, 0.001633731, 0.001644926, 0.001688099, 0.001750435, 
    0.001812569, 0.001881293, 0.001946454, 0.00214736, 0.001987186, 
    0.001720892, 0.001404346, 0.001098212, 0.0007497136, 0.0006495544,
  0.001706886, 0.001728236, 0.001745677, 0.001739178, 0.001771189, 
    0.001821802, 0.001869722, 0.002097195, 0.002059748, 0.001912389, 
    0.001650961, 0.001471064, 0.001241744, 0.0008969016, 0.0006326871,
  0.00179405, 0.00177456, 0.001767276, 0.001778896, 0.001802006, 0.00187317, 
    0.00211003, 0.002152956, 0.00215794, 0.001713887, 0.001594709, 
    0.001505308, 0.001361685, 0.001179339, 0.0006925558,
  0.000728547, 0.0008389141, 0.000802741, 0.0008535275, 0.0008588271, 
    0.0008752742, 0.0009984776, 0.001106636, 0.001154936, 0.001116903, 
    0.001047013, 0.001017584, 0.0008721931, 0.0006121976, 0.0002900136,
  0.001116366, 0.001150287, 0.001200538, 0.001118788, 0.0008724961, 
    0.0009117621, 0.001162086, 0.001244093, 0.001301431, 0.0012832, 
    0.001176197, 0.001230998, 0.001137654, 0.0005714473, 0.0002376136,
  0.001312441, 0.00134687, 0.001403043, 0.001394891, 0.001400566, 
    0.0009298103, 0.001299199, 0.001387226, 0.0014125, 0.001384244, 
    0.001394528, 0.001376385, 0.001226173, 0.0008873023, 0.0003446112,
  0.001321249, 0.001401057, 0.00146473, 0.001512083, 0.001539555, 
    0.001605565, 0.001002569, 0.001313777, 0.001464233, 0.001473395, 
    0.001469263, 0.001463591, 0.001330688, 0.0009449971, 0.0004005529,
  0.001389205, 0.001480517, 0.001522401, 0.00157069, 0.001640705, 
    0.001695211, 0.001807211, 0.001321521, 0.001406153, 0.001379345, 
    0.001523979, 0.001498216, 0.00132436, 0.0009915003, 0.0005099634,
  0.001503768, 0.001564141, 0.001622208, 0.001698762, 0.001771902, 
    0.001831229, 0.001875574, 0.001966004, 0.001779384, 0.001613056, 
    0.001549704, 0.001594511, 0.001403314, 0.001040868, 0.0005861561,
  0.001835385, 0.001881036, 0.001928149, 0.001969447, 0.002025402, 
    0.002080848, 0.002142184, 0.002152846, 0.002167171, 0.0020616, 
    0.001903404, 0.001776811, 0.001502109, 0.001031725, 0.0005960962,
  0.002269211, 0.002287496, 0.002308153, 0.002341062, 0.002367453, 
    0.002402682, 0.00238511, 0.002312532, 0.002258292, 0.002176277, 
    0.002004016, 0.001854323, 0.001592517, 0.001026506, 0.0005701969,
  0.002573137, 0.002552042, 0.002537875, 0.002568557, 0.00260155, 
    0.002596208, 0.002452173, 0.002267361, 0.002217629, 0.002190038, 
    0.002091617, 0.00201002, 0.001658197, 0.0009972638, 0.000545404,
  0.002650793, 0.002676548, 0.002703668, 0.002744016, 0.002733956, 
    0.00263714, 0.002328216, 0.002176527, 0.002150555, 0.002064756, 
    0.002153034, 0.002130338, 0.001722128, 0.001005196, 0.0005359699,
  0.000699554, 0.0008198161, 0.0008361782, 0.0008853439, 0.0008195323, 
    0.0008181051, 0.000883347, 0.0008547409, 0.0008305495, 0.0007374068, 
    0.0007580665, 0.0007650347, 0.000775832, 0.0008242911, 0.0005635891,
  0.001103955, 0.00116016, 0.001256764, 0.001118203, 0.0007946377, 
    0.000854279, 0.001019641, 0.000992397, 0.0009725541, 0.0009312031, 
    0.001030779, 0.001165821, 0.001213479, 0.0009968622, 0.0005728762,
  0.001478889, 0.001482619, 0.001514723, 0.001481982, 0.001361945, 
    0.001039262, 0.00120927, 0.001243707, 0.001250267, 0.001301238, 
    0.001429166, 0.001602229, 0.001565523, 0.001393116, 0.0006128948,
  0.00171345, 0.001668374, 0.001635794, 0.001658227, 0.001664144, 0.00157775, 
    0.0009832403, 0.001361276, 0.001631058, 0.001746622, 0.002015434, 
    0.002009296, 0.001853636, 0.001549823, 0.000540811,
  0.001994272, 0.001881796, 0.001812508, 0.001811242, 0.001836097, 
    0.001862434, 0.001961708, 0.00164447, 0.001737116, 0.002137845, 
    0.002390249, 0.002101635, 0.001945733, 0.001563852, 0.0005319812,
  0.002434041, 0.002215894, 0.002054477, 0.002009465, 0.002029703, 
    0.002105238, 0.002232598, 0.002381328, 0.002502173, 0.002582751, 
    0.002313078, 0.001903123, 0.001899005, 0.001529317, 0.0004932131,
  0.002907392, 0.002677176, 0.002422991, 0.002299126, 0.002297581, 
    0.002359516, 0.002482549, 0.002639697, 0.002756238, 0.002486657, 
    0.001970892, 0.001824371, 0.001895514, 0.001292284, 0.0004454981,
  0.003234242, 0.003057419, 0.002830182, 0.00264621, 0.002558755, 
    0.002564156, 0.002623181, 0.002708294, 0.002448575, 0.002137295, 
    0.001718504, 0.001788519, 0.001869629, 0.001053781, 0.0003830277,
  0.003356381, 0.003252131, 0.003094602, 0.002881117, 0.00269839, 
    0.002633526, 0.002683086, 0.002623501, 0.002344706, 0.002133796, 
    0.001705492, 0.001815623, 0.001631507, 0.0007619575, 0.0002886952,
  0.003487154, 0.003374263, 0.00320562, 0.003026349, 0.002852073, 
    0.002759614, 0.002686532, 0.002489035, 0.002242773, 0.001851196, 
    0.001875475, 0.00182678, 0.001329434, 0.0005718228, 0.0003013432,
  0.0005653467, 0.0006503145, 0.0005754103, 0.0005638853, 0.0004959096, 
    0.0005122497, 0.0005771958, 0.0005580473, 0.0005469393, 0.0004914161, 
    0.0005083476, 0.0005760791, 0.0006128071, 0.0007766383, 0.000987743,
  0.001030076, 0.001044545, 0.001059994, 0.0008369387, 0.0004932333, 
    0.0005926592, 0.0007051868, 0.0006460512, 0.0006164488, 0.0005918749, 
    0.0005968311, 0.0007296065, 0.0008902244, 0.001141711, 0.001135792,
  0.001998008, 0.001745371, 0.001678479, 0.001545426, 0.0009355238, 
    0.000542226, 0.0007909504, 0.0007964802, 0.0007483989, 0.000725998, 
    0.0007637213, 0.0009157605, 0.001201304, 0.00142039, 0.0007627523,
  0.002638689, 0.002391872, 0.002125182, 0.001960309, 0.001757931, 
    0.001212068, 0.0006723693, 0.0008147266, 0.0009070331, 0.0009265517, 
    0.0009868335, 0.001205382, 0.00139437, 0.001380577, 0.0005289999,
  0.003200987, 0.003043976, 0.00279311, 0.002489886, 0.002220431, 0.00192935, 
    0.001514868, 0.0008159127, 0.000802559, 0.0009957084, 0.001191048, 
    0.001418144, 0.001523184, 0.001340613, 0.0005363777,
  0.003429885, 0.003359039, 0.003257617, 0.003058162, 0.002816097, 
    0.002500387, 0.00214814, 0.0016953, 0.001145376, 0.001081984, 
    0.001227081, 0.001507372, 0.001608677, 0.00110805, 0.0004609544,
  0.003293086, 0.003307332, 0.003352431, 0.003295023, 0.003244393, 
    0.003045368, 0.002770844, 0.002371054, 0.001928779, 0.001441952, 
    0.001407541, 0.001577815, 0.001502238, 0.0008322605, 0.0004164633,
  0.003235451, 0.00316531, 0.003233959, 0.00328374, 0.003319487, 0.003235711, 
    0.003075318, 0.002828456, 0.002510644, 0.001888882, 0.001626289, 
    0.001666274, 0.00141767, 0.0006550042, 0.0003647048,
  0.002666799, 0.002672524, 0.002842701, 0.003022116, 0.003131397, 
    0.003161776, 0.003022793, 0.002877151, 0.002733193, 0.002229221, 
    0.001816058, 0.001750398, 0.001275474, 0.0005207355, 0.0002949758,
  0.002536069, 0.002536399, 0.002712088, 0.002916442, 0.003100101, 
    0.003193051, 0.003148705, 0.003011506, 0.002843312, 0.002465795, 
    0.002073945, 0.00179914, 0.001098369, 0.0004498032, 0.0003100481,
  0.0006801357, 0.000764827, 0.0005610632, 0.0005722246, 0.0004503362, 
    0.0004434017, 0.000516502, 0.0004648652, 0.0004188386, 0.0002663599, 
    0.0002680117, 0.0003179486, 0.0002580939, 0.0002807371, 0.0002758795,
  0.001049558, 0.001086708, 0.000945367, 0.000705266, 0.0004249398, 
    0.0005290616, 0.0006166216, 0.0005080157, 0.0004598014, 0.0003707023, 
    0.0003250674, 0.000412379, 0.0004102991, 0.0003074974, 0.0002285541,
  0.001850608, 0.001618847, 0.001565045, 0.00130702, 0.0006143142, 
    0.0004399866, 0.0007271691, 0.0006192874, 0.0005144798, 0.0004357111, 
    0.0004421151, 0.0004252936, 0.0004359834, 0.0004674838, 0.0003640762,
  0.002718682, 0.002060678, 0.001886634, 0.001752448, 0.001386986, 
    0.0008578105, 0.0005414248, 0.000676735, 0.0006611613, 0.0005672392, 
    0.0005167002, 0.0004708103, 0.0004728396, 0.0005408352, 0.0004600755,
  0.00333237, 0.002616994, 0.002153359, 0.00199256, 0.001728831, 0.001521341, 
    0.001164922, 0.0005888499, 0.0005898732, 0.0006959871, 0.0007058849, 
    0.0006350819, 0.0005539877, 0.0006149995, 0.0005679997,
  0.002877526, 0.002867276, 0.002380818, 0.002195499, 0.001975042, 
    0.001809442, 0.001658665, 0.001435444, 0.0009012813, 0.0007790829, 
    0.0007850325, 0.0007761691, 0.0006728346, 0.0006900053, 0.0005980527,
  0.002721866, 0.002625021, 0.002409217, 0.00230155, 0.002126652, 
    0.001988027, 0.001866289, 0.001770607, 0.001625708, 0.001210466, 
    0.0009925193, 0.0008704768, 0.0007629557, 0.0007669591, 0.000578968,
  0.002678064, 0.00272123, 0.002629659, 0.002528702, 0.002390665, 
    0.002308975, 0.002190161, 0.002102792, 0.001967083, 0.001609177, 
    0.001257107, 0.001019281, 0.0008545594, 0.0007943923, 0.0005433467,
  0.002208588, 0.002297543, 0.002408716, 0.00240745, 0.002344756, 
    0.002351286, 0.002465079, 0.002457506, 0.002364893, 0.002077708, 
    0.001589581, 0.001188856, 0.0009318095, 0.0008058015, 0.0004308886,
  0.001902439, 0.001891904, 0.001857515, 0.001862941, 0.001937144, 
    0.001984441, 0.002150239, 0.002356383, 0.002594274, 0.002475013, 
    0.001991077, 0.00141547, 0.001035514, 0.0007986691, 0.0004506409,
  0.0007295397, 0.0008324006, 0.0007061284, 0.0007345272, 0.0006288448, 
    0.0006408401, 0.0007649553, 0.0005519106, 0.0004788841, 0.0003008391, 
    0.0002717559, 0.0002970071, 0.0001777537, 0.0001662506, 9.81405e-05,
  0.0009889022, 0.001068711, 0.0009282262, 0.0007779954, 0.0005619676, 
    0.0007151836, 0.0007954491, 0.000574571, 0.000529778, 0.0004376115, 
    0.0003476395, 0.0004578891, 0.0004044951, 0.0001562303, 9.111016e-05,
  0.001559616, 0.001463871, 0.001380804, 0.001093641, 0.0007463832, 
    0.000564754, 0.0008020338, 0.0006118673, 0.0005529851, 0.0004999259, 
    0.0005360996, 0.0004666483, 0.0003984795, 0.0003146709, 0.0001519918,
  0.001850971, 0.001748496, 0.001657002, 0.001524613, 0.001275157, 
    0.0009494949, 0.0005738006, 0.0006191641, 0.0006027998, 0.0005305011, 
    0.0005232096, 0.000480603, 0.0004106072, 0.0003658515, 0.0002325363,
  0.002078286, 0.001903944, 0.001784254, 0.001702762, 0.001551712, 
    0.001443962, 0.001193492, 0.0005305298, 0.0004884254, 0.0005503827, 
    0.0005935581, 0.0005669403, 0.0004569535, 0.0004641544, 0.0003687094,
  0.002264915, 0.002052471, 0.001909533, 0.00182865, 0.001700823, 
    0.001627614, 0.00158425, 0.001329946, 0.0008181965, 0.0006770099, 
    0.0006700777, 0.0006690326, 0.0005338861, 0.0005071366, 0.0004356909,
  0.002311235, 0.002207427, 0.002020054, 0.001895097, 0.001786723, 
    0.001713606, 0.001657722, 0.001586745, 0.001425917, 0.0009973689, 
    0.0008172445, 0.0007382343, 0.0006130614, 0.0005416268, 0.000475291,
  0.002318952, 0.002239102, 0.002081084, 0.001986654, 0.001852466, 
    0.001778331, 0.001692434, 0.001647165, 0.001563011, 0.001206807, 
    0.0008886121, 0.0007708575, 0.0006733821, 0.0005550971, 0.0004640881,
  0.002308368, 0.002263878, 0.002165323, 0.00205551, 0.001927608, 
    0.001836539, 0.001736998, 0.00167619, 0.001546799, 0.001331366, 
    0.001003389, 0.0008694191, 0.0007358936, 0.0005753356, 0.0004258345,
  0.002041172, 0.00209274, 0.002067862, 0.002034053, 0.001957567, 
    0.001890552, 0.001809561, 0.001762569, 0.001619371, 0.001375315, 
    0.001225714, 0.0009864488, 0.0008175382, 0.0006413048, 0.0004758633,
  0.0006924176, 0.000785089, 0.0007415057, 0.0007232876, 0.0005653313, 
    0.000544225, 0.0005748299, 0.0003997071, 0.0003769669, 0.0002224255, 
    0.0001756261, 0.0002068886, 0.0001607106, 0.0001554543, 0.0001161939,
  0.0009938903, 0.001042548, 0.001007521, 0.0007563527, 0.0005404075, 
    0.0005860864, 0.0005418597, 0.0004260966, 0.0004065919, 0.0003578054, 
    0.0002842385, 0.0003627777, 0.000338151, 0.0001402639, 0.0001053811,
  0.001461687, 0.001361495, 0.001335145, 0.0009544346, 0.0007474078, 
    0.0004153663, 0.0005218023, 0.0004619775, 0.0004611704, 0.0004571723, 
    0.0004602894, 0.0003616413, 0.0003451021, 0.0003112165, 0.0001754105,
  0.001705227, 0.001631223, 0.001575283, 0.00144781, 0.001225383, 
    0.0008673404, 0.0003997506, 0.0004810041, 0.0004874336, 0.0004389953, 
    0.0004248263, 0.0003546767, 0.0003300109, 0.0003195394, 0.000300882,
  0.001829736, 0.00174327, 0.001665047, 0.001607806, 0.00150465, 0.00133652, 
    0.001044295, 0.0004342902, 0.0003684447, 0.0003980269, 0.0004751119, 
    0.000428449, 0.0003760955, 0.0003906198, 0.0003893851,
  0.001921491, 0.001818144, 0.001728896, 0.001645071, 0.001591721, 
    0.001505118, 0.001427005, 0.001197398, 0.0008058314, 0.0006718881, 
    0.0006067447, 0.0005806125, 0.0004580909, 0.000429121, 0.0003854443,
  0.002043021, 0.001928245, 0.001794532, 0.001698048, 0.001603407, 
    0.001559556, 0.001450502, 0.001351744, 0.001238666, 0.00098761, 
    0.0008171339, 0.0006992315, 0.0005495303, 0.0004834245, 0.0004098232,
  0.002148894, 0.002017749, 0.001860049, 0.001753366, 0.001650754, 
    0.001586144, 0.001504414, 0.001453628, 0.001350679, 0.001071228, 
    0.0008455387, 0.0006986639, 0.0005965147, 0.0004848515, 0.000404595,
  0.002197345, 0.00209347, 0.001970924, 0.001814062, 0.001699995, 
    0.001603049, 0.001558949, 0.001488519, 0.001359148, 0.0011325, 
    0.0008524375, 0.0007399777, 0.0006477156, 0.0005126146, 0.0004200353,
  0.002225563, 0.002109728, 0.001968168, 0.001863603, 0.001750124, 
    0.001653766, 0.001564936, 0.001485748, 0.00142708, 0.001069214, 
    0.001067875, 0.0008652624, 0.0007183675, 0.0006029613, 0.0004960757,
  0.0005856088, 0.0006542181, 0.0006054405, 0.0005714492, 0.0004502237, 
    0.0004115941, 0.000448596, 0.0004011734, 0.0004419372, 0.0003177136, 
    0.0002583889, 0.0003183697, 0.0002269185, 0.0001838898, 0.0001324752,
  0.0009595355, 0.0009130124, 0.0008729884, 0.0005684305, 0.0004269073, 
    0.000376967, 0.0004147608, 0.0004094234, 0.0004410677, 0.0004655865, 
    0.0003472005, 0.0004403875, 0.0004347783, 0.0002007242, 0.0001454669,
  0.001318085, 0.001170483, 0.001103017, 0.0006910622, 0.0005854084, 
    0.0002807908, 0.0004097836, 0.0004373883, 0.0004547601, 0.0004669891, 
    0.0004639566, 0.0004352486, 0.0004535422, 0.0004228121, 0.0002457704,
  0.00151722, 0.001440006, 0.001360184, 0.00113792, 0.001020543, 
    0.0006556257, 0.0003290131, 0.0004038284, 0.000432577, 0.0004195703, 
    0.000416479, 0.000413151, 0.0004371831, 0.000462166, 0.0004259939,
  0.001592805, 0.0014896, 0.001413063, 0.001321107, 0.00120365, 0.001066488, 
    0.0009455788, 0.0003461261, 0.0002796785, 0.0003870326, 0.000476735, 
    0.0004918539, 0.0004637253, 0.0004987291, 0.0005519452,
  0.001597805, 0.001503231, 0.001439677, 0.001360388, 0.001291887, 
    0.001209173, 0.001138792, 0.0009952913, 0.0007396303, 0.0006839994, 
    0.0005417907, 0.0005729682, 0.0005075648, 0.0004952345, 0.0005332779,
  0.001600043, 0.001516102, 0.001451074, 0.001377596, 0.001347307, 
    0.001291168, 0.001223658, 0.001111259, 0.001048288, 0.0008592383, 
    0.0007015942, 0.0006278704, 0.000564535, 0.0005177733, 0.0005041157,
  0.001620217, 0.001538604, 0.00146637, 0.001409505, 0.001375973, 
    0.001349368, 0.001287955, 0.001247152, 0.001074428, 0.0008601648, 
    0.0007181838, 0.000652898, 0.0006163655, 0.0005208545, 0.0005463911,
  0.001653038, 0.001571015, 0.001527611, 0.001445692, 0.001391886, 
    0.001369118, 0.001304432, 0.001250981, 0.001105719, 0.0008392819, 
    0.0007528021, 0.0007381953, 0.000696536, 0.0005850735, 0.0005862475,
  0.001663509, 0.001562643, 0.001510915, 0.001450657, 0.001397134, 
    0.00134126, 0.001270592, 0.001206954, 0.001079183, 0.000700467, 
    0.0008202506, 0.0008618213, 0.0007969311, 0.0006861088, 0.0006486044,
  0.0005718856, 0.0006575185, 0.000581726, 0.0005798685, 0.0004978992, 
    0.0004434825, 0.0004855823, 0.000452778, 0.0004439391, 0.000286967, 
    0.0002118449, 0.0002300698, 0.0002009032, 0.0002044125, 0.0001564908,
  0.000962219, 0.0008876296, 0.0007969941, 0.000594289, 0.0004487896, 
    0.0003780686, 0.0004909456, 0.0004998168, 0.0005144307, 0.0005024357, 
    0.0004056095, 0.0004557274, 0.0004740272, 0.0002956806, 0.0002305706,
  0.001332828, 0.001097304, 0.001045105, 0.0007215677, 0.0006638818, 
    0.0002905615, 0.000471285, 0.0005333505, 0.0005577914, 0.0005630927, 
    0.0005647501, 0.0005649414, 0.0005839382, 0.0005873004, 0.0004456201,
  0.001554049, 0.001409102, 0.001295386, 0.001108189, 0.001060434, 
    0.0007900883, 0.0003398995, 0.0005312208, 0.0006076843, 0.0005964773, 
    0.0005905885, 0.000625112, 0.0006765665, 0.0007384684, 0.0007092804,
  0.001653976, 0.001513857, 0.00140855, 0.001341148, 0.001234739, 
    0.001146543, 0.001217879, 0.0004293392, 0.000455818, 0.0006248479, 
    0.0006669543, 0.0007317648, 0.0007570075, 0.0008416215, 0.0008694509,
  0.001713462, 0.001582627, 0.001495232, 0.001422251, 0.001368435, 
    0.001339724, 0.001257881, 0.001132843, 0.0009529184, 0.0008073782, 
    0.0006767202, 0.0007712537, 0.0008301546, 0.0008903242, 0.0009823235,
  0.0017863, 0.001686725, 0.00155625, 0.001473905, 0.001424833, 0.001406805, 
    0.001379112, 0.001320676, 0.001168384, 0.0009218896, 0.000796016, 
    0.0007762514, 0.0008206377, 0.0008830959, 0.0009879469,
  0.001832729, 0.001716812, 0.001611666, 0.001521661, 0.001443346, 
    0.001420659, 0.00138205, 0.001347773, 0.001167099, 0.0009128304, 
    0.0008228784, 0.0007666813, 0.0007644899, 0.0008074811, 0.0009338213,
  0.001819699, 0.00174293, 0.001659033, 0.001552702, 0.001464309, 
    0.001408877, 0.001362894, 0.001293366, 0.001258953, 0.001017803, 
    0.0009370961, 0.0008281206, 0.0007402391, 0.0007579487, 0.0008346671,
  0.001780895, 0.001698511, 0.001640098, 0.001540311, 0.0014702, 0.001361023, 
    0.001278393, 0.001257438, 0.001207715, 0.000980781, 0.001076019, 
    0.0008929817, 0.0007392342, 0.0006933187, 0.000774834,
  0.0006187005, 0.0006576809, 0.0005988256, 0.0005145984, 0.000441419, 
    0.0003932725, 0.0003685628, 0.0003525113, 0.0003623695, 0.0002307781, 
    0.000202856, 0.0002700946, 0.0002514528, 0.0002700058, 0.0002093802,
  0.0008827003, 0.0007882376, 0.0007035334, 0.0005636833, 0.0004722332, 
    0.0003722064, 0.000455437, 0.0004257986, 0.0004215823, 0.0003921341, 
    0.0003131181, 0.0004162567, 0.0004505159, 0.0002473947, 0.0001795486,
  0.001139758, 0.0009596285, 0.0009475602, 0.0006904483, 0.000642782, 
    0.0002975216, 0.0005415981, 0.0005700586, 0.0005587896, 0.0005276586, 
    0.0005005422, 0.0005260546, 0.0005367108, 0.0005166429, 0.0003029112,
  0.001339609, 0.001263264, 0.001228132, 0.001083822, 0.001057791, 
    0.000837152, 0.0004386109, 0.0006647559, 0.0006985556, 0.0006202398, 
    0.000564122, 0.0005747019, 0.000580575, 0.0005753569, 0.0004347412,
  0.001440472, 0.001402037, 0.001425468, 0.001488343, 0.001399742, 
    0.001306242, 0.001198223, 0.000573448, 0.0005647462, 0.0006407632, 
    0.0007083645, 0.000676349, 0.0006772261, 0.0006839155, 0.0005588837,
  0.001574434, 0.001537906, 0.001545052, 0.001602249, 0.001653891, 
    0.001552669, 0.001421333, 0.001230917, 0.001044134, 0.0009565089, 
    0.0007746632, 0.0008407736, 0.000780293, 0.0007134754, 0.0006710378,
  0.001686243, 0.001661366, 0.001655966, 0.00168232, 0.001670577, 
    0.001708584, 0.001633301, 0.001464978, 0.001214125, 0.001075625, 
    0.001020806, 0.0009364937, 0.0008480718, 0.0007394461, 0.0007220028,
  0.001800049, 0.001739491, 0.00169577, 0.001690458, 0.001682626, 
    0.001676549, 0.001598556, 0.001466744, 0.001161866, 0.001073006, 
    0.001060551, 0.001043072, 0.001016147, 0.001044748, 0.001099097,
  0.001862204, 0.001783245, 0.001724745, 0.001685196, 0.001646061, 
    0.001629141, 0.001573864, 0.001428878, 0.001214002, 0.001070262, 
    0.001049793, 0.001041796, 0.001012451, 0.0009542105, 0.0009074672,
  0.001878266, 0.001775865, 0.001701103, 0.00163127, 0.001547736, 
    0.001516532, 0.001455474, 0.001383164, 0.001124563, 0.001004735, 
    0.0009698153, 0.0008945802, 0.0008738083, 0.0008339591, 0.0008403087,
  0.0005247268, 0.0005166846, 0.0004362356, 0.0004599867, 0.0004034601, 
    0.0004306459, 0.000509102, 0.0005583526, 0.0005952805, 0.0005120296, 
    0.0004786394, 0.0004708976, 0.000365667, 0.0003343772, 0.0002320368,
  0.0007512511, 0.00067175, 0.0005970386, 0.0005017136, 0.0004091033, 
    0.0003795661, 0.0005355185, 0.0005893821, 0.0006297979, 0.0006534199, 
    0.0005711545, 0.0006045422, 0.0005594786, 0.0003176811, 0.0002414889,
  0.001058288, 0.0008611314, 0.0008543879, 0.0005987749, 0.0005371646, 
    0.0002926128, 0.0005163579, 0.0005851996, 0.0006259656, 0.0006505011, 
    0.0006494515, 0.0006293396, 0.0006058646, 0.0004891727, 0.0003546571,
  0.001322816, 0.00120849, 0.00115602, 0.000923404, 0.0008615024, 
    0.0006656286, 0.0003646857, 0.0005181297, 0.000591674, 0.0005979706, 
    0.0006160634, 0.0006066205, 0.0005863518, 0.0005067084, 0.0004394632,
  0.001463922, 0.001421149, 0.001356309, 0.001262846, 0.001175242, 
    0.00105552, 0.001032866, 0.0004134533, 0.000372236, 0.000530567, 
    0.0006512934, 0.000672565, 0.0006680376, 0.000623363, 0.0005709312,
  0.001622652, 0.001604425, 0.001556579, 0.001479653, 0.001417674, 
    0.001280261, 0.001152468, 0.001089926, 0.0008878991, 0.0007254849, 
    0.0006813114, 0.0007465268, 0.0007227878, 0.0006958267, 0.0006727126,
  0.001783108, 0.001805619, 0.001741442, 0.001637089, 0.001563679, 
    0.001494439, 0.001358996, 0.001239676, 0.001082664, 0.0008601652, 
    0.0008037882, 0.0007434867, 0.000721026, 0.0006649557, 0.0006572898,
  0.001906366, 0.001897818, 0.001862454, 0.001761604, 0.001685654, 
    0.001573412, 0.00148202, 0.00142743, 0.001065721, 0.0008834114, 
    0.0008306673, 0.000792676, 0.0008215234, 0.0007718826, 0.000690217,
  0.001970042, 0.001888875, 0.001849998, 0.001803312, 0.00174351, 
    0.001640602, 0.001540977, 0.001437642, 0.001093965, 0.0009749447, 
    0.0009575898, 0.0009466455, 0.0008583429, 0.0007019087, 0.000591682,
  0.001969372, 0.001864054, 0.001827213, 0.001762563, 0.001694011, 
    0.001614165, 0.001536811, 0.001412467, 0.001089657, 0.001010443, 
    0.001014651, 0.0009541269, 0.0007618876, 0.0006473941, 0.0006275031,
  0.0004073874, 0.0005107169, 0.0004740721, 0.0005027748, 0.0004340613, 
    0.0005044807, 0.0006188334, 0.000599008, 0.0005433502, 0.0004235375, 
    0.0003992458, 0.0003560575, 0.0002565107, 0.0002085072, 0.000147591,
  0.0006541832, 0.0006702241, 0.0006318553, 0.0005459759, 0.000418003, 
    0.0004876664, 0.0006866258, 0.0006453819, 0.0006266379, 0.0005779359, 
    0.0004003131, 0.0004101819, 0.0003623016, 0.0002020372, 0.0001893421,
  0.0009999098, 0.0008748423, 0.0008717897, 0.0007165194, 0.0006760177, 
    0.0005079159, 0.0007202918, 0.000715833, 0.0006756208, 0.0005862821, 
    0.000501714, 0.0004573408, 0.0004207325, 0.0003758379, 0.0002813645,
  0.001226679, 0.001141382, 0.001111684, 0.001004678, 0.0009535495, 
    0.0008199952, 0.0005356367, 0.0006528233, 0.000603213, 0.0005578814, 
    0.0004979548, 0.0004475554, 0.0004138827, 0.0003930281, 0.0003847441,
  0.001315163, 0.001253072, 0.001234828, 0.001303126, 0.001311996, 
    0.001156464, 0.001065033, 0.0004814526, 0.0004228103, 0.0004726764, 
    0.0004907349, 0.0004482598, 0.0004385923, 0.000454229, 0.00045684,
  0.001427961, 0.001336003, 0.001347264, 0.001442376, 0.001484175, 
    0.001405685, 0.001287055, 0.001101972, 0.0008650123, 0.000652621, 
    0.0005190957, 0.0004920925, 0.0004804502, 0.0004933071, 0.0005077912,
  0.001579026, 0.001494256, 0.001479561, 0.001540067, 0.001588886, 
    0.001515774, 0.001426502, 0.001269408, 0.001033285, 0.0007253136, 
    0.0006055257, 0.0005441133, 0.000517192, 0.000497528, 0.0005207729,
  0.001731668, 0.001623924, 0.001585322, 0.001601228, 0.001616978, 
    0.001555127, 0.00153636, 0.00144524, 0.001002362, 0.0007510739, 
    0.0006286799, 0.0005876807, 0.0005415299, 0.0005082281, 0.0005263515,
  0.001903144, 0.001801499, 0.001742473, 0.001677367, 0.00165415, 0.00158608, 
    0.00155488, 0.001377153, 0.0009638484, 0.0007640557, 0.0006607713, 
    0.0006202154, 0.0005427513, 0.000517075, 0.0005337641,
  0.002030627, 0.001907552, 0.001804237, 0.001701253, 0.001654983, 
    0.00159922, 0.001496471, 0.001310767, 0.0008989641, 0.0007840237, 
    0.0007173171, 0.0006520152, 0.0005693614, 0.0005567972, 0.0005688053,
  0.0004303547, 0.0005326619, 0.0005326574, 0.0005586045, 0.0005672906, 
    0.0006011114, 0.0006316047, 0.000548024, 0.0004873729, 0.0003341761, 
    0.0002858212, 0.0002826518, 0.0002444095, 0.0002090949, 0.0001454625,
  0.0006786347, 0.0006983176, 0.0006924506, 0.0006323516, 0.0004721299, 
    0.0004894248, 0.0005655062, 0.0005047912, 0.0004580795, 0.0004165851, 
    0.0003427831, 0.0003741953, 0.00037416, 0.0001973809, 0.0001571866,
  0.001063292, 0.001005129, 0.0009631138, 0.0008463382, 0.0006772261, 
    0.0003279746, 0.00054142, 0.0004864706, 0.0004690681, 0.0004782249, 
    0.0004672509, 0.0004189939, 0.0004115146, 0.0003756038, 0.0002558292,
  0.001251503, 0.001249624, 0.001214031, 0.001114155, 0.001078113, 
    0.0008249928, 0.0003696456, 0.0004372478, 0.000457124, 0.0004684186, 
    0.0004530007, 0.0003985562, 0.0003967448, 0.0003607258, 0.0003565148,
  0.001354336, 0.001341466, 0.001349892, 0.001325526, 0.001329054, 
    0.001243493, 0.001000724, 0.0003344009, 0.0003012358, 0.0003811678, 
    0.0004263748, 0.0003920261, 0.0003969672, 0.0004059383, 0.0004262927,
  0.001458962, 0.001432228, 0.001424491, 0.001417033, 0.001395479, 
    0.00142582, 0.00119264, 0.0009944973, 0.0006853417, 0.0005314907, 
    0.0004457197, 0.0004134396, 0.000414441, 0.0004358093, 0.0004709706,
  0.001589975, 0.001554282, 0.001538829, 0.001518989, 0.001514671, 
    0.001499439, 0.001361248, 0.001151722, 0.000828848, 0.0005807749, 
    0.0005001341, 0.0004523921, 0.0004405593, 0.0004462778, 0.0004856369,
  0.001688718, 0.001659646, 0.001642105, 0.001627009, 0.001600607, 
    0.001539336, 0.001491547, 0.001342492, 0.0008895045, 0.0005810359, 
    0.000515798, 0.0004751439, 0.0004581274, 0.0004433861, 0.0004803547,
  0.00176017, 0.001748205, 0.001764371, 0.001727974, 0.001716216, 
    0.001592448, 0.001551704, 0.001441663, 0.000929083, 0.0005750755, 
    0.0005085748, 0.0004911426, 0.0004653758, 0.0004494547, 0.0004877269,
  0.001817578, 0.001813841, 0.001819916, 0.00175543, 0.001726169, 
    0.001603694, 0.001581057, 0.001558635, 0.000935591, 0.0006089162, 
    0.0005748129, 0.0005330728, 0.0004934762, 0.000498339, 0.0005160999,
  0.0005127306, 0.0005749416, 0.0006136285, 0.0006841084, 0.0006089194, 
    0.0005742068, 0.000535237, 0.000429338, 0.0003139288, 0.0001737405, 
    0.0001842047, 0.0002430909, 0.000240153, 0.0001845627, 0.0001208891,
  0.0006810588, 0.0007002176, 0.0007640107, 0.0008527758, 0.0005465564, 
    0.0004139814, 0.0005164683, 0.0004617228, 0.0003609374, 0.0003059128, 
    0.0002270492, 0.0003333046, 0.0004009366, 0.000175794, 0.0001179894,
  0.00115758, 0.001082612, 0.001010269, 0.001020879, 0.0008706738, 
    0.0003541229, 0.000433091, 0.0004750963, 0.0004071372, 0.0003671065, 
    0.0003308249, 0.000375557, 0.0004471321, 0.0003772949, 0.0002302658,
  0.001465496, 0.001395941, 0.001340597, 0.001261311, 0.001427426, 
    0.001050678, 0.0003086906, 0.0004182582, 0.0004326778, 0.0004176333, 
    0.0003659884, 0.0003633382, 0.0004275634, 0.0004008291, 0.0003045686,
  0.001580023, 0.001502439, 0.001463306, 0.001417994, 0.001453734, 
    0.001773983, 0.001152365, 0.0003285585, 0.0002882202, 0.000403541, 
    0.0003805824, 0.0003656714, 0.0004032585, 0.0004141425, 0.000374797,
  0.001705385, 0.001609118, 0.00153036, 0.00148323, 0.001472427, 0.001625243, 
    0.001664533, 0.001060917, 0.0006880607, 0.0006165573, 0.0004834192, 
    0.0004020072, 0.0003989803, 0.0003986054, 0.0003937005,
  0.001827581, 0.00171268, 0.001600359, 0.001549551, 0.001520419, 
    0.001551976, 0.001729217, 0.001586599, 0.001066657, 0.0007054508, 
    0.0005610836, 0.0004352505, 0.0004108092, 0.0003919176, 0.0003984916,
  0.001859566, 0.001733822, 0.001650438, 0.001605535, 0.001589191, 
    0.001584646, 0.001668806, 0.001726685, 0.001258229, 0.0007848954, 
    0.0005856288, 0.0004649977, 0.0004180476, 0.0003858688, 0.0003910066,
  0.0018702, 0.001752419, 0.001700523, 0.001668845, 0.001665621, 0.001667712, 
    0.0017311, 0.001796085, 0.001286869, 0.0007665904, 0.0005920796, 
    0.0004998082, 0.0004353566, 0.0003918699, 0.0003999998,
  0.001831736, 0.00172062, 0.001704715, 0.001718669, 0.001755595, 
    0.001824973, 0.001995602, 0.001977602, 0.001243934, 0.0008305419, 
    0.0007094428, 0.0005371905, 0.0004656737, 0.0004307771, 0.0004202875,
  0.0006322965, 0.0006231727, 0.0005519156, 0.0005999494, 0.0005706662, 
    0.0004112769, 0.0003251959, 0.0003335803, 0.0002884123, 0.0001565802, 
    0.0001812143, 0.0002466754, 0.0001911947, 0.0001567366, 9.944328e-05,
  0.0008096626, 0.0007615653, 0.0006914344, 0.0006693723, 0.0005338459, 
    0.0003507842, 0.0003428124, 0.0003357922, 0.0002942935, 0.0002578018, 
    0.0002560167, 0.0003415314, 0.0003455105, 0.0001487824, 9.119018e-05,
  0.001291418, 0.001138995, 0.0009557988, 0.0007771789, 0.0006309345, 
    0.0002707906, 0.0003394031, 0.0003394329, 0.0003040755, 0.0003157899, 
    0.0003358297, 0.0004445845, 0.0005018587, 0.0003350989, 0.0002077825,
  0.001808081, 0.001590736, 0.001435761, 0.001171531, 0.0009440146, 
    0.0005944336, 0.0002716359, 0.0003085485, 0.0003197436, 0.0003315659, 
    0.0003390249, 0.0004176011, 0.0005239177, 0.0004106844, 0.0002713884,
  0.001980488, 0.00182539, 0.001650825, 0.001490263, 0.001364868, 
    0.001173966, 0.0008764457, 0.0002887363, 0.0002322767, 0.0002995268, 
    0.0003464627, 0.0003860197, 0.0004957968, 0.0005034846, 0.0003391684,
  0.002058572, 0.001973154, 0.001786517, 0.001625386, 0.001506016, 
    0.001420674, 0.001297388, 0.0009788538, 0.0006643861, 0.0006118299, 
    0.000446722, 0.0004008396, 0.0004311253, 0.0004661773, 0.0004105966,
  0.002124534, 0.002082193, 0.001904556, 0.001739875, 0.001599889, 
    0.001513185, 0.001496438, 0.001420739, 0.00116432, 0.0008327502, 
    0.0005829454, 0.000435194, 0.0004209805, 0.0004322569, 0.0004081672,
  0.002159232, 0.002125997, 0.001952673, 0.001785281, 0.001656811, 
    0.001563771, 0.001516516, 0.001584591, 0.001513697, 0.001162049, 
    0.0007101358, 0.0004787908, 0.0004234045, 0.0003936396, 0.0003809863,
  0.002135344, 0.002128656, 0.002010815, 0.001823467, 0.001676293, 
    0.001587593, 0.001541808, 0.001581278, 0.001535262, 0.001362893, 
    0.001040132, 0.0006484551, 0.0004637388, 0.000386225, 0.000361999,
  0.002085827, 0.002098765, 0.002005548, 0.00183694, 0.001691083, 
    0.001606739, 0.001596637, 0.001723992, 0.001463401, 0.001317217, 
    0.001294283, 0.0009749298, 0.0006592514, 0.0004801042, 0.0003849557,
  0.00158845, 0.001377933, 0.0008541885, 0.0005373025, 0.0003824715, 
    0.0003146108, 0.000323176, 0.0003459796, 0.0003158007, 0.0001713678, 
    0.0001737625, 0.0001631344, 0.0001296445, 0.0001329196, 8.302342e-05,
  0.001874593, 0.001561322, 0.001051528, 0.0005817279, 0.0003722941, 
    0.000292436, 0.000326121, 0.0003456204, 0.0003299418, 0.0002641934, 
    0.0002339711, 0.0002589065, 0.0002442328, 0.0001212231, 8.409774e-05,
  0.002289322, 0.001972532, 0.001249155, 0.0006778628, 0.0004822811, 
    0.0002439988, 0.0003054616, 0.0003338121, 0.0003301409, 0.0003204297, 
    0.0003237636, 0.0003348644, 0.0003096777, 0.0002637092, 0.000178404,
  0.002478483, 0.002337811, 0.001775541, 0.001073807, 0.0007646697, 
    0.0005092127, 0.0002547379, 0.0002794756, 0.0003154978, 0.0003198836, 
    0.0003426086, 0.0003833497, 0.0003672465, 0.0003049737, 0.0002309412,
  0.002532377, 0.002489975, 0.002056215, 0.001545686, 0.001256097, 
    0.0009891891, 0.0007780224, 0.0002787478, 0.0002253275, 0.0002819333, 
    0.0003473227, 0.0004030042, 0.0004073649, 0.0003649933, 0.0002928606,
  0.002513417, 0.002525598, 0.002257532, 0.001726128, 0.001483816, 
    0.001301132, 0.001114577, 0.0008278551, 0.0005746404, 0.0005336804, 
    0.0004156426, 0.0004116021, 0.0004277247, 0.0003994276, 0.0003226194,
  0.002493319, 0.002495968, 0.00239591, 0.001847126, 0.001592779, 
    0.001435368, 0.001294059, 0.00103447, 0.0008246849, 0.0006852256, 
    0.0005418635, 0.0004400201, 0.000437693, 0.0004056235, 0.0003548785,
  0.002387463, 0.002432771, 0.002477369, 0.001989007, 0.001637984, 
    0.001528635, 0.001367236, 0.001255106, 0.0009848808, 0.0007482301, 
    0.000577055, 0.0004630541, 0.0004403637, 0.000393348, 0.0003616354,
  0.002228634, 0.002322911, 0.002481524, 0.002101625, 0.001716024, 
    0.001515864, 0.001419264, 0.001272161, 0.00101058, 0.000766686, 
    0.0006381872, 0.0005033936, 0.000449755, 0.0003854001, 0.0003442006,
  0.002056411, 0.002239886, 0.002405729, 0.002149654, 0.001777704, 
    0.001503761, 0.00135573, 0.001270329, 0.000978082, 0.0008158032, 
    0.0008165108, 0.0006756607, 0.0005218682, 0.0004325178, 0.0003647451,
  0.001788514, 0.002083512, 0.002064215, 0.001379205, 0.0007337383, 
    0.0004241287, 0.0003917962, 0.0003739761, 0.0002841234, 0.0001324584, 
    0.0001323175, 0.0001258613, 0.0001005381, 0.0001086667, 7.77211e-05,
  0.002280897, 0.002479991, 0.002305895, 0.001269693, 0.0005013824, 
    0.0003713685, 0.000363158, 0.0003495768, 0.0002770648, 0.0002186525, 
    0.0001616173, 0.0002000587, 0.0001900841, 9.789969e-05, 7.170482e-05,
  0.002570158, 0.002651348, 0.002378656, 0.001230249, 0.0005892372, 
    0.0002734232, 0.0003186292, 0.0003312869, 0.0002818084, 0.0002602013, 
    0.0002336933, 0.0002266548, 0.0002197879, 0.0001936639, 0.0001392066,
  0.002665909, 0.002745451, 0.00266172, 0.001554082, 0.0008924948, 
    0.0005761168, 0.0002488112, 0.0002677501, 0.0002747794, 0.0002601634, 
    0.0002407563, 0.0002396113, 0.0002294277, 0.0002101772, 0.0001883238,
  0.002612764, 0.002666098, 0.002758419, 0.002087655, 0.001323277, 0.0010004, 
    0.0007515568, 0.0002527315, 0.0001886493, 0.0002334275, 0.0002595131, 
    0.0002587342, 0.0002538525, 0.0002410527, 0.000231522,
  0.002556524, 0.002516488, 0.002750165, 0.002343241, 0.00167217, 
    0.001360676, 0.001068804, 0.0007332303, 0.0005039957, 0.0004524034, 
    0.000326003, 0.0002969279, 0.0002762744, 0.0002647685, 0.000242752,
  0.002448656, 0.002356928, 0.002635016, 0.002495634, 0.001820792, 
    0.001482749, 0.001214966, 0.0008595723, 0.000639924, 0.0005562777, 
    0.0004265732, 0.0003328327, 0.0003031396, 0.0002864437, 0.0002645411,
  0.002124674, 0.002171137, 0.002506094, 0.002552831, 0.001887156, 
    0.001531169, 0.001311573, 0.001111578, 0.0007839386, 0.0005395281, 
    0.000424881, 0.0003544182, 0.0003295632, 0.0003079343, 0.0002874906,
  0.001988614, 0.002119085, 0.002436906, 0.002571176, 0.001944025, 
    0.001515406, 0.001328809, 0.001195157, 0.0007543462, 0.0005386302, 
    0.0004450878, 0.0003857067, 0.0003606166, 0.0003277659, 0.0002993692,
  0.002107645, 0.002393509, 0.002553513, 0.002536366, 0.001902389, 
    0.00149546, 0.001263589, 0.001117065, 0.0006825865, 0.0005573121, 
    0.0005249615, 0.0004236083, 0.0003964195, 0.0003599145, 0.0003182816,
  0.0014721, 0.001507686, 0.001520399, 0.00162025, 0.001435081, 0.001073944, 
    0.0008217612, 0.000576797, 0.000339223, 0.0001588538, 0.0001528539, 
    0.0001399442, 0.0001159103, 0.0001203024, 8.000408e-05,
  0.001723359, 0.001677391, 0.001634382, 0.001678849, 0.00130113, 
    0.0008496913, 0.0006383686, 0.0004696124, 0.0003164354, 0.0002457236, 
    0.000181658, 0.0002154088, 0.000202649, 9.648546e-05, 6.521778e-05,
  0.00212047, 0.002068869, 0.001939861, 0.001813709, 0.001339113, 
    0.0005349072, 0.000442088, 0.000397558, 0.0002948052, 0.0002730586, 
    0.0002536751, 0.000245971, 0.000225632, 0.0001933391, 0.0001351125,
  0.002290971, 0.002257395, 0.002217982, 0.002115353, 0.00160935, 
    0.0008707701, 0.0003268787, 0.0002781323, 0.0002712007, 0.0002524453, 
    0.0002597742, 0.0002414861, 0.0002187049, 0.0001935934, 0.0001713781,
  0.002467302, 0.002431209, 0.002383968, 0.002365045, 0.001913374, 
    0.001271744, 0.0009206377, 0.0002718186, 0.0001918067, 0.0002185572, 
    0.0002555993, 0.0002451218, 0.0002220033, 0.0002071245, 0.0001972469,
  0.002457139, 0.002559354, 0.002547817, 0.002506684, 0.002215912, 
    0.001740774, 0.001341747, 0.0008794629, 0.0005413385, 0.0004347629, 
    0.0003212593, 0.0002675259, 0.0002322971, 0.0002060173, 0.000194373,
  0.002319959, 0.002519393, 0.002600126, 0.002592246, 0.002249224, 
    0.001799351, 0.001423892, 0.000940942, 0.0006402343, 0.0005589069, 
    0.0004159654, 0.0002851874, 0.0002408873, 0.000211045, 0.0001996041,
  0.002377447, 0.002466627, 0.002580328, 0.002604974, 0.002209782, 
    0.00178451, 0.001441664, 0.001114036, 0.0006937112, 0.000467519, 
    0.0003599089, 0.0002804305, 0.000241019, 0.0002142884, 0.0002098369,
  0.002183978, 0.002340618, 0.002465471, 0.002518597, 0.002118156, 
    0.00171053, 0.001404293, 0.001152458, 0.0005977495, 0.0003998225, 
    0.0003272045, 0.0002698214, 0.0002464637, 0.0002255907, 0.0002242257,
  0.002214205, 0.00232341, 0.002432878, 0.002434932, 0.001969228, 
    0.001570355, 0.001264045, 0.000937485, 0.000461581, 0.0004038838, 
    0.0003686268, 0.0002850552, 0.0002696054, 0.0002491255, 0.0002445522,
  0.001682732, 0.001637013, 0.001573536, 0.001514004, 0.001418405, 
    0.00132385, 0.001309588, 0.001134887, 0.0008546943, 0.0004394516, 
    0.000278323, 0.0002176622, 0.0001344137, 0.0001279439, 0.0001078438,
  0.002065493, 0.001952807, 0.001778976, 0.001628828, 0.001458698, 
    0.001328439, 0.00124336, 0.00103556, 0.0007671715, 0.0004976078, 
    0.0003122342, 0.0002924677, 0.0002446827, 0.0001138705, 8.886679e-05,
  0.002302187, 0.002275081, 0.002113603, 0.001784727, 0.001531687, 
    0.001039922, 0.001002856, 0.0008729914, 0.0006316206, 0.0004742864, 
    0.0003656188, 0.000334881, 0.0002887954, 0.0002416324, 0.0001799217,
  0.002351838, 0.0023164, 0.002280603, 0.002052877, 0.001708228, 0.00136983, 
    0.0005739869, 0.0004935617, 0.0004410739, 0.0003989936, 0.0003544728, 
    0.0003166939, 0.0002965113, 0.0002570392, 0.0002218883,
  0.002554665, 0.002550329, 0.002433244, 0.002210638, 0.001813459, 
    0.001562095, 0.001154278, 0.000371131, 0.0002830619, 0.0003026123, 
    0.000324561, 0.0003164102, 0.000295331, 0.0002671587, 0.0002432657,
  0.00239094, 0.002536242, 0.002603415, 0.002311832, 0.001904651, 
    0.001631405, 0.001461031, 0.0010268, 0.0007010218, 0.0005014083, 
    0.0003955241, 0.0003357001, 0.0002919812, 0.0002534097, 0.0002264192,
  0.002303933, 0.002341088, 0.002667683, 0.002386919, 0.001910156, 
    0.001659612, 0.001420807, 0.001166737, 0.0009215279, 0.0006842738, 
    0.0005194001, 0.0003404091, 0.0002818911, 0.0002345094, 0.0002211235,
  0.002495742, 0.002556324, 0.002700903, 0.002289371, 0.001924546, 
    0.001653782, 0.001481798, 0.00128762, 0.0008795908, 0.000556442, 
    0.0004503621, 0.0003206656, 0.0002716365, 0.0002224706, 0.0002203884,
  0.002694115, 0.002674519, 0.002573563, 0.002195125, 0.001862943, 
    0.001652143, 0.001574004, 0.001293028, 0.0006846573, 0.0004367235, 
    0.0003694253, 0.0002932709, 0.0002459498, 0.0002160875, 0.0002356524,
  0.002487849, 0.002401477, 0.002247307, 0.002023692, 0.001785313, 
    0.001646662, 0.001480209, 0.000820075, 0.0004333786, 0.0004049456, 
    0.0003876448, 0.0002880701, 0.0002561111, 0.0002353433, 0.0002663662,
  0.001388963, 0.001414516, 0.001342994, 0.001289736, 0.001190149, 
    0.001072975, 0.001081156, 0.001052365, 0.001031396, 0.000716695, 
    0.0006263231, 0.0005870977, 0.0004108562, 0.0003447016, 0.0002773058,
  0.002048249, 0.001826081, 0.001620185, 0.001446345, 0.001274716, 
    0.001188412, 0.001183155, 0.001098835, 0.001045177, 0.0009851148, 
    0.0007819667, 0.0007620232, 0.0005785798, 0.0002788048, 0.0002087615,
  0.002513092, 0.002522325, 0.002356638, 0.001954539, 0.001550898, 
    0.00111032, 0.001131791, 0.001079289, 0.0009477386, 0.0009374568, 
    0.000874248, 0.00075061, 0.0005664859, 0.0003852696, 0.0002522979,
  0.002599277, 0.002691265, 0.002756071, 0.002728193, 0.002217709, 
    0.00159661, 0.000864241, 0.0008034654, 0.0007419052, 0.0007506339, 
    0.0007370946, 0.0006392387, 0.0004887801, 0.0003422306, 0.0002578513,
  0.002463548, 0.002659298, 0.002767337, 0.002869544, 0.002749179, 
    0.002231137, 0.001593711, 0.0007453364, 0.0006505611, 0.000547498, 
    0.0006003301, 0.0005571686, 0.0004147899, 0.0003216909, 0.0002623099,
  0.002280655, 0.002509686, 0.002639315, 0.00287073, 0.002828708, 
    0.002301225, 0.001780605, 0.001347582, 0.001011422, 0.0008194334, 
    0.0006303372, 0.0004930773, 0.0003726489, 0.000288576, 0.0002420636,
  0.002170723, 0.002357901, 0.002712758, 0.0028019, 0.002517783, 0.001959955, 
    0.001531567, 0.001195132, 0.001011854, 0.0008831205, 0.0006940941, 
    0.0004496667, 0.0003369999, 0.0002671945, 0.0002289221,
  0.002009826, 0.002025074, 0.002054397, 0.002053303, 0.00181563, 
    0.001550847, 0.00138301, 0.001203043, 0.0008626697, 0.0007165617, 
    0.0005538819, 0.0003811897, 0.0003201945, 0.0002447026, 0.0002342846,
  0.001869195, 0.001780119, 0.001711967, 0.001627842, 0.001562279, 
    0.001442541, 0.001376767, 0.001145918, 0.0006703355, 0.000503657, 
    0.0004071661, 0.0003461873, 0.0002808864, 0.0002415118, 0.0002566103,
  0.001913085, 0.001798001, 0.001708533, 0.0016132, 0.001543768, 0.001483711, 
    0.001329945, 0.0007947728, 0.0004568266, 0.0004297218, 0.0004081008, 
    0.0003184665, 0.0002905878, 0.000278559, 0.0003277237,
  0.001633178, 0.001703297, 0.001558274, 0.00136955, 0.00113656, 
    0.0008154227, 0.0008043157, 0.0007251547, 0.0006392506, 0.0003546642, 
    0.000365503, 0.0004341379, 0.0003590252, 0.0003477817, 0.0002994717,
  0.002244129, 0.00222266, 0.002122467, 0.001873206, 0.001436732, 0.00115347, 
    0.000957703, 0.0007739895, 0.0006820089, 0.0005765987, 0.0004918765, 
    0.0005844228, 0.0005560868, 0.0003416044, 0.0002857016,
  0.002144144, 0.002421296, 0.002421959, 0.002247388, 0.001831129, 
    0.001230372, 0.001139484, 0.0009830699, 0.0007980962, 0.0007052155, 
    0.0006716324, 0.0006828617, 0.0006632307, 0.0005828509, 0.0003830774,
  0.001943731, 0.002149047, 0.00230976, 0.002511868, 0.002349092, 
    0.001725907, 0.001069632, 0.0008949384, 0.0008159694, 0.0007942463, 
    0.0007459503, 0.0007254554, 0.0006944022, 0.000618932, 0.0004291098,
  0.001848371, 0.002057046, 0.002173472, 0.002482216, 0.002503837, 
    0.002387535, 0.001598026, 0.0008226589, 0.0006935589, 0.0007783909, 
    0.0007712726, 0.0007682319, 0.0007167393, 0.0006255656, 0.0004646794,
  0.001714302, 0.001866553, 0.002034185, 0.002253935, 0.0024585, 0.002316548, 
    0.001831174, 0.001589166, 0.001343168, 0.001185896, 0.0009105777, 
    0.0008272383, 0.0007501284, 0.0005578988, 0.0004093362,
  0.001600531, 0.001647695, 0.001741822, 0.001798156, 0.00186022, 
    0.001854109, 0.001645617, 0.001490348, 0.001390704, 0.00133748, 
    0.001055671, 0.0008423261, 0.0006832257, 0.0004739259, 0.0003618706,
  0.001529175, 0.001509314, 0.001507278, 0.001496326, 0.001496301, 
    0.001478788, 0.001392712, 0.001294081, 0.001143751, 0.001110466, 
    0.0009168214, 0.0007406309, 0.0005734049, 0.0003956051, 0.0003145515,
  0.00157983, 0.001494688, 0.001463959, 0.001407707, 0.001388267, 
    0.001296814, 0.001217577, 0.001110805, 0.000714245, 0.0007108227, 
    0.0006824336, 0.0005868374, 0.0004192384, 0.0003079838, 0.0002490108,
  0.001640507, 0.001521979, 0.001446019, 0.001367549, 0.001317969, 
    0.001201844, 0.001035223, 0.000739312, 0.0005262051, 0.0004864633, 
    0.0005240488, 0.0004313963, 0.0003525126, 0.0002930302, 0.0002637699,
  0.001825624, 0.001970233, 0.001884324, 0.001883718, 0.001799833, 
    0.001628638, 0.00154712, 0.001303071, 0.0009683384, 0.0004642591, 
    0.0004352594, 0.0005026374, 0.0004316548, 0.0004116788, 0.0003708834,
  0.001862601, 0.001846504, 0.001741439, 0.001823272, 0.001762599, 
    0.001770384, 0.001655081, 0.001407683, 0.001170302, 0.0007039827, 
    0.0005388567, 0.0005775466, 0.0005175869, 0.0003317908, 0.0003114476,
  0.001569981, 0.001648873, 0.001843566, 0.001655465, 0.001671096, 
    0.001560741, 0.001531624, 0.001438145, 0.001275145, 0.001042104, 
    0.0007752518, 0.0006508117, 0.0005420355, 0.0004558194, 0.0003487959,
  0.001585949, 0.001493275, 0.001521697, 0.001620218, 0.001705728, 
    0.001673565, 0.001160805, 0.001027762, 0.0009809176, 0.0009608493, 
    0.0008045253, 0.0006467485, 0.000580003, 0.0004864785, 0.0003846252,
  0.001615025, 0.001448388, 0.001490684, 0.001525764, 0.001568582, 
    0.001572844, 0.001464087, 0.0006163863, 0.0008258751, 0.0008915081, 
    0.0008943029, 0.0007287987, 0.0006072329, 0.0005186225, 0.0004325546,
  0.001625673, 0.001465708, 0.00150165, 0.00155891, 0.001550337, 0.001482842, 
    0.001335792, 0.001178118, 0.001200199, 0.00129249, 0.001030901, 
    0.0008076152, 0.0006385343, 0.0005469909, 0.0004388696,
  0.001673672, 0.001549075, 0.001592668, 0.001642852, 0.001616161, 
    0.001522337, 0.001357075, 0.001080942, 0.001087925, 0.001296415, 
    0.001111949, 0.0007922358, 0.0006378445, 0.0005505322, 0.0004352457,
  0.00174568, 0.001653248, 0.001759408, 0.001776222, 0.001688324, 
    0.001573767, 0.001372368, 0.00110641, 0.0008940429, 0.001032962, 
    0.0009663888, 0.0007516131, 0.0006340744, 0.0005254907, 0.0004074726,
  0.00181253, 0.001810196, 0.001914657, 0.001905376, 0.001734367, 
    0.001552145, 0.001368537, 0.001050294, 0.0007910948, 0.0007781612, 
    0.0008525105, 0.0007092295, 0.0006165666, 0.0004448923, 0.000311205,
  0.001944996, 0.002070736, 0.002139593, 0.001941261, 0.00174155, 
    0.001548182, 0.001317045, 0.0009662181, 0.0006686266, 0.000520319, 
    0.0007445154, 0.0006573119, 0.0005431154, 0.0003804537, 0.0003145558,
  0.001472957, 0.001779011, 0.001209052, 0.001567627, 0.00131058, 
    0.001256714, 0.001427995, 0.001428504, 0.001394361, 0.0009766886, 
    0.0008474697, 0.0008306035, 0.0006451422, 0.0005696235, 0.0004716694,
  0.001714603, 0.001538663, 0.001405471, 0.00142028, 0.00117447, 0.001272243, 
    0.001426357, 0.001392908, 0.001403623, 0.001212161, 0.000984703, 
    0.0009689364, 0.0009061706, 0.0005844765, 0.0004516602,
  0.001694748, 0.001642511, 0.001836904, 0.001699717, 0.001483096, 
    0.001280977, 0.001463323, 0.001486243, 0.001409121, 0.001193517, 
    0.001064176, 0.001016967, 0.0008955913, 0.000755146, 0.0005445628,
  0.001824847, 0.001774293, 0.001883162, 0.002106875, 0.002219745, 
    0.002168302, 0.001829291, 0.001490546, 0.001317801, 0.001102575, 
    0.0008655043, 0.000812522, 0.0008006607, 0.0007157011, 0.0005687225,
  0.001981687, 0.002015285, 0.002148349, 0.002316578, 0.00250235, 
    0.002611069, 0.002487366, 0.001655164, 0.001166081, 0.0008692613, 
    0.0008170411, 0.0008128854, 0.0007812965, 0.0007417861, 0.0005695479,
  0.00199848, 0.002141278, 0.002343389, 0.002506057, 0.002595386, 
    0.002605857, 0.002483992, 0.002151479, 0.001492013, 0.001099722, 
    0.0008084027, 0.000821439, 0.000761422, 0.000676713, 0.0005264259,
  0.002158254, 0.002429411, 0.002552011, 0.002552578, 0.002568208, 
    0.002433668, 0.002140808, 0.001910331, 0.001545016, 0.001156262, 
    0.0008802086, 0.0006608785, 0.0006879788, 0.000635652, 0.0004923887,
  0.00242378, 0.002620025, 0.002661285, 0.002520511, 0.002448329, 
    0.002188114, 0.001748542, 0.001730407, 0.001422103, 0.0009764711, 
    0.0006948558, 0.0005453053, 0.0006412159, 0.0005553052, 0.0004550355,
  0.002689573, 0.002851184, 0.0027288, 0.002422562, 0.002320482, 0.00188613, 
    0.001523463, 0.001584294, 0.001231129, 0.0007952666, 0.0005794992, 
    0.0005495823, 0.0005819856, 0.0004701304, 0.0003760798,
  0.002989514, 0.003058385, 0.002739742, 0.00231746, 0.002188134, 
    0.001689314, 0.001355228, 0.001429447, 0.0009914414, 0.0005740112, 
    0.0005143, 0.000551186, 0.000520608, 0.0004038553, 0.000340298,
  0.001095661, 0.001275994, 0.001086177, 0.001304415, 0.00129309, 
    0.001303964, 0.001418369, 0.001392831, 0.001387196, 0.001288983, 
    0.001352431, 0.00144989, 0.001342688, 0.001191725, 0.0008221027,
  0.00149339, 0.001679571, 0.001594108, 0.001545159, 0.001437129, 
    0.001500426, 0.001513561, 0.001452901, 0.001369227, 0.001314632, 
    0.001408381, 0.001568717, 0.001475506, 0.0009608893, 0.0007112641,
  0.00199002, 0.002274055, 0.002318193, 0.002098051, 0.001785951, 
    0.001448883, 0.001534747, 0.001478943, 0.001344881, 0.001236083, 
    0.001353433, 0.00133978, 0.001146383, 0.000928239, 0.0006901833,
  0.002323939, 0.002566692, 0.002462053, 0.002235777, 0.002033039, 
    0.001546749, 0.001154212, 0.001201505, 0.001140958, 0.0009854981, 
    0.001000212, 0.0009821854, 0.0009080904, 0.0008624945, 0.0007501879,
  0.002603782, 0.002746935, 0.002461037, 0.002156901, 0.001865491, 
    0.001560786, 0.001392209, 0.0009408469, 0.0009155572, 0.0007535369, 
    0.000726137, 0.0007509474, 0.0007700869, 0.0008265372, 0.0008195732,
  0.002849808, 0.002852487, 0.00253362, 0.002180214, 0.001905473, 
    0.001544772, 0.001336011, 0.001278039, 0.0009975265, 0.0007634833, 
    0.0006175489, 0.0006762415, 0.0007756341, 0.0008630602, 0.0006907039,
  0.002947164, 0.002823755, 0.002581405, 0.002379274, 0.00205864, 
    0.001685799, 0.001426873, 0.001251774, 0.0009956722, 0.0007804204, 
    0.0006382219, 0.0005983187, 0.0006997176, 0.0006943263, 0.000525489,
  0.002922795, 0.002836222, 0.002638303, 0.002541164, 0.002209932, 
    0.001881453, 0.001572386, 0.00134701, 0.0009631332, 0.0007196489, 
    0.0005980846, 0.0005663016, 0.0005894932, 0.0004576457, 0.000424851,
  0.002874884, 0.002878371, 0.002680537, 0.002615247, 0.002356303, 
    0.001996623, 0.001741403, 0.001497311, 0.001052957, 0.0007103377, 
    0.0005609513, 0.0005030886, 0.0004708965, 0.0004122336, 0.000400987,
  0.002907881, 0.003164535, 0.002899154, 0.002707722, 0.002438292, 
    0.002133173, 0.001835675, 0.001613146, 0.001156596, 0.0006502434, 
    0.0004948576, 0.0004822298, 0.0004419921, 0.0003982688, 0.0003824709,
  0.001197677, 0.001367203, 0.001032372, 0.001107849, 0.0009416444, 
    0.0009975081, 0.001224684, 0.001134236, 0.000875624, 0.000538616, 
    0.0006449121, 0.0007816917, 0.0006717227, 0.0006297696, 0.0004957234,
  0.001721779, 0.001514848, 0.001166724, 0.001181929, 0.001033346, 
    0.001287794, 0.001371668, 0.001326521, 0.001028751, 0.0006690388, 
    0.0006384757, 0.0007671493, 0.0006882318, 0.0004462106, 0.0003786619,
  0.001921709, 0.001803494, 0.001793389, 0.001777189, 0.001513432, 
    0.001324677, 0.001639054, 0.001570825, 0.001293765, 0.0007197195, 
    0.0007008008, 0.0007671792, 0.0007075938, 0.000555385, 0.0004338996,
  0.002067305, 0.002056846, 0.002095214, 0.002265992, 0.002199524, 
    0.001982795, 0.001725738, 0.00160148, 0.001517973, 0.000904951, 
    0.000686351, 0.0007691569, 0.0007701837, 0.0005859516, 0.0004596287,
  0.002171226, 0.002197966, 0.002299535, 0.002366993, 0.002374392, 
    0.002600872, 0.002409377, 0.001816165, 0.001620059, 0.001292799, 
    0.0007036676, 0.0007206504, 0.000754267, 0.0006556228, 0.0006397484,
  0.002456779, 0.002649279, 0.002607343, 0.002472697, 0.002441725, 
    0.002634505, 0.002662151, 0.002481996, 0.002265503, 0.001836764, 
    0.0007642262, 0.0007389336, 0.000697626, 0.0005669484, 0.0004830077,
  0.002513648, 0.0025047, 0.002700668, 0.002863623, 0.002417533, 0.002569324, 
    0.002571733, 0.002655427, 0.002439778, 0.002148153, 0.001169086, 
    0.0007178773, 0.0006995433, 0.0004814119, 0.0003938702,
  0.002556482, 0.00255252, 0.00252687, 0.002731379, 0.002422567, 0.002511101, 
    0.002516737, 0.002663131, 0.00254026, 0.002317568, 0.001612485, 
    0.0008649575, 0.0006861278, 0.0004957649, 0.0003497594,
  0.00256506, 0.002492955, 0.002419111, 0.002630481, 0.002548064, 
    0.002670312, 0.002533951, 0.002581162, 0.002553971, 0.002404191, 
    0.001824761, 0.001113932, 0.0007553747, 0.0004515079, 0.0003721931,
  0.00251692, 0.002563526, 0.002627002, 0.002635289, 0.002672142, 
    0.002579404, 0.0025868, 0.002540952, 0.002559327, 0.002475011, 
    0.002007403, 0.001320984, 0.0008820249, 0.0005468515, 0.0004242188,
  0.001197214, 0.001355147, 0.001491584, 0.001934114, 0.00198742, 
    0.002089821, 0.002211505, 0.001881576, 0.0009305906, 0.0004042655, 
    0.0004558269, 0.0005422513, 0.0003705064, 0.0002797733, 0.0002449645,
  0.001444982, 0.001636731, 0.001857911, 0.002040151, 0.001918783, 
    0.002017945, 0.002123126, 0.001945465, 0.001542759, 0.0006650097, 
    0.0004300236, 0.0005784177, 0.0004907231, 0.0002291245, 0.0001887532,
  0.001857781, 0.001854562, 0.002111173, 0.002233587, 0.001925885, 
    0.001724076, 0.002024422, 0.002051316, 0.002117196, 0.001286299, 
    0.0007464121, 0.0006227792, 0.000531142, 0.0004808127, 0.0003642019,
  0.002008668, 0.002079617, 0.002058479, 0.002017011, 0.002141117, 
    0.002001902, 0.001789706, 0.001606881, 0.002180826, 0.002011778, 
    0.001197272, 0.0007688208, 0.0005788789, 0.000478075, 0.0004719683,
  0.002113499, 0.002106259, 0.002080799, 0.002016276, 0.001996096, 
    0.002094585, 0.002271587, 0.001854136, 0.002010396, 0.00224562, 
    0.001676544, 0.001250702, 0.0007151208, 0.000534448, 0.0005765051,
  0.002174111, 0.002215918, 0.002083083, 0.002018709, 0.002023786, 
    0.002086422, 0.002247155, 0.002355668, 0.002258444, 0.002310661, 
    0.002037317, 0.001702153, 0.001181243, 0.0006958183, 0.0005215818,
  0.002173523, 0.002286852, 0.002102131, 0.002114714, 0.002091902, 
    0.002164953, 0.002190666, 0.002324168, 0.002300048, 0.002278452, 
    0.002258629, 0.001897046, 0.001505223, 0.0009811496, 0.0005974316,
  0.002292191, 0.002376874, 0.002315252, 0.002320912, 0.002274765, 
    0.002327535, 0.002358803, 0.002377757, 0.002336503, 0.002260418, 
    0.00226263, 0.001998618, 0.001713606, 0.001254491, 0.0007880938,
  0.002539722, 0.002599395, 0.002612405, 0.002613745, 0.002680936, 
    0.002548986, 0.002605425, 0.00253823, 0.002409807, 0.002368011, 
    0.002316309, 0.002058317, 0.001847517, 0.001474163, 0.000988109,
  0.002650151, 0.002751037, 0.002951506, 0.002653825, 0.002591166, 
    0.002533094, 0.002527143, 0.002402727, 0.002417913, 0.002294425, 
    0.002311699, 0.002207031, 0.001895325, 0.001588009, 0.001171254,
  0.001593446, 0.001691067, 0.001627348, 0.001743715, 0.001767036, 
    0.001825449, 0.001870709, 0.001614079, 0.001296843, 0.0006878494, 
    0.000442366, 0.0004626252, 0.0002522281, 0.0002510417, 0.000220084,
  0.001818534, 0.00173924, 0.001774961, 0.001735633, 0.001558744, 
    0.001641261, 0.001563285, 0.001719643, 0.001690448, 0.001411006, 
    0.0008157885, 0.0007273052, 0.0005934549, 0.0003671588, 0.0002654229,
  0.001879734, 0.001810619, 0.001841015, 0.001796501, 0.001617912, 
    0.001274542, 0.001647446, 0.001722952, 0.001776667, 0.001719582, 
    0.001455952, 0.001190694, 0.0009654665, 0.0008246428, 0.0005868103,
  0.001908798, 0.00185153, 0.001802443, 0.001708305, 0.001816148, 
    0.001722345, 0.001529552, 0.001390313, 0.001492729, 0.001570522, 
    0.001605996, 0.001513018, 0.001336847, 0.001154325, 0.0009832438,
  0.001929536, 0.001846179, 0.001827133, 0.001834507, 0.001879059, 
    0.001934477, 0.002040659, 0.001764804, 0.001732081, 0.001675839, 
    0.001821429, 0.001863404, 0.001739217, 0.001472497, 0.001237363,
  0.001968476, 0.001928445, 0.001980172, 0.002009985, 0.002073796, 
    0.002162913, 0.002205192, 0.002342806, 0.002311826, 0.002250276, 
    0.002230828, 0.002067134, 0.002044392, 0.001881009, 0.001584682,
  0.002182157, 0.002203045, 0.002241403, 0.002288234, 0.002347143, 0.0023923, 
    0.00244018, 0.002537569, 0.002573333, 0.002493907, 0.002400056, 
    0.002230647, 0.002167428, 0.002080029, 0.001906935,
  0.0023926, 0.002449053, 0.002486793, 0.00260009, 0.002634332, 0.002669673, 
    0.002718527, 0.00282168, 0.002843264, 0.002788336, 0.002733844, 
    0.002505794, 0.002389273, 0.00227824, 0.002068375,
  0.002577102, 0.002662159, 0.002796532, 0.002858835, 0.00295013, 
    0.002887518, 0.002928641, 0.002991127, 0.003020156, 0.002986613, 
    0.00291494, 0.002767504, 0.002632319, 0.002370545, 0.002136943,
  0.002814104, 0.002919601, 0.003020798, 0.003077378, 0.00307386, 
    0.003098425, 0.003105165, 0.003088806, 0.003116458, 0.003083678, 
    0.003030586, 0.002930662, 0.002808811, 0.002522489, 0.002062878,
  0.001772866, 0.001402606, 0.001040889, 0.0009296859, 0.0007640691, 
    0.0007911069, 0.0009378688, 0.00104194, 0.001157236, 0.001084746, 
    0.001168077, 0.001255522, 0.00121886, 0.001192004, 0.00137395,
  0.001736543, 0.001541859, 0.001228013, 0.001035672, 0.0007643104, 
    0.0008898039, 0.001179414, 0.001225636, 0.001265939, 0.001255768, 
    0.001289026, 0.001513288, 0.001686879, 0.001609037, 0.001550981,
  0.001869081, 0.001685846, 0.001511011, 0.001246269, 0.0009318269, 
    0.0006911602, 0.00110331, 0.001242955, 0.001455963, 0.001579626, 
    0.001742211, 0.001980284, 0.002140824, 0.002143161, 0.002074207,
  0.002147491, 0.002056505, 0.001972743, 0.001874454, 0.001651724, 
    0.001234772, 0.001225879, 0.00149709, 0.001910407, 0.002133588, 
    0.002346538, 0.002487891, 0.00241279, 0.002305752, 0.002216694,
  0.002233656, 0.002138877, 0.002086326, 0.002061168, 0.002076982, 
    0.002139559, 0.002174383, 0.002019189, 0.002153972, 0.002416911, 
    0.002718423, 0.002677288, 0.002523999, 0.002411791, 0.002313168,
  0.002246875, 0.002210691, 0.002178535, 0.002190467, 0.002251314, 
    0.002329287, 0.00244531, 0.002550458, 0.002771603, 0.002989307, 
    0.002934063, 0.002619227, 0.002489393, 0.002391609, 0.00224623,
  0.002278314, 0.002305115, 0.002326653, 0.00233893, 0.002483877, 
    0.002593469, 0.002734248, 0.002928646, 0.003165699, 0.00309193, 
    0.002637065, 0.002453575, 0.002350894, 0.002242552, 0.002160781,
  0.002406995, 0.002447285, 0.00250544, 0.002600465, 0.00272791, 0.002855574, 
    0.003012174, 0.003180551, 0.0031747, 0.002580883, 0.002361587, 
    0.002230428, 0.002139952, 0.002049289, 0.002010199,
  0.002467615, 0.002598133, 0.002694768, 0.002779745, 0.002903272, 
    0.003030662, 0.003233615, 0.003239531, 0.002593408, 0.002190389, 
    0.002061267, 0.001945863, 0.001852684, 0.001822913, 0.001830328,
  0.002666582, 0.00277438, 0.002893725, 0.003008143, 0.00313591, 0.003286332, 
    0.00330771, 0.002538147, 0.002054518, 0.001770506, 0.001785299, 
    0.001709125, 0.001665755, 0.00166437, 0.001619376,
  0.001750855, 0.001598393, 0.001276566, 0.0010787, 0.0008386324, 
    0.0006914485, 0.000743359, 0.0006351423, 0.0005809816, 0.0005116706, 
    0.0006020249, 0.0008594726, 0.00114534, 0.001327774, 0.00105734,
  0.001935506, 0.001870246, 0.001501591, 0.001191292, 0.000827459, 
    0.0007384188, 0.0008289882, 0.0007131753, 0.0006897079, 0.0006646268, 
    0.0007517918, 0.001192625, 0.0014953, 0.001152159, 0.0008672056,
  0.002008689, 0.001959585, 0.001848724, 0.001527324, 0.0009636477, 
    0.000724673, 0.0009610312, 0.0009907881, 0.000952001, 0.0009066963, 
    0.001081674, 0.001458096, 0.001435402, 0.001134346, 0.00085743,
  0.00214138, 0.002200679, 0.00218685, 0.002100584, 0.001696112, 0.001036651, 
    0.0008593376, 0.0009763405, 0.001167889, 0.001210758, 0.001509643, 
    0.001658004, 0.001371972, 0.001209727, 0.0009835846,
  0.002221899, 0.002201303, 0.002205901, 0.002198073, 0.00219429, 
    0.002138321, 0.001683887, 0.001172503, 0.00112381, 0.001525934, 
    0.001929331, 0.001758089, 0.001523187, 0.001386886, 0.001219137,
  0.002220121, 0.002233843, 0.002252691, 0.002292186, 0.002302935, 
    0.002297713, 0.002277185, 0.002068288, 0.001869838, 0.002050433, 
    0.002138217, 0.001881287, 0.001712807, 0.001516737, 0.001267293,
  0.002249029, 0.002289985, 0.002272281, 0.002264506, 0.00227442, 
    0.002276799, 0.00230639, 0.002360515, 0.002369057, 0.002398715, 
    0.002223886, 0.001959434, 0.001762885, 0.001528219, 0.001278595,
  0.002232117, 0.002268502, 0.002265068, 0.002267782, 0.002305454, 
    0.002320343, 0.002362769, 0.002472159, 0.002454048, 0.00239874, 
    0.002203712, 0.001948179, 0.001721602, 0.001470249, 0.001251808,
  0.002293395, 0.002256599, 0.002267646, 0.002310849, 0.002351591, 
    0.002442947, 0.002492506, 0.002531758, 0.002554247, 0.002427534, 
    0.002221591, 0.001932882, 0.00170089, 0.001430484, 0.001234371,
  0.002376693, 0.002321689, 0.002294132, 0.002330602, 0.002461746, 
    0.002545764, 0.002508414, 0.00254305, 0.002509065, 0.002256683, 
    0.002154258, 0.001881943, 0.001610451, 0.001354296, 0.001160674,
  0.001960485, 0.001944831, 0.001922286, 0.001962247, 0.001853736, 
    0.001700818, 0.001652761, 0.001358963, 0.001062729, 0.0006040452, 
    0.0004800328, 0.0005064311, 0.0004173317, 0.0003749656, 0.0003461389,
  0.002023904, 0.002065046, 0.00205142, 0.002074284, 0.001913461, 
    0.001730885, 0.001712736, 0.001403375, 0.001077349, 0.0008645827, 
    0.0007105546, 0.0007028715, 0.0006466308, 0.0004630618, 0.0004558688,
  0.002089819, 0.002147558, 0.002239011, 0.002253696, 0.002099026, 
    0.001667182, 0.001758157, 0.001607037, 0.001173684, 0.001072775, 
    0.001042602, 0.001005401, 0.0009466298, 0.0009817573, 0.0009528702,
  0.002258996, 0.002286192, 0.002377956, 0.002457297, 0.002500994, 
    0.002067391, 0.001671364, 0.001525894, 0.001414592, 0.001376944, 
    0.001361405, 0.001335749, 0.001397205, 0.001263701, 0.001017184,
  0.002395622, 0.002437117, 0.002530087, 0.002629683, 0.002657337, 
    0.002711355, 0.002365196, 0.001574322, 0.001532683, 0.00166854, 
    0.001913792, 0.001804035, 0.001565951, 0.001140918, 0.001008547,
  0.00267457, 0.002722523, 0.002775104, 0.002765519, 0.002702647, 
    0.002599235, 0.002657761, 0.002396017, 0.002174356, 0.002099049, 
    0.002228572, 0.001974961, 0.001402621, 0.001120014, 0.00103162,
  0.003043597, 0.003010023, 0.002921917, 0.002782535, 0.00268445, 
    0.002531709, 0.002439101, 0.002552352, 0.002283718, 0.002372294, 
    0.002075938, 0.001508039, 0.001124136, 0.0009631194, 0.000906623,
  0.003321502, 0.003216061, 0.003025287, 0.002769663, 0.002695115, 
    0.002425398, 0.002442812, 0.002523849, 0.0025434, 0.002180337, 
    0.001476662, 0.001073287, 0.000883735, 0.0007847676, 0.0007593411,
  0.003524161, 0.003257733, 0.00304096, 0.002846039, 0.002643629, 
    0.002516338, 0.00241677, 0.002591808, 0.002289978, 0.001768746, 
    0.001326027, 0.0008870054, 0.0007161392, 0.0006264119, 0.0006236268,
  0.00342256, 0.003314827, 0.003068473, 0.002751345, 0.002627253, 
    0.002377786, 0.002450461, 0.002154013, 0.001714137, 0.001257628, 
    0.001129085, 0.0008380304, 0.0006295195, 0.0005318927, 0.0005016471,
  0.001588472, 0.001774826, 0.001774676, 0.002098376, 0.002137193, 
    0.002313338, 0.002519681, 0.002559268, 0.002417641, 0.001973553, 
    0.001568504, 0.001355379, 0.0009493666, 0.0007248968, 0.0005014867,
  0.001993761, 0.002074482, 0.002314406, 0.002575756, 0.002544312, 
    0.002740597, 0.00286771, 0.002747931, 0.002487748, 0.00196996, 
    0.001706284, 0.00154847, 0.001298228, 0.0008348296, 0.0006535889,
  0.002533752, 0.002765682, 0.002863808, 0.003004603, 0.003048887, 
    0.002982263, 0.002962776, 0.002834182, 0.002492107, 0.002057717, 
    0.001883059, 0.001708569, 0.001540821, 0.001362951, 0.00107536,
  0.002824835, 0.003230144, 0.003255719, 0.003272318, 0.003347853, 
    0.003313923, 0.00302131, 0.002759036, 0.002418464, 0.002150357, 
    0.001940264, 0.001800891, 0.001734328, 0.00160203, 0.001418969,
  0.003305302, 0.003396617, 0.003404716, 0.003481546, 0.003465274, 
    0.003399444, 0.003279729, 0.002640268, 0.002428049, 0.00219665, 
    0.00223483, 0.002159958, 0.001997365, 0.001790676, 0.001569078,
  0.003579899, 0.003648521, 0.003665603, 0.003607717, 0.003556737, 
    0.003409417, 0.003229641, 0.00297577, 0.002773766, 0.00254808, 
    0.002369616, 0.002268093, 0.002122728, 0.001876879, 0.001468046,
  0.003941685, 0.003963031, 0.003864956, 0.003663966, 0.003556926, 
    0.003322246, 0.003119535, 0.002961068, 0.002649402, 0.002420326, 
    0.002252298, 0.002257218, 0.002034086, 0.001622718, 0.001104079,
  0.004009501, 0.004026616, 0.003927781, 0.00367785, 0.003495376, 
    0.003248008, 0.003031377, 0.00288851, 0.002682655, 0.002529255, 
    0.002433971, 0.002202735, 0.001754963, 0.00111715, 0.0007829082,
  0.004198727, 0.004144677, 0.003959814, 0.003629117, 0.003351001, 
    0.003184733, 0.003032312, 0.002815964, 0.002619787, 0.002578524, 
    0.002474533, 0.001795717, 0.001100163, 0.0007645632, 0.0006283305,
  0.004123782, 0.003941381, 0.003715003, 0.003438132, 0.003262762, 
    0.003083427, 0.002856343, 0.002720001, 0.002718594, 0.002464062, 
    0.001949873, 0.001120284, 0.0007661739, 0.0005443532, 0.000448117,
  0.001047509, 0.001288099, 0.001364413, 0.001621857, 0.001772813, 
    0.002087987, 0.002313684, 0.002383074, 0.002251777, 0.002039941, 
    0.001972315, 0.002053547, 0.001888582, 0.001966638, 0.001907242,
  0.00155277, 0.001677634, 0.00176118, 0.001797771, 0.001927296, 0.002352315, 
    0.002433396, 0.002341313, 0.002240142, 0.002073635, 0.002005829, 
    0.002063125, 0.002170867, 0.0022024, 0.002143758,
  0.001928178, 0.002157965, 0.002280511, 0.002163662, 0.002415063, 
    0.002338186, 0.00255738, 0.002413387, 0.002272636, 0.002170541, 
    0.002256514, 0.002391959, 0.002598554, 0.002618704, 0.002463378,
  0.002178746, 0.002400769, 0.002566375, 0.002735169, 0.00270949, 
    0.002763308, 0.002640874, 0.002546361, 0.002448086, 0.002411182, 
    0.002545675, 0.002715121, 0.002784051, 0.002753249, 0.002246657,
  0.00243137, 0.002550601, 0.00269103, 0.002815981, 0.002905346, 0.002942261, 
    0.002964036, 0.002597491, 0.002552524, 0.002652856, 0.002830755, 
    0.002871684, 0.002896295, 0.002763978, 0.002056276,
  0.002632642, 0.002747111, 0.002889529, 0.002976718, 0.003079781, 
    0.003098352, 0.003105533, 0.00304594, 0.002954113, 0.002966054, 
    0.002915557, 0.002891133, 0.002915306, 0.002615465, 0.001741265,
  0.002952303, 0.003038112, 0.003118195, 0.00315968, 0.003171318, 
    0.003195748, 0.003171562, 0.00311522, 0.003036616, 0.00290769, 
    0.002825963, 0.002857188, 0.002886249, 0.002184664, 0.001261524,
  0.00314072, 0.003173252, 0.003248189, 0.003274191, 0.003294231, 
    0.003272262, 0.003188645, 0.003145796, 0.003039936, 0.002919001, 
    0.002837927, 0.002955772, 0.002657921, 0.00144657, 0.0007337006,
  0.003322209, 0.003405735, 0.003460829, 0.003450434, 0.003370269, 
    0.003281274, 0.003248629, 0.003158733, 0.003044214, 0.002947619, 
    0.002994221, 0.0029268, 0.001880427, 0.0007447009, 0.0004806179,
  0.003526863, 0.003518667, 0.003521134, 0.003416957, 0.003350389, 
    0.003273872, 0.003158616, 0.002982339, 0.002939658, 0.002894537, 
    0.003000979, 0.002452421, 0.000940351, 0.0004665662, 0.0003691338,
  0.0008801502, 0.001001508, 0.001005879, 0.001090868, 0.0009811004, 
    0.000972425, 0.001227312, 0.001324864, 0.001516275, 0.00166931, 
    0.001788269, 0.00193053, 0.001944254, 0.002003195, 0.002062151,
  0.001376716, 0.001422939, 0.001326226, 0.001211518, 0.001093285, 
    0.001433928, 0.001748564, 0.001787885, 0.001949251, 0.002034108, 
    0.002081443, 0.002112863, 0.002041577, 0.00202607, 0.002239654,
  0.001864826, 0.001947779, 0.002004821, 0.001951326, 0.002033918, 
    0.001938231, 0.00213525, 0.002188836, 0.002163102, 0.002110056, 
    0.00203874, 0.002074662, 0.002242444, 0.002565322, 0.0028116,
  0.00205062, 0.002190684, 0.00228543, 0.002327912, 0.002315867, 0.002290588, 
    0.002235152, 0.00231006, 0.002246781, 0.002025803, 0.002142826, 
    0.00236432, 0.002674421, 0.002882431, 0.002894473,
  0.002244209, 0.002288918, 0.002353252, 0.002387139, 0.002422053, 
    0.002492019, 0.002545631, 0.002298847, 0.00223646, 0.002386164, 
    0.002690165, 0.002816898, 0.002932451, 0.002972029, 0.002881972,
  0.002382588, 0.002430358, 0.002448343, 0.002458596, 0.002532599, 
    0.00264489, 0.002728842, 0.002765644, 0.002772581, 0.002846011, 
    0.002940095, 0.002998096, 0.003011358, 0.003007712, 0.002717651,
  0.002593942, 0.002608728, 0.002605445, 0.002655468, 0.002749395, 
    0.002823302, 0.002888463, 0.002967464, 0.003020797, 0.003051804, 
    0.003072675, 0.003072312, 0.003051559, 0.002990696, 0.00232737,
  0.002772795, 0.002772296, 0.002810969, 0.002909334, 0.003014968, 
    0.003078501, 0.003121079, 0.00316237, 0.003179231, 0.003173402, 
    0.003151679, 0.003124431, 0.003108229, 0.002801764, 0.002010711,
  0.003011542, 0.003040434, 0.003121624, 0.003163913, 0.003181742, 
    0.003197023, 0.003217041, 0.003232011, 0.003248667, 0.003251657, 
    0.003241901, 0.003186053, 0.003092036, 0.002529621, 0.001733446,
  0.003368257, 0.003356701, 0.003371887, 0.003319924, 0.00327297, 
    0.003251001, 0.003243379, 0.003238443, 0.003269994, 0.003296311, 
    0.00326756, 0.003222377, 0.002904851, 0.002252904, 0.001523831,
  0.0008100203, 0.0008952832, 0.0009323322, 0.0009914668, 0.000906995, 
    0.0009080417, 0.001018886, 0.0009500477, 0.0009801154, 0.001035106, 
    0.001167748, 0.001277723, 0.001377032, 0.001504743, 0.001611394,
  0.001318794, 0.001185859, 0.001060734, 0.001000163, 0.0008580679, 
    0.001087316, 0.001245199, 0.001292281, 0.001341114, 0.00141453, 
    0.001519589, 0.001638304, 0.001749614, 0.001778337, 0.001875827,
  0.001822979, 0.00195242, 0.001913018, 0.001717122, 0.001301007, 0.00127345, 
    0.001652239, 0.00174339, 0.001764977, 0.001760116, 0.001777395, 
    0.001863443, 0.001962574, 0.002045486, 0.002153202,
  0.001962075, 0.002059679, 0.002108631, 0.002171325, 0.002126143, 
    0.001797347, 0.00169773, 0.00191704, 0.001994479, 0.002028047, 
    0.002002182, 0.001957507, 0.002055024, 0.002139177, 0.002250352,
  0.002171496, 0.002181932, 0.002216537, 0.002272906, 0.002268782, 
    0.002350881, 0.002304538, 0.001991747, 0.001933358, 0.00204678, 
    0.0022561, 0.002128389, 0.002156018, 0.002294016, 0.002295026,
  0.002329641, 0.002347745, 0.002342887, 0.002312512, 0.002310451, 
    0.002319652, 0.002393399, 0.002430407, 0.002275598, 0.002286099, 
    0.00233805, 0.002286935, 0.002309131, 0.00241286, 0.002507863,
  0.002494061, 0.002489203, 0.002481912, 0.002431952, 0.002423706, 
    0.002406357, 0.002424648, 0.002516962, 0.002557571, 0.002490954, 
    0.002443166, 0.002411402, 0.00247475, 0.002541267, 0.002629094,
  0.002472667, 0.002486888, 0.002470376, 0.002502193, 0.002547694, 
    0.002547806, 0.002555714, 0.002581456, 0.002625669, 0.002591572, 
    0.002536954, 0.002517168, 0.002531239, 0.002561337, 0.002665637,
  0.002394536, 0.002415875, 0.002458399, 0.002570771, 0.00270569, 0.00277769, 
    0.002794588, 0.002780998, 0.002733167, 0.002723972, 0.002725287, 
    0.002636716, 0.002655662, 0.002669635, 0.002716418,
  0.002070188, 0.002079196, 0.002145875, 0.002305816, 0.002471309, 
    0.002668273, 0.002820028, 0.002950295, 0.002997495, 0.002950223, 
    0.002946792, 0.002926121, 0.002892, 0.002861783, 0.002836911,
  0.0008246755, 0.0008893264, 0.0009353479, 0.0009928164, 0.000849131, 
    0.0007936718, 0.0008583909, 0.0007366468, 0.0006071838, 0.000566079, 
    0.0005892422, 0.0006184601, 0.0005825044, 0.0005804308, 0.0005868389,
  0.00115782, 0.0009875314, 0.0009330808, 0.0008850403, 0.0007544952, 
    0.0009574367, 0.001034153, 0.0009207142, 0.0007377438, 0.0006556678, 
    0.000680143, 0.0007400432, 0.0007384444, 0.0006670719, 0.0007107087,
  0.001750788, 0.001715117, 0.001567614, 0.00129312, 0.0008112721, 
    0.0007363309, 0.001214637, 0.001237728, 0.001069593, 0.0008299568, 
    0.0008559303, 0.0008756873, 0.0008593259, 0.0008701875, 0.0009202625,
  0.00204233, 0.002035413, 0.002008862, 0.002005013, 0.001857375, 
    0.001129926, 0.001002416, 0.001371403, 0.001525366, 0.00139511, 
    0.00125346, 0.001249254, 0.001270684, 0.00133849, 0.001366016,
  0.00210382, 0.002213388, 0.002242836, 0.002225348, 0.002178255, 
    0.002170708, 0.001757788, 0.001321546, 0.001351233, 0.001554393, 
    0.001762245, 0.001768813, 0.001770743, 0.00180062, 0.001786079,
  0.001828849, 0.001962623, 0.002151127, 0.002257589, 0.002308823, 
    0.002370862, 0.002430414, 0.002232893, 0.001781031, 0.001753898, 
    0.001806478, 0.00195483, 0.002003382, 0.002033291, 0.002040034,
  0.001535335, 0.001520672, 0.001516003, 0.001539525, 0.001635645, 
    0.001750484, 0.001887824, 0.002078247, 0.002196247, 0.002089617, 
    0.002171755, 0.002207063, 0.002241612, 0.00223625, 0.002180899,
  0.00141805, 0.001344841, 0.001306063, 0.001294556, 0.001356332, 
    0.001485929, 0.001649091, 0.001846832, 0.002008264, 0.002018386, 
    0.002159987, 0.002205206, 0.002268927, 0.002299136, 0.002277666,
  0.001366389, 0.001264412, 0.001173152, 0.001096256, 0.001092338, 
    0.00118924, 0.0014406, 0.001733526, 0.001926292, 0.002048135, 
    0.002196193, 0.002223044, 0.002236057, 0.002224038, 0.002214779,
  0.001321925, 0.001205912, 0.001120222, 0.001042289, 0.000976963, 
    0.0009573312, 0.001009081, 0.001107625, 0.001583638, 0.001864772, 
    0.002168621, 0.002300651, 0.002141848, 0.002223133, 0.002283322,
  0.0009777204, 0.0009922357, 0.0010096, 0.001068382, 0.001030131, 
    0.001039245, 0.001094834, 0.0009636332, 0.0008454649, 0.0007253094, 
    0.000675974, 0.0007171768, 0.0006091589, 0.0005621969, 0.0004727418,
  0.001381529, 0.001135869, 0.001037232, 0.0009962376, 0.00089325, 
    0.001083333, 0.001125187, 0.001050117, 0.0008904628, 0.0008022611, 
    0.0007942883, 0.0008191938, 0.0007305196, 0.0005501655, 0.0004726195,
  0.002116481, 0.002057527, 0.00184094, 0.001445352, 0.001013503, 
    0.0008742471, 0.001190825, 0.001174345, 0.001066863, 0.0008577434, 
    0.0009086686, 0.0008512791, 0.0007646254, 0.0006441908, 0.0005369551,
  0.001828266, 0.001939877, 0.002087782, 0.002243678, 0.002014847, 
    0.001179744, 0.0009624924, 0.001248945, 0.00127586, 0.001171617, 
    0.001045071, 0.0009954328, 0.0008682815, 0.0008051965, 0.0006746216,
  0.001505742, 0.001551537, 0.001715002, 0.001870686, 0.002099599, 
    0.002181376, 0.001514756, 0.001036088, 0.0009970228, 0.001227543, 
    0.001413033, 0.001274461, 0.001064967, 0.0008964101, 0.0007596684,
  0.001454884, 0.00136734, 0.001414689, 0.001627589, 0.001786879, 
    0.001902737, 0.002055048, 0.001804877, 0.001410361, 0.001249282, 
    0.001383301, 0.001498165, 0.001537835, 0.00149346, 0.001397758,
  0.001455379, 0.001354475, 0.001291382, 0.0012865, 0.001313004, 0.001368963, 
    0.001548057, 0.001668056, 0.00177021, 0.001702451, 0.001732766, 
    0.001686848, 0.001707501, 0.001742187, 0.001761489,
  0.001525907, 0.001383812, 0.001265232, 0.001229882, 0.00118503, 
    0.001212742, 0.001176248, 0.001146552, 0.00117367, 0.001080053, 
    0.001017958, 0.0009365601, 0.000913711, 0.0009225557, 0.0009751134,
  0.00156496, 0.001426305, 0.001292589, 0.001183335, 0.001127522, 
    0.001079778, 0.001086587, 0.001059863, 0.000954217, 0.0008592362, 
    0.0009622464, 0.0008682274, 0.0008229208, 0.000777343, 0.0008224346,
  0.001553982, 0.00141275, 0.001270753, 0.001162036, 0.001080406, 
    0.0009893312, 0.0007876516, 0.0006332809, 0.0006365567, 0.0006158061, 
    0.0007633237, 0.0007142038, 0.000719753, 0.0007774472, 0.0009182403,
  0.001031637, 0.001078921, 0.001053107, 0.001071543, 0.0010248, 0.001063435, 
    0.00109149, 0.0010663, 0.0009849933, 0.0008165739, 0.0007795118, 
    0.0008028967, 0.0007651369, 0.0007258549, 0.0007035244,
  0.001647054, 0.001459637, 0.001228868, 0.001101321, 0.0009372259, 
    0.001095976, 0.001144442, 0.001108415, 0.001043928, 0.0009636599, 
    0.0009318426, 0.0008996411, 0.0008398609, 0.0007163387, 0.0006910202,
  0.002163815, 0.002196257, 0.002064571, 0.001769975, 0.001147023, 
    0.0009718311, 0.001240498, 0.00122292, 0.00117427, 0.001062473, 
    0.001067672, 0.0009926135, 0.0009017125, 0.0008322666, 0.0007494094,
  0.00211809, 0.001969862, 0.001934448, 0.002023401, 0.002041718, 
    0.001328098, 0.001071227, 0.001354568, 0.001380673, 0.00129725, 
    0.001250321, 0.001154025, 0.001035107, 0.0009432147, 0.0008435753,
  0.001977896, 0.001828498, 0.001735397, 0.001612781, 0.001658326, 
    0.002049331, 0.001693933, 0.001211065, 0.001186787, 0.001300899, 
    0.001458611, 0.001359443, 0.001238257, 0.001092543, 0.0009915996,
  0.001832272, 0.001710116, 0.001634319, 0.001548423, 0.001420212, 
    0.001420081, 0.001608435, 0.001719164, 0.00154898, 0.001276452, 
    0.001286283, 0.001311247, 0.001257947, 0.001224568, 0.001171076,
  0.001691649, 0.001628057, 0.001557416, 0.001407107, 0.001329884, 
    0.001324632, 0.001302527, 0.001317781, 0.00135855, 0.001418766, 
    0.001439241, 0.00143674, 0.001434823, 0.001353435, 0.001163656,
  0.001606051, 0.001522141, 0.001402568, 0.001309756, 0.001204515, 
    0.001178665, 0.001118663, 0.001075575, 0.000999607, 0.0008793192, 
    0.0009347954, 0.0008883191, 0.0008943662, 0.000872609, 0.0008111453,
  0.001498174, 0.001397945, 0.001290293, 0.001151064, 0.001021745, 
    0.0009367861, 0.0008688696, 0.000786986, 0.0006844208, 0.0006530259, 
    0.00070133, 0.0006297463, 0.0006832753, 0.000627748, 0.0005855297,
  0.001364119, 0.001203044, 0.001104122, 0.0009486931, 0.0007883804, 
    0.0006518768, 0.0005320814, 0.0004878597, 0.000485826, 0.00046201, 
    0.0005057855, 0.0004639231, 0.0004536689, 0.000435992, 0.0005245095,
  0.001124005, 0.001184177, 0.001127027, 0.001099218, 0.001008004, 
    0.0009615598, 0.001018064, 0.0009604082, 0.0008896826, 0.0006474645, 
    0.0007011953, 0.0007173775, 0.0006238603, 0.0005524, 0.0005091423,
  0.001798441, 0.001595143, 0.001356591, 0.001152974, 0.001026137, 
    0.001073494, 0.001093523, 0.0009982253, 0.0008828876, 0.0007495491, 
    0.0007935766, 0.0008337779, 0.0007726974, 0.0005935198, 0.0005811156,
  0.001956433, 0.002040443, 0.00205877, 0.001752255, 0.001196175, 
    0.0009549785, 0.001224809, 0.001162212, 0.001020735, 0.0007820245, 
    0.0008836493, 0.0008749249, 0.0008097648, 0.000742314, 0.0006470495,
  0.001730715, 0.001766109, 0.001990241, 0.002212265, 0.002112199, 
    0.001267125, 0.001042771, 0.001296148, 0.001288361, 0.001080241, 
    0.0009892273, 0.0009379369, 0.0008491293, 0.0008393113, 0.0007632701,
  0.001538926, 0.001616457, 0.001701765, 0.001854641, 0.002046308, 
    0.002057023, 0.00146854, 0.001117792, 0.001075643, 0.001204158, 
    0.001235842, 0.001106623, 0.0009858847, 0.0009102043, 0.000831659,
  0.001530808, 0.00147338, 0.001381856, 0.001428318, 0.001584399, 
    0.001710104, 0.001750985, 0.001626036, 0.001379075, 0.001274117, 
    0.001270792, 0.001224259, 0.001116193, 0.001019192, 0.0009187168,
  0.001501546, 0.001317317, 0.001125773, 0.001086937, 0.001156996, 
    0.001268087, 0.001361523, 0.001413152, 0.001329862, 0.001311294, 
    0.001302114, 0.00124221, 0.001215045, 0.001134148, 0.0010527,
  0.001435433, 0.001199428, 0.0009967335, 0.0008954843, 0.0008624331, 
    0.0008739527, 0.0008782568, 0.000867256, 0.0007282804, 0.0007116045, 
    0.0009463611, 0.0009955278, 0.001029279, 0.001011559, 0.0009894335,
  0.001438805, 0.001149261, 0.0009552732, 0.0008380873, 0.0007513899, 
    0.0006829017, 0.0006340738, 0.0005548009, 0.0004903829, 0.0004995267, 
    0.0006013149, 0.000595572, 0.0006433064, 0.0006683168, 0.0007205412,
  0.001531761, 0.001145021, 0.0009218964, 0.0007552583, 0.0006606437, 
    0.0005409879, 0.0004384156, 0.000381423, 0.0003593895, 0.0003951254, 
    0.0003990389, 0.0003586819, 0.0003600371, 0.0004120469, 0.0004813702,
  0.001513367, 0.001459134, 0.001321708, 0.001280318, 0.001092225, 
    0.001004572, 0.001009953, 0.0009071754, 0.0008565169, 0.0006424931, 
    0.000631003, 0.000641009, 0.000464669, 0.0004050213, 0.0003295533,
  0.00184346, 0.001682404, 0.001508933, 0.001379783, 0.001112532, 
    0.001211294, 0.001195704, 0.00102517, 0.0008816154, 0.0008020084, 
    0.0007408521, 0.0007720058, 0.0006690788, 0.0004420313, 0.0003696006,
  0.002231688, 0.002012162, 0.001893591, 0.001679561, 0.001362755, 
    0.00110365, 0.001323289, 0.00127458, 0.001066745, 0.0008352044, 
    0.0008961793, 0.0008616488, 0.0007546059, 0.0006460577, 0.0004815561,
  0.00235878, 0.002035244, 0.001769686, 0.001699915, 0.001886989, 0.00150206, 
    0.001164514, 0.001338573, 0.001321245, 0.001085547, 0.0009549256, 
    0.0009181504, 0.0008431481, 0.0007503408, 0.0006149282,
  0.002360238, 0.001982094, 0.001588808, 0.001271087, 0.001328758, 
    0.001743409, 0.001572792, 0.001162534, 0.0009261962, 0.001155164, 
    0.001207597, 0.001045168, 0.0009525534, 0.0008577945, 0.0006955179,
  0.002257422, 0.001884489, 0.0013773, 0.001096306, 0.001197373, 0.001302951, 
    0.001443614, 0.001361617, 0.001040083, 0.000919417, 0.001030425, 
    0.001110933, 0.001003543, 0.0009166485, 0.0007584455,
  0.002107692, 0.00179764, 0.001327329, 0.001035088, 0.0009496295, 
    0.00100475, 0.001079648, 0.001062638, 0.0008388747, 0.0007567674, 
    0.0009059209, 0.0009928219, 0.0009949782, 0.0009189517, 0.0008316161,
  0.00205895, 0.001690806, 0.001252141, 0.001083073, 0.00101323, 
    0.0009905124, 0.0009115019, 0.0007814025, 0.0005954111, 0.0005841488, 
    0.0006417083, 0.000780144, 0.0009804411, 0.0009222892, 0.0008476617,
  0.001925496, 0.001561921, 0.001248531, 0.001094768, 0.001076856, 
    0.0009720977, 0.0008009498, 0.000630435, 0.0004906472, 0.0004369125, 
    0.0005006593, 0.0005011008, 0.0007617266, 0.0009096746, 0.0008466841,
  0.00141365, 0.001240138, 0.001056993, 0.0008851796, 0.0007644636, 
    0.0005669782, 0.000440639, 0.0003769642, 0.0003227428, 0.0003183137, 
    0.0003547644, 0.0003599271, 0.000550886, 0.000844863, 0.0008592446,
  0.001826258, 0.001908918, 0.001801293, 0.001656003, 0.001351493, 
    0.001118346, 0.001133909, 0.0009926257, 0.001005993, 0.0007707268, 
    0.0007834131, 0.0007594606, 0.0005511739, 0.0004351646, 0.000330007,
  0.001831241, 0.001899765, 0.001835895, 0.0016522, 0.001323154, 0.001271521, 
    0.001218525, 0.001086951, 0.001018705, 0.0009946499, 0.000893696, 
    0.0008952506, 0.0007479794, 0.0004916351, 0.0003735546,
  0.001959231, 0.001951278, 0.001868728, 0.001707142, 0.001342921, 
    0.001090411, 0.001257786, 0.001206289, 0.001077756, 0.0009362994, 
    0.001065933, 0.001020845, 0.0008768063, 0.0006939523, 0.0005042367,
  0.002095855, 0.002053602, 0.001948363, 0.001851084, 0.001512274, 
    0.001158463, 0.0009941767, 0.001235649, 0.001234307, 0.001039193, 
    0.001008579, 0.0009948205, 0.000952181, 0.0008437853, 0.0006535426,
  0.00221815, 0.002055366, 0.001895056, 0.001797731, 0.001692708, 
    0.001500816, 0.001266031, 0.00104029, 0.001025851, 0.001119205, 
    0.00115601, 0.001026615, 0.0009408502, 0.0009249815, 0.0008114635,
  0.002214983, 0.001989402, 0.001826739, 0.001625427, 0.001446402, 
    0.00145774, 0.001582167, 0.001422358, 0.001080628, 0.001026541, 
    0.001020906, 0.001094446, 0.0009931289, 0.000890463, 0.0008166145,
  0.002127401, 0.001930876, 0.001717948, 0.001486867, 0.00134603, 
    0.001245398, 0.001351469, 0.001521529, 0.00133741, 0.001065181, 
    0.000839002, 0.0007307331, 0.0007865172, 0.000787377, 0.00077521,
  0.002140985, 0.001913104, 0.001673541, 0.001426211, 0.001292589, 
    0.001238636, 0.001274567, 0.001351313, 0.001227911, 0.0009232637, 
    0.0006937421, 0.000593739, 0.000509167, 0.0004786184, 0.0005389614,
  0.001889191, 0.001632558, 0.00135387, 0.001097598, 0.0009838481, 
    0.0009865612, 0.001214505, 0.001329983, 0.001135379, 0.0008360263, 
    0.0006330571, 0.0004894103, 0.0004011955, 0.0003563526, 0.0003892047,
  0.001378313, 0.001195898, 0.0009695489, 0.0006921684, 0.0005644907, 
    0.0005150688, 0.0006496388, 0.000821265, 0.0007343219, 0.0005881364, 
    0.0004411548, 0.0003468173, 0.0003225182, 0.0003300517, 0.0003895741,
  0.001292302, 0.001674844, 0.001760545, 0.001864769, 0.001851336, 
    0.001771941, 0.001709454, 0.001415967, 0.001171751, 0.0008575801, 
    0.0007151788, 0.0005971566, 0.0004186329, 0.0003904151, 0.0004069933,
  0.001495096, 0.00164677, 0.001740364, 0.001748915, 0.001642878, 
    0.001861636, 0.001857576, 0.001505168, 0.00121476, 0.0009464971, 
    0.0008044792, 0.0007752152, 0.0006304414, 0.0003608857, 0.0003829453,
  0.001506374, 0.001656317, 0.001759402, 0.001757629, 0.001671323, 
    0.001616084, 0.001808665, 0.001565497, 0.00125305, 0.001004395, 
    0.0009918716, 0.0008743986, 0.0006534662, 0.0005727668, 0.0004452399,
  0.001586739, 0.001683358, 0.001738191, 0.001831083, 0.001791379, 
    0.001600683, 0.001474559, 0.001463711, 0.001233546, 0.0009728086, 
    0.0009344465, 0.0009057774, 0.0007408706, 0.0006242748, 0.0005510382,
  0.001820665, 0.001793177, 0.001731958, 0.001686045, 0.001676727, 
    0.001639361, 0.001436773, 0.001014333, 0.0009021251, 0.0009252696, 
    0.0009088656, 0.0008924567, 0.0008347257, 0.0007513419, 0.0005824679,
  0.001868581, 0.001748483, 0.001644042, 0.001577846, 0.001538776, 
    0.001481712, 0.001503974, 0.001298713, 0.001031422, 0.0009400339, 
    0.0008850959, 0.0009160078, 0.0009309995, 0.0009047482, 0.0006672354,
  0.001826811, 0.001756098, 0.001660988, 0.001556777, 0.001482955, 
    0.001392601, 0.001290938, 0.001259773, 0.001290046, 0.001128579, 
    0.0009504523, 0.0008907028, 0.0009150573, 0.0009512226, 0.0008482409,
  0.001555766, 0.001455278, 0.001342344, 0.001222341, 0.001140481, 
    0.001073289, 0.0009678273, 0.0009189001, 0.0009963405, 0.001096747, 
    0.001072254, 0.0009330246, 0.0009029701, 0.0009092559, 0.0008916768,
  0.001230985, 0.001137925, 0.001050741, 0.0009538901, 0.0007975296, 
    0.000678191, 0.0006628201, 0.0006356242, 0.0006328046, 0.0007910933, 
    0.001128029, 0.001018218, 0.0008941265, 0.0008379885, 0.000791706,
  0.001015483, 0.0009309087, 0.0008533891, 0.0006196437, 0.0004752462, 
    0.0004227841, 0.0004245772, 0.0004585165, 0.0004925792, 0.0006832032, 
    0.0009711073, 0.0009782707, 0.0008450185, 0.0007891406, 0.0007794151,
  0.001150681, 0.001341942, 0.001240159, 0.001419108, 0.0014117, 0.001440032, 
    0.001415104, 0.00127047, 0.001008799, 0.0009408019, 0.0009089399, 
    0.0009184623, 0.0008894747, 0.0008656664, 0.0008116303,
  0.001499546, 0.001438049, 0.001419224, 0.001366088, 0.001332549, 
    0.001449706, 0.001522888, 0.001430257, 0.001171878, 0.001087105, 
    0.001055166, 0.001084587, 0.001007182, 0.0007892211, 0.0007543621,
  0.001695996, 0.001653507, 0.001591359, 0.001484925, 0.001290843, 
    0.001196956, 0.001530209, 0.001583139, 0.001454949, 0.001222012, 
    0.001247386, 0.001170377, 0.001028615, 0.0008971345, 0.0007342766,
  0.001668001, 0.001591536, 0.001675123, 0.001729849, 0.001624509, 
    0.001439832, 0.001301631, 0.001623763, 0.001590664, 0.001333484, 
    0.001264901, 0.001209983, 0.001036713, 0.0009083073, 0.0007545594,
  0.001611639, 0.001622773, 0.001646683, 0.001625759, 0.001762557, 
    0.001669168, 0.001596174, 0.001379015, 0.001307685, 0.001283005, 
    0.001295012, 0.001171659, 0.0009765766, 0.0008525467, 0.0007074815,
  0.001399476, 0.001421683, 0.001565447, 0.001646494, 0.001655513, 
    0.001664536, 0.001723068, 0.001685989, 0.001440208, 0.001388846, 
    0.001328265, 0.001200182, 0.0009653148, 0.000782607, 0.0006378187,
  0.001200629, 0.001197516, 0.001255539, 0.001378756, 0.001520584, 0.0015982, 
    0.001594886, 0.001611922, 0.001631897, 0.001480967, 0.001365649, 
    0.001142305, 0.0009006484, 0.0007061965, 0.0005402166,
  0.001033226, 0.0009861306, 0.0009910939, 0.00102877, 0.001051722, 
    0.001147547, 0.001155248, 0.001315465, 0.001344574, 0.001410181, 
    0.001280237, 0.001079084, 0.0008412617, 0.0006467658, 0.0005107562,
  0.0009988053, 0.0009430912, 0.0009157675, 0.0008742134, 0.0007801328, 
    0.0006949915, 0.0006758279, 0.0007053092, 0.0009440535, 0.001156201, 
    0.001190425, 0.001000415, 0.0007296153, 0.0005845652, 0.0004911806,
  0.001060416, 0.0009115685, 0.0007951865, 0.0006109793, 0.0004547451, 
    0.0004073704, 0.0004225858, 0.0004906275, 0.0005496104, 0.0007348044, 
    0.0009404558, 0.0008246137, 0.0006738613, 0.0005778368, 0.0005490076,
  0.001119773, 0.00128926, 0.001030732, 0.001262456, 0.001286535, 
    0.001131106, 0.001039471, 0.0009123924, 0.000877483, 0.0008126728, 
    0.0008937704, 0.001019348, 0.001029456, 0.00101287, 0.0009098376,
  0.001400711, 0.001303919, 0.001099588, 0.001206899, 0.00119159, 
    0.001155154, 0.001066447, 0.0009368692, 0.0008875334, 0.000936691, 
    0.0009815148, 0.0011007, 0.001118415, 0.0008747082, 0.0008054513,
  0.001574736, 0.001702324, 0.001398978, 0.001131198, 0.001115057, 
    0.0008297915, 0.001105841, 0.001016027, 0.0009898745, 0.001010576, 
    0.001094818, 0.001085572, 0.001012951, 0.0009580094, 0.0008269169,
  0.001435889, 0.001594324, 0.001677983, 0.001404153, 0.001230065, 
    0.001073101, 0.0009301979, 0.001075642, 0.001075601, 0.001067232, 
    0.001087592, 0.001060006, 0.0009408618, 0.0008917514, 0.0008690783,
  0.001242705, 0.001452039, 0.001626634, 0.001620628, 0.001431133, 
    0.001342693, 0.001136413, 0.0007777347, 0.0008333444, 0.001024515, 
    0.001086193, 0.001033342, 0.0009361758, 0.0009050407, 0.0008856294,
  0.001108668, 0.001192032, 0.001573083, 0.001618918, 0.001556608, 
    0.001523654, 0.001402457, 0.001218118, 0.001081964, 0.001093328, 
    0.001131675, 0.001069601, 0.000966835, 0.000882122, 0.0008418383,
  0.001019022, 0.001037708, 0.0012392, 0.001538923, 0.001567035, 0.001522479, 
    0.001487682, 0.001467257, 0.001292082, 0.001241763, 0.001187002, 
    0.001065181, 0.0009442242, 0.000880995, 0.0008755149,
  0.001007357, 0.0009726716, 0.0010228, 0.001189188, 0.001390634, 
    0.001456569, 0.001467454, 0.001509698, 0.001375524, 0.001226951, 
    0.001096468, 0.001076898, 0.0009834528, 0.0008982152, 0.0008868988,
  0.001030023, 0.0009459839, 0.0009376146, 0.0009452218, 0.0008595409, 
    0.0009716028, 0.001090004, 0.001211915, 0.001319275, 0.00122786, 
    0.001095039, 0.001102741, 0.001015364, 0.0009195401, 0.0008030375,
  0.000986967, 0.0008421813, 0.0007705322, 0.000612502, 0.0004821771, 
    0.0004673317, 0.0006431363, 0.0009510267, 0.001015336, 0.00103561, 
    0.001118207, 0.00114023, 0.001039776, 0.0009410867, 0.0007534442,
  0.001390358, 0.001501217, 0.001360177, 0.001506426, 0.001402244, 
    0.001268526, 0.001167357, 0.001135221, 0.001144363, 0.0008614194, 
    0.0008554411, 0.0009237347, 0.0007736135, 0.0007445771, 0.0006839352,
  0.00153096, 0.001608503, 0.001523456, 0.001525211, 0.001343394, 
    0.001114401, 0.001039788, 0.001096658, 0.001040366, 0.0009873824, 
    0.0009089131, 0.001029598, 0.001045702, 0.0006964196, 0.0006415643,
  0.00143486, 0.001581999, 0.001617108, 0.001519794, 0.001174232, 
    0.0007870342, 0.0009702298, 0.0009846864, 0.0009632005, 0.0009741849, 
    0.001019013, 0.001018731, 0.00103605, 0.0009902403, 0.0007427314,
  0.001385329, 0.00161932, 0.001600858, 0.00145138, 0.00119254, 0.0009016466, 
    0.000649146, 0.0008575417, 0.0009165077, 0.0009507945, 0.0009826575, 
    0.001002816, 0.0009911139, 0.0009734341, 0.0008818741,
  0.001348334, 0.001595224, 0.001614161, 0.001502928, 0.001326791, 
    0.001036794, 0.0009078312, 0.0006249087, 0.0006813305, 0.0008497216, 
    0.0009429863, 0.001001495, 0.0009790096, 0.0009767106, 0.000912035,
  0.001345119, 0.001570269, 0.001637695, 0.001569414, 0.001460156, 
    0.001303009, 0.001099016, 0.001000907, 0.0009805887, 0.001065807, 
    0.001093274, 0.001053602, 0.0009727369, 0.0008596587, 0.0007715569,
  0.001313738, 0.001499627, 0.001660436, 0.001638668, 0.001528327, 
    0.001462122, 0.001319026, 0.001203848, 0.001134988, 0.001169805, 
    0.00115477, 0.001039399, 0.0009007553, 0.0007504934, 0.0005929264,
  0.001299482, 0.001425258, 0.001570457, 0.001626245, 0.001605097, 
    0.001523312, 0.001401877, 0.001310519, 0.001206591, 0.001168063, 
    0.001036574, 0.0009278462, 0.0007435338, 0.000558676, 0.0004619062,
  0.001256595, 0.001359156, 0.001447721, 0.001400771, 0.001307296, 
    0.00134775, 0.001290299, 0.001230645, 0.001156735, 0.001012138, 
    0.0008621163, 0.0007444351, 0.0005938276, 0.0005261329, 0.0004999809,
  0.001119404, 0.001143706, 0.001122587, 0.0008847295, 0.0008840785, 
    0.001050537, 0.001113143, 0.001064424, 0.0008956454, 0.0008246301, 
    0.0007268554, 0.0006527665, 0.0005986193, 0.0005511029, 0.0005639835,
  0.001537543, 0.001781634, 0.001712083, 0.001485812, 0.001380445, 
    0.001505521, 0.001270214, 0.001034894, 0.000922363, 0.0007998899, 
    0.0008822234, 0.0008983836, 0.0008228428, 0.0007125082, 0.0006141741,
  0.001755777, 0.0016646, 0.001365983, 0.00102194, 0.0009412126, 0.00134763, 
    0.001316636, 0.001069582, 0.0009438088, 0.0008903826, 0.0008855583, 
    0.0009559113, 0.0009431236, 0.000622668, 0.0005298762,
  0.001606998, 0.001516556, 0.001259597, 0.0009446089, 0.0009351025, 
    0.001035538, 0.001247774, 0.001058327, 0.0009822886, 0.0009340504, 
    0.0009317723, 0.0009346124, 0.0008980136, 0.0007940062, 0.0005961107,
  0.001614352, 0.001496084, 0.001342597, 0.001179588, 0.001088682, 
    0.00112906, 0.0008962839, 0.0009748939, 0.0009580398, 0.0009144518, 
    0.0009011399, 0.000871475, 0.0008256586, 0.0008815777, 0.0007721047,
  0.001655116, 0.001531504, 0.001423516, 0.001307878, 0.001208792, 
    0.001106133, 0.001057327, 0.0006940116, 0.0007096997, 0.0007165204, 
    0.000808617, 0.0008057086, 0.0007784809, 0.0008635067, 0.0008621356,
  0.001689485, 0.001577926, 0.001469902, 0.001378843, 0.001342507, 
    0.001275105, 0.00108802, 0.0009859108, 0.0009370252, 0.0009286536, 
    0.0008012537, 0.000785849, 0.000773399, 0.0008149383, 0.0008128066,
  0.001708281, 0.001631232, 0.001525066, 0.001422549, 0.001367313, 
    0.001317637, 0.001252927, 0.001122727, 0.001047528, 0.00103461, 
    0.0009299916, 0.0007679053, 0.000758754, 0.0007558947, 0.0007222137,
  0.001777689, 0.001691832, 0.001573371, 0.001475324, 0.001418723, 
    0.001338933, 0.001277991, 0.001189306, 0.001024618, 0.0008902259, 
    0.000798544, 0.0007448134, 0.0006921132, 0.0006414647, 0.000548194,
  0.001776966, 0.001688705, 0.001588099, 0.001452916, 0.001319234, 
    0.001259846, 0.001198359, 0.001089327, 0.0008890619, 0.0006962285, 
    0.0006380381, 0.0007008233, 0.000600689, 0.0005166248, 0.0004567807,
  0.001476107, 0.001389846, 0.001333849, 0.001143689, 0.00109328, 
    0.001037735, 0.0009991238, 0.0009235775, 0.0007016764, 0.0005786828, 
    0.0005304811, 0.0005711301, 0.0004982231, 0.0004502238, 0.0004489468,
  0.001248508, 0.001219567, 0.001018534, 0.001063043, 0.0009009029, 
    0.0008609207, 0.0009629054, 0.0009775952, 0.000890159, 0.0005626698, 
    0.0005986087, 0.0009018746, 0.0008886118, 0.000869943, 0.001181401,
  0.001276013, 0.001156347, 0.001102016, 0.00103509, 0.0009484941, 
    0.001047879, 0.001070993, 0.0009831832, 0.0007605267, 0.0008688467, 
    0.0008284794, 0.001057971, 0.001026643, 0.0008056707, 0.0008668484,
  0.00144209, 0.001287118, 0.001178664, 0.001148325, 0.001101614, 
    0.0008984886, 0.000923562, 0.0008384815, 0.0008186367, 0.0008825391, 
    0.0009155108, 0.0009571592, 0.001012868, 0.0009609894, 0.0008584068,
  0.001504205, 0.001490825, 0.001438543, 0.001277312, 0.001044591, 
    0.0009328554, 0.0006600128, 0.000641721, 0.0007434404, 0.0008000587, 
    0.0008356635, 0.0008847598, 0.0009559576, 0.0009710098, 0.0009067976,
  0.001416616, 0.001413205, 0.001397824, 0.001341615, 0.001123613, 
    0.0009974929, 0.0009350016, 0.0004632602, 0.0005804804, 0.000729915, 
    0.0007897485, 0.0008372758, 0.0008989378, 0.0009967422, 0.0009386044,
  0.001412176, 0.001350625, 0.001327268, 0.001291696, 0.001238101, 0.0010943, 
    0.0009198358, 0.0008785078, 0.0007590157, 0.0007609452, 0.0007656016, 
    0.0008043321, 0.0009064105, 0.0009068316, 0.0008448118,
  0.001429282, 0.001338733, 0.001255423, 0.001221641, 0.001181421, 
    0.00113667, 0.001090998, 0.0008761383, 0.000806116, 0.0008023941, 
    0.0007466408, 0.0007374029, 0.0007877438, 0.0007925822, 0.0007420597,
  0.001444662, 0.001373963, 0.001288622, 0.001233073, 0.001194222, 
    0.001166324, 0.001109412, 0.0009326158, 0.00074176, 0.0007048444, 
    0.0006513527, 0.0006607374, 0.000645643, 0.0006259012, 0.000553315,
  0.001551493, 0.001456493, 0.001381139, 0.001231877, 0.00110937, 
    0.001038847, 0.0009803852, 0.0008420358, 0.0007138521, 0.0005641287, 
    0.0005079288, 0.0005359222, 0.0005119178, 0.000514988, 0.0005453617,
  0.001470941, 0.001356772, 0.001259541, 0.000975835, 0.0008783055, 
    0.000809159, 0.0007700078, 0.0007634776, 0.0006384858, 0.0004771789, 
    0.0004815481, 0.0005396588, 0.0005536377, 0.0005171645, 0.0005813757,
  0.0009020907, 0.0009367033, 0.0007864323, 0.0007844973, 0.0006257721, 
    0.0006359988, 0.0007526646, 0.0007982185, 0.0008329937, 0.0007845858, 
    0.0008583507, 0.001159275, 0.001146059, 0.00106756, 0.0009847258,
  0.00109148, 0.0009597733, 0.0008664211, 0.0007580524, 0.0006444335, 
    0.0006415929, 0.0007760911, 0.0007434114, 0.0007335758, 0.0008258015, 
    0.0008170918, 0.001074609, 0.001172077, 0.0009512314, 0.0008620259,
  0.001340134, 0.001089289, 0.0009617395, 0.0009064375, 0.0008163765, 
    0.0005018722, 0.0006779765, 0.0007119311, 0.0007446186, 0.0007236237, 
    0.0007885942, 0.0009177874, 0.001059646, 0.00109889, 0.0009738854,
  0.00129569, 0.001317026, 0.001237516, 0.001036373, 0.0008842243, 
    0.0008061365, 0.0004367381, 0.0004653325, 0.0005744679, 0.0006223764, 
    0.0006268548, 0.0008216393, 0.0008825937, 0.001001969, 0.0009947278,
  0.001213163, 0.001167675, 0.001162717, 0.001112162, 0.0009054122, 
    0.0008411473, 0.0008291461, 0.00049883, 0.0005684985, 0.0005813292, 
    0.000589602, 0.0006780695, 0.0007446253, 0.0009460734, 0.001022927,
  0.001216124, 0.001149347, 0.001080457, 0.001058564, 0.001011955, 
    0.000916763, 0.0007905338, 0.0007755546, 0.0007527891, 0.000700965, 
    0.0005732503, 0.0007366954, 0.0007586654, 0.0008949809, 0.0009322634,
  0.001322972, 0.001211502, 0.001095704, 0.001048618, 0.0009985243, 
    0.0009940432, 0.0009231191, 0.0007608363, 0.0007237767, 0.0006627347, 
    0.0005685399, 0.0007130982, 0.0008224678, 0.0009211147, 0.0008739953,
  0.001396201, 0.001290898, 0.001179021, 0.001156181, 0.001077399, 
    0.0009749516, 0.0009191326, 0.000785764, 0.0005980327, 0.0005093881, 
    0.0004861858, 0.0006567746, 0.0008561123, 0.000889616, 0.0007377327,
  0.001565599, 0.001426304, 0.001222224, 0.001077731, 0.001023428, 
    0.0009181585, 0.0008217912, 0.0006855927, 0.0005345994, 0.0004657251, 
    0.0004266863, 0.0004812531, 0.0006968397, 0.0007659394, 0.0006879277,
  0.001462692, 0.001322732, 0.001260882, 0.0008872684, 0.0008260815, 
    0.000692594, 0.0006969623, 0.0006902147, 0.0004732784, 0.0004029291, 
    0.0003456725, 0.0004263966, 0.0004722591, 0.0006204438, 0.0006346827,
  0.0007959139, 0.0008278707, 0.0007499365, 0.0008087077, 0.0007697158, 
    0.0007045017, 0.0007251283, 0.000719674, 0.0007588518, 0.0008469204, 
    0.0009707537, 0.001006758, 0.0007920092, 0.0007294178, 0.0008298266,
  0.001019865, 0.0009008486, 0.000867166, 0.0008536577, 0.0008304002, 
    0.0006156023, 0.0007322711, 0.0006980602, 0.0007650138, 0.0008728279, 
    0.00105334, 0.001124637, 0.0009396084, 0.000678622, 0.000672542,
  0.001108987, 0.001020433, 0.0009670351, 0.0009344861, 0.0008749817, 
    0.0005959937, 0.0007353437, 0.0006735315, 0.0007271938, 0.0008895612, 
    0.00110218, 0.001166774, 0.0009660999, 0.0008522857, 0.0007606078,
  0.001156829, 0.001033769, 0.0009930191, 0.0009436014, 0.0009389207, 
    0.0009092838, 0.0006815242, 0.0005678691, 0.0006552087, 0.0008530015, 
    0.001020845, 0.001088827, 0.0009468314, 0.0008677288, 0.0008657616,
  0.001294718, 0.001139726, 0.001068497, 0.0009931142, 0.0009351152, 
    0.0009662934, 0.0008807979, 0.0005339693, 0.0005495992, 0.0007475789, 
    0.0008886897, 0.0009350759, 0.0009002652, 0.0008902009, 0.0009098123,
  0.001664636, 0.001521832, 0.001350242, 0.001151961, 0.001043172, 
    0.001023424, 0.0008728153, 0.0007534691, 0.0006560004, 0.0007309137, 
    0.0007879969, 0.0008476507, 0.0008297626, 0.0008299477, 0.0008649663,
  0.00196688, 0.001875558, 0.001750451, 0.001579372, 0.001333742, 
    0.001054357, 0.001026757, 0.0008147209, 0.0006909305, 0.0006675959, 
    0.0007507769, 0.0007929906, 0.0007659638, 0.0007652989, 0.0007820574,
  0.002033851, 0.001903482, 0.00180613, 0.001597762, 0.00146523, 0.001169314, 
    0.001019777, 0.0008430178, 0.0005880365, 0.0005881807, 0.0006179316, 
    0.0007356987, 0.0007373016, 0.0007039838, 0.0006787834,
  0.002176214, 0.001990064, 0.001797579, 0.001517567, 0.001388821, 
    0.001248256, 0.000981768, 0.0006948082, 0.0005318859, 0.0005070095, 
    0.0004886934, 0.0005432263, 0.0006858638, 0.0006642923, 0.0007055941,
  0.002452204, 0.00215318, 0.001909796, 0.001540056, 0.00119771, 0.001021066, 
    0.0008995443, 0.00074064, 0.0004908129, 0.0004451608, 0.0003590433, 
    0.0004321272, 0.0004754027, 0.0005832507, 0.0006880375,
  0.0007588147, 0.0008599744, 0.0009153812, 0.0009825152, 0.0009743248, 
    0.0009341948, 0.0009665536, 0.0009263335, 0.0008902802, 0.0007467238, 
    0.0006180495, 0.0005993113, 0.0006273686, 0.0007752799, 0.0008247537,
  0.001170023, 0.001038611, 0.001030799, 0.001027169, 0.00102939, 
    0.000887874, 0.001020923, 0.0009510684, 0.0008668701, 0.0008306029, 
    0.0007226936, 0.0007580962, 0.0008195339, 0.0007403792, 0.0007499843,
  0.001599644, 0.00144435, 0.001420125, 0.001312734, 0.001314663, 
    0.001056704, 0.001152501, 0.0009158971, 0.0008385842, 0.0008452622, 
    0.0008039051, 0.0007802176, 0.0008150977, 0.0009494136, 0.0008775015,
  0.001605705, 0.001514139, 0.001452599, 0.001495652, 0.001630029, 
    0.001534781, 0.0007992656, 0.0007691326, 0.0008008351, 0.0008991141, 
    0.0008718648, 0.0008259561, 0.0007970626, 0.0009156633, 0.0009302878,
  0.001620389, 0.001496979, 0.001543731, 0.001669464, 0.001611421, 
    0.001165749, 0.0008206983, 0.0005320663, 0.000567553, 0.0008700428, 
    0.0008676708, 0.0007851627, 0.0007907608, 0.0009279551, 0.0009589278,
  0.001721564, 0.001602951, 0.001730446, 0.001757091, 0.001518904, 
    0.001055573, 0.0008334413, 0.0007648517, 0.0007979857, 0.0009213449, 
    0.0008018901, 0.0007448637, 0.0007786644, 0.0009485499, 0.0009361622,
  0.001856573, 0.001722543, 0.001802282, 0.001718343, 0.001468105, 
    0.001143911, 0.001009479, 0.0008754724, 0.0008864444, 0.0008598427, 
    0.0007790743, 0.0007230468, 0.0007791852, 0.0008982635, 0.0008860402,
  0.001927777, 0.001804153, 0.001836304, 0.001640692, 0.001406946, 
    0.001191608, 0.001056149, 0.0008846395, 0.0008137409, 0.0007560281, 
    0.0006822525, 0.0006692402, 0.0008116559, 0.0008379252, 0.0007384133,
  0.002011182, 0.001963532, 0.001854514, 0.001500266, 0.001122338, 
    0.0009425132, 0.0008255097, 0.0007279345, 0.0007024345, 0.0006578375, 
    0.000632196, 0.0006742512, 0.0007358841, 0.0007321155, 0.0006290278,
  0.002094554, 0.001970285, 0.001629522, 0.001011808, 0.0008029936, 
    0.0006903734, 0.0006445073, 0.0006284373, 0.0005459277, 0.0004922534, 
    0.0004782732, 0.000578059, 0.0006080359, 0.0005631063, 0.0005513872,
  0.0009770471, 0.0009416079, 0.0008803158, 0.0008095417, 0.000739452, 
    0.0007092837, 0.0007609021, 0.000721974, 0.0007295062, 0.0006894237, 
    0.0006736764, 0.0007354516, 0.0007318081, 0.0007144432, 0.0005979612,
  0.001136523, 0.00101087, 0.0009412069, 0.0008759109, 0.0007772172, 
    0.0007860491, 0.0008659492, 0.0008541182, 0.0008565372, 0.0009195675, 
    0.0008583619, 0.0008947222, 0.0009647377, 0.0006853217, 0.0005105183,
  0.00118615, 0.001045692, 0.0009819301, 0.0009352486, 0.000884773, 
    0.0007318124, 0.0009078397, 0.0009769684, 0.000992212, 0.001070524, 
    0.0009901325, 0.0008903714, 0.0009599624, 0.0009724534, 0.0006924202,
  0.001385666, 0.001342375, 0.001370026, 0.001324651, 0.001169282, 
    0.00113187, 0.0008429622, 0.0009306949, 0.001017711, 0.0009232527, 
    0.000813438, 0.0007213739, 0.0008798402, 0.0008302261, 0.0007167552,
  0.001475243, 0.001537002, 0.00149413, 0.001506527, 0.001168921, 
    0.001035124, 0.001163141, 0.0006825135, 0.0006036005, 0.0005564322, 
    0.0005758435, 0.0007593962, 0.0008461857, 0.0007757562, 0.0007063359,
  0.001467673, 0.001398994, 0.001333002, 0.001335834, 0.001240121, 
    0.001065572, 0.001089792, 0.0009486999, 0.0007982657, 0.0007901291, 
    0.0006633208, 0.0008233491, 0.0008097116, 0.0007510225, 0.0006585752,
  0.001473303, 0.001383792, 0.00132886, 0.001245368, 0.001186118, 
    0.001155298, 0.001090661, 0.000899142, 0.0008577092, 0.0008090224, 
    0.0007438433, 0.0006966428, 0.0006425941, 0.0005498342, 0.0005320327,
  0.001507652, 0.001442932, 0.001344395, 0.001267771, 0.001236169, 
    0.001204753, 0.001155397, 0.0009043369, 0.0007821356, 0.0006885321, 
    0.0006566272, 0.0006163934, 0.0005521618, 0.0004797131, 0.0004415567,
  0.001559165, 0.001501144, 0.001412512, 0.00125007, 0.001127878, 
    0.001052068, 0.0009325749, 0.0007929422, 0.0007068668, 0.000636872, 
    0.0006294586, 0.000614602, 0.0005650042, 0.0005200089, 0.0005318986,
  0.001531289, 0.001420555, 0.001222484, 0.0008489952, 0.0008306061, 
    0.0007823551, 0.0007337054, 0.0007172926, 0.0006539724, 0.0005890488, 
    0.0005795005, 0.0005953415, 0.0005903534, 0.0005207544, 0.0005596928,
  0.001082741, 0.001017632, 0.0009538549, 0.0009537684, 0.0008034174, 
    0.0006818417, 0.0007428267, 0.0006363709, 0.0005430976, 0.0003142463, 
    0.0003337042, 0.0003908947, 0.0003298467, 0.0003509618, 0.0003466005,
  0.001202655, 0.001102809, 0.001045433, 0.0009925644, 0.0008266486, 
    0.0007759575, 0.0007854326, 0.0006679785, 0.0006047484, 0.0005253815, 
    0.0004834991, 0.0005788236, 0.0006175407, 0.0004823738, 0.0004438057,
  0.001216008, 0.001036034, 0.001030205, 0.001039163, 0.0008889139, 
    0.0006899404, 0.0007766615, 0.0006904908, 0.0006022807, 0.0006372326, 
    0.0006664629, 0.0007261792, 0.0008174467, 0.0008677837, 0.0008499991,
  0.001083204, 0.001102029, 0.001199441, 0.00114102, 0.0009237305, 
    0.0008895134, 0.0006205906, 0.0006062184, 0.0006039311, 0.0006448353, 
    0.0007716069, 0.0008264898, 0.0009062712, 0.0009435913, 0.0009452845,
  0.001217311, 0.001163461, 0.001208748, 0.001251096, 0.0009820515, 
    0.0009455259, 0.0009622163, 0.0004876812, 0.0004338718, 0.0004734774, 
    0.0005156694, 0.0006989641, 0.0007567276, 0.0007440575, 0.0007652062,
  0.001372469, 0.001285243, 0.001259756, 0.001236421, 0.00117867, 
    0.001096402, 0.001019776, 0.001017253, 0.0008550216, 0.0007577292, 
    0.0005133243, 0.0005870583, 0.0005561797, 0.0005747034, 0.0006091971,
  0.001430465, 0.001364741, 0.00130962, 0.001244702, 0.001230041, 
    0.001237276, 0.001074743, 0.0009016237, 0.0007429132, 0.0005895031, 
    0.0005095061, 0.0004888137, 0.0004641767, 0.0004436454, 0.0004900029,
  0.001485167, 0.001427555, 0.001321736, 0.001311987, 0.001305645, 
    0.001270823, 0.001139719, 0.0007706865, 0.0005877159, 0.0004792941, 
    0.0004248209, 0.0004068023, 0.000400431, 0.0003930209, 0.0004096263,
  0.001538244, 0.001476913, 0.001448564, 0.001351246, 0.001216254, 
    0.001083665, 0.0008600367, 0.0006064564, 0.0005310505, 0.0004150589, 
    0.0003634578, 0.0003655943, 0.0003752216, 0.000410642, 0.0004092008,
  0.001618857, 0.00152617, 0.001345477, 0.0009557265, 0.0008689412, 
    0.0007321787, 0.0006708898, 0.0006108917, 0.0004751649, 0.0003268232, 
    0.000276361, 0.0003574005, 0.0003873791, 0.0004015279, 0.000415713,
  0.001108572, 0.001206161, 0.001151764, 0.001157695, 0.0009627831, 
    0.0008086499, 0.0008404998, 0.0006808156, 0.0005009954, 0.0003054441, 
    0.0003081355, 0.0003638522, 0.0002774343, 0.0002964442, 0.0002500317,
  0.001297451, 0.001216393, 0.001129071, 0.001103696, 0.0008106588, 
    0.0007984095, 0.0008067867, 0.0006142588, 0.0004882666, 0.0004169063, 
    0.0003683562, 0.0004880503, 0.0005215287, 0.0003720983, 0.0003482983,
  0.001613224, 0.001217965, 0.001026756, 0.0009905687, 0.0008506567, 
    0.0006382747, 0.0006728002, 0.0005373836, 0.0004592803, 0.0005136082, 
    0.0005481804, 0.0005794271, 0.0006374783, 0.000700767, 0.0006847883,
  0.001431559, 0.001287804, 0.001203846, 0.001102875, 0.0009409455, 
    0.0008602662, 0.0004501653, 0.0004555745, 0.0004254622, 0.0004744226, 
    0.000572951, 0.0006224292, 0.0006997235, 0.0007443849, 0.000736053,
  0.001365144, 0.001304393, 0.001286544, 0.001333799, 0.0009981568, 
    0.0009641431, 0.0009071147, 0.000413028, 0.0003268056, 0.0004445652, 
    0.0004723718, 0.000568315, 0.0006556978, 0.0006492913, 0.0006090511,
  0.001405829, 0.00137713, 0.001343892, 0.001337221, 0.001248411, 
    0.001100484, 0.0009327309, 0.0009318975, 0.0007495832, 0.000670723, 
    0.0003862058, 0.0005370085, 0.0005335225, 0.0005069676, 0.0005487896,
  0.00146952, 0.001431105, 0.001392801, 0.001332032, 0.001327052, 
    0.001267995, 0.001073542, 0.0009684042, 0.0006927985, 0.0005534294, 
    0.0004600151, 0.0004290574, 0.0004322092, 0.0004279163, 0.0004862879,
  0.001475846, 0.001400495, 0.001321806, 0.001278269, 0.001253751, 
    0.001235431, 0.001154643, 0.0008657611, 0.000561304, 0.0004563914, 
    0.0003993834, 0.0003911187, 0.0004075095, 0.0004322006, 0.0004858337,
  0.001494146, 0.00140213, 0.001327673, 0.001260075, 0.001178488, 
    0.001118155, 0.0009783359, 0.0006411453, 0.0004826605, 0.0003936906, 
    0.0003588674, 0.0003631783, 0.0003953537, 0.0004523667, 0.0004620464,
  0.001583705, 0.001524605, 0.001449187, 0.001179557, 0.00100865, 
    0.000818508, 0.0007614465, 0.000615009, 0.0004282775, 0.0002851952, 
    0.0002356774, 0.0003297899, 0.0003728092, 0.0003935049, 0.0004010651,
  0.0009781726, 0.0009871953, 0.0009741007, 0.0009885472, 0.0009328161, 
    0.0007728367, 0.0009857015, 0.0008271234, 0.0006940152, 0.0005813903, 
    0.0005122109, 0.0004757582, 0.0003551274, 0.0003149803, 0.0002367092,
  0.0011337, 0.001013778, 0.001084197, 0.001071126, 0.0007018996, 
    0.0007146806, 0.0007421414, 0.0006985838, 0.0006449798, 0.0006134629, 
    0.0005107575, 0.0005144039, 0.0004538537, 0.0002643706, 0.0002744727,
  0.001574817, 0.001272418, 0.001107973, 0.001038138, 0.0007760378, 
    0.0005157415, 0.0006120368, 0.0006092804, 0.0006051542, 0.0005924946, 
    0.0005404379, 0.0004972406, 0.0005236655, 0.000535211, 0.000543373,
  0.001320522, 0.001230282, 0.001185554, 0.0009885393, 0.0008099469, 
    0.0007366975, 0.0004061735, 0.0004657768, 0.0004685052, 0.0004304144, 
    0.0005213706, 0.0005473381, 0.0006112816, 0.0006176644, 0.0006248661,
  0.001371433, 0.001281428, 0.001283129, 0.001184952, 0.0008470022, 
    0.0008374313, 0.0008009743, 0.0003667693, 0.0002913841, 0.0003327101, 
    0.0003958281, 0.0005005851, 0.0005950238, 0.000593011, 0.0006290062,
  0.001389331, 0.001346341, 0.001324628, 0.001237403, 0.001074142, 
    0.000891683, 0.0008244085, 0.0008369664, 0.0007058925, 0.000535327, 
    0.0004000901, 0.0004806364, 0.0005379428, 0.0005779134, 0.0006177929,
  0.001356518, 0.001335276, 0.001289749, 0.001227701, 0.001208313, 
    0.001154217, 0.0009425708, 0.0007866902, 0.0006129178, 0.0005375383, 
    0.0004760008, 0.0004401173, 0.0004371923, 0.0004732376, 0.0005696358,
  0.001366192, 0.0013105, 0.001249379, 0.001184404, 0.001161985, 0.001163382, 
    0.001116904, 0.000689049, 0.0005126707, 0.0004457936, 0.0003918787, 
    0.000389392, 0.0003902134, 0.000439586, 0.0004879393,
  0.001468599, 0.001372139, 0.001275579, 0.001205577, 0.001183776, 
    0.001119274, 0.0009031068, 0.0005565797, 0.0004714675, 0.0003975846, 
    0.0003735356, 0.0003882587, 0.0004198042, 0.0004462633, 0.0004313198,
  0.00161566, 0.001517367, 0.001462267, 0.00134992, 0.001041695, 
    0.0008801417, 0.0007012562, 0.0005022381, 0.0004112757, 0.0003038025, 
    0.0003022074, 0.0003789594, 0.000395592, 0.000389771, 0.0004037582,
  0.001006736, 0.0009823011, 0.0008874878, 0.0007315426, 0.0006184022, 
    0.0005356625, 0.0006942084, 0.0007402005, 0.0007676345, 0.0005720399, 
    0.0004743141, 0.0005136624, 0.0004298514, 0.0003250871, 0.0002397101,
  0.001084617, 0.0009902683, 0.000792174, 0.0006713173, 0.0005153423, 
    0.0004821184, 0.0005546432, 0.0005939304, 0.0006490304, 0.0006551039, 
    0.000511672, 0.0005348908, 0.0005101548, 0.0002350139, 0.0001595515,
  0.001346509, 0.001011347, 0.0008044319, 0.0007302599, 0.0006105584, 
    0.0003623689, 0.0004475604, 0.0004969691, 0.0005599964, 0.0006301169, 
    0.0006274083, 0.0006034864, 0.0006189318, 0.0005587117, 0.000395723,
  0.001409433, 0.001261334, 0.001114473, 0.0008423994, 0.0007391425, 
    0.0007316986, 0.0002917075, 0.0003919668, 0.0004616416, 0.0005081396, 
    0.0006030259, 0.0006131324, 0.0006191154, 0.0005881498, 0.0005118567,
  0.001428873, 0.001249513, 0.001200358, 0.001065016, 0.0008064589, 
    0.000821251, 0.000804072, 0.0003258072, 0.0003164207, 0.0004214085, 
    0.0004891125, 0.0005445878, 0.0005570347, 0.0005311203, 0.0004789382,
  0.001461449, 0.001303449, 0.001175147, 0.00109004, 0.0009566693, 
    0.000853584, 0.0007723112, 0.0007406707, 0.00052466, 0.0004963193, 
    0.000429213, 0.0004876847, 0.0005102656, 0.0005055268, 0.0004747191,
  0.001488205, 0.001360382, 0.001208093, 0.001093737, 0.001074931, 
    0.001093902, 0.0007228786, 0.0005476631, 0.0004962853, 0.0004538521, 
    0.0004214401, 0.000414136, 0.0004379236, 0.0004425447, 0.0004849657,
  0.001488189, 0.001316328, 0.001189709, 0.001154589, 0.001176598, 
    0.00114725, 0.0009248391, 0.0005429522, 0.0004543608, 0.0004062059, 
    0.0003761995, 0.0003745249, 0.000388433, 0.0004217351, 0.0004576464,
  0.00149041, 0.001349246, 0.001286127, 0.001242493, 0.001162141, 
    0.0009549573, 0.0006337868, 0.000492281, 0.000416848, 0.0003772881, 
    0.0003509984, 0.0003622883, 0.0003787088, 0.0003953232, 0.0003987014,
  0.001554734, 0.001479088, 0.001403205, 0.0009271907, 0.0006806531, 
    0.00057799, 0.0005329731, 0.0004764055, 0.000387404, 0.0003026479, 
    0.0002889397, 0.0003605629, 0.0003604764, 0.0003598072, 0.0003797565,
  0.000815442, 0.0008080525, 0.0006601411, 0.000636693, 0.0005149605, 
    0.0004168105, 0.0005043528, 0.0005206161, 0.0006009801, 0.0004032758, 
    0.0003365766, 0.0004151254, 0.0003796435, 0.0002847764, 0.0002212644,
  0.0008552846, 0.0007416122, 0.000664587, 0.0005755597, 0.0004232028, 
    0.0003113548, 0.0003888155, 0.0004232192, 0.000487779, 0.0005130972, 
    0.0003851796, 0.0004726382, 0.0004767054, 0.0002448696, 0.0001634662,
  0.001111611, 0.0008411235, 0.0007828386, 0.000714715, 0.0006317958, 
    0.0002609754, 0.0003100012, 0.0003747315, 0.0004006842, 0.0004363623, 
    0.0004620081, 0.0004645016, 0.0004491427, 0.0004111839, 0.0002606832,
  0.001243675, 0.001139069, 0.001008268, 0.0008580562, 0.0008009616, 
    0.0008128871, 0.0002245405, 0.0003228473, 0.0003934147, 0.0003885679, 
    0.0004234854, 0.0004482013, 0.0004376528, 0.0003917114, 0.0002969306,
  0.001276826, 0.00107942, 0.001048217, 0.001051699, 0.0008740925, 
    0.0008180593, 0.0008010201, 0.0002483797, 0.0002801519, 0.0003567876, 
    0.0003935566, 0.0004182245, 0.0004451402, 0.0004251336, 0.0003956697,
  0.001334028, 0.001146922, 0.001086416, 0.001056286, 0.0009366604, 
    0.0007247217, 0.0006704648, 0.0006089559, 0.0004677011, 0.0004440974, 
    0.0003781649, 0.0004056222, 0.0004416755, 0.0004432807, 0.0004351067,
  0.00142139, 0.001198665, 0.001119733, 0.001088442, 0.00108936, 
    0.0009682815, 0.0006481112, 0.0005300141, 0.0004742463, 0.000441247, 
    0.0004113343, 0.0003885933, 0.0003852471, 0.0003939106, 0.0004372668,
  0.001459663, 0.001232189, 0.001173544, 0.00114831, 0.001126496, 
    0.001050126, 0.0008333417, 0.0005256619, 0.0004536333, 0.0004058556, 
    0.0003658168, 0.0003590616, 0.0003500679, 0.0003790727, 0.0004372428,
  0.001448672, 0.001326327, 0.001302855, 0.001226004, 0.001102891, 
    0.0008888337, 0.0006121858, 0.0005023406, 0.0004277102, 0.0003614656, 
    0.0003190647, 0.0003191986, 0.0003351055, 0.0003597747, 0.0003562193,
  0.001556367, 0.001537045, 0.001357904, 0.0007817216, 0.0005891986, 
    0.00054078, 0.000529752, 0.0004976285, 0.0003941773, 0.0002695176, 
    0.0002157287, 0.0002925751, 0.0002863934, 0.0002967532, 0.0003225438,
  0.0007792658, 0.0007978053, 0.0007073295, 0.0007094082, 0.000636753, 
    0.0005756925, 0.0005650753, 0.0005490176, 0.0005503531, 0.0003770168, 
    0.0003126809, 0.0003245716, 0.0002564679, 0.0002492509, 0.0001738773,
  0.0008090225, 0.0007351886, 0.0006696404, 0.0005967765, 0.0005022148, 
    0.0003653282, 0.000454962, 0.0004856481, 0.0005110267, 0.00046742, 
    0.0003157099, 0.0003949489, 0.0004236759, 0.0002442692, 0.0001749141,
  0.001073201, 0.0007696434, 0.0006821746, 0.0006013443, 0.0005177924, 
    0.0002720373, 0.0003255642, 0.0004010783, 0.0004283263, 0.0004460037, 
    0.0004023466, 0.0003995444, 0.0004349974, 0.0004628592, 0.0003387882,
  0.001197906, 0.001149292, 0.0009933759, 0.0007340589, 0.0006279324, 
    0.0006192905, 0.0002411612, 0.0003176743, 0.0003689053, 0.0003628729, 
    0.0003843466, 0.0004166499, 0.0004505158, 0.000436639, 0.0003410149,
  0.001170214, 0.001143075, 0.001138757, 0.0009882255, 0.0008004906, 
    0.0006707669, 0.000696309, 0.0002390708, 0.0001933152, 0.0002623137, 
    0.0003519757, 0.000413559, 0.0004425879, 0.0004078885, 0.0003754014,
  0.001182909, 0.001156283, 0.001119742, 0.001041204, 0.0008563318, 
    0.0007277254, 0.0006864177, 0.0007128517, 0.0005415883, 0.0004026037, 
    0.0003115328, 0.0003784746, 0.0004505824, 0.000457018, 0.0004158358,
  0.001260074, 0.001243743, 0.001153838, 0.001070734, 0.001044183, 
    0.0009278925, 0.0006774574, 0.0005910512, 0.000476715, 0.0004087875, 
    0.0003561393, 0.0003338977, 0.0003360062, 0.0003666945, 0.0004005918,
  0.001356293, 0.001291406, 0.001218307, 0.00112661, 0.001078342, 
    0.001038931, 0.0008073382, 0.0005442577, 0.0004388015, 0.0003415903, 
    0.0002945777, 0.0002942128, 0.0002814742, 0.0003114296, 0.0003682152,
  0.001354429, 0.001332435, 0.001322847, 0.00115425, 0.001069125, 
    0.0009779597, 0.0007031334, 0.0005195667, 0.0004197154, 0.0003004325, 
    0.0002761423, 0.0002737108, 0.0002754579, 0.0003154317, 0.0003794183,
  0.001580715, 0.001527839, 0.001355515, 0.0009719137, 0.0008251839, 
    0.0007299088, 0.0006067126, 0.0005202705, 0.0003737676, 0.0002331646, 
    0.0002078555, 0.000273221, 0.0002860063, 0.0003247862, 0.0003819149,
  0.0008180825, 0.0008213343, 0.0007751962, 0.0007903856, 0.0008291377, 
    0.0008151812, 0.0008514627, 0.0008601123, 0.0008762326, 0.0007276786, 
    0.0006566011, 0.0006460142, 0.0005502373, 0.0004983796, 0.0003677678,
  0.0009366769, 0.0008485586, 0.0008162688, 0.000793685, 0.0006996822, 
    0.0005886605, 0.0006674854, 0.0006924053, 0.0007161078, 0.0006950386, 
    0.0005686797, 0.0005924291, 0.0005461558, 0.0003245826, 0.0002489909,
  0.001164395, 0.0009264625, 0.0008505213, 0.000808205, 0.0006749147, 
    0.000406754, 0.0004565342, 0.0005121627, 0.0005425741, 0.0005671016, 
    0.0005365878, 0.0005070189, 0.0005008792, 0.0004533154, 0.0003218246,
  0.001198572, 0.00119472, 0.001064908, 0.0008273622, 0.0007266935, 
    0.000631541, 0.0003330561, 0.0003784074, 0.000395071, 0.0004136067, 
    0.0004671064, 0.0004721211, 0.0004826011, 0.0004665899, 0.0003946336,
  0.001200792, 0.001163553, 0.001136943, 0.0009499963, 0.000733779, 
    0.0006506806, 0.0006730625, 0.0002666424, 0.000220073, 0.000285416, 
    0.0003601979, 0.0004320757, 0.0004626038, 0.0004566531, 0.0004713353,
  0.001251942, 0.001156304, 0.001119548, 0.0009943915, 0.0008264941, 
    0.0007298416, 0.0006671858, 0.0006951952, 0.0005121151, 0.0003590183, 
    0.0002814598, 0.0003342451, 0.0003926606, 0.0004175387, 0.0004162028,
  0.001462818, 0.001269485, 0.001137362, 0.001028404, 0.0009576251, 
    0.0008611985, 0.0006506376, 0.0005510626, 0.0003953394, 0.0003511984, 
    0.0003249434, 0.0003123973, 0.0003218288, 0.0003276466, 0.0003687723,
  0.001876618, 0.001662223, 0.001450573, 0.001295374, 0.001043134, 
    0.0008977501, 0.0007296606, 0.0005402687, 0.0004402356, 0.0003847159, 
    0.0003290576, 0.0003028122, 0.0002724215, 0.0002769205, 0.0003626503,
  0.001949548, 0.001811755, 0.001703357, 0.001527064, 0.001233842, 
    0.0009458121, 0.0007186661, 0.0005766231, 0.0005220349, 0.0004635092, 
    0.0004247548, 0.0003900007, 0.0003554054, 0.000360786, 0.0003669768,
  0.001860698, 0.001750619, 0.001734375, 0.00140869, 0.0009594513, 
    0.0007563318, 0.0006289817, 0.0006048528, 0.0005704242, 0.000492131, 
    0.0005070035, 0.0005196314, 0.0004695216, 0.0004468874, 0.000422948,
  0.001022461, 0.001055812, 0.001008657, 0.0009472386, 0.0009328287, 
    0.0009613413, 0.001277146, 0.001404269, 0.001498591, 0.001368197, 
    0.001435451, 0.001616472, 0.001395327, 0.001219752, 0.0009888337,
  0.00110504, 0.001113675, 0.001073979, 0.00106408, 0.0008817837, 
    0.0007114915, 0.0008472382, 0.001154588, 0.001338743, 0.001418217, 
    0.00128914, 0.001455789, 0.001329706, 0.0009081534, 0.0007349025,
  0.001239235, 0.001174762, 0.00109946, 0.001085667, 0.0009388826, 
    0.0006094952, 0.0006124187, 0.0006991014, 0.0009170517, 0.001129563, 
    0.001199781, 0.00121155, 0.001157614, 0.001004344, 0.0007138519,
  0.001340996, 0.001311515, 0.001238323, 0.001050586, 0.000969241, 
    0.0008893372, 0.000495255, 0.000505869, 0.000508078, 0.000659899, 
    0.0008349406, 0.0008639639, 0.0008434071, 0.0007500855, 0.0006112217,
  0.001438931, 0.001341152, 0.001333925, 0.001261031, 0.0009565796, 
    0.0009311294, 0.0008971266, 0.0003418934, 0.0003007912, 0.0004172217, 
    0.0005303318, 0.0006390263, 0.0006798876, 0.0006322861, 0.0005788276,
  0.001635883, 0.0014833, 0.001381793, 0.001331848, 0.0009982716, 
    0.0009118152, 0.0008388027, 0.0007318854, 0.0005020377, 0.0004169452, 
    0.0003578543, 0.0004500708, 0.0005413783, 0.0005662742, 0.000534322,
  0.002009894, 0.001796728, 0.001517194, 0.001418977, 0.001260445, 
    0.001173802, 0.0008831957, 0.0006882718, 0.0005175858, 0.0004247949, 
    0.0003669481, 0.0003767691, 0.0003857167, 0.0004313163, 0.0004788921,
  0.002176474, 0.002055305, 0.001847862, 0.001553003, 0.00139848, 
    0.001310176, 0.00112329, 0.0008826027, 0.0007945755, 0.0005625237, 
    0.0004105573, 0.0003504374, 0.0003051471, 0.0003191053, 0.0004446536,
  0.00207685, 0.002019979, 0.001951881, 0.001626408, 0.001410067, 
    0.001189279, 0.0009790377, 0.0008279905, 0.0007807678, 0.0007368695, 
    0.0006128406, 0.0004476574, 0.000359972, 0.0003541067, 0.0003755324,
  0.001977966, 0.001852736, 0.001539825, 0.001182421, 0.001088137, 
    0.0009953824, 0.0009157652, 0.0007543843, 0.0006202045, 0.000533309, 
    0.0006683358, 0.0006616216, 0.000493212, 0.0004190254, 0.0004032513,
  0.001286084, 0.001614162, 0.001300476, 0.00119115, 0.001125455, 
    0.0008979059, 0.001075814, 0.001410669, 0.001510187, 0.001208218, 
    0.001257478, 0.001696936, 0.001385937, 0.001433805, 0.001144207,
  0.001436912, 0.001627913, 0.001444422, 0.001276987, 0.001117425, 
    0.0007853275, 0.0007973178, 0.001104362, 0.001594331, 0.001658259, 
    0.001425001, 0.00183953, 0.001721996, 0.001353106, 0.001095958,
  0.001789608, 0.001824406, 0.001632646, 0.001323527, 0.001188561, 
    0.0007457069, 0.0006830815, 0.0007222001, 0.0008871002, 0.001260499, 
    0.001613675, 0.001698183, 0.001726988, 0.001609374, 0.001218934,
  0.001780994, 0.001895779, 0.00203895, 0.00147329, 0.001272692, 0.001211383, 
    0.0005274396, 0.0005904481, 0.0006052454, 0.0006579369, 0.0009841735, 
    0.001285238, 0.001435885, 0.001409409, 0.001257179,
  0.001896313, 0.002024675, 0.002011105, 0.001940933, 0.001361128, 
    0.001324634, 0.001081175, 0.0003504598, 0.0003711884, 0.0004753399, 
    0.0005453885, 0.0008332562, 0.001000856, 0.001145516, 0.001189137,
  0.002045468, 0.002070188, 0.001978762, 0.001857229, 0.001647211, 
    0.001427625, 0.001109903, 0.0008346786, 0.0005664157, 0.0004654386, 
    0.0003862766, 0.0004899714, 0.0006719359, 0.0008301081, 0.0009206258,
  0.002051182, 0.002023276, 0.001942984, 0.001740955, 0.001499936, 
    0.001483921, 0.001127254, 0.0008872725, 0.0007053936, 0.0005298725, 
    0.0004319856, 0.0003685596, 0.0004056394, 0.0005284895, 0.0006829827,
  0.001903577, 0.002036653, 0.001995364, 0.001567888, 0.001498111, 
    0.001394181, 0.001038688, 0.0007584877, 0.0007179833, 0.00063156, 
    0.0005291625, 0.0003450981, 0.0003067057, 0.0003530065, 0.0004634905,
  0.0018204, 0.001920704, 0.001912998, 0.00167236, 0.001365858, 0.001036216, 
    0.0007739161, 0.0006583245, 0.0005352875, 0.0004803124, 0.0004638143, 
    0.0004256152, 0.0003602535, 0.0003309302, 0.0003372074,
  0.001750177, 0.001819137, 0.001766281, 0.00133048, 0.001010331, 
    0.0007093762, 0.0006283787, 0.0006157032, 0.0004578153, 0.0003560875, 
    0.0004798109, 0.000459754, 0.000366375, 0.0003243907, 0.0003251439,
  0.00111781, 0.001255709, 0.001310091, 0.001158166, 0.0009967927, 
    0.0005496881, 0.0006264641, 0.0008827169, 0.00124621, 0.001112587, 
    0.0008985429, 0.001151221, 0.001217854, 0.0009927083, 0.0009104236,
  0.001317111, 0.001280582, 0.001311975, 0.001492234, 0.001223312, 
    0.0004590916, 0.0005358015, 0.0006158284, 0.0008930475, 0.001106367, 
    0.001213307, 0.001570572, 0.001578072, 0.001069962, 0.0008973698,
  0.001808091, 0.001528183, 0.001474429, 0.00162762, 0.001521996, 
    0.0006892555, 0.0004818226, 0.0005052597, 0.000579291, 0.0006709707, 
    0.0009520277, 0.001223143, 0.001436836, 0.001500944, 0.001301369,
  0.001983375, 0.001920858, 0.001806155, 0.001759692, 0.001729712, 
    0.001575775, 0.0005603743, 0.0004814407, 0.0005244231, 0.0005031041, 
    0.0005537754, 0.0008224495, 0.001040511, 0.001168082, 0.001122892,
  0.002024458, 0.001961735, 0.001883381, 0.001951863, 0.00176889, 
    0.001781991, 0.001497917, 0.0004587717, 0.0003173932, 0.0004150133, 
    0.000439359, 0.0005118366, 0.000696922, 0.0008662255, 0.001015644,
  0.002050909, 0.002017063, 0.001936559, 0.001972088, 0.002017697, 
    0.001750838, 0.001455763, 0.001192424, 0.0007396257, 0.0004971298, 
    0.000365536, 0.0004159934, 0.0004626866, 0.0005900572, 0.0007303155,
  0.002051453, 0.002048595, 0.001997766, 0.001920981, 0.001986589, 
    0.002014553, 0.001298648, 0.0009712565, 0.0007182927, 0.0006042273, 
    0.0004644264, 0.0003679558, 0.0003688473, 0.0004279824, 0.0005311299,
  0.002054484, 0.002063713, 0.002048116, 0.001945387, 0.001860833, 
    0.001858885, 0.001281658, 0.0008693836, 0.0006644891, 0.0006125896, 
    0.0005108429, 0.0003622507, 0.0003126371, 0.0003577459, 0.0004305893,
  0.002080595, 0.002103183, 0.002099436, 0.001993829, 0.001820431, 
    0.001705031, 0.001130497, 0.0007735031, 0.0005926779, 0.0005121005, 
    0.0004482247, 0.0003780789, 0.0003141874, 0.0003206725, 0.0003692629,
  0.002109462, 0.002135679, 0.002159531, 0.0019408, 0.001462594, 0.001261047, 
    0.0009249378, 0.0007551391, 0.0005181837, 0.0004485158, 0.0005280533, 
    0.000374547, 0.0003052806, 0.0002922487, 0.0003265309,
  0.001230475, 0.001203414, 0.001203597, 0.001264527, 0.001138255, 
    0.0006815317, 0.0005595648, 0.0006225819, 0.0009751492, 0.001187163, 
    0.001226355, 0.001338986, 0.001215216, 0.0007791803, 0.0007118567,
  0.00172923, 0.001272071, 0.001296159, 0.001363962, 0.001158862, 
    0.0005959668, 0.0005420545, 0.0005585329, 0.0006650078, 0.000893132, 
    0.001174107, 0.001396803, 0.001308426, 0.001117904, 0.0008857357,
  0.002119131, 0.001560262, 0.00134131, 0.001463989, 0.001316777, 
    0.0007599687, 0.000545878, 0.0004885035, 0.000529058, 0.0005966622, 
    0.0006988025, 0.0008423495, 0.0009332428, 0.0009482253, 0.0009212002,
  0.002135239, 0.002122917, 0.001785622, 0.00157733, 0.001509647, 
    0.001305247, 0.0007575731, 0.0005131818, 0.0005149741, 0.0004827103, 
    0.0005809863, 0.000630582, 0.0006406901, 0.0006386392, 0.0006250623,
  0.002243398, 0.002183509, 0.002007984, 0.001743691, 0.001599617, 
    0.001564817, 0.001420164, 0.0008547282, 0.0007477304, 0.000446454, 
    0.0004692003, 0.000520591, 0.0005618276, 0.0005566038, 0.0005661027,
  0.002356319, 0.002285663, 0.002187089, 0.00190301, 0.001722428, 
    0.001678037, 0.001672695, 0.001589797, 0.00107523, 0.0006749837, 
    0.0004264342, 0.0004313, 0.0004313913, 0.0004861394, 0.000526095,
  0.002443274, 0.002382699, 0.002331797, 0.002124125, 0.001893936, 
    0.00183077, 0.001711191, 0.001414555, 0.0009811968, 0.0006341342, 
    0.0004842067, 0.0004209684, 0.0003721169, 0.0004108412, 0.0004974366,
  0.002401232, 0.002409314, 0.002395139, 0.002282013, 0.002017599, 
    0.001860389, 0.001853379, 0.001239212, 0.0007419903, 0.0005785726, 
    0.0004488661, 0.0003899981, 0.000304478, 0.0003652088, 0.0004813352,
  0.002277443, 0.002353478, 0.002395521, 0.00234675, 0.002126766, 
    0.002021969, 0.001728747, 0.001044531, 0.000639692, 0.0005380626, 
    0.0004149127, 0.0003802309, 0.0002787624, 0.0003315173, 0.0004453424,
  0.002226796, 0.002323685, 0.002464361, 0.002342869, 0.002042459, 
    0.001930092, 0.001481556, 0.0008215974, 0.0005509335, 0.000463242, 
    0.000421913, 0.0003388217, 0.0002657373, 0.0002849407, 0.0003868696,
  0.002017991, 0.001870029, 0.001459422, 0.001225164, 0.0009337231, 
    0.0008392639, 0.0009618272, 0.001132891, 0.00124507, 0.001200785, 
    0.001184019, 0.001172165, 0.001089993, 0.0008049131, 0.0006287515,
  0.002215037, 0.001957225, 0.001448684, 0.001100042, 0.0007706279, 
    0.0006684245, 0.0008785174, 0.001061039, 0.001204199, 0.001288189, 
    0.001302832, 0.001300818, 0.001191158, 0.0006028782, 0.0006041392,
  0.002451937, 0.002137207, 0.001484349, 0.001181403, 0.0009129557, 
    0.000537499, 0.0006738589, 0.0008412594, 0.001040383, 0.00111911, 
    0.001161401, 0.001086162, 0.0009086547, 0.000767834, 0.000504423,
  0.002389753, 0.002379254, 0.001712484, 0.001274924, 0.001081256, 
    0.0009357628, 0.0005663992, 0.0006828886, 0.0007594756, 0.0008349826, 
    0.0008698109, 0.0007485589, 0.000696534, 0.0006407787, 0.0005229144,
  0.002295776, 0.002362304, 0.001839933, 0.001492798, 0.001146557, 
    0.00110511, 0.0009668241, 0.0005538448, 0.0005624032, 0.000571379, 
    0.000651039, 0.00066213, 0.0006462955, 0.0005988895, 0.0005458863,
  0.002239395, 0.00241837, 0.001915001, 0.001572488, 0.001312818, 
    0.001174659, 0.001103383, 0.001094191, 0.001009285, 0.0007001462, 
    0.0005604736, 0.000558293, 0.0005330345, 0.0005016355, 0.000522305,
  0.002270832, 0.002441358, 0.002066532, 0.001667642, 0.001580383, 
    0.001426633, 0.001279454, 0.001342387, 0.0009961835, 0.0006920836, 
    0.0005915611, 0.0005065778, 0.0004314363, 0.0004327528, 0.000511064,
  0.002298185, 0.002455521, 0.002154669, 0.001787172, 0.001631165, 
    0.001562684, 0.001468127, 0.00119555, 0.0008151279, 0.0006054206, 
    0.0004917046, 0.000403042, 0.0003251312, 0.0004113762, 0.0005133692,
  0.002362747, 0.002491688, 0.00225159, 0.001885046, 0.001716661, 
    0.001643978, 0.001552633, 0.001084001, 0.0006744064, 0.00051825, 
    0.0004050641, 0.0003257227, 0.0002758867, 0.0003681307, 0.0004773526,
  0.002498278, 0.002592649, 0.002464388, 0.002132835, 0.001734303, 
    0.001724698, 0.001472503, 0.0008466794, 0.0005312057, 0.000430539, 
    0.0003587687, 0.0002921286, 0.0002525074, 0.0003073652, 0.000427264,
  0.001951266, 0.002049258, 0.002012427, 0.001709447, 0.001087262, 
    0.0005869581, 0.0007672379, 0.0009931793, 0.001049459, 0.0008875585, 
    0.0008304305, 0.0007771081, 0.000721704, 0.0006445663, 0.0004865573,
  0.002213022, 0.0021945, 0.002088708, 0.001529562, 0.0008752351, 
    0.0004941225, 0.0006847664, 0.0009513267, 0.001112066, 0.001086662, 
    0.0009876962, 0.000941917, 0.0008608068, 0.0005629021, 0.0005015853,
  0.002326432, 0.00234272, 0.002025749, 0.001452598, 0.001004952, 
    0.0004918188, 0.0006125927, 0.0008932625, 0.001121092, 0.001214008, 
    0.001147341, 0.001030609, 0.0009225996, 0.0008401438, 0.0006355738,
  0.002392712, 0.002424931, 0.002203015, 0.001382795, 0.001126124, 
    0.001007062, 0.0005398131, 0.0008093247, 0.000960212, 0.001083471, 
    0.001039768, 0.0009073435, 0.0008340388, 0.000742292, 0.0005687833,
  0.002443549, 0.002424401, 0.002117525, 0.001462073, 0.001061822, 
    0.001086317, 0.00104511, 0.0005522514, 0.0005423598, 0.0007527765, 
    0.0008072983, 0.0007446968, 0.0007241724, 0.0006678167, 0.0006081357,
  0.00252843, 0.002438741, 0.001968428, 0.001441915, 0.001175751, 
    0.0009787232, 0.00107133, 0.001119119, 0.0008668688, 0.0007195615, 
    0.0006515793, 0.0006446354, 0.0006379443, 0.0006329961, 0.0006086548,
  0.002525654, 0.002341371, 0.001819815, 0.001456494, 0.001354163, 
    0.001234253, 0.001099505, 0.0009648922, 0.0007830376, 0.0006865684, 
    0.0005988221, 0.0005603948, 0.0005646744, 0.0005776195, 0.0005698181,
  0.002428381, 0.002218348, 0.001717926, 0.001487015, 0.00142532, 
    0.001400517, 0.001013978, 0.0008348034, 0.000667141, 0.0005907334, 
    0.0005009044, 0.0004710081, 0.0004400183, 0.0004990011, 0.0005431903,
  0.002318941, 0.002055935, 0.001683423, 0.001539757, 0.001515653, 
    0.001321558, 0.0008717534, 0.0007335859, 0.0005550496, 0.0004630602, 
    0.000398468, 0.0003746646, 0.0003469823, 0.0004458477, 0.0004792541,
  0.002244136, 0.002017824, 0.001753278, 0.001680854, 0.001202228, 
    0.001052038, 0.0007566992, 0.0006142239, 0.0004645511, 0.0003726457, 
    0.0003263428, 0.0003224973, 0.0002952228, 0.0003689563, 0.0004286015,
  0.002377272, 0.002460612, 0.002472619, 0.002422248, 0.002331149, 
    0.002034876, 0.001662813, 0.0014164, 0.001189913, 0.0008449402, 
    0.0007990356, 0.0007953385, 0.000721753, 0.0007075733, 0.0005932546,
  0.00264369, 0.002610534, 0.002499936, 0.002345009, 0.002022746, 0.00122084, 
    0.001068612, 0.000937066, 0.0009074023, 0.0008866591, 0.0008570227, 
    0.0008983294, 0.0008618737, 0.0006291463, 0.0005290802,
  0.002607807, 0.002490164, 0.002268687, 0.002018384, 0.001470515, 
    0.0008402144, 0.0008859165, 0.0009341282, 0.0008918006, 0.000920364, 
    0.000924224, 0.0009298891, 0.0009353556, 0.0009276645, 0.0007182309,
  0.002322913, 0.002186685, 0.001980103, 0.001656647, 0.001332643, 
    0.001016366, 0.0006535868, 0.000754795, 0.0007146394, 0.0007841114, 
    0.0008163132, 0.000882169, 0.0009519254, 0.0009444479, 0.0007577699,
  0.002050645, 0.00194738, 0.001823999, 0.001512928, 0.001202449, 0.00113792, 
    0.001055053, 0.0005494541, 0.0004064198, 0.000667811, 0.0007843638, 
    0.0008619613, 0.0009360203, 0.0009128299, 0.0007732642,
  0.001916088, 0.001740558, 0.001580448, 0.001380378, 0.001188335, 
    0.00108881, 0.001058543, 0.001014496, 0.0008737723, 0.0007329892, 
    0.0007466403, 0.000839707, 0.0008792908, 0.0008330938, 0.0007409381,
  0.001782773, 0.001624968, 0.001480635, 0.001336702, 0.001231214, 
    0.001085834, 0.0009620049, 0.0008906795, 0.0007808362, 0.0007552212, 
    0.0007684331, 0.000794357, 0.0007925308, 0.0007422456, 0.0006938882,
  0.001695895, 0.001586156, 0.001453183, 0.00134903, 0.001291174, 
    0.001154706, 0.0008386388, 0.0007542982, 0.0006996089, 0.0006959334, 
    0.000699502, 0.0007135955, 0.0006946589, 0.0006822253, 0.0006386921,
  0.00171947, 0.001614927, 0.001488826, 0.001345778, 0.001213772, 
    0.0009532992, 0.0007005081, 0.000633059, 0.0005949749, 0.0005966555, 
    0.0006010482, 0.0006041003, 0.0005842394, 0.0005696241, 0.0004761631,
  0.001759125, 0.001642888, 0.001468306, 0.0009917313, 0.0007952874, 
    0.0007179255, 0.0006230433, 0.0005543083, 0.0004933972, 0.0004714997, 
    0.0004788772, 0.0004989338, 0.0004637418, 0.0004401315, 0.0004080656,
  0.00161198, 0.00152262, 0.001312623, 0.001191315, 0.001208979, 0.001007911, 
    0.0008731415, 0.0008795007, 0.0009421796, 0.0009443749, 0.0009305333, 
    0.0009375758, 0.001014129, 0.001152883, 0.001108293,
  0.001719968, 0.001512815, 0.001289079, 0.001114953, 0.001024709, 
    0.0008692474, 0.0007634101, 0.0006631343, 0.0007696607, 0.0008354838, 
    0.0007905397, 0.0008675578, 0.0008311736, 0.0006534219, 0.0008228389,
  0.001879052, 0.001518154, 0.001252199, 0.001141159, 0.001006713, 
    0.0007384457, 0.000714926, 0.0006778566, 0.0007440093, 0.0008285051, 
    0.0008880025, 0.0008919197, 0.0008549558, 0.0008880214, 0.0008760106,
  0.001841984, 0.001591951, 0.001338691, 0.001172734, 0.001005043, 
    0.000895082, 0.000588421, 0.0005787453, 0.000651709, 0.0007975307, 
    0.0009094933, 0.0009642822, 0.0008858835, 0.0008855279, 0.0008636959,
  0.001867131, 0.001589751, 0.001395866, 0.001178148, 0.001015249, 
    0.0008894111, 0.0008551871, 0.0004309434, 0.0004687386, 0.0007242825, 
    0.0008770856, 0.0009336999, 0.0009453263, 0.0009137665, 0.0008566302,
  0.001891735, 0.001617021, 0.001401353, 0.001199572, 0.001019216, 
    0.0008485071, 0.0007976954, 0.0007501081, 0.0007347471, 0.0008630308, 
    0.0008613874, 0.0009531502, 0.0009742467, 0.000910331, 0.0008197959,
  0.001909434, 0.001666584, 0.001457695, 0.001249832, 0.001150178, 
    0.0009284234, 0.0007180147, 0.0007119391, 0.0007676648, 0.0009099395, 
    0.0009631139, 0.0009573855, 0.0009430978, 0.0008706667, 0.0008028957,
  0.001943578, 0.001732538, 0.001491085, 0.001276562, 0.001196458, 
    0.001003821, 0.0006711011, 0.0006492372, 0.0006523965, 0.000766155, 
    0.0008761779, 0.0009087939, 0.0008714325, 0.0007931128, 0.0007439881,
  0.002009646, 0.001747329, 0.001510915, 0.001228465, 0.00104588, 
    0.0007776379, 0.0006319786, 0.0006154765, 0.0005992246, 0.0006091037, 
    0.0006712403, 0.0006949503, 0.0006713447, 0.0006250993, 0.0005346395,
  0.002078133, 0.001829791, 0.001477004, 0.0008949405, 0.0006769074, 
    0.0006157926, 0.000596309, 0.0005928189, 0.0005406184, 0.0005000343, 
    0.0005078209, 0.0005506317, 0.0005387895, 0.0005141385, 0.0004752348,
  0.001904575, 0.001700556, 0.001287191, 0.00108416, 0.0009447274, 
    0.0006763662, 0.0006448628, 0.0006191005, 0.0007220629, 0.0007156762, 
    0.0007778588, 0.0008913815, 0.0008847368, 0.0008311799, 0.0008909944,
  0.002344269, 0.001828219, 0.001437836, 0.001108119, 0.0008851351, 
    0.00058777, 0.0006379056, 0.0006104137, 0.0007178515, 0.0008459137, 
    0.0008527303, 0.001007385, 0.0009855507, 0.0006878111, 0.0008527417,
  0.00256523, 0.001918092, 0.001502559, 0.001128744, 0.0009282115, 
    0.0005211084, 0.0006008879, 0.0006799973, 0.000802343, 0.0009250853, 
    0.0009933783, 0.001020287, 0.001005198, 0.00102627, 0.001095871,
  0.002667002, 0.002239703, 0.001679251, 0.001221667, 0.001002215, 
    0.0007709306, 0.0004845785, 0.0005627354, 0.0007387408, 0.0009341124, 
    0.001016791, 0.001027416, 0.001022507, 0.001039054, 0.000974199,
  0.002917876, 0.002465901, 0.001899651, 0.001327826, 0.0009981729, 
    0.0007837531, 0.0007315332, 0.0003949188, 0.0005626506, 0.0008525462, 
    0.0009708612, 0.0009968219, 0.001001771, 0.0009830057, 0.00095339,
  0.003147508, 0.002784358, 0.002142752, 0.001516102, 0.001118258, 
    0.0007729478, 0.0006979538, 0.0006550129, 0.0007342866, 0.0008608249, 
    0.0008497908, 0.0009412091, 0.0009659376, 0.0009298858, 0.0008830112,
  0.003385325, 0.003097618, 0.002529769, 0.001737368, 0.001316929, 
    0.000951752, 0.0006597834, 0.0006422239, 0.0006759538, 0.0007763018, 
    0.000789923, 0.0008324093, 0.0008548695, 0.0008367079, 0.0007972993,
  0.003596723, 0.00335516, 0.002905269, 0.002036594, 0.00145263, 0.001060254, 
    0.0006450261, 0.0006031657, 0.0005746305, 0.0006202371, 0.0006498238, 
    0.0006853257, 0.0006827031, 0.0006819282, 0.000654544,
  0.003766105, 0.003558737, 0.003205968, 0.002463904, 0.001605036, 
    0.000929892, 0.0006382565, 0.000588619, 0.0005281198, 0.0004803443, 
    0.0004983115, 0.000524291, 0.00054322, 0.0005428261, 0.0005006506,
  0.00382983, 0.003648069, 0.003301458, 0.002690512, 0.001616765, 
    0.0008104254, 0.0006350463, 0.0005950925, 0.0004701588, 0.000362481, 
    0.0003663411, 0.0004523518, 0.0004681914, 0.000500483, 0.0005369979,
  0.003589258, 0.003069437, 0.002029315, 0.001210774, 0.0007384885, 
    0.0005005234, 0.0004490084, 0.0005136208, 0.0008047348, 0.0007747687, 
    0.000839164, 0.0008885839, 0.0007288604, 0.0006563858, 0.000500523,
  0.003625028, 0.002969195, 0.00191801, 0.001053109, 0.000651792, 
    0.0004477979, 0.0004870332, 0.00054799, 0.0007652032, 0.0008776246, 
    0.0008716864, 0.00103134, 0.0009579335, 0.0005902865, 0.0004078005,
  0.003570673, 0.002922822, 0.001850368, 0.001109867, 0.0008131618, 
    0.0004212557, 0.0004882502, 0.0006148732, 0.0008229468, 0.0009352501, 
    0.0009844017, 0.0009857184, 0.0009332309, 0.0008288722, 0.000736375,
  0.003720038, 0.003166733, 0.002159022, 0.001264341, 0.0009979189, 
    0.0008042902, 0.0003991735, 0.0005547234, 0.000694942, 0.000880677, 
    0.0009906451, 0.0009842854, 0.0009531521, 0.0009088552, 0.0008709874,
  0.003822675, 0.003216115, 0.00245388, 0.00147421, 0.001023002, 
    0.0009139127, 0.0008544769, 0.0004120239, 0.0005758793, 0.0007091288, 
    0.0008699928, 0.0009327912, 0.0009279074, 0.0008776907, 0.0008289074,
  0.003676945, 0.00330786, 0.002504741, 0.00162269, 0.001065352, 0.000874456, 
    0.0008162895, 0.000740419, 0.0006554796, 0.0007345562, 0.0007138686, 
    0.0008219648, 0.0008333994, 0.0008074583, 0.0007896387,
  0.003508082, 0.003200477, 0.002615046, 0.001760387, 0.001340842, 
    0.0009664918, 0.0007317612, 0.0006362522, 0.0006000409, 0.0006258981, 
    0.0006418684, 0.0007248248, 0.0007551207, 0.000767266, 0.0007697839,
  0.003315809, 0.003048013, 0.002655256, 0.001879591, 0.001520713, 
    0.001157071, 0.0006955708, 0.0006118018, 0.0005282519, 0.0004954804, 
    0.0005113464, 0.000575135, 0.0006151578, 0.0006743719, 0.0006763285,
  0.003145999, 0.002927236, 0.002667387, 0.001962037, 0.001554668, 
    0.001011364, 0.0006577063, 0.0005855576, 0.0004999475, 0.000443556, 
    0.0004513534, 0.0005097114, 0.000556592, 0.0006258979, 0.000646026,
  0.002995629, 0.002824452, 0.002532064, 0.00184049, 0.001230859, 
    0.0008026839, 0.0006711447, 0.0006146083, 0.0005056271, 0.0004044014, 
    0.0004185672, 0.0005290192, 0.0005805603, 0.0006428482, 0.0006841128,
  0.001255018, 0.0009093675, 0.0007445657, 0.0006883454, 0.0006342211, 
    0.0005935621, 0.0006615885, 0.0005099822, 0.0006022456, 0.000483344, 
    0.0005514912, 0.0006168347, 0.0005494026, 0.0004742463, 0.0004158733,
  0.001248007, 0.0009356985, 0.0008560162, 0.0007714835, 0.000677385, 
    0.000583168, 0.0006787112, 0.0005917646, 0.0006511435, 0.0006116066, 
    0.0005973116, 0.0007013446, 0.0006462407, 0.0003732153, 0.0003301636,
  0.001388733, 0.001021122, 0.0009411006, 0.0009312864, 0.0008539097, 
    0.0004942897, 0.0006235373, 0.0006826836, 0.0008045384, 0.00076551, 
    0.0007886252, 0.0007603976, 0.000675754, 0.0005783097, 0.0004708465,
  0.001570508, 0.001420249, 0.001180646, 0.001009395, 0.0009780327, 
    0.0008895074, 0.000571051, 0.0006410636, 0.0007263173, 0.0008260168, 
    0.0008818401, 0.0008681336, 0.0007855933, 0.0007050644, 0.0006010926,
  0.001646094, 0.001515618, 0.001424808, 0.001113197, 0.00100811, 
    0.0009694459, 0.0009238906, 0.000473456, 0.0005685543, 0.0007456848, 
    0.0008294933, 0.0008772094, 0.0008875646, 0.0008214274, 0.0007281164,
  0.001694029, 0.001557105, 0.001426508, 0.001228462, 0.001036852, 
    0.0008974667, 0.0008602149, 0.0007865605, 0.0007412031, 0.0007979457, 
    0.0007704106, 0.0008046225, 0.0008427865, 0.000857919, 0.0007976487,
  0.00173406, 0.001633845, 0.001526002, 0.001390398, 0.001313244, 
    0.0009627344, 0.0008235078, 0.0007834432, 0.0007741686, 0.0008062471, 
    0.0008518521, 0.0008414565, 0.0008217331, 0.0008414877, 0.0008434146,
  0.00176361, 0.001690138, 0.001590522, 0.001485878, 0.001413299, 
    0.001102946, 0.0008423148, 0.000801545, 0.0007563161, 0.0007653222, 
    0.0008421252, 0.0009205008, 0.0008941888, 0.0008680509, 0.0008665102,
  0.001789516, 0.001713494, 0.001583008, 0.001444705, 0.001281998, 
    0.0009890303, 0.0008792453, 0.0008440876, 0.0007770695, 0.0007419059, 
    0.00075232, 0.0009055078, 0.000966591, 0.0009598053, 0.0009460416,
  0.001761584, 0.001639823, 0.001425969, 0.001126218, 0.0009487774, 
    0.0009372723, 0.0009029029, 0.0008675854, 0.0007636906, 0.0006830014, 
    0.0006785047, 0.0007725714, 0.0009372034, 0.001019817, 0.001004726,
  0.00105142, 0.001036399, 0.0009677032, 0.0009397966, 0.0008138882, 
    0.000596525, 0.0005749064, 0.0005388296, 0.0005682071, 0.0003881711, 
    0.0004031649, 0.0005273013, 0.0005557218, 0.0005850081, 0.0006507518,
  0.001268767, 0.001119935, 0.001024377, 0.0009547278, 0.000810696, 
    0.0005867769, 0.0006269817, 0.0005881778, 0.0006586338, 0.0005254174, 
    0.0004205755, 0.0005650694, 0.0006580129, 0.000425585, 0.0004741231,
  0.001425364, 0.001313517, 0.001123072, 0.0009607191, 0.0008870423, 
    0.0005390471, 0.0006079383, 0.000643442, 0.0006980151, 0.0006979576, 
    0.0006112571, 0.0005737077, 0.0006347052, 0.0006614095, 0.0006142684,
  0.001515536, 0.001461024, 0.001314152, 0.001009537, 0.0009176117, 
    0.0007990326, 0.0005342376, 0.0005604847, 0.0006848972, 0.0007065622, 
    0.00073349, 0.0006226744, 0.0006106888, 0.0006532872, 0.0006028943,
  0.001596784, 0.001534377, 0.001437653, 0.001121622, 0.0009268043, 
    0.0008234644, 0.0007550019, 0.0004222323, 0.0005040216, 0.0006843514, 
    0.0006794287, 0.0006940038, 0.0006253918, 0.0006314315, 0.0006325062,
  0.001640476, 0.001574459, 0.001440885, 0.00121165, 0.001025685, 
    0.0007941153, 0.0007278734, 0.0006424772, 0.0006453866, 0.0008102487, 
    0.0006088343, 0.0007462534, 0.000691171, 0.000630661, 0.0006041096,
  0.001671516, 0.001602279, 0.001496779, 0.001292141, 0.00118244, 
    0.0008373785, 0.0007167908, 0.0006447837, 0.0006449363, 0.0008030799, 
    0.0007929649, 0.0007522337, 0.0007310984, 0.0006750022, 0.0006006518,
  0.001652518, 0.001576993, 0.001456988, 0.00133398, 0.001199241, 
    0.0008802766, 0.0007178247, 0.0006323771, 0.0005646136, 0.0006271283, 
    0.0008480641, 0.0008376854, 0.0007273451, 0.0007312993, 0.0006529929,
  0.001596109, 0.001504444, 0.001349463, 0.001167079, 0.000931591, 
    0.0007139514, 0.0007034824, 0.0006648615, 0.0005592393, 0.0005570815, 
    0.0006404204, 0.0009047274, 0.0008828918, 0.0008025714, 0.0007480159,
  0.001467225, 0.001331734, 0.001125628, 0.0007582949, 0.0006021328, 
    0.0006007156, 0.0006111335, 0.0006904941, 0.000551102, 0.0004845251, 
    0.0005119936, 0.0006951869, 0.0009361113, 0.0009386976, 0.0008438092,
  0.0009472769, 0.0009058112, 0.0008424453, 0.0008046235, 0.0006714729, 
    0.0004789553, 0.0004532833, 0.0004814663, 0.0005243015, 0.0004612073, 
    0.0004474945, 0.0004602661, 0.000416672, 0.0004531701, 0.0004300257,
  0.00112471, 0.0009686805, 0.0008872023, 0.0008194909, 0.0007276097, 
    0.0004358596, 0.0004582766, 0.0004797229, 0.0005439153, 0.0005509281, 
    0.0004791189, 0.0005384573, 0.0006020165, 0.0004414637, 0.0003884858,
  0.00140199, 0.00109804, 0.0009082519, 0.000804381, 0.0007485097, 
    0.0004695918, 0.0004710156, 0.0005055488, 0.0005579318, 0.0005857142, 
    0.0006084812, 0.000600192, 0.0006162696, 0.0006550269, 0.000628482,
  0.00132285, 0.001197729, 0.001000918, 0.0008055926, 0.0007281876, 
    0.0006571552, 0.0004065652, 0.0004602324, 0.0005362362, 0.000676411, 
    0.0006951056, 0.0006681572, 0.0006391446, 0.0006660682, 0.0006511753,
  0.001353053, 0.001233696, 0.001083071, 0.0008270033, 0.0007284746, 
    0.0006391299, 0.0005751328, 0.000309832, 0.0003766604, 0.0006317717, 
    0.0007270314, 0.0006767458, 0.0006201423, 0.0006552034, 0.0007209104,
  0.001360598, 0.001263699, 0.001091609, 0.0008984182, 0.0007661585, 
    0.0006157244, 0.0005821352, 0.0005096999, 0.0005301441, 0.0006710888, 
    0.0006482523, 0.0006057793, 0.0005827729, 0.0006467005, 0.0006788574,
  0.001359199, 0.001277826, 0.001165542, 0.001010634, 0.0009232913, 
    0.0006304019, 0.0005787765, 0.0005414042, 0.0005737385, 0.0007257247, 
    0.0007235698, 0.0005722637, 0.0005432994, 0.0005882472, 0.0006154954,
  0.00132912, 0.001263879, 0.001194058, 0.001113118, 0.0009737053, 
    0.0006447543, 0.0005652161, 0.0005435412, 0.0005463476, 0.0006801374, 
    0.0007100469, 0.0006055965, 0.0005138205, 0.0005269899, 0.0005548963,
  0.001300915, 0.00123129, 0.001137088, 0.0009781546, 0.0007016059, 
    0.0005299671, 0.0005474304, 0.0005598607, 0.0005416375, 0.000625092, 
    0.0007151364, 0.0006809713, 0.0005238838, 0.0005280161, 0.0005096583,
  0.001287223, 0.001142804, 0.0009277884, 0.0005823972, 0.0004725026, 
    0.0004545295, 0.0004774937, 0.0006295143, 0.000553059, 0.0005149716, 
    0.0006038379, 0.0007391288, 0.0006383123, 0.000526719, 0.0005142727,
  0.0007476927, 0.0007859663, 0.0007243161, 0.0006722991, 0.0005794151, 
    0.0004700169, 0.0004394657, 0.0003957782, 0.0004030085, 0.0003610807, 
    0.0004430497, 0.0004599231, 0.0003918952, 0.0003850904, 0.000369333,
  0.0008772985, 0.0007997387, 0.0007759221, 0.0007044197, 0.0005811552, 
    0.000392423, 0.0004231266, 0.0004138559, 0.0004204716, 0.0004597994, 
    0.000481745, 0.0004958143, 0.0004923136, 0.0004165353, 0.0003264058,
  0.001055908, 0.0008112363, 0.0007659335, 0.0007607116, 0.0006635159, 
    0.0003706959, 0.000429914, 0.000436849, 0.0004318441, 0.0005013405, 
    0.000580008, 0.0005806905, 0.0005503968, 0.0005022069, 0.0004237457,
  0.001133015, 0.00100067, 0.0008926823, 0.00073253, 0.0006857108, 
    0.0006099236, 0.0003562837, 0.0004682188, 0.0005028166, 0.0005793279, 
    0.0006636269, 0.0006931036, 0.0006602438, 0.0006173151, 0.000546707,
  0.001124468, 0.001067062, 0.0009670703, 0.0007803343, 0.0007031055, 
    0.0006193497, 0.0005807237, 0.0002927426, 0.0003763178, 0.0006228992, 
    0.0007076288, 0.0007009389, 0.0006982088, 0.0006936839, 0.0006728509,
  0.001132765, 0.001065169, 0.0009743075, 0.0008376734, 0.0007573247, 
    0.0006230649, 0.0005956122, 0.0005531119, 0.0005376263, 0.0006107982, 
    0.0006058226, 0.0006587427, 0.0006804266, 0.0006646266, 0.0006625896,
  0.00112009, 0.001097358, 0.001020247, 0.000943715, 0.0008894454, 
    0.0006396307, 0.0005764881, 0.0005511024, 0.0005448625, 0.0006082985, 
    0.0006070001, 0.0005457225, 0.0005634956, 0.0006059438, 0.0006135138,
  0.001155886, 0.001103839, 0.001071601, 0.001032795, 0.0009487614, 
    0.0006710792, 0.0005725309, 0.0005485864, 0.0005099563, 0.0005177518, 
    0.0005154228, 0.0005217538, 0.0005580965, 0.0006185339, 0.0006138132,
  0.001193975, 0.001103297, 0.001085614, 0.0009997139, 0.0007915088, 
    0.0006350927, 0.0005763255, 0.0005804567, 0.0005315288, 0.0004975469, 
    0.0004650951, 0.0005158656, 0.0005255165, 0.0006032545, 0.0005852731,
  0.00118562, 0.00112228, 0.001046482, 0.0008395472, 0.0007333658, 
    0.0006575939, 0.0005942706, 0.0007116654, 0.0005852801, 0.0004201838, 
    0.000348485, 0.000433802, 0.0004956418, 0.0005744825, 0.0005707838,
  0.0007127001, 0.0006903253, 0.0006112379, 0.0005912379, 0.0004889209, 
    0.000364624, 0.0003956069, 0.0004099735, 0.0004389174, 0.000367658, 
    0.0004260733, 0.0004977189, 0.0004751761, 0.0005105597, 0.0005422946,
  0.0007820532, 0.0007415753, 0.0007228855, 0.0007143551, 0.0006069371, 
    0.0004485995, 0.0004584765, 0.0004583816, 0.0004758557, 0.0004419604, 
    0.0004372821, 0.0004773112, 0.0005041888, 0.0004258989, 0.0004209753,
  0.001174847, 0.0009620452, 0.0008692938, 0.0008848684, 0.0008246343, 
    0.0004927136, 0.0005040477, 0.0005278556, 0.0004917044, 0.000513681, 
    0.0005369427, 0.0005216391, 0.0005084919, 0.000495391, 0.0004467555,
  0.001450406, 0.001485385, 0.001509691, 0.00125653, 0.001163609, 
    0.0009840134, 0.0006179939, 0.0006023913, 0.0005800461, 0.0006076497, 
    0.0006214461, 0.0006288015, 0.0006050807, 0.0005796887, 0.0005021132,
  0.001503986, 0.001583698, 0.001663161, 0.001616116, 0.001532139, 
    0.001361678, 0.001141666, 0.0006468134, 0.0005346916, 0.0006526398, 
    0.0006986875, 0.0006778962, 0.0006618379, 0.0006534968, 0.000624544,
  0.001710644, 0.001825034, 0.001816887, 0.001795855, 0.001715303, 
    0.001472826, 0.001245672, 0.00101565, 0.0008045602, 0.0006928645, 
    0.0006843804, 0.000677089, 0.0006554977, 0.0006639578, 0.0006567809,
  0.001976311, 0.001994282, 0.001877939, 0.001729865, 0.001582378, 
    0.001356972, 0.001128341, 0.0009661631, 0.0007745828, 0.0006677688, 
    0.0006008255, 0.0005979902, 0.0006128644, 0.000633633, 0.0006460434,
  0.002149164, 0.002027142, 0.001780328, 0.001625856, 0.001470273, 
    0.001204902, 0.0009845544, 0.0008297953, 0.0006940794, 0.0006096539, 
    0.0005598153, 0.0005239526, 0.000520355, 0.0005645634, 0.0005991564,
  0.002159569, 0.001916633, 0.001725595, 0.001535237, 0.001263131, 
    0.001022503, 0.0008232666, 0.0007380693, 0.0006503778, 0.0005685089, 
    0.0005113709, 0.0004831067, 0.0004801393, 0.0005155943, 0.0005538065,
  0.002066573, 0.001864755, 0.001642146, 0.001338032, 0.001067784, 
    0.0008521616, 0.0006818335, 0.000676254, 0.0006028894, 0.000503752, 
    0.0004498713, 0.0004416149, 0.000431073, 0.0004580593, 0.0004945492,
  0.001185783, 0.001180058, 0.001209894, 0.001183774, 0.0009628521, 
    0.0006526145, 0.000574505, 0.0005062557, 0.0004780627, 0.0003626005, 
    0.0003912115, 0.00043643, 0.0003744526, 0.0003965333, 0.0003531089,
  0.001402697, 0.001342749, 0.001352541, 0.001418527, 0.001174317, 
    0.001014004, 0.000931195, 0.0008380773, 0.0006875253, 0.0006052094, 
    0.000582164, 0.0005881114, 0.0005515824, 0.000430297, 0.00038688,
  0.00177664, 0.001674295, 0.001778335, 0.002042238, 0.001785716, 
    0.001571573, 0.001224819, 0.0009615127, 0.0008598232, 0.0007974796, 
    0.0007187006, 0.0007229695, 0.0006510311, 0.0005742349, 0.0004950191,
  0.001748419, 0.00205356, 0.002476169, 0.002496722, 0.002303728, 
    0.001834846, 0.00107548, 0.0009316236, 0.0008767149, 0.000810112, 
    0.0007984892, 0.0007530668, 0.0007014382, 0.0007134379, 0.0006523159,
  0.002035195, 0.00238526, 0.002642585, 0.00254891, 0.002024498, 0.001560354, 
    0.001178064, 0.0006472599, 0.0006172406, 0.0007296733, 0.0007707749, 
    0.0007395913, 0.0007070366, 0.0007044058, 0.0006922607,
  0.002473089, 0.002631937, 0.002649725, 0.002246372, 0.001830969, 
    0.001433512, 0.00124088, 0.0009586959, 0.0007108211, 0.0005440969, 
    0.0005843801, 0.000580802, 0.0005765079, 0.0005975054, 0.0006343157,
  0.002657731, 0.002543022, 0.002204242, 0.001830234, 0.001616372, 
    0.001307917, 0.0009939063, 0.0007434878, 0.0005823079, 0.0004802371, 
    0.0004625547, 0.000476183, 0.0004807632, 0.0004888787, 0.0005265286,
  0.002530755, 0.002232945, 0.001933358, 0.001634933, 0.001377143, 
    0.0008507821, 0.0005911979, 0.0005086185, 0.0004810452, 0.0004544097, 
    0.0004534351, 0.0004607714, 0.0004623398, 0.0004484611, 0.000472496,
  0.002265769, 0.002036655, 0.001718097, 0.00135856, 0.0009106269, 
    0.000589897, 0.0004814447, 0.0004895604, 0.000510965, 0.0004844301, 
    0.0004653594, 0.0004433124, 0.000430438, 0.0004112076, 0.0004181283,
  0.002097805, 0.001785024, 0.001443688, 0.0009189653, 0.0006385842, 
    0.0004615872, 0.0004153854, 0.0005207103, 0.0005031731, 0.0004320835, 
    0.0004422799, 0.0004319599, 0.0003824356, 0.000358322, 0.000374336,
  0.001134202, 0.001088975, 0.001119272, 0.001158469, 0.001435994, 
    0.001574167, 0.001944311, 0.001628883, 0.001299222, 0.0009334955, 
    0.0008560192, 0.0007961497, 0.0005869456, 0.0005205133, 0.0004621269,
  0.001195608, 0.001185746, 0.001190973, 0.001342269, 0.001567886, 
    0.001613091, 0.001946123, 0.00149253, 0.001341195, 0.001125935, 
    0.001008449, 0.001006146, 0.0009199283, 0.0007543216, 0.0006903257,
  0.001385427, 0.001440848, 0.001573476, 0.001976928, 0.002204719, 
    0.001924371, 0.001431606, 0.001213441, 0.001038908, 0.0009102431, 
    0.0008385472, 0.0009021432, 0.0008654587, 0.0008353696, 0.0007485675,
  0.001611964, 0.001851562, 0.002312985, 0.00248649, 0.002124323, 
    0.001317915, 0.0008679762, 0.0008255879, 0.000777462, 0.0007167021, 
    0.0007187008, 0.0007303948, 0.0007364224, 0.0007664124, 0.0007809128,
  0.001870797, 0.002306619, 0.002595197, 0.001964329, 0.001104985, 
    0.0008807656, 0.0008309454, 0.0005485353, 0.0005534069, 0.000632481, 
    0.0007003968, 0.0007033886, 0.0006830906, 0.0007017827, 0.0007510424,
  0.002454967, 0.002708749, 0.002411936, 0.001424142, 0.0009844011, 
    0.0006473728, 0.0005706962, 0.0005276168, 0.000485547, 0.0004189049, 
    0.0004908352, 0.0005646378, 0.0005660814, 0.0005964296, 0.0006276412,
  0.002750733, 0.002540268, 0.001782308, 0.001109686, 0.0009213192, 
    0.0006178207, 0.0005086307, 0.0004676901, 0.0004372009, 0.0004105709, 
    0.0004093241, 0.0004176408, 0.0004361186, 0.0004419606, 0.0004499367,
  0.002573509, 0.001784062, 0.001201117, 0.0009803547, 0.0008843828, 
    0.0005893902, 0.0005084023, 0.0004925668, 0.0004770661, 0.0004552006, 
    0.0004416632, 0.0004353325, 0.0004289931, 0.0004248405, 0.0004270697,
  0.002079122, 0.001363251, 0.001070751, 0.0008714659, 0.0005976395, 
    0.0005311367, 0.0005177338, 0.000535309, 0.0005259035, 0.0004993952, 
    0.0004663066, 0.0004379739, 0.0004510054, 0.0004660822, 0.0004449423,
  0.001651964, 0.0010983, 0.0008748528, 0.0005978745, 0.0005703925, 
    0.000545315, 0.0005473082, 0.0005794812, 0.0005394064, 0.0004486525, 
    0.0004245633, 0.0004255733, 0.0004677036, 0.0005030665, 0.0004380641,
  0.001173823, 0.00119557, 0.001140871, 0.001101278, 0.001034363, 
    0.001032407, 0.001252667, 0.001407561, 0.001259979, 0.0009098929, 
    0.000678023, 0.0005410404, 0.0004641312, 0.0004747481, 0.0004611165,
  0.001358565, 0.001282357, 0.00121462, 0.00116216, 0.001031109, 0.001060379, 
    0.001302572, 0.001103654, 0.0007865817, 0.0006507816, 0.0005122678, 
    0.0004980351, 0.0004827795, 0.0004167954, 0.0004369623,
  0.001852906, 0.001570006, 0.001385774, 0.001357027, 0.001393193, 
    0.00130767, 0.001150428, 0.0009021197, 0.0006937459, 0.0005906138, 
    0.0005338745, 0.0005098424, 0.0004948027, 0.0004710268, 0.0004486278,
  0.001886868, 0.0019993, 0.001970454, 0.001953598, 0.001875336, 0.001663873, 
    0.000938239, 0.0007219878, 0.0006154592, 0.0005836037, 0.0005657987, 
    0.0005317205, 0.0005004573, 0.0004792694, 0.000447111,
  0.001827663, 0.001915903, 0.00207039, 0.002097425, 0.001762756, 
    0.001509792, 0.00111828, 0.000559333, 0.0004620798, 0.0005507903, 
    0.0005734633, 0.0005242006, 0.0004832358, 0.0004661984, 0.0004536381,
  0.001850314, 0.001999489, 0.002165223, 0.002130813, 0.001827117, 
    0.001407937, 0.001132915, 0.0007287192, 0.0005377593, 0.0004077468, 
    0.0004047026, 0.0004706768, 0.0004666906, 0.0004511181, 0.0004350398,
  0.002068688, 0.002250417, 0.002287293, 0.002014319, 0.001774267, 
    0.001321366, 0.0007893017, 0.0005428245, 0.0004780211, 0.0004504058, 
    0.000485172, 0.0004775341, 0.0004621043, 0.0004287164, 0.0004137484,
  0.002532829, 0.002514478, 0.002244606, 0.001922373, 0.001662571, 
    0.0008440498, 0.0005806817, 0.000521721, 0.0005342234, 0.000523204, 
    0.0005145639, 0.0004725125, 0.0004233554, 0.0004003675, 0.0004215407,
  0.002985447, 0.002732621, 0.002267346, 0.001689137, 0.001011543, 
    0.000666698, 0.000572257, 0.0005824763, 0.000588234, 0.000569593, 
    0.0004777662, 0.0004020531, 0.0003873868, 0.0004070091, 0.0004294726,
  0.002764169, 0.002568285, 0.001867664, 0.001055234, 0.0006958539, 
    0.0006063593, 0.0005423889, 0.0005784211, 0.000569283, 0.0004351789, 
    0.0003553139, 0.0003244683, 0.0003446025, 0.0004239017, 0.0004339685,
  0.001618509, 0.001604786, 0.001487517, 0.001415475, 0.001253158, 
    0.001193861, 0.001180086, 0.001100894, 0.001047695, 0.001023205, 
    0.001083143, 0.001128339, 0.001056614, 0.001012707, 0.0008568307,
  0.001658055, 0.00160139, 0.001509568, 0.001333365, 0.001175835, 
    0.001166566, 0.001216133, 0.001123305, 0.001081953, 0.001085454, 
    0.001007585, 0.0009468025, 0.0008918149, 0.0008002875, 0.0007032616,
  0.001838436, 0.00165808, 0.001497888, 0.00136668, 0.00124948, 0.001016094, 
    0.001167057, 0.001202184, 0.001123833, 0.001110341, 0.001035319, 
    0.0009434809, 0.0008657224, 0.00078679, 0.0007147373,
  0.001929171, 0.00204947, 0.001957939, 0.001631191, 0.001352071, 
    0.001311686, 0.0009577252, 0.001144065, 0.001214845, 0.00118412, 
    0.001111364, 0.001011891, 0.0008989797, 0.0007875301, 0.0006976629,
  0.001883972, 0.002029584, 0.002137972, 0.001921485, 0.001491762, 
    0.001446876, 0.001302398, 0.0009985052, 0.001013209, 0.001137557, 
    0.001205806, 0.001084109, 0.0009207477, 0.00079284, 0.0006902132,
  0.001836425, 0.001944036, 0.002086684, 0.002086374, 0.001818502, 
    0.001552898, 0.001466429, 0.001277108, 0.001162065, 0.0009539077, 
    0.0008674543, 0.0008892867, 0.0007827507, 0.0006787395, 0.0005834097,
  0.00185273, 0.00186792, 0.002016623, 0.002134689, 0.002111814, 0.001834795, 
    0.00162038, 0.00138005, 0.001124318, 0.0008811448, 0.0007811615, 
    0.0007001345, 0.0006341015, 0.0005194715, 0.0004560074,
  0.001867293, 0.001860435, 0.001973574, 0.002110713, 0.002160166, 
    0.002017752, 0.001716639, 0.001392132, 0.001084377, 0.0007876011, 
    0.0006733639, 0.0005670505, 0.0004722803, 0.0004192212, 0.000396189,
  0.001987596, 0.001994076, 0.002039595, 0.002124196, 0.002283034, 
    0.001992721, 0.001683063, 0.001230333, 0.0009435075, 0.0007232427, 
    0.0005411694, 0.0004322024, 0.0003754695, 0.0003438595, 0.0003502296,
  0.002253911, 0.0025854, 0.002681162, 0.002279871, 0.00198514, 0.001536062, 
    0.001170157, 0.0008811866, 0.000652167, 0.0004423143, 0.0003101931, 
    0.0002860843, 0.0002848745, 0.0003115495, 0.0003538645,
  0.001562689, 0.001701102, 0.001711679, 0.001679516, 0.001616721, 
    0.001551795, 0.001514963, 0.00150219, 0.001364917, 0.001112548, 
    0.001078314, 0.001055852, 0.000893097, 0.0008973491, 0.0008493119,
  0.001910079, 0.001933343, 0.001885808, 0.001760861, 0.001601021, 
    0.001536433, 0.001480716, 0.001419628, 0.001345228, 0.001220963, 
    0.001145974, 0.001132723, 0.001015381, 0.0008630692, 0.0008304362,
  0.002113204, 0.002000569, 0.001886614, 0.001832683, 0.001710236, 
    0.001391507, 0.001455267, 0.001383555, 0.001345525, 0.001227694, 
    0.001164962, 0.001114347, 0.001024917, 0.000934526, 0.0009010791,
  0.002049562, 0.001899793, 0.001958428, 0.001913768, 0.001770066, 
    0.001598771, 0.001158437, 0.001262758, 0.001256026, 0.001195564, 
    0.001156474, 0.001116408, 0.001053469, 0.0009584053, 0.0009443772,
  0.00188011, 0.001815823, 0.001924326, 0.001831242, 0.001647601, 
    0.001638331, 0.001377166, 0.001007052, 0.0009724052, 0.001101474, 
    0.00122572, 0.001183374, 0.001087241, 0.00100804, 0.0009942539,
  0.001857204, 0.001764979, 0.001880895, 0.001844025, 0.00158372, 0.0015457, 
    0.001440487, 0.001201064, 0.001044267, 0.0009477453, 0.001025646, 
    0.001101812, 0.001051643, 0.001037343, 0.001018805,
  0.001867739, 0.001859515, 0.001885935, 0.001879117, 0.001700384, 
    0.001467458, 0.001325895, 0.001155028, 0.001017319, 0.0009706746, 
    0.0009599163, 0.0009267731, 0.0009541257, 0.0009285128, 0.0009106674,
  0.001993923, 0.001945191, 0.001960201, 0.00193593, 0.001816634, 
    0.001421507, 0.001283425, 0.001136089, 0.001005227, 0.0009202053, 
    0.0008913222, 0.00091406, 0.0008220714, 0.0006740401, 0.0006283196,
  0.002167981, 0.002081863, 0.002021398, 0.001902972, 0.001726331, 
    0.001442484, 0.001301582, 0.001134009, 0.0009526518, 0.0007472433, 
    0.000549793, 0.000482239, 0.0004282456, 0.0003659039, 0.0003244541,
  0.002150861, 0.002127594, 0.001842553, 0.001456689, 0.00125909, 
    0.001055366, 0.0009048677, 0.0007629891, 0.0005504694, 0.0003646627, 
    0.0002880031, 0.0002554972, 0.0002509417, 0.0002574939, 0.0002877158,
  0.00200915, 0.002070203, 0.002150425, 0.002089427, 0.001948756, 
    0.001850852, 0.001864424, 0.001853494, 0.001773389, 0.001570214, 
    0.001448747, 0.001437854, 0.00130942, 0.001205854, 0.001151374,
  0.002211966, 0.002221346, 0.002164452, 0.001979098, 0.001861907, 
    0.001836016, 0.001822261, 0.001730084, 0.001804243, 0.001692819, 
    0.001548458, 0.001499953, 0.001413906, 0.001172013, 0.001023164,
  0.002122905, 0.002030504, 0.001885233, 0.001771245, 0.001733249, 
    0.001589667, 0.001722582, 0.001711139, 0.001657532, 0.001636984, 
    0.001503404, 0.001373847, 0.001295426, 0.001195336, 0.001088483,
  0.001862706, 0.001811649, 0.001753754, 0.001624199, 0.001613721, 
    0.001679997, 0.001356046, 0.001519093, 0.001440101, 0.001403628, 
    0.001317985, 0.001260525, 0.001210046, 0.001217222, 0.001110154,
  0.001803054, 0.001732609, 0.001671449, 0.001462049, 0.001388535, 
    0.001492345, 0.001503535, 0.001047958, 0.00107993, 0.001254798, 
    0.001281883, 0.001238718, 0.001170778, 0.001131919, 0.001099919,
  0.001744068, 0.001654921, 0.001550041, 0.001376143, 0.001193166, 
    0.001142047, 0.001243343, 0.001241482, 0.001181405, 0.001176075, 
    0.001182992, 0.001195337, 0.001133702, 0.001098558, 0.001026196,
  0.001689053, 0.001594314, 0.00149514, 0.00134683, 0.001172892, 
    0.0008746026, 0.0008825044, 0.0009400795, 0.0009772929, 0.001000851, 
    0.0009982605, 0.0009904896, 0.0009789701, 0.0009451128, 0.0009304158,
  0.00162223, 0.001518408, 0.001405494, 0.00132454, 0.001168985, 
    0.0007509262, 0.0007113471, 0.0006682614, 0.000665142, 0.0006477133, 
    0.0006426886, 0.0006454756, 0.0006361104, 0.0006383155, 0.0006425383,
  0.001589321, 0.001482243, 0.001303271, 0.001035923, 0.0006988005, 
    0.0006260394, 0.0005932684, 0.0005505145, 0.0004738886, 0.0004054906, 
    0.0003617326, 0.0003778269, 0.0003850802, 0.0003815368, 0.0003646968,
  0.001595886, 0.001442637, 0.001147851, 0.000664936, 0.0005134764, 
    0.000492795, 0.0005416108, 0.0005757877, 0.0004383535, 0.0003248964, 
    0.0002894695, 0.0003040963, 0.0003132532, 0.0003236656, 0.0003222699,
  0.001616202, 0.001571653, 0.001619623, 0.001453465, 0.001207544, 
    0.001113968, 0.001163232, 0.00115739, 0.001227333, 0.001307968, 
    0.001411922, 0.001513218, 0.001547079, 0.001528378, 0.001483219,
  0.001755969, 0.001667908, 0.001590975, 0.001414354, 0.001082351, 
    0.001014156, 0.001015925, 0.0009976722, 0.001069352, 0.001204596, 
    0.001378511, 0.001514595, 0.001574023, 0.001446622, 0.001397114,
  0.001838899, 0.001789445, 0.001588689, 0.001377493, 0.001049414, 
    0.0007766407, 0.0008550165, 0.0008791732, 0.0009590176, 0.001091756, 
    0.001252769, 0.001328092, 0.001386823, 0.00140453, 0.001344504,
  0.001710678, 0.001682668, 0.001695778, 0.001531525, 0.001145949, 
    0.0008886408, 0.0005974848, 0.0006934214, 0.0007763283, 0.0008788479, 
    0.0009959341, 0.001064723, 0.001136139, 0.001191114, 0.001243792,
  0.001849945, 0.001753894, 0.001701026, 0.001557517, 0.001170053, 
    0.0008696842, 0.000776166, 0.0004406858, 0.0005404717, 0.0007295326, 
    0.0008143427, 0.0008397487, 0.0008318122, 0.0008763185, 0.0009823535,
  0.00214639, 0.001985301, 0.001853147, 0.001644715, 0.001147585, 
    0.0007461557, 0.0006716647, 0.0006025126, 0.0005841639, 0.0005911464, 
    0.0005930309, 0.0006472765, 0.0006659396, 0.0007031218, 0.0007563367,
  0.002425057, 0.002294166, 0.002100929, 0.001808033, 0.00108677, 
    0.0006513441, 0.0005588297, 0.0005388401, 0.0005294294, 0.0005174655, 
    0.0004967056, 0.0004974261, 0.0005094977, 0.0005453097, 0.0006028753,
  0.002513856, 0.002479003, 0.002397169, 0.001732689, 0.001018104, 
    0.0006072327, 0.000506134, 0.0004758833, 0.0004722553, 0.0004442276, 
    0.0004180599, 0.0004391308, 0.000413207, 0.0004423693, 0.0004680846,
  0.002530378, 0.002445946, 0.002273294, 0.001485265, 0.0007753439, 
    0.0005946782, 0.0005316663, 0.0005233305, 0.0004660634, 0.0004085689, 
    0.0003758151, 0.0003838979, 0.0003614342, 0.0003768636, 0.0004076173,
  0.002389014, 0.002236757, 0.001928914, 0.001066398, 0.0006185776, 
    0.0005253216, 0.0005125692, 0.0005347712, 0.0004479248, 0.0003669451, 
    0.0003318708, 0.0003337054, 0.0003159243, 0.0003321831, 0.000355861,
  0.001855302, 0.001854481, 0.001732974, 0.001718594, 0.001550595, 
    0.001544665, 0.001665865, 0.001427633, 0.001231246, 0.001069057, 
    0.0009526201, 0.0008787776, 0.0007493514, 0.00068748, 0.0006553045,
  0.001680919, 0.001697893, 0.00171695, 0.001649395, 0.001526028, 
    0.001550788, 0.001486561, 0.001331054, 0.001183697, 0.001013698, 
    0.0009222465, 0.0008972461, 0.000776857, 0.0006229254, 0.0005537752,
  0.002134283, 0.001950938, 0.001649024, 0.00158552, 0.001386198, 0.00119833, 
    0.001303293, 0.001223762, 0.001060871, 0.001060044, 0.001036161, 
    0.0009214581, 0.0008296453, 0.0006990618, 0.000590514,
  0.001999314, 0.002090076, 0.002220287, 0.001948074, 0.00152587, 
    0.001427013, 0.001168743, 0.001202725, 0.001173876, 0.001005336, 
    0.0008652417, 0.0007437536, 0.0006798116, 0.0006172088, 0.000535182,
  0.002092271, 0.002035652, 0.002049127, 0.002060506, 0.001799362, 
    0.001873001, 0.001717727, 0.0008550609, 0.0005249445, 0.0006026519, 
    0.0006053452, 0.0005514427, 0.000525881, 0.0005036715, 0.0004909175,
  0.002475859, 0.002306752, 0.002081894, 0.001734473, 0.001422671, 
    0.001189084, 0.0008856113, 0.0006751373, 0.0005182089, 0.0004201543, 
    0.0003918975, 0.0004201351, 0.0004173164, 0.0004109128, 0.0004063049,
  0.002285682, 0.002094972, 0.001733978, 0.00126984, 0.0008836339, 
    0.000627514, 0.0005665803, 0.0004909714, 0.0004201322, 0.0003943295, 
    0.0003796548, 0.0003665536, 0.0003602002, 0.0003387986, 0.000337124,
  0.001937518, 0.001729091, 0.001492241, 0.001198793, 0.0008635374, 
    0.0005275501, 0.0004606892, 0.0004047815, 0.0003865637, 0.0003692772, 
    0.0003374303, 0.0003282063, 0.0002980219, 0.0003010376, 0.0003213861,
  0.001614163, 0.001448871, 0.001235784, 0.0009362221, 0.0005476989, 
    0.0004611766, 0.0004209042, 0.0004021406, 0.0003789979, 0.0003470253, 
    0.0003092822, 0.0002832384, 0.0002698074, 0.0002629448, 0.0002885758,
  0.0013947, 0.001227537, 0.0009444089, 0.0005306888, 0.0004514824, 
    0.0004293965, 0.0004155081, 0.0004220959, 0.0003815812, 0.0003086889, 
    0.0002878938, 0.0002783665, 0.0002583197, 0.0002496631, 0.0002646917,
  0.001932382, 0.001915655, 0.001834995, 0.001847892, 0.002122976, 
    0.002407313, 0.002506752, 0.002281505, 0.002095731, 0.001996711, 
    0.001885997, 0.001774678, 0.001625026, 0.001501591, 0.001325781,
  0.001972555, 0.001860923, 0.001787912, 0.001757113, 0.001711429, 
    0.001791282, 0.001958616, 0.001970024, 0.001920601, 0.00186793, 
    0.001735943, 0.001734376, 0.001588343, 0.001367504, 0.001228755,
  0.002096205, 0.001878737, 0.001733198, 0.001629255, 0.00148463, 
    0.001296064, 0.00140976, 0.00148897, 0.00156546, 0.001683839, 
    0.001693445, 0.001593295, 0.001486867, 0.001398088, 0.001254077,
  0.001972758, 0.002007284, 0.001944187, 0.001707951, 0.001427422, 
    0.001351848, 0.001211518, 0.001234843, 0.001243384, 0.00124668, 
    0.001196343, 0.001064278, 0.001009215, 0.0009128819, 0.0007688146,
  0.001983418, 0.001955418, 0.001917113, 0.001703513, 0.001395912, 
    0.001475684, 0.001358256, 0.0008129185, 0.0006479567, 0.0007083039, 
    0.0007568595, 0.0006577411, 0.0006191734, 0.0005738689, 0.0005244827,
  0.001796468, 0.001647751, 0.001485174, 0.001049733, 0.0008957943, 
    0.0008718789, 0.001000045, 0.0008812759, 0.0005933025, 0.0004803043, 
    0.0004456273, 0.0004759349, 0.0004415752, 0.000419398, 0.0003889808,
  0.001394043, 0.001294516, 0.001181058, 0.000770357, 0.0006970257, 
    0.0006086418, 0.0005941417, 0.0005484516, 0.000464637, 0.0004569755, 
    0.0004226055, 0.0003888772, 0.0003883868, 0.0003793274, 0.0003650816,
  0.001297012, 0.001205849, 0.001111315, 0.001003079, 0.0007982653, 
    0.0005397465, 0.000466812, 0.0004588169, 0.0004628115, 0.0004417224, 
    0.0004107972, 0.0003958303, 0.0003823647, 0.0003800735, 0.0003799452,
  0.001452232, 0.0013247, 0.001215851, 0.001061784, 0.0008992367, 
    0.0007304939, 0.0006251661, 0.0005717028, 0.0005406583, 0.0005349024, 
    0.0005256911, 0.0004878241, 0.0004654549, 0.0004462535, 0.0004191874,
  0.001676923, 0.001581049, 0.001422356, 0.001179871, 0.0009518731, 
    0.0008107287, 0.0006846017, 0.0006490113, 0.000647894, 0.0006303781, 
    0.0006723742, 0.0006308866, 0.0005710219, 0.0005657126, 0.0005358551,
  0.001501272, 0.001468065, 0.001520379, 0.001691663, 0.002348869, 
    0.002632697, 0.002823007, 0.002610797, 0.002766546, 0.002586555, 
    0.002484446, 0.002471447, 0.002397998, 0.002252834, 0.002188146,
  0.001610277, 0.001484912, 0.001498085, 0.001559053, 0.001798494, 
    0.002387932, 0.002719926, 0.002715463, 0.002756947, 0.002603479, 
    0.002496376, 0.002448273, 0.002334193, 0.002038314, 0.001953908,
  0.001628826, 0.001561156, 0.001528754, 0.001493815, 0.00155266, 
    0.001672618, 0.002357549, 0.002665851, 0.002711715, 0.002609442, 
    0.002509073, 0.002381782, 0.002248758, 0.002077942, 0.001798557,
  0.001620253, 0.001639907, 0.001669426, 0.001395267, 0.001434594, 
    0.001675793, 0.001785884, 0.002200027, 0.002413416, 0.002448658, 
    0.002420413, 0.002274133, 0.002150404, 0.001940036, 0.001641816,
  0.001577991, 0.001549921, 0.001644168, 0.001265737, 0.001207611, 
    0.001411592, 0.001707601, 0.001525521, 0.001486324, 0.002063721, 
    0.002193887, 0.002038965, 0.001937664, 0.001776971, 0.001555255,
  0.001584949, 0.001503318, 0.001545821, 0.001149422, 0.001055737, 
    0.001099864, 0.001273808, 0.00150531, 0.001536054, 0.001706961, 
    0.001772494, 0.001725873, 0.001670488, 0.00152999, 0.001320002,
  0.00171584, 0.001664452, 0.001577746, 0.001229304, 0.001013318, 
    0.0009102435, 0.0009763828, 0.001087834, 0.001312922, 0.001421757, 
    0.001406677, 0.001399077, 0.001368997, 0.001250788, 0.001046517,
  0.002048686, 0.001994323, 0.001941269, 0.001900124, 0.001264256, 
    0.000736066, 0.0007457, 0.0007848819, 0.000863355, 0.001040953, 
    0.001127656, 0.001114106, 0.001076723, 0.0009844197, 0.0008363031,
  0.002484252, 0.002380886, 0.002300918, 0.002208272, 0.001711428, 
    0.00092887, 0.0006938152, 0.0006595371, 0.0006984565, 0.000762736, 
    0.0008478194, 0.0008732556, 0.0008206152, 0.0007236667, 0.000622944,
  0.002909424, 0.002874445, 0.002817933, 0.002566969, 0.002232545, 
    0.001281854, 0.0007318272, 0.0006059899, 0.0005954569, 0.0005959725, 
    0.000701244, 0.00068583, 0.0006568912, 0.0006265602, 0.0005880228,
  0.001289906, 0.001255658, 0.001251492, 0.001595095, 0.001830421, 
    0.001962928, 0.00189761, 0.001626033, 0.001552858, 0.00182938, 
    0.001697461, 0.001985888, 0.002057586, 0.002054602, 0.001951292,
  0.001573623, 0.001485245, 0.001520146, 0.001813475, 0.001818821, 
    0.001914305, 0.001909669, 0.001558476, 0.001956345, 0.001884834, 
    0.001907609, 0.00216096, 0.002321516, 0.002235024, 0.001930478,
  0.002224303, 0.002054595, 0.001912797, 0.001919986, 0.001746428, 
    0.001944972, 0.002199905, 0.00181204, 0.002386512, 0.00240952, 
    0.002330519, 0.002296508, 0.002452688, 0.002387648, 0.002031932,
  0.00237501, 0.002272707, 0.002068495, 0.002058427, 0.001771274, 
    0.002045379, 0.001994814, 0.002091449, 0.002491836, 0.002538375, 
    0.002483061, 0.002347054, 0.002342816, 0.002126389, 0.001769356,
  0.002543003, 0.002380069, 0.002156141, 0.001943914, 0.001697778, 
    0.00190243, 0.00252789, 0.002225748, 0.002199574, 0.00245976, 
    0.002503055, 0.002265293, 0.002194421, 0.001873813, 0.001688511,
  0.002477386, 0.002349134, 0.002226893, 0.002000301, 0.001750335, 
    0.001695185, 0.002058839, 0.00231239, 0.002321468, 0.002363299, 
    0.002329949, 0.002278249, 0.001987127, 0.00160413, 0.00145682,
  0.002356744, 0.002303641, 0.002230599, 0.002212103, 0.001938253, 
    0.001559828, 0.001893553, 0.002145078, 0.002315389, 0.002380318, 
    0.002246492, 0.002182683, 0.001860562, 0.001547213, 0.001259693,
  0.002225541, 0.002213982, 0.002226747, 0.002294888, 0.002231118, 
    0.001370148, 0.001464265, 0.001736484, 0.002081525, 0.002231043, 
    0.002163038, 0.002115139, 0.001811119, 0.001433294, 0.001074302,
  0.001953676, 0.002037951, 0.002178127, 0.002396503, 0.002405486, 
    0.001702303, 0.001251206, 0.001596122, 0.001731258, 0.001955174, 
    0.002131807, 0.002056559, 0.001739202, 0.001269499, 0.0009575327,
  0.001474228, 0.001493304, 0.001566984, 0.001827142, 0.002434531, 
    0.001940074, 0.001269059, 0.001266229, 0.001484436, 0.001684483, 
    0.001950309, 0.001974977, 0.001644497, 0.001182686, 0.0009947596,
  0.001469133, 0.00147512, 0.001416744, 0.001427157, 0.001574161, 
    0.001395431, 0.001538369, 0.00154228, 0.00150291, 0.001449893, 
    0.001345726, 0.001523169, 0.001608673, 0.001590411, 0.00145265,
  0.001737019, 0.001648888, 0.00157771, 0.001523532, 0.001622669, 
    0.001335237, 0.001444849, 0.001431347, 0.001479243, 0.001247412, 
    0.001311454, 0.001571891, 0.001640227, 0.001597754, 0.00123431,
  0.001651511, 0.001746121, 0.001593882, 0.001557365, 0.001598157, 
    0.001386722, 0.001254685, 0.001159653, 0.00153002, 0.001463314, 
    0.001668728, 0.001792178, 0.001797274, 0.001743416, 0.001592195,
  0.001483597, 0.001595821, 0.001776655, 0.001796652, 0.001746238, 
    0.001743673, 0.001405112, 0.001314959, 0.001763823, 0.001821912, 
    0.001514651, 0.001637785, 0.001737708, 0.00186529, 0.001767373,
  0.001383469, 0.001404441, 0.0015902, 0.001640895, 0.001706095, 0.001877217, 
    0.001988612, 0.001676593, 0.00135326, 0.001593197, 0.001695068, 
    0.001778644, 0.001812488, 0.001854177, 0.00184993,
  0.00133017, 0.001272746, 0.001364724, 0.001528029, 0.00167064, 0.001887232, 
    0.002006815, 0.001887602, 0.001788595, 0.001911115, 0.00158323, 
    0.00171256, 0.001845838, 0.001920575, 0.001669098,
  0.001278256, 0.001210683, 0.001270369, 0.001393377, 0.001627917, 
    0.001757209, 0.001942873, 0.001589509, 0.001938684, 0.002037727, 
    0.00177111, 0.001751644, 0.001881697, 0.001673229, 0.001047367,
  0.001220783, 0.001194826, 0.00126751, 0.001423284, 0.001809582, 
    0.001630377, 0.001490707, 0.001752826, 0.001852543, 0.001961508, 
    0.001700129, 0.001747459, 0.001567974, 0.0009734753, 0.0005819513,
  0.001164704, 0.001189338, 0.001258757, 0.001214982, 0.001780295, 
    0.001894406, 0.001532192, 0.001649875, 0.001898079, 0.001810114, 
    0.001654196, 0.001548006, 0.0009925236, 0.0006347705, 0.0005317213,
  0.001054384, 0.001050233, 0.0009150985, 0.0008040927, 0.001570102, 
    0.001965982, 0.001687334, 0.001863836, 0.001671803, 0.001646563, 
    0.001486935, 0.001140509, 0.0007454238, 0.000621621, 0.0005720523,
  0.001366898, 0.001223002, 0.001072734, 0.001069749, 0.001285273, 
    0.001426008, 0.001262013, 0.001337208, 0.001395087, 0.001368782, 
    0.001421681, 0.001706009, 0.001556527, 0.001432359, 0.001362663,
  0.001595916, 0.001284278, 0.001158499, 0.001111875, 0.001235791, 
    0.001340474, 0.001408947, 0.001340795, 0.00145978, 0.001396867, 
    0.001316084, 0.001501994, 0.001506061, 0.001265824, 0.00110189,
  0.001622151, 0.001497368, 0.001295491, 0.00118165, 0.001141067, 
    0.001326708, 0.001299751, 0.001233293, 0.00119718, 0.001267695, 
    0.001364939, 0.001420215, 0.001397821, 0.001305944, 0.0009463158,
  0.001662177, 0.001620048, 0.001495635, 0.001367477, 0.001299495, 
    0.001485891, 0.001333454, 0.00117502, 0.001324963, 0.001441567, 
    0.001357645, 0.00134548, 0.00129403, 0.001137329, 0.0009040036,
  0.001690353, 0.001667194, 0.00164192, 0.001589173, 0.001509267, 
    0.001596516, 0.001742253, 0.0009969342, 0.001100532, 0.001243537, 
    0.001374345, 0.001339017, 0.001205726, 0.001057466, 0.0008863715,
  0.001683862, 0.001705018, 0.00173247, 0.001793041, 0.001778983, 
    0.001688812, 0.001776498, 0.00169512, 0.001418158, 0.00138699, 
    0.00127061, 0.001241017, 0.001105423, 0.0009175675, 0.000765547,
  0.001684148, 0.001730607, 0.001805892, 0.001872835, 0.001930677, 
    0.001609289, 0.001618392, 0.001517586, 0.001456057, 0.001366385, 
    0.001269602, 0.001139453, 0.0009057822, 0.0006810474, 0.0005831618,
  0.001641391, 0.001715352, 0.001798058, 0.00189769, 0.001983923, 
    0.001586007, 0.001417987, 0.001424843, 0.00129125, 0.001278426, 
    0.001102422, 0.0008350561, 0.0006123064, 0.000511993, 0.0004757053,
  0.001477172, 0.001518802, 0.001542234, 0.001442519, 0.00161681, 
    0.001629639, 0.001340487, 0.001321671, 0.001339649, 0.001062094, 
    0.0007937021, 0.0005978481, 0.0005054623, 0.0004879786, 0.0004895558,
  0.001250486, 0.001173395, 0.001036173, 0.000968173, 0.001238186, 
    0.001424755, 0.001389673, 0.001278979, 0.001158521, 0.0008588617, 
    0.0006194782, 0.0005086628, 0.0004917104, 0.0004990507, 0.0005351671,
  0.001701227, 0.001480503, 0.001329678, 0.001411367, 0.001322328, 
    0.001113446, 0.001037366, 0.001101859, 0.001194715, 0.00113643, 
    0.001078901, 0.001145563, 0.00105594, 0.0009325731, 0.0008364317,
  0.001997185, 0.001620613, 0.001509209, 0.001443892, 0.00125568, 
    0.0009745678, 0.0009884943, 0.001025568, 0.001021317, 0.001057311, 
    0.0009923457, 0.001086506, 0.001068076, 0.0008772452, 0.0008228284,
  0.00204276, 0.001916123, 0.0015966, 0.00151104, 0.001190495, 0.0009941995, 
    0.0008588873, 0.0009291168, 0.0008892458, 0.0009184621, 0.0009088746, 
    0.0009862023, 0.001042324, 0.00101074, 0.00087924,
  0.002000821, 0.0018915, 0.001728661, 0.001494418, 0.001281166, 0.001138585, 
    0.000737514, 0.0007679374, 0.0008050974, 0.0007943293, 0.000768607, 
    0.0008122115, 0.0009104088, 0.0009581269, 0.0009229483,
  0.001992926, 0.001838807, 0.001725049, 0.001454243, 0.001245386, 0.0011631, 
    0.001055663, 0.0006469615, 0.0006471236, 0.0007046797, 0.0006871711, 
    0.0006813119, 0.0007382489, 0.0007943358, 0.000855657,
  0.001967907, 0.001848037, 0.001706345, 0.001602102, 0.001354051, 
    0.001057793, 0.0009927112, 0.000916268, 0.0007500554, 0.0007131583, 
    0.00061602, 0.0006269886, 0.0006174822, 0.0006515139, 0.000725576,
  0.002030521, 0.001836901, 0.00178049, 0.001705862, 0.001479307, 
    0.0009688846, 0.0008003513, 0.0007472837, 0.0007008163, 0.000643192, 
    0.0005874408, 0.0005699864, 0.0005660331, 0.0005612036, 0.0005916686,
  0.002086368, 0.001845943, 0.001771703, 0.001796788, 0.001657562, 
    0.001041603, 0.0007386934, 0.0006247454, 0.0005628231, 0.000529632, 
    0.0004976849, 0.000514213, 0.0005204238, 0.0005310808, 0.000532061,
  0.002171193, 0.001870255, 0.001712812, 0.00144756, 0.001458305, 
    0.001363915, 0.0007914605, 0.0006184523, 0.000510825, 0.0004583677, 
    0.0004469074, 0.000468133, 0.0004757746, 0.0005093632, 0.0005419841,
  0.002306292, 0.001893607, 0.001544019, 0.001262419, 0.001212088, 
    0.001178715, 0.0008875637, 0.0006788526, 0.0005187768, 0.0004200174, 
    0.0004202041, 0.0004328925, 0.0004356935, 0.0004724289, 0.0005291961,
  0.002426483, 0.002184019, 0.001840585, 0.001756373, 0.001506625, 
    0.001160634, 0.0009979656, 0.0008786447, 0.0008275257, 0.0007846206, 
    0.0007819207, 0.0008875486, 0.0008174957, 0.0008072017, 0.0008634331,
  0.002813528, 0.00258749, 0.002201971, 0.001951502, 0.001679039, 
    0.001338503, 0.001141654, 0.0009908675, 0.0008975088, 0.0008664833, 
    0.0007694621, 0.0008644203, 0.0009052259, 0.0007156596, 0.0006721846,
  0.003087261, 0.002948059, 0.002559418, 0.002134769, 0.001702018, 
    0.001277189, 0.001145488, 0.0009845475, 0.0009060364, 0.000853295, 
    0.0007971501, 0.000812948, 0.0008956388, 0.000891675, 0.0007106186,
  0.003352122, 0.002988839, 0.002734477, 0.002282422, 0.001837267, 
    0.001469068, 0.001054167, 0.0009299014, 0.0008752279, 0.0008241546, 
    0.0007822719, 0.0007442016, 0.0008018165, 0.0008566714, 0.0008019963,
  0.003559967, 0.003024275, 0.002677623, 0.002268113, 0.001841787, 
    0.001476103, 0.001246002, 0.0007968053, 0.0006848703, 0.0007767662, 
    0.0007526199, 0.0007288347, 0.0007075435, 0.0007615671, 0.0008236152,
  0.003593361, 0.003052925, 0.002561921, 0.002210115, 0.001837872, 
    0.001475038, 0.001230718, 0.001133239, 0.001016297, 0.0009534345, 
    0.0007805986, 0.0007404403, 0.0006667647, 0.000667126, 0.0007245081,
  0.003528399, 0.002996152, 0.00245715, 0.00207941, 0.001748664, 0.001429942, 
    0.001218504, 0.001126906, 0.001056712, 0.0009651357, 0.0008343706, 
    0.0007577246, 0.0006647861, 0.0006149907, 0.0006559378,
  0.003272598, 0.002787567, 0.002292146, 0.001950787, 0.001652138, 
    0.001376276, 0.001195378, 0.001150362, 0.00108424, 0.001009643, 
    0.0009241706, 0.0007962871, 0.0006532774, 0.0005717099, 0.0005731959,
  0.002961244, 0.002499798, 0.002091164, 0.001669614, 0.001366597, 
    0.001194276, 0.00115329, 0.001192812, 0.001145913, 0.001069315, 
    0.0009738471, 0.0008267818, 0.0006480992, 0.0005664915, 0.0005642948,
  0.002588017, 0.002118487, 0.001656611, 0.001331012, 0.001109571, 
    0.0009948834, 0.001041744, 0.001200572, 0.001209131, 0.001088001, 
    0.0009785679, 0.0007978298, 0.0006202321, 0.0005579722, 0.0005643357,
  0.002381458, 0.002311113, 0.002025817, 0.001674186, 0.001397396, 
    0.001198036, 0.00115109, 0.001075659, 0.001022958, 0.0009479533, 
    0.0009206752, 0.0008544806, 0.0008302217, 0.00088703, 0.0008796356,
  0.002433849, 0.002189519, 0.001837226, 0.001427702, 0.001179524, 
    0.00099627, 0.0009881257, 0.0009592862, 0.000939671, 0.0009577281, 
    0.0008294196, 0.0008315044, 0.0008625963, 0.0008168729, 0.0008040164,
  0.002313565, 0.002049342, 0.001751827, 0.001308597, 0.001079469, 
    0.000906371, 0.0009240297, 0.0009409822, 0.0009138558, 0.0008542598, 
    0.0008321815, 0.0008246762, 0.0008501893, 0.0009144586, 0.0009322269,
  0.002148106, 0.001978993, 0.001720666, 0.001290945, 0.001063624, 
    0.0009434544, 0.0008390659, 0.0008963691, 0.00091502, 0.0009201762, 
    0.0008315232, 0.0008668842, 0.0008710459, 0.0009895741, 0.0009926412,
  0.002053336, 0.001878101, 0.00161551, 0.00120264, 0.0010418, 0.0009806207, 
    0.0009732083, 0.0008019479, 0.0008001304, 0.0009300669, 0.0008523688, 
    0.0008771872, 0.0009845401, 0.001010324, 0.0009846435,
  0.001998852, 0.001739231, 0.001483983, 0.001159166, 0.001031733, 
    0.0009993664, 0.001030801, 0.00105012, 0.001035453, 0.0009594786, 
    0.0007946916, 0.0008706744, 0.0009701864, 0.000985979, 0.0009612843,
  0.00202366, 0.001652123, 0.001475791, 0.001251077, 0.00103534, 
    0.0009450775, 0.001015663, 0.001057079, 0.001056952, 0.0009917065, 
    0.000864203, 0.0008662505, 0.0008943175, 0.0008750522, 0.0008353967,
  0.002187214, 0.001670753, 0.001465037, 0.001296831, 0.001067375, 
    0.0008850504, 0.0009409111, 0.0009973509, 0.0009886189, 0.0009664124, 
    0.0008463783, 0.0008507207, 0.0008097368, 0.000754579, 0.0007192733,
  0.002395898, 0.00178818, 0.001490186, 0.001040103, 0.0008926989, 
    0.0008304134, 0.0008794756, 0.000939025, 0.0009271708, 0.0008862674, 
    0.0008310952, 0.0007873147, 0.0007157063, 0.0006340183, 0.000580975,
  0.002500471, 0.00176265, 0.001303878, 0.0009665323, 0.0008685227, 
    0.0008005587, 0.0008029251, 0.0008999658, 0.0008502303, 0.0007340249, 
    0.0006664183, 0.0006656045, 0.0006041757, 0.0005829994, 0.0005629144,
  0.001807843, 0.00171226, 0.001494837, 0.00131263, 0.001256056, 0.001031374, 
    0.0009519373, 0.0009292764, 0.0008751422, 0.0008195394, 0.0009075223, 
    0.0007721221, 0.0006467634, 0.0006735134, 0.0006650802,
  0.002266464, 0.002076031, 0.001838311, 0.001542399, 0.001384671, 
    0.001122819, 0.001080238, 0.001004251, 0.0009311665, 0.0008983368, 
    0.0007891905, 0.000929145, 0.0009195214, 0.0007498228, 0.0006368427,
  0.002646487, 0.002457574, 0.002283731, 0.00193512, 0.001565538, 
    0.001179065, 0.001156416, 0.001080988, 0.0009843427, 0.0008943279, 
    0.0008632608, 0.000912889, 0.000951436, 0.0009559045, 0.0008162921,
  0.002966271, 0.002775615, 0.002631192, 0.002332673, 0.001972545, 
    0.001528078, 0.001147976, 0.001062424, 0.001039017, 0.0009403707, 
    0.0008446135, 0.0009097848, 0.0009357763, 0.0009585242, 0.0008994003,
  0.003336979, 0.003064611, 0.00292443, 0.00262837, 0.002311978, 0.001906152, 
    0.001435492, 0.000948988, 0.0008718135, 0.0009436118, 0.0008349803, 
    0.0007965808, 0.0008562281, 0.000895219, 0.0009248104,
  0.003730808, 0.003463379, 0.003164757, 0.002909397, 0.002619534, 
    0.002283076, 0.001838535, 0.001392983, 0.001148205, 0.0009625413, 
    0.0007863138, 0.0007294673, 0.0007140276, 0.0007539876, 0.000816178,
  0.004050678, 0.003808398, 0.003456576, 0.003122356, 0.002848433, 
    0.002519388, 0.002163731, 0.001785705, 0.001430624, 0.001099593, 
    0.0008437177, 0.0007288761, 0.0006585187, 0.000638188, 0.0006701946,
  0.004109637, 0.003937975, 0.003633127, 0.003314558, 0.003084707, 
    0.002762973, 0.002388754, 0.002066372, 0.001716985, 0.001327983, 
    0.0009201385, 0.0007219902, 0.0006357325, 0.0005859432, 0.0005937112,
  0.003981696, 0.003823163, 0.003696515, 0.003472788, 0.003238712, 
    0.002934335, 0.002611575, 0.00230042, 0.001965035, 0.00152579, 
    0.001046378, 0.0007485606, 0.0006158624, 0.0005499253, 0.0005613679,
  0.00373886, 0.003627535, 0.00357647, 0.003513188, 0.003306511, 0.003061768, 
    0.002747466, 0.002453114, 0.002139477, 0.001551147, 0.001037008, 
    0.0007409096, 0.0005788876, 0.0005012218, 0.0005484797,
  0.003039782, 0.003143935, 0.003230782, 0.003309397, 0.00327543, 
    0.003125571, 0.002939464, 0.002630468, 0.00216753, 0.00155164, 
    0.001417281, 0.001234595, 0.0009784758, 0.000855198, 0.0007424272,
  0.003199445, 0.003243058, 0.003364628, 0.003496706, 0.003502046, 
    0.003356119, 0.003183174, 0.002976918, 0.002661617, 0.002031914, 
    0.001602686, 0.001399206, 0.001213913, 0.0009695702, 0.0007992818,
  0.003257701, 0.003198595, 0.003293161, 0.003496765, 0.003602256, 
    0.003354675, 0.003255255, 0.003190382, 0.002935613, 0.00259175, 
    0.002086842, 0.001681851, 0.00138562, 0.001176427, 0.001007372,
  0.003284625, 0.003211682, 0.003208604, 0.00333975, 0.003510488, 0.00353364, 
    0.003245892, 0.003091688, 0.002897322, 0.002686673, 0.002308662, 
    0.001939571, 0.001573287, 0.001301151, 0.001116066,
  0.003280476, 0.003079166, 0.003084642, 0.00318459, 0.003296315, 
    0.003347311, 0.003354593, 0.002884774, 0.002728093, 0.002815018, 
    0.002707321, 0.002301766, 0.001824667, 0.001418756, 0.001165836,
  0.003224189, 0.002988904, 0.002904675, 0.002986986, 0.003034901, 
    0.003034179, 0.003086317, 0.003079589, 0.00305838, 0.002994138, 
    0.00281614, 0.002515943, 0.002038478, 0.001539976, 0.001182709,
  0.003184866, 0.002908331, 0.002784241, 0.002733841, 0.002744976, 
    0.002731574, 0.002756186, 0.002798702, 0.002829911, 0.002843668, 
    0.002700465, 0.002428773, 0.001904947, 0.001424226, 0.001104573,
  0.003145357, 0.002866529, 0.002666241, 0.00250769, 0.002436653, 
    0.002424855, 0.002459604, 0.002478877, 0.002462708, 0.002542973, 
    0.002495658, 0.002133447, 0.001532157, 0.001140925, 0.000974283,
  0.003120731, 0.002827301, 0.00254629, 0.002205284, 0.002078995, 
    0.002129753, 0.002142668, 0.002157434, 0.002135629, 0.002123259, 
    0.00197217, 0.001494478, 0.001095014, 0.0008993087, 0.0007654267,
  0.003034913, 0.002717449, 0.002294231, 0.001986517, 0.00179137, 
    0.001768697, 0.001754026, 0.001794661, 0.001733598, 0.001529932, 
    0.001308289, 0.0009828423, 0.0008018341, 0.00069244, 0.0006107542,
  0.003290345, 0.003113189, 0.002970607, 0.002680254, 0.002324362, 
    0.002101452, 0.002057592, 0.002221119, 0.002630728, 0.002663226, 
    0.0026674, 0.002463366, 0.00178674, 0.001335128, 0.001063517,
  0.00348314, 0.003247089, 0.003012241, 0.002675972, 0.002159468, 
    0.001780881, 0.001753255, 0.001835693, 0.00203182, 0.002244659, 
    0.002351667, 0.002432908, 0.002122417, 0.001490719, 0.001174407,
  0.003554555, 0.003258161, 0.0030493, 0.002755369, 0.002150547, 0.001515765, 
    0.001560203, 0.001507989, 0.001597456, 0.001907233, 0.002127567, 
    0.002353149, 0.002378064, 0.001982576, 0.001447893,
  0.003837175, 0.003533461, 0.003242569, 0.002858867, 0.002281076, 
    0.001654004, 0.001205862, 0.001309693, 0.001308664, 0.00147665, 
    0.001775212, 0.002155951, 0.002375337, 0.002331305, 0.001771063,
  0.004085165, 0.003684605, 0.003392687, 0.002988678, 0.002413993, 
    0.001702443, 0.001332475, 0.0009503568, 0.001049253, 0.001258852, 
    0.001558299, 0.001944292, 0.002279773, 0.002432766, 0.002214478,
  0.004314541, 0.00391165, 0.003466369, 0.003095657, 0.002642644, 
    0.001973698, 0.001406595, 0.001148761, 0.001002583, 0.001098995, 
    0.001348876, 0.00177244, 0.002132548, 0.002412803, 0.002237656,
  0.004481693, 0.00413052, 0.003690057, 0.003237618, 0.00282846, 0.00226195, 
    0.00165627, 0.00122131, 0.001009272, 0.0009745385, 0.001126235, 
    0.001485941, 0.001860042, 0.001929643, 0.001649989,
  0.00451214, 0.004207946, 0.003817244, 0.003381487, 0.002995802, 
    0.002482658, 0.001906655, 0.001367443, 0.001021784, 0.0008540834, 
    0.0009394719, 0.0009755394, 0.001082, 0.001121029, 0.001046193,
  0.004439234, 0.004174737, 0.003850784, 0.003441398, 0.003039799, 
    0.002575943, 0.002085807, 0.001572386, 0.001140725, 0.000876486, 
    0.0007988815, 0.0008655968, 0.0008007089, 0.0007620329, 0.000704928,
  0.004150582, 0.003930656, 0.003640061, 0.00329745, 0.002966932, 
    0.002620379, 0.002231156, 0.001803442, 0.00135993, 0.0009393427, 
    0.0007237231, 0.000689726, 0.0006633883, 0.000625178, 0.0006256519,
  0.003876847, 0.003589261, 0.003548523, 0.003654256, 0.003546953, 
    0.002952364, 0.002587354, 0.001988325, 0.001467971, 0.001409209, 
    0.001162834, 0.001463207, 0.001815837, 0.00188757, 0.001741795,
  0.003775412, 0.00349999, 0.003435762, 0.003525936, 0.003549115, 
    0.003065452, 0.002652216, 0.00205089, 0.001472416, 0.001357997, 
    0.001365385, 0.001511023, 0.001616865, 0.001712518, 0.001586549,
  0.003796358, 0.003374635, 0.003292936, 0.003362597, 0.003551943, 
    0.003054237, 0.002658116, 0.002200262, 0.001650481, 0.001464233, 
    0.001334151, 0.001474194, 0.001574416, 0.001846434, 0.001853191,
  0.003973646, 0.003560633, 0.003314929, 0.003221027, 0.003414456, 
    0.003455916, 0.002721781, 0.002139705, 0.001785131, 0.001582342, 
    0.001406944, 0.001324306, 0.001471221, 0.001711217, 0.001998225,
  0.004050054, 0.003580577, 0.003247915, 0.003088603, 0.003182963, 
    0.003373086, 0.003158822, 0.002146025, 0.00176124, 0.001858051, 
    0.001647323, 0.001386287, 0.001481641, 0.001601248, 0.001900605,
  0.004105685, 0.003687938, 0.003112264, 0.002900378, 0.002952159, 
    0.003093388, 0.003128912, 0.002869149, 0.002427235, 0.001950287, 
    0.00162577, 0.00143305, 0.001332489, 0.001517763, 0.001801864,
  0.004103205, 0.003741449, 0.003104147, 0.002703728, 0.002669055, 
    0.002743158, 0.002857841, 0.00284454, 0.00260294, 0.002149198, 
    0.001717938, 0.001419231, 0.001260192, 0.001339593, 0.001578777,
  0.004091356, 0.003697101, 0.003051713, 0.002552861, 0.00231704, 
    0.002374944, 0.002520517, 0.002616245, 0.00253084, 0.002148377, 
    0.00176327, 0.001461944, 0.001219653, 0.001061479, 0.001307776,
  0.00399728, 0.003615759, 0.002982126, 0.002287228, 0.002024538, 
    0.002016578, 0.002147352, 0.002244485, 0.002250283, 0.001979951, 
    0.001672085, 0.001458371, 0.001295087, 0.001069159, 0.0009389014,
  0.00381568, 0.003384754, 0.002768342, 0.002089716, 0.00172478, 0.001626145, 
    0.001764938, 0.001835079, 0.00186376, 0.001679825, 0.001474185, 
    0.001372483, 0.001262294, 0.001130617, 0.0009346181,
  0.003571734, 0.003316985, 0.00314422, 0.002750717, 0.00240088, 0.002484387, 
    0.00270734, 0.003053278, 0.00279535, 0.002232094, 0.001565275, 
    0.001385791, 0.001120465, 0.001470955, 0.001870107,
  0.003558639, 0.003361169, 0.00308127, 0.002541964, 0.002003448, 
    0.002047195, 0.002390611, 0.002772039, 0.002827407, 0.002438905, 
    0.001972489, 0.001659344, 0.001272951, 0.001198198, 0.001645613,
  0.003500998, 0.003272867, 0.002978675, 0.002412696, 0.001814874, 
    0.001791365, 0.002091391, 0.002425956, 0.002535632, 0.002385169, 
    0.002150039, 0.001967701, 0.001579317, 0.00133208, 0.001443357,
  0.003487808, 0.003274466, 0.002943645, 0.002264089, 0.001665194, 
    0.001655894, 0.001782764, 0.001915025, 0.002023682, 0.00209598, 
    0.00206391, 0.002062382, 0.001933185, 0.001580617, 0.001480198,
  0.003380563, 0.003123377, 0.002861609, 0.002125512, 0.001519271, 
    0.001419189, 0.001602834, 0.001476387, 0.001483834, 0.001807519, 
    0.001984891, 0.002017051, 0.002081044, 0.001911102, 0.001629503,
  0.003248968, 0.002982107, 0.002673606, 0.001985599, 0.001375065, 
    0.001163693, 0.00127083, 0.00132979, 0.001388074, 0.001449729, 
    0.001542696, 0.001664996, 0.001785393, 0.001901915, 0.001796752,
  0.003141603, 0.002835838, 0.002516739, 0.001839317, 0.001220549, 
    0.001006886, 0.0009940437, 0.0009951729, 0.001003334, 0.001023751, 
    0.001057374, 0.00119328, 0.001383047, 0.001545751, 0.00172424,
  0.003012037, 0.002633022, 0.002313109, 0.001605442, 0.00109624, 
    0.0008812035, 0.0008397801, 0.0007931886, 0.0007617666, 0.0007417716, 
    0.0007438876, 0.0008345159, 0.001024061, 0.001279636, 0.001487123,
  0.002820328, 0.002491243, 0.00207251, 0.001253147, 0.0009064778, 
    0.0008184955, 0.000775018, 0.0007334251, 0.0006794692, 0.0006521214, 
    0.0006132985, 0.0006418448, 0.0007421927, 0.001016258, 0.001231109,
  0.002544786, 0.002249935, 0.001694813, 0.001083715, 0.000853806, 
    0.0007574818, 0.0007248382, 0.0006756171, 0.0006131597, 0.0005458441, 
    0.0005124791, 0.0005417839, 0.0005891242, 0.0007818033, 0.001002458,
  0.001644808, 0.001305958, 0.001049229, 0.0009811468, 0.0009680468, 
    0.0009295014, 0.0008908338, 0.0009862294, 0.001120047, 0.001221972, 
    0.001373493, 0.001599346, 0.00167826, 0.001538307, 0.001363247,
  0.001841619, 0.001411724, 0.00105779, 0.0009232163, 0.0008502901, 
    0.0007121126, 0.0007502104, 0.0007685352, 0.0008001725, 0.000857058, 
    0.001018541, 0.001369725, 0.001472905, 0.001400027, 0.001312193,
  0.001800334, 0.001524498, 0.001303046, 0.0009317927, 0.0008141127, 
    0.0006227801, 0.0006685999, 0.0006436678, 0.00062056, 0.0006385393, 
    0.0006935248, 0.000972163, 0.00126503, 0.00138174, 0.001493831,
  0.001802726, 0.001524164, 0.001354987, 0.0009829275, 0.0008546578, 
    0.0007056865, 0.0005346184, 0.0005747867, 0.0005842895, 0.0005790457, 
    0.0005712454, 0.0006793141, 0.0009595053, 0.001234657, 0.001452172,
  0.001807857, 0.00152158, 0.001335564, 0.001026935, 0.0009307024, 
    0.0007196388, 0.0006386363, 0.000424308, 0.0004499831, 0.0005486591, 
    0.0005403392, 0.0005510286, 0.0006529355, 0.0009565349, 0.001330714,
  0.001815931, 0.001545394, 0.0013288, 0.001110489, 0.0009698277, 
    0.000755766, 0.0006586661, 0.0005790835, 0.0005028787, 0.000439567, 
    0.0004216223, 0.0004717033, 0.0005347132, 0.0006636381, 0.001063469,
  0.001811165, 0.001566654, 0.001351053, 0.001149694, 0.000968953, 
    0.0007781312, 0.0007025022, 0.0006317506, 0.000569412, 0.0004916659, 
    0.0004369909, 0.000434387, 0.0004872418, 0.0005428554, 0.0007575863,
  0.001797881, 0.001596456, 0.001371787, 0.001149502, 0.0009710077, 
    0.0008304517, 0.0007454034, 0.0006598338, 0.0005873609, 0.0005290566, 
    0.0004592189, 0.0004250442, 0.0004371836, 0.0004814427, 0.0006604188,
  0.001757639, 0.001600139, 0.001357507, 0.001112767, 0.0009663706, 
    0.0008443494, 0.0007258898, 0.000624066, 0.0005710716, 0.000516897, 
    0.000461027, 0.000412797, 0.0003962998, 0.0004478593, 0.0005854227,
  0.001699945, 0.00149644, 0.001247903, 0.001113616, 0.0009640587, 
    0.0008285373, 0.000695843, 0.0005904722, 0.0005358367, 0.0004473961, 
    0.0004146062, 0.0003999943, 0.0003701199, 0.0004180591, 0.0005290944,
  0.00190767, 0.00182861, 0.001697497, 0.001632659, 0.001613826, 0.001337132, 
    0.0009230187, 0.0006232899, 0.0005525102, 0.0004767743, 0.0004410334, 
    0.000535895, 0.0007844092, 0.001143021, 0.001534709,
  0.002257218, 0.00204217, 0.001819479, 0.001750365, 0.001661486, 
    0.001310462, 0.0008945783, 0.0006593763, 0.000596532, 0.0005623176, 
    0.0004302333, 0.0005033229, 0.0006014645, 0.0007145106, 0.001103414,
  0.002048596, 0.001879252, 0.001837254, 0.001800752, 0.001719477, 
    0.001125013, 0.0009817644, 0.0007794544, 0.0006875502, 0.0006003589, 
    0.0005360468, 0.0004748456, 0.0005619074, 0.0006809899, 0.0009284851,
  0.001913762, 0.001773174, 0.001695133, 0.001647163, 0.00167526, 
    0.001267494, 0.0008982548, 0.0008489216, 0.0007748932, 0.0007301033, 
    0.0006304782, 0.0004984356, 0.0004919597, 0.0005727548, 0.0007571938,
  0.001789882, 0.001638667, 0.001573689, 0.001518887, 0.001509258, 
    0.001413622, 0.001059746, 0.000735841, 0.0006216324, 0.0007595575, 
    0.0007268983, 0.0005726449, 0.0004562205, 0.0005060395, 0.0006219874,
  0.00168202, 0.0015039, 0.001397583, 0.001282385, 0.001236769, 0.001187584, 
    0.001133742, 0.0009214043, 0.0007659352, 0.0006488687, 0.0006246876, 
    0.0005681597, 0.0004708053, 0.000460681, 0.0005708817,
  0.001571119, 0.001411784, 0.001252448, 0.001091423, 0.000943481, 
    0.0009023575, 0.0009240006, 0.00080673, 0.0007262913, 0.000653553, 
    0.0006427145, 0.0005694383, 0.000488464, 0.0004363049, 0.0005362103,
  0.00150006, 0.001318227, 0.001131161, 0.0009193073, 0.0008082752, 
    0.0007301595, 0.0006835712, 0.0006710234, 0.0006208202, 0.0006082536, 
    0.0006097342, 0.0005626608, 0.0004918571, 0.0004310742, 0.0005238682,
  0.001423039, 0.001232773, 0.0009885681, 0.0007758633, 0.0007462507, 
    0.0006527046, 0.0006168975, 0.0005998996, 0.0005671842, 0.0005405249, 
    0.0005749537, 0.0005392884, 0.0004757093, 0.0004322263, 0.0004894037,
  0.001272057, 0.001023981, 0.0008254665, 0.0007081704, 0.0006733424, 
    0.0006270459, 0.0005900778, 0.0005750564, 0.0005391904, 0.0005120735, 
    0.0005369482, 0.0005064388, 0.0004410576, 0.0004097887, 0.000451037,
  0.001400018, 0.00139149, 0.001259903, 0.001213929, 0.001277425, 
    0.001494759, 0.001556923, 0.001348207, 0.001112914, 0.0008542673, 
    0.0007070147, 0.0005589618, 0.0006642734, 0.001032161, 0.001647825,
  0.00152797, 0.0013999, 0.001281855, 0.001181653, 0.001338838, 0.001490079, 
    0.001372477, 0.001164063, 0.0009669877, 0.0007418655, 0.000593851, 
    0.0005700403, 0.00073637, 0.001018405, 0.00151486,
  0.00134989, 0.001195028, 0.001122857, 0.001158699, 0.001357898, 
    0.001157956, 0.001141974, 0.0009173836, 0.0007485735, 0.0006342258, 
    0.0005890948, 0.0005704362, 0.0007377066, 0.001130308, 0.001601721,
  0.001274819, 0.001128968, 0.001047278, 0.001025297, 0.001128588, 
    0.001077511, 0.0007702378, 0.0007286791, 0.0006255739, 0.0005892835, 
    0.0005521876, 0.0005855267, 0.0007680571, 0.001100852, 0.001468016,
  0.001203559, 0.001042816, 0.0009380149, 0.0008270773, 0.0009391172, 
    0.0009655415, 0.0008659541, 0.0005795921, 0.0004815386, 0.0005954275, 
    0.0005803498, 0.0005697064, 0.0007155468, 0.00104457, 0.001367149,
  0.00118802, 0.00102883, 0.0008982109, 0.0007144334, 0.0007308106, 
    0.0008996845, 0.0009670362, 0.0008156862, 0.0006702113, 0.0006415723, 
    0.0005505196, 0.0005701453, 0.000675539, 0.0009978685, 0.001292989,
  0.001158669, 0.001060347, 0.0009726989, 0.0008350351, 0.0008264756, 
    0.0009409014, 0.001018211, 0.0008912592, 0.0007624577, 0.0006778945, 
    0.00063133, 0.0005899985, 0.0007143412, 0.001012572, 0.001299137,
  0.001151163, 0.001079287, 0.001006391, 0.0009089863, 0.0009404841, 
    0.0009768406, 0.0009571888, 0.0008404463, 0.0007062397, 0.0006545089, 
    0.0006007717, 0.0005957836, 0.0007421511, 0.001000811, 0.001255763,
  0.001106896, 0.001022819, 0.0008690823, 0.0007824085, 0.0009055233, 
    0.0009260441, 0.0008737325, 0.000745683, 0.0006563104, 0.0005941071, 
    0.0005493627, 0.0005736793, 0.0006984943, 0.0009704908, 0.001165337,
  0.0009945076, 0.000804599, 0.0007192523, 0.0006957232, 0.0007768238, 
    0.0008263242, 0.0007776055, 0.0007237532, 0.0006055292, 0.0005074374, 
    0.0005002827, 0.0005376404, 0.0006321866, 0.0009065329, 0.00118516,
  0.001034401, 0.001055592, 0.0009596502, 0.0008412446, 0.0008794856, 
    0.0008796429, 0.0008714689, 0.0008637072, 0.001063479, 0.001409666, 
    0.00161258, 0.001377993, 0.001169014, 0.00101096, 0.0008229619,
  0.001238875, 0.001148734, 0.001027727, 0.0008702846, 0.0009099949, 
    0.0009227512, 0.001038971, 0.001016089, 0.001188695, 0.001441363, 
    0.001502745, 0.001299668, 0.001139406, 0.0008379028, 0.0007645772,
  0.001237273, 0.001167428, 0.001089737, 0.0009076091, 0.0008843861, 
    0.0008201971, 0.001070736, 0.001119587, 0.001236216, 0.001423151, 
    0.001366949, 0.001199162, 0.001091724, 0.0009122733, 0.0008714764,
  0.001238869, 0.001194188, 0.00113326, 0.0009157935, 0.000881592, 
    0.0008376971, 0.0007500318, 0.0009447588, 0.00110769, 0.001233355, 
    0.001120166, 0.001054821, 0.00104808, 0.0009882838, 0.001009783,
  0.001240056, 0.001184394, 0.001120812, 0.0008967721, 0.0008516276, 
    0.0008370466, 0.0008078321, 0.0005567301, 0.0005761823, 0.0008904942, 
    0.0009217422, 0.0007665027, 0.0009419784, 0.001132901, 0.001153922,
  0.001249354, 0.00121533, 0.001122808, 0.0009330978, 0.0008497242, 
    0.0007687519, 0.0007451077, 0.0007404902, 0.0006085008, 0.0005823851, 
    0.0005713984, 0.0007236112, 0.001097428, 0.001278338, 0.001282173,
  0.001243348, 0.001221582, 0.001177367, 0.0009829332, 0.0008517843, 
    0.0007261246, 0.0006715029, 0.0006438607, 0.0006137009, 0.0005444862, 
    0.00063122, 0.0009619766, 0.001353006, 0.001495736, 0.001453166,
  0.001245347, 0.001239428, 0.00115243, 0.0009566618, 0.0007977359, 
    0.0007069603, 0.0006484597, 0.0006223857, 0.0005948172, 0.000679738, 
    0.0008896512, 0.001326223, 0.001555436, 0.001592943, 0.001588374,
  0.001155579, 0.001115378, 0.0009710206, 0.0008263192, 0.0007573419, 
    0.0006772476, 0.0006834587, 0.0006920794, 0.0007251316, 0.0008472528, 
    0.001162155, 0.001522094, 0.001595051, 0.001532747, 0.001486298,
  0.00102505, 0.0008584465, 0.0007708358, 0.0007497828, 0.0007291737, 
    0.0006973778, 0.0007198097, 0.0008167292, 0.0009016356, 0.0009919099, 
    0.001165804, 0.001385948, 0.001425983, 0.001464705, 0.001525458,
  0.001400537, 0.001130762, 0.0009126462, 0.0008348114, 0.0009494098, 
    0.001112406, 0.001350562, 0.001403357, 0.001378253, 0.001329444, 
    0.001313142, 0.001440554, 0.001617566, 0.001584261, 0.00156544,
  0.001621519, 0.00126982, 0.001001821, 0.0008828363, 0.0009582398, 
    0.001092337, 0.001360674, 0.001452238, 0.00151263, 0.001578733, 
    0.001763652, 0.001925451, 0.001841345, 0.001632531, 0.001652476,
  0.001491602, 0.001257436, 0.001105424, 0.0009100071, 0.0009303685, 
    0.0009886986, 0.001224161, 0.001340848, 0.001418798, 0.00145748, 
    0.001495443, 0.001601002, 0.001680644, 0.001696824, 0.001641309,
  0.001385191, 0.001206329, 0.001114854, 0.0009130169, 0.0009319472, 
    0.001028884, 0.00110198, 0.001180638, 0.001192288, 0.001239553, 
    0.001236226, 0.001272394, 0.00137108, 0.001460005, 0.001510655,
  0.00126401, 0.001171602, 0.001082409, 0.000899911, 0.0009131963, 
    0.0009641332, 0.001118504, 0.0009058382, 0.0009178494, 0.001122701, 
    0.001092402, 0.001029341, 0.001073889, 0.001175911, 0.001313361,
  0.001259493, 0.001176664, 0.001053731, 0.00093238, 0.0009225672, 
    0.0009143528, 0.0009626435, 0.0009458924, 0.0007828056, 0.0008486368, 
    0.0008829923, 0.0009648051, 0.0009874178, 0.0009996864, 0.001088727,
  0.00127878, 0.001200202, 0.001104464, 0.0009737898, 0.0009097174, 
    0.0009265571, 0.000941578, 0.0008734871, 0.0008049695, 0.000764017, 
    0.0007736592, 0.0008832732, 0.0009526635, 0.0009604666, 0.00104769,
  0.00125759, 0.001199468, 0.001107566, 0.0009508182, 0.0009088139, 
    0.000959714, 0.00105661, 0.001090862, 0.0009989265, 0.0008281903, 
    0.0008092371, 0.0007924899, 0.0008673089, 0.001006345, 0.001068001,
  0.001232714, 0.001152436, 0.0009533829, 0.0008569018, 0.0008802523, 
    0.0009283614, 0.001099031, 0.001191192, 0.001180597, 0.001084005, 
    0.001125232, 0.001110449, 0.001126133, 0.001085576, 0.001206647,
  0.001126584, 0.0009195128, 0.0008619379, 0.0008160305, 0.0008216816, 
    0.0008552846, 0.001074977, 0.001334811, 0.001416734, 0.001443293, 
    0.001496613, 0.001435477, 0.001423885, 0.001310806, 0.001331111,
  0.001249313, 0.001257483, 0.001153896, 0.001125771, 0.001229582, 
    0.001076905, 0.0009795481, 0.0009682788, 0.001126018, 0.001328143, 
    0.001338999, 0.001034625, 0.0007495118, 0.0008262652, 0.0008276614,
  0.001555387, 0.001476521, 0.001291156, 0.001159214, 0.001177554, 
    0.001018545, 0.0009814291, 0.0009433152, 0.0009921457, 0.001205993, 
    0.001328904, 0.001306093, 0.0008819611, 0.000720128, 0.0007491629,
  0.001521306, 0.001500939, 0.001444671, 0.001176944, 0.001051857, 
    0.000925357, 0.0009678291, 0.0009421946, 0.0009627182, 0.001014917, 
    0.001137851, 0.001443507, 0.00119267, 0.0009241049, 0.0008173009,
  0.001570038, 0.001527684, 0.001453408, 0.001209515, 0.001090627, 
    0.0009901354, 0.0008898249, 0.0008974616, 0.000956822, 0.001004654, 
    0.000961808, 0.001260574, 0.001544482, 0.001243409, 0.000996485,
  0.001599668, 0.001532565, 0.001433837, 0.001226271, 0.001126588, 
    0.001019011, 0.001019011, 0.0008436634, 0.0008880103, 0.001056124, 
    0.0009472661, 0.001056706, 0.00139599, 0.001429227, 0.001292743,
  0.001625134, 0.001555111, 0.001475515, 0.00131612, 0.00115666, 0.00103363, 
    0.001023357, 0.001102204, 0.001203041, 0.001106169, 0.0009101456, 
    0.0009771342, 0.001224922, 0.001480924, 0.001437394,
  0.00167946, 0.001651968, 0.001586126, 0.00140906, 0.001171784, 0.00104822, 
    0.001026136, 0.001141989, 0.001351707, 0.001223688, 0.0009932544, 
    0.0009561126, 0.001151123, 0.001406565, 0.001535985,
  0.001865505, 0.001846657, 0.0017643, 0.001478177, 0.001236918, 0.001036793, 
    0.000983173, 0.001160284, 0.001448185, 0.001375754, 0.001088568, 
    0.001000722, 0.001096562, 0.001326061, 0.001473071,
  0.002302455, 0.002209106, 0.001967799, 0.001582551, 0.001253256, 
    0.0009929057, 0.0009362854, 0.001159316, 0.001455396, 0.001514607, 
    0.001276609, 0.001103299, 0.001152156, 0.001291686, 0.001316047,
  0.00270017, 0.002395989, 0.002078322, 0.001639964, 0.001352292, 
    0.0009300431, 0.0008748749, 0.001138592, 0.001448575, 0.001617, 
    0.00144046, 0.001218242, 0.00128827, 0.001338915, 0.001346911,
  0.001284378, 0.001568092, 0.001744971, 0.001742869, 0.001675705, 
    0.001632506, 0.001539956, 0.001308693, 0.001065109, 0.001212723, 
    0.001116331, 0.001016268, 0.0009282693, 0.0009883634, 0.001035925,
  0.002169358, 0.002270683, 0.002164775, 0.002067037, 0.001998119, 
    0.001837339, 0.001720852, 0.001342084, 0.001003664, 0.001235298, 
    0.001161457, 0.001084816, 0.001016676, 0.0009105866, 0.0009474595,
  0.002510078, 0.002663171, 0.002654094, 0.002335898, 0.002089278, 
    0.001967084, 0.001874831, 0.001379339, 0.0009784348, 0.00129457, 
    0.001180998, 0.001187587, 0.001076083, 0.001099208, 0.0009871003,
  0.002914312, 0.002881221, 0.002760867, 0.002537093, 0.002432807, 
    0.002310597, 0.001834066, 0.00113217, 0.000911614, 0.001226493, 
    0.001217834, 0.001237748, 0.001159939, 0.001073361, 0.0009541531,
  0.003185764, 0.003051563, 0.002860496, 0.002693129, 0.002567156, 
    0.00223355, 0.001681461, 0.0007767713, 0.0007946956, 0.001172188, 
    0.001265256, 0.001291576, 0.001324086, 0.001106598, 0.001043228,
  0.003177981, 0.003085364, 0.002897626, 0.002744904, 0.00247161, 
    0.001958281, 0.001223891, 0.0009135256, 0.000949936, 0.001212212, 
    0.001246706, 0.001304081, 0.001479472, 0.001406849, 0.001211838,
  0.003175076, 0.003138476, 0.002974945, 0.002640017, 0.002175937, 
    0.001486321, 0.001061235, 0.001006868, 0.001082231, 0.001373188, 
    0.001260724, 0.001312767, 0.001483083, 0.001581136, 0.001535005,
  0.003296023, 0.003160228, 0.002917278, 0.002300079, 0.001725942, 
    0.001151911, 0.001015059, 0.001028723, 0.00112753, 0.001441296, 
    0.001271372, 0.001287644, 0.001403664, 0.001508903, 0.001612737,
  0.003352856, 0.00296998, 0.002641053, 0.00183779, 0.001370882, 0.001033843, 
    0.0009707122, 0.001079646, 0.001232314, 0.001425296, 0.001293534, 
    0.00130927, 0.001368242, 0.001467972, 0.001485913,
  0.003374136, 0.002752101, 0.002322861, 0.001759847, 0.001412822, 
    0.000924892, 0.0009329832, 0.001141986, 0.00128556, 0.001375769, 
    0.001295805, 0.001340687, 0.001432607, 0.001563936, 0.001447234,
  0.001998475, 0.002314961, 0.002556758, 0.002540882, 0.00248721, 
    0.002484994, 0.002559658, 0.002477501, 0.002158856, 0.001381967, 
    0.001031212, 0.001232639, 0.001222166, 0.00118544, 0.001146239,
  0.002932234, 0.002871537, 0.002628975, 0.002382956, 0.002099084, 
    0.002165242, 0.002333462, 0.002183055, 0.001719001, 0.001131991, 
    0.00103071, 0.001287189, 0.001280928, 0.00115736, 0.001136445,
  0.003112193, 0.002818367, 0.002496885, 0.002024746, 0.00182134, 
    0.001691838, 0.001802474, 0.001574978, 0.001135978, 0.001030647, 
    0.001191919, 0.001284089, 0.001329351, 0.001354576, 0.001331224,
  0.003061235, 0.002572264, 0.002249012, 0.001717596, 0.001502747, 
    0.001396901, 0.00116488, 0.001126714, 0.00091627, 0.001012909, 
    0.001116561, 0.001276416, 0.001322556, 0.001414155, 0.00136852,
  0.002956212, 0.002375514, 0.0019967, 0.001432494, 0.001271739, 0.001048106, 
    0.001029161, 0.0007515305, 0.0007205075, 0.001005924, 0.001163737, 
    0.001290554, 0.00134895, 0.001430978, 0.001529053,
  0.003035051, 0.00233738, 0.001893496, 0.001526291, 0.001334551, 
    0.001067003, 0.0009300863, 0.0009627963, 0.0009962447, 0.001044413, 
    0.001198598, 0.001274217, 0.001407, 0.001518862, 0.001538701,
  0.003229211, 0.002582107, 0.002152237, 0.001684969, 0.001435791, 
    0.001101285, 0.0009430086, 0.001002117, 0.001177998, 0.001253902, 
    0.00128788, 0.001391993, 0.001543464, 0.001614135, 0.001461962,
  0.003423722, 0.002751032, 0.002464822, 0.001970819, 0.00162273, 
    0.001136543, 0.000932932, 0.0010661, 0.001332735, 0.001374673, 
    0.001451472, 0.001552107, 0.001697867, 0.001671358, 0.001444669,
  0.003541504, 0.003165876, 0.002806206, 0.002298226, 0.001828848, 
    0.001207936, 0.0009220462, 0.001123178, 0.001398083, 0.001536121, 
    0.001584042, 0.001709006, 0.00174799, 0.001649103, 0.001539108,
  0.003675838, 0.003341851, 0.002839515, 0.002638722, 0.001956707, 
    0.001084597, 0.0008805208, 0.001212411, 0.00148187, 0.001571179, 
    0.00172617, 0.001812155, 0.001750797, 0.001606184, 0.001576289,
  0.002023255, 0.00156714, 0.001505291, 0.001352354, 0.001212348, 
    0.001175889, 0.001057032, 0.001149139, 0.001233234, 0.001295885, 
    0.001247931, 0.001269383, 0.001249059, 0.001192911, 0.001185439,
  0.002459365, 0.001984647, 0.001887767, 0.001723398, 0.00150707, 
    0.001182432, 0.00107554, 0.0009526468, 0.001046175, 0.001152562, 
    0.001197117, 0.001203155, 0.001149873, 0.001022776, 0.001053969,
  0.002725532, 0.002460827, 0.002437987, 0.002139937, 0.001836214, 
    0.001334287, 0.001050396, 0.0009954441, 0.001102077, 0.001209085, 
    0.001307325, 0.001334185, 0.001291022, 0.001265074, 0.001252035,
  0.003143962, 0.002956377, 0.002786584, 0.002444387, 0.002226264, 
    0.001725416, 0.001125923, 0.0009390645, 0.001147905, 0.001367634, 
    0.001456737, 0.001482422, 0.00145214, 0.001534939, 0.001603282,
  0.003673364, 0.003373599, 0.002933776, 0.002718107, 0.002455305, 
    0.001948854, 0.001156953, 0.0009456789, 0.001074393, 0.001503126, 
    0.001534402, 0.001531995, 0.001476295, 0.001517579, 0.001545466,
  0.004035862, 0.003568753, 0.002902469, 0.00292909, 0.002426534, 
    0.001874286, 0.001237738, 0.001325985, 0.001506072, 0.001610407, 
    0.001528266, 0.001486505, 0.001486655, 0.001431756, 0.001444416,
  0.004063688, 0.003353891, 0.002742673, 0.002918403, 0.002221111, 
    0.001583233, 0.001232001, 0.00144507, 0.001660802, 0.001579242, 
    0.001482416, 0.001480072, 0.001450513, 0.001487756, 0.001552948,
  0.003867687, 0.003105125, 0.002503014, 0.002644158, 0.001937414, 
    0.001351057, 0.001304501, 0.001587403, 0.001600618, 0.001474668, 
    0.001387623, 0.001412118, 0.001467121, 0.0015969, 0.001701906,
  0.003683982, 0.002988225, 0.002309989, 0.002213222, 0.001489916, 
    0.001156166, 0.001381414, 0.001621702, 0.001552125, 0.00137987, 
    0.00130355, 0.001348019, 0.001455705, 0.00161325, 0.001738066,
  0.003833327, 0.002932535, 0.002094037, 0.00186018, 0.001163545, 
    0.001145064, 0.001441595, 0.001645076, 0.001507482, 0.00127444, 
    0.001209779, 0.001285896, 0.001388901, 0.001533413, 0.001673669,
  0.002391356, 0.002624394, 0.00267193, 0.002402879, 0.002146144, 
    0.001896047, 0.001395901, 0.001289257, 0.001259055, 0.001331127, 
    0.001332062, 0.001379311, 0.001395414, 0.001206638, 0.0010891,
  0.002976497, 0.002997434, 0.002595461, 0.00224038, 0.002055267, 
    0.001598444, 0.001415577, 0.001157205, 0.001183074, 0.00122419, 
    0.001340362, 0.001384927, 0.001421232, 0.00131442, 0.001213562,
  0.003265969, 0.002817159, 0.002324073, 0.002158189, 0.001817216, 
    0.00148409, 0.001306112, 0.001220545, 0.001254023, 0.001304184, 
    0.001319208, 0.001352084, 0.001378661, 0.001328887, 0.001304108,
  0.003424564, 0.002719976, 0.002071502, 0.00202805, 0.001645992, 
    0.001400016, 0.001135199, 0.001199209, 0.001260131, 0.001307525, 
    0.001296729, 0.001348895, 0.001372512, 0.001373015, 0.001344785,
  0.003422529, 0.002532559, 0.00196223, 0.001897656, 0.001484763, 
    0.001357727, 0.001300355, 0.001006838, 0.001052418, 0.001268604, 
    0.001326761, 0.00138725, 0.001473137, 0.001530742, 0.001443243,
  0.003550394, 0.002436428, 0.001834546, 0.001836773, 0.001450569, 
    0.001321492, 0.001340733, 0.001250569, 0.001167518, 0.001204263, 
    0.001278947, 0.00142815, 0.001578106, 0.001612906, 0.001625269,
  0.003586102, 0.002437671, 0.001702973, 0.001775732, 0.001427899, 0.0013506, 
    0.001326216, 0.001240181, 0.00120937, 0.00123474, 0.00127775, 
    0.001414539, 0.00153822, 0.001657763, 0.001656834,
  0.003577456, 0.002505054, 0.001728736, 0.001582648, 0.001389392, 
    0.001471937, 0.00129899, 0.001226468, 0.001249312, 0.00126383, 
    0.001253236, 0.001349048, 0.001463529, 0.001602181, 0.001576254,
  0.003693986, 0.002737247, 0.001799097, 0.001424386, 0.001327593, 
    0.001415759, 0.001286364, 0.001265121, 0.001303656, 0.001293631, 
    0.001212656, 0.001263138, 0.001381033, 0.001551295, 0.001549174,
  0.003939443, 0.002864618, 0.001907922, 0.001514651, 0.00131124, 
    0.001414165, 0.001335373, 0.001339029, 0.001304406, 0.001148264, 
    0.001116435, 0.001206294, 0.001315865, 0.001509126, 0.001598881,
  0.001813841, 0.001673155, 0.001604198, 0.001214347, 0.001062315, 
    0.001014812, 0.000942568, 0.000973176, 0.001030535, 0.001106765, 
    0.001099233, 0.001076101, 0.001233467, 0.001212606, 0.00114514,
  0.002261061, 0.001868877, 0.001728663, 0.001337949, 0.001171186, 
    0.001054152, 0.001018593, 0.001038519, 0.001082849, 0.001086776, 
    0.001054364, 0.001089493, 0.001141719, 0.001165287, 0.001128158,
  0.002754187, 0.002226085, 0.001964876, 0.00146257, 0.001284166, 
    0.001095751, 0.001107941, 0.001098263, 0.001105138, 0.001164208, 
    0.001129727, 0.001107378, 0.001178474, 0.00119412, 0.001222799,
  0.003170833, 0.002677941, 0.002246505, 0.001790871, 0.001519443, 
    0.001332292, 0.001107432, 0.001148975, 0.001170891, 0.001204519, 
    0.001183136, 0.001123667, 0.001169567, 0.001186846, 0.00120774,
  0.003508218, 0.003108826, 0.002622003, 0.002193057, 0.001833153, 
    0.001528028, 0.001423411, 0.001042557, 0.001007011, 0.001242013, 
    0.001248181, 0.001173039, 0.001161256, 0.001147202, 0.001245497,
  0.003804522, 0.003453966, 0.002826938, 0.002506927, 0.002165718, 
    0.001839248, 0.001545916, 0.001399336, 0.001289748, 0.001259781, 
    0.001226734, 0.001190279, 0.001186192, 0.001145842, 0.001257964,
  0.004207509, 0.003882814, 0.003139538, 0.002741941, 0.002389005, 
    0.002017962, 0.001724042, 0.001583946, 0.001472315, 0.001426453, 
    0.001361657, 0.001251329, 0.001168959, 0.001167283, 0.001276913,
  0.004265041, 0.00397795, 0.003340093, 0.002900003, 0.002581197, 0.00231364, 
    0.002084364, 0.00188994, 0.001804825, 0.001705278, 0.001527816, 
    0.001307214, 0.001160203, 0.001194785, 0.00126086,
  0.004111379, 0.003888241, 0.003414546, 0.00307112, 0.002807352, 
    0.002594536, 0.002377647, 0.002238694, 0.002107314, 0.001925709, 
    0.001654679, 0.001341003, 0.00120226, 0.001179926, 0.001251903,
  0.00383683, 0.003575038, 0.003516774, 0.003360188, 0.003051528, 
    0.002866803, 0.002643678, 0.002534908, 0.002286805, 0.001978721, 
    0.001592398, 0.001275414, 0.001110811, 0.001144366, 0.001234491,
  0.002527491, 0.002457368, 0.002415891, 0.002236841, 0.002068738, 
    0.001718172, 0.001472396, 0.001307873, 0.00133375, 0.001294091, 
    0.001278337, 0.001088368, 0.001047212, 0.0009443313, 0.000808906,
  0.003113473, 0.002953666, 0.002709788, 0.002389435, 0.002058698, 
    0.001936346, 0.001572671, 0.001537516, 0.001578349, 0.00145545, 
    0.001443601, 0.001278873, 0.001182455, 0.00103791, 0.0009440678,
  0.003493187, 0.003356352, 0.003132513, 0.002586344, 0.002417365, 
    0.00202123, 0.002035638, 0.001995678, 0.001948176, 0.001891423, 
    0.001816872, 0.001664548, 0.001512131, 0.001296396, 0.001171717,
  0.003798401, 0.003701091, 0.003487866, 0.003041219, 0.002837692, 
    0.002314449, 0.002163875, 0.002252431, 0.002208471, 0.002179102, 
    0.002054609, 0.001876672, 0.001730429, 0.001617936, 0.00140694,
  0.004125405, 0.003773956, 0.003542385, 0.003285918, 0.003214238, 
    0.003114416, 0.002935791, 0.002444467, 0.002374289, 0.002576141, 
    0.002599271, 0.002495531, 0.002299577, 0.002087654, 0.001788216,
  0.004191882, 0.00394336, 0.003491971, 0.003292907, 0.003310276, 
    0.003387864, 0.003379035, 0.003309284, 0.003214867, 0.003098657, 
    0.00290982, 0.002730318, 0.002597849, 0.002469605, 0.002294212,
  0.004246153, 0.004002531, 0.003601486, 0.003366591, 0.0033944, 0.003457692, 
    0.003477975, 0.003348493, 0.00303218, 0.002771251, 0.002645263, 
    0.002575063, 0.002534931, 0.002462453, 0.002373618,
  0.004430218, 0.00411248, 0.003638614, 0.00348252, 0.003513137, 0.003480121, 
    0.003217819, 0.00275185, 0.002516235, 0.002449537, 0.002400849, 
    0.002306992, 0.002159549, 0.002078023, 0.002037905,
  0.004511569, 0.004070032, 0.003529842, 0.003503077, 0.003345692, 
    0.003002811, 0.002494274, 0.002230708, 0.00215098, 0.002033212, 
    0.001736051, 0.00167223, 0.001706582, 0.001701029, 0.001703236,
  0.004190269, 0.00358775, 0.003459896, 0.003268478, 0.002888601, 
    0.002246081, 0.0019602, 0.001837028, 0.001639183, 0.001321082, 
    0.001331301, 0.001449348, 0.001547823, 0.001552124, 0.001553173,
  0.003089791, 0.003062344, 0.003291399, 0.003169173, 0.003069167, 
    0.003006847, 0.002741517, 0.002364795, 0.002158037, 0.001968549, 
    0.002007035, 0.002125217, 0.00208184, 0.002038803, 0.001833428,
  0.003450035, 0.003378873, 0.003332552, 0.003238891, 0.003172205, 
    0.003122513, 0.002826588, 0.002516588, 0.002275845, 0.002162606, 
    0.002219636, 0.002317388, 0.002344375, 0.002130825, 0.001925909,
  0.003725162, 0.003534386, 0.003425117, 0.003197744, 0.00322898, 
    0.002824391, 0.002756483, 0.002602887, 0.002377816, 0.002374464, 
    0.00246907, 0.00265409, 0.002744669, 0.002712364, 0.002369458,
  0.00390259, 0.003661952, 0.003392256, 0.003103507, 0.003027616, 
    0.002712601, 0.002317614, 0.002245307, 0.002251758, 0.002324692, 
    0.002372374, 0.002527531, 0.002574861, 0.002560711, 0.002456039,
  0.004016749, 0.003503195, 0.003148127, 0.00279655, 0.002615192, 
    0.002442608, 0.002301953, 0.00188818, 0.001857546, 0.001965235, 
    0.001876703, 0.001788289, 0.00162483, 0.001576677, 0.001706136,
  0.00393835, 0.003396646, 0.002804197, 0.002457205, 0.002247379, 
    0.002019321, 0.001912359, 0.001870909, 0.001732385, 0.001330995, 
    0.001146833, 0.001079162, 0.001067226, 0.001057085, 0.001141633,
  0.003751064, 0.003147446, 0.002579495, 0.002073105, 0.001793469, 
    0.001542619, 0.001371736, 0.001290779, 0.00119742, 0.001121669, 
    0.001074792, 0.001019074, 0.001083054, 0.001049364, 0.001055211,
  0.003417548, 0.002800073, 0.002154458, 0.001631673, 0.00136346, 
    0.001187696, 0.001112101, 0.001116036, 0.001114423, 0.001076048, 
    0.001072708, 0.001097995, 0.001113584, 0.001098184, 0.001069541,
  0.002994095, 0.002392636, 0.001656274, 0.001237887, 0.001169352, 
    0.001108531, 0.001085862, 0.001148131, 0.001130524, 0.001082655, 
    0.001145249, 0.00114136, 0.001170747, 0.001146762, 0.001145797,
  0.002573732, 0.001962332, 0.001372958, 0.001161373, 0.001116759, 
    0.001088269, 0.001081124, 0.001169185, 0.001155029, 0.001119566, 
    0.001208185, 0.00119579, 0.001176507, 0.001136245, 0.001086292,
  0.002275156, 0.002163805, 0.002072692, 0.001930306, 0.001897784, 
    0.00172484, 0.001523917, 0.001434153, 0.001385237, 0.001442881, 
    0.001517997, 0.00163543, 0.001798438, 0.002037131, 0.002349679,
  0.002257053, 0.001985563, 0.001712458, 0.001604098, 0.001581147, 
    0.001364836, 0.001232469, 0.001180308, 0.001161088, 0.001195427, 
    0.001355339, 0.001474365, 0.001637766, 0.001778407, 0.002064809,
  0.00217343, 0.001935809, 0.001646587, 0.001280974, 0.001203475, 
    0.001046083, 0.001041243, 0.001068503, 0.001069015, 0.001079721, 
    0.001115754, 0.001195414, 0.00131184, 0.001525972, 0.001954511,
  0.002130368, 0.001886377, 0.001676706, 0.0012813, 0.00115919, 0.001034708, 
    0.0009119933, 0.0009372996, 0.001015363, 0.001088291, 0.001100053, 
    0.001080107, 0.001073384, 0.001185127, 0.001446238,
  0.002236358, 0.001940224, 0.001735382, 0.001363812, 0.001177444, 
    0.001098984, 0.000992923, 0.0008111458, 0.0009034763, 0.001099267, 
    0.001131737, 0.001060188, 0.001053995, 0.001036095, 0.001074252,
  0.002385544, 0.002146279, 0.001849164, 0.001481424, 0.001237177, 
    0.001117657, 0.001052883, 0.001087539, 0.001155409, 0.00108946, 
    0.00108897, 0.001033923, 0.001079639, 0.001039648, 0.00102211,
  0.002602299, 0.002354901, 0.001999134, 0.001580847, 0.001273019, 
    0.001128834, 0.001028907, 0.001113956, 0.001192561, 0.001176762, 
    0.001172967, 0.001097999, 0.001140206, 0.001154881, 0.001175266,
  0.002969422, 0.002685553, 0.002151284, 0.001665771, 0.001368999, 
    0.001237982, 0.001027783, 0.001101449, 0.001226221, 0.001217516, 
    0.001223686, 0.001137151, 0.001206649, 0.001267463, 0.001192394,
  0.003328756, 0.002960913, 0.002257935, 0.001838244, 0.0015319, 0.001331775, 
    0.001107182, 0.001170467, 0.00122252, 0.001216979, 0.001188269, 
    0.001146398, 0.001195814, 0.001228653, 0.001279751,
  0.003535126, 0.003018563, 0.002497492, 0.002189647, 0.001825214, 
    0.001499765, 0.001151378, 0.001192042, 0.001244309, 0.001197562, 
    0.001118049, 0.001105091, 0.001153351, 0.001246107, 0.001325401,
  0.002088611, 0.001889082, 0.001732109, 0.001644355, 0.001601057, 
    0.001556586, 0.001331683, 0.001146242, 0.001105627, 0.001146978, 
    0.001184955, 0.001039756, 0.001086657, 0.001209996, 0.001446452,
  0.002635509, 0.002422628, 0.002214942, 0.002055699, 0.001990179, 
    0.001794801, 0.001585154, 0.001357618, 0.001187353, 0.001122458, 
    0.00108771, 0.000972158, 0.001001475, 0.001179717, 0.001160617,
  0.002997889, 0.002778581, 0.002697467, 0.002478009, 0.002347904, 
    0.001993436, 0.001751881, 0.001527469, 0.001311625, 0.001172619, 
    0.001072314, 0.001018955, 0.00104181, 0.001192926, 0.001161464,
  0.003353157, 0.00317244, 0.00309931, 0.002962675, 0.002768512, 0.002437456, 
    0.001863447, 0.001494503, 0.001285308, 0.001194485, 0.001097431, 
    0.001005544, 0.001051017, 0.001186185, 0.001138107,
  0.003713883, 0.003501497, 0.003433964, 0.003285828, 0.003084493, 
    0.002767953, 0.002292796, 0.001506111, 0.001170783, 0.001205656, 
    0.001106254, 0.001006045, 0.00104705, 0.001198999, 0.001196657,
  0.003985651, 0.003818033, 0.003565831, 0.003447981, 0.003334455, 
    0.003042431, 0.00262265, 0.002106308, 0.001552897, 0.00123728, 
    0.001040177, 0.0009825873, 0.001019721, 0.001114572, 0.001262554,
  0.004215085, 0.004162035, 0.003857358, 0.0035711, 0.00347675, 0.003122103, 
    0.002724112, 0.002226562, 0.001532929, 0.001235048, 0.001067032, 
    0.00104947, 0.001025755, 0.001139157, 0.00125129,
  0.004340478, 0.004115218, 0.003866612, 0.003662394, 0.003514477, 
    0.003112758, 0.002672875, 0.002120843, 0.001526172, 0.001310537, 
    0.001142135, 0.00108764, 0.001073934, 0.001148304, 0.001183939,
  0.004394445, 0.00411048, 0.00365996, 0.003685364, 0.003416157, 0.002955082, 
    0.002643596, 0.002031868, 0.00154368, 0.001287581, 0.001110445, 
    0.001034306, 0.001042477, 0.001102298, 0.001123183,
  0.004054082, 0.003720462, 0.003642159, 0.003508436, 0.003146996, 
    0.002825821, 0.002478607, 0.001907096, 0.00142915, 0.00117037, 
    0.000943625, 0.0009712526, 0.0009741951, 0.001053143, 0.001098591,
  0.003316605, 0.003242862, 0.003205954, 0.003043729, 0.002915078, 
    0.002825421, 0.002774165, 0.002818791, 0.002687682, 0.002362258, 
    0.002162179, 0.001789002, 0.001409121, 0.001078899, 0.0009332568,
  0.003614429, 0.003479273, 0.003411839, 0.003311128, 0.003211683, 
    0.003067709, 0.002855476, 0.002840157, 0.002802695, 0.002527319, 
    0.002296814, 0.001915542, 0.001401177, 0.00105512, 0.0009192184,
  0.003872746, 0.003616328, 0.003453614, 0.003324543, 0.003169668, 
    0.002959545, 0.002909113, 0.002807936, 0.002643291, 0.002284567, 
    0.002053266, 0.001829657, 0.001336475, 0.001080282, 0.001033758,
  0.00409523, 0.003711479, 0.003480831, 0.003182641, 0.002928709, 
    0.002906713, 0.002595793, 0.002399398, 0.002145684, 0.001977051, 
    0.001836924, 0.001518738, 0.001198971, 0.001054074, 0.0009883011,
  0.004252407, 0.003624606, 0.003314298, 0.002907768, 0.002718565, 
    0.002646763, 0.002402562, 0.001819829, 0.001658491, 0.001680228, 
    0.001483047, 0.001285812, 0.001149878, 0.001024709, 0.0009891465,
  0.004174334, 0.003541705, 0.002991602, 0.002634201, 0.002441998, 
    0.002255805, 0.0020203, 0.001848633, 0.001532855, 0.001356212, 
    0.001292134, 0.001162513, 0.001113636, 0.001030223, 0.000981398,
  0.003996512, 0.003326204, 0.002831928, 0.002431377, 0.002215598, 
    0.001862157, 0.001671637, 0.001439824, 0.001296197, 0.001139879, 
    0.001102191, 0.001133841, 0.001098921, 0.001047604, 0.001035315,
  0.003794323, 0.003106876, 0.002609574, 0.002228387, 0.001859457, 
    0.001619915, 0.00148291, 0.001286793, 0.00121256, 0.001163115, 
    0.001094166, 0.001092502, 0.001131661, 0.001126762, 0.001066606,
  0.003512857, 0.00296363, 0.002248737, 0.001808619, 0.001562875, 
    0.001437893, 0.001346778, 0.001243431, 0.001198044, 0.001146145, 
    0.001066206, 0.001027543, 0.0009846304, 0.001036402, 0.001006943,
  0.003086281, 0.002482834, 0.001855139, 0.00151699, 0.001303939, 
    0.001168165, 0.001133308, 0.001167298, 0.001122908, 0.001009758, 
    0.0008898739, 0.0008993532, 0.0008513692, 0.0008725924, 0.0009107482,
  0.002112158, 0.002025351, 0.00199209, 0.001991922, 0.001804552, 
    0.001442884, 0.001308641, 0.001364847, 0.001515829, 0.00169786, 
    0.001927882, 0.002162898, 0.002252889, 0.002202434, 0.001924394,
  0.002213786, 0.0019155, 0.001719664, 0.001642483, 0.001626287, 0.001207977, 
    0.00111091, 0.001126486, 0.001202984, 0.001417874, 0.001751764, 
    0.002395248, 0.002420152, 0.002107078, 0.001833839,
  0.002215345, 0.001879044, 0.001662513, 0.001416462, 0.00133742, 
    0.001123555, 0.001045272, 0.00104386, 0.001100293, 0.001296857, 
    0.001605791, 0.002153061, 0.002511815, 0.002099404, 0.001725631,
  0.00220403, 0.001852011, 0.001641401, 0.001305677, 0.001199859, 
    0.001125003, 0.0009302668, 0.0009520866, 0.001012139, 0.001175334, 
    0.001445466, 0.001869816, 0.002021194, 0.001811325, 0.001604962,
  0.002195518, 0.001814386, 0.001627241, 0.001276664, 0.001183686, 
    0.001147424, 0.001128625, 0.0008704488, 0.0008685838, 0.001098815, 
    0.001248664, 0.001505821, 0.001652768, 0.001676182, 0.001662399,
  0.002249534, 0.001842345, 0.0015711, 0.001330138, 0.001167903, 0.001122033, 
    0.001107283, 0.001087512, 0.001010937, 0.001083683, 0.001144234, 
    0.001294004, 0.001443268, 0.00146719, 0.001419132,
  0.002188366, 0.001881118, 0.001562556, 0.001330525, 0.001143112, 
    0.001108559, 0.001115392, 0.001101837, 0.001117151, 0.001082114, 
    0.001101523, 0.001144501, 0.001167317, 0.001217375, 0.00120898,
  0.002055878, 0.001850958, 0.001509493, 0.00121781, 0.001123229, 
    0.001090585, 0.001096406, 0.001103805, 0.001100294, 0.00111279, 
    0.001063702, 0.001122186, 0.001111585, 0.001074134, 0.001054958,
  0.001914492, 0.001801158, 0.001368627, 0.001208049, 0.001117554, 
    0.001079565, 0.001107253, 0.001142058, 0.001161555, 0.001156429, 
    0.001104349, 0.001077056, 0.00104664, 0.001085487, 0.001012648,
  0.001732987, 0.001588756, 0.001414314, 0.001285519, 0.001146353, 
    0.001074743, 0.001089128, 0.001145332, 0.001150055, 0.001119274, 
    0.001059913, 0.0009797105, 0.0009745049, 0.000983621, 0.001023851,
  0.001679172, 0.001780919, 0.001763241, 0.001655435, 0.001516254, 
    0.001180697, 0.001038385, 0.0009391616, 0.000961786, 0.00109271, 
    0.001217247, 0.001498506, 0.001682949, 0.001789105, 0.001850318,
  0.002017917, 0.002043611, 0.001892881, 0.00172742, 0.001492274, 
    0.001144601, 0.001061305, 0.001008771, 0.0009871792, 0.001045103, 
    0.001256008, 0.001611962, 0.00187217, 0.001882194, 0.001808438,
  0.002122894, 0.002101155, 0.001964199, 0.001712205, 0.001417849, 
    0.001161212, 0.001033959, 0.001060092, 0.001008907, 0.001103056, 
    0.001267507, 0.001683382, 0.002063753, 0.002030218, 0.001998395,
  0.002184621, 0.00213365, 0.00195426, 0.00171077, 0.001432589, 0.001168063, 
    0.000929179, 0.0009950628, 0.001030483, 0.00113587, 0.00122307, 
    0.001587643, 0.002156883, 0.002257828, 0.002139231,
  0.002266129, 0.002145958, 0.001927171, 0.00163654, 0.001415567, 
    0.001178297, 0.001060827, 0.0008596627, 0.0008810684, 0.001106195, 
    0.001170049, 0.001375842, 0.00180469, 0.002196679, 0.002196921,
  0.002304009, 0.002159676, 0.001874744, 0.001611467, 0.001410088, 
    0.001219795, 0.001078297, 0.001086531, 0.001045468, 0.001074033, 
    0.001111134, 0.001198873, 0.001367457, 0.001647701, 0.001842292,
  0.002344368, 0.002175437, 0.001861978, 0.001561204, 0.001385767, 
    0.001213452, 0.001093246, 0.001103285, 0.001083104, 0.001059547, 
    0.001095768, 0.001149626, 0.001215679, 0.001272944, 0.001358372,
  0.002356185, 0.002184846, 0.001814315, 0.001528045, 0.001364583, 
    0.001202239, 0.001135946, 0.001121759, 0.001111621, 0.001062975, 
    0.001044737, 0.001077571, 0.001170244, 0.001216416, 0.001261017,
  0.00241369, 0.002146902, 0.001740605, 0.001495152, 0.00134824, 0.001193293, 
    0.001147731, 0.00111769, 0.001124391, 0.001089169, 0.001040789, 
    0.001032359, 0.001100803, 0.001188036, 0.001279438,
  0.002387988, 0.00207011, 0.001720521, 0.00144877, 0.00130935, 0.001179261, 
    0.0011719, 0.001135518, 0.001150108, 0.001122801, 0.001071163, 
    0.001040273, 0.001051586, 0.001140214, 0.001292879,
  0.002513873, 0.002019904, 0.001494236, 0.001362816, 0.001316584, 
    0.001178481, 0.0009689892, 0.0009492526, 0.0009257091, 0.001059558, 
    0.001111491, 0.001171298, 0.001325354, 0.001638255, 0.002319196,
  0.002856578, 0.001966121, 0.001483622, 0.001284458, 0.001248119, 
    0.001061839, 0.0009741609, 0.0009923939, 0.0009856843, 0.000969036, 
    0.00108708, 0.001226756, 0.001390542, 0.001480873, 0.001764344,
  0.002788247, 0.001847394, 0.001480999, 0.001232771, 0.001143947, 
    0.001031945, 0.000983858, 0.001048906, 0.00107165, 0.001095958, 
    0.001111416, 0.001320398, 0.001447933, 0.001529124, 0.001588603,
  0.002675972, 0.001800342, 0.001454622, 0.001183063, 0.001163282, 
    0.001010616, 0.000910688, 0.001015262, 0.00108037, 0.00118359, 
    0.001228863, 0.001297792, 0.001474046, 0.001692746, 0.001610446,
  0.002535899, 0.001703167, 0.001414929, 0.001171876, 0.001131305, 
    0.001104724, 0.001016128, 0.0008869951, 0.0009368843, 0.00119089, 
    0.001295642, 0.001367456, 0.001442706, 0.001692899, 0.001899888,
  0.002380907, 0.001736355, 0.001368934, 0.001192774, 0.001088912, 
    0.001140061, 0.001125127, 0.001139718, 0.001185254, 0.001239235, 
    0.001323538, 0.001486391, 0.001489011, 0.001454965, 0.001827017,
  0.002317294, 0.001776998, 0.001397994, 0.001096426, 0.001064089, 
    0.001130338, 0.00116449, 0.001179067, 0.001237883, 0.001278466, 
    0.001361794, 0.001553543, 0.001735025, 0.001528315, 0.001472588,
  0.002315565, 0.00174034, 0.001285327, 0.001065308, 0.001059695, 
    0.001120517, 0.001207852, 0.001217677, 0.001246427, 0.001283475, 
    0.001362625, 0.001595727, 0.001881753, 0.001928199, 0.00164336,
  0.002376448, 0.00168685, 0.001190006, 0.001060377, 0.001074791, 
    0.001129219, 0.001239163, 0.001249817, 0.001272326, 0.001283139, 
    0.001365865, 0.001581501, 0.00192424, 0.002221371, 0.00198861,
  0.002341127, 0.001643556, 0.00122997, 0.001058908, 0.001073046, 
    0.001170115, 0.00124712, 0.001280236, 0.001300511, 0.001281986, 
    0.001352875, 0.001532073, 0.001831562, 0.002246997, 0.002473737,
  0.002545594, 0.001973592, 0.001334874, 0.001106348, 0.0009596135, 
    0.001036458, 0.001144084, 0.001283406, 0.001305224, 0.001349244, 
    0.001346905, 0.001307174, 0.001403751, 0.001767377, 0.00254773,
  0.002521872, 0.001706239, 0.001282613, 0.001104207, 0.001080704, 
    0.001041221, 0.001252958, 0.00131847, 0.001339242, 0.001195192, 
    0.001314774, 0.001434882, 0.001405521, 0.001607577, 0.002257475,
  0.00234039, 0.001745107, 0.001370355, 0.001193699, 0.001092609, 
    0.001042142, 0.001263085, 0.001406889, 0.001427427, 0.001443578, 
    0.00137303, 0.001548441, 0.001482924, 0.001582883, 0.002204563,
  0.002127491, 0.001648354, 0.00139211, 0.001151705, 0.001156335, 0.00117889, 
    0.001207837, 0.001328975, 0.001382257, 0.001556683, 0.001640862, 
    0.001681907, 0.001580736, 0.001412424, 0.001985078,
  0.001940224, 0.001533414, 0.001345312, 0.00115997, 0.001183195, 
    0.001256459, 0.001330745, 0.001152625, 0.001189043, 0.001593252, 
    0.001855679, 0.001941612, 0.001713806, 0.001305563, 0.001809848,
  0.001823569, 0.001523036, 0.001283528, 0.001161015, 0.001172055, 
    0.001256349, 0.001312617, 0.001367062, 0.001432377, 0.001661927, 
    0.001957875, 0.002090184, 0.001829187, 0.00151951, 0.001664354,
  0.001823901, 0.001522593, 0.001304742, 0.001102851, 0.001173982, 
    0.001239272, 0.001283118, 0.001363279, 0.001451257, 0.001686074, 
    0.002000308, 0.002205826, 0.00194824, 0.001593145, 0.001535404,
  0.001830714, 0.001499363, 0.001235619, 0.001067548, 0.00117606, 
    0.001255796, 0.001265635, 0.001279355, 0.001356204, 0.001580551, 
    0.001920978, 0.00218701, 0.002130589, 0.00170481, 0.001561729,
  0.00188642, 0.001538226, 0.001102449, 0.001057876, 0.001158063, 
    0.001260272, 0.001258052, 0.00126495, 0.001334358, 0.001523204, 
    0.00177858, 0.002085257, 0.002321579, 0.00198175, 0.001505485,
  0.001867031, 0.001427026, 0.001100454, 0.001054694, 0.001147041, 
    0.00124091, 0.001215285, 0.00122684, 0.001260031, 0.001378825, 
    0.001633417, 0.00188525, 0.002225895, 0.002452051, 0.001735073,
  0.001754438, 0.001623175, 0.001374, 0.001190187, 0.001184169, 0.001096533, 
    0.001207395, 0.001313829, 0.001511873, 0.001683138, 0.001825141, 
    0.001850044, 0.001801091, 0.001786592, 0.001792526,
  0.001694921, 0.001495331, 0.00134004, 0.001272886, 0.001247138, 
    0.001175779, 0.001333977, 0.001505283, 0.001662763, 0.001616128, 
    0.001916132, 0.001946086, 0.00187844, 0.001652287, 0.001774404,
  0.001689009, 0.001566485, 0.001423216, 0.001360094, 0.001255261, 
    0.001147688, 0.00137181, 0.001526546, 0.001699106, 0.001925117, 
    0.002028772, 0.001911236, 0.00178589, 0.001695176, 0.002031141,
  0.00159135, 0.001566428, 0.001473104, 0.001354554, 0.001262813, 0.00123712, 
    0.001245872, 0.001403145, 0.00162145, 0.001952306, 0.002063203, 
    0.001781819, 0.001632783, 0.001708499, 0.002409449,
  0.001539334, 0.001518982, 0.001439188, 0.001339688, 0.001266435, 
    0.001251617, 0.001307539, 0.001280674, 0.001405679, 0.001924203, 
    0.002076892, 0.001742901, 0.001667241, 0.001789544, 0.002547764,
  0.001522279, 0.001460436, 0.001336548, 0.001300726, 0.00124962, 
    0.001192917, 0.001320469, 0.001440622, 0.001657228, 0.00189388, 
    0.002067877, 0.001875038, 0.001703861, 0.001768082, 0.002391333,
  0.001514845, 0.001408388, 0.001270613, 0.001238305, 0.001272904, 
    0.001155816, 0.001268135, 0.001455491, 0.001651444, 0.001862697, 
    0.002068417, 0.002176638, 0.00177064, 0.001743314, 0.002168298,
  0.001621736, 0.00143907, 0.001226724, 0.001135665, 0.001281627, 
    0.001139787, 0.001208672, 0.001367887, 0.001490148, 0.001711667, 
    0.00192962, 0.002223822, 0.002102086, 0.001771787, 0.001960519,
  0.001831956, 0.001643232, 0.001225927, 0.001060708, 0.001249847, 
    0.001167831, 0.00115615, 0.001334402, 0.001440742, 0.00163609, 
    0.001743845, 0.002167606, 0.002304062, 0.00195307, 0.001836708,
  0.002013956, 0.001812481, 0.001352715, 0.001098165, 0.001264888, 
    0.001161796, 0.001113571, 0.001299222, 0.001389716, 0.00150288, 
    0.001551488, 0.001868941, 0.002340611, 0.002298365, 0.001861758,
  0.001388551, 0.001505456, 0.001276594, 0.001291201, 0.001247565, 
    0.001217105, 0.001310702, 0.001539989, 0.001687688, 0.001824756, 
    0.002046461, 0.002094951, 0.002059091, 0.002028173, 0.002021491,
  0.001596097, 0.001471848, 0.001383978, 0.001309269, 0.001321911, 
    0.001174316, 0.001272956, 0.001566103, 0.001715528, 0.001962889, 
    0.002194639, 0.002150392, 0.002032161, 0.001755002, 0.00173863,
  0.00150469, 0.001578144, 0.001476404, 0.001295032, 0.001236967, 
    0.001159251, 0.001253647, 0.001435236, 0.001731603, 0.002027756, 
    0.002213765, 0.002221867, 0.00212472, 0.001938474, 0.001890858,
  0.001507211, 0.001557362, 0.001477515, 0.001268299, 0.00122821, 
    0.001128274, 0.00120426, 0.001318271, 0.001575727, 0.001934717, 
    0.002197785, 0.002367454, 0.002209906, 0.002210809, 0.002288174,
  0.001555467, 0.001453196, 0.001427962, 0.001258241, 0.0012242, 0.00120807, 
    0.001356148, 0.001251403, 0.001347575, 0.001865428, 0.002166291, 
    0.002421328, 0.002296819, 0.00233169, 0.002445943,
  0.00169005, 0.00143273, 0.001366832, 0.001274916, 0.001240156, 0.001215507, 
    0.001344181, 0.001482294, 0.001605364, 0.001866956, 0.002108982, 
    0.002429314, 0.002385304, 0.002392491, 0.002523474,
  0.001872012, 0.001511327, 0.001384919, 0.001291914, 0.001274547, 
    0.001233188, 0.001323784, 0.001392436, 0.001539914, 0.001787303, 
    0.0020108, 0.002386874, 0.002442475, 0.002428113, 0.002523311,
  0.002002601, 0.001647045, 0.001549969, 0.001233745, 0.001322917, 
    0.001240794, 0.001328988, 0.001358104, 0.001400416, 0.001604478, 
    0.001830293, 0.002286974, 0.002445864, 0.002440813, 0.002487547,
  0.002184042, 0.002035712, 0.001815891, 0.001270673, 0.001308924, 
    0.001243393, 0.001331362, 0.001332028, 0.001354833, 0.001499181, 
    0.00164946, 0.002106472, 0.002456869, 0.002457601, 0.002443557,
  0.002231391, 0.002170874, 0.00197717, 0.001343492, 0.001321885, 
    0.001233349, 0.001287897, 0.001325112, 0.001351401, 0.001403854, 
    0.001500691, 0.001857982, 0.002420267, 0.002487344, 0.002386904,
  0.001440078, 0.001404061, 0.00132272, 0.001260634, 0.001254234, 0.0012669, 
    0.001396281, 0.001473744, 0.001613952, 0.001790549, 0.001903077, 
    0.002172774, 0.002293942, 0.002268721, 0.002154613,
  0.001697205, 0.001548634, 0.001386146, 0.001249958, 0.001267781, 
    0.001282144, 0.001331414, 0.001351487, 0.001428477, 0.001680937, 
    0.001830138, 0.002077535, 0.002271851, 0.002251128, 0.002278413,
  0.001794402, 0.001552887, 0.001447256, 0.00125272, 0.001243006, 
    0.001193852, 0.001235941, 0.00123386, 0.001411545, 0.001568971, 
    0.001683352, 0.001991133, 0.002264789, 0.002396884, 0.002480916,
  0.001892911, 0.001501484, 0.001449506, 0.001259722, 0.001293118, 
    0.001273225, 0.001214721, 0.001169018, 0.00127399, 0.001449022, 0.001558, 
    0.001880322, 0.002242765, 0.002347331, 0.002425221,
  0.001909934, 0.001525729, 0.001511657, 0.001280192, 0.001308055, 
    0.001269035, 0.001332774, 0.001118805, 0.001134627, 0.001355854, 
    0.001479291, 0.001842478, 0.002253419, 0.002349209, 0.002455231,
  0.001887224, 0.001624256, 0.001572895, 0.001306962, 0.001333907, 
    0.001295337, 0.001310291, 0.001299758, 0.00129189, 0.001305247, 
    0.001435683, 0.001854372, 0.002299951, 0.00243024, 0.002547793,
  0.001829054, 0.001742486, 0.001771572, 0.001351198, 0.001308715, 
    0.001297232, 0.00130253, 0.001300444, 0.001288966, 0.001272883, 
    0.001460197, 0.001879651, 0.002309193, 0.00242779, 0.002384828,
  0.001878253, 0.00181284, 0.001871888, 0.001328798, 0.001287618, 
    0.001361217, 0.001316514, 0.001286053, 0.001285427, 0.001255677, 
    0.001451292, 0.00189804, 0.002278408, 0.002284669, 0.002328118,
  0.00202726, 0.002050986, 0.00202924, 0.001516111, 0.001418155, 0.001350267, 
    0.00133455, 0.001285236, 0.001268694, 0.001288836, 0.001420157, 
    0.001906476, 0.002193102, 0.002066734, 0.002079407,
  0.002125619, 0.002503971, 0.002385214, 0.00198944, 0.001784726, 
    0.001514317, 0.001335777, 0.001305886, 0.001270279, 0.001292226, 
    0.001377489, 0.001901194, 0.002093125, 0.002010829, 0.001936219,
  0.001311359, 0.001511692, 0.001458227, 0.001362395, 0.001336358, 
    0.001272215, 0.001288709, 0.001338776, 0.001264551, 0.001307256, 
    0.001261907, 0.001281035, 0.00147457, 0.001752198, 0.001861808,
  0.001525287, 0.001687084, 0.001611582, 0.001506172, 0.001449068, 
    0.00134374, 0.001293219, 0.001159259, 0.001130683, 0.001189915, 
    0.001233333, 0.001284029, 0.00145974, 0.001762803, 0.001782924,
  0.001702139, 0.001836882, 0.001829605, 0.001704393, 0.001566153, 
    0.001367825, 0.001280494, 0.001276766, 0.00119272, 0.001251529, 
    0.001166938, 0.001315132, 0.001562402, 0.00182436, 0.00188755,
  0.001879156, 0.00199826, 0.0020591, 0.001927633, 0.001900622, 0.001681905, 
    0.00135252, 0.001254537, 0.001219188, 0.001239058, 0.001261161, 
    0.001329522, 0.001571877, 0.001776458, 0.001906984,
  0.002103442, 0.002225493, 0.002384912, 0.002246974, 0.002175655, 
    0.002002321, 0.001713762, 0.001281398, 0.001110848, 0.001232014, 
    0.001251241, 0.001335897, 0.001565512, 0.001773419, 0.001841143,
  0.002293093, 0.002460646, 0.002631168, 0.002509723, 0.002307774, 
    0.002114308, 0.001951856, 0.001749182, 0.001487324, 0.001328981, 
    0.001298853, 0.001387539, 0.001620369, 0.001758499, 0.001828743,
  0.002498336, 0.002635718, 0.002724601, 0.002524015, 0.002224687, 
    0.002027552, 0.002040465, 0.001968179, 0.001739032, 0.001448232, 
    0.00136885, 0.001425295, 0.001683308, 0.001806112, 0.001814256,
  0.002600493, 0.002636755, 0.002660742, 0.002458276, 0.002124839, 
    0.001987939, 0.002037103, 0.002149695, 0.001861939, 0.001529641, 
    0.001367889, 0.001486962, 0.00171596, 0.001838392, 0.001862557,
  0.002581225, 0.002552029, 0.002511112, 0.002334769, 0.002147647, 
    0.001981076, 0.001955638, 0.001931446, 0.001591842, 0.001290013, 
    0.001326679, 0.00154049, 0.001817088, 0.001887657, 0.001942235,
  0.002543729, 0.002509487, 0.002312508, 0.002138451, 0.001979929, 
    0.001777528, 0.001660947, 0.00162785, 0.001370388, 0.001394057, 
    0.001391683, 0.001725423, 0.001962541, 0.001993269, 0.001890307,
  0.001906782, 0.001830231, 0.001864227, 0.001825281, 0.001853968, 
    0.001865446, 0.001810727, 0.001764514, 0.001741763, 0.001664461, 
    0.001522696, 0.001316569, 0.001217773, 0.001273726, 0.001507055,
  0.002470227, 0.002236012, 0.002274169, 0.002246827, 0.002221713, 
    0.002199733, 0.002090932, 0.001999959, 0.001852515, 0.001728073, 
    0.00159012, 0.001371225, 0.001124321, 0.00121067, 0.001311725,
  0.002550818, 0.002525014, 0.002485837, 0.002451391, 0.002498969, 
    0.002390408, 0.002490086, 0.002448282, 0.002278842, 0.002040741, 
    0.001723368, 0.001508642, 0.001181121, 0.001235579, 0.001304064,
  0.002543184, 0.002455402, 0.002355102, 0.002255727, 0.002208402, 
    0.002259207, 0.002158771, 0.002309873, 0.002315689, 0.002342709, 
    0.002132752, 0.001761269, 0.001300844, 0.001233181, 0.001256708,
  0.002404244, 0.002287747, 0.002097333, 0.001916755, 0.00183701, 
    0.001804136, 0.001835205, 0.001680505, 0.001635747, 0.002111934, 
    0.002208162, 0.001945984, 0.001398198, 0.001219218, 0.001165676,
  0.002211533, 0.002022807, 0.001806864, 0.001686313, 0.001641887, 
    0.001574242, 0.001566156, 0.001674359, 0.001682647, 0.001717551, 
    0.002005524, 0.001981422, 0.001568055, 0.001251668, 0.001207848,
  0.002044145, 0.001853331, 0.001681904, 0.001667564, 0.001673401, 
    0.001668886, 0.001635688, 0.001769842, 0.001850759, 0.001860693, 
    0.001943173, 0.001928721, 0.001606075, 0.001352899, 0.001358152,
  0.001989601, 0.001854166, 0.001696965, 0.00168173, 0.001719844, 
    0.001809451, 0.001838609, 0.001839659, 0.001848031, 0.002045308, 
    0.001977653, 0.001873197, 0.001622894, 0.001456255, 0.001369423,
  0.0020127, 0.001874682, 0.001680608, 0.001711951, 0.001804484, 0.001952731, 
    0.00203989, 0.001860971, 0.001699882, 0.001805551, 0.00199973, 
    0.001812335, 0.001614138, 0.001455109, 0.001461051,
  0.002031485, 0.001808722, 0.001707896, 0.001744129, 0.001855318, 
    0.002058005, 0.002190574, 0.002103554, 0.001763923, 0.001667017, 
    0.001870482, 0.001765646, 0.001592329, 0.0014772, 0.001516607,
  0.00200172, 0.001953771, 0.002029005, 0.001767777, 0.001626447, 
    0.001569257, 0.00166801, 0.00184507, 0.00172704, 0.00158777, 0.001632718, 
    0.001591914, 0.001370718, 0.001223088, 0.001308082,
  0.002237373, 0.002233316, 0.002124147, 0.002004982, 0.001938686, 
    0.001873392, 0.001861463, 0.001948738, 0.001933177, 0.001720536, 
    0.001686775, 0.001716178, 0.001519041, 0.001256585, 0.001249344,
  0.00249395, 0.002510954, 0.002467394, 0.002262686, 0.00208086, 0.001809851, 
    0.001650498, 0.001693147, 0.001919956, 0.002002852, 0.001830022, 
    0.001827996, 0.001643469, 0.00139585, 0.001295497,
  0.002576485, 0.002561276, 0.002532324, 0.002420996, 0.002253534, 
    0.002041241, 0.001546665, 0.00141987, 0.001381034, 0.001875237, 
    0.001996502, 0.002001997, 0.001825994, 0.001533563, 0.001322734,
  0.002618742, 0.002530977, 0.002380219, 0.002344699, 0.002099684, 
    0.002044635, 0.001855113, 0.001413723, 0.001158478, 0.001331658, 
    0.002030829, 0.002160708, 0.001930147, 0.001662611, 0.001179442,
  0.002561791, 0.002356553, 0.002160701, 0.00188873, 0.001792006, 
    0.001787652, 0.001947663, 0.001840536, 0.001488342, 0.001346414, 
    0.001920773, 0.002274311, 0.002061842, 0.001543, 0.001366846,
  0.002395535, 0.002200241, 0.001908767, 0.001806692, 0.001813824, 
    0.001975658, 0.002109727, 0.002149805, 0.001909147, 0.001458367, 
    0.001723835, 0.00228295, 0.002047526, 0.001544554, 0.001597816,
  0.002284847, 0.002074895, 0.001840017, 0.001883482, 0.002047171, 
    0.002165333, 0.002147694, 0.00211743, 0.001960456, 0.001732269, 
    0.001704475, 0.002269149, 0.0019473, 0.001542883, 0.001551463,
  0.002186301, 0.002025059, 0.001935925, 0.001992344, 0.002137063, 
    0.002115067, 0.002242164, 0.002164955, 0.001975255, 0.001697372, 
    0.00176974, 0.002200078, 0.001770945, 0.001545463, 0.001493711,
  0.002126352, 0.001963023, 0.002002775, 0.002116185, 0.002233787, 
    0.002306802, 0.002250907, 0.002147868, 0.001765297, 0.001695851, 
    0.001965204, 0.002092794, 0.001618871, 0.001515768, 0.001480387,
  0.002731265, 0.002619199, 0.00263968, 0.002519478, 0.002236102, 0.00195299, 
    0.001874754, 0.001849145, 0.001893126, 0.00202457, 0.001927974, 
    0.001666776, 0.001539113, 0.001456468, 0.001644586,
  0.002960655, 0.00272424, 0.002610682, 0.002662415, 0.002593947, 
    0.002490932, 0.002214093, 0.001901004, 0.001886526, 0.00208364, 
    0.002048323, 0.001818138, 0.001510742, 0.001267347, 0.001452964,
  0.003198608, 0.003175918, 0.003037738, 0.002987043, 0.002917289, 
    0.002624895, 0.002518019, 0.00225779, 0.001911123, 0.002103854, 
    0.002028234, 0.001878573, 0.001642326, 0.001347431, 0.001410164,
  0.002946944, 0.002825385, 0.002719252, 0.00272666, 0.002665004, 0.00278169, 
    0.002454627, 0.002354852, 0.001893426, 0.001930105, 0.001973178, 
    0.001850693, 0.001662808, 0.00138484, 0.001279752,
  0.002617569, 0.002386675, 0.002201091, 0.002305317, 0.001915307, 
    0.002107133, 0.002107263, 0.002053159, 0.001642778, 0.001794343, 
    0.001996579, 0.001837902, 0.001653077, 0.00143253, 0.001312066,
  0.002319793, 0.002195982, 0.002099389, 0.002054803, 0.001840425, 
    0.001515008, 0.002044375, 0.002101025, 0.001778027, 0.001713395, 
    0.001830231, 0.001825617, 0.001701485, 0.001427539, 0.00134647,
  0.002157904, 0.002089851, 0.001952455, 0.002117065, 0.001922829, 
    0.001631423, 0.001943081, 0.002041942, 0.001814238, 0.001739082, 
    0.001830707, 0.0018107, 0.001676798, 0.001491188, 0.001694851,
  0.002028905, 0.001978681, 0.001971716, 0.002020248, 0.002012055, 
    0.00194497, 0.001873905, 0.002039815, 0.001792559, 0.001751006, 
    0.001808643, 0.001819496, 0.001677641, 0.00161861, 0.001677964,
  0.00195167, 0.001961101, 0.001946871, 0.001892772, 0.002080162, 
    0.001929267, 0.002037975, 0.001975434, 0.001852239, 0.001742325, 
    0.001807627, 0.001842809, 0.001647659, 0.001604913, 0.001611027,
  0.00191601, 0.001951924, 0.001999406, 0.00198842, 0.001963122, 0.001998028, 
    0.001992024, 0.001959434, 0.001821324, 0.001747878, 0.001881635, 
    0.001848942, 0.001635688, 0.001574872, 0.001605632,
  0.002824596, 0.002573733, 0.002592213, 0.002692037, 0.002734389, 
    0.002520383, 0.002259867, 0.002266794, 0.00218491, 0.002190778, 
    0.001882776, 0.001689413, 0.00200946, 0.002151057, 0.002507075,
  0.003199606, 0.002936634, 0.002756564, 0.002942208, 0.002861652, 
    0.002558805, 0.002414187, 0.002236443, 0.001975478, 0.00187499, 
    0.002048989, 0.001773953, 0.001938576, 0.002001511, 0.002398997,
  0.003441923, 0.003343159, 0.003145196, 0.002723549, 0.002625641, 
    0.002444801, 0.002471843, 0.002277846, 0.002046126, 0.002051213, 
    0.002029652, 0.001759975, 0.001947656, 0.00198182, 0.002221292,
  0.002610645, 0.002536662, 0.002436037, 0.002446767, 0.00243902, 
    0.002585121, 0.002511439, 0.00247233, 0.002091985, 0.002147483, 
    0.001972159, 0.001719445, 0.00180455, 0.001891874, 0.002044271,
  0.002351731, 0.002292547, 0.002247797, 0.002473661, 0.002399371, 
    0.002445709, 0.002693755, 0.002238276, 0.001999887, 0.002083178, 
    0.001908812, 0.001780669, 0.001791784, 0.001859206, 0.002003899,
  0.002046726, 0.001985728, 0.001976926, 0.002180671, 0.002174712, 
    0.00183328, 0.002291204, 0.002545824, 0.002166771, 0.00209962, 
    0.001930225, 0.001727331, 0.00176472, 0.001803013, 0.002003407,
  0.001920014, 0.001820943, 0.001740584, 0.001892946, 0.002086407, 
    0.00183547, 0.00178869, 0.002454577, 0.002281629, 0.002067549, 
    0.001903546, 0.001711991, 0.001707649, 0.001881421, 0.001961573,
  0.001823191, 0.001740749, 0.001642041, 0.001795958, 0.002035643, 
    0.001828307, 0.001761536, 0.002321171, 0.002210373, 0.001957784, 
    0.001808365, 0.001665178, 0.001736474, 0.001848949, 0.001890999,
  0.001829254, 0.001859679, 0.001954539, 0.001948118, 0.001984794, 
    0.001853217, 0.002106452, 0.002318311, 0.002187463, 0.001864065, 
    0.001697455, 0.001633953, 0.001699718, 0.001756869, 0.001755886,
  0.0018634, 0.001913692, 0.00201083, 0.00201487, 0.002019849, 0.002095333, 
    0.002229255, 0.002247765, 0.002009658, 0.001758338, 0.001578032, 
    0.001581961, 0.001652751, 0.001621688, 0.001636288,
  0.002734944, 0.002676569, 0.002596698, 0.002664851, 0.002596716, 
    0.00242672, 0.002423208, 0.002638163, 0.002704879, 0.002600323, 
    0.002204874, 0.002097062, 0.002040705, 0.002049474, 0.002427476,
  0.003204499, 0.003033279, 0.002763306, 0.002761211, 0.002848053, 
    0.002602069, 0.002586406, 0.002654612, 0.002547096, 0.002381089, 
    0.002174214, 0.002051754, 0.002043383, 0.002191209, 0.002630858,
  0.003504223, 0.003432278, 0.003231781, 0.002699608, 0.002846774, 
    0.002297511, 0.002281255, 0.002369333, 0.002331894, 0.002227363, 
    0.001920792, 0.001919304, 0.002035157, 0.002383599, 0.002859922,
  0.002526416, 0.00254034, 0.002560595, 0.002528345, 0.002278156, 
    0.002301725, 0.002295151, 0.002161909, 0.00224657, 0.001979527, 
    0.001743094, 0.001795896, 0.002215204, 0.00260838, 0.002941728,
  0.002311178, 0.002279616, 0.002205046, 0.002421451, 0.00218344, 
    0.002299107, 0.002477921, 0.001890256, 0.001664512, 0.002033034, 
    0.0018176, 0.00209548, 0.002455124, 0.002789532, 0.002835104,
  0.002096906, 0.001969527, 0.0019408, 0.002130298, 0.002099616, 0.002099564, 
    0.002310376, 0.00207697, 0.001923933, 0.001880943, 0.001938638, 
    0.002358107, 0.002685306, 0.002781934, 0.002691064,
  0.001948626, 0.001812294, 0.001730975, 0.001905898, 0.002002438, 
    0.002043153, 0.002466943, 0.002230457, 0.002043319, 0.002079967, 
    0.002304673, 0.002584951, 0.002683759, 0.00268583, 0.002586325,
  0.001826928, 0.001719858, 0.001598315, 0.0017712, 0.002019831, 0.002132558, 
    0.002406639, 0.002317656, 0.002065063, 0.002195147, 0.002353643, 
    0.002508462, 0.002531963, 0.002454016, 0.002382868,
  0.001769534, 0.001841331, 0.00192443, 0.001909037, 0.002004003, 
    0.002179477, 0.002392738, 0.002226323, 0.002050382, 0.002107662, 
    0.002217878, 0.002355136, 0.002332712, 0.002291068, 0.002237295,
  0.001806281, 0.00189857, 0.00200195, 0.00201909, 0.002199989, 0.002293164, 
    0.002284325, 0.00208571, 0.001955686, 0.001967445, 0.002048206, 
    0.002114446, 0.002144661, 0.002136238, 0.002143058,
  0.003391913, 0.003078708, 0.002851414, 0.002973518, 0.002713574, 
    0.002793904, 0.002875512, 0.002813631, 0.002607765, 0.002508506, 
    0.002440069, 0.002498238, 0.002491093, 0.00233314, 0.002199048,
  0.003254837, 0.002871041, 0.002800258, 0.00278551, 0.00293335, 0.002925461, 
    0.002913898, 0.00281304, 0.002640944, 0.002614526, 0.002482193, 
    0.002566846, 0.002550289, 0.002263231, 0.002165418,
  0.003332175, 0.003168056, 0.003175384, 0.002829632, 0.002795817, 
    0.002171393, 0.00221543, 0.002330012, 0.002378163, 0.002346016, 
    0.00232464, 0.002469276, 0.002385431, 0.002179815, 0.002065124,
  0.002678859, 0.0025674, 0.00262425, 0.00278924, 0.002198262, 0.00217991, 
    0.001940771, 0.00193085, 0.002115678, 0.002310389, 0.002289619, 
    0.002322193, 0.002192558, 0.002157916, 0.002268657,
  0.002474341, 0.002504354, 0.002360073, 0.002253168, 0.001842857, 
    0.001903843, 0.001974195, 0.001725778, 0.001586954, 0.001836259, 
    0.002135439, 0.002137106, 0.002117351, 0.002162529, 0.002445225,
  0.002437293, 0.002178502, 0.002020857, 0.001985265, 0.001779541, 
    0.001866331, 0.001947757, 0.001875028, 0.002005376, 0.001845015, 
    0.001909974, 0.002120088, 0.00223856, 0.002499665, 0.002472577,
  0.002090647, 0.001977775, 0.001675646, 0.001896504, 0.001903741, 
    0.001984758, 0.002083124, 0.001972543, 0.002132751, 0.002194581, 
    0.002311186, 0.002438062, 0.002546408, 0.002511389, 0.002398413,
  0.001922684, 0.001837944, 0.001723551, 0.001956762, 0.0020645, 0.002232926, 
    0.002142491, 0.00207448, 0.00215654, 0.002394115, 0.002545159, 
    0.002590794, 0.002514793, 0.002323573, 0.002214138,
  0.001837051, 0.001915672, 0.001953477, 0.002033751, 0.002123364, 
    0.002181084, 0.002186187, 0.002231851, 0.002372328, 0.002615398, 
    0.002626361, 0.002504725, 0.002357894, 0.00225863, 0.002295586,
  0.001874138, 0.001962027, 0.002091979, 0.002137359, 0.002175625, 
    0.002231944, 0.002264365, 0.002425315, 0.002594329, 0.002543672, 
    0.002432246, 0.002340466, 0.002284741, 0.00234398, 0.002435311,
  0.003531136, 0.00321705, 0.002984217, 0.002831341, 0.002750177, 
    0.002730081, 0.002613311, 0.002532524, 0.002407073, 0.002394612, 
    0.002480321, 0.002156527, 0.002218322, 0.002181174, 0.002158443,
  0.003360159, 0.003104165, 0.002977428, 0.00283891, 0.002771107, 
    0.002787609, 0.002598628, 0.002481026, 0.002362166, 0.002408199, 
    0.002516364, 0.002394935, 0.002227834, 0.002196421, 0.001966532,
  0.003553107, 0.003385102, 0.003206841, 0.003007474, 0.00278242, 
    0.002285813, 0.002143886, 0.002020833, 0.002059803, 0.002159778, 
    0.002282287, 0.002493079, 0.002429808, 0.002138785, 0.002095814,
  0.003550994, 0.00317796, 0.003068236, 0.002906023, 0.0025497, 0.002181162, 
    0.001662799, 0.001637521, 0.001664653, 0.00178161, 0.002109147, 
    0.002427822, 0.002527791, 0.002402748, 0.002245904,
  0.00335608, 0.003198749, 0.00301792, 0.002616455, 0.002098302, 0.001961374, 
    0.001830122, 0.001664311, 0.001333841, 0.001652872, 0.001940208, 
    0.002248809, 0.002506145, 0.002306556, 0.002161145,
  0.003063365, 0.002721605, 0.0024776, 0.002286443, 0.00198719, 0.002007678, 
    0.002042573, 0.001966382, 0.001834775, 0.001649729, 0.001788494, 
    0.001939687, 0.002203152, 0.002276729, 0.002267129,
  0.00251198, 0.002247629, 0.002165582, 0.002006088, 0.001952784, 
    0.002063211, 0.002083174, 0.002031934, 0.00210335, 0.001886, 0.00193038, 
    0.002125052, 0.002260752, 0.002180371, 0.002157247,
  0.002116586, 0.001947662, 0.001997052, 0.001977195, 0.002086469, 
    0.002110714, 0.001993877, 0.002037999, 0.001881658, 0.0017839, 
    0.00192912, 0.002085232, 0.002123077, 0.002074165, 0.002084632,
  0.001886245, 0.001963888, 0.002051824, 0.002098551, 0.002221064, 
    0.001984169, 0.001990326, 0.001963626, 0.002050078, 0.001989295, 
    0.001836957, 0.002067347, 0.002088835, 0.00204747, 0.002061815,
  0.001918517, 0.002051726, 0.002057036, 0.002246133, 0.002160162, 
    0.002384724, 0.002247503, 0.002289043, 0.002216695, 0.002085817, 
    0.002010845, 0.002072966, 0.002067962, 0.002051473, 0.002100481,
  0.004959674, 0.004561756, 0.004189422, 0.004137703, 0.004001113, 
    0.003866927, 0.003680406, 0.003508057, 0.003311618, 0.003124717, 
    0.002957867, 0.002721703, 0.002585319, 0.002464193, 0.002292778,
  0.004237161, 0.004242615, 0.004126579, 0.00405054, 0.004093833, 
    0.003778156, 0.003614246, 0.003414956, 0.003186044, 0.002910224, 
    0.002728421, 0.002462743, 0.002416602, 0.002259146, 0.002062888,
  0.004337595, 0.004214833, 0.004119747, 0.004017307, 0.003793592, 
    0.003493165, 0.003140354, 0.002962394, 0.002782914, 0.002538878, 
    0.002375202, 0.002242532, 0.002309451, 0.00221965, 0.002219553,
  0.004433058, 0.004305761, 0.004050106, 0.003764012, 0.003527277, 
    0.003134392, 0.002476783, 0.002490696, 0.002390817, 0.00224439, 
    0.002192059, 0.002059411, 0.002052349, 0.002250432, 0.002200806,
  0.004334421, 0.003946872, 0.003673169, 0.003257334, 0.002891787, 
    0.002546321, 0.002234375, 0.001970866, 0.001769884, 0.002033701, 
    0.001840028, 0.00179151, 0.001894787, 0.002179377, 0.002258763,
  0.003533775, 0.003359257, 0.003072273, 0.002752913, 0.002418095, 
    0.002213818, 0.002049811, 0.002019951, 0.001990389, 0.001909556, 
    0.001789449, 0.001875394, 0.002012091, 0.002199575, 0.00229976,
  0.003082713, 0.002918495, 0.002754851, 0.002329799, 0.0021746, 0.002101423, 
    0.002006616, 0.001969388, 0.001926296, 0.001860251, 0.001696602, 
    0.001800261, 0.002198636, 0.002299677, 0.002319966,
  0.002660815, 0.002557287, 0.002472941, 0.002170375, 0.002073016, 
    0.002170706, 0.001989474, 0.001949895, 0.001861398, 0.001881193, 
    0.001828525, 0.00205768, 0.0022797, 0.002340186, 0.002196321,
  0.002420616, 0.002308698, 0.002328857, 0.002152261, 0.002246598, 
    0.002064756, 0.00196754, 0.001893784, 0.001817596, 0.001789706, 
    0.001911324, 0.002001267, 0.002080275, 0.001970814, 0.001833236,
  0.002284222, 0.002225419, 0.002261413, 0.002304624, 0.002110266, 
    0.002056317, 0.001963242, 0.001883958, 0.001791237, 0.00179798, 
    0.001834584, 0.001825008, 0.00186587, 0.001889344, 0.001791963,
  0.002871404, 0.003009218, 0.003090433, 0.003195695, 0.003332098, 
    0.003444728, 0.003515763, 0.003617904, 0.003697127, 0.003737071, 
    0.003788857, 0.003794538, 0.003834636, 0.003718592, 0.00360619,
  0.00308782, 0.002999297, 0.003050629, 0.003257009, 0.003457591, 
    0.003547277, 0.003631682, 0.00369851, 0.00374244, 0.003788386, 
    0.003825273, 0.003834197, 0.003769991, 0.003595484, 0.003449925,
  0.002912948, 0.002911244, 0.00309582, 0.003355165, 0.003550736, 
    0.003594583, 0.003602111, 0.00322915, 0.003286134, 0.003388281, 
    0.00347593, 0.00354103, 0.003513319, 0.00341593, 0.003268068,
  0.002764647, 0.002927485, 0.003128518, 0.003285419, 0.003378775, 
    0.003302019, 0.002635228, 0.002609214, 0.002673659, 0.002902573, 
    0.002978899, 0.003106391, 0.003187902, 0.003112479, 0.002937182,
  0.002662622, 0.002784583, 0.002840529, 0.002755682, 0.002656622, 
    0.002576087, 0.002343288, 0.00213813, 0.002084834, 0.002573227, 
    0.002685253, 0.002748575, 0.002810586, 0.002775377, 0.002643337,
  0.00246574, 0.002451628, 0.0024006, 0.002279837, 0.002180122, 0.002133803, 
    0.002128458, 0.002221185, 0.002296062, 0.002362117, 0.002437869, 
    0.002473982, 0.002491581, 0.002477647, 0.00241156,
  0.00228001, 0.00228056, 0.002107463, 0.00202306, 0.001984037, 0.00195409, 
    0.001930489, 0.001957913, 0.002041458, 0.002185332, 0.002247502, 
    0.002252835, 0.00227235, 0.002267234, 0.002230168,
  0.002188874, 0.002122457, 0.001945798, 0.001944703, 0.001920967, 0.0019863, 
    0.001975819, 0.001975637, 0.001966314, 0.001997265, 0.002151529, 
    0.002156111, 0.002181153, 0.002160901, 0.002044022,
  0.002097467, 0.002008321, 0.001796096, 0.001774511, 0.001771384, 
    0.001827012, 0.001905724, 0.001993373, 0.002046649, 0.002113397, 
    0.002142394, 0.002196164, 0.002133088, 0.002079467, 0.00199634,
  0.002014015, 0.001896868, 0.001793839, 0.001752328, 0.001723169, 
    0.001721659, 0.001765844, 0.001886143, 0.001937422, 0.002063683, 
    0.002133004, 0.002170175, 0.002046812, 0.002064807, 0.002240119,
  0.003036485, 0.002960595, 0.002712046, 0.002496848, 0.002596266, 
    0.002620983, 0.00255431, 0.002288973, 0.00225708, 0.002417391, 
    0.002624766, 0.002790074, 0.002955321, 0.003088265, 0.003267163,
  0.003236259, 0.002882221, 0.002590109, 0.002446299, 0.002524889, 
    0.002384384, 0.002314241, 0.002133378, 0.002094308, 0.002228135, 
    0.00247005, 0.002738438, 0.002959603, 0.00312862, 0.003358426,
  0.00321478, 0.002833379, 0.00252995, 0.002381035, 0.002360302, 0.002130867, 
    0.002139947, 0.001995057, 0.001950353, 0.002065517, 0.002227075, 
    0.002567488, 0.002913305, 0.003271034, 0.003488355,
  0.003232092, 0.002788051, 0.002456238, 0.002385881, 0.002212103, 
    0.002140306, 0.001871932, 0.001834277, 0.001868541, 0.002013305, 
    0.002111823, 0.002433856, 0.002904205, 0.003367217, 0.003574556,
  0.002936405, 0.00248336, 0.002305601, 0.002280927, 0.002071444, 
    0.001961399, 0.001996963, 0.001830009, 0.001762119, 0.001982777, 
    0.002022027, 0.002321729, 0.002859123, 0.003384472, 0.003613438,
  0.002505494, 0.002197164, 0.002048425, 0.002121851, 0.001935948, 
    0.001907858, 0.002075926, 0.002191115, 0.002198694, 0.002089853, 
    0.001952639, 0.002298989, 0.002760999, 0.003120102, 0.003407759,
  0.002242049, 0.002027906, 0.001795915, 0.001826082, 0.001791091, 
    0.001826857, 0.001838898, 0.002094347, 0.002117237, 0.002084207, 
    0.001934915, 0.002318327, 0.002731356, 0.002907516, 0.003032737,
  0.002135522, 0.001941503, 0.001647382, 0.001565415, 0.001602057, 
    0.001674689, 0.001756949, 0.00194282, 0.002041024, 0.001906729, 
    0.001917337, 0.002363391, 0.002728704, 0.002764583, 0.002736981,
  0.002167732, 0.001820542, 0.001523432, 0.001562913, 0.001624264, 
    0.001691911, 0.001773907, 0.001910418, 0.001927584, 0.001872828, 
    0.001905477, 0.00237626, 0.00270361, 0.002766082, 0.002663642,
  0.00209949, 0.001694227, 0.001560377, 0.001682605, 0.001787669, 
    0.001755042, 0.001756955, 0.001868758, 0.001807456, 0.001773068, 
    0.00196746, 0.002460742, 0.002651273, 0.00278475, 0.002697166,
  0.002573714, 0.00284328, 0.003044419, 0.003178172, 0.00329392, 0.003357753, 
    0.003310783, 0.003101841, 0.002825846, 0.002613286, 0.002343944, 
    0.002158509, 0.002037704, 0.001875845, 0.001874504,
  0.002836562, 0.002865471, 0.003032455, 0.003197944, 0.003354081, 
    0.003352409, 0.003270859, 0.002934209, 0.002639829, 0.002365935, 
    0.002229192, 0.002105698, 0.0018637, 0.001796615, 0.00191041,
  0.002812607, 0.002856326, 0.002989712, 0.003106394, 0.003230453, 
    0.003024355, 0.002908268, 0.002595616, 0.002378886, 0.002186799, 
    0.002101387, 0.002008836, 0.001823678, 0.001907076, 0.002312079,
  0.002739505, 0.002712792, 0.002826351, 0.002874346, 0.002854664, 
    0.002635809, 0.002296978, 0.002336806, 0.002176974, 0.002065359, 
    0.001941077, 0.00181975, 0.00185153, 0.002305985, 0.002839345,
  0.002534883, 0.002404668, 0.002466304, 0.002401675, 0.002450099, 
    0.002380461, 0.002203726, 0.001807877, 0.001693291, 0.001907015, 
    0.001789239, 0.001758428, 0.002147626, 0.002803797, 0.003399314,
  0.002420977, 0.002165508, 0.002091216, 0.002021186, 0.002082887, 
    0.002121782, 0.002101845, 0.002005251, 0.001898291, 0.001852338, 
    0.001841392, 0.002056704, 0.002575017, 0.003225514, 0.003623799,
  0.002320967, 0.001949372, 0.001794892, 0.001808851, 0.00177855, 
    0.001763941, 0.001805944, 0.001809184, 0.001755951, 0.001810857, 
    0.001873021, 0.002425211, 0.002817526, 0.003344471, 0.003621182,
  0.002235171, 0.001861281, 0.001613803, 0.001645465, 0.001613996, 
    0.001594708, 0.001655069, 0.001735177, 0.001794049, 0.001816614, 
    0.002150044, 0.00265568, 0.002889959, 0.003079507, 0.003232169,
  0.002290579, 0.001949125, 0.001708159, 0.001730622, 0.001745449, 
    0.001772116, 0.001744097, 0.001721105, 0.001810631, 0.001989743, 
    0.002442425, 0.002900854, 0.002877439, 0.002907173, 0.002880882,
  0.002360272, 0.00214057, 0.002051874, 0.002088235, 0.002063059, 
    0.001723967, 0.001780219, 0.001865612, 0.001789729, 0.002072513, 
    0.002658308, 0.002786209, 0.002667798, 0.002578195, 0.002496309,
  0.002418474, 0.002757654, 0.002750803, 0.002235527, 0.002049491, 
    0.002140473, 0.002310459, 0.002623141, 0.002933291, 0.003144855, 
    0.00321737, 0.002943604, 0.002757254, 0.002550314, 0.002466793,
  0.003080705, 0.002978142, 0.002645446, 0.00203655, 0.001942358, 
    0.002022705, 0.002150564, 0.002420021, 0.002707676, 0.002838474, 
    0.002781389, 0.002645891, 0.002469671, 0.002290667, 0.002194968,
  0.003361106, 0.003079877, 0.002504826, 0.001926088, 0.001834176, 
    0.001947145, 0.001986661, 0.002159609, 0.002349169, 0.002486279, 
    0.002431355, 0.002345336, 0.002219306, 0.00215918, 0.00221612,
  0.003657049, 0.003192865, 0.002416593, 0.001834276, 0.001778582, 
    0.001977774, 0.001885387, 0.001953651, 0.002105386, 0.002361627, 
    0.002420821, 0.002350674, 0.002262287, 0.002275012, 0.002460032,
  0.003821093, 0.003131284, 0.002374048, 0.001762521, 0.001751461, 
    0.001885568, 0.001952163, 0.001751638, 0.001800817, 0.002375476, 
    0.002500708, 0.002603076, 0.002744845, 0.003007339, 0.003346464,
  0.003646143, 0.003158202, 0.002442162, 0.001949837, 0.00181507, 
    0.001802343, 0.001877745, 0.001971564, 0.002069298, 0.00239092, 
    0.002557351, 0.002750125, 0.003096333, 0.003473622, 0.003522421,
  0.003090973, 0.002944192, 0.002694549, 0.002313792, 0.002012052, 
    0.001863096, 0.001807908, 0.001914411, 0.002039065, 0.002442828, 
    0.002703075, 0.002868321, 0.00326316, 0.003552625, 0.003593133,
  0.003007893, 0.002940309, 0.002903856, 0.00263641, 0.002335757, 
    0.001980274, 0.001823903, 0.00192589, 0.002023546, 0.002339556, 
    0.002677063, 0.002881281, 0.003236926, 0.003509584, 0.003474351,
  0.002703535, 0.002703639, 0.00283423, 0.002780547, 0.002589434, 
    0.002152262, 0.001899893, 0.002034523, 0.002058484, 0.002330167, 
    0.002656244, 0.002821025, 0.003009475, 0.003103015, 0.003070511,
  0.002554796, 0.002575903, 0.002547175, 0.00258774, 0.002670499, 0.00233974, 
    0.002075366, 0.002036885, 0.002035749, 0.002340244, 0.002556516, 
    0.002499107, 0.002538446, 0.002674597, 0.002661488,
  0.002710751, 0.002951732, 0.003104002, 0.002889334, 0.002125857, 
    0.001695266, 0.001580208, 0.001885345, 0.002300781, 0.002803326, 
    0.003083937, 0.003109811, 0.003032975, 0.002937348, 0.002943339,
  0.003253463, 0.003268241, 0.003180719, 0.002629034, 0.002033367, 
    0.001657507, 0.00155013, 0.001842325, 0.002157208, 0.002874146, 
    0.003180349, 0.003208359, 0.003104038, 0.002968894, 0.003044778,
  0.003570339, 0.003360891, 0.002972529, 0.002367876, 0.001858263, 
    0.001656684, 0.001621183, 0.001766025, 0.002097559, 0.00277953, 
    0.003129342, 0.003330385, 0.003252276, 0.003214041, 0.003203623,
  0.003941755, 0.003504055, 0.002898637, 0.002275631, 0.001674337, 
    0.00168706, 0.001686209, 0.001730392, 0.001944963, 0.002532874, 
    0.003006456, 0.003356806, 0.003351429, 0.003287336, 0.003224224,
  0.003779327, 0.003562752, 0.003133258, 0.002353411, 0.001907647, 
    0.001866546, 0.001882688, 0.001720623, 0.0017521, 0.002376553, 
    0.002883156, 0.003292551, 0.003299107, 0.003178626, 0.00308579,
  0.003124209, 0.003199336, 0.003373412, 0.002887908, 0.002432037, 
    0.002148918, 0.002068734, 0.002088851, 0.002015017, 0.00238474, 
    0.002821827, 0.003186997, 0.003188532, 0.003002964, 0.00291268,
  0.002688199, 0.002604238, 0.003074434, 0.003054723, 0.002930712, 
    0.00276664, 0.002600995, 0.002246226, 0.001972966, 0.002338246, 
    0.002759867, 0.003029335, 0.003037256, 0.002880418, 0.002814291,
  0.002780729, 0.002772294, 0.002673182, 0.002715526, 0.002736546, 
    0.003059311, 0.0028724, 0.002119358, 0.001990968, 0.002265603, 
    0.002657857, 0.002851111, 0.002861559, 0.002784917, 0.002804552,
  0.002494816, 0.00227766, 0.002418784, 0.002559683, 0.002678508, 0.00297775, 
    0.002576107, 0.002093187, 0.001998374, 0.002172098, 0.002643651, 
    0.002737991, 0.002757816, 0.002769265, 0.00286738,
  0.00239171, 0.002197917, 0.002373899, 0.002556996, 0.002608607, 
    0.002673414, 0.002284388, 0.002001127, 0.001976922, 0.002175828, 
    0.002589823, 0.002659172, 0.002750507, 0.002824224, 0.002918272,
  0.003265034, 0.002980269, 0.002780332, 0.002376633, 0.002042274, 
    0.00185576, 0.001690286, 0.00166534, 0.00194005, 0.002469371, 
    0.002816829, 0.002988331, 0.00296519, 0.00287344, 0.002909556,
  0.003112296, 0.002873871, 0.002583227, 0.002273401, 0.002058994, 
    0.001848033, 0.001720753, 0.001717787, 0.001782079, 0.002372779, 
    0.002758482, 0.002941702, 0.002966673, 0.002768767, 0.002767349,
  0.003069937, 0.002822377, 0.002583559, 0.002327859, 0.002089329, 
    0.001909353, 0.001892041, 0.001971241, 0.001844812, 0.002325921, 
    0.00273264, 0.002936862, 0.003004249, 0.002892104, 0.002854384,
  0.003051797, 0.0027369, 0.002512722, 0.002338189, 0.002021871, 0.002092227, 
    0.002034748, 0.001991373, 0.001949682, 0.002321465, 0.002730877, 
    0.002948167, 0.003065316, 0.003030465, 0.002959403,
  0.002891892, 0.002565102, 0.002456974, 0.002587033, 0.002146845, 
    0.002252596, 0.002338309, 0.001952935, 0.001860259, 0.002298156, 
    0.002740274, 0.00294346, 0.003125679, 0.003175161, 0.003163982,
  0.002851636, 0.002790059, 0.002731506, 0.00284178, 0.00280624, 0.002545942, 
    0.002388739, 0.002328486, 0.002306153, 0.002469436, 0.002759886, 
    0.002971173, 0.003187539, 0.003311363, 0.00337779,
  0.002676947, 0.002541467, 0.002447708, 0.002486606, 0.002532179, 
    0.002520903, 0.002439327, 0.002277919, 0.002335442, 0.002521435, 
    0.002693038, 0.002939893, 0.003230914, 0.003388482, 0.003454695,
  0.002615896, 0.002452395, 0.00229231, 0.002336269, 0.002263836, 
    0.002300979, 0.00227474, 0.002392534, 0.00246663, 0.002468599, 
    0.002707275, 0.003024542, 0.003292036, 0.003389986, 0.003426751,
  0.002530542, 0.002384949, 0.002293798, 0.00226228, 0.002216947, 
    0.002167653, 0.002254795, 0.002383888, 0.002503956, 0.002493916, 
    0.002708562, 0.003092132, 0.003347592, 0.003364993, 0.003369103,
  0.002487239, 0.002289496, 0.002170341, 0.002113475, 0.002103643, 
    0.002147322, 0.002249257, 0.002353961, 0.002407038, 0.002499379, 
    0.002719104, 0.003153334, 0.003385012, 0.003413421, 0.003369755,
  0.002207838, 0.002449317, 0.002341141, 0.002248066, 0.002181201, 
    0.002024016, 0.001978991, 0.002070284, 0.002298067, 0.002508626, 
    0.002763843, 0.002998057, 0.003151234, 0.003039989, 0.003076684,
  0.002515745, 0.002513797, 0.002376181, 0.00230853, 0.00220692, 0.002132029, 
    0.002091375, 0.002207581, 0.002290531, 0.002528305, 0.002798982, 
    0.003089727, 0.003149147, 0.002998833, 0.003064496,
  0.00262854, 0.002543915, 0.002362828, 0.002211583, 0.002112074, 
    0.002048803, 0.002137614, 0.002312502, 0.00241608, 0.002528176, 
    0.002774062, 0.003058744, 0.003114375, 0.003187139, 0.003201746,
  0.002700802, 0.002638995, 0.002368008, 0.002174154, 0.002083241, 
    0.002124572, 0.002134447, 0.002200717, 0.002380768, 0.002473041, 
    0.002731812, 0.003024821, 0.0030786, 0.003164216, 0.003215525,
  0.002709616, 0.002415138, 0.002201826, 0.00219722, 0.002116809, 
    0.002146652, 0.002243345, 0.002099082, 0.002105422, 0.002430572, 
    0.00277636, 0.002969438, 0.003108478, 0.003199837, 0.003259045,
  0.002612262, 0.002292328, 0.002103707, 0.002079365, 0.002092649, 
    0.002220256, 0.00229593, 0.00238302, 0.002502695, 0.002632244, 
    0.002838423, 0.002977364, 0.003158116, 0.003259907, 0.00334271,
  0.002589083, 0.002215137, 0.002011084, 0.002030775, 0.002096066, 
    0.002240649, 0.002287489, 0.00233144, 0.0025481, 0.002698909, 
    0.002811162, 0.003069288, 0.003253155, 0.003316981, 0.003404229,
  0.002485674, 0.002079157, 0.00197617, 0.002045644, 0.002145236, 0.00224253, 
    0.002223239, 0.002254459, 0.002531571, 0.002668697, 0.002815099, 
    0.003128214, 0.003284708, 0.003343535, 0.003391952,
  0.002325961, 0.001974074, 0.001995035, 0.002051635, 0.002200408, 
    0.002218626, 0.002136875, 0.002190439, 0.002465502, 0.00260693, 
    0.002808558, 0.003140115, 0.003307843, 0.003363174, 0.003372821,
  0.002185455, 0.001971949, 0.002033713, 0.002057929, 0.002204464, 
    0.002160463, 0.002058756, 0.002104485, 0.002381139, 0.002524486, 
    0.002815001, 0.003107992, 0.003298836, 0.003413716, 0.003412788,
  0.002306184, 0.002450043, 0.00222531, 0.00214091, 0.002132559, 0.002177465, 
    0.002159858, 0.002322519, 0.002423563, 0.002567429, 0.002635158, 
    0.00273052, 0.002879266, 0.002935005, 0.003011807,
  0.00245036, 0.002282623, 0.002114893, 0.002057691, 0.002153145, 
    0.002173588, 0.002178412, 0.002390604, 0.002481546, 0.002586848, 
    0.002681387, 0.002827789, 0.003032672, 0.003024529, 0.003101076,
  0.002476807, 0.002200748, 0.002120845, 0.002082671, 0.002169388, 
    0.002039466, 0.002116248, 0.002344007, 0.002461678, 0.00257708, 
    0.002700248, 0.003005545, 0.003145144, 0.00325433, 0.003338289,
  0.002428544, 0.002250782, 0.00216592, 0.002143171, 0.002169506, 
    0.002136183, 0.002068453, 0.002189402, 0.002339698, 0.002541919, 
    0.002760936, 0.003168309, 0.00325609, 0.003263393, 0.003420681,
  0.002358465, 0.002073506, 0.002182458, 0.002127144, 0.002152526, 
    0.002141628, 0.002135094, 0.001968577, 0.002056734, 0.002520142, 
    0.00289506, 0.003304311, 0.003304879, 0.003275581, 0.003396024,
  0.002216307, 0.002071857, 0.002133016, 0.002139475, 0.002166017, 
    0.002121464, 0.00218267, 0.002365491, 0.002579915, 0.002715833, 
    0.003124714, 0.003462652, 0.00331511, 0.003181322, 0.003256258,
  0.002181379, 0.002122381, 0.002146587, 0.002179489, 0.00218548, 
    0.002088232, 0.002158837, 0.002443011, 0.002672874, 0.002896452, 
    0.003297279, 0.003525177, 0.003354644, 0.003175974, 0.00316891,
  0.002181367, 0.002176163, 0.002200021, 0.002178806, 0.002172481, 
    0.00210845, 0.002239757, 0.002522555, 0.00275897, 0.003019642, 
    0.003382039, 0.003537731, 0.003439214, 0.00332735, 0.003128359,
  0.002172557, 0.00226441, 0.002317, 0.002210936, 0.002154676, 0.002135995, 
    0.002329239, 0.002639425, 0.002855468, 0.003137419, 0.003423454, 
    0.003522333, 0.003470945, 0.003385975, 0.003224138,
  0.002286327, 0.002423199, 0.002432583, 0.002224104, 0.002207943, 
    0.002184815, 0.002442233, 0.002719256, 0.002975466, 0.003288507, 
    0.003441965, 0.003498978, 0.003464213, 0.003437372, 0.003287548,
  0.002256578, 0.002276199, 0.002310039, 0.002221901, 0.002207727, 
    0.00224553, 0.002285959, 0.002399335, 0.002513106, 0.002654342, 
    0.002760304, 0.002993797, 0.003061201, 0.003045981, 0.003267521,
  0.002317671, 0.00226842, 0.002284801, 0.002285579, 0.002309972, 
    0.002249344, 0.002317439, 0.002340667, 0.002467022, 0.002611269, 
    0.002756803, 0.002893408, 0.002957143, 0.002949665, 0.003137326,
  0.002333709, 0.002273941, 0.002397284, 0.002374233, 0.002367689, 
    0.002255487, 0.002333226, 0.002439442, 0.002552477, 0.002590253, 
    0.002675464, 0.002777805, 0.002852679, 0.002913189, 0.003102561,
  0.002258245, 0.002368552, 0.002464043, 0.002464668, 0.00247525, 
    0.002504532, 0.002407587, 0.002543673, 0.002546377, 0.002549987, 
    0.002652354, 0.00276347, 0.002916429, 0.002979347, 0.003081287,
  0.002322477, 0.002360505, 0.002561784, 0.002631168, 0.002593806, 
    0.00268841, 0.002786976, 0.002368473, 0.002323807, 0.002602609, 
    0.002700266, 0.002800357, 0.003018673, 0.003075256, 0.003139021,
  0.002348225, 0.002584861, 0.002680226, 0.002765071, 0.002663542, 
    0.002818871, 0.00296681, 0.003017218, 0.002982841, 0.002939556, 
    0.002914529, 0.00289246, 0.003030347, 0.003125956, 0.003118671,
  0.002526627, 0.002775792, 0.002812827, 0.002757396, 0.002768843, 
    0.002983663, 0.003070636, 0.003102719, 0.003083334, 0.003075292, 
    0.003042683, 0.003024307, 0.003102005, 0.003041231, 0.003041961,
  0.002798613, 0.002942185, 0.002805126, 0.002736501, 0.00286277, 
    0.003079234, 0.003129396, 0.003149221, 0.003136446, 0.003116847, 
    0.003093333, 0.003160833, 0.003173101, 0.003108122, 0.003157013,
  0.002938342, 0.002895312, 0.002843451, 0.002787946, 0.002937333, 
    0.003151576, 0.003173678, 0.00320752, 0.003215858, 0.003213862, 
    0.003280644, 0.003322072, 0.003147613, 0.003216104, 0.003299203,
  0.002968598, 0.002959898, 0.002849669, 0.002922276, 0.003003101, 
    0.003195047, 0.003210735, 0.003244349, 0.003277004, 0.003322544, 
    0.003361032, 0.003383445, 0.003291557, 0.00332915, 0.003309417,
  0.002471925, 0.002394755, 0.002398608, 0.0025822, 0.00278426, 0.002829636, 
    0.002897623, 0.002999858, 0.00303608, 0.003065129, 0.003025466, 
    0.00288775, 0.002886131, 0.002640844, 0.002858354,
  0.00237379, 0.002253649, 0.0025139, 0.002917731, 0.002925445, 0.002937276, 
    0.003002374, 0.003083153, 0.0031592, 0.003174939, 0.003171207, 
    0.003009113, 0.002899311, 0.002747128, 0.002865823,
  0.002448348, 0.002497849, 0.002756667, 0.002976901, 0.003000017, 
    0.002858121, 0.003048546, 0.003122517, 0.003237084, 0.003246392, 
    0.003212977, 0.003118714, 0.002943912, 0.002895291, 0.002880416,
  0.002487587, 0.002782538, 0.00285017, 0.003003567, 0.003066036, 
    0.003212094, 0.002944679, 0.003020072, 0.003151698, 0.003237488, 
    0.003239935, 0.003154795, 0.002943554, 0.002911857, 0.002943591,
  0.002708793, 0.002938158, 0.002823213, 0.003013257, 0.003118876, 
    0.003281735, 0.003255186, 0.002796243, 0.002761941, 0.003212223, 
    0.003350019, 0.003236092, 0.003007597, 0.002926809, 0.002962194,
  0.00306221, 0.00301807, 0.002829915, 0.003027122, 0.003165883, 0.003315033, 
    0.003330175, 0.003349105, 0.003340118, 0.003402288, 0.003452537, 
    0.003318397, 0.003073576, 0.002933806, 0.002972787,
  0.003158541, 0.002977568, 0.002817749, 0.003093679, 0.003251469, 
    0.003367853, 0.003367646, 0.003380367, 0.003385243, 0.003406608, 
    0.003504227, 0.003362258, 0.003098388, 0.002894572, 0.002911668,
  0.003078138, 0.002878987, 0.002745174, 0.00315866, 0.003322063, 
    0.003401094, 0.003424625, 0.003413325, 0.003373453, 0.003391496, 
    0.00353637, 0.003472543, 0.003179577, 0.002882414, 0.002856987,
  0.002983755, 0.002839809, 0.002814402, 0.00319732, 0.003353338, 
    0.003431705, 0.003464672, 0.003434168, 0.003371078, 0.003366271, 
    0.003448798, 0.003561868, 0.003161101, 0.00286325, 0.002826223,
  0.003100547, 0.002984029, 0.002912493, 0.003195547, 0.003337994, 
    0.003416346, 0.003474729, 0.00345392, 0.003419936, 0.003363149, 
    0.003429078, 0.003538172, 0.003253599, 0.002877578, 0.00281063,
  0.002562635, 0.00266767, 0.002656814, 0.002740099, 0.002912275, 
    0.002956842, 0.002991586, 0.003033574, 0.003093434, 0.00317306, 
    0.003195219, 0.003076688, 0.00289202, 0.002646262, 0.002749063,
  0.00272404, 0.002674916, 0.0026936, 0.00294565, 0.003076816, 0.003085479, 
    0.003095877, 0.003064551, 0.003059247, 0.003210894, 0.003233102, 
    0.003044782, 0.002871585, 0.002715693, 0.002730932,
  0.002894665, 0.002788013, 0.002716824, 0.00306354, 0.003273907, 
    0.003022113, 0.003168069, 0.003157785, 0.003073054, 0.003160451, 
    0.003224621, 0.003262652, 0.002937808, 0.002887073, 0.003008947,
  0.00301369, 0.002818561, 0.002859307, 0.003187122, 0.003355525, 
    0.003434861, 0.003119157, 0.003192475, 0.003045876, 0.003175055, 
    0.003323434, 0.003333531, 0.00297599, 0.002913565, 0.002903228,
  0.003066532, 0.002869869, 0.002966693, 0.003245753, 0.003416622, 
    0.003539702, 0.003545298, 0.002968313, 0.002646232, 0.003226569, 
    0.003395263, 0.003330254, 0.003005598, 0.002925144, 0.002880287,
  0.003078318, 0.002987675, 0.00303598, 0.003319098, 0.003463228, 
    0.003568849, 0.003613455, 0.003349121, 0.00312424, 0.00336322, 
    0.003429473, 0.003290659, 0.003048141, 0.003025674, 0.00299172,
  0.003061262, 0.003044043, 0.003150855, 0.003353181, 0.003447382, 
    0.003546298, 0.003512667, 0.003357921, 0.003334677, 0.00343368, 
    0.003416036, 0.003284299, 0.003126091, 0.003109096, 0.003044132,
  0.003068221, 0.00303397, 0.003238934, 0.003355484, 0.0034005, 0.003437988, 
    0.00337626, 0.003315104, 0.003428521, 0.003452137, 0.003426154, 
    0.003259432, 0.003152597, 0.00314718, 0.003105293,
  0.003038942, 0.003052511, 0.003257606, 0.003335504, 0.003391002, 
    0.003398198, 0.003385744, 0.003353491, 0.003383136, 0.003459902, 
    0.003408845, 0.003232385, 0.003181284, 0.003159871, 0.003134084,
  0.003080571, 0.003143964, 0.003294265, 0.003362272, 0.003418553, 
    0.003434316, 0.00344401, 0.003383345, 0.003409063, 0.003432621, 
    0.003382582, 0.003219596, 0.003174707, 0.003137086, 0.003112121,
  0.002573937, 0.002620959, 0.002766988, 0.002873074, 0.003034233, 
    0.003124151, 0.003311723, 0.003273132, 0.003006808, 0.00295158, 
    0.002815667, 0.002700639, 0.002820674, 0.002679696, 0.00304904,
  0.002708938, 0.002938489, 0.002855056, 0.00288427, 0.003071458, 
    0.003339879, 0.003440145, 0.003444245, 0.003185993, 0.003041744, 
    0.002916954, 0.002707161, 0.00246824, 0.002616462, 0.003162451,
  0.002928107, 0.002841309, 0.002694135, 0.002813021, 0.003179424, 
    0.00321055, 0.003439014, 0.003474508, 0.003207321, 0.003118633, 
    0.002950542, 0.002805679, 0.002369002, 0.002677703, 0.003344872,
  0.002883743, 0.002746144, 0.00269283, 0.002987617, 0.003430422, 
    0.003510182, 0.003155324, 0.003372889, 0.003146295, 0.003096231, 
    0.002980058, 0.002850358, 0.002682089, 0.003019463, 0.003380679,
  0.002869524, 0.002722902, 0.002773697, 0.003248412, 0.003542124, 
    0.00344644, 0.003360078, 0.002711192, 0.002530564, 0.003050954, 
    0.003003963, 0.00296358, 0.0030052, 0.003178566, 0.003396162,
  0.002908185, 0.002782287, 0.002954452, 0.003358629, 0.003371029, 
    0.003436256, 0.003320026, 0.002952382, 0.002917374, 0.003009137, 
    0.003082597, 0.003115235, 0.003244602, 0.003300887, 0.003459573,
  0.002911642, 0.002817493, 0.003071112, 0.003329798, 0.003167813, 
    0.003061612, 0.002969672, 0.00292931, 0.003058899, 0.003159964, 
    0.003231383, 0.00329451, 0.003342067, 0.003382889, 0.00345165,
  0.002909183, 0.002842889, 0.003266771, 0.003304482, 0.003315463, 
    0.003262473, 0.003236176, 0.003217062, 0.003223481, 0.003269083, 
    0.003269595, 0.003301692, 0.003328663, 0.003333068, 0.003388734,
  0.002958573, 0.00308905, 0.003346157, 0.003324444, 0.003318371, 0.00331779, 
    0.003287435, 0.003289168, 0.003286386, 0.003256264, 0.003268282, 
    0.00328681, 0.003302473, 0.003330722, 0.003354979,
  0.002975588, 0.003270624, 0.003401895, 0.003415711, 0.00340182, 
    0.003364217, 0.003340338, 0.003276268, 0.00322324, 0.003205603, 
    0.003246147, 0.003266623, 0.003269901, 0.003284988, 0.003311233,
  0.003506077, 0.003263942, 0.003216129, 0.002974885, 0.002796155, 
    0.002744895, 0.002838403, 0.003131792, 0.003159787, 0.002694519, 
    0.003141455, 0.002746979, 0.002513786, 0.002657252, 0.003059604,
  0.003316854, 0.003197215, 0.003008078, 0.002728265, 0.002658505, 
    0.002908026, 0.003046867, 0.00314237, 0.00316704, 0.003085011, 
    0.00305424, 0.002560437, 0.002344328, 0.002700398, 0.003050724,
  0.003347398, 0.003085616, 0.002725889, 0.002575105, 0.002688332, 
    0.002776424, 0.003333796, 0.003385308, 0.003318135, 0.002999924, 
    0.002926561, 0.002706191, 0.002325919, 0.002595474, 0.003248278,
  0.003285831, 0.002906822, 0.002562158, 0.002495905, 0.002798946, 
    0.003135808, 0.002836044, 0.003399677, 0.003312672, 0.003068683, 
    0.002972432, 0.002751399, 0.002477792, 0.002789515, 0.003473098,
  0.003050679, 0.002674889, 0.00250277, 0.002642256, 0.002989069, 0.00333089, 
    0.003370112, 0.00278021, 0.002542247, 0.002833385, 0.002873232, 
    0.002559915, 0.002682985, 0.003268594, 0.003669228,
  0.002885628, 0.002641088, 0.002565376, 0.002875376, 0.003062733, 
    0.003226082, 0.003261471, 0.002882983, 0.002744124, 0.002710552, 
    0.00260341, 0.002707534, 0.003203498, 0.003632962, 0.003704047,
  0.002814965, 0.002654382, 0.002650853, 0.002864578, 0.0030422, 0.003090674, 
    0.003018314, 0.002861387, 0.002723453, 0.00271292, 0.002946013, 
    0.003161405, 0.003527372, 0.003685059, 0.00369938,
  0.002813979, 0.002771555, 0.003040542, 0.002840183, 0.002975409, 
    0.00301172, 0.003027136, 0.003040458, 0.003087596, 0.003220626, 
    0.003257994, 0.003492128, 0.00364154, 0.003660254, 0.003638204,
  0.002910682, 0.003069099, 0.003158536, 0.003090671, 0.003077411, 
    0.003141308, 0.003227646, 0.003295814, 0.003339075, 0.003366187, 
    0.00352392, 0.003623334, 0.003634743, 0.003617229, 0.00358338,
  0.00301599, 0.003124356, 0.003204226, 0.003117073, 0.00314893, 0.00318242, 
    0.003153742, 0.003225541, 0.003384922, 0.003515659, 0.003607733, 
    0.003619674, 0.003598568, 0.003564528, 0.003518612,
  0.005352847, 0.004075862, 0.004393763, 0.003480387, 0.003288331, 
    0.003106636, 0.002867039, 0.002814926, 0.00282716, 0.002945787, 
    0.002825507, 0.002619939, 0.002510667, 0.002720712, 0.002973268,
  0.003962945, 0.003780751, 0.003606422, 0.003291894, 0.003206281, 
    0.002982687, 0.002851569, 0.002808731, 0.002899359, 0.002875023, 
    0.002699086, 0.0022876, 0.002471191, 0.002671859, 0.002997274,
  0.0039211, 0.003697131, 0.003449706, 0.003193506, 0.003068339, 0.002806898, 
    0.002776313, 0.002754319, 0.002853138, 0.002664399, 0.002560091, 
    0.002474276, 0.002702703, 0.002801397, 0.003307965,
  0.003879969, 0.003600946, 0.003338838, 0.00313195, 0.002951382, 
    0.002817354, 0.002627777, 0.002828929, 0.002946039, 0.002710918, 
    0.002669649, 0.002742057, 0.002740853, 0.003001237, 0.003530554,
  0.00364225, 0.003341876, 0.003137452, 0.002931045, 0.002820287, 
    0.002823041, 0.002844522, 0.002594255, 0.002435644, 0.002605187, 
    0.002621052, 0.002644266, 0.0027878, 0.003353381, 0.003659302,
  0.003155299, 0.002981215, 0.002823217, 0.002739453, 0.002745362, 
    0.002888557, 0.002964922, 0.002791998, 0.002626257, 0.002588474, 
    0.002654796, 0.002708867, 0.003126743, 0.003599838, 0.003685518,
  0.002736859, 0.002629075, 0.002520424, 0.002775156, 0.002925149, 
    0.003016158, 0.003100445, 0.002876563, 0.00263626, 0.002692142, 
    0.002642434, 0.002912019, 0.003512057, 0.003661284, 0.003682178,
  0.002519367, 0.002428485, 0.002926224, 0.002714227, 0.002943009, 
    0.00309017, 0.003181738, 0.00291268, 0.00271803, 0.002642236, 
    0.002808661, 0.003391061, 0.003631738, 0.003653685, 0.003686272,
  0.002627661, 0.002717112, 0.002988507, 0.002990994, 0.003033933, 
    0.003073001, 0.003195641, 0.003064016, 0.002623232, 0.002728348, 
    0.003169744, 0.003616043, 0.003633587, 0.003634277, 0.003634014,
  0.002770915, 0.002878002, 0.003050266, 0.002930796, 0.003049689, 
    0.003120498, 0.003080896, 0.002901271, 0.002873187, 0.003186044, 
    0.003627679, 0.003640628, 0.003610621, 0.003596763, 0.003568919,
  0.006419483, 0.004975914, 0.00557236, 0.004152661, 0.003862522, 
    0.003630489, 0.003425476, 0.003266354, 0.003134561, 0.003107334, 
    0.003025692, 0.002871685, 0.002757013, 0.00261023, 0.00273182,
  0.004763334, 0.004494915, 0.004173465, 0.003743554, 0.003688925, 
    0.003527537, 0.00334156, 0.003123543, 0.002973644, 0.002925095, 
    0.002805662, 0.002614876, 0.002493304, 0.002543924, 0.002727112,
  0.004530817, 0.004267276, 0.003838796, 0.003574731, 0.003468917, 
    0.003293794, 0.0031068, 0.002928806, 0.002758063, 0.002601657, 
    0.002507356, 0.002511796, 0.002597889, 0.002697997, 0.003146299,
  0.004519406, 0.004163117, 0.003752665, 0.00353491, 0.003323048, 0.00305448, 
    0.002786336, 0.002806717, 0.002625797, 0.002440088, 0.002382611, 
    0.002565253, 0.002739976, 0.003135547, 0.003533738,
  0.004444832, 0.003989377, 0.003708069, 0.00343275, 0.003236209, 
    0.002918397, 0.002710371, 0.002376672, 0.002211547, 0.002332663, 
    0.002444687, 0.002839654, 0.00330354, 0.003596833, 0.003699113,
  0.00431719, 0.003878986, 0.003527679, 0.003273792, 0.00311576, 0.002839869, 
    0.002698651, 0.002572581, 0.002601813, 0.002634944, 0.002731732, 
    0.00323301, 0.003591022, 0.003683442, 0.003698276,
  0.004091286, 0.003775207, 0.003380009, 0.003166693, 0.003006664, 
    0.002841146, 0.002752896, 0.002615723, 0.002589101, 0.002671598, 
    0.002997923, 0.003518516, 0.003652902, 0.003679711, 0.003712332,
  0.003760995, 0.003527789, 0.003173695, 0.003033383, 0.002884412, 
    0.002792062, 0.002778868, 0.002623249, 0.00249427, 0.002560846, 
    0.003251465, 0.0035879, 0.003635475, 0.003685565, 0.003715061,
  0.003452953, 0.003233477, 0.003005784, 0.002946465, 0.002828314, 
    0.002777227, 0.002795215, 0.002517379, 0.002339333, 0.002843722, 
    0.003440412, 0.003619384, 0.003631884, 0.003653977, 0.003672163,
  0.003231653, 0.003094976, 0.002966075, 0.002899292, 0.002823171, 
    0.002784317, 0.002829885, 0.002833377, 0.002778661, 0.00315398, 
    0.003566989, 0.003638133, 0.003612374, 0.003593338, 0.00356362,
  0.005527923, 0.004640535, 0.005188029, 0.004399619, 0.004319856, 
    0.004320093, 0.004106665, 0.003828174, 0.003626247, 0.003615435, 
    0.003528295, 0.003165987, 0.002933834, 0.00277885, 0.002630771,
  0.004241121, 0.004172189, 0.004173533, 0.004071536, 0.004233961, 
    0.003904311, 0.003854664, 0.003697007, 0.00358587, 0.003480091, 
    0.003269344, 0.002950547, 0.002661899, 0.002714539, 0.002879363,
  0.004378444, 0.004238581, 0.004065173, 0.004065818, 0.003809539, 
    0.003845559, 0.003687249, 0.00359451, 0.003430421, 0.003184247, 
    0.002964657, 0.00269079, 0.002502498, 0.002518424, 0.002961508,
  0.004461398, 0.004205644, 0.003983141, 0.003875128, 0.003669377, 
    0.003567413, 0.003306711, 0.003233282, 0.003111482, 0.00294083, 
    0.002671855, 0.002504635, 0.002764026, 0.002988273, 0.003224314,
  0.00451884, 0.004111383, 0.003951444, 0.003764544, 0.003649911, 
    0.003403071, 0.003194683, 0.002914199, 0.002517659, 0.002671448, 
    0.002608275, 0.002815411, 0.003106195, 0.003391636, 0.003543759,
  0.004533597, 0.004092967, 0.003774056, 0.003635007, 0.003494804, 
    0.003227867, 0.003047894, 0.002928255, 0.002732686, 0.002703584, 
    0.00271521, 0.00315049, 0.003473347, 0.003637982, 0.003678482,
  0.00447678, 0.004072579, 0.003636207, 0.003379453, 0.003070842, 
    0.002806175, 0.002754973, 0.002714337, 0.002701702, 0.002941674, 
    0.00334742, 0.003595961, 0.003661358, 0.003650697, 0.003616828,
  0.004434214, 0.003952415, 0.003397162, 0.00305709, 0.002833228, 
    0.002778169, 0.002855222, 0.002967367, 0.003122425, 0.003497354, 
    0.003641023, 0.003650772, 0.003638328, 0.003637788, 0.003624247,
  0.004150697, 0.003593055, 0.003073267, 0.002859626, 0.002828127, 0.0028384, 
    0.002917382, 0.003073447, 0.003344213, 0.003608086, 0.003654805, 
    0.003649087, 0.003644496, 0.003640056, 0.003637178,
  0.00381239, 0.00330701, 0.002997048, 0.002861677, 0.002869977, 0.002899863, 
    0.002983541, 0.003188381, 0.003400497, 0.0036125, 0.00364365, 0.00363095, 
    0.003606032, 0.003588875, 0.003554419,
  0.004095216, 0.00370648, 0.004172163, 0.003919837, 0.00399834, 0.003978968, 
    0.003916197, 0.003938984, 0.004082974, 0.003974371, 0.003811656, 
    0.003595053, 0.003444513, 0.003634907, 0.003718552,
  0.004113457, 0.003790418, 0.00379076, 0.003745425, 0.003914812, 
    0.003802566, 0.00381149, 0.003931057, 0.003974709, 0.00391496, 
    0.003725973, 0.00353297, 0.003415331, 0.003437587, 0.003453018,
  0.004362618, 0.004089459, 0.003870755, 0.003725586, 0.003780709, 
    0.003865069, 0.00374342, 0.003848863, 0.003922985, 0.003902039, 
    0.003706367, 0.003531266, 0.003361706, 0.003302443, 0.003255328,
  0.004440519, 0.004211539, 0.003953911, 0.003826609, 0.003730212, 
    0.003731019, 0.003965269, 0.003843471, 0.003875703, 0.003790623, 
    0.003686828, 0.003486321, 0.003408711, 0.003265161, 0.003107914,
  0.004458425, 0.004143961, 0.003999481, 0.003847419, 0.003807564, 
    0.003597839, 0.003644582, 0.003910865, 0.003706448, 0.003704183, 
    0.003625032, 0.003502016, 0.003294843, 0.003140175, 0.003101652,
  0.004383679, 0.004135876, 0.003897518, 0.003823935, 0.003810931, 
    0.003834722, 0.003783426, 0.003654449, 0.003527049, 0.003497506, 
    0.003445115, 0.003338378, 0.003208036, 0.003158984, 0.003235784,
  0.004245054, 0.004045694, 0.003750835, 0.003691411, 0.003663405, 
    0.003603609, 0.003538864, 0.003419689, 0.003319774, 0.003287817, 
    0.00326634, 0.003246904, 0.003276592, 0.003365579, 0.003422188,
  0.004020405, 0.003813236, 0.003484487, 0.003410263, 0.00339789, 
    0.003357713, 0.003281318, 0.003258784, 0.003236843, 0.003295586, 
    0.003366045, 0.003409427, 0.003485244, 0.003539931, 0.003546404,
  0.003703748, 0.003476171, 0.003277384, 0.003303793, 0.00333729, 
    0.003360178, 0.003384158, 0.003439849, 0.003544512, 0.00357496, 
    0.003566786, 0.003591212, 0.003612407, 0.003600611, 0.003584682,
  0.003561139, 0.003400465, 0.003296678, 0.003349188, 0.003482438, 
    0.003578622, 0.003639172, 0.00362954, 0.003668967, 0.003671747, 
    0.003669213, 0.003615381, 0.003479292, 0.00327793, 0.00340197,
  0.004577772, 0.004018121, 0.004355425, 0.003972348, 0.003875495, 
    0.003971213, 0.00392131, 0.003851247, 0.003781231, 0.003796627, 
    0.003984944, 0.003879256, 0.003812062, 0.00398943, 0.003971563,
  0.003993856, 0.003823977, 0.003802353, 0.00376048, 0.003841701, 
    0.003881025, 0.003885631, 0.003816816, 0.003736178, 0.003722272, 
    0.00381624, 0.003801961, 0.003750767, 0.003947758, 0.003889849,
  0.004212066, 0.004061363, 0.003914405, 0.003700516, 0.003768937, 
    0.003864372, 0.003849174, 0.003792631, 0.003780164, 0.003703214, 
    0.003734603, 0.003743112, 0.003685725, 0.003839007, 0.003768678,
  0.004326959, 0.004141533, 0.003963287, 0.003809733, 0.003706312, 
    0.003812286, 0.003937217, 0.003868839, 0.003819016, 0.003781791, 
    0.003743362, 0.003694304, 0.003619296, 0.003785633, 0.003691998,
  0.004392824, 0.004064004, 0.003924957, 0.003751608, 0.003757241, 
    0.003770059, 0.003817619, 0.004028707, 0.003929878, 0.003827085, 
    0.003763839, 0.003662435, 0.003699958, 0.003702495, 0.003602243,
  0.004352686, 0.004066572, 0.003831753, 0.003717409, 0.003728528, 
    0.003788194, 0.003786933, 0.003752233, 0.003763689, 0.003766812, 
    0.003773813, 0.003708658, 0.003677643, 0.00363601, 0.003559669,
  0.004329206, 0.004095177, 0.003755212, 0.003684125, 0.003708854, 
    0.003716838, 0.003730165, 0.003739126, 0.003747339, 0.003740234, 
    0.003740231, 0.003692644, 0.003617893, 0.003521527, 0.003445684,
  0.004184198, 0.003929361, 0.003646911, 0.003607558, 0.003641099, 
    0.003671836, 0.003682391, 0.003697367, 0.003701276, 0.003697479, 
    0.003663113, 0.003588716, 0.003488896, 0.003402669, 0.003368798,
  0.003977186, 0.003781708, 0.003556854, 0.003551945, 0.003563548, 
    0.003573032, 0.003590703, 0.003594719, 0.003601589, 0.003599282, 
    0.003556496, 0.003510351, 0.003456013, 0.003453292, 0.003478991,
  0.003879569, 0.003758856, 0.003594476, 0.003580739, 0.003563931, 
    0.003552637, 0.003536957, 0.003540478, 0.003596399, 0.003607374, 
    0.003579453, 0.00350443, 0.003445049, 0.003457369, 0.003581242,
  0.004317152, 0.00398067, 0.004445626, 0.004023666, 0.004055714, 
    0.004405046, 0.004211536, 0.004006306, 0.004153015, 0.003730841, 
    0.003895445, 0.00405925, 0.004006664, 0.004093372, 0.004022195,
  0.004007159, 0.003866175, 0.003846607, 0.003756748, 0.003872087, 
    0.003996195, 0.004032813, 0.003890364, 0.003864457, 0.003546306, 
    0.00371449, 0.003914732, 0.003976148, 0.004066919, 0.003947868,
  0.004164326, 0.004097636, 0.003984497, 0.003692859, 0.003775004, 
    0.003932491, 0.003930435, 0.003840405, 0.003816568, 0.003489369, 
    0.003653127, 0.003830735, 0.00389926, 0.003943107, 0.003846948,
  0.004074844, 0.003984732, 0.003927835, 0.003814843, 0.003716295, 
    0.003805553, 0.003930227, 0.003760698, 0.003703421, 0.003505626, 
    0.003701715, 0.003799413, 0.003795248, 0.00388409, 0.003794706,
  0.003924906, 0.003867961, 0.003841036, 0.00375792, 0.003728265, 0.00375333, 
    0.003817082, 0.00392073, 0.003860109, 0.003609046, 0.003714954, 
    0.00378048, 0.003782782, 0.003846907, 0.0038668,
  0.003817841, 0.003830642, 0.00377073, 0.003657811, 0.003714004, 
    0.003754117, 0.003804781, 0.003731028, 0.003728393, 0.003673384, 
    0.003722268, 0.003765983, 0.00376635, 0.00381959, 0.00381292,
  0.00373009, 0.003791478, 0.003718395, 0.003654317, 0.003701611, 0.00376203, 
    0.003810661, 0.003758056, 0.003699627, 0.003629721, 0.003673865, 
    0.003675584, 0.003739316, 0.003811101, 0.003750171,
  0.003634324, 0.003702805, 0.003624951, 0.003669, 0.003718747, 0.003775891, 
    0.003772006, 0.003743508, 0.003701734, 0.003613905, 0.003630196, 
    0.00362447, 0.003703556, 0.003716701, 0.003650578,
  0.003484901, 0.003510553, 0.003503283, 0.003641015, 0.003735327, 
    0.00376666, 0.003738907, 0.003654582, 0.003605261, 0.003626899, 
    0.003715702, 0.003624249, 0.0036712, 0.003675255, 0.003641885,
  0.003312474, 0.003284479, 0.003364612, 0.003518698, 0.003661979, 
    0.003703272, 0.003657736, 0.003620238, 0.00362495, 0.003659979, 
    0.003608948, 0.003635683, 0.003615428, 0.003606881, 0.003617145,
  0.004017376, 0.003728673, 0.003898028, 0.003658428, 0.003743894, 
    0.003885835, 0.00379466, 0.003760903, 0.003857755, 0.003805212, 
    0.004086569, 0.004072133, 0.00395415, 0.004068504, 0.004020636,
  0.003882137, 0.003715515, 0.003673499, 0.003583245, 0.003694941, 
    0.003718453, 0.003726827, 0.003726784, 0.003749799, 0.003732353, 
    0.00394848, 0.003922866, 0.003946194, 0.004010011, 0.003986678,
  0.003844634, 0.003755188, 0.003727192, 0.003581643, 0.003656742, 
    0.00369926, 0.003746296, 0.003775641, 0.003784765, 0.003685263, 
    0.00367342, 0.003739315, 0.003903314, 0.003958145, 0.003979824,
  0.003951812, 0.003915233, 0.003860228, 0.003751668, 0.003666076, 
    0.003697522, 0.003715442, 0.003703279, 0.003786366, 0.003605111, 
    0.003695829, 0.003789471, 0.00387956, 0.003905153, 0.003841358,
  0.004034906, 0.003964266, 0.003917701, 0.003771702, 0.003736542, 
    0.003691747, 0.003682792, 0.003750677, 0.003990491, 0.003635402, 
    0.003645429, 0.003787551, 0.003856586, 0.003891964, 0.003931068,
  0.004067614, 0.004009947, 0.003890082, 0.003706903, 0.003728251, 
    0.003719199, 0.003715601, 0.003683015, 0.003717191, 0.003606913, 
    0.003747207, 0.003793027, 0.003843577, 0.003856929, 0.003842615,
  0.004057255, 0.00408119, 0.003835494, 0.003596677, 0.00365957, 0.003698497, 
    0.00372132, 0.003735279, 0.003646491, 0.003598605, 0.003714545, 
    0.003787953, 0.003807101, 0.003777683, 0.003711094,
  0.004089961, 0.004014657, 0.003664046, 0.003576278, 0.003645486, 
    0.003688793, 0.003701624, 0.003710938, 0.003671749, 0.003646782, 
    0.003725498, 0.003742008, 0.003746546, 0.003680649, 0.003628526,
  0.003974634, 0.003926645, 0.003656902, 0.003669611, 0.003681615, 
    0.003705068, 0.003696301, 0.003679474, 0.003672734, 0.003659782, 
    0.00373025, 0.003707092, 0.003705522, 0.003674492, 0.003666236,
  0.003857675, 0.003912207, 0.003765777, 0.00374277, 0.003724763, 
    0.003711639, 0.003654299, 0.003634853, 0.003654998, 0.003698232, 
    0.00367519, 0.0036874, 0.003684616, 0.003659198, 0.003662176,
  0.005225115, 0.004439325, 0.004885283, 0.004091873, 0.003995848, 
    0.004167886, 0.003864588, 0.003744609, 0.003663691, 0.003592907, 
    0.003712787, 0.003738593, 0.003720863, 0.003750117, 0.003697298,
  0.004310056, 0.00401032, 0.004044116, 0.003767733, 0.003899463, 
    0.003990655, 0.003824504, 0.003745253, 0.0036711, 0.003620469, 
    0.003721163, 0.003725723, 0.003720827, 0.003797182, 0.003865519,
  0.004322732, 0.004117075, 0.00389953, 0.003589005, 0.003649232, 
    0.003706954, 0.003647225, 0.003677393, 0.003671647, 0.003624532, 
    0.00363026, 0.003696595, 0.003708771, 0.003750275, 0.00381832,
  0.004085425, 0.004004641, 0.003911672, 0.00380678, 0.003666534, 
    0.003699852, 0.003694057, 0.003688128, 0.003624372, 0.003640221, 
    0.003661508, 0.003695382, 0.003717584, 0.003720125, 0.003755274,
  0.004101302, 0.00411399, 0.004045532, 0.003832079, 0.003788905, 0.00374761, 
    0.003733135, 0.003479643, 0.003431128, 0.003625123, 0.003629656, 
    0.003714254, 0.003748298, 0.003737635, 0.003803155,
  0.004358937, 0.004248704, 0.004049819, 0.003741979, 0.003740364, 
    0.003752433, 0.003744869, 0.003614471, 0.003588168, 0.003613062, 
    0.003689026, 0.00366293, 0.00365263, 0.003713379, 0.003793334,
  0.004433581, 0.004272909, 0.003836646, 0.003520786, 0.003572743, 
    0.003665821, 0.003717029, 0.003708779, 0.003623699, 0.003539205, 
    0.003585749, 0.003632672, 0.003683517, 0.003681564, 0.003711364,
  0.004330311, 0.003859418, 0.003624454, 0.003485213, 0.003594313, 
    0.003664124, 0.003685941, 0.00365505, 0.003617452, 0.003634899, 
    0.003638204, 0.003687085, 0.003687503, 0.00365676, 0.003632079,
  0.004015577, 0.003869516, 0.003613665, 0.003646438, 0.003664023, 
    0.00368339, 0.003663947, 0.003613045, 0.003656716, 0.003698698, 
    0.003729407, 0.003701608, 0.003669989, 0.003633809, 0.003591408,
  0.003965264, 0.003860351, 0.003724774, 0.003701794, 0.003688221, 
    0.003667859, 0.003618967, 0.003557749, 0.00369661, 0.003752948, 
    0.003749351, 0.003691938, 0.003641135, 0.003590642, 0.003521488,
  0.006779321, 0.005142569, 0.005927658, 0.004443092, 0.004358677, 
    0.004907922, 0.004252255, 0.003984889, 0.004144134, 0.004758029, 
    0.004586207, 0.004264683, 0.00366784, 0.003741747, 0.003687793,
  0.00505955, 0.004660718, 0.004621404, 0.004121403, 0.004622187, 
    0.004865791, 0.003914837, 0.00379615, 0.003889195, 0.004219634, 
    0.003987107, 0.003703974, 0.003608104, 0.003530452, 0.003588706,
  0.004621478, 0.004485135, 0.004185619, 0.003892804, 0.004090715, 
    0.004096819, 0.003763991, 0.003667128, 0.003634596, 0.003615023, 
    0.003432221, 0.003448001, 0.003482326, 0.003531145, 0.003644202,
  0.004277708, 0.004200398, 0.00403059, 0.003929795, 0.003764968, 
    0.003821156, 0.00377376, 0.003565766, 0.003459903, 0.003385419, 
    0.003366387, 0.003413593, 0.003470119, 0.003516747, 0.003652421,
  0.00419755, 0.0041037, 0.003995244, 0.003766144, 0.003718772, 0.003680384, 
    0.003687945, 0.003724983, 0.003592358, 0.00335384, 0.003368203, 
    0.003373991, 0.003505519, 0.003531158, 0.00357225,
  0.004327164, 0.004225425, 0.003934636, 0.003649937, 0.003673212, 0.0037056, 
    0.003681754, 0.00366186, 0.003587724, 0.003476776, 0.003425515, 
    0.003408471, 0.003239624, 0.003506703, 0.003562019,
  0.004375311, 0.004314355, 0.003904435, 0.003601145, 0.003553986, 
    0.003641594, 0.00368813, 0.003705048, 0.003660801, 0.003498167, 
    0.003583145, 0.003512563, 0.003266441, 0.003499931, 0.003436625,
  0.004440296, 0.004228078, 0.003819734, 0.003633258, 0.003614704, 
    0.003631022, 0.003643676, 0.003648952, 0.003681099, 0.003626132, 
    0.00360752, 0.003479991, 0.003314551, 0.003461615, 0.003318906,
  0.004323624, 0.004101267, 0.003757518, 0.003722172, 0.003693939, 
    0.003675542, 0.003653776, 0.003657503, 0.003693342, 0.00369124, 
    0.003592697, 0.003429657, 0.003472095, 0.003499897, 0.003254799,
  0.004189234, 0.004038902, 0.003826181, 0.003761722, 0.003717867, 
    0.003683522, 0.003627555, 0.003623528, 0.003688587, 0.003675482, 
    0.003549737, 0.003443113, 0.003575601, 0.003464645, 0.003165409,
  0.004797311, 0.004591998, 0.005549639, 0.004272943, 0.004522379, 
    0.004897947, 0.004234114, 0.00421886, 0.004682174, 0.005663034, 
    0.00502969, 0.004205684, 0.003757468, 0.003630539, 0.003804195,
  0.004274101, 0.004387013, 0.004512896, 0.004321691, 0.004947383, 
    0.004744755, 0.004038999, 0.004082529, 0.004211407, 0.004466791, 
    0.004183263, 0.003528035, 0.003292959, 0.003379778, 0.003685762,
  0.00439127, 0.004511352, 0.004324462, 0.0041536, 0.00424961, 0.004020671, 
    0.003947197, 0.003841301, 0.003833243, 0.003637712, 0.00346665, 
    0.003280777, 0.003219166, 0.003508525, 0.003677287,
  0.00433214, 0.004390488, 0.004296163, 0.004176734, 0.003933277, 
    0.004006227, 0.003897837, 0.003766798, 0.00361874, 0.003417987, 
    0.003318158, 0.00324237, 0.00321471, 0.003437595, 0.003579085,
  0.00424604, 0.004182588, 0.004158094, 0.003961439, 0.003895193, 0.00387839, 
    0.003866448, 0.003939265, 0.003659312, 0.003402361, 0.003303362, 
    0.003226198, 0.003167051, 0.003360372, 0.003484132,
  0.004144898, 0.004079465, 0.003885134, 0.00373461, 0.003772134, 
    0.003841082, 0.003810189, 0.003724258, 0.003626433, 0.00344796, 
    0.00327332, 0.003166443, 0.003127942, 0.003252079, 0.003397017,
  0.004040016, 0.00402952, 0.0037159, 0.003582298, 0.003606562, 0.003790606, 
    0.003823849, 0.003715027, 0.003524993, 0.003377635, 0.003309368, 
    0.003115452, 0.002980613, 0.002928345, 0.002992298,
  0.004179524, 0.003850871, 0.003700726, 0.003595924, 0.003647693, 
    0.003746418, 0.003749481, 0.003619488, 0.003490871, 0.00346413, 
    0.003369247, 0.003185489, 0.002938938, 0.002860625, 0.002783315,
  0.004263597, 0.003807824, 0.00363674, 0.003722352, 0.003729795, 
    0.003743174, 0.00371995, 0.003631265, 0.003584778, 0.003553041, 
    0.003409743, 0.003056723, 0.002904914, 0.00279737, 0.0027214,
  0.004198238, 0.003920384, 0.003714445, 0.003736897, 0.003749542, 
    0.003736197, 0.003691946, 0.003633653, 0.003637934, 0.003601142, 
    0.003389983, 0.003019732, 0.002935508, 0.002752542, 0.002603386,
  0.003663004, 0.003788437, 0.004396066, 0.003841618, 0.004213545, 
    0.004442162, 0.003995018, 0.00414126, 0.004320701, 0.005022061, 
    0.005107011, 0.004613657, 0.004163635, 0.004022573, 0.004134074,
  0.003772837, 0.003917601, 0.004055291, 0.003939236, 0.004510188, 
    0.004385501, 0.00389936, 0.003937828, 0.004003893, 0.004165758, 
    0.004452001, 0.003818069, 0.003700931, 0.0036541, 0.003786535,
  0.003972259, 0.004062309, 0.004106872, 0.003896768, 0.004024317, 
    0.003876689, 0.003813941, 0.003747132, 0.003715794, 0.003643613, 
    0.003579869, 0.003530995, 0.003566619, 0.003711377, 0.003755905,
  0.004148727, 0.004076741, 0.004093442, 0.003967358, 0.003664797, 
    0.003732446, 0.003626279, 0.00353498, 0.003389232, 0.003401155, 
    0.003436575, 0.00346521, 0.003472072, 0.003543558, 0.003470018,
  0.004226859, 0.004014644, 0.004025347, 0.003859944, 0.003700488, 
    0.003624757, 0.003565877, 0.003382508, 0.002923619, 0.003276244, 
    0.003292202, 0.003249548, 0.003159194, 0.003180006, 0.003092516,
  0.004282606, 0.00402614, 0.003882759, 0.003757674, 0.003685588, 
    0.003644893, 0.003518837, 0.003402057, 0.003276994, 0.003153969, 
    0.003142625, 0.00303277, 0.002909831, 0.002786257, 0.002795663,
  0.004297456, 0.004108677, 0.0037422, 0.003624691, 0.003585065, 0.003616424, 
    0.003528292, 0.003398557, 0.003210346, 0.003103254, 0.003046454, 
    0.002855653, 0.002659914, 0.002625499, 0.002561667,
  0.004178014, 0.004124686, 0.00356871, 0.003540706, 0.003579398, 
    0.003630735, 0.003459726, 0.003315536, 0.003112443, 0.003007608, 
    0.002884988, 0.002616307, 0.002492561, 0.002406268, 0.002379506,
  0.004420948, 0.004057494, 0.003586331, 0.00365448, 0.003661117, 0.00365293, 
    0.003435899, 0.003270665, 0.003087058, 0.00297547, 0.002713851, 
    0.002544272, 0.002448017, 0.002404144, 0.002433505,
  0.00445765, 0.004051869, 0.003719359, 0.003750788, 0.003743307, 
    0.003679271, 0.003394109, 0.003261576, 0.003039806, 0.002848955, 
    0.002628804, 0.002528028, 0.002432629, 0.002371121, 0.002453376,
  0.005853028, 0.004310134, 0.00463291, 0.003892678, 0.004087208, 
    0.004399817, 0.003968023, 0.004130744, 0.004366331, 0.005293381, 
    0.00517423, 0.004765355, 0.004605495, 0.00450968, 0.00442926,
  0.004419203, 0.004142478, 0.004186285, 0.003948925, 0.00456107, 
    0.004320932, 0.003877302, 0.003926256, 0.003921362, 0.004259254, 
    0.004450481, 0.00404704, 0.003904115, 0.003738046, 0.003909385,
  0.004521651, 0.004274802, 0.004154145, 0.003926228, 0.004331545, 
    0.003837966, 0.003807031, 0.00372776, 0.003733019, 0.003691751, 
    0.003803033, 0.003575078, 0.003503979, 0.003482125, 0.003393803,
  0.004599418, 0.004364075, 0.004157765, 0.004023421, 0.003792324, 
    0.003776699, 0.003710056, 0.003631323, 0.003626846, 0.003642953, 
    0.003609651, 0.00345356, 0.003275035, 0.003167728, 0.003103575,
  0.004532485, 0.004253005, 0.004131925, 0.003891869, 0.003675224, 
    0.003629655, 0.003627535, 0.003331305, 0.003181813, 0.003576174, 
    0.003421772, 0.003062405, 0.002861684, 0.002841055, 0.002934158,
  0.004454643, 0.004202331, 0.003996707, 0.003701456, 0.003612146, 
    0.003626566, 0.003537756, 0.003416239, 0.003400752, 0.003355443, 
    0.003077338, 0.002749939, 0.00265007, 0.002619589, 0.002756467,
  0.004380819, 0.004188192, 0.003796852, 0.003582665, 0.003543033, 
    0.003548545, 0.003534937, 0.003361244, 0.003292121, 0.003029105, 
    0.002803107, 0.002612757, 0.002535854, 0.002472328, 0.002661997,
  0.004300545, 0.004078026, 0.003598072, 0.003514207, 0.003498524, 
    0.003515675, 0.00338238, 0.003317478, 0.003147189, 0.002858264, 
    0.002560144, 0.002431949, 0.002289902, 0.002486414, 0.002792762,
  0.004252626, 0.003876944, 0.003520142, 0.003562152, 0.003571418, 
    0.003536889, 0.003346133, 0.003234541, 0.002974481, 0.002694041, 
    0.002463048, 0.002332424, 0.002379881, 0.002808249, 0.003136676,
  0.004294202, 0.003904822, 0.003644444, 0.003679612, 0.003670902, 
    0.003548342, 0.003254489, 0.003093967, 0.002866569, 0.002557038, 
    0.002398103, 0.002352141, 0.002541754, 0.003015813, 0.003267439,
  0.004651412, 0.003974164, 0.004232773, 0.003774706, 0.004150323, 
    0.00447804, 0.004041263, 0.003963464, 0.004178569, 0.005855378, 
    0.005635452, 0.004752561, 0.004464049, 0.004185088, 0.004144765,
  0.003977223, 0.003846189, 0.003806909, 0.003709936, 0.004137252, 
    0.004236963, 0.003866463, 0.003913113, 0.003948994, 0.00458177, 
    0.00520255, 0.004409042, 0.003889269, 0.003508599, 0.00356225,
  0.003968964, 0.003864472, 0.003740528, 0.003599783, 0.003764995, 
    0.00363753, 0.003799123, 0.003827536, 0.003881744, 0.003979273, 
    0.00436048, 0.003949197, 0.003620218, 0.003278836, 0.003233419,
  0.003859699, 0.003843043, 0.003678062, 0.003696886, 0.003582262, 
    0.003691157, 0.003620993, 0.003675976, 0.003735898, 0.003832164, 
    0.003893199, 0.003716753, 0.00337172, 0.003124437, 0.003078873,
  0.003645729, 0.003626011, 0.003641182, 0.003582121, 0.003512276, 
    0.003511278, 0.00368554, 0.003534575, 0.003544625, 0.003784693, 
    0.003739335, 0.00354599, 0.003236367, 0.003032596, 0.003014948,
  0.003620132, 0.003647493, 0.003655936, 0.003511527, 0.003477886, 
    0.003543543, 0.003620464, 0.003615555, 0.003606891, 0.00364851, 
    0.003591746, 0.003366055, 0.00309458, 0.002907549, 0.00303193,
  0.004014716, 0.003992471, 0.003722949, 0.003511009, 0.003484266, 
    0.003495716, 0.003614116, 0.003632787, 0.003587936, 0.003539426, 
    0.003408467, 0.003164991, 0.002897528, 0.002769571, 0.002753141,
  0.004144042, 0.004026317, 0.003656528, 0.003496232, 0.003462713, 
    0.003500608, 0.003591717, 0.003580174, 0.003570342, 0.003518101, 
    0.003280558, 0.002956922, 0.002748806, 0.002703466, 0.002781146,
  0.004071941, 0.003825642, 0.003581631, 0.003523861, 0.003492948, 
    0.003534228, 0.003590858, 0.003596156, 0.003573106, 0.003404017, 
    0.003038697, 0.00281498, 0.002735224, 0.002934718, 0.003010811,
  0.004061535, 0.003902613, 0.003620504, 0.003603724, 0.003644962, 
    0.003631821, 0.003588185, 0.003526682, 0.003395526, 0.003070162, 
    0.002772018, 0.002702198, 0.003054029, 0.003352098, 0.003469491,
  0.006528313, 0.00526787, 0.006091077, 0.004491266, 0.004406638, 
    0.004444389, 0.0041456, 0.004095568, 0.004384747, 0.005541279, 
    0.006305137, 0.006005729, 0.005834167, 0.004920316, 0.004343819,
  0.004256694, 0.004182772, 0.004113325, 0.0039147, 0.004095772, 0.003830702, 
    0.003698929, 0.003760457, 0.003801082, 0.004105416, 0.005065346, 
    0.004737635, 0.004801223, 0.004499238, 0.004239298,
  0.004117718, 0.004017309, 0.003861938, 0.003707784, 0.00377665, 
    0.003358073, 0.003343109, 0.003290634, 0.003516922, 0.003595208, 
    0.003899058, 0.003977385, 0.004010956, 0.00409036, 0.004020117,
  0.003953766, 0.003774997, 0.003580177, 0.003441629, 0.003331664, 
    0.003329653, 0.003104954, 0.003158053, 0.003263071, 0.00332229, 
    0.003553327, 0.003711967, 0.003820917, 0.003841335, 0.003755915,
  0.00360228, 0.003469837, 0.003421544, 0.003397403, 0.003321832, 
    0.003263413, 0.003147263, 0.002912031, 0.002866863, 0.003249204, 
    0.003231746, 0.00350401, 0.003728668, 0.003701167, 0.003596552,
  0.003557546, 0.003606831, 0.003603383, 0.00346614, 0.003384326, 
    0.003429625, 0.003472789, 0.003422934, 0.003317625, 0.003202993, 
    0.003201464, 0.003384435, 0.003637643, 0.003622391, 0.003492506,
  0.003675473, 0.003729044, 0.003628377, 0.003471536, 0.003450444, 
    0.003423989, 0.003521452, 0.003576518, 0.003559545, 0.003438844, 
    0.003394204, 0.003450501, 0.003610282, 0.003539144, 0.003421667,
  0.003857005, 0.003608497, 0.003611489, 0.003519512, 0.003468557, 
    0.003441432, 0.003536551, 0.003602629, 0.003607588, 0.003604402, 
    0.003542873, 0.003542195, 0.003590715, 0.003439088, 0.003222986,
  0.003509229, 0.003816601, 0.003643135, 0.003581417, 0.003455492, 
    0.003493522, 0.003567609, 0.003635272, 0.003661984, 0.003629792, 
    0.003592377, 0.003594813, 0.003541498, 0.003285243, 0.003102438,
  0.003687562, 0.003879077, 0.003761601, 0.003550166, 0.003564735, 
    0.003625246, 0.003551885, 0.003635004, 0.003672707, 0.003630876, 
    0.003599564, 0.003551626, 0.003403991, 0.003174417, 0.003077863,
  0.003797268, 0.003768719, 0.00428535, 0.003933571, 0.00406978, 0.004521029, 
    0.004296311, 0.004246464, 0.004345674, 0.005834336, 0.006568232, 
    0.006531525, 0.007065004, 0.00680187, 0.005909367,
  0.003824772, 0.003811854, 0.003893779, 0.003786735, 0.004276691, 
    0.004328167, 0.004041849, 0.004056883, 0.004062954, 0.004449677, 
    0.005355439, 0.004845622, 0.005095398, 0.005693929, 0.005630817,
  0.003897174, 0.00386021, 0.003795813, 0.003746842, 0.004101778, 
    0.003853149, 0.003928494, 0.0038764, 0.003877855, 0.003907633, 
    0.004176721, 0.004090431, 0.004099742, 0.00442567, 0.004814136,
  0.003772102, 0.00368972, 0.003584573, 0.003621996, 0.00361039, 0.003862736, 
    0.003590423, 0.003659681, 0.003611026, 0.003643752, 0.003675866, 
    0.003666993, 0.003801126, 0.003903294, 0.004064377,
  0.003680364, 0.003575217, 0.00343858, 0.003416253, 0.003340037, 
    0.003419536, 0.003531603, 0.003321982, 0.003120666, 0.003428919, 
    0.003412595, 0.00336554, 0.003526542, 0.003766593, 0.003882392,
  0.003791316, 0.003474897, 0.003450199, 0.003373202, 0.003324304, 
    0.003355903, 0.00341718, 0.003426072, 0.003378577, 0.003249917, 
    0.00317999, 0.003141838, 0.003322686, 0.003702252, 0.003752034,
  0.003739352, 0.003434288, 0.003509094, 0.003394401, 0.003386662, 
    0.00338942, 0.003413571, 0.003398827, 0.003391803, 0.00324474, 
    0.003209475, 0.003181953, 0.003266077, 0.003621038, 0.0037362,
  0.003744011, 0.003528888, 0.003541989, 0.003421327, 0.003382198, 
    0.003432039, 0.003411111, 0.003358061, 0.003464996, 0.003360403, 
    0.003368237, 0.003412163, 0.003556643, 0.003667732, 0.003684111,
  0.0034511, 0.003659027, 0.003527536, 0.003474434, 0.003446637, 0.003456572, 
    0.003534402, 0.003601565, 0.00362511, 0.00361475, 0.003598635, 
    0.003573923, 0.003599278, 0.003579868, 0.00343827,
  0.003389167, 0.003651994, 0.003570351, 0.003512242, 0.003577911, 
    0.003554711, 0.003464933, 0.003449074, 0.003576697, 0.003618674, 
    0.003574216, 0.003563882, 0.003536892, 0.00337072, 0.00320932,
  0.003733405, 0.003605075, 0.003602934, 0.003319036, 0.003425287, 
    0.003528783, 0.003366405, 0.003352433, 0.003426629, 0.003798881, 
    0.00402482, 0.004093037, 0.004298054, 0.004656576, 0.005217423,
  0.003709339, 0.003552347, 0.003385196, 0.003301159, 0.003395648, 
    0.003384573, 0.003259423, 0.003345854, 0.003405832, 0.003596157, 
    0.003907762, 0.003927755, 0.003968508, 0.004121465, 0.004470911,
  0.00380134, 0.003462567, 0.003313386, 0.003208558, 0.003166625, 
    0.003090569, 0.003243809, 0.00334046, 0.003392398, 0.003397319, 
    0.003576059, 0.003807105, 0.003821456, 0.003893076, 0.004151531,
  0.004075019, 0.003645386, 0.003484328, 0.003131071, 0.003196563, 
    0.003079101, 0.003115917, 0.003272906, 0.00322922, 0.003326416, 
    0.003636717, 0.003796761, 0.003809989, 0.00381616, 0.003913225,
  0.004197241, 0.003972064, 0.003378728, 0.003102351, 0.003141875, 
    0.003299714, 0.003218172, 0.003004161, 0.00296821, 0.003372368, 
    0.003732172, 0.003825726, 0.003814204, 0.003798617, 0.003849152,
  0.004286928, 0.004108909, 0.003590101, 0.003407062, 0.003362402, 
    0.003378297, 0.003405674, 0.003167744, 0.003124773, 0.003477318, 
    0.003777725, 0.003811812, 0.003801339, 0.003847765, 0.003898275,
  0.004177825, 0.003889229, 0.003612535, 0.003434359, 0.003422202, 
    0.003394906, 0.003396441, 0.003309485, 0.003359962, 0.003558249, 
    0.003706011, 0.00375459, 0.003725548, 0.00374225, 0.003731537,
  0.004015086, 0.003364007, 0.003428434, 0.003446886, 0.003453798, 
    0.003431936, 0.003472481, 0.003406643, 0.003522576, 0.003629529, 
    0.003736774, 0.003720136, 0.003650817, 0.003626627, 0.003606127,
  0.003653858, 0.003522151, 0.003512588, 0.00349022, 0.003490684, 
    0.003456989, 0.003522073, 0.003523329, 0.003580209, 0.003666971, 
    0.003726478, 0.003698716, 0.003600632, 0.003525403, 0.003469937,
  0.003666021, 0.003514032, 0.003568191, 0.003534216, 0.003493497, 
    0.003500598, 0.003446056, 0.00350593, 0.003419542, 0.003626061, 
    0.003679344, 0.003651808, 0.003550004, 0.003446834, 0.003431701,
  0.004837724, 0.004692601, 0.006111139, 0.004626386, 0.004693931, 
    0.005593006, 0.004472414, 0.004112347, 0.004094479, 0.004654168, 
    0.004473598, 0.004045814, 0.003989719, 0.004057277, 0.004223429,
  0.003977145, 0.00408721, 0.004301192, 0.004217466, 0.004936396, 
    0.004617619, 0.003890807, 0.003802735, 0.003756912, 0.003913513, 
    0.0040734, 0.003813071, 0.003706226, 0.003818189, 0.004064944,
  0.003873046, 0.003990192, 0.003989534, 0.003930838, 0.004129092, 
    0.003669231, 0.003659521, 0.003582219, 0.003522594, 0.003505645, 
    0.003628293, 0.003686792, 0.003549779, 0.003634477, 0.003948524,
  0.00364435, 0.003692391, 0.003667753, 0.00366451, 0.003610672, 0.003603637, 
    0.003353795, 0.003410565, 0.003358395, 0.003395263, 0.003627887, 
    0.003609745, 0.003396054, 0.003587947, 0.003897787,
  0.003509503, 0.003437229, 0.003356514, 0.00338165, 0.003391364, 
    0.003480557, 0.003341467, 0.003061729, 0.002913338, 0.003392623, 
    0.00362847, 0.003524791, 0.00336545, 0.003566266, 0.003618636,
  0.003475478, 0.00334505, 0.003331879, 0.003344346, 0.00331229, 0.003342269, 
    0.003395281, 0.00319466, 0.003225733, 0.003539335, 0.003522871, 
    0.003533294, 0.003394705, 0.003548868, 0.003537155,
  0.003461898, 0.003307765, 0.003309801, 0.003315689, 0.003317915, 
    0.003332324, 0.003323993, 0.003373385, 0.003449676, 0.003511597, 
    0.003534186, 0.003520784, 0.003418922, 0.00345906, 0.003473134,
  0.003505071, 0.003221611, 0.003321157, 0.003296124, 0.003289122, 
    0.003247411, 0.003184507, 0.003160188, 0.003472193, 0.003545571, 
    0.003588906, 0.003480007, 0.003398788, 0.00350488, 0.003448412,
  0.003621781, 0.00349292, 0.003460904, 0.003439093, 0.003349918, 
    0.003276612, 0.003171873, 0.00316572, 0.003465204, 0.00359694, 
    0.003494621, 0.003407879, 0.003478816, 0.003509799, 0.00345942,
  0.003582309, 0.003544456, 0.003534077, 0.003508355, 0.003388566, 
    0.003364061, 0.003084685, 0.003167444, 0.003429565, 0.003295234, 
    0.003450447, 0.003420065, 0.003265726, 0.003458113, 0.00333579,
  0.003855289, 0.003945656, 0.004564035, 0.004004606, 0.004329359, 
    0.005993624, 0.005129867, 0.005063323, 0.00551952, 0.00931668, 
    0.00861134, 0.006841415, 0.00583503, 0.00507152, 0.004798797,
  0.003755238, 0.003883244, 0.003986083, 0.00391839, 0.005060511, 
    0.006224781, 0.00443305, 0.00445823, 0.004643641, 0.006141597, 
    0.007954011, 0.00550977, 0.004678096, 0.004703329, 0.00458598,
  0.003638122, 0.003818526, 0.004013005, 0.003912694, 0.004809811, 
    0.004648738, 0.004461102, 0.004075918, 0.004161717, 0.004563871, 
    0.005082532, 0.004516353, 0.004135147, 0.003996288, 0.004130342,
  0.003489723, 0.003679475, 0.003811918, 0.00397632, 0.003993939, 
    0.004951133, 0.004218844, 0.004053088, 0.003985474, 0.004059883, 
    0.004108961, 0.003975621, 0.003794435, 0.003693335, 0.003944161,
  0.003377462, 0.003465407, 0.003653508, 0.00372458, 0.003692659, 
    0.003956163, 0.004197345, 0.004318238, 0.004376594, 0.004428461, 
    0.003906073, 0.00383046, 0.003631303, 0.003605479, 0.003702424,
  0.00326587, 0.003382175, 0.003430818, 0.003571256, 0.003574607, 
    0.003709141, 0.003909198, 0.004055106, 0.004439919, 0.004023845, 
    0.003816549, 0.00365453, 0.003546176, 0.003534647, 0.003422322,
  0.003290004, 0.003323911, 0.003268599, 0.003424658, 0.003529276, 
    0.003572982, 0.003663416, 0.003866889, 0.003852171, 0.003701698, 
    0.003671698, 0.003600375, 0.003497001, 0.00342697, 0.003311712,
  0.003458063, 0.003299872, 0.003184594, 0.003329211, 0.003418531, 
    0.003504819, 0.003554154, 0.003670917, 0.003663389, 0.003631869, 
    0.003583187, 0.00348914, 0.003453467, 0.003371556, 0.003329176,
  0.00361955, 0.003302894, 0.003165669, 0.003232981, 0.003302942, 
    0.003373879, 0.003541681, 0.003640155, 0.003612692, 0.003564109, 
    0.00347511, 0.003393287, 0.003328393, 0.003333658, 0.003443307,
  0.003663944, 0.003517177, 0.003129216, 0.003178922, 0.003222178, 
    0.003288272, 0.003396096, 0.003498699, 0.003503521, 0.003428845, 
    0.003314585, 0.003232606, 0.00316272, 0.003266587, 0.003405401,
  0.003685011, 0.003879458, 0.004269832, 0.003945498, 0.004605622, 
    0.005713613, 0.004925458, 0.004945342, 0.005555459, 0.01079451, 
    0.01104336, 0.009472773, 0.009699243, 0.008324606, 0.007469548,
  0.003593748, 0.003619878, 0.00370472, 0.003870196, 0.004932858, 
    0.005224013, 0.004013399, 0.004271525, 0.004294327, 0.006143617, 
    0.01034843, 0.007922011, 0.006907204, 0.008235756, 0.007086581,
  0.003408382, 0.003469625, 0.003605745, 0.003610117, 0.003935212, 
    0.00393946, 0.004282555, 0.003988026, 0.004043411, 0.004287405, 
    0.005557167, 0.005189542, 0.004904166, 0.00557052, 0.005966696,
  0.00333759, 0.003310634, 0.00336197, 0.003520059, 0.003471625, 0.003904599, 
    0.003913743, 0.0042893, 0.00399452, 0.004017107, 0.00425638, 0.004499582, 
    0.004201565, 0.004719961, 0.005239985,
  0.00336465, 0.003188058, 0.003210372, 0.003414421, 0.003364896, 
    0.003419853, 0.003707448, 0.003980679, 0.004379422, 0.004789571, 
    0.003982256, 0.004113233, 0.004090056, 0.004178906, 0.004316712,
  0.003406653, 0.003240013, 0.003143536, 0.003378296, 0.003313791, 
    0.00334976, 0.00343273, 0.003577499, 0.004063977, 0.00404483, 
    0.004431411, 0.004001676, 0.003951963, 0.003940624, 0.004011942,
  0.003598749, 0.003390792, 0.003115222, 0.003355924, 0.003321134, 
    0.003337053, 0.003374861, 0.003497845, 0.003586513, 0.003697615, 
    0.003840206, 0.003934927, 0.003876776, 0.003843362, 0.003861466,
  0.003656671, 0.003521736, 0.003104179, 0.003329327, 0.003294171, 
    0.003331043, 0.003377794, 0.003489336, 0.00359736, 0.003712142, 
    0.003780954, 0.003831114, 0.003837934, 0.003794062, 0.003784593,
  0.003816271, 0.003412215, 0.003076857, 0.003337678, 0.003331289, 
    0.003266655, 0.00340015, 0.003568341, 0.003680429, 0.003761227, 
    0.003792219, 0.003798687, 0.003788329, 0.003747658, 0.003748578,
  0.003905533, 0.003383199, 0.003130707, 0.003325296, 0.003336754, 
    0.003308287, 0.003363923, 0.003532497, 0.003673096, 0.003765515, 
    0.003802769, 0.003767986, 0.003732257, 0.003704884, 0.003748195,
  0.003850346, 0.00404425, 0.004991103, 0.004737658, 0.005380753, 
    0.006601301, 0.0051316, 0.005030091, 0.006580524, 0.01119078, 0.01150998, 
    0.01029137, 0.01129228, 0.01041108, 0.01013341,
  0.003724327, 0.003785484, 0.004031555, 0.004642287, 0.006404015, 
    0.006151134, 0.004434456, 0.004538123, 0.005075237, 0.006889544, 
    0.01095957, 0.007584006, 0.006963092, 0.0108165, 0.01017104,
  0.003672775, 0.003730277, 0.003788477, 0.003958452, 0.004822031, 
    0.00426187, 0.00440153, 0.004223675, 0.004430359, 0.004668441, 
    0.005612204, 0.005422794, 0.004791189, 0.005706744, 0.008170893,
  0.003591676, 0.00359688, 0.003567605, 0.003661535, 0.00384321, 0.004609004, 
    0.004086253, 0.004298786, 0.004022995, 0.00406803, 0.004144238, 
    0.004114322, 0.004123753, 0.004546187, 0.006688714,
  0.003594699, 0.003467497, 0.003422292, 0.003405982, 0.003402457, 
    0.003693526, 0.004222478, 0.004179848, 0.004007407, 0.004106039, 
    0.003904185, 0.003903655, 0.003927322, 0.003938755, 0.004456148,
  0.003626887, 0.003518897, 0.003260115, 0.003253625, 0.003257057, 
    0.003346866, 0.00349209, 0.003652036, 0.003707305, 0.003712484, 
    0.003912199, 0.003731989, 0.003805955, 0.003813225, 0.003878187,
  0.003713483, 0.00383728, 0.003324896, 0.003183759, 0.0031215, 0.003179289, 
    0.003248258, 0.00335573, 0.003370908, 0.003422009, 0.003502179, 
    0.003663321, 0.003696759, 0.003728866, 0.003760961,
  0.004015473, 0.004182907, 0.003642043, 0.003144759, 0.003014605, 
    0.003065328, 0.003077911, 0.003186986, 0.003243014, 0.003391919, 
    0.003470297, 0.003590264, 0.003618427, 0.003627426, 0.003705938,
  0.00405049, 0.003755702, 0.003515343, 0.003346521, 0.002894508, 
    0.002828786, 0.002941168, 0.003039374, 0.003142113, 0.003232021, 
    0.003354044, 0.00347393, 0.003510299, 0.003562666, 0.003640904,
  0.004198946, 0.004055617, 0.003681662, 0.003423079, 0.003183301, 
    0.002851529, 0.002824774, 0.002898844, 0.002985392, 0.003094113, 
    0.003191799, 0.003284679, 0.003347973, 0.003431258, 0.003565686,
  0.004023871, 0.004105258, 0.004351567, 0.004038975, 0.004611154, 
    0.005942853, 0.005094214, 0.005190107, 0.006138201, 0.01105648, 
    0.01121232, 0.01028356, 0.01120334, 0.01036802, 0.01037729,
  0.003910614, 0.00403764, 0.0040758, 0.004021073, 0.005849987, 0.00656944, 
    0.00450231, 0.004893174, 0.00546834, 0.006829595, 0.01086233, 
    0.007792918, 0.00812799, 0.01080112, 0.01069372,
  0.00395435, 0.004088139, 0.00413138, 0.004159377, 0.005885946, 0.004599595, 
    0.004713749, 0.00448954, 0.004879147, 0.005244444, 0.00642986, 
    0.00669763, 0.005803511, 0.006139253, 0.009217522,
  0.00392467, 0.003927086, 0.004067918, 0.004331164, 0.004671389, 
    0.005613855, 0.004473573, 0.00502964, 0.004633381, 0.004676378, 
    0.004865831, 0.005042133, 0.004738844, 0.005077135, 0.007078908,
  0.003795662, 0.00372616, 0.003796139, 0.003916365, 0.003987591, 
    0.004591019, 0.004985896, 0.004778714, 0.005001607, 0.005257593, 
    0.00456077, 0.004595912, 0.004515543, 0.004467403, 0.004932785,
  0.003938273, 0.003597276, 0.00354519, 0.003569922, 0.003685047, 
    0.003989304, 0.004477633, 0.00472686, 0.005789388, 0.005105447, 
    0.004993484, 0.00437089, 0.004280351, 0.004184009, 0.004182503,
  0.003929187, 0.00354265, 0.003365789, 0.003367235, 0.003555988, 
    0.003697169, 0.003935373, 0.004272341, 0.004529286, 0.004218505, 
    0.004224596, 0.004133691, 0.00409587, 0.004058583, 0.00401845,
  0.00386844, 0.00356233, 0.00329054, 0.003249667, 0.003355109, 0.003573809, 
    0.003612873, 0.003890421, 0.00406429, 0.00403075, 0.004034976, 
    0.003951485, 0.003920003, 0.003869516, 0.003955847,
  0.003811145, 0.003679619, 0.003362873, 0.003177135, 0.0031367, 0.003303402, 
    0.003515891, 0.003697933, 0.003792387, 0.003822026, 0.003842022, 
    0.00379274, 0.003733392, 0.003678499, 0.003758931,
  0.00402038, 0.003992262, 0.003465307, 0.003323159, 0.003123809, 
    0.003073641, 0.003269169, 0.003459828, 0.00357319, 0.003633407, 
    0.003647032, 0.003586128, 0.00352853, 0.003474938, 0.003514434,
  0.003866677, 0.00391637, 0.004193766, 0.003958089, 0.004047876, 
    0.004213444, 0.003865599, 0.004004826, 0.004466728, 0.01091296, 
    0.01079896, 0.009519359, 0.01001713, 0.009369325, 0.009040846,
  0.003861233, 0.003895503, 0.004031448, 0.003939218, 0.004246192, 
    0.004353972, 0.0039759, 0.004067258, 0.004268444, 0.006494997, 
    0.01044801, 0.008033818, 0.007955531, 0.009642051, 0.009411842,
  0.003862004, 0.003986234, 0.004136659, 0.003949569, 0.004265129, 
    0.003950498, 0.004240151, 0.0041195, 0.004114913, 0.005277447, 
    0.006928584, 0.006891948, 0.005837682, 0.005365967, 0.008551666,
  0.003781697, 0.003848037, 0.004058294, 0.004099178, 0.004035166, 
    0.00457739, 0.004228771, 0.004576492, 0.004151735, 0.00460432, 
    0.004982912, 0.004954162, 0.004810101, 0.005079193, 0.007121265,
  0.003710749, 0.003687725, 0.00377256, 0.003994837, 0.003893207, 
    0.003965132, 0.004650872, 0.004510793, 0.00467959, 0.005180036, 
    0.00455155, 0.004537554, 0.004587272, 0.004525877, 0.004733809,
  0.00398071, 0.00357186, 0.003593774, 0.003603137, 0.003757707, 0.003799586, 
    0.003935449, 0.004277907, 0.005588823, 0.005216605, 0.005238127, 
    0.004420199, 0.004364324, 0.004396567, 0.004218682,
  0.003664025, 0.00347523, 0.003482223, 0.003479981, 0.00361751, 0.00375302, 
    0.00385537, 0.004004628, 0.00429818, 0.004175764, 0.00434884, 
    0.004338165, 0.00424852, 0.004287458, 0.004174955,
  0.003511115, 0.003403017, 0.003359486, 0.003412195, 0.003488892, 
    0.003621625, 0.003696038, 0.003881705, 0.004055026, 0.004130019, 
    0.004161078, 0.004233522, 0.004173432, 0.004230306, 0.00419153,
  0.003577895, 0.003389717, 0.00330505, 0.003299642, 0.003354367, 
    0.003473219, 0.003659618, 0.003852679, 0.004001212, 0.004088083, 
    0.004113615, 0.004112953, 0.004141281, 0.004141227, 0.004180904,
  0.003801725, 0.003451837, 0.003317756, 0.003286403, 0.003297613, 
    0.003354308, 0.003638913, 0.003793674, 0.003924753, 0.004021948, 
    0.004113134, 0.004074271, 0.004051307, 0.003994623, 0.004133043,
  0.003909171, 0.003728815, 0.003930378, 0.003840366, 0.003752419, 
    0.003893807, 0.003725272, 0.003675812, 0.003747024, 0.006361892, 
    0.008897002, 0.008174461, 0.007903298, 0.007708987, 0.007782138,
  0.003905132, 0.003797938, 0.00376686, 0.003762352, 0.003880844, 
    0.003908335, 0.003722216, 0.003702999, 0.003682997, 0.004656288, 
    0.0083287, 0.007118522, 0.0068936, 0.007750343, 0.008034582,
  0.003994422, 0.003933364, 0.00391358, 0.003814889, 0.003954625, 
    0.003748467, 0.003931739, 0.003789994, 0.003778189, 0.00412533, 
    0.0060497, 0.006499897, 0.005392725, 0.005108977, 0.00753658,
  0.004122571, 0.003875389, 0.003809693, 0.003859311, 0.003846598, 
    0.004070425, 0.003856268, 0.004115009, 0.003970113, 0.004146488, 
    0.004513535, 0.00446529, 0.004198572, 0.005049737, 0.007027236,
  0.004120284, 0.003712169, 0.00371992, 0.003926433, 0.003759906, 
    0.003854691, 0.004321751, 0.004103151, 0.004297956, 0.004772096, 
    0.004122849, 0.004106523, 0.003979817, 0.004336783, 0.004707993,
  0.004218637, 0.003573445, 0.00359999, 0.003685929, 0.003733861, 
    0.003735736, 0.003725303, 0.00400801, 0.005006844, 0.0050496, 
    0.004773432, 0.00407314, 0.003987845, 0.004074575, 0.004129449,
  0.004041937, 0.003445518, 0.003485426, 0.003509095, 0.00370388, 
    0.003750538, 0.003670094, 0.003694767, 0.003955889, 0.004177605, 
    0.004076072, 0.003972908, 0.004051998, 0.004062969, 0.004086233,
  0.003882741, 0.003373286, 0.00341171, 0.003478165, 0.003548617, 0.00370028, 
    0.003549418, 0.003603323, 0.003839894, 0.004020141, 0.004002954, 
    0.004062068, 0.004086454, 0.003997829, 0.003922372,
  0.003933262, 0.003317531, 0.003333692, 0.003419057, 0.003441741, 
    0.003501674, 0.00348403, 0.003644736, 0.003832595, 0.003957141, 
    0.003953471, 0.004055496, 0.004047768, 0.00406031, 0.004135339,
  0.004019734, 0.003424104, 0.003283049, 0.003303637, 0.003422029, 
    0.003444012, 0.003555438, 0.003656062, 0.003797261, 0.003868585, 
    0.003997931, 0.004008973, 0.003983081, 0.003980203, 0.004209472,
  0.004064866, 0.003875114, 0.004095922, 0.003716289, 0.003636429, 
    0.003557174, 0.003346733, 0.003353163, 0.003468577, 0.004216614, 
    0.005545596, 0.007156952, 0.007971506, 0.007918334, 0.007907867,
  0.003979325, 0.003852707, 0.003837878, 0.003702823, 0.003651657, 
    0.003544864, 0.003320152, 0.003381945, 0.003436325, 0.003922211, 
    0.005138685, 0.006587908, 0.00716678, 0.007776647, 0.007951519,
  0.004075447, 0.004073229, 0.004020643, 0.003720186, 0.003667325, 
    0.003440979, 0.003302024, 0.003367505, 0.003506302, 0.003702638, 
    0.004761968, 0.006250926, 0.005770283, 0.005487892, 0.007124272,
  0.004306993, 0.004236782, 0.004041594, 0.003810883, 0.003533963, 
    0.003393579, 0.003289989, 0.003551132, 0.00351246, 0.003849357, 
    0.003875281, 0.004169865, 0.004402518, 0.00518429, 0.00646593,
  0.004459398, 0.004266905, 0.003871469, 0.003502465, 0.003308592, 
    0.003302228, 0.00340531, 0.003160332, 0.003365658, 0.004119575, 
    0.003914501, 0.003758822, 0.004161495, 0.004660011, 0.005063234,
  0.004567116, 0.004130423, 0.003596196, 0.003357707, 0.003299495, 
    0.003299413, 0.003363166, 0.003381141, 0.003570936, 0.003905605, 
    0.004117053, 0.003670906, 0.003961579, 0.004301138, 0.004579076,
  0.004390055, 0.003948854, 0.003656586, 0.003489124, 0.003510689, 
    0.003499595, 0.003437543, 0.003373174, 0.003353406, 0.003458925, 
    0.003618838, 0.003683021, 0.003951904, 0.004166996, 0.004289485,
  0.004226296, 0.004075443, 0.003756311, 0.003585269, 0.003540652, 
    0.003546117, 0.003462834, 0.003419703, 0.003368813, 0.003464537, 
    0.003580344, 0.003713115, 0.003941125, 0.004065525, 0.004116254,
  0.004338141, 0.004168054, 0.003723569, 0.00352681, 0.003461333, 
    0.003423512, 0.003353768, 0.003491334, 0.003487228, 0.003573862, 
    0.003614001, 0.003724499, 0.003857281, 0.004002362, 0.004241135,
  0.004436906, 0.004290433, 0.003685254, 0.003436793, 0.003469037, 
    0.003359029, 0.003391381, 0.003474202, 0.003474073, 0.003697004, 
    0.003712084, 0.003750931, 0.003839497, 0.003950357, 0.004315779,
  0.003914619, 0.003871237, 0.003867427, 0.003653501, 0.003575881, 
    0.003343848, 0.003227726, 0.003412024, 0.003680477, 0.004690233, 
    0.006939432, 0.007945639, 0.00873948, 0.009152628, 0.009537729,
  0.004039139, 0.003869885, 0.003802045, 0.003612559, 0.00369036, 
    0.003416413, 0.003252866, 0.003267246, 0.003551546, 0.00404494, 
    0.006220207, 0.007215368, 0.007461271, 0.008960775, 0.009362794,
  0.004157203, 0.004035825, 0.003987421, 0.003730637, 0.003601213, 
    0.00326656, 0.003254301, 0.003243784, 0.00341423, 0.003700785, 
    0.004852145, 0.006441742, 0.006070239, 0.00535595, 0.007699552,
  0.004434297, 0.004212331, 0.003997938, 0.003950467, 0.003688953, 
    0.003321735, 0.003038352, 0.003180022, 0.003224182, 0.003433061, 
    0.003610718, 0.004015783, 0.004141239, 0.00485939, 0.006756961,
  0.004585173, 0.004341973, 0.004037062, 0.003828758, 0.003518979, 
    0.003366826, 0.003158514, 0.002978744, 0.002953495, 0.003230783, 
    0.003463991, 0.003615703, 0.00396694, 0.004412157, 0.005089546,
  0.004504573, 0.004377133, 0.004123049, 0.003832836, 0.003620841, 
    0.003477279, 0.003334162, 0.003164869, 0.003141739, 0.003138134, 
    0.003265288, 0.003450186, 0.00375384, 0.004052563, 0.004675598,
  0.004287852, 0.004310204, 0.003964846, 0.003752275, 0.003724232, 
    0.003698251, 0.003560559, 0.003346474, 0.003286002, 0.003110623, 
    0.00306238, 0.003301208, 0.003628566, 0.003885286, 0.004177291,
  0.003900056, 0.004050318, 0.003802713, 0.003645574, 0.003625094, 
    0.003683025, 0.00361888, 0.003533996, 0.003448843, 0.003306027, 
    0.003142396, 0.003195352, 0.003532556, 0.003760111, 0.003965139,
  0.003708094, 0.003716772, 0.003618621, 0.003543385, 0.003482637, 
    0.003504047, 0.003484118, 0.003543298, 0.003575483, 0.003412887, 
    0.003241214, 0.003194373, 0.003409244, 0.003693517, 0.004018453,
  0.003672285, 0.003650319, 0.003556414, 0.003528291, 0.003512886, 
    0.003417205, 0.003394474, 0.003506209, 0.003546659, 0.003530687, 
    0.003397214, 0.003247583, 0.003393465, 0.003651729, 0.004123297 ;

 land_mask =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  1.541242e-05, 2.149244e-05, 1.789696e-05, 3.449073e-05, 2.898845e-05, 
    1.512394e-05, 1.853227e-05, 2.058743e-05, 1.964916e-05, 5.417909e-06, 
    6.469748e-06, 8.294474e-06, 4.556026e-06, 4.174302e-06, 8.112652e-07,
  3.304964e-05, 2.855557e-05, 2.48103e-05, 3.996154e-05, 2.033398e-05, 
    1.540473e-05, 2.119337e-05, 1.839629e-05, 2.010591e-05, 1.204061e-05, 
    9.248628e-06, 1.643999e-05, 1.432952e-05, 3.740712e-06, 6.340566e-07,
  2.534045e-05, 2.754723e-05, 3.171658e-05, 3.572768e-05, 2.471734e-05, 
    2.096064e-06, 1.998213e-05, 1.67057e-05, 1.929956e-05, 1.896231e-05, 
    1.636189e-05, 2.006903e-05, 2.098643e-05, 1.281043e-05, 5.704926e-06,
  3.098029e-05, 2.329577e-05, 2.966183e-05, 3.702644e-05, 3.815746e-05, 
    1.704895e-05, 2.312034e-06, 1.615273e-05, 2.379888e-05, 1.880619e-05, 
    1.717348e-05, 2.036215e-05, 2.227437e-05, 1.931813e-05, 1.215085e-05,
  5.019759e-05, 3.128999e-05, 3.013168e-05, 3.177963e-05, 3.684043e-05, 
    3.744761e-05, 2.050868e-05, 3.039537e-06, 6.722388e-06, 9.672612e-06, 
    1.475029e-05, 1.818954e-05, 2.200485e-05, 2.437644e-05, 1.912651e-05,
  5.403291e-05, 4.348331e-05, 3.468652e-05, 3.491564e-05, 3.3709e-05, 
    3.53848e-05, 3.447505e-05, 2.461184e-05, 1.636995e-05, 1.600544e-05, 
    1.260528e-05, 1.895299e-05, 2.190742e-05, 2.607091e-05, 2.208986e-05,
  5.01689e-05, 4.673811e-05, 3.903202e-05, 3.838182e-05, 3.828103e-05, 
    3.800392e-05, 3.834345e-05, 3.748023e-05, 3.334786e-05, 3.21458e-05, 
    2.53297e-05, 2.12881e-05, 2.228568e-05, 2.52427e-05, 2.482493e-05,
  5.790083e-05, 4.494716e-05, 3.954942e-05, 4.051331e-05, 3.755954e-05, 
    3.961224e-05, 4.153988e-05, 3.96587e-05, 3.895505e-05, 3.826829e-05, 
    3.429255e-05, 2.26958e-05, 2.379993e-05, 2.567318e-05, 2.399821e-05,
  4.721759e-05, 4.113105e-05, 3.815673e-05, 4.024105e-05, 3.708599e-05, 
    3.644662e-05, 3.709995e-05, 4.082697e-05, 4.040192e-05, 4.171166e-05, 
    3.637889e-05, 2.57895e-05, 2.530864e-05, 2.473353e-05, 1.735654e-05,
  3.364938e-05, 3.401121e-05, 3.603425e-05, 3.531952e-05, 3.373628e-05, 
    3.501731e-05, 3.616545e-05, 3.476049e-05, 2.928733e-05, 1.872777e-05, 
    2.544651e-05, 2.473375e-05, 2.280703e-05, 2.2938e-05, 1.901704e-05,
  1.76077e-05, 2.864065e-05, 1.776834e-05, 3.148875e-05, 1.508937e-05, 
    7.106938e-06, 2.181913e-05, 2.782342e-05, 3.137803e-05, 3.520778e-05, 
    4.732734e-05, 6.401946e-05, 5.233364e-05, 2.89776e-05, 2.358943e-05,
  4.307582e-05, 4.057435e-05, 4.180562e-05, 2.543804e-05, 5.837779e-06, 
    3.058517e-06, 2.23636e-05, 2.730484e-05, 2.95197e-05, 3.580458e-05, 
    4.368949e-05, 6.172113e-05, 5.117038e-05, 2.675562e-05, 1.987387e-05,
  5.131335e-05, 5.417901e-05, 5.288439e-05, 4.300658e-05, 1.343086e-05, 
    3.457004e-07, 1.25697e-05, 2.788672e-05, 3.400298e-05, 3.627205e-05, 
    4.337105e-05, 5.520205e-05, 4.9348e-05, 2.86029e-05, 1.637547e-05,
  4.812831e-05, 5.133654e-05, 5.419298e-05, 5.286975e-05, 4.325551e-05, 
    1.41237e-05, 1.120472e-06, 1.395564e-05, 2.853648e-05, 3.594159e-05, 
    4.130859e-05, 4.7857e-05, 4.391781e-05, 3.278372e-05, 1.785635e-05,
  4.53042e-05, 5.034003e-05, 4.927324e-05, 4.875718e-05, 4.662075e-05, 
    4.112302e-05, 1.465915e-05, 1.945829e-06, 1.149936e-05, 2.568054e-05, 
    3.628296e-05, 4.258106e-05, 3.871245e-05, 2.953047e-05, 1.993626e-05,
  4.317964e-05, 4.63599e-05, 4.774864e-05, 4.832307e-05, 4.654443e-05, 
    4.591968e-05, 4.397864e-05, 3.67497e-05, 2.601861e-05, 2.856782e-05, 
    2.572462e-05, 3.661433e-05, 3.543294e-05, 2.57325e-05, 1.911987e-05,
  4.269351e-05, 4.499312e-05, 4.432832e-05, 4.543574e-05, 4.369643e-05, 
    4.319287e-05, 4.12421e-05, 3.823872e-05, 4.36662e-05, 4.025041e-05, 
    3.021921e-05, 3.083509e-05, 3.223219e-05, 2.487799e-05, 1.796996e-05,
  4.032556e-05, 4.450034e-05, 4.252103e-05, 4.576749e-05, 4.338922e-05, 
    4.022404e-05, 3.970858e-05, 3.855252e-05, 4.279742e-05, 4.217462e-05, 
    2.867606e-05, 2.352637e-05, 2.6028e-05, 2.34745e-05, 1.773227e-05,
  3.680445e-05, 3.8561e-05, 3.932453e-05, 4.008911e-05, 4.10592e-05, 
    4.242024e-05, 4.183842e-05, 4.25545e-05, 4.257812e-05, 4.113019e-05, 
    2.809104e-05, 1.796148e-05, 1.856431e-05, 1.771724e-05, 1.29635e-05,
  2.843303e-05, 3.07888e-05, 3.418518e-05, 3.619152e-05, 3.659911e-05, 
    3.608476e-05, 3.940264e-05, 4.082692e-05, 3.383959e-05, 2.009884e-05, 
    2.079521e-05, 1.416753e-05, 1.292397e-05, 1.170525e-05, 8.398287e-06,
  7.106108e-06, 3.670168e-05, 2.88846e-05, 2.202875e-05, 5.372665e-06, 
    1.350819e-06, 7.190079e-06, 1.132825e-05, 6.466976e-06, 3.321941e-06, 
    4.574737e-06, 5.205121e-06, 2.596597e-06, 2.163669e-06, 1.301985e-06,
  4.009838e-05, 3.509641e-05, 3.697587e-05, 2.820417e-05, 6.392709e-06, 
    6.295394e-07, 1.232776e-05, 1.453577e-05, 6.511846e-06, 7.562039e-06, 
    6.278542e-06, 1.045935e-05, 9.465883e-06, 1.30805e-06, 6.833992e-07,
  3.503971e-05, 3.417911e-05, 3.774076e-05, 3.748374e-05, 1.579207e-05, 
    1.184036e-06, 5.742508e-06, 1.46137e-05, 1.241755e-05, 1.337688e-05, 
    1.188243e-05, 1.271275e-05, 1.296508e-05, 4.735341e-06, 5.874992e-07,
  3.529558e-05, 3.386871e-05, 3.967529e-05, 4.145858e-05, 4.401032e-05, 
    1.389758e-05, 2.564483e-06, 8.944627e-06, 1.747162e-05, 1.942495e-05, 
    1.542892e-05, 1.26918e-05, 1.172026e-05, 8.336124e-06, 1.337085e-06,
  3.723596e-05, 3.666956e-05, 3.789528e-05, 4.137732e-05, 4.707062e-05, 
    4.249486e-05, 7.523884e-06, 2.050615e-06, 5.395336e-06, 1.15063e-05, 
    1.527645e-05, 1.421404e-05, 1.145178e-05, 7.691116e-06, 2.805901e-06,
  3.648175e-05, 3.707033e-05, 3.878397e-05, 4.180503e-05, 4.775535e-05, 
    4.881659e-05, 3.888029e-05, 2.997961e-05, 1.846556e-05, 2.206802e-05, 
    1.332975e-05, 1.529024e-05, 1.224978e-05, 6.190134e-06, 2.958833e-06,
  3.925908e-05, 4.129323e-05, 4.056869e-05, 4.317392e-05, 4.581196e-05, 
    4.981386e-05, 4.843214e-05, 4.989196e-05, 4.048089e-05, 3.314703e-05, 
    2.424715e-05, 1.76877e-05, 1.319223e-05, 6.311184e-06, 2.774854e-06,
  4.088867e-05, 4.21737e-05, 4.627809e-05, 4.676771e-05, 4.444002e-05, 
    4.957293e-05, 4.8714e-05, 5.927267e-05, 5.232033e-05, 4.109531e-05, 
    3.365188e-05, 2.267609e-05, 1.833405e-05, 7.386638e-06, 3.835118e-06,
  3.886756e-05, 4.237497e-05, 4.564897e-05, 4.671698e-05, 4.964941e-05, 
    4.870181e-05, 4.883225e-05, 5.750599e-05, 5.689275e-05, 4.763461e-05, 
    3.870661e-05, 2.895994e-05, 2.243406e-05, 1.501851e-05, 7.439327e-06,
  3.417029e-05, 4.132056e-05, 4.452689e-05, 4.569264e-05, 4.866045e-05, 
    5.059425e-05, 5.060138e-05, 5.159399e-05, 4.085731e-05, 3.639381e-05, 
    3.66254e-05, 2.962897e-05, 2.69435e-05, 2.110098e-05, 9.786656e-06,
  1.412738e-05, 3.444016e-05, 1.635069e-05, 2.225159e-05, 7.356462e-06, 
    8.719302e-07, 2.014427e-06, 3.486881e-06, 3.841482e-06, 2.111431e-06, 
    7.175692e-07, 9.108653e-07, 5.561317e-07, 1.272681e-07, 2.690871e-07,
  3.631439e-05, 3.37885e-05, 2.48995e-05, 1.747194e-05, 6.427564e-06, 
    2.510525e-07, 2.213334e-06, 3.22136e-06, 4.88044e-06, 3.200353e-06, 
    1.247699e-06, 2.836145e-06, 3.682734e-06, 3.42205e-08, 2.658369e-07,
  3.351846e-05, 2.381559e-05, 1.586314e-05, 1.812548e-05, 1.985387e-05, 
    7.334171e-07, 4.118428e-06, 7.266663e-06, 8.08518e-06, 7.848668e-06, 
    3.929903e-06, 3.392017e-06, 5.330818e-06, 3.87821e-06, 8.943454e-07,
  2.953811e-05, 1.496253e-05, 1.609937e-05, 1.831245e-05, 1.645817e-05, 
    5.183783e-06, 4.002048e-06, 5.362692e-06, 9.015164e-06, 9.118558e-06, 
    5.044044e-06, 4.002778e-06, 4.895315e-06, 5.037329e-06, 3.294717e-06,
  2.186925e-05, 1.425226e-05, 1.705011e-05, 1.835076e-05, 1.859686e-05, 
    2.50432e-05, 5.595197e-06, 2.7204e-06, 9.917804e-06, 3.8406e-06, 
    4.141937e-06, 4.583349e-06, 4.039588e-06, 3.886976e-06, 4.157724e-06,
  1.979912e-05, 1.518336e-05, 1.828795e-05, 1.711965e-05, 1.453967e-05, 
    2.846233e-05, 3.653477e-05, 1.00077e-05, 6.513677e-06, 1.137004e-05, 
    5.253334e-06, 4.09401e-06, 5.057036e-06, 3.682434e-06, 3.60486e-06,
  1.880611e-05, 1.776303e-05, 2.077824e-05, 1.521339e-05, 1.3767e-05, 
    2.771851e-05, 5.454841e-05, 3.307261e-05, 1.870485e-05, 1.397699e-05, 
    8.859436e-06, 5.220707e-06, 5.089776e-06, 4.91151e-06, 3.609422e-06,
  1.919027e-05, 2.068648e-05, 2.025739e-05, 1.960491e-05, 2.162403e-05, 
    3.15303e-05, 4.929882e-05, 3.467216e-05, 3.201815e-05, 2.176693e-05, 
    1.196053e-05, 5.668135e-06, 4.68384e-06, 5.203618e-06, 3.816795e-06,
  2.018142e-05, 2.152686e-05, 2.57855e-05, 2.41367e-05, 3.20894e-05, 
    3.495532e-05, 5.013483e-05, 3.623669e-05, 3.930576e-05, 1.867432e-05, 
    1.438282e-05, 6.87781e-06, 5.442775e-06, 5.600813e-06, 2.671478e-06,
  2.019565e-05, 2.283523e-05, 2.839691e-05, 3.400622e-05, 3.5409e-05, 
    3.545139e-05, 4.125768e-05, 3.571088e-05, 3.149284e-05, 2.456321e-05, 
    1.221603e-05, 7.44139e-06, 7.482104e-06, 5.503097e-06, 5.564933e-06,
  1.752341e-05, 2.099896e-05, 1.537613e-05, 2.173466e-05, 1.152757e-05, 
    4.971685e-06, 8.514819e-06, 3.574243e-06, 4.631477e-06, 2.614068e-06, 
    5.756787e-09, 1.016617e-06, 1.46572e-07, 7.788366e-08, 4.55008e-07,
  3.061757e-05, 2.768067e-05, 3.024626e-05, 3.695185e-05, 8.30832e-06, 
    5.380177e-06, 3.86527e-06, 3.439745e-06, 3.274955e-06, 3.304777e-06, 
    1.389057e-06, 2.84804e-06, 3.301066e-06, 4.41918e-07, 4.752208e-07,
  3.105542e-05, 2.622523e-05, 3.109545e-05, 4.069283e-05, 8.007421e-06, 
    6.22273e-06, 4.159048e-06, 5.101505e-06, 5.051807e-06, 4.263374e-06, 
    3.349738e-06, 2.779153e-06, 3.054392e-06, 2.109542e-06, 8.564373e-07,
  3.300374e-05, 2.806824e-05, 3.036661e-05, 3.879301e-05, 1.479754e-05, 
    7.166243e-07, 2.507696e-06, 5.116882e-06, 5.82435e-06, 4.166865e-06, 
    4.020592e-06, 2.532243e-06, 2.008002e-06, 1.417135e-06, 1.42629e-06,
  2.952376e-05, 3.114973e-05, 2.870732e-05, 4.113417e-05, 3.194893e-05, 
    6.580437e-06, 3.053424e-06, 1.463493e-07, 4.589897e-07, 2.77236e-07, 
    2.504381e-06, 2.519391e-06, 1.699709e-06, 1.717649e-06, 8.326155e-07,
  3.040198e-05, 3.231596e-05, 2.802285e-05, 3.641824e-05, 3.444136e-05, 
    2.795694e-05, 1.914651e-05, 2.357668e-06, 1.994413e-06, 7.307915e-06, 
    2.920713e-06, 2.248071e-06, 1.920849e-06, 1.234466e-06, 6.787951e-07,
  3.705618e-05, 3.34023e-05, 2.648386e-05, 3.159286e-05, 2.955497e-05, 
    3.914058e-05, 4.522553e-05, 2.220027e-05, 1.431991e-05, 1.110772e-05, 
    7.127015e-06, 2.768784e-06, 1.492566e-06, 1.24927e-06, 1.350831e-06,
  4.43046e-05, 3.436562e-05, 2.547515e-05, 2.70438e-05, 2.904631e-05, 
    3.622569e-05, 5.217173e-05, 3.874659e-05, 2.584917e-05, 2.092771e-05, 
    7.549831e-06, 2.63617e-06, 1.563876e-06, 1.645815e-06, 1.122549e-06,
  4.909705e-05, 3.40258e-05, 2.259159e-05, 2.231401e-05, 3.134281e-05, 
    3.785728e-05, 4.238695e-05, 3.91304e-05, 3.061182e-05, 2.232408e-05, 
    8.190901e-06, 2.533904e-06, 1.856204e-06, 2.396991e-06, 3.132101e-06,
  3.687808e-05, 1.86409e-05, 1.733961e-05, 2.4629e-05, 3.290036e-05, 
    3.397434e-05, 4.087497e-05, 3.626336e-05, 3.247584e-05, 1.804245e-05, 
    6.740474e-06, 2.608029e-06, 2.544454e-06, 3.917464e-06, 6.270015e-06,
  1.06478e-05, 1.431573e-05, 1.048107e-05, 1.287163e-05, 8.986055e-06, 
    3.892292e-06, 5.378562e-06, 5.099647e-06, 3.920752e-06, 1.090905e-06, 
    3.419457e-08, 4.124352e-07, 7.587582e-07, 6.906409e-07, 8.059101e-07,
  2.322648e-05, 2.387119e-05, 2.105791e-05, 2.240594e-05, 7.293786e-06, 
    4.666224e-06, 1.010588e-05, 5.663745e-06, 2.341855e-06, 1.705447e-06, 
    1.930042e-07, 1.168953e-06, 2.023119e-06, 8.371455e-07, 9.026458e-07,
  2.722425e-05, 2.825668e-05, 2.752863e-05, 3.183777e-05, 1.555354e-05, 
    4.297801e-06, 6.535015e-06, 4.288318e-06, 2.284601e-06, 1.688399e-06, 
    1.023505e-06, 9.42911e-07, 2.250051e-06, 2.393114e-06, 1.134731e-06,
  2.423591e-05, 2.654565e-05, 2.616609e-05, 3.669896e-05, 3.767787e-05, 
    6.328013e-06, 4.746244e-07, 2.228652e-06, 2.463529e-06, 1.141557e-06, 
    7.768962e-07, 4.356372e-07, 1.210966e-06, 1.795753e-06, 1.612568e-06,
  2.541812e-05, 2.563124e-05, 2.424826e-05, 3.129381e-05, 5.206249e-05, 
    2.070494e-05, 4.979934e-06, 3.150046e-07, 9.220792e-08, 2.429744e-08, 
    4.534852e-07, 2.158743e-07, 2.189301e-07, 1.826514e-06, 1.97209e-06,
  2.623544e-05, 2.377849e-05, 2.629076e-05, 3.276596e-05, 5.077579e-05, 
    3.031946e-05, 1.871367e-05, 4.494448e-06, 8.86356e-07, 2.825796e-06, 
    6.070585e-07, 2.16035e-07, 1.053637e-06, 2.217998e-06, 2.640924e-06,
  2.611388e-05, 2.659559e-05, 2.698322e-05, 3.540641e-05, 4.149429e-05, 
    3.658383e-05, 2.976739e-05, 2.127413e-05, 6.560479e-06, 7.505824e-06, 
    3.391236e-06, 4.457638e-07, 1.212298e-06, 2.147879e-06, 3.505626e-06,
  2.536511e-05, 2.712699e-05, 2.609855e-05, 3.842176e-05, 4.020065e-05, 
    3.068848e-05, 3.327176e-05, 3.605329e-05, 1.481386e-05, 1.677567e-05, 
    4.358502e-06, 6.029626e-07, 8.503265e-07, 3.121112e-06, 4.146217e-06,
  2.986007e-05, 2.917002e-05, 2.750625e-05, 4.146071e-05, 3.331664e-05, 
    2.649478e-05, 3.601538e-05, 3.18672e-05, 2.210747e-05, 2.143873e-05, 
    4.501671e-06, 6.521493e-07, 1.623643e-06, 3.246793e-06, 5.409243e-06,
  2.728973e-05, 2.489198e-05, 2.680654e-05, 3.519013e-05, 2.789481e-05, 
    2.304223e-05, 3.286481e-05, 3.442131e-05, 3.024768e-05, 1.269489e-05, 
    3.570869e-06, 9.656679e-07, 1.508252e-06, 2.905624e-06, 7.819478e-06,
  4.998793e-06, 7.65902e-06, 3.412169e-06, 5.245841e-06, 1.887118e-06, 
    3.041168e-06, 2.700231e-06, 1.53128e-06, 2.201577e-06, 1.532195e-06, 
    2.772602e-06, 2.358015e-06, 1.968987e-06, 1.393593e-06, 1.307008e-06,
  1.048298e-05, 1.494318e-05, 8.433472e-06, 1.12313e-05, 3.928435e-06, 
    2.583957e-06, 3.48558e-06, 1.506647e-06, 1.299753e-06, 1.85045e-06, 
    1.890599e-06, 3.966035e-06, 2.525848e-06, 1.577959e-06, 1.676463e-06,
  1.574986e-05, 1.802609e-05, 1.966399e-05, 1.5598e-05, 7.55392e-06, 
    2.757856e-06, 2.666781e-06, 1.407077e-06, 1.142679e-06, 2.308755e-06, 
    3.943802e-06, 5.13705e-06, 4.847727e-06, 3.3568e-06, 2.285886e-06,
  2.000883e-05, 2.696049e-05, 2.660057e-05, 2.720395e-05, 1.49541e-05, 
    7.735958e-06, 1.541842e-06, 6.129939e-08, 2.055062e-07, 1.060487e-06, 
    3.512821e-06, 3.0753e-06, 4.193606e-06, 3.231095e-06, 2.976665e-06,
  3.209926e-05, 3.366826e-05, 3.286461e-05, 3.452356e-05, 2.742427e-05, 
    1.319695e-05, 8.371133e-06, 2.66236e-06, 1.021162e-07, 8.98469e-07, 
    2.482654e-06, 3.033358e-06, 2.114281e-06, 4.35885e-06, 2.454068e-06,
  4.051539e-05, 3.744676e-05, 3.468842e-05, 3.213275e-05, 2.28083e-05, 
    2.252959e-05, 1.985927e-05, 3.177517e-06, 3.540291e-07, 1.222648e-06, 
    1.473193e-06, 2.277684e-06, 5.624359e-06, 5.522311e-06, 3.157246e-06,
  4.382286e-05, 4.7232e-05, 4.083032e-05, 3.308685e-05, 2.111509e-05, 
    2.485146e-05, 2.244575e-05, 1.488162e-05, 4.853005e-06, 2.868445e-06, 
    3.056387e-06, 2.302619e-06, 5.624697e-06, 5.441173e-06, 4.637694e-06,
  4.151858e-05, 4.808913e-05, 4.182328e-05, 3.613642e-05, 2.255305e-05, 
    2.105529e-05, 2.2509e-05, 1.880564e-05, 1.032971e-05, 9.882336e-06, 
    2.043281e-06, 1.114972e-06, 4.888148e-06, 6.157805e-06, 4.842219e-06,
  3.775155e-05, 4.475031e-05, 4.698021e-05, 3.4487e-05, 2.676021e-05, 
    1.937849e-05, 2.003453e-05, 1.896481e-05, 1.745352e-05, 9.744554e-06, 
    9.523638e-07, 5.158356e-07, 3.645368e-06, 6.140134e-06, 7.993112e-06,
  3.182033e-05, 3.316294e-05, 3.472876e-05, 3.111656e-05, 2.43347e-05, 
    1.740456e-05, 1.843311e-05, 2.499783e-05, 1.114864e-05, 1.293708e-06, 
    1.353442e-06, 2.360391e-07, 2.384027e-06, 5.382725e-06, 6.969449e-06,
  2.201507e-05, 1.809655e-05, 6.276631e-06, 4.392483e-06, 1.773554e-06, 
    3.522572e-07, 2.985092e-06, 3.576798e-06, 3.250454e-06, 1.637118e-06, 
    6.088225e-07, 5.360899e-07, 3.553882e-07, 3.413656e-07, 3.519811e-07,
  3.060243e-05, 2.574447e-05, 8.256703e-06, 7.890771e-06, 4.376517e-07, 
    2.342886e-07, 2.353646e-06, 3.394885e-06, 3.146197e-06, 3.260209e-06, 
    9.100903e-07, 6.487885e-07, 6.094171e-07, 2.671719e-07, 3.834202e-07,
  4.093137e-05, 3.442397e-05, 2.035385e-05, 1.302207e-05, 8.551165e-06, 
    1.589394e-06, 4.515638e-07, 2.731658e-06, 3.210897e-06, 3.269002e-06, 
    2.351889e-06, 9.835214e-07, 9.463446e-07, 8.064054e-07, 4.170828e-07,
  5.214785e-05, 5.47898e-05, 2.735289e-05, 1.727798e-05, 9.651163e-06, 
    5.410365e-06, 9.002266e-07, 1.128709e-06, 3.122523e-06, 3.695787e-06, 
    2.372291e-06, 2.122253e-06, 1.566494e-06, 1.36032e-06, 1.479317e-06,
  5.418365e-05, 5.748347e-05, 4.547316e-05, 3.379874e-05, 1.807458e-05, 
    1.40257e-05, 3.988113e-06, 1.506978e-06, 1.02718e-06, 2.171234e-06, 
    1.89155e-06, 2.688308e-06, 1.763245e-06, 1.491348e-06, 1.757153e-06,
  3.756225e-05, 4.828137e-05, 4.496732e-05, 2.878976e-05, 2.324308e-05, 
    1.919061e-05, 1.539657e-05, 3.142015e-06, 3.77586e-06, 6.24622e-06, 
    1.4737e-06, 3.344171e-06, 2.063058e-06, 1.89221e-06, 1.441565e-06,
  2.610262e-05, 3.746607e-05, 3.324546e-05, 2.733076e-05, 2.37115e-05, 
    1.929271e-05, 1.602088e-05, 1.237449e-05, 1.2518e-05, 1.268021e-05, 
    7.825873e-06, 4.13014e-06, 2.702758e-06, 2.788162e-06, 1.222801e-06,
  2.029222e-05, 2.43429e-05, 3.141717e-05, 2.648073e-05, 2.091228e-05, 
    1.893462e-05, 1.608677e-05, 1.236809e-05, 1.574148e-05, 1.338636e-05, 
    5.001908e-06, 4.503632e-06, 3.543877e-06, 3.268252e-06, 1.967328e-06,
  8.996947e-06, 2.023147e-05, 2.726487e-05, 2.325203e-05, 2.016671e-05, 
    2.030799e-05, 1.67495e-05, 1.475029e-05, 1.595659e-05, 1.249616e-05, 
    3.418822e-06, 4.661791e-06, 4.598432e-06, 4.292406e-06, 4.844431e-06,
  2.144176e-05, 1.019784e-05, 1.625401e-05, 2.199205e-05, 2.184052e-05, 
    1.500472e-05, 1.59726e-05, 1.647582e-05, 1.311972e-05, 6.501938e-06, 
    4.372801e-06, 4.185934e-06, 5.550366e-06, 5.267158e-06, 6.328429e-06,
  1.552007e-05, 3.279196e-05, 1.370485e-05, 8.230774e-06, 2.403046e-06, 
    8.947109e-07, 1.663719e-06, 8.984823e-07, 1.229593e-06, 1.472535e-07, 
    3.174239e-07, 2.630269e-07, 5.619775e-07, 2.567926e-07, 7.792533e-07,
  2.421359e-05, 3.86815e-05, 2.454916e-05, 1.695308e-05, 1.341209e-06, 
    1.254033e-06, 2.704043e-06, 1.537179e-06, 7.978408e-07, 4.93708e-07, 
    1.059226e-07, 2.118677e-07, 6.316327e-07, 3.901215e-07, 1.216401e-06,
  2.741767e-05, 4.107391e-05, 3.547553e-05, 2.119417e-05, 8.721006e-06, 
    1.180394e-06, 2.486973e-06, 1.630487e-06, 1.247308e-06, 8.813684e-07, 
    3.092141e-07, 4.067542e-07, 8.323493e-07, 2.190784e-06, 7.534626e-07,
  2.744207e-05, 4.211738e-05, 4.095511e-05, 2.377037e-05, 1.835674e-05, 
    5.369346e-06, 1.370283e-06, 3.709432e-07, 1.667814e-06, 6.972698e-07, 
    5.018362e-07, 2.880515e-07, 5.973994e-07, 1.463312e-06, 9.065301e-07,
  2.284937e-05, 3.670134e-05, 4.997773e-05, 4.136192e-05, 2.322079e-05, 
    1.769195e-05, 7.016017e-06, 2.258523e-06, 4.250411e-07, 4.471919e-08, 
    3.521147e-08, 2.757708e-07, 3.592066e-07, 7.00389e-07, 1.468963e-06,
  2.335516e-05, 3.570079e-05, 4.022707e-05, 3.551592e-05, 2.828414e-05, 
    2.462839e-05, 1.969481e-05, 4.573005e-06, 8.507042e-07, 1.222012e-06, 
    4.956352e-07, 7.572601e-07, 4.662857e-07, 6.920789e-07, 1.485584e-06,
  2.261596e-05, 3.085616e-05, 3.557306e-05, 2.797346e-05, 2.644337e-05, 
    2.269312e-05, 2.088257e-05, 1.707859e-05, 1.13213e-05, 4.805464e-06, 
    2.944914e-06, 7.601024e-07, 4.24443e-07, 8.518285e-07, 1.064457e-06,
  1.988127e-05, 2.709284e-05, 2.639515e-05, 2.546435e-05, 2.357973e-05, 
    2.106262e-05, 1.666488e-05, 1.682527e-05, 1.765642e-05, 1.282993e-05, 
    1.899801e-06, 1.1608e-06, 7.788253e-07, 5.764144e-07, 1.000481e-06,
  1.376657e-05, 2.070619e-05, 2.594516e-05, 1.944798e-05, 1.980348e-05, 
    1.977199e-05, 1.586107e-05, 1.47847e-05, 1.512546e-05, 1.247751e-05, 
    8.04066e-07, 1.315696e-06, 1.701364e-06, 1.089701e-06, 1.391836e-06,
  3.671504e-06, 1.172106e-05, 1.630736e-05, 1.800432e-05, 1.712807e-05, 
    1.66588e-05, 1.598885e-05, 1.19165e-05, 1.022398e-05, 1.910326e-06, 
    4.367544e-06, 3.755144e-06, 2.373468e-06, 2.344985e-06, 2.321552e-06,
  6.763263e-06, 1.193236e-05, 4.016117e-06, 5.889353e-06, 2.006802e-06, 
    1.824046e-07, 1.653464e-06, 1.690532e-06, 2.986036e-06, 1.192861e-06, 
    2.274012e-06, 2.820745e-06, 3.623316e-06, 2.152836e-06, 2.280014e-06,
  1.507645e-05, 1.987646e-05, 1.448813e-05, 1.055448e-05, 6.766785e-07, 
    3.750407e-08, 1.038627e-06, 1.217686e-06, 1.708718e-06, 1.056225e-06, 
    1.646769e-06, 1.809791e-06, 3.045232e-06, 3.113802e-06, 4.344904e-06,
  2.854803e-05, 2.438236e-05, 2.519524e-05, 1.568382e-05, 7.015562e-06, 
    7.744748e-07, 3.287183e-07, 6.237069e-07, 6.195275e-07, 8.705326e-07, 
    8.790709e-07, 1.731053e-06, 3.850345e-06, 8.319124e-06, 6.266853e-06,
  2.974493e-05, 2.911567e-05, 2.081978e-05, 2.096066e-05, 1.544463e-05, 
    5.639313e-06, 1.076971e-06, 5.464229e-08, 1.409378e-07, 4.800496e-07, 
    6.21204e-07, 1.140652e-06, 2.09036e-06, 3.95188e-06, 5.831717e-06,
  2.417445e-05, 2.594568e-05, 3.245455e-05, 2.746467e-05, 1.945025e-05, 
    1.164788e-05, 7.303208e-06, 1.635235e-06, 1.241921e-06, 4.352215e-07, 
    2.099072e-07, 7.629641e-07, 2.811809e-06, 3.222392e-06, 5.185057e-06,
  2.326039e-05, 2.246878e-05, 2.423201e-05, 2.413371e-05, 2.001474e-05, 
    1.708748e-05, 1.441458e-05, 7.062131e-06, 3.527574e-07, 5.240665e-08, 
    5.170422e-08, 4.927804e-07, 2.434387e-06, 3.86817e-06, 4.873932e-06,
  2.139024e-05, 2.055767e-05, 2.072162e-05, 1.950318e-05, 1.982272e-05, 
    1.549715e-05, 1.57318e-05, 1.518067e-05, 9.437919e-06, 4.229087e-06, 
    2.046076e-06, 1.040996e-06, 2.193831e-06, 3.765578e-06, 4.774584e-06,
  1.69181e-05, 1.869241e-05, 1.911675e-05, 2.028047e-05, 2.037645e-05, 
    1.756121e-05, 1.538677e-05, 1.662589e-05, 1.082312e-05, 7.717204e-06, 
    1.214045e-06, 7.056334e-07, 1.491254e-06, 3.159153e-06, 5.621006e-06,
  9.246479e-06, 1.707221e-05, 2.131385e-05, 1.804964e-05, 1.809993e-05, 
    1.867384e-05, 1.666229e-05, 1.303839e-05, 1.443538e-05, 6.680256e-06, 
    1.866727e-07, 1.458878e-06, 1.334596e-06, 2.027285e-06, 3.585908e-06,
  9.913512e-06, 1.039814e-05, 1.431267e-05, 1.641205e-05, 1.797968e-05, 
    1.775134e-05, 1.67597e-05, 1.452126e-05, 7.855944e-06, 3.512758e-07, 
    1.781435e-06, 9.459179e-07, 5.452825e-07, 8.063911e-07, 2.016058e-06,
  2.77858e-06, 9.419674e-06, 2.142617e-06, 2.541194e-06, 1.89134e-06, 
    1.493924e-07, 1.037957e-06, 1.316604e-06, 2.918207e-06, 3.523624e-06, 
    4.458025e-06, 4.154181e-06, 4.087705e-06, 2.058804e-06, 2.825804e-06,
  1.023586e-05, 1.42337e-05, 1.245857e-05, 8.123897e-06, 1.162887e-06, 
    7.344101e-07, 2.430932e-07, 8.809419e-07, 1.705374e-06, 2.201768e-06, 
    3.744961e-06, 3.802121e-06, 1.829889e-06, 1.834353e-06, 3.39151e-06,
  2.081403e-05, 1.777669e-05, 1.532809e-05, 1.088033e-05, 2.15391e-06, 
    1.316271e-06, 4.087682e-07, 9.756868e-07, 2.420961e-06, 2.750422e-06, 
    2.691783e-06, 2.678114e-06, 5.093994e-06, 7.743492e-06, 5.120096e-06,
  1.788367e-05, 1.616439e-05, 1.473468e-05, 1.127074e-05, 1.139116e-05, 
    3.990029e-06, 1.548335e-06, 6.877104e-07, 1.793219e-06, 2.044437e-06, 
    3.00058e-06, 3.223289e-06, 2.705224e-06, 6.07837e-06, 3.919945e-06,
  1.672238e-05, 1.412579e-05, 1.355057e-05, 1.13089e-05, 1.068416e-05, 
    1.32228e-05, 2.66206e-06, 1.851501e-06, 2.677953e-06, 2.751166e-06, 
    4.567738e-06, 4.180816e-06, 2.142131e-06, 1.130754e-06, 6.58646e-06,
  1.304478e-05, 1.41927e-05, 1.432241e-05, 1.290115e-05, 1.213267e-05, 
    1.227119e-05, 1.035767e-05, 6.177894e-06, 2.799416e-07, 2.981608e-06, 
    6.013041e-06, 4.284357e-06, 3.238332e-06, 2.675579e-06, 2.933871e-06,
  1.318736e-05, 1.355458e-05, 1.397682e-05, 1.39412e-05, 1.412605e-05, 
    1.340062e-05, 1.066852e-05, 6.673246e-06, 8.591696e-06, 7.852006e-06, 
    4.248632e-06, 7.661565e-06, 6.757009e-06, 4.037841e-06, 3.630639e-06,
  1.30427e-05, 1.397821e-05, 1.415083e-05, 1.51775e-05, 1.649977e-05, 
    1.531894e-05, 1.175805e-05, 8.198056e-06, 8.165056e-06, 8.254695e-06, 
    3.11807e-06, 7.598513e-06, 5.741099e-06, 5.305281e-06, 5.286512e-06,
  5.634334e-05, 6.461261e-05, 5.697446e-05, 3.629631e-05, 1.920628e-05, 
    1.465611e-05, 1.419324e-05, 1.307266e-05, 7.863641e-06, 8.484423e-06, 
    6.945814e-07, 4.438205e-06, 4.735038e-06, 4.875713e-06, 4.020088e-06,
  8.764693e-05, 9.081877e-05, 7.929967e-05, 5.120238e-05, 2.561474e-05, 
    1.086447e-05, 1.1126e-05, 1.095444e-05, 5.071305e-06, 8.579331e-07, 
    1.310499e-06, 5.619085e-06, 4.340158e-06, 3.291143e-06, 1.183014e-05,
  2.225269e-06, 2.892379e-06, 1.524403e-07, 2.587593e-07, 1.4203e-06, 
    4.082505e-07, 7.31055e-07, 1.978219e-06, 2.103851e-06, 3.176472e-06, 
    4.301305e-06, 5.661399e-06, 6.743454e-06, 6.832377e-06, 1.163252e-05,
  6.275816e-06, 1.153149e-05, 1.233574e-05, 9.573107e-06, 3.546137e-06, 
    1.007009e-06, 1.127512e-07, 7.43574e-07, 1.108131e-06, 1.508472e-06, 
    3.397086e-06, 4.136726e-06, 5.733872e-06, 5.125845e-06, 1.056169e-05,
  1.398998e-05, 1.686552e-05, 1.240102e-05, 1.395197e-05, 5.842602e-06, 
    3.481336e-06, 1.837889e-07, 8.079307e-07, 1.254941e-06, 1.008941e-06, 
    1.18998e-06, 2.280234e-06, 6.541944e-06, 1.13755e-05, 9.984505e-06,
  1.642843e-05, 1.560874e-05, 1.395927e-05, 1.774874e-05, 1.723473e-05, 
    4.412449e-06, 1.570061e-06, 4.230978e-07, 4.742667e-07, 6.092508e-07, 
    1.160475e-06, 1.199646e-06, 2.543686e-06, 9.145764e-06, 5.537893e-06,
  1.343384e-05, 1.610334e-05, 2.10746e-05, 1.955415e-05, 1.785224e-05, 
    8.190154e-06, 2.515264e-06, 1.601185e-06, 2.78612e-06, 4.826368e-07, 
    7.500761e-07, 4.484262e-07, 7.928239e-07, 1.734219e-06, 7.445217e-06,
  6.418928e-06, 1.359723e-05, 2.084397e-05, 2.069545e-05, 2.023797e-05, 
    1.348001e-05, 5.161909e-06, 1.313146e-06, 9.728076e-08, 1.206034e-06, 
    2.032461e-06, 1.084246e-07, 3.531841e-07, 8.079149e-07, 5.904346e-06,
  2.030655e-05, 1.592009e-05, 1.266675e-05, 1.38811e-05, 1.582172e-05, 
    1.279312e-05, 9.994381e-06, 1.198962e-05, 4.209625e-06, 6.300318e-06, 
    2.737486e-08, 3.153783e-08, 1.358806e-07, 2.956658e-07, 7.475192e-07,
  4.62646e-05, 4.615689e-05, 4.006907e-05, 2.395116e-05, 1.465185e-05, 
    1.483932e-05, 9.728508e-06, 5.051705e-06, 9.058657e-06, 5.880824e-06, 
    7.000906e-09, 2.054156e-08, 5.71902e-08, 9.548418e-08, 1.915701e-07,
  2.893395e-05, 4.288947e-05, 4.876393e-05, 2.644561e-05, 2.074928e-05, 
    1.257386e-05, 7.321855e-06, 9.229324e-06, 9.628874e-06, 1.031796e-05, 
    1.032004e-07, 9.538481e-09, 3.657588e-08, 1.171627e-07, 9.138574e-07,
  3.507137e-06, 6.316194e-06, 8.916379e-06, 1.373738e-05, 1.765994e-05, 
    9.046523e-06, 5.955465e-06, 9.681086e-06, 8.563119e-06, 7.126378e-07, 
    4.589815e-07, 2.777547e-08, 1.406318e-08, 1.534899e-07, 3.418753e-06,
  2.361968e-06, 3.679297e-06, 2.085587e-06, 3.434955e-06, 1.410155e-06, 
    1.70226e-06, 3.074804e-06, 1.657314e-06, 3.391615e-07, 1.906705e-06, 
    3.151204e-06, 4.471759e-06, 6.487726e-06, 7.042913e-06, 1.132477e-05,
  5.276638e-06, 9.756613e-06, 1.247526e-05, 1.653389e-05, 4.717509e-06, 
    2.333068e-06, 1.183522e-06, 2.662659e-06, 2.372444e-07, 2.39283e-07, 
    1.819876e-06, 2.833425e-06, 3.935127e-06, 6.545625e-06, 9.150286e-06,
  1.39207e-05, 1.50208e-05, 1.410074e-05, 2.709829e-05, 1.042501e-05, 
    5.898223e-06, 1.091277e-06, 5.368198e-07, 2.822784e-08, 4.807691e-08, 
    2.407708e-07, 1.355583e-06, 7.46391e-06, 8.867955e-06, 1.162883e-05,
  2.274672e-05, 1.789954e-05, 1.490572e-05, 1.252749e-05, 1.834064e-05, 
    3.37133e-06, 4.493654e-06, 9.762273e-08, 2.547351e-08, 2.409576e-08, 
    4.38705e-07, 6.636859e-07, 6.102874e-06, 1.285677e-05, 9.443009e-06,
  2.284157e-05, 2.201252e-05, 1.832084e-05, 1.23559e-05, 1.784549e-05, 
    1.392559e-05, 3.124778e-06, 2.783818e-06, 1.426091e-06, 6.602233e-07, 
    1.407351e-06, 1.405652e-07, 6.726287e-07, 3.153521e-06, 8.483963e-06,
  1.815807e-05, 1.964586e-05, 2.132296e-05, 1.423461e-05, 1.491237e-05, 
    1.445729e-05, 9.55023e-06, 9.831979e-07, 1.648672e-06, 7.1541e-08, 
    9.583993e-07, 2.696834e-07, 3.577169e-07, 8.888104e-07, 5.442631e-06,
  1.40147e-05, 1.849571e-05, 1.84875e-05, 1.516381e-05, 1.237466e-05, 
    9.604869e-06, 1.064506e-05, 1.108241e-05, 4.955933e-06, 1.563534e-06, 
    1.997664e-07, 5.593478e-07, 7.249608e-07, 2.865512e-07, 1.055049e-06,
  1.777885e-05, 2.076536e-05, 1.941081e-05, 1.364058e-05, 1.273982e-05, 
    9.239765e-06, 1.195238e-05, 1.058354e-05, 7.609872e-06, 6.026878e-06, 
    2.968357e-06, 1.642873e-06, 1.740739e-06, 5.166535e-07, 6.40182e-07,
  2.041461e-05, 2.299178e-05, 1.754985e-05, 1.447968e-05, 9.408461e-06, 
    9.41249e-06, 8.721047e-06, 8.900474e-06, 8.728232e-06, 4.757491e-06, 
    2.414378e-06, 2.254914e-06, 1.993671e-06, 1.325261e-06, 2.110409e-06,
  1.013169e-05, 1.205676e-05, 1.29036e-05, 1.10453e-05, 7.653897e-06, 
    4.354697e-06, 4.902782e-06, 4.732983e-06, 5.208041e-07, 9.67793e-08, 
    1.361636e-06, 1.846944e-06, 1.388528e-06, 1.041733e-06, 8.092092e-07,
  1.679785e-05, 1.295379e-05, 4.541805e-06, 2.673489e-06, 3.623758e-06, 
    3.10659e-06, 3.240261e-06, 2.89048e-06, 1.864396e-07, 1.887635e-06, 
    2.698043e-06, 1.879677e-06, 3.736282e-06, 4.596312e-06, 8.190429e-06,
  1.778411e-05, 1.503239e-05, 9.274941e-06, 9.292849e-06, 1.732097e-06, 
    2.774492e-06, 2.820868e-06, 2.870109e-06, 5.473509e-07, 3.807248e-07, 
    1.508642e-06, 1.584461e-06, 2.310973e-06, 5.929754e-06, 8.255264e-06,
  2.834806e-05, 2.55667e-05, 2.716348e-05, 1.71766e-05, 6.664808e-06, 
    1.691246e-06, 3.884079e-07, 3.474756e-06, 5.310843e-07, 5.584491e-07, 
    7.826204e-07, 1.856303e-06, 3.733137e-06, 7.965262e-06, 1.032341e-05,
  3.623783e-05, 3.662251e-05, 3.352518e-05, 2.847776e-05, 1.51221e-05, 
    3.517984e-06, 3.094873e-06, 7.119495e-07, 2.181694e-07, 3.51844e-07, 
    3.508667e-07, 2.338775e-06, 4.633009e-06, 8.765182e-06, 9.793521e-06,
  4.321398e-05, 3.531141e-05, 2.605879e-05, 1.969615e-05, 1.853898e-05, 
    1.429836e-05, 5.719566e-06, 9.184429e-06, 7.521792e-06, 1.453436e-06, 
    8.814479e-07, 3.578764e-06, 6.279165e-06, 9.542036e-06, 1.164057e-05,
  4.115492e-05, 3.426007e-05, 2.410801e-05, 1.625662e-05, 1.280413e-05, 
    1.002139e-05, 9.484224e-06, 6.920191e-06, 2.248738e-06, 3.626084e-06, 
    3.923686e-06, 5.483984e-06, 8.837703e-06, 1.00932e-05, 1.176014e-05,
  3.794126e-05, 3.155717e-05, 2.443832e-05, 1.784052e-05, 1.34026e-05, 
    1.019956e-05, 1.010665e-05, 7.963862e-06, 2.957097e-06, 3.776676e-06, 
    5.659197e-06, 6.578452e-06, 9.363164e-06, 9.934309e-06, 1.176835e-05,
  2.879559e-05, 2.663204e-05, 2.356624e-05, 1.919951e-05, 1.440352e-05, 
    1.111596e-05, 9.514882e-06, 9.452988e-06, 6.545205e-06, 1.674366e-06, 
    2.841098e-06, 3.948043e-06, 5.329572e-06, 1.005735e-05, 1.258036e-05,
  2.08936e-05, 2.035832e-05, 2.101844e-05, 1.667817e-05, 1.388909e-05, 
    1.172051e-05, 9.25818e-06, 7.254724e-06, 6.270389e-06, 5.410525e-07, 
    3.376672e-07, 6.817547e-07, 2.54626e-06, 7.395258e-06, 1.251245e-05,
  1.259752e-05, 1.474983e-05, 1.407852e-05, 1.204776e-05, 9.447641e-06, 
    7.271488e-06, 7.311155e-06, 4.853964e-06, 9.683804e-07, 4.104438e-07, 
    5.032321e-07, 2.907997e-06, 6.463425e-06, 7.351309e-06, 1.016837e-05,
  1.019132e-05, 1.429162e-05, 7.18898e-06, 4.190149e-06, 2.855155e-06, 
    4.730629e-07, 8.679834e-07, 6.944843e-07, 1.480787e-06, 1.767908e-06, 
    2.002815e-06, 3.654836e-06, 1.133303e-05, 2.055789e-05, 1.681869e-05,
  1.971646e-05, 2.52029e-05, 1.563731e-05, 8.502132e-06, 1.796802e-06, 
    5.143004e-07, 1.665328e-06, 1.715135e-06, 1.407405e-06, 1.799293e-06, 
    1.969346e-06, 3.838713e-06, 1.116106e-05, 2.34181e-05, 1.536804e-05,
  3.900062e-05, 3.768644e-05, 2.615728e-05, 1.564158e-05, 4.830132e-06, 
    1.119975e-06, 1.112553e-07, 1.926906e-06, 2.876144e-06, 9.439881e-07, 
    2.224371e-06, 5.046015e-06, 1.199461e-05, 2.207496e-05, 1.270153e-05,
  4.952309e-05, 4.725549e-05, 3.580248e-05, 2.157031e-05, 5.419633e-06, 
    3.06757e-06, 1.818912e-06, 2.172987e-06, 2.039958e-06, 2.059983e-06, 
    4.639509e-06, 6.24634e-06, 1.203247e-05, 2.29471e-05, 1.076451e-05,
  5.44633e-05, 5.451138e-05, 4.606473e-05, 2.828587e-05, 1.716509e-05, 
    5.091977e-06, 2.341503e-06, 2.144214e-06, 5.867833e-06, 6.944091e-06, 
    6.395433e-06, 7.277795e-06, 9.896517e-06, 1.829534e-05, 1.094894e-05,
  5.131691e-05, 5.078133e-05, 4.452249e-05, 3.326208e-05, 1.73707e-05, 
    1.08669e-05, 7.237678e-06, 1.171141e-06, 3.042656e-06, 5.521682e-06, 
    5.905438e-06, 6.807515e-06, 8.688965e-06, 1.405308e-05, 1.410963e-05,
  5.229908e-05, 4.786335e-05, 3.821086e-05, 2.862693e-05, 2.051821e-05, 
    1.156676e-05, 1.186177e-05, 1.050138e-05, 5.680392e-06, 2.581159e-06, 
    2.876499e-06, 4.14987e-06, 6.37824e-06, 1.211233e-05, 1.56442e-05,
  4.63158e-05, 4.14145e-05, 3.598603e-05, 2.839445e-05, 2.295552e-05, 
    1.682359e-05, 1.218047e-05, 9.986374e-06, 8.661502e-06, 8.260026e-07, 
    7.839676e-07, 1.221917e-06, 4.202304e-06, 9.894963e-06, 1.623417e-05,
  3.763423e-05, 3.663676e-05, 3.184832e-05, 2.337728e-05, 1.812362e-05, 
    1.500236e-05, 1.120729e-05, 1.089025e-05, 9.619418e-06, 4.656197e-07, 
    5.644252e-07, 1.814748e-06, 6.220171e-06, 8.070889e-06, 1.331984e-05,
  2.805151e-05, 2.205809e-05, 1.853048e-05, 1.738057e-05, 1.329053e-05, 
    1.064093e-05, 1.022843e-05, 9.525797e-06, 2.149165e-06, 1.910092e-07, 
    9.586181e-07, 2.941222e-06, 4.891826e-06, 5.536183e-06, 9.570052e-06,
  2.420271e-06, 1.002945e-06, 3.389465e-07, 3.312222e-07, 7.199221e-07, 
    8.650488e-08, 2.890324e-07, 7.456234e-07, 1.693031e-06, 3.693009e-06, 
    4.518564e-06, 5.597477e-06, 5.721421e-06, 6.457637e-06, 8.82586e-06,
  7.509135e-06, 4.081869e-06, 5.199538e-06, 1.41148e-06, 3.083072e-07, 
    3.392402e-07, 2.539348e-07, 4.442673e-07, 9.218161e-07, 4.043176e-06, 
    6.082799e-06, 7.19323e-06, 6.111098e-06, 7.830624e-06, 1.137367e-05,
  1.621273e-05, 1.184945e-05, 7.478134e-06, 7.02918e-06, 3.037742e-06, 
    8.3124e-07, 3.009641e-07, 4.297036e-07, 1.636061e-06, 4.318609e-06, 
    6.736758e-06, 7.384607e-06, 6.998866e-06, 8.246197e-06, 1.053737e-05,
  2.165582e-05, 1.82455e-05, 1.686122e-05, 1.536254e-05, 7.523749e-06, 
    3.138747e-06, 1.260253e-06, 4.536065e-07, 7.49977e-07, 4.742897e-06, 
    7.113646e-06, 7.291883e-06, 6.750661e-06, 8.621471e-06, 9.830972e-06,
  2.451051e-05, 2.061811e-05, 2.15798e-05, 2.262256e-05, 1.61751e-05, 
    5.451211e-06, 1.864828e-06, 1.197806e-06, 3.939598e-06, 5.73594e-06, 
    6.638948e-06, 6.588614e-06, 6.712099e-06, 6.80788e-06, 9.339647e-06,
  2.789911e-05, 2.295696e-05, 2.283804e-05, 2.638529e-05, 2.591391e-05, 
    1.805915e-05, 7.482464e-06, 4.628711e-07, 5.913032e-07, 5.342659e-06, 
    6.468746e-06, 6.387842e-06, 5.55564e-06, 5.919002e-06, 8.388273e-06,
  2.863616e-05, 2.966729e-05, 2.758128e-05, 2.681372e-05, 2.71814e-05, 
    1.930936e-05, 1.434495e-05, 6.86964e-06, 3.509128e-06, 2.515147e-06, 
    5.752485e-06, 5.646635e-06, 5.189911e-06, 6.28566e-06, 7.515919e-06,
  3.45758e-05, 3.548714e-05, 3.371477e-05, 3.386008e-05, 3.071837e-05, 
    2.488208e-05, 1.673439e-05, 1.553962e-05, 1.550162e-05, 7.05091e-07, 
    1.132615e-06, 2.256493e-06, 2.879923e-06, 4.371236e-06, 7.79269e-06,
  3.332357e-05, 3.648308e-05, 3.961209e-05, 3.514978e-05, 2.816588e-05, 
    2.512722e-05, 2.085533e-05, 1.700093e-05, 1.344615e-05, 2.012654e-06, 
    1.617111e-07, 5.43757e-08, 4.829727e-07, 2.202753e-06, 4.587263e-06,
  2.530439e-05, 2.734741e-05, 2.694391e-05, 2.673512e-05, 2.574527e-05, 
    2.346001e-05, 2.082595e-05, 1.399853e-05, 6.455556e-06, 7.681368e-07, 
    1.901549e-07, 9.609745e-08, 4.16773e-07, 1.674094e-06, 4.197016e-06,
  1.720687e-06, 9.915171e-07, 7.302187e-07, 1.368717e-07, 1.37194e-07, 
    4.226952e-07, 2.212581e-06, 2.699999e-06, 3.959523e-06, 6.292029e-06, 
    7.356979e-06, 9.507394e-06, 1.625483e-05, 1.749035e-05, 1.273559e-05,
  6.986319e-06, 5.907416e-06, 6.189685e-06, 1.186788e-06, 6.586768e-08, 
    2.119105e-07, 2.066933e-07, 1.711378e-06, 1.700322e-06, 4.155101e-06, 
    6.379914e-06, 8.464649e-06, 1.258742e-05, 1.692286e-05, 1.298179e-05,
  1.520141e-05, 1.251777e-05, 9.096638e-06, 5.997574e-06, 3.8975e-06, 
    5.474674e-07, 3.487833e-07, 7.440032e-07, 1.496901e-06, 3.16432e-06, 
    4.747621e-06, 6.217695e-06, 1.223832e-05, 1.62746e-05, 1.427351e-05,
  2.38569e-05, 1.70512e-05, 1.616338e-05, 1.313991e-05, 9.923037e-06, 
    2.743128e-06, 2.994015e-06, 8.409573e-07, 3.322271e-07, 2.384102e-06, 
    3.81233e-06, 6.099342e-06, 1.22123e-05, 1.685415e-05, 1.487616e-05,
  2.950269e-05, 1.479674e-05, 1.403407e-05, 1.651181e-05, 1.785694e-05, 
    1.633741e-05, 5.356012e-06, 5.610401e-06, 1.099156e-06, 1.27361e-06, 
    3.051626e-06, 4.131256e-06, 9.338899e-06, 1.328868e-05, 1.400152e-05,
  2.929006e-05, 2.280487e-05, 2.264352e-05, 2.235397e-05, 2.097896e-05, 
    2.103296e-05, 1.97846e-05, 4.556274e-06, 1.573348e-06, 1.756465e-06, 
    2.055083e-06, 2.385766e-06, 6.028403e-06, 1.243947e-05, 1.431996e-05,
  2.740443e-05, 2.41747e-05, 2.159867e-05, 1.93778e-05, 2.017259e-05, 
    2.126551e-05, 2.263021e-05, 1.524948e-05, 6.542926e-06, 1.949131e-06, 
    1.134831e-06, 1.406908e-06, 3.701305e-06, 1.018199e-05, 1.444127e-05,
  2.743059e-05, 2.302405e-05, 1.950187e-05, 1.988472e-05, 1.851487e-05, 
    1.947337e-05, 1.951334e-05, 1.909185e-05, 1.20168e-05, 2.09389e-06, 
    1.516444e-06, 8.128459e-07, 1.479639e-06, 5.251607e-06, 1.206442e-05,
  2.249177e-05, 2.378021e-05, 2.566028e-05, 2.152541e-05, 1.883411e-05, 
    2.024529e-05, 1.542031e-05, 1.567495e-05, 1.358881e-05, 1.617355e-06, 
    1.13481e-06, 6.243171e-07, 2.510206e-07, 1.657021e-06, 1.122954e-05,
  1.906133e-05, 2.056616e-05, 2.510234e-05, 2.899638e-05, 2.612138e-05, 
    2.378261e-05, 2.301912e-05, 1.739239e-05, 8.930825e-06, 2.990115e-06, 
    2.28923e-06, 8.021394e-07, 2.844052e-07, 2.370533e-07, 7.402016e-06,
  4.38411e-07, 1.67716e-06, 1.665448e-06, 6.461823e-08, 5.82079e-07, 
    6.220338e-07, 9.366979e-07, 1.790739e-06, 1.424283e-06, 1.074343e-06, 
    2.523721e-06, 4.573515e-06, 8.630541e-07, 3.085891e-08, 8.929901e-08,
  7.017721e-06, 1.245286e-05, 9.157158e-06, 1.675363e-06, 1.67544e-07, 
    6.254828e-07, 9.128062e-07, 2.56023e-06, 2.031304e-06, 9.497741e-07, 
    2.631765e-06, 4.530889e-06, 8.548363e-07, 3.588297e-08, 4.757691e-08,
  1.452641e-05, 1.777485e-05, 1.71487e-05, 9.84588e-06, 3.361682e-06, 
    2.107524e-06, 9.163303e-07, 6.84764e-06, 7.822085e-06, 1.084105e-06, 
    1.35635e-06, 3.609963e-06, 8.114611e-07, 9.630833e-07, 1.55404e-07,
  1.802359e-05, 1.767656e-05, 1.507476e-05, 1.465118e-05, 1.751153e-05, 
    8.239923e-06, 2.518504e-06, 7.945687e-06, 9.045046e-06, 4.970079e-06, 
    8.788862e-07, 2.057881e-06, 1.183631e-06, 8.978193e-07, 7.437217e-07,
  2.136916e-05, 1.591574e-05, 1.554368e-05, 1.485878e-05, 1.70911e-05, 
    1.637649e-05, 2.073669e-05, 9.295667e-06, 1.24919e-05, 7.357884e-06, 
    1.060381e-06, 1.413313e-06, 1.412179e-06, 4.965866e-07, 6.253246e-07,
  2.011425e-05, 1.526475e-05, 1.547843e-05, 1.561834e-05, 1.669218e-05, 
    2.338361e-05, 1.689074e-05, 9.387047e-06, 3.330074e-06, 5.865343e-06, 
    1.365608e-06, 8.407962e-07, 2.404515e-06, 4.227545e-07, 3.996568e-07,
  1.980259e-05, 2.156249e-05, 1.862725e-05, 1.628166e-05, 2.117784e-05, 
    2.544279e-05, 2.599592e-05, 1.802276e-05, 1.039455e-05, 2.476559e-06, 
    1.882746e-06, 6.88501e-07, 3.806047e-06, 8.385411e-07, 4.332983e-07,
  1.996472e-05, 2.112027e-05, 1.990349e-05, 2.038105e-05, 2.351382e-05, 
    2.248088e-05, 1.58135e-05, 1.227577e-05, 7.205235e-06, 1.336139e-06, 
    2.985456e-06, 1.00515e-06, 1.650165e-06, 2.606996e-06, 2.200362e-07,
  2.434849e-05, 2.746887e-05, 2.59307e-05, 2.391366e-05, 2.127541e-05, 
    1.754971e-05, 1.049784e-05, 1.011976e-05, 9.440493e-06, 9.332725e-07, 
    1.471202e-06, 6.200959e-07, 4.963056e-07, 4.782186e-06, 1.702597e-06,
  2.321937e-05, 2.001971e-05, 1.694103e-05, 1.445459e-05, 1.010794e-05, 
    7.040107e-06, 8.518131e-06, 1.448038e-05, 5.035609e-06, 3.301286e-06, 
    1.926825e-06, 7.346143e-07, 3.52854e-07, 1.047857e-06, 3.945687e-06,
  1.516913e-06, 8.239923e-08, 2.581756e-10, 2.231725e-09, 2.844952e-07, 
    1.87156e-06, 1.706787e-05, 1.122739e-05, 1.751535e-06, 3.084805e-07, 
    8.003174e-08, 2.520468e-08, 3.045683e-07, 3.413798e-07, 1.390794e-06,
  1.147556e-05, 8.338392e-06, 1.349617e-06, 3.970079e-08, 2.929791e-07, 
    4.31442e-07, 1.133363e-05, 1.252288e-05, 2.075102e-06, 1.306427e-06, 
    3.425369e-07, 5.211479e-07, 2.116771e-07, 6.600342e-07, 1.779291e-06,
  1.957787e-05, 1.13514e-05, 7.043172e-06, 5.108544e-06, 2.202856e-07, 
    1.885953e-06, 4.600724e-06, 1.412171e-05, 9.645621e-06, 2.21012e-06, 
    1.369624e-06, 3.146798e-07, 1.567769e-07, 4.181463e-07, 1.590939e-06,
  1.986166e-05, 1.08413e-05, 9.169778e-06, 1.257795e-05, 1.539692e-05, 
    8.560031e-06, 9.810551e-06, 1.322464e-05, 1.193209e-05, 5.834429e-06, 
    1.52991e-06, 3.820314e-07, 1.179862e-07, 5.333941e-07, 1.130075e-06,
  2.096957e-05, 1.27376e-05, 1.05563e-05, 1.104291e-05, 2.223866e-05, 
    2.857326e-05, 1.900484e-05, 1.507734e-05, 1.128167e-05, 2.60068e-06, 
    7.352668e-07, 5.644448e-08, 6.762643e-08, 3.276992e-07, 1.296354e-06,
  2.309719e-05, 1.834346e-05, 1.597187e-05, 1.409378e-05, 2.445394e-05, 
    2.956753e-05, 2.225094e-05, 7.814523e-06, 9.260028e-07, 1.072765e-06, 
    1.456579e-06, 3.894836e-07, 5.505185e-08, 1.838108e-07, 1.266771e-06,
  2.176537e-05, 1.966818e-05, 1.64994e-05, 1.876371e-05, 2.343288e-05, 
    2.168384e-05, 1.614148e-05, 1.010603e-05, 2.700652e-06, 9.386067e-07, 
    2.299684e-06, 3.646672e-07, 2.784558e-07, 2.251251e-07, 6.935503e-07,
  2.077392e-05, 2.124612e-05, 1.92902e-05, 1.886455e-05, 2.25543e-05, 
    1.753712e-05, 9.46561e-06, 8.829628e-06, 6.347862e-06, 4.441195e-06, 
    5.434812e-06, 2.078072e-06, 6.554079e-07, 6.47703e-07, 5.08523e-07,
  1.609646e-05, 2.016982e-05, 2.068162e-05, 1.765802e-05, 1.85114e-05, 
    1.251905e-05, 7.90888e-06, 6.676141e-06, 9.282283e-06, 6.08155e-06, 
    6.800586e-06, 4.955837e-06, 3.084803e-06, 2.531189e-06, 4.189246e-07,
  2.148743e-05, 1.927221e-05, 1.6584e-05, 1.356815e-05, 1.108919e-05, 
    6.819135e-06, 5.94451e-06, 9.537712e-06, 7.251434e-06, 6.818907e-06, 
    8.850903e-06, 8.929336e-06, 6.051358e-06, 3.252666e-06, 1.049695e-06,
  1.786156e-06, 7.566111e-07, 8.355103e-07, 9.464239e-07, 6.918989e-08, 
    2.448829e-06, 7.757296e-06, 2.240316e-06, 1.634962e-06, 3.870071e-06, 
    6.457278e-06, 8.822904e-06, 7.238436e-06, 5.333779e-06, 5.424189e-06,
  5.092377e-06, 3.45888e-06, 4.764355e-06, 3.207106e-07, 1.936408e-08, 
    6.954681e-07, 1.831928e-06, 8.46382e-07, 9.156275e-07, 2.757125e-06, 
    5.50525e-06, 8.863612e-06, 7.123725e-06, 5.463524e-06, 6.344337e-06,
  1.092712e-05, 1.075936e-05, 1.326279e-05, 1.489504e-05, 7.377046e-07, 
    1.975972e-06, 2.797502e-07, 1.467832e-06, 2.206071e-06, 4.136064e-06, 
    6.302214e-06, 7.975711e-06, 7.387626e-06, 6.120313e-06, 7.618251e-06,
  1.8346e-05, 2.217593e-05, 1.960682e-05, 1.82465e-05, 1.385918e-05, 
    2.671441e-06, 8.612859e-07, 1.786928e-06, 1.501696e-06, 2.601482e-06, 
    8.801257e-06, 8.18821e-06, 7.602389e-06, 5.929284e-06, 7.097375e-06,
  3.143772e-05, 2.657136e-05, 2.126952e-05, 1.702488e-05, 2.053999e-05, 
    2.113798e-05, 1.585999e-05, 8.574366e-06, 9.980178e-06, 3.61523e-06, 
    1.103004e-05, 9.8193e-06, 8.927305e-06, 4.426821e-06, 6.628848e-06,
  3.180317e-05, 2.816008e-05, 2.15683e-05, 1.654928e-05, 1.964123e-05, 
    2.334628e-05, 1.87631e-05, 4.802107e-06, 3.731929e-06, 7.688977e-06, 
    1.302225e-05, 1.148125e-05, 9.571459e-06, 3.779211e-06, 5.849648e-06,
  3.328741e-05, 2.738107e-05, 2.336301e-05, 2.185489e-05, 1.933665e-05, 
    1.666956e-05, 1.961949e-05, 1.368678e-05, 4.006573e-06, 5.541144e-06, 
    1.035405e-05, 1.16807e-05, 8.4745e-06, 3.445447e-06, 4.358356e-06,
  2.519741e-05, 2.835957e-05, 2.568187e-05, 2.343929e-05, 2.146817e-05, 
    1.819345e-05, 1.780016e-05, 1.740474e-05, 5.024447e-06, 5.1125e-06, 
    7.78751e-06, 9.21228e-06, 7.563617e-06, 3.722954e-06, 3.493279e-06,
  2.499749e-05, 2.863413e-05, 2.72618e-05, 2.058027e-05, 2.003493e-05, 
    1.895485e-05, 1.512995e-05, 9.581368e-06, 1.829679e-05, 6.448705e-06, 
    5.458979e-06, 6.154036e-06, 6.142579e-06, 4.730866e-06, 2.635524e-06,
  2.047012e-05, 2.031241e-05, 1.759104e-05, 1.396208e-05, 1.283725e-05, 
    6.678508e-06, 2.990557e-06, 1.032636e-05, 8.04331e-06, 7.877687e-06, 
    7.765108e-06, 5.838626e-06, 5.302623e-06, 6.694871e-06, 1.723812e-06,
  9.294788e-06, 5.740592e-06, 4.055748e-06, 2.263421e-06, 1.17433e-06, 
    8.964182e-07, 7.44204e-07, 9.900297e-07, 1.578103e-06, 2.440797e-06, 
    2.225877e-06, 4.935137e-06, 1.278752e-05, 2.294654e-05, 1.788398e-05,
  1.265502e-05, 8.21773e-06, 7.093321e-06, 2.499281e-06, 9.339585e-07, 
    4.719262e-07, 4.551272e-07, 8.745171e-07, 1.916179e-06, 3.11917e-06, 
    3.160189e-06, 5.471063e-06, 1.343699e-05, 2.306222e-05, 1.874291e-05,
  2.320087e-05, 1.75364e-05, 2.130457e-05, 2.160958e-05, 2.163746e-06, 
    1.688529e-06, 1.712901e-07, 5.582117e-07, 2.265781e-06, 3.315169e-06, 
    4.444675e-06, 6.206546e-06, 1.524769e-05, 2.220246e-05, 2.091346e-05,
  2.57492e-05, 2.550523e-05, 2.67732e-05, 3.095067e-05, 2.720648e-05, 
    1.301551e-06, 8.082632e-07, 2.399517e-07, 4.189421e-07, 1.122515e-06, 
    4.960079e-06, 7.570431e-06, 1.589122e-05, 2.36309e-05, 2.289235e-05,
  2.269676e-05, 2.493074e-05, 2.233956e-05, 2.518628e-05, 2.536989e-05, 
    2.127062e-05, 1.042751e-05, 4.274701e-06, 4.035893e-06, 1.898802e-06, 
    5.725107e-06, 8.600417e-06, 1.702437e-05, 2.53964e-05, 2.366808e-05,
  1.679301e-05, 1.776438e-05, 1.862263e-05, 1.95958e-05, 2.276614e-05, 
    2.425206e-05, 2.854917e-05, 1.864409e-05, 1.464821e-05, 1.071626e-05, 
    1.231022e-05, 1.372182e-05, 2.226736e-05, 3.077446e-05, 2.137819e-05,
  1.748345e-05, 1.764549e-05, 2.085743e-05, 1.908371e-05, 2.383705e-05, 
    2.49619e-05, 3.664997e-05, 3.516992e-05, 2.489639e-05, 1.867622e-05, 
    1.652955e-05, 1.955823e-05, 3.155662e-05, 3.730317e-05, 1.868592e-05,
  1.99654e-05, 2.347804e-05, 2.505792e-05, 2.209529e-05, 2.449393e-05, 
    3.36563e-05, 3.308253e-05, 4.057371e-05, 1.632113e-05, 1.27715e-05, 
    1.422634e-05, 2.380483e-05, 4.114206e-05, 4.372064e-05, 1.602162e-05,
  2.511337e-05, 2.857622e-05, 3.193465e-05, 2.686151e-05, 3.51518e-05, 
    4.290594e-05, 3.39882e-05, 1.652732e-05, 2.204836e-05, 7.94173e-06, 
    9.938655e-06, 2.784829e-05, 4.868542e-05, 4.593512e-05, 1.35518e-05,
  2.00553e-05, 1.682523e-05, 2.159703e-05, 3.509543e-05, 3.799444e-05, 
    2.557807e-05, 1.626788e-05, 2.430983e-05, 1.306464e-05, 9.032186e-06, 
    1.487042e-05, 3.406893e-05, 4.824257e-05, 4.258291e-05, 1.360451e-05,
  3.441804e-06, 2.248602e-06, 2.13347e-06, 1.339033e-06, 5.473066e-07, 
    3.461908e-07, 1.643129e-07, 1.852453e-07, 2.764124e-07, 1.322685e-06, 
    1.797255e-06, 9.53166e-06, 3.270667e-05, 4.797104e-05, 5.487775e-05,
  8.206268e-06, 7.924887e-06, 5.633647e-06, 2.110813e-06, 2.989478e-07, 
    5.600141e-07, 8.136473e-07, 3.463855e-08, 1.412054e-07, 7.810838e-07, 
    9.284461e-06, 3.316314e-05, 4.603568e-05, 5.651926e-05, 6.719239e-05,
  1.536484e-05, 1.228569e-05, 1.521725e-05, 1.617552e-05, 1.44311e-06, 
    5.366752e-06, 2.715583e-07, 1.995776e-07, 2.242061e-06, 1.323949e-05, 
    3.788839e-05, 5.015494e-05, 3.478992e-05, 4.387964e-05, 7.542977e-05,
  1.765446e-05, 1.765128e-05, 1.879385e-05, 2.18802e-05, 1.82896e-05, 
    2.545962e-06, 2.573609e-06, 1.242096e-06, 5.578131e-06, 3.099021e-05, 
    6.561174e-05, 4.511387e-05, 2.278236e-05, 3.438175e-05, 7.172494e-05,
  2.340587e-05, 1.561691e-05, 1.608593e-05, 1.788854e-05, 2.196848e-05, 
    1.842094e-05, 1.476652e-05, 3.160589e-05, 4.142001e-05, 4.240819e-05, 
    5.919157e-05, 3.242374e-05, 1.963552e-05, 2.973429e-05, 5.989166e-05,
  2.972039e-05, 2.500016e-05, 1.635494e-05, 1.066704e-05, 1.228032e-05, 
    1.945243e-05, 3.611052e-05, 5.224088e-05, 7.312319e-05, 5.738284e-05, 
    3.057516e-05, 1.585257e-05, 1.542073e-05, 3.892674e-05, 5.57297e-05,
  2.786353e-05, 2.893061e-05, 2.495116e-05, 1.523405e-05, 1.223975e-05, 
    1.785093e-05, 3.425019e-05, 5.262253e-05, 5.321305e-05, 3.064218e-05, 
    1.596557e-05, 7.882101e-06, 1.427411e-05, 4.558187e-05, 4.708474e-05,
  2.456331e-05, 3.136875e-05, 3.336933e-05, 3.01795e-05, 1.850014e-05, 
    1.571459e-05, 2.214899e-05, 2.846047e-05, 2.450304e-05, 1.730599e-05, 
    1.098878e-05, 5.244992e-06, 1.462732e-05, 4.26252e-05, 3.123375e-05,
  2.613647e-05, 3.212157e-05, 4.024597e-05, 3.979907e-05, 3.202761e-05, 
    2.220535e-05, 1.83707e-05, 2.252407e-05, 1.964896e-05, 1.354765e-05, 
    7.595691e-06, 4.111536e-06, 1.397441e-05, 3.476398e-05, 1.453811e-05,
  3.189611e-05, 3.482134e-05, 4.223435e-05, 4.670258e-05, 4.342954e-05, 
    3.391573e-05, 2.497582e-05, 2.078951e-05, 1.762332e-05, 1.25958e-05, 
    6.32571e-06, 4.054081e-06, 1.797185e-05, 2.416468e-05, 6.888646e-06,
  1.390293e-05, 5.922469e-06, 3.293599e-06, 1.814476e-06, 1.328199e-07, 
    1.01259e-07, 4.813183e-07, 2.42518e-08, 9.602798e-08, 3.086985e-07, 
    3.456261e-07, 8.815678e-07, 1.034376e-05, 2.6197e-05, 4.000246e-05,
  3.665836e-05, 1.686222e-05, 1.248481e-05, 8.154074e-06, 1.032544e-06, 
    1.490382e-06, 9.019711e-07, 1.275445e-08, 1.016865e-08, 1.285926e-07, 
    2.044929e-07, 3.030663e-06, 1.98068e-05, 3.03539e-05, 2.227765e-05,
  4.032458e-05, 2.947237e-05, 1.804263e-05, 1.951051e-05, 7.682414e-06, 
    1.872583e-06, 8.003541e-07, 1.124607e-08, 6.137686e-09, 1.376276e-08, 
    3.556088e-07, 6.392653e-06, 2.275281e-05, 2.565727e-05, 1.427486e-05,
  4.780438e-05, 4.137945e-05, 3.393898e-05, 2.255439e-05, 2.461684e-05, 
    9.73592e-06, 3.390202e-06, 1.631019e-06, 1.914837e-06, 1.798134e-07, 
    2.462024e-06, 8.638266e-06, 1.691965e-05, 1.53267e-05, 9.415715e-06,
  4.863353e-05, 4.947363e-05, 4.025216e-05, 4.310551e-05, 4.486044e-05, 
    3.241612e-05, 1.244216e-05, 9.424442e-06, 1.497496e-06, 2.796873e-07, 
    4.868403e-06, 9.781922e-06, 1.182257e-05, 5.004738e-06, 5.561863e-06,
  4.825626e-05, 5.495115e-05, 4.832256e-05, 4.540909e-05, 4.682012e-05, 
    4.183661e-05, 3.603e-05, 1.219801e-05, 3.475983e-06, 2.356314e-06, 
    5.651351e-06, 1.007941e-05, 8.219785e-06, 5.229451e-06, 3.407461e-06,
  3.744841e-05, 5.453671e-05, 5.752804e-05, 5.830581e-05, 5.442773e-05, 
    4.760119e-05, 4.217146e-05, 4.258644e-05, 2.190766e-05, 9.08081e-06, 
    6.472112e-06, 1.088073e-05, 6.693135e-06, 6.266546e-06, 2.632731e-06,
  2.51399e-05, 2.266732e-05, 2.611514e-05, 3.163944e-05, 4.406465e-05, 
    4.389333e-05, 3.582659e-05, 3.284128e-05, 2.939561e-05, 2.242893e-05, 
    1.165638e-05, 1.094609e-05, 7.316155e-06, 5.311213e-06, 8.855538e-07,
  1.039104e-05, 1.465953e-05, 1.568413e-05, 1.583832e-05, 2.442549e-05, 
    3.608549e-05, 3.994476e-05, 3.569485e-05, 3.310678e-05, 3.459826e-05, 
    1.9844e-05, 1.237048e-05, 7.834827e-06, 3.790357e-06, 5.833718e-07,
  1.15347e-05, 1.529635e-05, 1.504481e-05, 1.388915e-05, 2.364015e-05, 
    3.724746e-05, 4.664895e-05, 4.983898e-05, 4.522369e-05, 4.381343e-05, 
    3.087224e-05, 1.522457e-05, 1.113167e-05, 6.540736e-06, 8.549744e-07,
  5.008507e-05, 2.516355e-05, 5.985595e-06, 4.089868e-06, 2.018773e-07, 
    1.633976e-08, 1.277063e-07, 2.627375e-08, 1.183735e-08, 1.796471e-08, 
    9.892455e-09, 8.199066e-08, 5.190209e-07, 2.157452e-06, 2.456286e-06,
  6.572218e-05, 5.117661e-05, 2.21608e-05, 7.776404e-06, 2.062726e-06, 
    1.901454e-06, 1.068064e-06, 1.216191e-08, 1.255635e-09, 7.366933e-11, 
    3.760066e-10, 9.398064e-08, 3.537266e-07, 1.839663e-06, 1.800069e-06,
  5.256108e-05, 6.051718e-05, 4.837662e-05, 2.648294e-05, 3.394129e-06, 
    5.692092e-07, 2.941088e-06, 1.674436e-06, 6.610885e-09, 9.409886e-12, 
    5.578776e-09, 3.017779e-08, 2.011351e-07, 1.316871e-06, 1.340122e-06,
  4.776864e-05, 6.915266e-05, 6.651314e-05, 3.472735e-05, 2.642589e-05, 
    3.512146e-06, 7.449457e-07, 3.40775e-06, 1.552858e-06, 1.402689e-08, 
    9.464841e-08, 2.332445e-08, 1.505013e-07, 1.047064e-06, 2.205838e-06,
  4.104929e-05, 8.459441e-05, 9.332711e-05, 6.644207e-05, 3.607185e-05, 
    2.517694e-05, 9.052481e-06, 1.295685e-06, 3.422612e-07, 5.395985e-09, 
    1.10703e-07, 5.9478e-08, 6.068162e-07, 1.197715e-06, 1.587351e-06,
  2.721829e-05, 7.468125e-05, 0.0001051132, 9.326907e-05, 6.273211e-05, 
    3.290532e-05, 2.392613e-05, 5.715423e-06, 7.297054e-07, 1.117709e-06, 
    7.503197e-07, 1.365034e-06, 2.023574e-06, 7.784187e-07, 1.132989e-06,
  3.153306e-05, 5.052637e-05, 9.130991e-05, 0.0001031852, 8.340398e-05, 
    4.832354e-05, 3.111623e-05, 2.28002e-05, 1.318877e-05, 5.089928e-06, 
    2.677283e-06, 2.243297e-06, 2.059552e-06, 6.512782e-07, 1.178354e-06,
  4.964078e-05, 4.695082e-05, 5.558258e-05, 7.478884e-05, 7.961268e-05, 
    6.257987e-05, 4.736431e-05, 3.271292e-05, 2.964822e-05, 1.117349e-05, 
    1.028506e-05, 6.259453e-06, 1.287659e-06, 1.066104e-06, 1.004596e-06,
  3.152233e-05, 3.521531e-05, 4.358233e-05, 4.098921e-05, 3.93182e-05, 
    4.250389e-05, 3.725691e-05, 3.041326e-05, 2.140937e-05, 1.661277e-05, 
    1.610321e-05, 9.625493e-06, 1.785761e-06, 2.144602e-06, 1.438753e-06,
  2.001548e-05, 1.71332e-05, 2.427856e-05, 2.056175e-05, 2.059799e-05, 
    1.780399e-05, 1.548716e-05, 1.714022e-05, 1.364261e-05, 1.640029e-05, 
    1.984144e-05, 1.201296e-05, 5.06038e-06, 2.767102e-06, 1.892e-06,
  1.192025e-05, 1.118469e-05, 6.876136e-06, 4.501471e-06, 1.113498e-06, 
    9.16724e-07, 1.6619e-06, 9.654567e-07, 8.24483e-07, 1.481353e-07, 
    3.347818e-07, 3.311857e-07, 3.571999e-07, 2.972883e-07, 3.59013e-07,
  1.687769e-05, 1.562489e-05, 1.098047e-05, 5.462571e-06, 2.060704e-06, 
    2.496768e-06, 2.256316e-06, 6.313729e-07, 1.78022e-07, 5.537667e-07, 
    1.728941e-07, 2.349667e-07, 2.87035e-07, 2.065316e-07, 1.944958e-07,
  2.66876e-05, 2.393276e-05, 2.144577e-05, 1.452289e-05, 4.440001e-07, 
    1.24517e-06, 9.459379e-07, 1.106821e-06, 2.309884e-07, 1.21338e-07, 
    3.707239e-07, 1.062347e-07, 1.060135e-07, 2.302253e-07, 1.091142e-07,
  3.147129e-05, 3.268941e-05, 3.235709e-05, 1.635549e-05, 1.42777e-05, 
    2.29406e-07, 1.269497e-06, 1.144945e-06, 7.2558e-07, 2.323677e-07, 
    1.205476e-07, 6.194976e-08, 6.939617e-08, 1.170986e-07, 5.368636e-07,
  4.072974e-05, 3.640669e-05, 3.574968e-05, 2.538344e-05, 1.821802e-05, 
    7.957979e-06, 2.614119e-06, 1.452516e-07, 3.836137e-08, 1.386532e-08, 
    2.503565e-07, 7.731126e-08, 4.980705e-08, 1.379862e-07, 2.215762e-07,
  5.722153e-05, 5.68361e-05, 4.961972e-05, 3.695234e-05, 2.480486e-05, 
    1.601458e-05, 8.328122e-06, 6.932445e-07, 1.109989e-09, 6.967645e-08, 
    7.664775e-07, 4.046304e-07, 4.333443e-08, 8.932794e-08, 2.828334e-08,
  5.442121e-05, 4.968644e-05, 4.606237e-05, 4.111139e-05, 3.245896e-05, 
    2.337871e-05, 2.20285e-05, 7.275855e-06, 1.201524e-06, 4.275213e-07, 
    1.592233e-07, 2.393513e-08, 3.419503e-08, 7.699099e-08, 4.348799e-08,
  5.882966e-05, 6.276659e-05, 5.913381e-05, 5.74509e-05, 4.122294e-05, 
    3.194021e-05, 2.412949e-05, 1.762999e-05, 1.524436e-05, 2.97157e-06, 
    3.641538e-07, 7.146139e-08, 4.08794e-08, 6.285274e-08, 5.016123e-08,
  5.158884e-05, 5.186469e-05, 5.253405e-05, 5.230794e-05, 5.179057e-05, 
    4.312865e-05, 3.205866e-05, 2.466595e-05, 2.260085e-05, 1.658788e-06, 
    2.07627e-07, 1.166821e-07, 1.270187e-07, 1.195522e-07, 9.099423e-08,
  3.945362e-05, 3.685265e-05, 3.816534e-05, 4.158928e-05, 4.091776e-05, 
    3.605875e-05, 2.696873e-05, 2.181022e-05, 5.577454e-06, 9.116752e-07, 
    2.03774e-06, 2.891715e-06, 1.456368e-06, 2.866678e-07, 3.433331e-07,
  3.073241e-06, 2.366558e-06, 1.513007e-06, 8.516952e-07, 5.995163e-07, 
    3.736895e-07, 1.955763e-07, 1.161762e-06, 1.189717e-06, 3.610666e-07, 
    8.801287e-08, 2.624878e-07, 8.70703e-08, 6.145421e-08, 9.720491e-08,
  5.187781e-06, 1.940839e-06, 2.177657e-06, 9.129253e-07, 4.323082e-07, 
    2.591953e-07, 7.577924e-07, 4.669051e-07, 4.979319e-07, 1.1911e-06, 
    5.982418e-08, 2.624593e-07, 4.138929e-07, 3.535759e-08, 5.840014e-08,
  1.168266e-05, 4.497601e-06, 5.076377e-06, 2.998086e-06, 6.149458e-07, 
    9.007721e-07, 5.028592e-07, 8.547692e-07, 6.800364e-07, 2.233143e-07, 
    1.900817e-07, 5.358361e-07, 3.469773e-08, 1.265555e-07, 4.027825e-08,
  1.454388e-05, 1.05434e-05, 7.835542e-06, 5.008073e-06, 2.347955e-06, 
    1.438945e-06, 4.8838e-07, 5.371515e-07, 2.523361e-07, 4.29697e-07, 
    9.644338e-08, 4.795116e-08, 5.770566e-08, 1.361887e-07, 1.209629e-07,
  2.17361e-05, 1.759371e-05, 1.24456e-05, 9.091703e-06, 7.483006e-06, 
    4.992925e-06, 3.459793e-06, 2.256041e-07, 2.236122e-07, 1.043666e-07, 
    6.728895e-09, 2.544681e-08, 1.023638e-08, 2.503271e-08, 7.734219e-08,
  2.59555e-05, 2.338458e-05, 1.789666e-05, 1.364557e-05, 1.116113e-05, 
    8.394745e-06, 4.250986e-06, 1.929266e-08, 4.877134e-09, 1.328534e-06, 
    5.783215e-08, 6.298198e-09, 2.389151e-09, 1.724529e-08, 8.390368e-09,
  2.974792e-05, 2.780215e-05, 2.352615e-05, 1.813051e-05, 1.398375e-05, 
    1.318976e-05, 7.266092e-06, 1.072143e-06, 2.903366e-07, 6.913799e-07, 
    4.148361e-07, 1.47799e-08, 9.012204e-09, 2.545121e-08, 2.195858e-08,
  3.963355e-05, 3.178267e-05, 2.699436e-05, 2.167427e-05, 1.633227e-05, 
    1.314862e-05, 1.266015e-05, 1.136738e-05, 5.885985e-06, 2.389195e-07, 
    1.185863e-07, 5.247317e-08, 1.474106e-08, 4.049233e-08, 6.313906e-08,
  4.190197e-05, 3.371961e-05, 3.025317e-05, 2.144376e-05, 1.801519e-05, 
    1.595782e-05, 1.356431e-05, 1.111443e-05, 6.96232e-06, 7.474874e-08, 
    3.373891e-08, 1.920361e-08, 2.033487e-08, 3.577927e-08, 6.564395e-08,
  3.296701e-05, 2.684479e-05, 2.593209e-05, 1.668336e-05, 1.848476e-05, 
    1.548354e-05, 1.193177e-05, 1.052453e-05, 8.915218e-07, 4.809379e-08, 
    2.736487e-07, 1.539635e-08, 2.319605e-08, 2.949299e-08, 4.393018e-08,
  7.335825e-06, 2.02987e-06, 1.58116e-06, 1.901392e-06, 4.837169e-07, 
    2.397131e-07, 7.034442e-07, 7.840907e-07, 9.993695e-07, 3.328494e-07, 
    5.465503e-07, 6.989419e-07, 8.008675e-07, 4.564703e-07, 4.134204e-07,
  1.04633e-05, 5.246503e-06, 6.98223e-06, 2.933819e-06, 5.045604e-09, 
    1.281859e-07, 5.505484e-07, 2.736058e-07, 3.176395e-07, 1.014791e-06, 
    6.984603e-07, 3.876747e-07, 1.157049e-06, 2.163073e-07, 4.310191e-07,
  2.280469e-05, 1.071666e-05, 9.202932e-06, 3.853037e-06, 1.116923e-06, 
    3.109111e-07, 1.417894e-07, 2.037499e-07, 2.913e-07, 1.020897e-07, 
    1.38829e-07, 2.030249e-07, 1.723715e-07, 6.239115e-07, 9.100618e-07,
  3.179514e-05, 2.362019e-05, 1.433156e-05, 1.269374e-05, 9.309621e-06, 
    8.299148e-07, 1.605672e-07, 2.922552e-08, 1.952631e-08, 1.393334e-07, 
    1.860825e-07, 3.525809e-07, 4.992326e-07, 8.581627e-07, 1.689423e-06,
  3.070411e-05, 1.971953e-05, 1.723733e-05, 1.798418e-05, 1.516318e-05, 
    8.193481e-06, 1.270704e-06, 7.044861e-09, 1.402071e-07, 5.012828e-07, 
    2.582908e-07, 2.940715e-07, 4.476748e-07, 6.075943e-07, 2.174946e-06,
  3.937306e-05, 3.314107e-05, 1.905828e-05, 1.934116e-05, 1.727497e-05, 
    1.390737e-05, 5.299637e-06, 3.750081e-09, 3.104486e-08, 4.130384e-07, 
    2.15935e-07, 5.240127e-08, 1.995053e-07, 3.161062e-07, 9.322849e-07,
  5.793567e-05, 4.875657e-05, 3.709278e-05, 2.227954e-05, 1.671234e-05, 
    1.366384e-05, 8.546269e-06, 2.95694e-06, 9.126514e-07, 4.193653e-07, 
    3.188558e-07, 6.234861e-08, 2.099005e-07, 2.041399e-07, 5.566478e-07,
  5.075933e-05, 4.012495e-05, 3.315638e-05, 2.603462e-05, 2.338939e-05, 
    1.754119e-05, 1.144027e-05, 7.938213e-06, 5.819967e-07, 5.940872e-07, 
    1.2432e-07, 7.105508e-07, 3.543229e-07, 3.537544e-07, 4.255529e-07,
  4.466638e-05, 4.264106e-05, 3.610233e-05, 2.793587e-05, 2.134959e-05, 
    1.944736e-05, 1.772488e-05, 9.936564e-06, 8.524823e-07, 2.43423e-07, 
    7.076497e-07, 1.344197e-06, 1.22533e-06, 7.964857e-07, 4.855149e-07,
  3.939582e-05, 3.510565e-05, 2.920582e-05, 2.117453e-05, 1.971162e-05, 
    1.741952e-05, 1.491604e-05, 7.813216e-06, 7.797183e-08, 1.144967e-06, 
    1.944267e-06, 5.039594e-07, 1.119898e-06, 1.837563e-06, 7.033552e-07,
  1.252771e-06, 8.375124e-07, 9.3792e-07, 1.503598e-06, 7.599083e-07, 
    3.280479e-07, 1.143104e-06, 1.485617e-06, 2.555762e-06, 9.023498e-07, 
    9.647041e-07, 1.59505e-06, 1.656455e-06, 1.540151e-06, 1.921917e-06,
  2.338542e-06, 1.919642e-06, 1.679138e-06, 2.362573e-06, 2.031077e-08, 
    2.912851e-07, 9.587612e-07, 9.722777e-07, 9.879318e-07, 3.750803e-06, 
    2.809023e-06, 5.20709e-06, 6.776093e-06, 3.939165e-06, 5.880247e-06,
  9.569389e-06, 4.506298e-06, 5.269639e-06, 3.244941e-06, 2.13405e-06, 
    1.967828e-07, 3.779172e-07, 3.531833e-06, 6.911312e-06, 7.568825e-06, 
    8.75402e-06, 1.005502e-05, 1.152926e-05, 1.235299e-05, 1.490097e-05,
  1.677307e-05, 1.185334e-05, 7.969613e-06, 5.816825e-06, 3.251364e-06, 
    1.832129e-06, 4.181825e-07, 2.510408e-06, 6.046925e-06, 1.278769e-05, 
    1.522248e-05, 1.637108e-05, 1.725318e-05, 1.636214e-05, 1.673411e-05,
  2.395245e-05, 1.534704e-05, 1.283377e-05, 1.245132e-05, 7.376029e-06, 
    4.732473e-06, 1.288454e-06, 5.236937e-07, 2.723011e-06, 9.305335e-06, 
    1.458918e-05, 1.661452e-05, 1.806539e-05, 1.242161e-05, 1.091379e-05,
  2.667155e-05, 1.242287e-05, 1.175075e-05, 1.595041e-05, 1.029429e-05, 
    1.147909e-05, 6.743927e-06, 4.692341e-06, 3.900989e-06, 7.821217e-06, 
    8.927003e-06, 1.266375e-05, 1.416046e-05, 1.08354e-05, 9.019418e-06,
  3.295262e-05, 2.141258e-05, 1.76644e-05, 1.398386e-05, 1.360033e-05, 
    1.261355e-05, 1.098141e-05, 1.020948e-05, 5.755858e-06, 5.445556e-06, 
    5.296864e-06, 7.723022e-06, 9.092464e-06, 9.926157e-06, 8.83274e-06,
  4.780712e-05, 3.235445e-05, 1.997912e-05, 2.031132e-05, 1.758835e-05, 
    1.688655e-05, 1.314818e-05, 5.174766e-06, 2.971013e-06, 2.576548e-06, 
    2.946382e-06, 4.040191e-06, 5.664944e-06, 7.620935e-06, 8.764647e-06,
  5.419815e-05, 3.658526e-05, 3.073385e-05, 1.984753e-05, 1.909718e-05, 
    1.852e-05, 1.158098e-05, 5.595784e-06, 1.065061e-06, 4.384083e-07, 
    1.332644e-06, 1.674156e-06, 2.325124e-06, 3.971503e-06, 4.927203e-06,
  4.593025e-05, 3.283632e-05, 2.477263e-05, 2.0165e-05, 1.656241e-05, 
    1.764775e-05, 1.171203e-05, 3.293611e-06, 6.247342e-08, 5.798095e-07, 
    4.933594e-07, 3.970437e-07, 5.934147e-07, 8.263447e-07, 1.484829e-06,
  1.112142e-06, 3.54557e-06, 4.605015e-07, 1.347457e-06, 2.331187e-06, 
    9.062121e-08, 4.828525e-07, 8.532039e-07, 1.1012e-06, 8.320613e-07, 
    2.103137e-06, 4.063877e-06, 3.783547e-06, 3.04504e-06, 2.513623e-06,
  6.126196e-06, 6.069471e-06, 5.665604e-06, 3.32812e-06, 1.184071e-07, 
    7.417203e-07, 1.507697e-06, 1.326708e-06, 1.254134e-06, 1.607961e-06, 
    1.712898e-06, 2.888592e-06, 3.964086e-06, 2.277851e-06, 1.635985e-06,
  1.414197e-05, 1.169379e-05, 9.327058e-06, 5.701193e-06, 4.938374e-06, 
    1.963227e-07, 7.047632e-07, 6.021728e-06, 6.706148e-06, 4.325289e-06, 
    2.558274e-06, 1.773424e-06, 2.48168e-06, 2.588106e-06, 1.509239e-06,
  1.977463e-05, 1.876228e-05, 1.517132e-05, 1.200371e-05, 1.628599e-05, 
    1.035115e-05, 2.416938e-06, 8.543631e-06, 1.070636e-05, 7.303572e-06, 
    3.288449e-06, 1.016724e-06, 1.157626e-06, 2.082306e-06, 2.222744e-06,
  2.086907e-05, 2.005091e-05, 1.94728e-05, 1.780784e-05, 1.92016e-05, 
    2.360513e-05, 2.014606e-05, 2.449528e-06, 4.046029e-06, 7.049384e-06, 
    5.444609e-06, 1.285588e-06, 8.863589e-07, 2.509549e-06, 1.307088e-06,
  2.119036e-05, 1.884613e-05, 2.122908e-05, 2.257399e-05, 2.248086e-05, 
    2.081177e-05, 2.171321e-05, 1.280129e-05, 1.135616e-05, 1.090607e-05, 
    6.94369e-06, 2.897674e-06, 2.602607e-06, 1.877568e-06, 7.656055e-08,
  2.360382e-05, 2.20822e-05, 2.421967e-05, 2.343425e-05, 2.707424e-05, 
    2.434795e-05, 1.958339e-05, 1.90195e-05, 1.718931e-05, 1.598262e-05, 
    1.229451e-05, 6.855072e-06, 3.498935e-06, 1.965772e-06, 2.935236e-07,
  2.959487e-05, 2.745985e-05, 2.672564e-05, 2.300825e-05, 2.468788e-05, 
    2.267422e-05, 1.965038e-05, 1.670421e-05, 1.443252e-05, 1.308129e-05, 
    1.249658e-05, 9.792674e-06, 5.40615e-06, 3.17512e-06, 2.959017e-06,
  2.950479e-05, 2.791048e-05, 3.334332e-05, 2.677176e-05, 2.082134e-05, 
    1.833197e-05, 1.599642e-05, 1.490201e-05, 1.476985e-05, 1.183649e-05, 
    1.063082e-05, 1.078421e-05, 7.229082e-06, 4.800391e-06, 2.698701e-06,
  2.570229e-05, 2.408132e-05, 2.541181e-05, 1.723715e-05, 1.778953e-05, 
    1.584948e-05, 1.265581e-05, 7.782138e-06, 7.052859e-06, 6.477689e-06, 
    8.239122e-06, 6.1356e-06, 4.855363e-06, 2.701922e-06, 1.236199e-06,
  2.552458e-06, 2.15915e-06, 1.798905e-06, 2.365765e-06, 4.843896e-06, 
    7.345443e-06, 9.850912e-06, 1.247477e-05, 1.165399e-05, 7.167692e-06, 
    3.968814e-06, 2.483094e-06, 2.584634e-06, 1.71713e-06, 1.229449e-06,
  7.695605e-06, 5.262685e-06, 4.70759e-06, 4.684219e-06, 6.122481e-06, 
    9.172004e-06, 1.583769e-05, 1.223481e-05, 8.351922e-06, 6.898809e-06, 
    3.270043e-06, 3.587377e-06, 3.107248e-06, 1.651845e-06, 8.097142e-07,
  1.537914e-05, 8.776921e-06, 1.005283e-05, 7.317123e-06, 1.093442e-05, 
    7.540401e-06, 1.357538e-05, 1.548327e-05, 1.108905e-05, 7.927496e-06, 
    4.640857e-06, 2.441388e-06, 2.903883e-06, 2.125654e-06, 4.374718e-07,
  2.155918e-05, 1.598148e-05, 1.708644e-05, 1.13782e-05, 1.569884e-05, 
    1.263227e-05, 6.775562e-06, 8.431654e-06, 8.983206e-06, 9.890299e-06, 
    4.309178e-06, 1.612541e-06, 1.514312e-06, 1.744063e-06, 9.030067e-07,
  2.178261e-05, 1.760431e-05, 1.921961e-05, 1.741105e-05, 1.611788e-05, 
    1.874971e-05, 1.234345e-05, 1.099162e-06, 1.750882e-06, 4.536674e-06, 
    3.689266e-06, 1.926766e-06, 1.355238e-06, 1.272187e-06, 7.951882e-07,
  1.931619e-05, 1.662285e-05, 1.765597e-05, 1.855838e-05, 1.697806e-05, 
    1.50701e-05, 1.358719e-05, 5.955847e-06, 3.331436e-06, 4.310376e-06, 
    2.911676e-06, 2.245661e-06, 2.251877e-06, 9.027752e-07, 1.408403e-07,
  2.308085e-05, 2.226843e-05, 1.991893e-05, 1.8259e-05, 1.767766e-05, 
    1.536686e-05, 1.158688e-05, 9.785806e-06, 7.270974e-06, 4.455776e-06, 
    4.325909e-06, 3.233569e-06, 1.986676e-06, 3.148243e-07, 1.884659e-07,
  2.831535e-05, 2.86454e-05, 2.356997e-05, 2.069365e-05, 1.927904e-05, 
    1.879985e-05, 1.468801e-05, 1.123609e-05, 6.235552e-06, 4.131061e-06, 
    4.314956e-06, 3.284491e-06, 1.641875e-06, 5.555129e-07, 1.749388e-07,
  3.034073e-05, 2.875175e-05, 3.194662e-05, 2.533752e-05, 2.113211e-05, 
    1.921649e-05, 1.644496e-05, 1.153368e-05, 6.250107e-06, 4.253925e-06, 
    4.389092e-06, 3.186372e-06, 1.953152e-06, 9.16301e-07, 1.430723e-07,
  2.405831e-05, 1.997682e-05, 2.47583e-05, 2.443882e-05, 2.144922e-05, 
    1.684965e-05, 1.315336e-05, 1.001868e-05, 6.659676e-06, 4.224592e-06, 
    6.751591e-06, 2.749673e-06, 9.513836e-07, 1.918721e-07, 2.39006e-08,
  1.347232e-06, 1.014448e-06, 2.557354e-07, 1.458039e-06, 4.032937e-07, 
    1.263928e-06, 2.128506e-06, 2.557943e-06, 3.963738e-06, 2.77404e-06, 
    2.673295e-06, 3.436824e-06, 2.091077e-06, 6.008461e-07, 3.483736e-07,
  4.061891e-06, 3.778237e-06, 4.207242e-06, 3.237249e-06, 1.845034e-06, 
    1.895464e-06, 2.777415e-06, 2.63453e-06, 2.728123e-06, 3.256454e-06, 
    1.235441e-06, 2.527102e-06, 1.230744e-06, 4.493284e-08, 1.104442e-07,
  1.256123e-05, 8.516502e-06, 1.110963e-05, 8.409015e-06, 9.539342e-06, 
    2.5892e-06, 2.257342e-06, 4.237612e-06, 4.184744e-06, 3.067157e-06, 
    2.13256e-06, 1.496265e-06, 1.281501e-06, 5.072346e-07, 1.228846e-08,
  2.147782e-05, 1.997599e-05, 2.113416e-05, 1.958014e-05, 1.865577e-05, 
    9.521503e-06, 2.414902e-06, 2.234632e-06, 2.22406e-06, 2.550655e-06, 
    8.7508e-07, 1.595376e-07, 4.614181e-07, 3.125099e-07, 2.100055e-08,
  2.521423e-05, 2.280263e-05, 2.46775e-05, 2.648572e-05, 2.498798e-05, 
    2.298889e-05, 1.136911e-05, 1.026843e-06, 1.157843e-06, 1.397946e-06, 
    6.2328e-07, 1.195163e-07, 2.927995e-08, 3.387267e-08, 2.06562e-11,
  2.460203e-05, 2.22305e-05, 2.50402e-05, 2.884415e-05, 2.869389e-05, 
    2.536679e-05, 2.238742e-05, 5.932524e-06, 1.707397e-06, 5.421876e-06, 
    6.481553e-07, 2.555888e-07, 1.033083e-08, 3.421521e-10, 7.490733e-11,
  2.62968e-05, 2.229375e-05, 2.40784e-05, 2.549287e-05, 3.072757e-05, 
    2.725783e-05, 2.102322e-05, 1.55967e-05, 9.307252e-06, 4.677515e-06, 
    2.796464e-06, 5.754954e-07, 1.140426e-09, 7.17395e-12, 7.941422e-11,
  2.776776e-05, 1.828416e-05, 2.062798e-05, 2.257918e-05, 2.393556e-05, 
    2.515766e-05, 2.065335e-05, 1.498998e-05, 8.437606e-06, 2.945273e-06, 
    2.083955e-06, 2.917063e-07, 1.297842e-09, 6.280661e-11, 2.32873e-10,
  3.045973e-05, 1.835553e-05, 2.214342e-05, 2.20918e-05, 2.077199e-05, 
    2.056131e-05, 1.958847e-05, 1.546222e-05, 6.250671e-06, 2.578156e-06, 
    1.357401e-06, 3.39172e-07, 1.852274e-09, 1.772703e-10, 8.727929e-09,
  2.465724e-05, 1.582496e-05, 1.846385e-05, 1.576286e-05, 1.919098e-05, 
    1.684388e-05, 1.587764e-05, 1.221861e-05, 5.494327e-06, 4.76079e-06, 
    3.144693e-06, 3.268055e-07, 3.082157e-09, 2.344748e-10, 5.643008e-10,
  2.358616e-07, 8.165462e-07, 5.380934e-07, 3.924926e-06, 6.501504e-06, 
    6.183597e-06, 5.321049e-06, 6.272162e-06, 7.25333e-06, 4.014978e-06, 
    2.372261e-06, 1.828642e-06, 8.024061e-07, 1.859351e-07, 1.710504e-07,
  2.558028e-06, 1.589662e-06, 2.056513e-06, 2.050737e-06, 4.153948e-06, 
    4.795448e-06, 6.086398e-06, 4.677413e-06, 5.318506e-06, 5.471278e-06, 
    2.702618e-06, 2.507168e-06, 1.907453e-06, 8.743522e-08, 5.300605e-08,
  9.141938e-06, 7.563072e-06, 7.763216e-06, 3.416749e-06, 4.576954e-06, 
    1.889539e-06, 2.16689e-06, 5.076333e-06, 6.095445e-06, 5.945201e-06, 
    4.007608e-06, 1.682742e-06, 1.491973e-06, 7.605752e-07, 8.250384e-08,
  1.852392e-05, 1.830183e-05, 1.721621e-05, 1.332704e-05, 8.324745e-06, 
    6.477175e-06, 1.612869e-06, 2.127661e-06, 4.59142e-06, 4.593286e-06, 
    2.976635e-06, 1.437665e-07, 2.205412e-08, 5.873448e-07, 2.527457e-07,
  2.367655e-05, 2.212014e-05, 1.776443e-05, 2.069008e-05, 1.947086e-05, 
    1.074002e-05, 1.27926e-05, 1.376854e-06, 8.181371e-07, 2.046013e-06, 
    1.195057e-06, 8.580746e-08, 9.973472e-09, 1.596534e-07, 7.087739e-08,
  2.696196e-05, 2.666415e-05, 2.238567e-05, 2.173985e-05, 2.148462e-05, 
    1.619419e-05, 1.634643e-05, 4.333019e-06, 1.836162e-06, 4.790576e-06, 
    6.573726e-07, 1.4337e-08, 5.633503e-09, 2.283632e-09, 2.073326e-09,
  3.515388e-05, 3.121447e-05, 2.318072e-05, 1.838692e-05, 1.784801e-05, 
    2.121026e-05, 1.826877e-05, 1.284254e-05, 7.944062e-06, 3.86668e-06, 
    1.965474e-06, 4.474676e-07, 1.928864e-09, 1.275504e-09, 9.323098e-10,
  3.504107e-05, 3.170142e-05, 2.609515e-05, 1.931303e-05, 1.729518e-05, 
    2.107061e-05, 2.20039e-05, 1.792671e-05, 7.369346e-06, 1.27106e-06, 
    3.496119e-07, 1.262207e-07, 5.20471e-09, 9.545341e-09, 1.00648e-08,
  3.067935e-05, 3.093492e-05, 2.887694e-05, 1.954079e-05, 1.595342e-05, 
    1.802334e-05, 1.858544e-05, 1.510136e-05, 3.206382e-06, 1.018466e-07, 
    2.497503e-08, 3.393588e-09, 7.038428e-09, 9.34663e-09, 6.292087e-08,
  2.511361e-05, 2.324422e-05, 2.274147e-05, 1.484809e-05, 1.206e-05, 
    1.287164e-05, 1.136386e-05, 5.989634e-06, 1.194798e-06, 3.214727e-07, 
    2.89878e-06, 2.508068e-07, 4.820589e-09, 5.52944e-09, 1.514979e-08,
  3.934951e-07, 6.524153e-07, 2.234211e-07, 2.490402e-06, 2.919966e-06, 
    2.019521e-06, 1.926113e-06, 1.004136e-06, 9.735878e-07, 2.806279e-07, 
    5.691753e-08, 1.121515e-06, 1.311436e-06, 2.905879e-08, 3.016254e-08,
  2.17624e-06, 1.697974e-06, 2.512345e-06, 3.217137e-07, 2.500318e-06, 
    1.971847e-06, 1.072272e-06, 1.163562e-06, 8.787337e-07, 9.577633e-07, 
    3.668963e-07, 1.746148e-06, 2.322454e-06, 6.511851e-08, 6.502736e-08,
  7.84705e-06, 5.687995e-06, 4.559824e-06, 3.074165e-06, 5.536202e-06, 
    2.004235e-06, 4.04592e-07, 1.717216e-06, 1.39425e-06, 1.087664e-06, 
    6.86765e-07, 1.053573e-06, 1.507292e-06, 9.026316e-07, 8.861392e-08,
  1.606399e-05, 1.450124e-05, 1.417532e-05, 1.277952e-05, 8.033511e-06, 
    1.367236e-05, 1.772106e-06, 1.074514e-06, 2.424573e-06, 5.944769e-07, 
    1.176258e-07, 2.723675e-07, 4.531439e-07, 1.480822e-06, 8.903053e-07,
  2.115738e-05, 1.806476e-05, 1.439847e-05, 1.406802e-05, 1.656427e-05, 
    1.286967e-05, 1.951705e-05, 1.454745e-06, 2.762176e-07, 3.018973e-07, 
    4.132153e-08, 2.397336e-08, 2.275477e-07, 6.511359e-07, 8.683891e-07,
  2.931543e-05, 2.125483e-05, 1.910811e-05, 1.7223e-05, 1.608443e-05, 
    1.89952e-05, 1.532852e-05, 7.289399e-06, 3.476653e-07, 2.358852e-06, 
    2.256171e-06, 4.453416e-07, 2.871559e-08, 7.924129e-08, 3.104552e-08,
  4.239439e-05, 4.290642e-05, 2.507352e-05, 1.837322e-05, 1.558391e-05, 
    1.451543e-05, 1.988629e-05, 8.43683e-06, 1.00753e-05, 4.554372e-06, 
    3.094627e-06, 2.928435e-07, 1.485874e-09, 4.729543e-08, 1.632183e-08,
  6.147671e-05, 5.632774e-05, 3.214338e-05, 2.206984e-05, 1.659191e-05, 
    1.522864e-05, 1.506203e-05, 1.915707e-05, 9.749261e-06, 1.820049e-06, 
    2.017071e-07, 1.459645e-07, 3.034831e-08, 1.113901e-07, 6.938789e-08,
  7.563406e-05, 5.382991e-05, 3.638635e-05, 2.306803e-05, 1.802358e-05, 
    1.257249e-05, 1.328666e-05, 1.024797e-05, 3.353842e-06, 1.392007e-06, 
    2.62087e-07, 6.272787e-07, 2.372734e-07, 2.055447e-07, 1.334594e-07,
  6.154044e-05, 4.402497e-05, 2.696583e-05, 2.39472e-05, 1.642149e-05, 
    6.159868e-06, 3.448923e-06, 3.776082e-06, 3.192862e-06, 1.88696e-06, 
    2.60605e-06, 2.69449e-06, 5.120091e-07, 1.092759e-06, 5.619226e-08,
  3.686472e-05, 2.733292e-05, 1.363675e-05, 4.560141e-06, 2.866656e-06, 
    1.184041e-06, 7.614792e-07, 5.597404e-07, 6.211265e-07, 6.142898e-08, 
    1.496363e-07, 1.727356e-07, 2.426687e-07, 1.070902e-07, 8.748647e-08,
  3.906028e-05, 2.919574e-05, 1.919998e-05, 7.50029e-06, 2.114379e-06, 
    1.489987e-06, 5.162856e-07, 2.43053e-07, 7.210308e-07, 7.037502e-07, 
    1.01088e-07, 1.117096e-06, 9.282923e-07, 8.084503e-08, 1.228752e-07,
  4.601111e-05, 3.717118e-05, 2.751089e-05, 1.282675e-05, 3.580954e-06, 
    1.25989e-06, 5.407072e-07, 4.223533e-07, 3.669296e-07, 3.866951e-07, 
    8.344631e-07, 1.934337e-07, 2.929111e-07, 6.599143e-07, 2.465422e-07,
  5.537603e-05, 4.564738e-05, 3.732232e-05, 1.829582e-05, 1.539754e-05, 
    2.033031e-06, 5.787447e-07, 4.094491e-07, 9.331018e-08, 2.583601e-08, 
    6.216057e-08, 2.118923e-07, 1.291421e-06, 1.079532e-06, 7.948938e-07,
  6.473818e-05, 5.806355e-05, 4.112702e-05, 2.62338e-05, 2.331941e-05, 
    1.276604e-05, 7.58483e-06, 4.534107e-07, 2.253688e-08, 1.424144e-09, 
    3.327331e-09, 1.170286e-07, 7.886405e-07, 1.138015e-06, 7.32434e-07,
  7.598235e-05, 7.4142e-05, 5.721115e-05, 3.497636e-05, 2.618595e-05, 
    2.290206e-05, 1.615013e-05, 6.69227e-06, 2.78449e-07, 1.220176e-06, 
    2.727195e-06, 1.184523e-06, 1.801614e-07, 6.880236e-07, 4.459478e-07,
  7.135195e-05, 8.860392e-05, 6.474989e-05, 4.768377e-05, 3.387695e-05, 
    2.207626e-05, 2.106329e-05, 1.130463e-05, 9.950125e-06, 1.854864e-06, 
    1.540732e-06, 1.091959e-08, 1.237548e-08, 5.098772e-07, 2.727248e-07,
  6.901781e-05, 8.672155e-05, 8.351902e-05, 5.343434e-05, 3.436144e-05, 
    3.063527e-05, 2.111181e-05, 2.021228e-05, 7.632048e-06, 3.295808e-06, 
    4.47746e-07, 1.674789e-07, 1.152751e-08, 2.676243e-07, 3.17143e-07,
  7.130524e-05, 9.820643e-05, 7.831037e-05, 5.447262e-05, 4.555431e-05, 
    2.77862e-05, 2.118167e-05, 1.145065e-05, 1.90642e-06, 3.047608e-06, 
    1.981309e-06, 2.081708e-06, 4.196041e-07, 3.27136e-07, 2.862672e-07,
  5.921522e-05, 6.407696e-05, 6.117031e-05, 3.616198e-05, 2.757736e-05, 
    1.666769e-05, 1.356218e-05, 1.83475e-06, 8.002511e-07, 2.039206e-06, 
    3.313122e-06, 4.314722e-06, 3.846195e-06, 1.606849e-06, 3.029924e-07,
  1.727584e-05, 1.783226e-05, 2.151484e-05, 1.766621e-05, 8.247745e-06, 
    1.5377e-06, 1.051282e-06, 9.220714e-07, 1.554286e-06, 1.062714e-06, 
    4.048704e-07, 7.868399e-07, 1.96453e-07, 1.002768e-07, 9.349038e-08,
  2.20351e-05, 2.049738e-05, 1.992336e-05, 1.761146e-05, 7.209318e-06, 
    1.574534e-06, 4.511884e-07, 5.680934e-07, 1.506001e-06, 2.161879e-06, 
    9.131718e-07, 1.397488e-06, 1.071451e-06, 8.888932e-08, 1.87324e-07,
  2.236166e-05, 2.506173e-05, 1.997754e-05, 1.754086e-05, 5.440923e-06, 
    9.418457e-07, 5.361485e-07, 1.326528e-06, 1.952712e-06, 2.79702e-06, 
    2.103157e-06, 1.191515e-06, 1.5544e-06, 5.945546e-07, 2.949643e-07,
  3.605475e-05, 3.27434e-05, 2.538863e-05, 2.365433e-05, 1.367126e-05, 
    7.889697e-07, 3.962339e-07, 7.545084e-07, 9.369029e-07, 2.15505e-06, 
    1.574619e-06, 6.823528e-07, 7.229659e-07, 1.020455e-06, 7.383022e-07,
  3.242931e-05, 3.664857e-05, 3.455882e-05, 2.964278e-05, 3.186969e-05, 
    1.533349e-05, 3.93238e-06, 1.324823e-07, 1.04793e-07, 3.44336e-07, 
    7.935907e-07, 1.023225e-06, 4.110543e-07, 9.040271e-07, 9.481369e-07,
  2.681882e-05, 5.018283e-05, 3.554521e-05, 4.811304e-05, 2.954745e-05, 
    2.11076e-05, 1.714936e-05, 1.968622e-06, 8.026054e-08, 1.698067e-06, 
    2.345081e-06, 1.764408e-06, 3.76234e-07, 4.560492e-07, 6.788222e-07,
  3.128219e-05, 5.530247e-05, 5.172516e-05, 4.173264e-05, 4.930487e-05, 
    2.958704e-05, 3.037651e-05, 1.007337e-05, 3.891791e-06, 2.066825e-06, 
    1.963652e-06, 4.632722e-07, 6.839986e-07, 4.793139e-07, 5.261955e-07,
  3.140712e-05, 4.882808e-05, 6.843861e-05, 3.361714e-05, 5.364511e-05, 
    3.89557e-05, 2.347362e-05, 2.218176e-05, 7.136221e-06, 3.095183e-07, 
    5.021635e-07, 3.805798e-07, 4.186221e-07, 5.666041e-07, 5.682443e-07,
  2.97787e-05, 4.41751e-05, 7.808138e-05, 3.566123e-05, 3.694383e-05, 
    5.154208e-05, 3.183902e-05, 2.133209e-05, 8.109664e-07, 1.923197e-07, 
    2.449694e-07, 8.835124e-07, 4.341543e-07, 4.930349e-07, 4.935568e-07,
  1.505346e-05, 2.628838e-05, 5.054371e-05, 3.035276e-05, 2.541264e-05, 
    3.408323e-05, 3.409186e-05, 9.106197e-06, 4.313129e-07, 2.886059e-07, 
    4.665609e-06, 2.611712e-06, 2.081787e-06, 3.090098e-07, 3.480739e-07,
  9.011866e-06, 1.793589e-05, 2.077088e-05, 2.263558e-05, 1.413072e-05, 
    4.156075e-06, 3.637418e-06, 2.04815e-06, 1.147807e-06, 6.105938e-07, 
    2.837343e-07, 7.971755e-07, 7.00962e-07, 3.847209e-07, 4.301484e-07,
  8.489352e-06, 1.491329e-05, 2.296259e-05, 2.77654e-05, 1.744183e-05, 
    4.993592e-06, 2.608664e-06, 1.283856e-06, 1.62824e-06, 1.742678e-06, 
    9.394223e-07, 1.267733e-06, 9.738752e-07, 6.661848e-08, 2.911068e-07,
  1.083249e-05, 1.299019e-05, 2.084839e-05, 2.845617e-05, 1.479491e-05, 
    3.486934e-06, 1.848393e-06, 2.404198e-06, 2.85022e-06, 3.285332e-06, 
    2.01258e-06, 1.57169e-06, 1.361628e-06, 6.309712e-07, 3.868558e-07,
  2.495086e-05, 2.256849e-05, 2.295624e-05, 2.804057e-05, 2.264438e-05, 
    3.024682e-06, 5.790187e-07, 1.617377e-06, 2.011133e-06, 3.226436e-06, 
    1.892884e-06, 1.18052e-06, 1.139964e-06, 1.226692e-06, 7.949953e-07,
  2.65964e-05, 2.681798e-05, 3.302272e-05, 3.020379e-05, 3.422012e-05, 
    2.125945e-05, 3.826875e-06, 1.129427e-07, 1.776686e-07, 3.225518e-07, 
    6.000564e-07, 1.060113e-06, 8.716748e-07, 1.048126e-06, 1.013789e-06,
  2.939174e-05, 3.039322e-05, 4.157834e-05, 3.505901e-05, 3.847757e-05, 
    3.110303e-05, 2.036248e-05, 3.448411e-06, 6.010942e-07, 3.407709e-06, 
    3.01777e-06, 1.488925e-06, 1.119851e-06, 8.137294e-07, 1.009279e-06,
  2.529943e-05, 2.292465e-05, 4.371961e-05, 3.980236e-05, 4.676701e-05, 
    3.140205e-05, 2.870442e-05, 1.210662e-05, 5.472923e-06, 6.111432e-06, 
    3.88523e-06, 1.321862e-06, 1.109346e-06, 7.006325e-07, 8.806687e-07,
  1.52487e-05, 1.552281e-05, 3.189369e-05, 5.586964e-05, 4.305723e-05, 
    4.191393e-05, 1.986225e-05, 1.928362e-05, 9.035795e-06, 2.7633e-06, 
    1.925863e-06, 1.142101e-06, 7.73368e-07, 6.878609e-07, 9.164867e-07,
  9.701825e-06, 1.503796e-05, 3.037109e-05, 6.073593e-05, 3.734962e-05, 
    3.971306e-05, 4.406432e-05, 2.025502e-05, 4.933118e-06, 9.353214e-08, 
    2.432108e-07, 1.093841e-06, 8.966994e-07, 9.409017e-07, 1.004302e-06,
  1.227696e-05, 2.340704e-05, 2.730312e-05, 4.57008e-05, 2.926296e-05, 
    2.603796e-05, 3.080857e-05, 9.716446e-06, 1.080989e-07, 2.023652e-07, 
    4.729926e-06, 2.057284e-06, 1.66888e-06, 1.624348e-06, 1.362701e-06,
  3.439972e-05, 3.397624e-05, 2.684644e-05, 2.280473e-05, 2.062031e-05, 
    2.033759e-05, 1.461812e-05, 1.043485e-05, 4.143083e-06, 5.538785e-07, 
    2.945768e-08, 3.956561e-07, 2.066254e-07, 1.647521e-07, 4.825998e-07,
  4.205255e-05, 3.320817e-05, 3.279222e-05, 2.67196e-05, 2.682936e-05, 
    2.59862e-05, 1.554594e-05, 1.097291e-05, 5.85083e-06, 2.18375e-06, 
    9.14774e-07, 1.150905e-06, 9.578766e-07, 2.653498e-08, 2.169097e-07,
  5.118552e-05, 3.956469e-05, 3.390251e-05, 3.208868e-05, 3.02592e-05, 
    2.640777e-05, 1.327358e-05, 8.861181e-06, 6.477785e-06, 3.759488e-06, 
    1.466129e-06, 1.283794e-06, 1.138488e-06, 7.62153e-07, 3.868608e-07,
  5.862736e-05, 5.202702e-05, 3.73052e-05, 2.982024e-05, 3.586995e-05, 
    1.828423e-05, 7.936607e-06, 3.378991e-06, 3.522752e-06, 3.61322e-06, 
    2.144294e-06, 1.040322e-06, 8.775048e-07, 1.094588e-06, 8.079011e-07,
  4.65959e-05, 5.286422e-05, 5.120499e-05, 4.041467e-05, 4.009539e-05, 
    3.241794e-05, 9.96052e-06, 1.112204e-06, 8.639267e-07, 8.309071e-07, 
    8.046028e-07, 9.128798e-07, 9.382392e-07, 8.208407e-07, 8.780677e-07,
  2.500949e-05, 4.279265e-05, 6.222274e-05, 5.937513e-05, 5.380376e-05, 
    3.592588e-05, 2.397249e-05, 3.695163e-06, 7.891102e-07, 3.072846e-06, 
    2.46654e-06, 1.450807e-06, 1.193941e-06, 7.647931e-07, 7.005365e-07,
  1.483599e-05, 2.867696e-05, 5.545914e-05, 7.618361e-05, 5.368235e-05, 
    4.23256e-05, 2.559114e-05, 1.048902e-05, 5.327532e-06, 7.509484e-06, 
    3.989585e-06, 1.922968e-06, 1.292183e-06, 6.773727e-07, 4.107363e-07,
  2.681781e-05, 3.750298e-05, 5.957041e-05, 7.313056e-05, 4.638968e-05, 
    3.764127e-05, 2.868476e-05, 1.215743e-05, 6.26225e-06, 4.906891e-06, 
    2.115077e-06, 1.72745e-06, 1.313342e-06, 6.217955e-07, 2.807333e-07,
  3.409578e-05, 4.470529e-05, 6.006728e-05, 5.937005e-05, 3.856579e-05, 
    3.13372e-05, 3.123286e-05, 1.559247e-05, 2.33431e-06, 4.332318e-08, 
    8.337719e-08, 1.344109e-06, 1.064435e-06, 5.713242e-07, 2.889131e-07,
  2.877379e-05, 2.949757e-05, 4.626719e-05, 3.395131e-05, 3.079095e-05, 
    2.480513e-05, 2.192289e-05, 9.878159e-06, 3.808024e-07, 1.140714e-07, 
    3.968062e-06, 1.638429e-06, 1.525093e-06, 1.300395e-06, 1.261077e-06,
  3.489617e-05, 3.76153e-05, 3.64857e-05, 4.214638e-05, 3.955129e-05, 
    3.220703e-05, 2.483277e-05, 2.028901e-05, 1.759011e-05, 1.334821e-05, 
    7.723666e-06, 4.607462e-06, 2.078176e-06, 7.702874e-07, 2.244778e-06,
  4.938705e-05, 3.365944e-05, 3.632316e-05, 3.885182e-05, 3.751439e-05, 
    3.01804e-05, 2.631177e-05, 2.342472e-05, 1.874908e-05, 1.569845e-05, 
    8.212217e-06, 4.613676e-06, 1.434909e-06, 1.70415e-07, 8.029832e-07,
  3.48266e-05, 1.927679e-05, 2.25842e-05, 2.436517e-05, 2.40804e-05, 
    1.855825e-05, 2.596744e-05, 2.783251e-05, 2.232192e-05, 1.814861e-05, 
    8.73673e-06, 3.942042e-06, 1.342691e-06, 1.854465e-07, 3.111084e-07,
  2.054638e-05, 2.139738e-05, 2.390952e-05, 2.345662e-05, 2.521404e-05, 
    1.294438e-05, 1.572842e-05, 1.35932e-05, 1.315301e-05, 1.378168e-05, 
    8.211482e-06, 2.040712e-06, 3.860051e-07, 2.08223e-07, 1.70478e-07,
  2.562251e-05, 2.236375e-05, 3.402064e-05, 3.666865e-05, 2.771881e-05, 
    2.454395e-05, 1.025637e-05, 1.539959e-06, 1.597272e-06, 5.919272e-06, 
    5.022483e-06, 6.332379e-07, 1.283055e-07, 1.028282e-07, 1.211856e-07,
  2.428652e-05, 2.78834e-05, 3.906164e-05, 4.862956e-05, 3.999077e-05, 
    3.487193e-05, 2.06227e-05, 4.739618e-06, 4.375791e-06, 9.755244e-06, 
    5.667634e-06, 2.032888e-06, 6.817284e-07, 5.506618e-08, 6.617213e-08,
  1.588411e-05, 2.451831e-05, 6.551806e-05, 4.307999e-05, 4.267272e-05, 
    3.978976e-05, 3.008568e-05, 1.038271e-05, 1.032227e-05, 1.203132e-05, 
    8.092633e-06, 2.483627e-06, 8.451972e-07, 3.799842e-08, 4.362499e-09,
  2.461108e-05, 3.808535e-05, 6.015057e-05, 5.069119e-05, 4.737731e-05, 
    4.009156e-05, 2.354779e-05, 1.590921e-05, 8.01531e-06, 4.875297e-06, 
    3.281822e-06, 1.843857e-06, 4.592706e-07, 1.241687e-07, 3.542796e-08,
  6.680486e-05, 7.180852e-05, 8.518304e-05, 6.108966e-05, 4.781898e-05, 
    3.368383e-05, 1.934181e-05, 1.567175e-05, 1.85009e-06, 1.522786e-06, 
    1.286063e-06, 1.25735e-06, 8.388487e-07, 4.353774e-07, 1.473516e-07,
  4.943025e-05, 4.836696e-05, 4.701743e-05, 3.97577e-05, 3.565191e-05, 
    3.298939e-05, 1.39644e-05, 9.618408e-06, 3.109581e-06, 1.240445e-06, 
    5.317542e-06, 2.280449e-06, 1.65508e-06, 9.791851e-07, 5.215867e-07,
  1.406451e-05, 1.109358e-05, 1.132208e-05, 1.183235e-05, 1.135346e-05, 
    1.321232e-05, 1.220186e-05, 1.205615e-05, 1.082208e-05, 8.041744e-06, 
    8.592227e-06, 1.28508e-05, 1.62025e-05, 1.655742e-05, 1.624797e-05,
  2.47321e-05, 1.840508e-05, 2.340351e-05, 2.801609e-05, 2.576329e-05, 
    1.364234e-05, 9.737825e-06, 1.244401e-05, 9.844811e-06, 1.057979e-05, 
    1.200492e-05, 1.405387e-05, 1.293133e-05, 8.445063e-06, 1.003183e-05,
  2.123641e-05, 1.292402e-05, 2.71319e-05, 4.069007e-05, 3.450618e-05, 
    1.312558e-05, 1.501109e-05, 2.471553e-05, 1.301798e-05, 8.915944e-06, 
    1.063845e-05, 1.127804e-05, 1.082102e-05, 8.649772e-06, 7.484937e-06,
  1.812652e-05, 1.857316e-05, 2.40834e-05, 2.142298e-05, 3.62408e-05, 
    2.446789e-05, 2.570682e-05, 2.208178e-05, 7.597278e-06, 6.447975e-06, 
    9.0437e-06, 8.554561e-06, 8.48986e-06, 7.41965e-06, 4.173972e-06,
  2.365997e-05, 2.17471e-05, 2.32396e-05, 3.059255e-05, 2.845824e-05, 
    5.389034e-05, 2.960989e-05, 1.125112e-05, 4.18922e-06, 6.943175e-06, 
    8.746532e-06, 6.344747e-06, 5.932595e-06, 2.923701e-06, 1.790649e-06,
  1.831407e-05, 1.90504e-05, 2.241578e-05, 3.864246e-05, 6.308366e-05, 
    4.765758e-05, 2.979364e-05, 1.011425e-05, 5.777769e-06, 8.174936e-06, 
    6.479737e-06, 6.698757e-06, 5.039654e-06, 2.524303e-06, 6.201022e-07,
  2.100928e-05, 3.096402e-05, 4.84101e-05, 7.972237e-05, 5.030916e-05, 
    3.05408e-05, 2.260294e-05, 1.211199e-05, 8.089026e-06, 1.140052e-05, 
    1.112606e-05, 8.535675e-06, 4.532767e-06, 1.954024e-06, 1.810541e-08,
  2.070288e-05, 2.997324e-05, 4.435879e-05, 3.64572e-05, 3.300522e-05, 
    2.350392e-05, 2.041471e-05, 1.436458e-05, 6.440078e-06, 5.023591e-06, 
    9.011676e-06, 7.629958e-06, 3.330706e-06, 1.120391e-06, 9.677117e-09,
  2.973454e-05, 2.526979e-05, 2.859136e-05, 3.118788e-05, 2.204823e-05, 
    2.143289e-05, 1.993034e-05, 1.358394e-05, 1.430732e-06, 1.888889e-06, 
    4.514154e-06, 4.771494e-06, 2.395519e-06, 3.465383e-07, 2.179551e-07,
  2.654372e-05, 3.056698e-05, 3.305851e-05, 3.377455e-05, 3.195368e-05, 
    2.00747e-05, 1.116953e-05, 7.332625e-06, 2.527977e-06, 1.47781e-06, 
    5.32051e-06, 4.285611e-06, 2.070791e-06, 3.210569e-07, 2.85799e-07,
  3.702089e-06, 5.316386e-06, 8.134696e-06, 9.880708e-06, 7.71784e-06, 
    8.378558e-06, 6.056211e-06, 3.094808e-06, 1.87618e-06, 1.442737e-06, 
    1.252986e-06, 3.730044e-06, 6.585742e-06, 7.173988e-06, 8.781169e-06,
  5.491135e-07, 1.297026e-06, 3.645077e-06, 9.370394e-06, 1.434763e-05, 
    1.302154e-05, 9.565899e-06, 6.345537e-06, 3.138733e-06, 2.712168e-06, 
    2.861397e-06, 4.542607e-06, 5.935146e-06, 4.643411e-06, 9.436762e-06,
  7.501195e-06, 4.1526e-06, 1.261207e-06, 3.51954e-06, 1.120214e-05, 
    1.830454e-05, 1.591342e-05, 2.120201e-05, 1.039518e-05, 5.051635e-06, 
    4.566521e-06, 6.242083e-06, 7.528526e-06, 8.074334e-06, 1.118539e-05,
  9.532765e-06, 1.519606e-05, 2.033014e-05, 1.195482e-05, 6.602255e-06, 
    1.76656e-05, 2.815549e-05, 2.05478e-05, 7.683001e-06, 5.195987e-06, 
    6.703314e-06, 6.506468e-06, 7.03689e-06, 8.66882e-06, 8.450774e-06,
  1.051666e-05, 1.502439e-05, 1.770276e-05, 2.006637e-05, 1.093982e-05, 
    3.022703e-05, 3.484886e-05, 1.196552e-05, 3.067248e-06, 8.290608e-06, 
    1.209116e-05, 5.799917e-06, 6.121054e-06, 4.724157e-06, 5.633834e-06,
  1.243222e-05, 1.830521e-05, 1.947173e-05, 2.839124e-05, 2.952539e-05, 
    3.771895e-05, 3.798479e-05, 1.81028e-05, 1.619271e-05, 1.801281e-05, 
    1.357307e-05, 8.645372e-06, 6.685264e-06, 4.34907e-06, 3.475976e-06,
  1.147816e-05, 1.917309e-05, 2.489706e-05, 2.315261e-05, 3.020949e-05, 
    2.570678e-05, 2.454752e-05, 1.456551e-05, 1.121658e-05, 1.44736e-05, 
    1.764078e-05, 1.524612e-05, 8.505617e-06, 4.86495e-06, 2.685023e-06,
  8.670674e-06, 1.35259e-05, 1.824345e-05, 2.02683e-05, 2.216991e-05, 
    2.570376e-05, 2.125676e-05, 1.499697e-05, 3.63184e-06, 8.663346e-06, 
    1.813621e-05, 1.932859e-05, 1.221384e-05, 6.789165e-06, 2.288173e-06,
  8.572915e-06, 1.35397e-05, 1.932437e-05, 2.183153e-05, 2.198497e-05, 
    1.96532e-05, 2.175673e-05, 1.041424e-05, 2.117773e-06, 4.249642e-06, 
    1.2229e-05, 1.682965e-05, 1.508828e-05, 7.77727e-06, 2.064816e-06,
  6.384933e-06, 7.575529e-06, 9.064763e-06, 1.372657e-05, 1.58603e-05, 
    1.402123e-05, 1.35477e-05, 6.030598e-06, 5.063089e-07, 1.367403e-06, 
    7.968646e-06, 1.318931e-05, 1.324243e-05, 7.464216e-06, 1.803955e-06,
  8.289644e-07, 7.007809e-07, 6.888297e-07, 1.615258e-06, 5.666602e-06, 
    8.036859e-06, 6.879828e-06, 5.436042e-06, 7.580825e-06, 7.099869e-06, 
    6.588001e-06, 1.27537e-05, 1.859074e-05, 1.840098e-05, 1.858907e-05,
  1.616263e-06, 8.272864e-07, 1.814098e-07, 6.34089e-07, 3.42037e-06, 
    3.88218e-06, 7.966351e-06, 8.293431e-06, 6.721066e-06, 6.738658e-06, 
    7.115314e-06, 9.549673e-06, 1.168925e-05, 1.10303e-05, 1.483263e-05,
  5.264164e-06, 1.407364e-06, 1.571957e-06, 6.180837e-07, 2.678555e-06, 
    6.83841e-06, 3.898973e-06, 8.143034e-06, 9.400233e-06, 6.307909e-06, 
    9.64041e-06, 8.25882e-06, 8.784646e-06, 1.113661e-05, 1.20989e-05,
  4.482179e-06, 5.934816e-06, 1.203102e-05, 1.073086e-05, 3.782816e-06, 
    5.235527e-06, 8.451763e-06, 5.188392e-06, 5.922101e-06, 9.711183e-06, 
    9.935281e-06, 8.179031e-06, 8.676204e-06, 1.025675e-05, 8.409771e-06,
  5.189285e-06, 3.133978e-06, 7.934519e-06, 1.394247e-05, 1.68763e-05, 
    1.044989e-05, 7.225355e-06, 3.682685e-06, 7.284091e-06, 9.561639e-06, 
    1.208672e-05, 9.404761e-06, 1.006637e-05, 7.937929e-06, 7.326594e-06,
  6.465806e-06, 1.926752e-06, 6.110867e-06, 1.184229e-05, 2.19456e-05, 
    2.13057e-05, 1.470221e-05, 8.452249e-06, 4.949762e-06, 7.644197e-06, 
    1.045898e-05, 1.16133e-05, 1.130219e-05, 7.859155e-06, 7.039637e-06,
  5.032562e-06, 8.666032e-07, 4.619363e-06, 1.524816e-05, 2.731483e-05, 
    2.73635e-05, 1.790781e-05, 9.307273e-06, 4.098586e-06, 4.397996e-06, 
    9.264057e-06, 1.281051e-05, 1.027744e-05, 7.329088e-06, 5.591999e-06,
  1.543892e-06, 4.406258e-07, 5.446673e-06, 2.549504e-05, 2.699219e-05, 
    2.541678e-05, 2.021176e-05, 1.338456e-05, 3.306794e-06, 1.589081e-06, 
    6.699666e-06, 1.168189e-05, 1.049995e-05, 6.630195e-06, 4.514463e-06,
  4.509641e-08, 1.994129e-06, 2.672062e-05, 2.990481e-05, 2.320801e-05, 
    2.24842e-05, 2.220149e-05, 1.218231e-05, 9.086611e-07, 9.100586e-07, 
    4.877825e-06, 1.257866e-05, 1.07143e-05, 6.391929e-06, 3.92431e-06,
  1.392881e-06, 9.823711e-06, 3.464685e-05, 2.867158e-05, 1.883768e-05, 
    1.836418e-05, 1.791954e-05, 9.746563e-06, 7.073533e-07, 9.153269e-07, 
    4.108676e-06, 1.261236e-05, 1.459621e-05, 6.995367e-06, 3.426071e-06,
  2.220159e-07, 9.962987e-09, 1.078995e-06, 1.702152e-07, 1.624054e-07, 
    4.956371e-06, 9.950752e-06, 9.833201e-06, 1.144849e-05, 1.245333e-05, 
    1.06143e-05, 7.033677e-06, 5.96899e-06, 8.989075e-06, 1.163649e-05,
  1.998692e-07, 5.283034e-07, 2.531892e-07, 6.669298e-08, 8.71907e-07, 
    6.06555e-06, 8.207062e-06, 1.095042e-05, 1.442474e-05, 1.167142e-05, 
    9.168855e-06, 6.515394e-06, 5.329205e-06, 7.341366e-06, 1.052793e-05,
  2.555571e-06, 2.120239e-06, 3.229511e-07, 4.010183e-07, 4.71204e-06, 
    1.915889e-05, 1.430923e-05, 1.639514e-05, 2.075566e-05, 1.350837e-05, 
    5.539191e-06, 3.82291e-06, 4.420071e-06, 6.518093e-06, 9.31973e-06,
  8.872266e-06, 3.014391e-06, 5.691183e-06, 8.124619e-06, 2.19815e-05, 
    4.193878e-05, 6.437553e-05, 3.129306e-05, 2.290476e-05, 1.470651e-05, 
    5.254887e-06, 2.648723e-06, 3.594505e-06, 3.782092e-06, 6.184581e-06,
  8.701762e-06, 2.521491e-06, 1.108294e-05, 2.789657e-05, 3.922057e-05, 
    6.04499e-05, 7.471373e-05, 7.350511e-05, 2.497858e-05, 1.116605e-05, 
    5.247013e-06, 2.459394e-06, 2.937269e-06, 2.937628e-06, 4.181695e-06,
  1.013314e-05, 1.205645e-05, 2.909222e-05, 4.553007e-05, 6.344027e-05, 
    6.634876e-05, 6.02891e-05, 3.286357e-05, 9.586854e-06, 4.772727e-06, 
    3.000034e-06, 2.651104e-06, 3.375197e-06, 4.229985e-06, 4.278144e-06,
  8.53138e-06, 2.453381e-05, 4.030217e-05, 5.719629e-05, 6.132155e-05, 
    5.365003e-05, 3.464637e-05, 1.07376e-05, 8.488998e-06, 6.08112e-06, 
    7.752091e-07, 1.804819e-06, 2.366471e-06, 5.652723e-06, 6.059721e-06,
  9.320142e-06, 3.219198e-05, 5.002724e-05, 7.214243e-05, 5.520819e-05, 
    3.62847e-05, 1.815911e-05, 1.231918e-05, 1.011096e-05, 6.388157e-06, 
    4.899663e-07, 4.549615e-07, 2.435181e-06, 5.608891e-06, 6.049672e-06,
  2.082663e-05, 4.797346e-05, 7.172948e-05, 6.336974e-05, 3.825034e-05, 
    2.483939e-05, 1.618033e-05, 8.405081e-06, 8.989292e-06, 3.723625e-06, 
    3.621409e-07, 4.538068e-07, 2.722681e-06, 5.277758e-06, 6.109025e-06,
  1.259752e-05, 4.447536e-05, 6.461157e-05, 3.842339e-05, 2.99312e-05, 
    1.549117e-05, 1.161401e-05, 5.111019e-06, 7.701544e-06, 3.149441e-06, 
    2.786404e-07, 5.794819e-07, 3.596968e-06, 5.539459e-06, 6.128178e-06,
  9.103151e-09, 3.006169e-08, 3.624728e-07, 2.331765e-06, 1.480528e-05, 
    2.823537e-05, 3.443325e-05, 3.335945e-05, 2.458758e-05, 1.432006e-05, 
    1.383314e-05, 2.436355e-05, 3.888299e-05, 3.647128e-05, 2.484101e-05,
  8.253664e-08, 5.902563e-07, 1.352691e-06, 1.186848e-05, 2.749601e-05, 
    3.389488e-05, 3.529957e-05, 3.02077e-05, 1.836705e-05, 1.251079e-05, 
    1.553272e-05, 3.552154e-05, 4.018565e-05, 2.771713e-05, 1.989628e-05,
  1.825735e-06, 3.662918e-06, 8.6978e-06, 2.784856e-05, 4.640118e-05, 
    4.667748e-05, 1.806248e-05, 9.482486e-06, 1.010845e-05, 1.276471e-05, 
    1.90433e-05, 3.308578e-05, 2.516349e-05, 1.577658e-05, 1.10355e-05,
  6.477885e-06, 9.1332e-06, 2.450744e-05, 3.955951e-05, 3.831352e-05, 
    2.423264e-05, 8.379351e-06, 8.105015e-07, 3.150469e-06, 1.52141e-05, 
    2.217358e-05, 1.346944e-05, 9.664843e-06, 8.505643e-06, 4.023127e-06,
  7.504396e-06, 1.259823e-05, 2.570375e-05, 2.772193e-05, 1.745269e-05, 
    8.337417e-06, 9.013831e-07, 4.565653e-06, 1.223369e-05, 1.217714e-05, 
    1.112661e-05, 3.728944e-06, 3.292245e-06, 6.051499e-06, 3.988021e-06,
  8.311964e-06, 1.208483e-05, 1.478451e-05, 1.250235e-05, 1.339184e-05, 
    1.11384e-05, 1.006156e-05, 5.98938e-06, 7.560522e-06, 4.618983e-06, 
    1.69549e-06, 3.78406e-06, 4.138778e-06, 2.690395e-06, 2.523497e-06,
  1.280033e-05, 1.177401e-05, 8.830548e-06, 9.371782e-06, 1.131046e-05, 
    1.258436e-05, 1.668327e-05, 1.093664e-05, 7.339535e-06, 3.045266e-06, 
    1.301797e-06, 2.035781e-06, 4.396074e-06, 2.428345e-06, 2.178498e-06,
  1.298553e-05, 1.111667e-05, 9.631355e-06, 6.564061e-06, 1.389128e-05, 
    1.250935e-05, 1.93537e-05, 2.165386e-05, 1.476224e-05, 7.023774e-06, 
    1.653341e-06, 1.526268e-06, 2.767335e-07, 1.425867e-06, 1.469566e-06,
  1.244257e-05, 9.312165e-06, 1.042935e-05, 4.072294e-06, 6.966881e-06, 
    1.310316e-05, 2.079944e-05, 2.999415e-05, 2.858485e-05, 1.598845e-05, 
    3.848954e-06, 1.57523e-07, 1.192964e-07, 8.706759e-07, 1.426598e-06,
  4.098054e-06, 1.350621e-06, 3.770014e-06, 2.215678e-06, 4.11388e-06, 
    1.134369e-05, 2.075708e-05, 3.230749e-05, 4.208825e-05, 3.489195e-05, 
    1.112414e-05, 9.351494e-07, 7.192879e-08, 7.441059e-07, 1.386478e-06,
  3.136083e-07, 4.36748e-08, 1.123629e-06, 4.831843e-08, 1.361153e-06, 
    2.511899e-06, 4.617649e-06, 1.772212e-05, 1.70348e-05, 3.321075e-06, 
    1.759764e-06, 3.766545e-06, 8.472547e-06, 9.110274e-06, 1.037367e-05,
  3.610735e-07, 1.978539e-08, 2.049245e-08, 1.184164e-06, 2.504539e-06, 
    1.751202e-06, 5.930091e-06, 2.6387e-05, 2.437749e-05, 4.628578e-06, 
    7.527083e-07, 2.129902e-06, 3.567428e-06, 3.405366e-06, 5.395387e-06,
  1.645386e-06, 3.423919e-08, 1.085683e-06, 3.161858e-06, 3.269787e-06, 
    3.553182e-06, 5.994488e-06, 2.948733e-05, 4.029698e-05, 1.203333e-05, 
    1.166112e-06, 3.533545e-07, 8.537708e-07, 2.786932e-06, 2.850941e-06,
  5.616435e-06, 4.849217e-06, 5.915319e-06, 6.983494e-06, 4.299879e-06, 
    2.54512e-06, 1.350179e-05, 1.319488e-05, 2.359855e-05, 2.761132e-05, 
    3.31081e-06, 1.671996e-06, 1.718781e-07, 6.945857e-07, 1.422378e-06,
  1.103956e-05, 7.938179e-06, 7.403465e-06, 1.047274e-05, 7.778284e-06, 
    4.783901e-06, 9.445932e-06, 4.22807e-05, 7.050742e-05, 4.689557e-05, 
    1.366547e-05, 2.687279e-06, 1.659396e-06, 8.921779e-07, 2.652908e-06,
  9.666919e-06, 6.285429e-06, 5.762002e-06, 7.253442e-06, 1.319805e-05, 
    8.687037e-06, 1.203526e-05, 2.375715e-05, 4.751861e-05, 6.43372e-05, 
    2.992956e-05, 6.29281e-06, 7.363496e-07, 7.719977e-07, 2.652049e-07,
  1.291634e-05, 6.832656e-06, 5.61222e-06, 3.45776e-06, 1.050025e-05, 
    8.80537e-06, 1.258555e-05, 2.282569e-05, 4.602762e-05, 5.408252e-05, 
    4.389939e-05, 1.520232e-05, 2.279292e-06, 1.397257e-07, 1.255042e-08,
  1.125615e-05, 5.042686e-06, 3.83943e-06, 2.499133e-06, 8.268416e-06, 
    2.511463e-06, 6.258192e-06, 9.448077e-06, 2.892392e-05, 4.962902e-05, 
    5.160133e-05, 2.475426e-05, 7.540863e-06, 1.530209e-06, 1.517251e-07,
  9.146428e-06, 4.767401e-06, 6.862194e-06, 3.692609e-06, 2.978913e-06, 
    7.994743e-07, 2.981452e-06, 6.310661e-06, 1.898384e-05, 4.280595e-05, 
    4.735558e-05, 3.007516e-05, 1.342045e-05, 3.608221e-06, 4.000964e-07,
  2.872244e-06, 2.254556e-06, 3.771516e-06, 2.982839e-06, 1.366918e-06, 
    3.91797e-07, 1.348262e-06, 4.737565e-06, 1.139685e-05, 3.785559e-05, 
    4.830309e-05, 3.516272e-05, 1.568882e-05, 6.922751e-06, 1.400895e-06,
  5.43162e-06, 4.53087e-07, 1.829019e-06, 1.511549e-06, 3.310053e-06, 
    3.53077e-06, 3.303739e-06, 2.332888e-06, 1.583588e-06, 5.862355e-07, 
    7.961636e-07, 8.909325e-07, 6.417694e-07, 8.469675e-07, 1.238395e-06,
  1.80418e-06, 7.212079e-07, 2.164482e-06, 8.936128e-07, 2.333845e-06, 
    1.946686e-06, 1.358514e-06, 1.377732e-06, 3.993222e-06, 1.452955e-06, 
    7.794916e-07, 1.671092e-06, 1.459907e-06, 7.060956e-07, 1.180569e-06,
  1.443278e-06, 1.086436e-05, 3.280293e-06, 2.306007e-06, 1.819908e-06, 
    4.98378e-06, 4.589315e-07, 2.046529e-06, 5.113882e-06, 6.311802e-06, 
    2.125727e-06, 8.398129e-07, 7.335757e-07, 2.489921e-06, 1.801225e-06,
  7.377897e-06, 2.100001e-05, 1.156159e-05, 1.003322e-05, 5.270091e-06, 
    2.436779e-06, 2.43077e-06, 2.61154e-06, 3.987415e-06, 1.176777e-05, 
    7.254119e-06, 2.221338e-06, 1.757653e-07, 1.135268e-06, 2.075314e-06,
  1.457415e-05, 1.27813e-05, 1.234659e-05, 1.020064e-05, 9.061151e-06, 
    6.931661e-06, 3.924995e-06, 1.194374e-05, 2.39942e-05, 1.374913e-05, 
    1.440314e-05, 8.983438e-06, 2.177754e-06, 3.872221e-07, 2.223245e-07,
  2.041478e-05, 1.157937e-05, 1.098081e-05, 8.521866e-06, 9.062239e-06, 
    1.076616e-05, 8.23723e-06, 6.603816e-06, 6.967476e-06, 8.030245e-06, 
    1.315227e-05, 1.11308e-05, 6.71714e-06, 2.507977e-06, 1.154066e-06,
  1.115361e-05, 9.157489e-06, 8.648502e-06, 5.935877e-06, 8.922526e-06, 
    1.069046e-05, 1.314843e-05, 9.563917e-06, 8.825115e-06, 7.855914e-06, 
    1.013591e-05, 9.838822e-06, 8.425873e-06, 4.045454e-06, 2.416526e-06,
  1.114412e-05, 7.456606e-06, 5.072513e-06, 2.715633e-06, 6.688608e-06, 
    8.360802e-06, 8.330771e-06, 8.135973e-06, 9.476177e-06, 7.909855e-06, 
    8.22871e-06, 8.239339e-06, 8.001903e-06, 6.539075e-06, 3.7467e-06,
  1.031732e-05, 1.018037e-05, 6.647133e-06, 4.811503e-06, 4.77377e-06, 
    6.781916e-06, 7.6956e-06, 5.693767e-06, 6.990095e-06, 6.439692e-06, 
    5.653622e-06, 6.46086e-06, 6.611536e-06, 6.770356e-06, 6.577907e-06,
  7.481814e-06, 3.257478e-06, 2.313796e-06, 2.045518e-06, 4.253384e-06, 
    5.024192e-06, 5.550867e-06, 3.391972e-06, 3.168517e-06, 3.381658e-06, 
    3.969048e-06, 4.108098e-06, 4.705422e-06, 6.540973e-06, 7.487288e-06,
  5.981321e-06, 6.948021e-07, 1.114121e-06, 2.498622e-07, 4.662008e-07, 
    8.280001e-07, 2.729798e-06, 5.41349e-06, 5.702573e-06, 2.852047e-06, 
    1.691639e-06, 1.467793e-06, 1.203987e-06, 1.228763e-06, 1.639641e-06,
  1.382994e-06, 1.585203e-06, 3.747993e-07, 9.418427e-08, 3.10572e-07, 
    1.347702e-06, 2.19812e-06, 3.396134e-06, 4.000971e-06, 4.98609e-06, 
    1.894154e-06, 2.258894e-06, 2.33891e-06, 2.967754e-06, 2.678454e-06,
  1.302903e-05, 1.084788e-05, 7.540336e-07, 9.474717e-08, 1.681247e-07, 
    1.082542e-06, 9.925232e-07, 2.7118e-06, 4.077122e-06, 4.984808e-06, 
    5.309566e-06, 5.250402e-06, 4.054824e-06, 3.47583e-06, 4.243256e-06,
  1.675573e-05, 1.624859e-05, 1.488246e-05, 7.798611e-06, 7.824999e-07, 
    9.237692e-07, 3.370505e-06, 1.839397e-06, 3.469034e-06, 5.265322e-06, 
    6.732447e-06, 8.57031e-06, 9.418284e-06, 1.005973e-05, 1.065313e-05,
  1.365596e-05, 1.203704e-05, 1.116285e-05, 9.207786e-06, 9.087644e-06, 
    6.904885e-06, 4.313001e-06, 9.165409e-06, 7.223346e-06, 4.96443e-06, 
    1.191711e-05, 1.366836e-05, 1.760404e-05, 2.069319e-05, 2.22523e-05,
  9.861689e-06, 8.005465e-06, 6.863038e-06, 8.413298e-06, 9.607954e-06, 
    5.384192e-06, 6.54395e-06, 8.237545e-06, 1.568175e-05, 2.247923e-05, 
    2.774575e-05, 2.831835e-05, 3.063422e-05, 3.474173e-05, 3.630744e-05,
  5.041693e-06, 7.277337e-06, 9.064072e-06, 6.424777e-06, 6.656059e-06, 
    5.963632e-06, 8.301714e-06, 1.861717e-05, 3.265906e-05, 3.125618e-05, 
    3.212578e-05, 3.524614e-05, 3.910042e-05, 4.064905e-05, 3.595277e-05,
  4.990898e-06, 6.863751e-06, 6.548036e-06, 2.419575e-06, 3.595575e-06, 
    5.325363e-06, 1.017482e-05, 2.039777e-05, 3.044615e-05, 3.622803e-05, 
    3.977385e-05, 4.140881e-05, 4.26409e-05, 4.232711e-05, 3.651512e-05,
  4.283218e-06, 4.290524e-06, 4.678221e-06, 4.790177e-06, 7.79253e-06, 
    1.101172e-05, 1.247264e-05, 1.896155e-05, 3.152972e-05, 3.466142e-05, 
    3.166043e-05, 3.326069e-05, 3.794338e-05, 4.174203e-05, 4.118079e-05,
  2.182552e-06, 4.169981e-06, 8.991585e-06, 1.801752e-05, 2.593175e-05, 
    2.593871e-05, 1.855103e-05, 2.17878e-05, 3.346959e-05, 3.779163e-05, 
    3.76522e-05, 4.085355e-05, 4.615076e-05, 4.913911e-05, 4.655766e-05,
  3.563034e-06, 3.974244e-06, 2.260103e-06, 4.259969e-07, 7.640682e-08, 
    1.222187e-07, 1.365549e-07, 4.636722e-07, 1.165042e-06, 2.805366e-06, 
    5.432577e-06, 1.279287e-05, 2.292187e-05, 2.847344e-05, 3.260748e-05,
  7.277794e-06, 3.852615e-06, 2.801604e-06, 4.368831e-07, 1.117547e-06, 
    1.493607e-07, 8.849337e-08, 2.063577e-07, 7.139902e-07, 2.548505e-06, 
    6.550359e-06, 1.659869e-05, 3.022136e-05, 4.3868e-05, 4.35654e-05,
  7.0109e-06, 6.042768e-06, 4.664692e-06, 1.72401e-06, 2.487013e-06, 
    1.165444e-06, 4.999892e-08, 5.081504e-07, 3.302091e-06, 1.184349e-05, 
    1.725673e-05, 2.173995e-05, 3.164302e-05, 4.004495e-05, 5.42499e-05,
  7.27919e-06, 6.008964e-06, 5.165936e-06, 3.810994e-06, 2.738492e-06, 
    8.317819e-07, 1.728456e-06, 8.911722e-07, 4.294864e-06, 1.51637e-05, 
    2.824302e-05, 2.521682e-05, 2.707565e-05, 3.250225e-05, 4.960516e-05,
  9.662532e-06, 5.882052e-06, 5.387394e-06, 3.930629e-06, 4.635594e-06, 
    3.749562e-06, 9.710576e-07, 8.956865e-06, 5.140247e-06, 7.279932e-06, 
    2.000816e-05, 1.981949e-05, 2.012622e-05, 2.156639e-05, 3.065107e-05,
  2.046303e-05, 9.940803e-06, 5.668974e-06, 3.75678e-06, 3.223375e-06, 
    2.727303e-06, 2.075514e-06, 4.32789e-06, 1.403911e-05, 1.966437e-05, 
    1.663313e-05, 1.298786e-05, 1.158603e-05, 1.249194e-05, 1.703436e-05,
  2.284935e-05, 1.694077e-05, 8.398665e-06, 5.007224e-06, 2.361965e-06, 
    1.786195e-06, 2.507406e-06, 8.233796e-06, 2.054578e-05, 1.239387e-05, 
    4.73454e-06, 3.719329e-06, 3.424817e-06, 4.56272e-06, 6.796795e-06,
  2.067193e-05, 1.537942e-05, 8.00352e-06, 4.590871e-06, 1.69864e-06, 
    1.925428e-06, 5.625437e-06, 1.489116e-05, 1.175363e-05, 5.219465e-06, 
    2.137026e-06, 1.444478e-06, 1.555089e-06, 1.932302e-06, 4.439916e-06,
  1.63178e-05, 1.218995e-05, 7.775515e-06, 4.84931e-06, 3.940135e-06, 
    5.598866e-06, 1.766371e-05, 1.599458e-05, 9.024575e-06, 3.685598e-06, 
    1.970203e-06, 6.753179e-07, 7.333138e-07, 1.502487e-06, 6.254442e-06,
  1.24938e-05, 7.632641e-06, 5.809557e-06, 5.050472e-06, 6.74684e-06, 
    1.659516e-05, 1.952463e-05, 1.184554e-05, 8.905676e-06, 3.159764e-06, 
    2.965948e-06, 3.775429e-07, 6.904727e-07, 3.669631e-06, 1.447341e-05,
  5.33387e-06, 3.71014e-06, 6.078503e-06, 6.3353e-06, 4.491275e-06, 
    3.411763e-06, 2.411645e-06, 8.322525e-07, 3.965886e-07, 3.592548e-07, 
    1.90834e-07, 1.054763e-06, 2.601449e-06, 1.705538e-06, 2.188187e-06,
  8.592951e-06, 6.591795e-06, 6.561503e-06, 6.378342e-06, 5.599831e-06, 
    3.963729e-06, 3.319368e-06, 1.435075e-06, 6.242867e-07, 3.717214e-07, 
    3.677501e-07, 1.402955e-06, 2.043462e-06, 2.624488e-06, 2.513468e-06,
  1.428433e-05, 1.106095e-05, 9.224145e-06, 9.361261e-06, 8.674685e-06, 
    6.363687e-06, 2.428886e-06, 2.439404e-06, 2.016972e-06, 1.344153e-06, 
    1.053694e-06, 2.410805e-06, 2.423831e-06, 2.492203e-06, 3.411199e-06,
  1.737762e-05, 2.127654e-05, 2.247908e-05, 1.895879e-05, 1.82999e-05, 
    8.576911e-06, 8.504107e-06, 2.356872e-06, 7.614999e-07, 5.558351e-07, 
    2.100157e-06, 2.736383e-06, 4.068543e-06, 5.50397e-06, 6.972972e-06,
  1.745599e-05, 2.241989e-05, 2.517188e-05, 2.838702e-05, 2.75827e-05, 
    1.871857e-05, 1.814261e-05, 1.374698e-05, 1.350368e-06, 2.411807e-06, 
    4.831918e-06, 5.032079e-06, 7.769529e-06, 1.049216e-05, 1.292547e-05,
  1.907644e-05, 2.115146e-05, 2.349561e-05, 2.569381e-05, 2.763707e-05, 
    2.579832e-05, 2.46279e-05, 1.248257e-05, 5.389917e-06, 6.909037e-06, 
    1.121319e-05, 1.22035e-05, 1.56414e-05, 1.72352e-05, 1.964158e-05,
  1.992592e-05, 2.638543e-05, 2.541506e-05, 2.153262e-05, 2.066399e-05, 
    1.976275e-05, 1.856636e-05, 1.106818e-05, 4.624759e-06, 5.38172e-06, 
    8.712937e-06, 1.399208e-05, 1.782045e-05, 1.755467e-05, 1.84101e-05,
  1.822978e-05, 2.264945e-05, 2.129475e-05, 1.985566e-05, 1.768897e-05, 
    1.721233e-05, 1.107094e-05, 6.389252e-06, 3.081909e-06, 6.538218e-06, 
    1.14944e-05, 1.705006e-05, 2.02614e-05, 2.116157e-05, 2.271824e-05,
  2.294974e-05, 2.46819e-05, 2.725845e-05, 1.887197e-05, 1.20918e-05, 
    9.106185e-06, 1.134745e-05, 4.318433e-06, 6.244141e-06, 1.356244e-05, 
    1.789402e-05, 2.268352e-05, 2.618843e-05, 2.999685e-05, 3.510633e-05,
  2.196498e-05, 1.726756e-05, 1.396841e-05, 7.395427e-06, 4.798083e-06, 
    2.458852e-06, 3.300554e-06, 5.916845e-06, 1.26568e-05, 2.242422e-05, 
    3.157185e-05, 3.535731e-05, 4.14553e-05, 4.685473e-05, 5.04373e-05,
  2.712642e-06, 2.504274e-06, 3.579719e-06, 5.346666e-06, 7.105124e-06, 
    8.576723e-06, 8.134809e-06, 8.759289e-06, 1.116917e-05, 1.331619e-05, 
    1.28581e-05, 1.48405e-05, 1.191335e-05, 6.145695e-06, 4.09722e-06,
  1.492207e-06, 1.96541e-06, 3.018567e-06, 4.52094e-06, 7.032009e-06, 
    7.037098e-06, 1.237309e-05, 1.021539e-05, 8.271759e-06, 1.272623e-05, 
    1.48874e-05, 1.401423e-05, 1.093774e-05, 6.750673e-06, 5.97998e-06,
  5.817978e-06, 2.025145e-06, 2.900636e-06, 5.839815e-06, 8.246787e-06, 
    1.454343e-05, 1.49512e-05, 2.199853e-05, 1.220297e-05, 7.744551e-06, 
    9.60533e-06, 1.224461e-05, 1.200896e-05, 1.193108e-05, 1.145783e-05,
  5.971286e-06, 1.261621e-05, 1.086802e-05, 9.126166e-06, 1.523385e-05, 
    1.552657e-05, 1.631287e-05, 1.512292e-05, 1.309674e-05, 1.283317e-05, 
    9.393785e-06, 8.222629e-06, 8.918064e-06, 7.838382e-06, 9.697856e-06,
  6.168431e-06, 8.68995e-06, 9.329316e-06, 1.034836e-05, 1.799174e-05, 
    2.010018e-05, 1.93857e-05, 1.924238e-05, 1.004189e-05, 1.829017e-05, 
    1.397069e-05, 6.604368e-06, 5.757168e-06, 4.191476e-06, 5.749197e-06,
  6.25074e-06, 8.111992e-06, 9.470894e-06, 1.213045e-05, 1.734173e-05, 
    1.87572e-05, 2.022345e-05, 1.423963e-05, 7.259486e-06, 9.900919e-06, 
    9.718047e-06, 5.925979e-06, 3.757532e-06, 2.640196e-06, 2.827012e-06,
  1.29298e-05, 1.490355e-05, 1.151165e-05, 1.249911e-05, 1.317221e-05, 
    1.148895e-05, 1.472467e-05, 1.32134e-05, 6.217043e-06, 5.747735e-06, 
    5.408411e-06, 5.409712e-06, 4.030728e-06, 2.490973e-06, 2.341857e-06,
  2.241913e-05, 1.951883e-05, 8.094334e-06, 6.377691e-06, 6.39e-06, 
    1.201066e-05, 1.038766e-05, 9.352418e-06, 4.328457e-06, 6.020576e-06, 
    4.823441e-06, 3.70417e-06, 3.371722e-06, 2.537541e-06, 2.280394e-06,
  2.711447e-05, 1.679235e-05, 1.417654e-05, 4.194528e-06, 5.175074e-06, 
    7.478294e-06, 9.207594e-06, 7.309583e-06, 5.207409e-06, 4.179194e-06, 
    4.411095e-06, 4.102176e-06, 3.678515e-06, 3.171141e-06, 3.401224e-06,
  1.077321e-05, 9.221157e-06, 6.229514e-06, 4.773986e-06, 2.208194e-06, 
    6.647461e-06, 6.14332e-06, 6.804597e-06, 5.360828e-06, 4.266468e-06, 
    8.117017e-06, 8.572208e-06, 8.42255e-06, 7.386209e-06, 5.828303e-06,
  3.840651e-07, 1.765217e-07, 5.016885e-07, 2.158577e-07, 2.755755e-07, 
    2.731399e-06, 5.635671e-06, 4.660318e-06, 4.853614e-06, 5.691588e-06, 
    6.83401e-06, 8.844111e-06, 1.266345e-05, 1.273384e-05, 1.350209e-05,
  2.686668e-07, 1.592988e-07, 4.955518e-07, 6.663742e-07, 7.976369e-07, 
    2.060684e-06, 3.31113e-06, 3.602022e-06, 3.698011e-06, 3.418512e-06, 
    4.942668e-06, 8.145415e-06, 8.706125e-06, 9.244292e-06, 1.189582e-05,
  2.894509e-07, 2.935364e-07, 1.895864e-06, 7.498243e-07, 1.865556e-06, 
    2.549988e-05, 3.410013e-06, 3.109001e-06, 3.578021e-06, 4.211789e-06, 
    3.23098e-06, 5.502576e-06, 7.715413e-06, 1.091668e-05, 1.323828e-05,
  3.591529e-07, 5.297837e-07, 1.743816e-06, 1.097864e-06, 4.781115e-06, 
    1.220283e-05, 3.6594e-05, 3.434049e-06, 2.397522e-06, 3.987534e-06, 
    3.476195e-06, 3.424311e-06, 7.758799e-06, 1.123136e-05, 1.59747e-05,
  3.451283e-08, 3.15816e-07, 1.8288e-06, 3.400241e-06, 8.33154e-06, 
    9.546772e-06, 1.442898e-05, 4.223632e-05, 2.302089e-05, 4.758042e-06, 
    5.617811e-06, 4.937669e-06, 7.627167e-06, 1.040086e-05, 1.329435e-05,
  8.107126e-08, 2.467277e-07, 1.548116e-06, 3.943253e-06, 5.827784e-06, 
    5.83744e-06, 6.236033e-06, 9.81627e-06, 1.037317e-05, 9.782036e-06, 
    9.607021e-06, 6.763169e-06, 8.364426e-06, 1.064783e-05, 1.130418e-05,
  6.320101e-07, 2.675765e-07, 7.242904e-07, 3.348845e-06, 3.138067e-06, 
    4.063263e-06, 7.781719e-06, 1.029891e-05, 1.007911e-05, 1.129834e-05, 
    1.150554e-05, 1.097657e-05, 1.138877e-05, 1.542771e-05, 1.1721e-05,
  6.514675e-07, 1.624939e-06, 1.407355e-06, 1.92435e-06, 2.69985e-06, 
    5.080071e-06, 3.771346e-06, 8.133315e-06, 9.333871e-06, 1.402643e-05, 
    1.742339e-05, 1.710889e-05, 1.516334e-05, 1.157016e-05, 1.104205e-05,
  1.984006e-07, 6.799395e-07, 1.425269e-06, 1.877181e-06, 2.202686e-06, 
    3.050543e-06, 2.840426e-06, 6.70761e-06, 1.315804e-05, 2.090417e-05, 
    2.523594e-05, 2.295158e-05, 1.413607e-05, 1.06767e-05, 1.146895e-05,
  2.967785e-07, 1.349351e-06, 2.500939e-06, 2.536453e-06, 3.580121e-06, 
    5.506372e-06, 6.415374e-06, 1.230625e-05, 2.327991e-05, 3.264334e-05, 
    3.476553e-05, 2.560448e-05, 1.3006e-05, 1.097292e-05, 9.279913e-06,
  5.022125e-07, 4.876343e-07, 1.062837e-06, 4.850242e-07, 3.267139e-07, 
    6.219394e-07, 1.885552e-06, 2.705644e-06, 3.019082e-06, 4.849731e-06, 
    2.75113e-06, 3.043571e-06, 6.725968e-06, 1.435761e-05, 2.517514e-05,
  4.016132e-07, 3.772312e-07, 4.621212e-07, 2.815753e-07, 9.123709e-07, 
    1.148074e-06, 6.598507e-07, 1.378646e-06, 1.961181e-06, 2.452124e-06, 
    2.492878e-06, 4.277445e-06, 1.051829e-05, 2.622551e-05, 4.020839e-05,
  2.264533e-07, 3.874864e-07, 1.598073e-06, 2.23153e-06, 3.297949e-06, 
    9.837577e-06, 1.008509e-06, 6.928692e-07, 1.18603e-06, 3.096911e-06, 
    4.164699e-06, 6.841676e-06, 1.56947e-05, 2.970239e-05, 4.861616e-05,
  1.843367e-07, 4.927851e-07, 2.524438e-07, 2.123757e-07, 1.392009e-06, 
    5.207421e-06, 1.648233e-05, 2.023581e-06, 5.036795e-07, 1.569087e-06, 
    4.786316e-06, 7.453794e-06, 1.568088e-05, 3.30658e-05, 4.551437e-05,
  1.573882e-07, 3.051139e-07, 2.451435e-07, 5.112502e-07, 2.106649e-06, 
    5.548179e-06, 1.140413e-05, 3.838804e-05, 1.852233e-05, 2.186193e-06, 
    5.655804e-06, 1.033994e-05, 2.016591e-05, 3.591408e-05, 3.777352e-05,
  6.613329e-07, 5.819042e-07, 1.482848e-06, 2.337759e-06, 3.771004e-06, 
    5.430515e-06, 1.017163e-05, 1.028141e-05, 7.66242e-06, 8.093003e-06, 
    1.347548e-05, 1.802318e-05, 3.031482e-05, 3.590551e-05, 3.865415e-05,
  2.487742e-06, 3.956594e-06, 6.075561e-06, 3.650489e-06, 4.406945e-06, 
    5.727687e-06, 7.746574e-06, 9.19652e-06, 8.902977e-06, 9.618183e-06, 
    1.315907e-05, 1.992603e-05, 3.243521e-05, 3.91902e-05, 4.234448e-05,
  6.481514e-06, 9.834132e-06, 4.447188e-06, 2.8288e-06, 3.838249e-06, 
    5.740615e-06, 6.856819e-06, 7.655614e-06, 7.824059e-06, 7.942662e-06, 
    1.030448e-05, 2.000276e-05, 3.929298e-05, 4.290049e-05, 3.689745e-05,
  8.48614e-06, 4.971517e-06, 5.817016e-06, 4.623883e-06, 3.728993e-06, 
    4.990351e-06, 6.634426e-06, 7.468645e-06, 9.18925e-06, 8.314199e-06, 
    1.070243e-05, 2.366803e-05, 4.164073e-05, 3.686777e-05, 2.134641e-05,
  2.574814e-06, 5.173451e-06, 5.039382e-06, 5.391473e-06, 4.323024e-06, 
    3.787897e-06, 4.361867e-06, 5.852812e-06, 8.783e-06, 1.084559e-05, 
    1.60847e-05, 3.2495e-05, 3.777056e-05, 2.067564e-05, 7.316914e-06,
  2.21388e-07, 2.541748e-07, 2.37368e-07, 2.059799e-07, 2.62354e-07, 
    4.811828e-07, 8.85836e-07, 2.31068e-06, 4.563209e-06, 7.720011e-06, 
    9.047901e-06, 8.855822e-06, 1.345618e-05, 1.299247e-05, 1.213876e-05,
  3.60802e-07, 3.790773e-07, 2.690031e-07, 2.421861e-07, 1.457086e-06, 
    3.034585e-06, 1.66721e-06, 3.539144e-06, 4.926539e-06, 5.479312e-06, 
    6.67131e-06, 6.41728e-06, 8.483119e-06, 1.988072e-05, 1.771877e-05,
  5.496339e-07, 9.799041e-07, 8.564597e-07, 2.066082e-06, 3.765361e-06, 
    1.065513e-05, 2.8121e-06, 2.829704e-06, 5.110999e-06, 5.725082e-06, 
    3.513081e-06, 2.257312e-06, 5.048377e-06, 1.319488e-05, 2.323947e-05,
  4.370918e-06, 5.893289e-06, 8.869832e-06, 9.257677e-06, 3.220494e-06, 
    3.778436e-06, 1.67778e-05, 4.611047e-06, 1.68679e-06, 1.959426e-06, 
    3.156106e-06, 3.547464e-06, 8.928056e-06, 1.465905e-05, 2.542795e-05,
  6.804135e-06, 1.052275e-05, 1.111852e-05, 1.327433e-05, 1.725229e-05, 
    1.280708e-05, 7.161326e-06, 3.596271e-05, 2.190336e-05, 3.14309e-06, 
    6.999227e-06, 9.306063e-06, 1.170886e-05, 1.513894e-05, 2.207549e-05,
  5.50231e-06, 1.045981e-05, 1.357653e-05, 1.495061e-05, 1.89088e-05, 
    1.605894e-05, 1.515364e-05, 9.228651e-06, 9.438689e-06, 1.184062e-05, 
    1.510001e-05, 1.238953e-05, 1.382647e-05, 1.658368e-05, 2.261197e-05,
  9.769252e-06, 1.51503e-05, 1.540138e-05, 1.187947e-05, 1.372791e-05, 
    1.190106e-05, 1.361532e-05, 1.216061e-05, 1.057867e-05, 1.051357e-05, 
    1.16565e-05, 1.21783e-05, 1.328576e-05, 1.71514e-05, 2.228936e-05,
  1.329461e-05, 1.516577e-05, 1.263922e-05, 6.788394e-06, 5.2654e-06, 
    8.044203e-06, 1.032769e-05, 9.858147e-06, 9.342401e-06, 1.164043e-05, 
    1.339007e-05, 1.193345e-05, 1.360508e-05, 2.016733e-05, 2.529125e-05,
  2.075547e-05, 1.368477e-05, 1.300195e-05, 8.597317e-06, 9.277812e-06, 
    1.029244e-05, 1.234626e-05, 1.277916e-05, 1.318694e-05, 1.43206e-05, 
    1.144037e-05, 1.204444e-05, 1.608627e-05, 2.284793e-05, 3.579233e-05,
  2.858484e-05, 2.508447e-05, 2.388624e-05, 1.989809e-05, 1.565431e-05, 
    1.30195e-05, 1.151986e-05, 1.083856e-05, 1.07139e-05, 9.165125e-06, 
    9.106899e-06, 9.815093e-06, 1.638264e-05, 3.135344e-05, 4.371831e-05,
  3.99376e-08, 6.108696e-08, 1.24767e-07, 1.756948e-07, 2.116063e-07, 
    2.778291e-07, 4.132345e-07, 7.247399e-07, 1.661385e-06, 3.685432e-06, 
    5.111272e-06, 5.59421e-06, 9.200289e-06, 1.142072e-05, 1.081102e-05,
  5.389086e-07, 7.139918e-07, 9.445865e-07, 1.105934e-06, 1.213961e-06, 
    1.33079e-06, 1.52204e-06, 1.964904e-06, 2.68348e-06, 4.100815e-06, 
    5.658878e-06, 8.469759e-06, 1.074279e-05, 1.724444e-05, 1.239649e-05,
  1.680995e-06, 1.786492e-06, 1.766143e-06, 1.922582e-06, 2.346866e-06, 
    4.482462e-06, 1.97239e-06, 2.518579e-06, 4.530018e-06, 4.662596e-06, 
    4.070663e-06, 4.585329e-06, 7.493186e-06, 9.390167e-06, 1.254977e-05,
  6.112529e-06, 3.962197e-06, 2.725314e-06, 2.928829e-06, 4.418564e-06, 
    5.742394e-06, 9.227163e-06, 3.337674e-06, 1.993071e-06, 5.089389e-06, 
    6.707646e-06, 4.41081e-06, 5.776598e-06, 8.42971e-06, 1.275858e-05,
  2.145859e-05, 1.987347e-05, 2.134094e-05, 2.621114e-05, 3.762413e-05, 
    2.840435e-05, 2.03073e-05, 2.183995e-05, 1.891009e-05, 8.452536e-06, 
    1.544321e-05, 6.134293e-06, 4.858897e-06, 7.783591e-06, 1.359895e-05,
  2.964655e-05, 3.541809e-05, 3.598825e-05, 3.848875e-05, 3.669945e-05, 
    2.969666e-05, 2.967243e-05, 1.557203e-05, 3.756122e-06, 8.021007e-06, 
    1.506153e-05, 9.244418e-06, 7.643915e-06, 8.359727e-06, 1.132218e-05,
  3.552568e-05, 3.247815e-05, 2.854158e-05, 2.766014e-05, 2.317514e-05, 
    1.736047e-05, 2.048677e-05, 2.125581e-05, 8.941094e-06, 7.351142e-06, 
    8.729132e-06, 1.060648e-05, 1.117123e-05, 9.978974e-06, 9.468687e-06,
  3.28032e-05, 2.763646e-05, 2.791094e-05, 1.973728e-05, 1.681809e-05, 
    1.697302e-05, 8.756057e-06, 6.221011e-06, 2.567554e-06, 3.755209e-06, 
    7.790414e-06, 9.515114e-06, 9.072823e-06, 9.437438e-06, 9.732744e-06,
  4.737316e-05, 4.430607e-05, 4.050917e-05, 3.308164e-05, 2.907871e-05, 
    2.438668e-05, 2.047354e-05, 1.573738e-05, 1.176487e-05, 8.524093e-06, 
    5.665393e-06, 6.783766e-06, 1.040341e-05, 1.264823e-05, 1.457223e-05,
  4.288847e-05, 4.057396e-05, 3.738966e-05, 3.376731e-05, 3.523496e-05, 
    3.98864e-05, 4.364654e-05, 4.364772e-05, 3.561191e-05, 2.446151e-05, 
    1.421363e-05, 1.345277e-05, 1.821972e-05, 1.938287e-05, 1.807407e-05,
  3.076706e-07, 2.613732e-06, 3.738907e-07, 5.518625e-07, 8.919779e-07, 
    8.532185e-07, 6.771242e-07, 3.589223e-07, 2.635633e-07, 3.283233e-07, 
    1.415088e-07, 1.625562e-07, 2.872985e-07, 4.43296e-07, 7.537236e-07,
  5.843681e-06, 2.202196e-06, 1.539816e-07, 4.317191e-07, 1.138872e-06, 
    7.595706e-07, 1.325699e-06, 4.447053e-07, 4.587274e-07, 3.14851e-07, 
    2.657289e-07, 2.095146e-07, 3.802615e-07, 1.012443e-06, 1.183865e-06,
  1.700381e-05, 7.431627e-06, 4.641727e-06, 1.699834e-06, 2.24362e-06, 
    1.292367e-06, 1.735072e-07, 2.752202e-07, 5.795746e-07, 3.394312e-07, 
    2.268833e-07, 2.750318e-07, 6.152689e-07, 1.916537e-06, 4.580392e-06,
  4.135493e-05, 2.763361e-05, 1.908494e-05, 1.50719e-05, 5.833544e-06, 
    4.843499e-06, 3.582637e-06, 7.285391e-07, 4.169605e-07, 2.424181e-07, 
    1.505892e-06, 2.143077e-06, 2.58146e-06, 5.447389e-06, 1.021302e-05,
  4.162294e-05, 4.122565e-05, 4.720215e-05, 5.318121e-05, 4.943652e-05, 
    2.736783e-05, 1.761099e-05, 1.661221e-05, 5.350209e-06, 1.069006e-06, 
    6.249666e-06, 3.207416e-06, 1.788335e-06, 4.528611e-06, 8.724636e-06,
  2.069525e-05, 2.141578e-05, 2.519459e-05, 2.918135e-05, 3.827305e-05, 
    4.901372e-05, 5.302395e-05, 3.04258e-05, 8.193886e-06, 1.175344e-05, 
    9.240052e-06, 4.096635e-06, 3.586321e-06, 6.115865e-06, 8.081334e-06,
  1.982664e-05, 1.484911e-05, 9.78657e-06, 7.012738e-06, 9.27594e-06, 
    1.122249e-05, 1.988496e-05, 2.365506e-05, 1.40003e-05, 4.531436e-06, 
    4.425793e-06, 5.581861e-06, 7.691438e-06, 1.002105e-05, 1.138633e-05,
  3.459427e-05, 2.651498e-05, 1.938177e-05, 1.472673e-05, 1.335445e-05, 
    1.638307e-05, 1.359567e-05, 8.856251e-06, 9.369944e-06, 2.293032e-06, 
    5.623784e-06, 6.515153e-06, 6.556168e-06, 8.134001e-06, 1.013577e-05,
  3.163177e-05, 3.230822e-05, 3.087076e-05, 2.633795e-05, 2.158091e-05, 
    1.886013e-05, 1.456324e-05, 9.130246e-06, 9.81886e-06, 7.003363e-06, 
    7.687046e-06, 6.725973e-06, 9.728024e-06, 1.139985e-05, 1.247789e-05,
  3.136e-05, 2.937903e-05, 3.246044e-05, 2.763657e-05, 1.926949e-05, 
    1.239243e-05, 6.120215e-06, 4.077523e-06, 1.190619e-05, 1.82357e-05, 
    2.476963e-05, 2.462787e-05, 2.735809e-05, 2.853524e-05, 3.22389e-05,
  5.580314e-06, 1.018319e-05, 7.312902e-06, 9.036933e-06, 4.877723e-06, 
    4.928887e-06, 4.444114e-06, 1.85424e-06, 2.919305e-06, 3.636683e-06, 
    2.567854e-06, 2.709181e-06, 4.30108e-06, 3.729281e-06, 3.125452e-06,
  1.172744e-05, 6.493171e-06, 1.845406e-06, 3.349855e-06, 5.955961e-06, 
    3.238957e-06, 1.359465e-05, 1.422912e-06, 2.194432e-06, 2.783975e-06, 
    2.589696e-06, 3.49795e-06, 5.111611e-06, 4.558991e-06, 2.089199e-06,
  1.337203e-05, 1.366415e-05, 2.262834e-05, 2.13572e-05, 1.852256e-05, 
    9.036547e-06, 4.951658e-06, 6.633722e-06, 4.057227e-06, 2.982903e-06, 
    2.450635e-06, 2.583969e-06, 3.818737e-06, 3.074518e-06, 3.332567e-06,
  2.837044e-05, 3.190703e-05, 2.907468e-05, 2.300585e-05, 2.262209e-05, 
    1.923715e-05, 1.467136e-05, 7.423662e-06, 6.4601e-06, 8.900789e-07, 
    2.895024e-06, 3.399142e-06, 4.14448e-06, 5.248791e-06, 7.409958e-06,
  1.634134e-05, 1.31304e-05, 1.716735e-05, 2.549909e-05, 3.586694e-05, 
    2.118099e-05, 3.100502e-05, 2.290093e-05, 4.95527e-06, 2.844263e-06, 
    4.959097e-06, 3.541711e-06, 3.290022e-06, 3.790158e-06, 4.477632e-06,
  2.036548e-05, 1.276506e-05, 1.223558e-05, 1.975603e-05, 2.012873e-05, 
    2.508864e-05, 4.426536e-05, 3.061244e-05, 1.559266e-05, 1.424377e-05, 
    6.149046e-06, 6.070788e-06, 1.021462e-05, 1.148559e-05, 1.497694e-05,
  2.495079e-05, 2.230756e-05, 1.560898e-05, 1.060681e-05, 9.505251e-06, 
    1.2751e-05, 1.806529e-05, 2.104975e-05, 1.848365e-05, 4.46252e-06, 
    1.972397e-06, 4.495121e-06, 4.959329e-06, 5.418674e-06, 7.151718e-06,
  2.329841e-05, 2.342032e-05, 1.956859e-05, 1.781234e-05, 1.406216e-05, 
    1.391065e-05, 1.1883e-05, 1.086926e-05, 6.435097e-06, 9.800109e-07, 
    8.820581e-07, 1.035522e-06, 4.378936e-07, 7.435826e-07, 8.217403e-07,
  2.186119e-05, 2.118791e-05, 2.111896e-05, 1.958266e-05, 1.90615e-05, 
    1.580654e-05, 1.096367e-05, 1.050553e-05, 8.701548e-06, 6.781045e-06, 
    1.143064e-05, 1.056245e-06, 5.512788e-07, 5.998613e-07, 1.311605e-06,
  1.676279e-05, 1.624359e-05, 1.581949e-05, 1.39396e-05, 1.46959e-05, 
    1.052609e-05, 5.941972e-06, 4.162531e-06, 3.865061e-06, 4.216454e-06, 
    8.568078e-06, 5.004872e-06, 3.07095e-06, 3.183286e-06, 6.583835e-06,
  3.568265e-06, 6.630577e-06, 6.300366e-06, 1.046613e-05, 5.064956e-06, 
    5.595305e-06, 8.997989e-06, 3.458402e-06, 7.031003e-06, 7.212685e-06, 
    4.814411e-06, 7.363697e-06, 1.17497e-05, 1.152628e-05, 6.951102e-06,
  7.751715e-06, 7.542379e-06, 4.008501e-06, 2.975512e-06, 4.202318e-06, 
    6.782427e-06, 1.334895e-05, 2.972282e-06, 4.543936e-06, 6.3944e-06, 
    7.244479e-06, 1.252587e-05, 1.421664e-05, 9.533675e-06, 5.433914e-06,
  2.802572e-05, 9.888328e-06, 1.273364e-05, 1.575854e-05, 1.793148e-05, 
    9.606872e-06, 7.524045e-06, 1.941877e-05, 1.104683e-05, 7.010698e-06, 
    5.704051e-06, 8.957979e-06, 1.244694e-05, 1.137125e-05, 1.367022e-05,
  4.383597e-05, 4.56715e-05, 3.561965e-05, 3.536737e-05, 1.39903e-05, 
    1.939846e-05, 1.141623e-05, 1.128625e-05, 9.847271e-06, 2.256627e-06, 
    7.15223e-06, 9.838568e-06, 1.198142e-05, 1.967145e-05, 2.462064e-05,
  3.260334e-05, 2.238513e-05, 2.429815e-05, 2.529522e-05, 3.270152e-05, 
    1.06272e-05, 2.862905e-05, 3.18705e-05, 1.157491e-05, 1.30079e-06, 
    5.283827e-06, 6.42504e-06, 9.594321e-06, 1.591751e-05, 2.066633e-05,
  3.043081e-05, 2.689e-05, 2.722449e-05, 2.167959e-05, 1.827173e-05, 
    2.559198e-05, 3.230468e-05, 1.313118e-05, 8.478103e-06, 8.221421e-06, 
    7.055124e-06, 5.727885e-06, 9.762592e-06, 1.2987e-05, 1.499764e-05,
  3.061816e-05, 3.234331e-05, 3.05859e-05, 2.230706e-05, 1.864404e-05, 
    1.771286e-05, 1.97111e-05, 2.270607e-05, 1.340603e-05, 3.839635e-06, 
    2.938917e-06, 6.152762e-06, 1.064091e-05, 1.00263e-05, 9.926863e-06,
  3.332934e-05, 3.403701e-05, 3.407001e-05, 2.516096e-05, 2.441115e-05, 
    2.238048e-05, 1.873613e-05, 1.417917e-05, 6.550285e-06, 1.649805e-06, 
    1.736823e-06, 3.536629e-06, 4.251148e-06, 5.783532e-06, 6.249614e-06,
  3.227837e-05, 3.725358e-05, 3.869264e-05, 2.79078e-05, 2.241462e-05, 
    1.829851e-05, 1.662803e-05, 1.204544e-05, 6.14469e-06, 4.231255e-06, 
    6.094985e-06, 8.955165e-07, 1.5159e-06, 2.833894e-06, 3.271397e-06,
  2.112007e-05, 2.359346e-05, 2.909814e-05, 2.067833e-05, 1.456658e-05, 
    1.105219e-05, 7.087957e-06, 6.149265e-06, 5.882649e-06, 2.731406e-06, 
    6.061031e-06, 1.459681e-06, 1.338535e-06, 1.762714e-06, 2.083945e-06,
  1.21951e-05, 9.970094e-06, 1.125878e-05, 1.184364e-05, 4.685462e-06, 
    3.788193e-06, 8.37284e-06, 4.16701e-06, 4.617024e-06, 4.84069e-06, 
    3.826625e-06, 4.614615e-06, 5.763905e-06, 5.605177e-06, 4.565331e-06,
  9.652812e-06, 8.546115e-06, 8.810194e-06, 5.950043e-06, 4.717644e-06, 
    1.251134e-05, 1.323813e-05, 4.309903e-06, 2.892195e-06, 4.270714e-06, 
    4.889191e-06, 7.435454e-06, 7.027097e-06, 4.727892e-06, 4.007893e-06,
  2.526126e-05, 1.585629e-05, 1.771357e-05, 1.827459e-05, 1.610512e-05, 
    1.187675e-05, 4.743673e-06, 4.355838e-06, 2.261469e-06, 1.921934e-06, 
    3.270646e-06, 4.148853e-06, 5.121152e-06, 5.260849e-06, 8.515711e-06,
  2.406459e-05, 2.65559e-05, 3.182537e-05, 3.792911e-05, 3.1349e-05, 
    2.333542e-05, 2.603485e-05, 1.314301e-05, 2.058494e-06, 1.123669e-06, 
    2.423764e-06, 2.962452e-06, 3.346505e-06, 7.968379e-06, 1.160736e-05,
  1.924642e-05, 1.70644e-05, 2.16656e-05, 2.835803e-05, 4.33171e-05, 
    4.941746e-05, 5.24043e-05, 3.963527e-05, 1.563851e-05, 1.239445e-06, 
    5.389544e-06, 6.048129e-06, 2.793023e-06, 6.203823e-06, 9.404684e-06,
  2.520214e-05, 2.006432e-05, 1.657294e-05, 1.860112e-05, 2.992947e-05, 
    4.383936e-05, 5.666413e-05, 3.670377e-05, 1.845244e-05, 1.767719e-05, 
    7.825043e-06, 1.83897e-06, 3.563865e-06, 6.652613e-06, 8.737001e-06,
  2.723043e-05, 2.222284e-05, 1.333214e-05, 1.654583e-05, 1.96775e-05, 
    2.516105e-05, 3.552268e-05, 3.812843e-05, 3.213017e-05, 2.3934e-05, 
    1.341293e-05, 7.783088e-06, 6.309546e-06, 6.573769e-06, 7.548867e-06,
  1.831582e-05, 1.740827e-05, 1.462403e-05, 1.749837e-05, 1.833015e-05, 
    2.109617e-05, 1.600808e-05, 1.264986e-05, 4.365928e-06, 6.331158e-06, 
    1.51338e-05, 1.996994e-05, 1.399775e-05, 9.099787e-06, 7.28193e-06,
  1.536406e-05, 1.52274e-05, 1.708686e-05, 1.760757e-05, 1.73991e-05, 
    1.565182e-05, 1.341209e-05, 9.53629e-06, 4.569225e-06, 5.008696e-06, 
    6.44103e-06, 1.069577e-05, 1.240378e-05, 1.080577e-05, 7.960326e-06,
  2.934844e-05, 1.214242e-05, 1.43362e-05, 1.38436e-05, 1.123007e-05, 
    7.831944e-06, 5.253338e-06, 4.262636e-06, 4.454429e-06, 2.51918e-06, 
    2.066276e-06, 2.05112e-06, 4.501399e-06, 4.78894e-06, 5.36687e-06,
  1.726794e-05, 1.361447e-05, 8.810215e-06, 1.044078e-05, 7.563349e-06, 
    7.10169e-06, 5.457326e-06, 1.890182e-06, 2.833369e-06, 3.794354e-06, 
    3.641313e-06, 4.715539e-06, 4.99275e-06, 3.987637e-06, 3.070571e-06,
  3.478982e-05, 2.470152e-05, 1.322908e-05, 1.389166e-05, 1.528264e-05, 
    1.173802e-05, 8.906609e-06, 2.960178e-06, 3.142663e-06, 2.926072e-06, 
    4.644201e-06, 8.433564e-06, 6.864108e-06, 4.554705e-06, 3.244765e-06,
  3.882687e-05, 4.185108e-05, 3.248525e-05, 1.947543e-05, 1.712518e-05, 
    1.559787e-05, 9.634991e-06, 1.044612e-05, 8.006269e-06, 4.555801e-06, 
    4.725719e-06, 7.906272e-06, 7.234786e-06, 6.985223e-06, 7.364358e-06,
  4.595118e-05, 3.361172e-05, 2.290675e-05, 1.436894e-05, 1.007407e-05, 
    1.014397e-05, 1.879811e-05, 1.985595e-05, 1.394851e-05, 6.580628e-06, 
    6.270385e-06, 5.936372e-06, 6.732026e-06, 9.949935e-06, 1.127233e-05,
  4.15718e-05, 2.311572e-05, 5.537352e-06, 9.5007e-06, 1.505661e-05, 
    1.82387e-05, 1.306498e-05, 2.096061e-05, 1.114009e-05, 1.202148e-05, 
    1.328105e-05, 6.163222e-06, 5.961147e-06, 8.617349e-06, 1.038881e-05,
  3.701841e-05, 1.1285e-05, 1.029344e-06, 4.521829e-06, 1.429976e-05, 
    2.738965e-05, 3.159625e-05, 8.215036e-06, 7.079916e-06, 1.019738e-05, 
    8.069128e-06, 6.814507e-06, 6.334636e-06, 6.777739e-06, 9.510956e-06,
  3.501832e-05, 1.387928e-05, 4.785323e-06, 5.265224e-06, 1.223272e-05, 
    2.206524e-05, 2.957881e-05, 1.999864e-05, 3.974304e-06, 2.425425e-06, 
    4.12338e-06, 7.019328e-06, 7.602669e-06, 5.751854e-06, 7.079163e-06,
  8.669456e-05, 4.286025e-05, 1.369377e-05, 1.771688e-05, 2.793329e-05, 
    3.184427e-05, 2.192597e-05, 1.022785e-05, 2.282846e-06, 8.393633e-07, 
    5.993393e-07, 5.779737e-06, 8.232157e-06, 7.628558e-06, 7.318808e-06,
  0.000113129, 4.351574e-05, 2.235454e-05, 2.63927e-05, 3.264225e-05, 
    3.303308e-05, 2.453807e-05, 1.307554e-05, 2.594948e-06, 3.948196e-06, 
    2.727197e-06, 3.420046e-06, 9.03857e-06, 1.035308e-05, 8.527365e-06,
  4.058194e-05, 2.552566e-05, 2.032095e-05, 1.891474e-05, 1.432643e-05, 
    7.280537e-06, 6.440712e-06, 3.937231e-06, 2.82073e-06, 1.370105e-06, 
    1.84626e-06, 1.998196e-06, 8.804999e-06, 1.473813e-05, 1.398986e-05,
  3.046773e-05, 2.912692e-05, 2.437296e-05, 1.756803e-05, 1.271595e-05, 
    8.504755e-06, 7.574607e-06, 2.325484e-06, 2.663611e-06, 4.124756e-06, 
    2.330102e-06, 1.876508e-06, 2.795973e-06, 3.623851e-06, 5.305765e-06,
  1.831821e-05, 2.629041e-05, 2.219061e-05, 1.92172e-05, 1.899452e-05, 
    1.667046e-05, 1.287764e-05, 4.232314e-06, 3.403675e-06, 4.141798e-06, 
    5.131345e-06, 5.53012e-06, 3.08906e-06, 2.642438e-06, 3.305082e-06,
  2.780463e-05, 2.895119e-05, 2.678732e-05, 1.521256e-05, 1.496814e-05, 
    1.177697e-05, 1.411966e-05, 1.511249e-05, 1.089622e-05, 5.540082e-06, 
    6.59057e-06, 5.936362e-06, 4.053482e-06, 2.197938e-06, 2.445336e-06,
  4.921764e-05, 4.463702e-05, 3.785638e-05, 2.750148e-05, 1.538866e-05, 
    8.75058e-06, 1.185755e-05, 1.656792e-05, 1.043704e-05, 7.144717e-06, 
    7.594652e-06, 5.704402e-06, 5.260397e-06, 4.420908e-06, 4.366958e-06,
  6.131966e-05, 4.369192e-05, 3.245121e-05, 3.229139e-05, 2.308422e-05, 
    2.09415e-05, 1.016442e-05, 1.212206e-05, 8.401584e-06, 3.101882e-06, 
    9.50899e-06, 7.485654e-06, 6.91255e-06, 5.277844e-06, 4.601406e-06,
  4.531816e-05, 2.441487e-05, 2.429748e-05, 2.103072e-05, 1.983637e-05, 
    1.738043e-05, 2.163481e-05, 6.235668e-06, 2.417768e-06, 5.346315e-06, 
    5.698912e-06, 6.134522e-06, 8.135667e-06, 7.142005e-06, 5.951656e-06,
  3.038153e-05, 2.341926e-05, 2.35487e-05, 2.248992e-05, 1.535363e-05, 
    1.313138e-05, 2.322866e-05, 1.965932e-05, 4.420694e-06, 3.128412e-06, 
    1.691039e-06, 2.61893e-06, 5.40754e-06, 6.747217e-06, 7.006117e-06,
  8.139233e-05, 5.205841e-05, 3.260065e-05, 2.100719e-05, 1.879807e-05, 
    1.970261e-05, 2.945697e-05, 2.606462e-05, 3.929483e-06, 2.485749e-06, 
    2.054518e-06, 2.024634e-06, 2.16405e-06, 2.200837e-06, 3.924537e-06,
  0.00011925, 6.398658e-05, 2.798241e-05, 1.287008e-05, 1.312123e-05, 
    1.170019e-05, 2.277989e-05, 4.029545e-05, 2.531429e-05, 1.124401e-05, 
    3.484107e-06, 1.340461e-06, 7.92075e-07, 6.104147e-07, 1.125018e-06,
  4.299207e-05, 2.44804e-05, 1.134082e-05, 1.055109e-05, 7.69019e-06, 
    6.664029e-06, 1.590584e-05, 3.742243e-05, 4.134321e-05, 3.078369e-05, 
    1.051989e-05, 1.872592e-06, 3.042517e-07, 1.550502e-07, 7.026804e-07,
  5.866977e-06, 1.277197e-05, 1.533523e-05, 2.13543e-05, 2.750404e-05, 
    2.723825e-05, 2.058691e-05, 9.562445e-06, 4.190881e-06, 3.258809e-06, 
    2.776021e-06, 2.167914e-06, 2.521228e-06, 3.483304e-06, 7.59003e-06,
  2.980862e-06, 8.574632e-06, 1.570768e-05, 2.011897e-05, 2.838331e-05, 
    2.641607e-05, 2.302622e-05, 1.752528e-05, 1.218343e-05, 7.843484e-06, 
    3.632969e-06, 3.0143e-06, 1.403333e-06, 1.969694e-06, 5.502703e-06,
  7.817965e-06, 1.622334e-05, 1.806938e-05, 1.8772e-05, 1.646416e-05, 
    2.174721e-05, 2.206231e-05, 2.685835e-05, 2.254885e-05, 1.492209e-05, 
    8.372655e-06, 4.984683e-06, 1.773048e-06, 1.241375e-06, 3.80689e-06,
  2.852659e-05, 4.591803e-05, 4.387434e-05, 3.106477e-05, 1.866039e-05, 
    1.072678e-05, 2.214375e-05, 2.619059e-05, 2.243646e-05, 1.561975e-05, 
    9.43168e-06, 4.469458e-06, 1.822034e-06, 1.971888e-06, 2.293457e-06,
  5.841381e-05, 5.591639e-05, 4.575165e-05, 4.012682e-05, 3.701903e-05, 
    2.429189e-05, 1.261101e-05, 1.218129e-05, 1.096423e-05, 5.699339e-06, 
    5.203757e-06, 2.036133e-06, 2.457349e-06, 2.480267e-06, 1.726099e-06,
  5.420929e-05, 3.486199e-05, 3.504971e-05, 3.706834e-05, 3.890053e-05, 
    4.002617e-05, 2.595053e-05, 1.308529e-05, 6.449236e-06, 6.458316e-06, 
    2.176598e-06, 6.405665e-07, 2.163675e-06, 2.712383e-06, 1.659625e-06,
  5.301091e-05, 4.639283e-05, 4.101628e-05, 3.592556e-05, 3.315708e-05, 
    3.041739e-05, 2.606589e-05, 2.501202e-05, 1.286612e-05, 6.751879e-06, 
    1.16366e-06, 1.825293e-06, 2.80293e-06, 2.301924e-06, 2.141325e-06,
  5.66676e-05, 5.240634e-05, 3.862749e-05, 3.077725e-05, 2.431395e-05, 
    2.113943e-05, 1.454954e-05, 1.161517e-05, 4.043912e-06, 5.459186e-06, 
    6.508935e-06, 5.612314e-06, 4.141719e-06, 2.646005e-06, 2.889871e-06,
  4.524839e-05, 4.334838e-05, 4.029241e-05, 2.503583e-05, 1.319617e-05, 
    9.985339e-06, 8.282725e-06, 6.596882e-06, 2.203941e-06, 1.461652e-06, 
    6.132853e-06, 6.399839e-06, 4.91572e-06, 3.161143e-06, 3.102548e-06,
  2.784846e-05, 3.037666e-05, 2.264767e-05, 9.578094e-06, 5.639591e-06, 
    5.065674e-06, 5.116042e-06, 5.307032e-06, 3.96382e-06, 1.708347e-06, 
    3.605384e-06, 5.667682e-06, 5.832377e-06, 4.63118e-06, 3.296218e-06,
  2.230954e-06, 1.983851e-06, 1.596967e-06, 2.740012e-06, 2.219149e-06, 
    3.148536e-06, 2.838648e-06, 1.95312e-06, 9.155815e-07, 1.142656e-06, 
    1.505601e-06, 2.254616e-06, 3.159747e-06, 3.933077e-06, 4.392729e-06,
  6.21698e-06, 4.596799e-06, 4.306203e-06, 5.32448e-06, 7.893709e-06, 
    9.228653e-06, 5.412831e-06, 3.363365e-06, 2.312606e-06, 2.565033e-06, 
    2.650913e-06, 4.188122e-06, 5.367323e-06, 3.009484e-06, 3.385014e-06,
  9.013596e-06, 1.101226e-05, 9.725253e-06, 5.79372e-06, 8.494966e-06, 
    8.905677e-06, 9.340602e-06, 1.333732e-05, 1.132949e-05, 7.664496e-06, 
    4.941177e-06, 3.800862e-06, 3.178838e-06, 3.380311e-06, 5.173967e-06,
  4.462645e-05, 3.132409e-05, 3.628789e-05, 1.916722e-05, 8.976848e-06, 
    7.819944e-06, 1.29105e-05, 1.654806e-05, 1.476682e-05, 1.065049e-05, 
    7.750008e-06, 5.698814e-06, 6.29551e-06, 6.359821e-06, 6.33533e-06,
  5.111007e-05, 4.415593e-05, 5.169122e-05, 3.965834e-05, 3.188848e-05, 
    2.62369e-05, 1.535698e-05, 1.957085e-05, 1.65549e-05, 5.247752e-06, 
    1.026705e-05, 6.570717e-06, 7.496072e-06, 5.937809e-06, 4.126695e-06,
  4.875611e-05, 4.45322e-05, 5.613244e-05, 5.976858e-05, 6.805267e-05, 
    5.648512e-05, 3.931066e-05, 1.485137e-05, 8.362393e-06, 1.198181e-05, 
    1.086596e-05, 7.009657e-06, 8.645434e-06, 6.092421e-06, 5.29909e-06,
  4.274205e-05, 4.292443e-05, 3.763827e-05, 4.30545e-05, 4.677424e-05, 
    4.495781e-05, 3.937364e-05, 3.565418e-05, 2.325311e-05, 1.891167e-05, 
    1.293882e-05, 1.099899e-05, 9.318615e-06, 6.023538e-06, 4.75241e-06,
  2.807795e-05, 4.152516e-05, 4.00004e-05, 2.845212e-05, 2.524388e-05, 
    2.270116e-05, 1.87504e-05, 2.018739e-05, 1.757079e-05, 1.553735e-05, 
    1.78159e-05, 1.699364e-05, 1.229666e-05, 7.573897e-06, 4.579656e-06,
  2.075901e-05, 3.869065e-05, 4.221686e-05, 3.098447e-05, 1.320565e-05, 
    8.497696e-06, 8.051783e-06, 1.197878e-05, 1.755895e-05, 2.044306e-05, 
    2.322222e-05, 2.033427e-05, 1.537949e-05, 9.877311e-06, 4.338161e-06,
  1.249722e-05, 2.019136e-05, 2.442008e-05, 1.107827e-05, 4.771007e-06, 
    4.632812e-06, 4.529563e-06, 5.523545e-06, 1.271892e-05, 1.610969e-05, 
    2.175384e-05, 2.222773e-05, 1.639341e-05, 9.063961e-06, 3.498764e-06,
  3.668737e-06, 2.530715e-06, 2.364348e-06, 2.329917e-06, 1.041667e-05, 
    1.315888e-05, 1.78967e-05, 1.757368e-05, 1.687441e-05, 1.429895e-05, 
    1.52618e-05, 1.815478e-05, 1.645375e-05, 1.223125e-05, 1.15655e-05,
  7.097921e-06, 1.248767e-06, 2.462885e-06, 1.234573e-06, 8.119626e-06, 
    1.181808e-05, 2.053951e-05, 1.677395e-05, 1.425449e-05, 1.849218e-05, 
    1.340823e-05, 1.650496e-05, 1.333907e-05, 7.825968e-06, 3.329933e-06,
  4.211209e-05, 1.257918e-05, 1.83991e-06, 5.708673e-07, 3.942881e-06, 
    5.273338e-06, 1.503314e-05, 2.293698e-05, 2.229204e-05, 2.116296e-05, 
    2.237862e-05, 1.804723e-05, 1.925104e-05, 1.092496e-05, 3.364416e-06,
  4.100969e-05, 6.011146e-05, 2.503239e-05, 1.154352e-05, 2.313172e-06, 
    5.562143e-06, 7.450498e-06, 1.475149e-05, 2.280428e-05, 2.724973e-05, 
    2.067518e-05, 1.768206e-05, 2.045225e-05, 1.449821e-05, 5.485299e-06,
  2.717459e-05, 5.165634e-05, 6.136546e-05, 2.732684e-05, 1.638057e-05, 
    9.1419e-06, 6.817955e-06, 1.794765e-06, 8.551877e-06, 1.901353e-05, 
    1.925894e-05, 1.441428e-05, 1.280955e-05, 8.750286e-06, 3.97168e-06,
  1.645563e-05, 4.377124e-05, 6.541172e-05, 4.869594e-05, 3.458444e-05, 
    2.518062e-05, 2.164878e-05, 9.649612e-06, 6.589878e-06, 1.350003e-05, 
    1.40746e-05, 1.319749e-05, 8.036625e-06, 3.357041e-06, 2.242428e-06,
  2.700808e-05, 3.65748e-05, 4.703565e-05, 5.303884e-05, 4.924081e-05, 
    3.712191e-05, 2.267826e-05, 2.029523e-05, 1.442872e-05, 1.339805e-05, 
    1.362252e-05, 1.105495e-05, 5.712034e-06, 2.791634e-06, 2.48068e-06,
  4.250103e-05, 4.41885e-05, 3.808317e-05, 3.98594e-05, 3.44157e-05, 
    3.407906e-05, 2.079693e-05, 1.242265e-05, 8.726824e-06, 9.749434e-06, 
    1.052638e-05, 1.024219e-05, 4.813386e-06, 3.45351e-06, 4.175528e-06,
  4.897351e-05, 4.943293e-05, 4.238148e-05, 2.255443e-05, 1.383106e-05, 
    1.257154e-05, 1.090441e-05, 7.778933e-06, 6.981464e-06, 8.010765e-06, 
    7.877193e-06, 6.886567e-06, 4.953535e-06, 6.03862e-06, 6.966564e-06,
  3.274261e-05, 3.534878e-05, 2.382463e-05, 8.920401e-06, 3.870369e-06, 
    3.469729e-06, 4.418179e-06, 6.301088e-06, 6.843102e-06, 6.618459e-06, 
    6.614979e-06, 5.976761e-06, 6.766949e-06, 9.750543e-06, 1.015241e-05,
  2.838422e-07, 2.339664e-06, 3.770786e-06, 1.211539e-05, 2.664841e-05, 
    3.936296e-05, 3.492589e-05, 2.132201e-05, 1.767775e-05, 1.040291e-05, 
    5.103002e-06, 3.3895e-06, 4.373248e-06, 4.592567e-06, 4.33749e-06,
  3.630637e-06, 1.099585e-06, 5.037138e-06, 1.363636e-05, 2.794571e-05, 
    3.492305e-05, 2.679159e-05, 1.664249e-05, 1.208505e-05, 9.479327e-06, 
    3.634144e-06, 5.759815e-06, 3.630088e-06, 2.71721e-06, 3.590481e-06,
  3.819317e-05, 1.56581e-05, 6.456773e-06, 1.297056e-05, 1.985779e-05, 
    1.205459e-05, 1.249748e-05, 1.506318e-05, 1.222107e-05, 8.713091e-06, 
    7.570491e-06, 2.548877e-06, 2.633127e-06, 4.164306e-06, 7.241117e-06,
  4.215604e-05, 5.867104e-05, 4.859871e-05, 2.111079e-05, 1.704838e-05, 
    1.013673e-05, 3.720763e-06, 7.595226e-06, 1.31221e-05, 1.08317e-05, 
    4.622508e-06, 2.653502e-06, 4.980557e-06, 9.705665e-06, 1.286862e-05,
  4.985067e-05, 5.874125e-05, 4.715277e-05, 2.915205e-05, 2.282018e-05, 
    1.78065e-05, 7.377109e-06, 1.013058e-06, 6.100913e-06, 6.53108e-06, 
    4.769706e-06, 5.742393e-06, 6.862619e-06, 7.464476e-06, 1.129112e-05,
  5.913063e-05, 5.685071e-05, 6.094461e-05, 4.285351e-05, 2.732052e-05, 
    2.45806e-05, 1.891126e-05, 5.910363e-06, 2.867641e-06, 9.109681e-06, 
    4.983144e-06, 5.621534e-06, 6.133954e-06, 5.259737e-06, 6.197562e-06,
  6.498343e-05, 6.375746e-05, 5.882223e-05, 4.882981e-05, 4.351318e-05, 
    3.460089e-05, 2.380343e-05, 2.173621e-05, 1.677662e-05, 1.611231e-05, 
    1.217132e-05, 6.104934e-06, 4.256038e-06, 3.864657e-06, 4.077563e-06,
  6.061849e-05, 5.83397e-05, 5.19253e-05, 3.96357e-05, 4.261967e-05, 
    3.593651e-05, 2.970032e-05, 2.215832e-05, 9.681215e-06, 7.725078e-06, 
    9.14928e-06, 6.974675e-06, 4.024774e-06, 2.623807e-06, 1.793547e-06,
  5.212054e-05, 4.839282e-05, 3.844353e-05, 2.842766e-05, 2.241937e-05, 
    2.347956e-05, 2.183919e-05, 1.756183e-05, 1.329128e-05, 1.257055e-05, 
    1.21063e-05, 7.659367e-06, 2.795538e-06, 1.365089e-06, 1.209071e-06,
  2.468251e-05, 1.552409e-05, 1.453626e-05, 1.145001e-05, 1.238339e-05, 
    1.144473e-05, 1.289017e-05, 1.655876e-05, 1.671345e-05, 1.161657e-05, 
    1.112834e-05, 6.342078e-06, 2.297309e-06, 8.388911e-07, 8.596539e-07,
  1.507717e-05, 2.21523e-05, 2.184138e-05, 1.617219e-05, 1.527377e-05, 
    2.615277e-05, 3.239099e-05, 9.393028e-06, 5.632238e-06, 4.47815e-06, 
    9.629677e-06, 1.460721e-05, 1.276595e-05, 1.06459e-05, 6.326707e-06,
  2.451115e-05, 1.10562e-05, 9.463226e-06, 4.538835e-06, 3.050313e-06, 
    2.220774e-05, 4.304878e-05, 1.602754e-05, 2.760082e-06, 7.98937e-06, 
    5.198445e-06, 9.113991e-06, 6.743033e-06, 3.701446e-06, 3.210432e-06,
  4.733371e-05, 1.742376e-05, 7.448386e-06, 3.2636e-06, 2.869447e-06, 
    1.620339e-05, 3.611185e-05, 2.580496e-05, 9.387883e-06, 8.36147e-06, 
    3.604346e-06, 2.418909e-06, 4.368642e-06, 2.312845e-06, 1.912495e-06,
  5.326469e-05, 5.056736e-05, 3.846442e-05, 2.265826e-05, 9.977407e-06, 
    6.248177e-06, 1.885965e-05, 2.168439e-05, 1.821114e-05, 7.73488e-06, 
    2.851864e-06, 6.620654e-07, 2.685503e-06, 2.984616e-06, 3.208592e-06,
  5.550749e-05, 5.289581e-05, 4.268056e-05, 3.637037e-05, 2.937465e-05, 
    1.530157e-05, 2.603641e-06, 4.923012e-06, 1.131974e-05, 4.516426e-06, 
    2.1913e-06, 1.901321e-06, 3.422036e-06, 4.369498e-06, 3.332323e-06,
  5.808794e-05, 5.151614e-05, 4.587306e-05, 4.175426e-05, 3.886547e-05, 
    2.921758e-05, 7.546519e-06, 4.827109e-07, 1.435964e-06, 5.344197e-06, 
    3.883355e-06, 5.548676e-06, 3.704225e-06, 3.37028e-06, 3.378772e-06,
  6.413024e-05, 5.80821e-05, 5.037379e-05, 4.213331e-05, 3.820646e-05, 
    3.44857e-05, 2.365046e-05, 1.115417e-05, 5.242963e-06, 9.307096e-06, 
    5.236863e-06, 4.746805e-06, 3.241744e-06, 2.128623e-06, 5.349939e-06,
  6.624966e-05, 5.632803e-05, 4.584897e-05, 3.632365e-05, 3.624291e-05, 
    2.793498e-05, 2.053448e-05, 1.389285e-05, 1.867077e-06, 1.920125e-06, 
    3.949694e-06, 2.118148e-06, 2.696506e-06, 5.447984e-06, 7.45973e-06,
  3.200039e-05, 3.980783e-05, 3.768355e-05, 2.587813e-05, 1.457905e-05, 
    1.50246e-05, 1.127121e-05, 5.598314e-06, 1.778315e-06, 7.897085e-07, 
    1.793589e-06, 3.383428e-06, 6.12664e-06, 6.188542e-06, 4.860869e-06,
  9.571145e-06, 1.595594e-05, 1.702411e-05, 9.682951e-06, 2.84143e-06, 
    1.869138e-06, 2.1484e-06, 5.929905e-06, 3.247972e-06, 1.232803e-06, 
    2.064168e-06, 3.155228e-06, 4.013461e-06, 2.266824e-06, 1.275988e-06,
  1.90656e-06, 2.003751e-06, 1.018725e-06, 2.239429e-06, 1.451484e-06, 
    3.360807e-06, 8.148457e-06, 1.06938e-05, 4.189583e-06, 4.392552e-07, 
    1.920342e-06, 9.405805e-06, 1.079723e-05, 1.440727e-05, 2.117596e-05,
  9.904272e-06, 2.990836e-06, 1.010896e-06, 1.758977e-06, 5.391896e-06, 
    1.22032e-05, 1.826765e-05, 6.96155e-06, 9.829089e-07, 4.515972e-06, 
    6.557453e-06, 1.792756e-05, 1.987769e-05, 1.571243e-05, 1.703798e-05,
  3.413814e-05, 2.227202e-05, 1.417289e-05, 9.903154e-06, 7.322018e-06, 
    1.020702e-05, 8.733945e-06, 5.772662e-06, 3.111963e-06, 6.050629e-06, 
    1.040681e-05, 1.544972e-05, 2.056474e-05, 1.873644e-05, 1.493008e-05,
  5.845852e-05, 5.14165e-05, 3.352e-05, 2.427579e-05, 1.225598e-05, 
    4.447661e-06, 1.68545e-06, 6.93972e-07, 2.359366e-06, 3.610582e-06, 
    4.617766e-06, 1.005777e-05, 1.699121e-05, 1.778356e-05, 1.655892e-05,
  4.330989e-05, 3.993617e-05, 3.237615e-05, 2.447751e-05, 1.525494e-05, 
    9.187738e-06, 1.218849e-06, 6.438558e-07, 5.909857e-06, 2.077677e-06, 
    3.465787e-06, 7.570029e-06, 1.323985e-05, 1.35977e-05, 1.540051e-05,
  3.179314e-05, 3.38469e-05, 2.824724e-05, 2.150578e-05, 1.868318e-05, 
    1.376341e-05, 7.531445e-06, 3.202227e-06, 1.600003e-06, 9.334111e-06, 
    5.585906e-06, 8.526404e-06, 1.181795e-05, 1.114888e-05, 1.044481e-05,
  2.592294e-05, 2.612079e-05, 2.824623e-05, 2.575485e-05, 2.740987e-05, 
    2.394927e-05, 1.58033e-05, 6.906374e-06, 8.779075e-06, 9.166852e-06, 
    5.299576e-06, 8.980387e-06, 1.132549e-05, 1.089766e-05, 8.183588e-06,
  2.110494e-05, 2.226965e-05, 2.039804e-05, 2.044957e-05, 2.485173e-05, 
    2.345119e-05, 1.78211e-05, 9.977897e-06, 3.889463e-06, 2.120466e-06, 
    1.837756e-06, 4.491058e-06, 6.702468e-06, 9.675072e-06, 9.637094e-06,
  1.723015e-05, 1.922536e-05, 1.782725e-05, 1.737745e-05, 1.128621e-05, 
    1.042554e-05, 1.109574e-05, 3.842024e-06, 8.45639e-07, 6.880022e-07, 
    9.732947e-07, 1.37004e-06, 2.772825e-06, 4.308197e-06, 5.946879e-06,
  1.37263e-05, 1.201134e-05, 8.593532e-06, 5.817982e-06, 3.61721e-06, 
    1.668001e-06, 1.942727e-06, 2.739657e-06, 7.245622e-07, 1.118227e-06, 
    1.433126e-06, 1.687574e-06, 1.922017e-06, 2.686681e-06, 3.417105e-06,
  3.665684e-06, 4.333014e-06, 2.300186e-06, 1.791015e-06, 3.071311e-06, 
    2.787089e-06, 4.904712e-06, 6.914939e-06, 8.894489e-06, 1.672865e-05, 
    3.212727e-05, 4.073312e-05, 3.531041e-05, 2.140876e-05, 8.780714e-06,
  1.103639e-05, 5.803375e-06, 3.823584e-06, 3.506689e-06, 3.525496e-06, 
    2.050121e-06, 2.339445e-06, 2.807609e-06, 5.558122e-06, 1.132388e-05, 
    2.022625e-05, 3.120803e-05, 2.300856e-05, 1.669272e-05, 1.008139e-05,
  1.790405e-05, 9.705592e-06, 8.270405e-06, 2.955152e-06, 2.378204e-06, 
    8.885028e-07, 1.355124e-06, 1.101332e-06, 1.157746e-06, 5.356306e-06, 
    1.060792e-05, 1.72096e-05, 1.731927e-05, 1.335079e-05, 9.006916e-06,
  3.668553e-05, 2.867011e-05, 2.103992e-05, 1.330965e-05, 6.356652e-06, 
    1.415214e-06, 1.289539e-06, 1.282677e-07, 2.474274e-07, 1.79604e-06, 
    4.852363e-06, 8.267999e-06, 1.058319e-05, 9.43846e-06, 6.454365e-06,
  2.199734e-05, 2.303494e-05, 2.114234e-05, 1.645375e-05, 8.761335e-06, 
    8.439891e-06, 4.617186e-06, 1.450117e-06, 3.851993e-06, 8.390465e-07, 
    2.993364e-06, 3.02965e-06, 6.423608e-06, 5.240972e-06, 5.229163e-06,
  1.498516e-05, 1.462722e-05, 1.517373e-05, 1.610392e-05, 1.409507e-05, 
    1.123191e-05, 6.637371e-06, 7.987488e-06, 2.81249e-06, 5.261258e-06, 
    1.232199e-06, 2.353818e-06, 2.817409e-06, 4.353649e-06, 3.768565e-06,
  1.265065e-05, 1.204526e-05, 1.131511e-05, 1.197692e-05, 1.50874e-05, 
    1.43468e-05, 1.191919e-05, 8.814197e-06, 5.475826e-06, 4.818284e-06, 
    2.417963e-06, 3.546363e-06, 3.049285e-06, 2.841323e-06, 3.632918e-06,
  1.040995e-05, 1.144951e-05, 9.238341e-06, 9.449583e-06, 1.179027e-05, 
    1.638896e-05, 1.064452e-05, 7.73827e-06, 1.705226e-06, 1.729792e-06, 
    1.982712e-06, 3.217423e-06, 4.030181e-06, 3.649394e-06, 3.968859e-06,
  9.206597e-06, 1.007361e-05, 1.28317e-05, 1.172311e-05, 6.649374e-06, 
    5.030916e-06, 5.661207e-06, 1.593846e-06, 1.311626e-06, 1.779431e-06, 
    1.404293e-06, 2.503524e-06, 4.846328e-06, 4.891397e-06, 5.668162e-06,
  8.762277e-06, 7.273047e-06, 2.962308e-06, 1.487943e-06, 1.596883e-06, 
    1.883632e-08, 5.962014e-08, 1.290789e-08, 1.64862e-06, 1.903686e-06, 
    1.088639e-06, 1.360305e-06, 3.179612e-06, 5.663256e-06, 6.405639e-06,
  1.151508e-06, 3.640921e-06, 2.037256e-06, 2.336164e-06, 4.992077e-06, 
    3.068752e-06, 5.945686e-06, 7.240499e-06, 2.080856e-05, 2.520629e-05, 
    2.372311e-05, 1.75379e-05, 1.287238e-05, 6.023639e-06, 2.847979e-06,
  2.90139e-06, 1.698479e-06, 2.11424e-06, 2.462057e-06, 1.245741e-06, 
    9.889171e-07, 3.616352e-06, 5.573621e-06, 1.500533e-05, 2.94589e-05, 
    2.423169e-05, 2.240959e-05, 1.515749e-05, 1.6252e-06, 1.654695e-06,
  1.482794e-05, 4.286951e-06, 3.304678e-06, 9.21513e-07, 6.763691e-08, 
    1.506791e-06, 1.237068e-06, 8.940148e-06, 1.852768e-05, 3.569293e-05, 
    2.567393e-05, 2.262839e-05, 1.436363e-05, 9.55047e-07, 5.441113e-07,
  1.601696e-05, 1.426253e-05, 1.236541e-05, 8.107813e-06, 3.733251e-07, 
    1.601662e-06, 1.841193e-06, 2.60516e-06, 7.607234e-06, 2.280499e-05, 
    2.559853e-05, 2.019985e-05, 1.089847e-05, 2.27083e-06, 8.426193e-07,
  1.151882e-05, 5.375689e-06, 6.773046e-06, 8.761472e-06, 5.302788e-06, 
    5.739016e-06, 3.198443e-06, 1.618633e-06, 1.156353e-05, 2.02772e-05, 
    2.370845e-05, 1.735132e-05, 8.649565e-06, 1.470302e-06, 2.71688e-06,
  1.941927e-05, 1.207827e-05, 1.233359e-05, 9.996123e-06, 1.096167e-05, 
    8.947633e-06, 7.215014e-06, 1.079195e-05, 1.920172e-05, 2.337904e-05, 
    1.72624e-05, 1.361703e-05, 6.800018e-06, 1.764848e-06, 1.207859e-06,
  2.692647e-05, 2.738044e-05, 2.344705e-05, 2.413862e-05, 1.917783e-05, 
    9.705392e-06, 9.431326e-06, 1.035796e-05, 1.412705e-05, 1.534571e-05, 
    1.369122e-05, 1.033256e-05, 6.48945e-06, 3.003239e-06, 1.082695e-06,
  2.069416e-05, 2.4089e-05, 2.533751e-05, 2.145389e-05, 1.393524e-05, 
    8.276269e-06, 4.972043e-06, 6.276777e-06, 6.874454e-06, 9.724362e-06, 
    1.008496e-05, 8.258463e-06, 5.874098e-06, 3.851778e-06, 2.461019e-06,
  1.744002e-05, 2.204204e-05, 1.94373e-05, 7.925743e-06, 6.076847e-06, 
    9.228289e-07, 1.007529e-06, 1.333074e-06, 3.913332e-06, 6.861683e-06, 
    6.557375e-06, 5.664885e-06, 4.668766e-06, 3.177769e-06, 3.14949e-06,
  2.043505e-05, 1.995807e-05, 1.685773e-05, 2.874379e-06, 5.098785e-07, 
    6.486128e-08, 2.535454e-08, 4.489933e-07, 1.407638e-06, 2.973362e-06, 
    2.917719e-06, 3.186633e-06, 2.579466e-06, 2.26088e-06, 2.200894e-06,
  3.467455e-06, 2.335257e-06, 3.378676e-06, 2.084284e-06, 3.852399e-06, 
    3.094285e-06, 7.881607e-06, 1.17976e-05, 1.436697e-05, 6.674846e-06, 
    1.379967e-06, 1.699604e-06, 6.531374e-06, 7.166725e-06, 6.274015e-06,
  6.744394e-06, 3.126057e-06, 1.931918e-06, 1.970646e-06, 6.970665e-07, 
    6.772717e-06, 1.866693e-05, 1.87696e-05, 1.26186e-05, 7.815188e-06, 
    4.155255e-06, 3.380988e-06, 4.955246e-06, 5.034762e-06, 5.588744e-06,
  2.000204e-05, 4.789829e-06, 1.61335e-06, 8.871928e-07, 1.08216e-05, 
    3.220479e-05, 2.679425e-05, 2.442425e-05, 1.187514e-05, 8.739311e-06, 
    7.052502e-06, 5.61387e-06, 4.724897e-06, 5.062506e-06, 5.866867e-06,
  3.033933e-05, 1.884449e-05, 1.348785e-05, 1.931524e-05, 3.798205e-05, 
    3.239881e-05, 1.361536e-05, 1.176557e-05, 1.052202e-05, 7.16431e-06, 
    7.52138e-06, 3.125202e-06, 3.472075e-06, 4.382749e-06, 7.49537e-06,
  1.651476e-05, 8.767088e-06, 2.293867e-05, 3.704724e-05, 3.816115e-05, 
    1.557928e-05, 6.46728e-06, 1.001512e-06, 5.18665e-06, 7.001535e-06, 
    4.011131e-06, 2.087812e-06, 2.207265e-06, 2.727512e-06, 7.054235e-06,
  1.87999e-05, 1.637729e-05, 2.223204e-05, 4.913741e-05, 3.88448e-05, 
    1.373545e-05, 9.647176e-06, 8.662489e-06, 8.004344e-06, 4.899833e-06, 
    3.260084e-06, 1.84632e-06, 2.614888e-06, 3.740084e-06, 4.007768e-06,
  2.436882e-05, 1.897019e-05, 3.674007e-05, 4.847477e-05, 3.361295e-05, 
    2.353213e-05, 2.218938e-05, 1.664195e-05, 1.010837e-05, 3.376206e-06, 
    2.29119e-06, 1.748214e-06, 2.387848e-06, 3.692248e-06, 2.406113e-06,
  2.453719e-05, 2.940593e-05, 4.350132e-05, 3.274206e-05, 2.665585e-05, 
    2.530854e-05, 2.210118e-05, 1.355742e-05, 4.567381e-06, 2.59913e-06, 
    2.109627e-06, 2.443178e-06, 2.67146e-06, 3.8536e-06, 3.447851e-06,
  2.433486e-05, 3.350383e-05, 3.195435e-05, 1.179191e-05, 1.083527e-05, 
    1.245766e-05, 1.210979e-05, 5.194849e-06, 3.815383e-06, 2.222991e-06, 
    2.357536e-06, 2.579578e-06, 3.427128e-06, 3.342354e-06, 4.688454e-06,
  2.047907e-05, 2.239933e-05, 1.026245e-05, 4.615849e-06, 5.130528e-06, 
    1.948617e-06, 2.113593e-06, 3.802673e-06, 2.716995e-06, 2.046297e-06, 
    2.315752e-06, 2.082608e-06, 2.111224e-06, 2.423505e-06, 2.400981e-06,
  4.691558e-05, 4.307595e-05, 3.081175e-05, 1.751258e-05, 7.125682e-06, 
    3.614528e-06, 2.651105e-06, 1.267748e-06, 4.228614e-06, 8.231788e-06, 
    8.506322e-06, 8.277048e-06, 1.025133e-05, 1.154524e-05, 1.282026e-05,
  1.756733e-05, 2.033837e-05, 2.599692e-05, 1.999283e-05, 1.23518e-05, 
    5.655928e-06, 2.894732e-06, 4.560548e-06, 8.947231e-06, 1.425795e-05, 
    1.362041e-05, 1.09703e-05, 1.11978e-05, 8.014487e-06, 8.817999e-06,
  1.664507e-05, 9.970067e-06, 1.516947e-05, 1.5178e-05, 1.066515e-05, 
    9.602027e-06, 4.606859e-06, 9.43961e-06, 1.040925e-05, 1.097501e-05, 
    8.69361e-06, 4.461168e-06, 6.306677e-06, 7.254322e-06, 6.584558e-06,
  1.132625e-05, 1.406776e-05, 1.898201e-05, 2.138339e-05, 2.093038e-05, 
    1.098832e-05, 8.977063e-06, 1.114078e-05, 9.647515e-06, 7.294685e-06, 
    2.235081e-06, 1.020009e-06, 4.88368e-06, 5.622652e-06, 5.927773e-06,
  3.1199e-05, 2.809352e-05, 3.063928e-05, 3.093912e-05, 1.756831e-05, 
    8.284223e-06, 5.262346e-06, 4.060782e-06, 7.514525e-06, 2.93576e-06, 
    1.478275e-06, 2.568445e-06, 6.161961e-06, 5.664024e-06, 5.521984e-06,
  4.855455e-05, 4.085842e-05, 3.669698e-05, 3.499665e-05, 2.243068e-05, 
    1.434656e-05, 8.527553e-06, 1.740008e-06, 1.21626e-06, 1.729256e-06, 
    1.697496e-06, 4.724089e-06, 6.091983e-06, 5.356354e-06, 3.906921e-06,
  5.22822e-05, 5.410182e-05, 4.765428e-05, 4.384309e-05, 4.146797e-05, 
    3.434117e-05, 2.30982e-05, 1.24186e-05, 2.982549e-06, 1.330453e-06, 
    4.005004e-06, 4.973072e-06, 4.065983e-06, 3.219603e-06, 1.695328e-06,
  6.350696e-05, 6.299395e-05, 5.824623e-05, 4.982144e-05, 4.912876e-05, 
    4.564021e-05, 1.582497e-05, 1.151509e-05, 1.281836e-06, 2.036919e-06, 
    3.297089e-06, 2.840163e-06, 1.508986e-06, 1.030022e-06, 1.113692e-06,
  7.275477e-05, 6.347682e-05, 5.02268e-05, 3.430249e-05, 2.208066e-05, 
    1.976398e-05, 1.360307e-05, 6.934708e-06, 9.263194e-07, 3.024388e-06, 
    1.918586e-06, 3.165858e-06, 1.7024e-06, 1.51851e-06, 1.586679e-06,
  3.752568e-05, 2.574893e-05, 1.140874e-05, 1.023914e-05, 7.441503e-06, 
    2.663153e-07, 4.028789e-07, 8.191711e-06, 1.192964e-06, 3.268748e-06, 
    2.450213e-06, 1.993654e-06, 2.23649e-06, 2.004477e-06, 1.686122e-06,
  8.933483e-06, 2.509235e-05, 2.781023e-05, 1.689653e-05, 4.706574e-06, 
    1.168286e-06, 1.136177e-06, 8.12252e-07, 6.836239e-07, 4.842211e-07, 
    2.078872e-07, 1.108474e-07, 3.93784e-07, 8.211426e-07, 1.788685e-06,
  7.860543e-06, 1.070956e-05, 2.368824e-05, 2.387819e-05, 1.281845e-05, 
    5.35522e-06, 2.521991e-06, 1.908965e-06, 1.521961e-06, 1.023817e-06, 
    7.325286e-07, 1.211554e-06, 2.386985e-06, 3.339147e-06, 3.838054e-06,
  1.651113e-05, 1.290652e-05, 1.564565e-05, 2.392114e-05, 1.636488e-05, 
    7.290098e-06, 3.879988e-06, 3.294011e-06, 2.375798e-06, 1.513146e-06, 
    1.431852e-06, 2.191663e-06, 5.237232e-06, 7.285252e-06, 8.930862e-06,
  2.317319e-05, 2.500118e-05, 3.11281e-05, 3.300421e-05, 2.330489e-05, 
    6.751255e-06, 5.011928e-06, 3.495034e-06, 2.066569e-06, 1.348494e-06, 
    1.274789e-06, 1.147899e-06, 4.845491e-06, 8.987171e-06, 1.05092e-05,
  3.412975e-05, 3.821254e-05, 5.123162e-05, 3.243583e-05, 2.187504e-05, 
    9.549216e-06, 2.609435e-06, 1.841557e-06, 1.347821e-06, 5.94664e-07, 
    1.05779e-06, 1.072344e-06, 4.364434e-06, 6.331518e-06, 5.757581e-06,
  4.544576e-05, 4.792206e-05, 4.84852e-05, 3.693768e-05, 2.238588e-05, 
    1.303645e-05, 2.925339e-06, 2.108539e-07, 5.27258e-08, 1.922233e-06, 
    8.238027e-07, 1.919228e-06, 3.308294e-06, 3.150513e-06, 3.661055e-06,
  4.896145e-05, 5.367171e-05, 4.274222e-05, 3.600477e-05, 2.98923e-05, 
    1.711189e-05, 8.79493e-06, 4.745412e-06, 2.085059e-06, 1.015055e-06, 
    1.284331e-06, 1.578117e-06, 1.820827e-06, 1.907049e-06, 2.053116e-06,
  5.825617e-05, 5.113159e-05, 4.482604e-05, 4.08915e-05, 3.783337e-05, 
    2.538212e-05, 1.18247e-05, 4.845545e-06, 1.383314e-06, 9.874818e-07, 
    6.476076e-07, 7.417222e-07, 7.252219e-07, 7.542839e-07, 1.157977e-06,
  5.157898e-05, 5.910188e-05, 4.393524e-05, 2.612343e-05, 1.926116e-05, 
    1.601563e-05, 7.362559e-06, 2.967481e-06, 9.800765e-07, 2.920236e-07, 
    5.515444e-07, 6.130683e-07, 5.605029e-07, 5.447444e-07, 3.016456e-07,
  2.719991e-05, 2.185773e-05, 9.702884e-06, 3.410054e-06, 5.963408e-07, 
    1.493662e-06, 1.733193e-07, 1.840566e-06, 7.575222e-07, 4.089921e-07, 
    9.855005e-07, 9.685486e-07, 7.348568e-07, 6.633277e-07, 3.277092e-07,
  2.278139e-06, 6.299737e-06, 1.029713e-05, 1.324107e-05, 1.357707e-05, 
    1.306913e-05, 1.263794e-05, 7.307987e-06, 1.931318e-06, 6.401115e-07, 
    3.295868e-07, 2.213435e-07, 4.396371e-07, 4.731679e-07, 1.07344e-06,
  2.489017e-06, 3.275365e-06, 9.148525e-06, 1.467306e-05, 1.561249e-05, 
    1.172481e-05, 1.245315e-05, 5.897631e-06, 7.50609e-07, 3.335174e-07, 
    4.458052e-07, 7.213084e-07, 5.935049e-07, 1.324982e-06, 2.669978e-06,
  1.317355e-05, 7.975004e-06, 9.71626e-06, 1.694802e-05, 1.235794e-05, 
    4.868827e-06, 7.007438e-06, 3.301629e-06, 7.390067e-07, 3.470305e-07, 
    6.817282e-07, 6.739552e-07, 1.120015e-06, 2.620539e-06, 5.209028e-06,
  3.542606e-05, 2.295579e-05, 2.566222e-05, 2.078235e-05, 1.401216e-05, 
    2.051448e-06, 1.162161e-06, 1.194289e-06, 7.766965e-07, 8.312508e-07, 
    4.575514e-07, 7.439182e-07, 1.153846e-06, 5.505855e-06, 7.104932e-06,
  3.264797e-05, 2.687586e-05, 3.28753e-05, 2.44926e-05, 1.031471e-05, 
    2.859747e-06, 9.670538e-07, 6.632132e-07, 4.195998e-07, 2.789502e-07, 
    4.132827e-07, 4.092286e-07, 2.191326e-06, 2.356798e-06, 4.26302e-06,
  4.050886e-05, 3.61394e-05, 3.264516e-05, 2.638178e-05, 1.411294e-05, 
    5.66096e-06, 8.866497e-07, 1.015861e-07, 4.489445e-08, 1.477463e-07, 
    9.596129e-07, 4.647247e-07, 1.455092e-06, 1.277547e-06, 1.129626e-06,
  4.27583e-05, 4.184149e-05, 3.5837e-05, 2.891089e-05, 1.796569e-05, 
    7.125836e-06, 4.506878e-06, 2.362076e-07, 2.815538e-07, 1.288382e-07, 
    2.578793e-07, 7.105639e-07, 9.035077e-07, 9.787129e-07, 1.25366e-06,
  4.39901e-05, 3.983081e-05, 3.377431e-05, 2.71229e-05, 2.74175e-05, 
    1.809932e-05, 8.397777e-06, 5.287057e-06, 1.370149e-06, 3.292182e-07, 
    7.177838e-07, 7.715793e-07, 8.527622e-07, 8.640694e-07, 1.078835e-06,
  3.639225e-05, 3.835045e-05, 3.297274e-05, 2.48581e-05, 1.927826e-05, 
    1.363823e-05, 5.836133e-06, 8.66894e-07, 8.206516e-07, 8.107176e-07, 
    7.940715e-07, 9.873671e-07, 8.64297e-07, 5.994629e-07, 6.955583e-07,
  2.374634e-05, 1.795555e-05, 4.559719e-06, 5.470313e-07, 7.190997e-07, 
    9.854582e-07, 1.888632e-06, 2.330868e-07, 7.559794e-07, 7.921176e-07, 
    9.610749e-07, 9.794575e-07, 9.216565e-07, 6.287814e-07, 2.139869e-07,
  3.414702e-06, 4.253316e-06, 4.968169e-06, 2.485471e-06, 2.593448e-06, 
    3.652501e-06, 9.497204e-06, 2.141896e-05, 2.088893e-05, 1.507372e-05, 
    9.829269e-06, 7.450378e-06, 3.844262e-06, 1.33201e-06, 7.983639e-07,
  4.228306e-06, 6.424157e-07, 2.049045e-06, 1.960248e-06, 2.148161e-06, 
    3.539635e-06, 2.095309e-05, 2.086486e-05, 1.411998e-05, 9.952053e-06, 
    3.071206e-06, 1.507307e-06, 5.117121e-07, 3.115979e-07, 5.222121e-07,
  1.028885e-05, 5.076567e-06, 3.955885e-06, 1.787723e-06, 2.401529e-06, 
    2.626703e-06, 1.269648e-05, 1.571622e-05, 7.588694e-06, 2.506649e-06, 
    2.748141e-07, 1.461297e-07, 3.629722e-08, 4.760994e-07, 1.831054e-06,
  1.927155e-05, 2.137852e-05, 1.740783e-05, 1.040741e-05, 6.511628e-06, 
    4.359419e-06, 1.794339e-06, 2.476348e-06, 1.684982e-06, 9.212746e-07, 
    4.127372e-07, 1.691219e-07, 4.566498e-07, 1.470242e-06, 2.875555e-06,
  2.269331e-05, 2.283902e-05, 2.232342e-05, 1.633655e-05, 3.803068e-06, 
    5.470489e-06, 5.348087e-07, 5.13353e-08, 2.427896e-07, 4.690617e-07, 
    9.07686e-07, 7.496168e-07, 3.784905e-07, 1.424032e-06, 3.100979e-06,
  2.321537e-05, 2.57975e-05, 2.488574e-05, 1.374734e-05, 6.894581e-06, 
    1.255e-06, 1.893534e-07, 3.297451e-09, 2.608452e-08, 8.623273e-07, 
    7.593064e-07, 5.268296e-07, 8.501927e-07, 3.089616e-07, 2.4658e-06,
  2.283913e-05, 2.508023e-05, 2.443865e-05, 1.969748e-05, 1.116366e-05, 
    4.30336e-06, 1.073895e-06, 1.393383e-06, 8.314694e-07, 4.283274e-07, 
    8.506993e-08, 3.509772e-07, 3.052202e-07, 8.064145e-07, 4.774596e-07,
  2.209625e-05, 2.691289e-05, 2.436774e-05, 2.12846e-05, 2.042689e-05, 
    1.177073e-05, 8.773084e-06, 3.055498e-06, 1.084705e-06, 3.381583e-07, 
    3.253494e-07, 3.554684e-07, 4.209214e-07, 5.49119e-07, 3.412595e-07,
  3.097482e-05, 3.096693e-05, 2.77431e-05, 2.510835e-05, 1.742223e-05, 
    1.013482e-05, 6.33829e-06, 2.190515e-06, 1.423391e-06, 8.91169e-07, 
    6.535089e-07, 7.220158e-07, 7.711855e-07, 5.584062e-07, 6.369968e-07,
  3.810339e-05, 3.637878e-05, 1.338626e-05, 1.146227e-06, 5.698261e-07, 
    8.214113e-07, 2.259204e-06, 1.501404e-06, 6.813667e-07, 6.505707e-07, 
    9.564334e-07, 7.144233e-07, 6.165907e-07, 4.62242e-07, 3.309516e-07,
  2.229688e-06, 4.099081e-06, 2.895998e-06, 1.994349e-06, 7.308973e-07, 
    1.218212e-06, 3.159109e-06, 4.894784e-06, 5.373329e-06, 3.346826e-06, 
    1.664645e-06, 1.627435e-06, 2.075956e-06, 8.716909e-07, 1.159128e-06,
  4.707055e-06, 1.250511e-06, 1.893235e-06, 1.046368e-06, 5.370115e-07, 
    8.706325e-07, 3.506557e-06, 4.445576e-06, 4.296523e-06, 4.798381e-06, 
    1.426178e-06, 8.358986e-07, 4.657297e-07, 1.953667e-07, 2.488336e-07,
  1.076287e-05, 4.015008e-06, 2.543728e-06, 7.744647e-07, 4.706827e-07, 
    1.501431e-07, 8.337095e-07, 2.566989e-06, 2.184829e-06, 1.232051e-06, 
    1.403627e-06, 3.675111e-07, 2.569194e-07, 1.855808e-07, 8.592108e-07,
  1.7491e-05, 1.405089e-05, 9.990049e-06, 3.990743e-06, 4.921109e-07, 
    1.58562e-07, 3.108452e-07, 5.197024e-07, 3.19141e-07, 1.399898e-06, 
    1.315075e-06, 1.09347e-06, 1.671676e-06, 2.347505e-06, 4.099407e-07,
  2.337597e-05, 1.931214e-05, 1.639929e-05, 5.677717e-06, 3.446192e-08, 
    1.17116e-07, 4.594254e-08, 8.878649e-08, 1.321249e-06, 1.781677e-06, 
    1.542589e-06, 1.072241e-06, 1.373e-06, 1.504574e-06, 1.990978e-06,
  3.09816e-05, 1.950466e-05, 1.686775e-05, 1.028955e-05, 4.048681e-06, 
    2.61841e-06, 2.045805e-06, 2.438496e-06, 1.745914e-06, 2.084689e-06, 
    1.010736e-06, 6.533656e-07, 9.539676e-07, 4.489558e-07, 1.400674e-06,
  3.389299e-05, 2.406127e-05, 1.979958e-05, 1.807578e-05, 1.408929e-05, 
    1.27768e-05, 4.012485e-06, 2.416852e-06, 1.956221e-06, 1.799412e-06, 
    1.117455e-06, 9.632171e-07, 8.324523e-07, 4.95639e-07, 4.12246e-07,
  3.380329e-05, 3.166603e-05, 2.423289e-05, 1.964312e-05, 2.469109e-05, 
    1.73292e-05, 1.007946e-05, 2.753512e-06, 1.813749e-06, 8.266804e-07, 
    8.981982e-07, 1.162662e-06, 1.121155e-06, 8.525396e-07, 1.148381e-06,
  2.959201e-05, 3.332751e-05, 3.091682e-05, 2.337055e-05, 1.795414e-05, 
    1.075573e-05, 3.894243e-06, 1.882529e-06, 1.960933e-06, 6.494491e-07, 
    6.764088e-07, 9.790483e-07, 1.253062e-06, 1.187013e-06, 1.949341e-06,
  2.845599e-05, 2.672494e-05, 4.397818e-06, 3.922944e-06, 1.801196e-06, 
    1.585691e-06, 9.717656e-07, 1.758854e-06, 6.717023e-07, 5.103592e-07, 
    7.375048e-07, 6.563591e-07, 7.299367e-07, 8.086366e-07, 9.090737e-07,
  5.809568e-06, 4.087439e-06, 2.774716e-06, 2.119651e-06, 1.317067e-06, 
    6.140615e-07, 6.466643e-07, 5.361229e-07, 3.52975e-07, 1.721379e-07, 
    2.948648e-07, 1.964983e-07, 5.846107e-07, 4.498428e-07, 6.555498e-07,
  3.933382e-06, 1.334871e-06, 1.154554e-06, 1.826267e-06, 3.348599e-07, 
    1.722632e-07, 1.42491e-07, 3.283332e-07, 3.141062e-07, 9.264447e-07, 
    1.700607e-07, 9.190904e-08, 3.958489e-07, 2.480575e-07, 2.108914e-07,
  6.905189e-06, 2.827781e-06, 1.645036e-06, 1.122858e-06, 5.927272e-07, 
    2.438546e-07, 1.78902e-07, 4.503198e-07, 4.678782e-07, 6.199394e-07, 
    5.409112e-07, 5.653649e-07, 8.302437e-07, 6.872815e-07, 2.549461e-07,
  1.52603e-05, 1.164257e-05, 8.854139e-06, 6.370071e-06, 3.575092e-06, 
    2.792135e-07, 4.830258e-07, 5.20588e-07, 5.032426e-07, 1.061719e-07, 
    4.855278e-07, 5.330878e-07, 1.061891e-06, 8.577397e-07, 6.468526e-07,
  1.959613e-05, 1.712739e-05, 1.577334e-05, 1.15842e-05, 1.277221e-07, 
    3.450918e-06, 1.037262e-06, 4.351475e-07, 6.124787e-07, 8.772062e-07, 
    5.227411e-07, 2.840709e-07, 1.111696e-06, 1.290544e-06, 2.202974e-06,
  2.314723e-05, 1.812664e-05, 1.618189e-05, 1.24041e-05, 7.872067e-06, 
    3.499266e-06, 2.422338e-06, 2.70616e-06, 1.412963e-06, 2.66292e-06, 
    1.04402e-06, 7.373698e-07, 6.488388e-07, 1.008601e-06, 1.090938e-06,
  3.024438e-05, 1.824765e-05, 2.015715e-05, 1.969e-05, 1.807663e-05, 
    1.196534e-05, 3.714676e-06, 2.651365e-06, 2.778905e-06, 2.361074e-06, 
    1.669692e-06, 1.031361e-06, 4.454437e-07, 4.6057e-07, 1.679271e-07,
  3.428408e-05, 2.354149e-05, 2.319416e-05, 2.078432e-05, 2.019322e-05, 
    1.514352e-05, 8.483341e-06, 2.662222e-06, 2.231855e-06, 1.720883e-06, 
    1.752183e-06, 1.453893e-06, 6.731636e-07, 4.37937e-07, 2.127566e-07,
  3.248472e-05, 2.735995e-05, 2.971741e-05, 1.979996e-05, 1.31354e-05, 
    9.044379e-06, 3.58424e-06, 2.661619e-06, 2.550254e-06, 1.756897e-06, 
    1.328713e-06, 1.147801e-06, 1.074435e-06, 4.707385e-07, 6.734886e-08,
  3.033988e-05, 1.313729e-05, 5.996134e-06, 3.119784e-06, 2.199662e-06, 
    2.35879e-06, 2.841597e-06, 2.675009e-06, 1.444954e-06, 9.266566e-07, 
    8.399709e-07, 5.681823e-07, 5.203959e-07, 2.830384e-07, 8.893672e-08,
  1.198659e-05, 1.98838e-05, 2.394551e-05, 2.525161e-05, 2.313836e-05, 
    1.930085e-05, 1.603508e-05, 1.109463e-05, 6.074131e-06, 2.27829e-06, 
    7.707893e-07, 2.751254e-07, 2.833386e-07, 1.570762e-07, 2.979888e-07,
  5.007153e-06, 5.266357e-06, 6.75067e-06, 8.34589e-06, 5.259332e-06, 
    4.144538e-06, 4.179273e-06, 2.420898e-06, 8.920208e-07, 7.550473e-07, 
    2.783318e-07, 8.846528e-08, 6.578352e-09, 3.911628e-07, 5.277763e-07,
  9.252285e-06, 3.141567e-06, 2.722941e-06, 3.283577e-06, 1.835873e-06, 
    5.964416e-07, 1.030166e-06, 9.955653e-07, 5.080336e-07, 4.105086e-08, 
    2.475572e-07, 3.197083e-07, 4.512859e-07, 3.60369e-08, 4.531787e-07,
  2.086224e-05, 1.795343e-05, 1.104268e-05, 4.377793e-06, 2.001781e-06, 
    2.600204e-06, 5.446585e-07, 4.743996e-07, 5.484594e-07, 3.456824e-07, 
    6.474711e-08, 3.39053e-07, 1.645353e-08, 2.427249e-07, 8.183169e-07,
  2.358494e-05, 2.127078e-05, 1.856041e-05, 1.299608e-05, 3.869291e-08, 
    3.048865e-06, 2.596223e-06, 7.335164e-07, 3.872864e-07, 2.410918e-07, 
    3.683124e-07, 2.221854e-07, 1.606563e-07, 5.959909e-07, 7.414725e-07,
  1.963389e-05, 1.617664e-05, 1.637152e-05, 1.094039e-05, 7.164296e-06, 
    1.10812e-06, 3.16994e-06, 1.074135e-06, 4.665639e-09, 1.207409e-07, 
    3.508936e-07, 2.57543e-07, 2.900785e-07, 8.183646e-08, 2.258773e-08,
  2.304129e-05, 1.505641e-05, 1.544996e-05, 1.250042e-05, 1.384463e-05, 
    1.107842e-05, 4.041509e-06, 1.828053e-06, 1.10304e-06, 4.072631e-07, 
    1.014642e-07, 1.20191e-07, 2.441663e-07, 4.906233e-07, 8.885134e-08,
  2.863199e-05, 2.504204e-05, 2.440547e-05, 1.733676e-05, 1.915041e-05, 
    1.581932e-05, 8.459705e-06, 1.740535e-06, 7.63945e-07, 1.938883e-07, 
    1.403715e-07, 1.501356e-07, 2.600847e-07, 4.542035e-07, 6.536509e-07,
  1.910925e-05, 2.003335e-05, 2.392938e-05, 1.789904e-05, 1.537679e-05, 
    9.70657e-06, 3.306081e-06, 1.376015e-06, 3.600571e-07, 2.70637e-07, 
    1.787649e-07, 3.308938e-07, 7.725192e-07, 1.177078e-06, 1.001646e-06,
  2.018858e-05, 2.038868e-05, 9.464126e-06, 3.956206e-06, 3.187581e-06, 
    1.883678e-06, 7.847332e-07, 4.043358e-07, 2.794567e-07, 3.407937e-07, 
    8.426778e-07, 2.470072e-06, 5.963811e-06, 1.058871e-05, 1.278093e-05,
  2.247338e-05, 5.497442e-05, 6.487512e-05, 7.69682e-05, 8.256343e-05, 
    7.477737e-05, 6.342655e-05, 5.135422e-05, 3.873288e-05, 2.527641e-05, 
    1.710361e-05, 1.519041e-05, 1.542377e-05, 1.408392e-05, 1.108349e-05,
  9.481085e-06, 2.200011e-05, 3.813907e-05, 5.656371e-05, 4.951813e-05, 
    4.482274e-05, 5.206445e-05, 3.889872e-05, 2.717896e-05, 1.795305e-05, 
    9.519747e-06, 9.343456e-06, 9.176719e-06, 7.903537e-06, 5.73744e-06,
  7.394661e-06, 4.39625e-06, 7.5491e-06, 1.060352e-05, 9.747168e-06, 
    1.025674e-05, 1.297766e-05, 1.475848e-05, 1.169604e-05, 6.820172e-06, 
    3.730247e-06, 2.455343e-06, 2.949311e-06, 3.422921e-06, 1.908014e-06,
  2.520586e-05, 1.878973e-05, 8.879405e-06, 3.700886e-06, 2.858244e-06, 
    2.055236e-06, 1.744975e-06, 1.909014e-06, 1.527687e-06, 1.802853e-06, 
    4.403115e-07, 2.051673e-07, 2.914799e-07, 6.226022e-07, 4.439495e-07,
  1.898505e-05, 2.216171e-05, 1.80613e-05, 8.048169e-06, 1.369201e-06, 
    1.599058e-06, 7.491616e-07, 2.314609e-07, 3.650434e-07, 6.357157e-07, 
    5.888836e-07, 7.834977e-07, 4.875553e-08, 5.657664e-09, 9.695563e-09,
  1.072721e-05, 1.386127e-05, 1.679449e-05, 1.042802e-05, 7.003775e-06, 
    1.049008e-06, 2.503493e-06, 4.17013e-07, 3.342607e-09, 3.530589e-07, 
    4.349263e-07, 5.111453e-07, 1.071795e-07, 2.872376e-08, 2.465306e-08,
  9.419412e-06, 4.052482e-06, 8.765036e-06, 1.160826e-05, 1.461285e-05, 
    8.948038e-06, 2.996527e-06, 9.173634e-07, 3.962265e-07, 3.642869e-07, 
    2.724397e-07, 1.020833e-07, 2.60515e-07, 7.341396e-07, 2.290924e-07,
  4.530495e-05, 1.59008e-05, 1.415644e-05, 1.573885e-05, 1.253798e-05, 
    1.221583e-05, 3.821303e-06, 6.295296e-07, 1.361731e-07, 3.761324e-07, 
    3.160394e-07, 3.713703e-07, 5.458016e-07, 5.199722e-07, 2.418919e-07,
  6.979654e-05, 5.408105e-05, 4.486703e-05, 3.237692e-05, 8.748232e-06, 
    5.132181e-06, 1.53119e-06, 1.433282e-06, 2.131558e-06, 3.131672e-06, 
    3.593023e-06, 4.065197e-06, 4.4706e-06, 3.692668e-06, 1.482655e-06,
  1.86878e-05, 2.828561e-05, 1.496186e-05, 1.251759e-06, 9.543738e-07, 
    4.161297e-06, 8.768383e-06, 1.226116e-05, 1.319164e-05, 1.749725e-05, 
    2.570595e-05, 3.276149e-05, 3.288817e-05, 2.477531e-05, 1.11593e-05,
  2.084849e-06, 1.713065e-05, 4.200431e-05, 7.705107e-05, 9.335952e-05, 
    7.666548e-05, 6.117464e-05, 5.001589e-05, 3.914263e-05, 2.600627e-05, 
    2.519197e-05, 3.721104e-05, 4.363648e-05, 3.65191e-05, 2.795077e-05,
  6.899076e-07, 4.683283e-06, 1.743525e-05, 5.876632e-05, 8.204049e-05, 
    6.83589e-05, 7.762278e-05, 5.677858e-05, 4.182164e-05, 3.146217e-05, 
    2.414873e-05, 3.524589e-05, 4.080439e-05, 3.544439e-05, 3.318064e-05,
  7.414491e-06, 1.879704e-06, 5.034423e-06, 1.118701e-05, 1.527519e-05, 
    1.626297e-05, 1.957157e-05, 3.794494e-05, 3.546348e-05, 2.695273e-05, 
    2.136301e-05, 2.85413e-05, 3.992558e-05, 4.421669e-05, 3.575453e-05,
  1.807606e-05, 1.947175e-05, 8.966237e-06, 3.396979e-06, 3.666546e-06, 
    2.877337e-06, 9.36874e-07, 1.392501e-06, 3.865251e-06, 1.307741e-05, 
    1.169614e-05, 1.417179e-05, 2.093745e-05, 2.615259e-05, 2.291756e-05,
  1.794967e-05, 1.560407e-05, 1.489286e-05, 2.660413e-06, 6.389815e-07, 
    5.870043e-07, 1.258894e-07, 1.792656e-08, 3.345789e-07, 1.248027e-06, 
    2.685251e-06, 3.957063e-06, 5.737561e-06, 7.505084e-06, 1.050662e-05,
  2.325135e-05, 1.570479e-05, 9.888739e-06, 6.826252e-06, 1.134057e-06, 
    3.516849e-07, 1.920114e-07, 1.131516e-08, 1.112802e-07, 6.783527e-08, 
    6.424603e-07, 7.72041e-07, 1.426232e-06, 2.261329e-06, 3.774397e-06,
  6.708279e-05, 2.538239e-05, 5.237781e-06, 1.028744e-05, 1.170444e-05, 
    6.63607e-06, 1.957796e-07, 9.655134e-09, 7.109553e-08, 4.26839e-07, 
    2.15741e-07, 3.535022e-07, 8.95669e-07, 1.277151e-06, 1.180052e-06,
  7.299881e-05, 3.473553e-05, 2.504417e-05, 1.519707e-05, 7.840908e-06, 
    6.418344e-06, 4.713171e-06, 8.214049e-07, 3.246736e-06, 2.761902e-06, 
    1.13395e-06, 3.340384e-07, 5.39261e-07, 6.717866e-07, 9.250273e-07,
  3.027802e-05, 2.613423e-05, 2.084891e-05, 8.61244e-06, 5.619894e-06, 
    7.22531e-06, 5.875721e-06, 5.63458e-06, 7.545102e-06, 1.264743e-05, 
    1.551386e-05, 1.106167e-05, 3.558099e-06, 9.614512e-07, 7.888593e-07,
  1.371416e-05, 8.144068e-06, 3.897225e-06, 3.098846e-06, 4.167006e-06, 
    7.992925e-06, 9.559688e-06, 7.896024e-06, 7.845911e-06, 1.043459e-05, 
    1.651973e-05, 2.220478e-05, 1.904536e-05, 9.423285e-06, 3.337988e-06,
  3.704431e-07, 4.745986e-07, 1.317223e-06, 7.916789e-06, 2.035666e-05, 
    2.179884e-05, 1.691894e-05, 7.042021e-06, 5.420142e-06, 9.143184e-06, 
    1.215574e-05, 1.140678e-05, 7.168139e-06, 4.33764e-06, 4.028371e-06,
  6.840273e-07, 5.98123e-07, 5.953858e-07, 3.650065e-06, 9.324032e-06, 
    1.166197e-05, 1.715612e-05, 1.942563e-05, 1.613294e-05, 1.712916e-05, 
    1.913247e-05, 1.909018e-05, 1.490773e-05, 7.361266e-06, 6.403727e-06,
  1.610424e-06, 1.360959e-06, 8.334713e-07, 1.411829e-06, 1.889955e-06, 
    1.818362e-06, 5.473657e-06, 1.924984e-05, 2.553122e-05, 2.345994e-05, 
    2.095543e-05, 2.172812e-05, 2.185604e-05, 1.942151e-05, 1.711482e-05,
  2.657823e-06, 1.163094e-05, 1.106097e-05, 1.180364e-06, 1.339177e-06, 
    1.161123e-06, 6.607388e-07, 2.140319e-06, 4.202658e-06, 1.072971e-05, 
    1.428911e-05, 1.588159e-05, 2.068638e-05, 2.593094e-05, 2.30701e-05,
  1.463285e-06, 7.435142e-06, 1.028162e-05, 2.781951e-06, 1.697861e-06, 
    1.849492e-06, 4.553574e-07, 2.628965e-08, 8.446047e-08, 5.514052e-07, 
    2.276698e-06, 3.949911e-06, 1.035331e-05, 1.654339e-05, 2.468448e-05,
  4.537449e-06, 1.475776e-05, 3.355188e-06, 5.237712e-06, 3.28806e-06, 
    2.463152e-06, 2.164488e-06, 1.962705e-07, 4.130217e-08, 1.167604e-07, 
    2.247622e-07, 2.86492e-07, 8.793272e-07, 4.681766e-06, 1.590597e-05,
  1.628279e-05, 1.520209e-05, 7.974718e-06, 3.069415e-06, 7.452529e-06, 
    3.984482e-06, 2.885123e-06, 1.277442e-06, 2.732253e-06, 8.536127e-07, 
    6.245489e-08, 9.433543e-08, 3.540201e-07, 1.152044e-06, 3.422219e-06,
  1.596676e-05, 1.990455e-05, 1.422348e-05, 7.092973e-06, 9.88748e-06, 
    9.243703e-06, 3.638552e-06, 2.219278e-06, 2.465634e-06, 2.974081e-06, 
    8.812981e-07, 9.321166e-08, 2.152305e-07, 6.0433e-07, 1.266203e-06,
  1.63579e-05, 2.274414e-05, 1.877287e-05, 4.629973e-06, 4.101745e-06, 
    2.192974e-06, 9.597397e-07, 8.791233e-09, 1.28773e-06, 1.745118e-06, 
    6.535606e-07, 7.478744e-07, 1.061108e-06, 4.86961e-07, 6.49579e-07,
  1.640768e-05, 1.599999e-05, 6.777202e-06, 2.612357e-06, 1.126879e-06, 
    7.716174e-07, 5.424218e-07, 9.212624e-09, 8.073079e-07, 1.296904e-06, 
    8.764292e-07, 7.961344e-07, 1.5584e-06, 1.588168e-06, 1.045431e-06,
  3.738094e-06, 1.743475e-06, 1.042703e-06, 1.043415e-06, 2.828069e-07, 
    2.373975e-07, 6.905639e-07, 2.683772e-06, 3.301845e-06, 4.560316e-06, 
    4.164035e-06, 3.677985e-06, 3.432438e-06, 1.341483e-06, 1.420442e-06,
  5.080967e-06, 2.454479e-06, 1.739459e-06, 1.17977e-06, 1.343112e-06, 
    6.679763e-07, 4.782628e-07, 1.866478e-07, 1.936055e-06, 3.974634e-06, 
    4.991648e-06, 5.164352e-06, 4.971861e-06, 5.041555e-06, 3.550169e-06,
  5.735102e-06, 3.245739e-06, 2.443895e-06, 1.704405e-06, 1.171373e-06, 
    2.930367e-06, 8.104163e-07, 5.370582e-07, 5.949875e-07, 1.430944e-06, 
    1.819624e-06, 3.924525e-06, 4.507045e-06, 5.287633e-06, 4.351044e-06,
  1.694653e-05, 8.987953e-06, 3.809652e-06, 2.025714e-06, 1.068555e-06, 
    7.67241e-07, 2.682374e-06, 7.363229e-07, 1.734278e-07, 3.500582e-07, 
    8.930646e-07, 2.510007e-07, 1.255146e-06, 2.573346e-06, 4.726818e-06,
  2.656949e-05, 1.870987e-05, 1.225796e-05, 3.214316e-06, 1.615452e-06, 
    1.451653e-06, 1.526284e-06, 3.154029e-06, 4.373047e-07, 2.639032e-07, 
    2.244248e-07, 3.24726e-07, 3.411205e-07, 2.503605e-07, 2.405729e-06,
  4.325556e-05, 3.100582e-05, 1.942591e-05, 9.368125e-06, 1.448506e-06, 
    2.325952e-06, 2.561251e-06, 1.654121e-06, 7.066637e-07, 3.104794e-07, 
    1.272527e-07, 3.308991e-08, 2.009311e-07, 2.104369e-07, 7.750074e-07,
  4.645477e-05, 4.379969e-05, 2.831888e-05, 1.118861e-05, 5.660671e-06, 
    4.310426e-06, 3.789582e-06, 2.006663e-06, 1.65986e-06, 1.502262e-06, 
    1.634783e-07, 9.395175e-09, 9.084583e-08, 1.703691e-07, 4.076244e-07,
  4.470369e-05, 4.100278e-05, 3.02665e-05, 1.437437e-05, 1.345012e-05, 
    1.494728e-05, 4.416102e-06, 2.119628e-06, 1.713269e-06, 2.368293e-06, 
    1.032276e-06, 2.282564e-08, 6.386973e-08, 7.896102e-08, 2.208626e-08,
  4.248709e-05, 3.833165e-05, 2.842392e-05, 1.166927e-05, 6.550031e-06, 
    2.537269e-06, 2.158926e-06, 2.095207e-06, 2.135181e-06, 1.357547e-06, 
    1.077097e-06, 2.94852e-07, 5.689801e-08, 7.476635e-08, 4.239399e-08,
  3.878346e-05, 3.295146e-05, 1.082113e-05, 3.138174e-06, 2.218989e-06, 
    2.335668e-06, 3.120203e-06, 3.124299e-06, 1.790188e-06, 1.686173e-06, 
    1.486743e-06, 5.510808e-07, 7.737781e-08, 1.003662e-07, 7.487069e-08,
  1.002261e-05, 1.300508e-05, 2.123673e-05, 2.415569e-05, 1.54745e-05, 
    6.550293e-06, 2.761349e-06, 1.942022e-06, 3.137825e-06, 5.349551e-06, 
    6.510968e-06, 6.274766e-06, 4.432273e-06, 2.20082e-06, 2.459282e-06,
  7.809961e-06, 7.152735e-06, 1.258237e-05, 1.781876e-05, 1.386598e-05, 
    4.991332e-06, 2.108462e-06, 1.511657e-06, 1.234424e-06, 2.690159e-06, 
    3.328312e-06, 6.128702e-06, 3.912153e-06, 3.254523e-06, 3.453968e-06,
  5.763479e-06, 6.282279e-06, 8.341337e-06, 1.417084e-05, 1.026841e-05, 
    4.502827e-06, 1.904857e-06, 1.394821e-06, 7.519715e-07, 6.138328e-07, 
    8.53786e-07, 1.053163e-06, 1.933304e-06, 4.08877e-06, 2.012356e-06,
  1.691516e-05, 1.123402e-05, 1.014305e-05, 1.219704e-05, 1.039716e-05, 
    4.706012e-06, 3.910392e-06, 1.535459e-06, 8.194655e-07, 2.993788e-07, 
    2.456751e-07, 2.466351e-07, 4.577115e-07, 7.192464e-07, 4.716583e-07,
  2.213007e-05, 1.886514e-05, 1.731329e-05, 1.36614e-05, 1.020585e-05, 
    7.483199e-06, 4.296412e-06, 5.258951e-06, 3.344277e-06, 9.270949e-07, 
    2.851637e-07, 8.894482e-08, 1.595475e-07, 3.239537e-07, 6.779746e-07,
  3.355317e-05, 2.749858e-05, 1.550251e-05, 1.542412e-05, 1.05349e-05, 
    6.560779e-06, 5.324903e-06, 5.658895e-06, 2.961576e-06, 4.083936e-07, 
    3.699186e-07, 1.112359e-07, 1.207115e-07, 3.015309e-07, 5.515066e-07,
  5.636282e-05, 4.732815e-05, 3.24291e-05, 1.37804e-05, 1.46927e-05, 
    9.929533e-06, 4.060797e-06, 4.736636e-06, 2.885778e-06, 1.957268e-06, 
    7.909385e-07, 1.058534e-07, 3.232547e-08, 9.238666e-08, 2.767914e-07,
  5.332501e-05, 5.166496e-05, 3.715577e-05, 1.888223e-05, 1.871002e-05, 
    1.891944e-05, 3.759762e-06, 4.143548e-06, 2.545458e-06, 2.43444e-06, 
    1.335827e-06, 7.035648e-07, 1.798498e-07, 1.270514e-07, 1.465116e-08,
  2.853686e-05, 3.322267e-05, 3.33967e-05, 1.998371e-05, 1.636182e-05, 
    6.128267e-06, 4.548167e-06, 3.666117e-06, 2.183562e-06, 2.676299e-06, 
    1.509904e-06, 1.102972e-06, 1.519856e-07, 1.951129e-07, 5.717125e-08,
  2.032275e-05, 1.794341e-05, 9.37396e-06, 5.72431e-06, 5.376611e-06, 
    5.018314e-06, 5.249626e-06, 4.95162e-06, 2.188923e-06, 2.344216e-06, 
    2.241896e-06, 5.431074e-07, 1.972284e-07, 2.454506e-07, 1.991233e-07,
  3.918236e-06, 1.630734e-06, 3.278267e-06, 4.753313e-06, 8.10136e-06, 
    1.138696e-05, 1.750577e-05, 2.758828e-05, 3.171087e-05, 2.547738e-05, 
    1.640234e-05, 9.914282e-06, 4.78198e-06, 4.815191e-06, 3.059838e-06,
  2.262394e-06, 1.810061e-06, 2.392478e-06, 4.806646e-06, 7.15236e-06, 
    7.795821e-06, 1.587894e-05, 2.156379e-05, 2.236606e-05, 2.144505e-05, 
    1.38785e-05, 1.129622e-05, 5.472916e-06, 1.188586e-06, 3.473401e-06,
  2.597837e-06, 1.629152e-06, 3.686995e-06, 7.268598e-06, 5.699285e-06, 
    5.544183e-06, 1.057216e-05, 2.014336e-05, 2.144018e-05, 1.782343e-05, 
    1.286005e-05, 7.17363e-06, 4.262272e-06, 2.161533e-06, 5.391542e-07,
  1.145168e-05, 1.063569e-05, 6.393755e-06, 7.335982e-06, 7.550377e-06, 
    8.438966e-06, 6.657797e-06, 1.210788e-05, 1.51401e-05, 1.573932e-05, 
    9.370006e-06, 3.639532e-06, 1.632167e-06, 6.097247e-07, 5.247261e-08,
  1.447172e-05, 1.63811e-05, 1.436229e-05, 9.578325e-06, 5.726391e-06, 
    9.332061e-06, 8.870295e-06, 2.113522e-06, 1.974792e-06, 6.726129e-06, 
    4.410128e-06, 1.299115e-06, 5.946002e-07, 9.163808e-08, 1.517707e-08,
  1.899771e-05, 2.01811e-05, 1.631627e-05, 1.375128e-05, 7.469602e-06, 
    5.668726e-06, 1.04996e-05, 9.880395e-06, 6.402741e-06, 4.209071e-06, 
    1.695805e-06, 9.293067e-07, 2.6313e-07, 2.436168e-08, 1.430506e-08,
  1.751487e-05, 2.947107e-05, 1.515043e-05, 1.36219e-05, 1.495119e-05, 
    1.136922e-05, 7.382664e-06, 9.621207e-06, 7.170947e-06, 4.246391e-06, 
    1.752399e-06, 5.644319e-07, 2.056386e-07, 2.396253e-07, 1.094312e-08,
  1.305878e-05, 2.340616e-05, 1.357658e-05, 1.341585e-05, 2.000244e-05, 
    1.952168e-05, 7.884069e-06, 5.205297e-06, 3.8424e-06, 2.802563e-06, 
    1.833672e-06, 8.567601e-07, 2.909796e-07, 2.200761e-07, 4.179592e-09,
  1.400284e-05, 2.279945e-05, 1.218394e-05, 8.782249e-06, 1.591799e-05, 
    9.480282e-06, 5.026709e-06, 4.552455e-06, 3.565377e-06, 2.726267e-06, 
    1.745247e-06, 5.0515e-07, 3.18843e-07, 2.148452e-07, 2.60554e-08,
  1.475727e-05, 1.99706e-05, 9.587568e-06, 3.626408e-06, 1.825503e-06, 
    2.536648e-06, 4.931187e-06, 4.499249e-06, 3.080037e-06, 2.656844e-06, 
    1.408623e-06, 3.379045e-07, 3.383187e-07, 4.319981e-07, 4.886247e-07,
  1.02661e-05, 6.481072e-06, 7.314729e-06, 7.715804e-06, 4.447549e-06, 
    3.010789e-06, 2.596185e-06, 4.690359e-06, 9.778532e-06, 1.640989e-05, 
    2.182371e-05, 1.999979e-05, 1.276732e-05, 3.911226e-06, 1.735047e-06,
  1.203702e-05, 8.32177e-06, 1.079413e-05, 1.049386e-05, 6.387526e-06, 
    3.556489e-06, 1.439387e-06, 4.313099e-06, 1.002005e-05, 1.885415e-05, 
    2.634994e-05, 2.437782e-05, 1.538023e-05, 3.192836e-06, 1.548861e-06,
  1.712569e-05, 1.451124e-05, 1.673554e-05, 1.55166e-05, 8.164289e-06, 
    2.025733e-06, 1.11976e-06, 5.122464e-06, 1.078169e-05, 2.036364e-05, 
    2.916608e-05, 2.677645e-05, 1.787345e-05, 7.05408e-06, 2.687206e-06,
  2.906211e-05, 3.023279e-05, 2.21431e-05, 1.786725e-05, 6.653544e-06, 
    1.647868e-06, 2.60052e-06, 3.581652e-06, 9.76525e-06, 1.926818e-05, 
    2.412031e-05, 2.394354e-05, 1.603064e-05, 7.906152e-06, 2.618192e-06,
  4.599498e-05, 4.539936e-05, 3.648326e-05, 1.536203e-05, 1.853719e-06, 
    1.26651e-06, 4.652468e-06, 1.56686e-06, 4.368445e-06, 1.211893e-05, 
    1.519855e-05, 1.550053e-05, 1.105418e-05, 5.199694e-06, 1.991128e-06,
  6.184679e-05, 5.268906e-05, 2.20933e-05, 1.208598e-05, 1.421496e-06, 
    7.004965e-07, 4.486201e-06, 8.772382e-06, 1.08612e-05, 1.087341e-05, 
    9.592977e-06, 9.278818e-06, 6.524303e-06, 3.544512e-06, 4.08107e-07,
  7.456303e-05, 4.08968e-05, 2.301297e-05, 1.405381e-05, 8.979438e-06, 
    8.456907e-06, 5.286231e-06, 1.103277e-05, 1.224828e-05, 9.106844e-06, 
    8.801632e-06, 7.330701e-06, 3.176512e-06, 1.149125e-06, 1.029395e-07,
  5.088366e-05, 3.066545e-05, 2.286633e-05, 1.642029e-05, 1.710276e-05, 
    1.303432e-05, 7.478015e-06, 6.280446e-06, 7.005077e-06, 6.671843e-06, 
    5.950906e-06, 4.109958e-06, 1.502585e-06, 5.101936e-07, 3.757414e-08,
  2.932997e-05, 2.128541e-05, 2.021781e-05, 2.136692e-05, 1.659944e-05, 
    8.382111e-06, 5.255194e-06, 5.91722e-06, 5.453644e-06, 4.114646e-06, 
    3.513745e-06, 1.752811e-06, 7.16507e-07, 2.993449e-07, 2.100603e-08,
  1.555406e-05, 7.394597e-06, 7.806731e-06, 3.764953e-07, 1.024057e-07, 
    2.053942e-06, 3.130464e-06, 3.990162e-06, 3.494605e-06, 2.537706e-06, 
    1.815186e-06, 9.404219e-07, 5.935387e-07, 5.057615e-07, 1.302866e-07,
  7.500432e-06, 6.276397e-06, 9.686873e-06, 1.186457e-05, 1.621335e-05, 
    2.316682e-05, 2.54918e-05, 3.009324e-05, 3.071205e-05, 2.684601e-05, 
    2.264406e-05, 1.807772e-05, 1.512922e-05, 9.408494e-06, 7.041894e-06,
  2.029599e-06, 2.277784e-06, 4.419565e-06, 1.109387e-05, 1.910815e-05, 
    3.313061e-05, 3.479791e-05, 2.913418e-05, 2.396856e-05, 1.831239e-05, 
    1.363726e-05, 1.17603e-05, 1.164785e-05, 6.111868e-06, 7.885887e-06,
  2.882682e-06, 2.465515e-06, 6.392329e-06, 1.783007e-05, 3.221219e-05, 
    3.974924e-05, 3.027392e-05, 2.109661e-05, 1.327985e-05, 7.667522e-06, 
    5.886417e-06, 6.849648e-06, 1.316818e-05, 1.457786e-05, 1.484811e-05,
  1.25783e-05, 1.407898e-05, 1.650421e-05, 2.679464e-05, 3.436295e-05, 
    1.896481e-05, 1.207677e-05, 1.141167e-05, 5.786248e-06, 3.376701e-06, 
    3.246004e-06, 8.364134e-06, 1.796407e-05, 2.052852e-05, 1.596666e-05,
  1.910347e-05, 2.437037e-05, 2.798059e-05, 2.208933e-05, 1.550651e-05, 
    1.12715e-05, 5.963661e-06, 3.891077e-06, 1.721341e-06, 2.235362e-06, 
    4.491907e-06, 1.327103e-05, 2.162529e-05, 1.883666e-05, 1.624404e-05,
  2.662209e-05, 2.801894e-05, 2.386016e-05, 1.43765e-05, 1.137532e-05, 
    6.638287e-06, 6.226e-06, 5.163729e-06, 2.68192e-06, 3.914221e-06, 
    7.749346e-06, 1.633876e-05, 2.297385e-05, 2.238568e-05, 1.614264e-05,
  2.79868e-05, 2.824463e-05, 2.838491e-05, 2.374069e-05, 1.990947e-05, 
    1.397134e-05, 6.524056e-06, 5.485941e-06, 5.52637e-06, 7.298049e-06, 
    1.264435e-05, 1.876028e-05, 2.128714e-05, 2.054624e-05, 1.348991e-05,
  2.54805e-05, 2.846113e-05, 3.169584e-05, 2.104206e-05, 2.270032e-05, 
    1.623183e-05, 6.725594e-06, 5.435504e-06, 7.118705e-06, 1.000851e-05, 
    1.519139e-05, 1.748473e-05, 1.70643e-05, 1.373863e-05, 9.106657e-06,
  1.661746e-05, 2.298328e-05, 1.923476e-05, 1.634393e-05, 1.573469e-05, 
    1.044251e-05, 5.838257e-06, 8.045972e-06, 9.66631e-06, 1.08556e-05, 
    1.182265e-05, 1.23911e-05, 1.036308e-05, 7.420772e-06, 3.56383e-06,
  9.793564e-06, 8.977941e-06, 4.01507e-06, 2.199294e-06, 3.876281e-07, 
    4.261337e-06, 5.697485e-06, 6.894397e-06, 7.44917e-06, 7.440951e-06, 
    7.10952e-06, 6.583027e-06, 4.887634e-06, 2.814894e-06, 1.314346e-06,
  1.465965e-06, 6.21954e-07, 4.488605e-07, 1.069178e-06, 3.988895e-06, 
    3.216951e-06, 3.614449e-06, 2.982127e-06, 6.103458e-06, 7.964066e-06, 
    8.877403e-06, 1.128938e-05, 1.869366e-05, 2.509514e-05, 2.709818e-05,
  3.915974e-06, 5.423079e-07, 6.744094e-08, 5.318657e-06, 4.194224e-06, 
    1.833396e-06, 3.009242e-06, 2.194523e-06, 1.776645e-06, 4.314571e-06, 
    4.800116e-06, 8.828812e-06, 1.285068e-05, 1.876489e-05, 2.553723e-05,
  7.672255e-06, 8.889693e-07, 3.837896e-07, 2.599234e-06, 4.230523e-06, 
    1.996916e-06, 1.666152e-06, 7.054029e-06, 4.628785e-06, 1.629025e-06, 
    2.810186e-06, 5.835046e-06, 1.012714e-05, 1.810517e-05, 1.918484e-05,
  1.922769e-05, 1.895546e-05, 8.435586e-06, 4.433317e-06, 7.520426e-06, 
    7.195339e-06, 2.012606e-06, 1.852155e-06, 2.047414e-06, 1.383837e-06, 
    2.061012e-06, 4.420805e-06, 8.050122e-06, 1.456048e-05, 1.276262e-05,
  2.032015e-05, 1.459773e-05, 1.961146e-05, 1.158763e-05, 3.0559e-06, 
    1.037855e-05, 9.227243e-06, 1.687829e-06, 2.14584e-06, 2.784339e-06, 
    3.951252e-06, 3.972805e-06, 7.599303e-06, 9.828771e-06, 1.118859e-05,
  2.270099e-05, 1.60068e-05, 1.969465e-05, 1.791925e-05, 8.992979e-06, 
    8.115885e-06, 1.089874e-05, 1.143769e-05, 9.196466e-06, 7.01063e-06, 
    4.782364e-06, 4.499675e-06, 5.585126e-06, 6.244267e-06, 5.262765e-06,
  2.385942e-05, 1.801114e-05, 2.093212e-05, 1.966529e-05, 2.32998e-05, 
    1.509428e-05, 7.39292e-06, 8.526657e-06, 7.351793e-06, 5.66489e-06, 
    5.6875e-06, 6.262261e-06, 5.703084e-06, 5.861928e-06, 5.146781e-06,
  2.263777e-05, 1.941481e-05, 1.788681e-05, 1.791216e-05, 2.386957e-05, 
    1.626531e-05, 6.009393e-06, 5.62708e-06, 7.106192e-06, 7.624613e-06, 
    7.396301e-06, 7.571454e-06, 7.23396e-06, 9.764952e-06, 1.109576e-05,
  2.322378e-05, 1.85846e-05, 1.33608e-05, 7.698451e-06, 1.077314e-05, 
    7.651593e-06, 4.695394e-06, 5.340069e-06, 6.693395e-06, 7.437671e-06, 
    8.270659e-06, 1.041144e-05, 1.106889e-05, 1.059733e-05, 7.102509e-06,
  2.184197e-05, 1.218207e-05, 8.711478e-06, 2.514586e-06, 9.863611e-07, 
    1.471378e-06, 2.148703e-06, 2.588908e-06, 2.781677e-06, 3.609101e-06, 
    5.94764e-06, 8.659257e-06, 8.570541e-06, 6.2402e-06, 3.603171e-06,
  2.330482e-05, 7.670861e-06, 1.541746e-06, 6.880825e-07, 1.531325e-06, 
    2.524191e-06, 1.52616e-06, 1.401784e-06, 2.802648e-06, 3.430477e-06, 
    5.912229e-06, 9.117658e-06, 1.256891e-05, 1.139843e-05, 9.187956e-06,
  2.777975e-05, 8.493864e-06, 1.682397e-06, 1.788343e-07, 1.71558e-06, 
    7.085832e-07, 1.200717e-06, 1.199454e-06, 1.763713e-06, 2.736565e-06, 
    5.651933e-06, 8.248034e-06, 1.154465e-05, 1.000433e-05, 9.524196e-06,
  3.943063e-05, 1.532194e-05, 3.905258e-06, 2.836666e-07, 2.518962e-06, 
    4.798524e-07, 2.562938e-07, 5.586401e-06, 5.850955e-06, 5.211981e-06, 
    5.960464e-06, 7.868308e-06, 8.342846e-06, 8.592656e-06, 1.034784e-05,
  5.460326e-05, 3.471784e-05, 1.523437e-05, 1.181574e-06, 5.016772e-06, 
    2.568703e-06, 5.209785e-07, 2.386732e-06, 2.635081e-06, 5.269239e-06, 
    8.850811e-06, 8.653848e-06, 7.790601e-06, 7.220422e-06, 9.30483e-06,
  6.643739e-05, 4.894125e-05, 2.605669e-05, 7.2119e-06, 1.626073e-06, 
    4.280874e-06, 3.606587e-06, 6.233872e-07, 4.755762e-06, 7.303273e-06, 
    9.744679e-06, 9.053348e-06, 8.886236e-06, 5.464107e-06, 8.208337e-06,
  7.618195e-05, 6.569538e-05, 4.167958e-05, 9.576251e-06, 3.911701e-06, 
    4.599705e-06, 5.661767e-06, 4.467712e-06, 5.390471e-06, 9.695054e-06, 
    6.3471e-06, 6.869147e-06, 7.189444e-06, 3.853641e-06, 3.205971e-06,
  8.460083e-05, 8.360187e-05, 5.935109e-05, 1.60484e-05, 7.250846e-06, 
    6.065704e-06, 3.457653e-06, 2.43328e-06, 3.087699e-06, 3.913538e-06, 
    3.019168e-06, 3.904529e-06, 4.225626e-06, 2.759758e-06, 1.672761e-06,
  8.837183e-05, 9.56881e-05, 7.528481e-05, 3.114056e-05, 6.760357e-06, 
    5.914074e-06, 2.065501e-06, 1.597724e-06, 1.429879e-06, 1.26408e-06, 
    1.863349e-06, 1.957597e-06, 2.506782e-06, 2.375029e-06, 1.647495e-06,
  9.854021e-05, 0.0001034592, 9.047279e-05, 5.684164e-05, 7.260568e-06, 
    1.574511e-06, 1.776064e-06, 8.20609e-07, 7.000588e-07, 6.198237e-07, 
    9.389245e-07, 1.450374e-06, 1.669475e-06, 1.127634e-06, 5.565163e-07,
  0.0001002569, 0.0001031726, 8.961857e-05, 7.790478e-05, 2.472395e-05, 
    7.863225e-07, 3.751956e-07, 5.695377e-07, 4.113091e-07, 2.378432e-07, 
    4.913866e-07, 8.277875e-07, 9.324611e-07, 6.032565e-07, 3.010057e-07,
  8.346894e-05, 8.520084e-05, 4.378451e-05, 1.69686e-06, 7.531766e-07, 
    1.271977e-06, 1.197663e-06, 2.941062e-06, 6.552918e-06, 7.871186e-06, 
    7.843612e-06, 7.849076e-06, 6.99077e-06, 4.552373e-06, 2.422817e-06,
  8.342534e-05, 7.842143e-05, 3.653023e-05, 1.789353e-06, 7.080303e-07, 
    1.28401e-06, 1.136621e-06, 1.394136e-06, 3.212193e-06, 6.221606e-06, 
    6.919135e-06, 7.683828e-06, 7.31979e-06, 3.290456e-06, 1.201776e-06,
  7.617329e-05, 7.68613e-05, 3.959262e-05, 1.728615e-06, 6.233783e-07, 
    1.334967e-06, 7.065544e-07, 2.94286e-06, 7.724323e-06, 6.739822e-06, 
    4.917105e-06, 4.615119e-06, 3.130067e-06, 1.290331e-06, 1.185098e-06,
  6.216995e-05, 7.6207e-05, 5.206746e-05, 2.768907e-06, 1.81455e-06, 
    1.985059e-07, 1.022425e-06, 2.339721e-06, 3.137269e-06, 8.762342e-06, 
    5.831669e-06, 2.672703e-06, 2.311768e-06, 2.096993e-06, 4.076026e-06,
  4.584041e-05, 7.747547e-05, 7.415206e-05, 7.589092e-06, 3.019535e-06, 
    3.192879e-06, 4.958005e-07, 8.672862e-07, 4.262285e-06, 8.737335e-06, 
    7.856104e-06, 5.295424e-06, 7.920959e-06, 9.927136e-06, 1.378568e-05,
  3.295397e-05, 5.700791e-05, 8.271032e-05, 1.784947e-05, 4.789771e-06, 
    5.150137e-06, 4.551979e-06, 2.875574e-06, 2.767773e-06, 7.972891e-06, 
    5.019493e-06, 4.74468e-06, 8.663947e-06, 1.011144e-05, 1.109858e-05,
  2.549784e-05, 3.523669e-05, 7.207553e-05, 2.842172e-05, 8.114507e-06, 
    7.233625e-06, 4.477253e-06, 2.566751e-06, 1.890506e-06, 2.396163e-06, 
    2.342544e-06, 3.800514e-06, 6.932552e-06, 9.961757e-06, 1.272095e-05,
  2.122107e-05, 2.236886e-05, 5.391936e-05, 3.469976e-05, 1.215068e-05, 
    8.966001e-06, 4.071103e-06, 1.738159e-06, 7.747362e-07, 1.025233e-06, 
    1.783627e-06, 3.286376e-06, 6.120503e-06, 9.79573e-06, 1.394318e-05,
  2.122872e-05, 2.214413e-05, 3.817843e-05, 3.803272e-05, 8.776588e-06, 
    6.448665e-06, 3.084116e-06, 1.522437e-06, 7.618314e-07, 7.716606e-07, 
    1.530714e-06, 3.049075e-06, 5.607119e-06, 9.315502e-06, 1.510954e-05,
  1.896386e-05, 2.232265e-05, 2.774505e-05, 3.864215e-05, 6.677767e-06, 
    3.02125e-06, 1.086349e-06, 1.568551e-06, 1.117854e-06, 1.202373e-06, 
    1.907597e-06, 2.830702e-06, 4.441009e-06, 7.927294e-06, 1.408851e-05,
  1.037417e-05, 5.223651e-06, 1.089607e-06, 1.840369e-06, 1.871359e-06, 
    3.1431e-06, 3.306606e-06, 1.790352e-06, 1.655179e-06, 1.244997e-06, 
    1.637978e-06, 2.002346e-06, 2.057684e-06, 1.515947e-06, 1.329775e-06,
  4.966552e-06, 2.419493e-06, 9.848313e-07, 1.197218e-06, 1.810503e-06, 
    2.730501e-06, 3.155516e-06, 2.280835e-06, 1.340712e-06, 6.121189e-07, 
    7.562411e-07, 1.174018e-06, 1.358728e-06, 6.756191e-07, 6.077585e-07,
  9.869738e-06, 2.563723e-06, 1.752074e-06, 1.734649e-06, 6.261181e-07, 
    2.110878e-06, 2.951625e-06, 8.628619e-06, 9.479334e-06, 2.594601e-06, 
    9.041263e-07, 1.404319e-06, 6.910819e-07, 3.300496e-07, 5.741829e-07,
  1.836387e-05, 1.464449e-05, 1.084703e-05, 3.725003e-06, 6.697519e-06, 
    5.532411e-06, 4.401249e-06, 8.19414e-06, 8.960184e-06, 9.577771e-06, 
    7.197315e-06, 3.178608e-06, 2.018705e-06, 2.881469e-06, 1.943898e-06,
  2.335363e-05, 1.74718e-05, 1.432307e-05, 9.898404e-06, 6.59879e-06, 
    1.034265e-05, 5.831996e-06, 2.422272e-06, 6.431058e-06, 1.650575e-05, 
    1.673008e-05, 1.149776e-05, 8.559875e-06, 5.90938e-06, 5.006256e-06,
  2.587642e-05, 1.951905e-05, 1.601471e-05, 1.336233e-05, 8.883638e-06, 
    8.191531e-06, 1.200315e-05, 1.975838e-05, 2.924082e-05, 2.813866e-05, 
    2.016764e-05, 1.65841e-05, 1.408708e-05, 1.084733e-05, 8.287136e-06,
  2.806521e-05, 2.64901e-05, 2.181145e-05, 2.044863e-05, 1.516905e-05, 
    9.457375e-06, 1.001383e-05, 1.761366e-05, 2.451482e-05, 2.436516e-05, 
    2.316776e-05, 2.150528e-05, 1.801324e-05, 1.436975e-05, 1.06376e-05,
  3.415694e-05, 2.887066e-05, 1.878901e-05, 1.972972e-05, 1.689345e-05, 
    1.069989e-05, 9.166148e-06, 1.03574e-05, 1.464694e-05, 1.736564e-05, 
    2.208761e-05, 2.330075e-05, 2.118765e-05, 1.759571e-05, 1.335048e-05,
  3.657789e-05, 2.274739e-05, 2.299594e-05, 1.669717e-05, 1.436694e-05, 
    1.022549e-05, 7.240347e-06, 3.328927e-06, 6.573459e-06, 1.143655e-05, 
    1.784145e-05, 2.347145e-05, 2.259819e-05, 2.088569e-05, 1.839794e-05,
  2.549213e-05, 1.834999e-05, 1.372072e-05, 1.132664e-05, 9.381365e-06, 
    6.635712e-06, 9.179916e-07, 3.938805e-06, 3.641198e-06, 4.107123e-06, 
    1.030321e-05, 1.834849e-05, 2.320004e-05, 2.269155e-05, 2.296344e-05,
  3.031824e-06, 2.933662e-06, 5.595495e-06, 4.657883e-06, 6.380658e-07, 
    2.451401e-06, 1.764407e-06, 1.549201e-06, 1.189145e-06, 1.020952e-06, 
    6.553028e-07, 1.209138e-06, 2.293415e-06, 3.576677e-06, 1.212976e-05,
  5.19617e-07, 3.414178e-07, 3.718049e-06, 2.828177e-06, 1.379741e-06, 
    1.877263e-06, 2.315551e-06, 1.121912e-06, 1.134381e-06, 7.070686e-07, 
    5.315616e-07, 7.185871e-07, 1.598149e-06, 2.534093e-06, 7.964442e-06,
  8.513694e-06, 1.50441e-06, 1.321666e-06, 5.773779e-06, 2.790356e-06, 
    6.519353e-07, 1.427638e-06, 4.693366e-06, 5.122143e-06, 1.897854e-06, 
    9.723968e-07, 7.580389e-07, 9.246012e-07, 3.674612e-06, 6.890335e-06,
  2.354956e-05, 2.429684e-05, 1.231774e-05, 7.273635e-06, 8.68393e-06, 
    5.216858e-06, 2.542226e-06, 3.384e-06, 4.54139e-06, 3.237654e-06, 
    2.994757e-06, 1.637432e-06, 9.371807e-07, 2.955646e-06, 4.940441e-06,
  2.634454e-05, 2.731902e-05, 2.193062e-05, 1.036776e-05, 8.757954e-06, 
    8.9788e-06, 6.236626e-06, 1.576643e-06, 4.485081e-06, 3.656542e-06, 
    2.949774e-06, 1.822088e-06, 1.808173e-06, 1.693477e-06, 3.439902e-06,
  3.158868e-05, 2.081706e-05, 2.149045e-05, 1.829165e-05, 1.424295e-05, 
    8.105604e-06, 9.77303e-06, 1.095963e-05, 1.302269e-05, 9.554073e-06, 
    1.982322e-06, 6.990244e-07, 2.200479e-06, 1.337688e-06, 2.139734e-06,
  2.57734e-05, 3.086436e-05, 1.934433e-05, 2.308184e-05, 2.140263e-05, 
    9.95026e-06, 7.782482e-06, 1.04761e-05, 1.47868e-05, 1.094759e-05, 
    3.59576e-06, 1.753938e-06, 2.995803e-07, 2.984402e-07, 1.333208e-06,
  2.819819e-05, 1.91967e-05, 2.356379e-05, 1.724796e-05, 1.549885e-05, 
    1.134525e-05, 7.611474e-06, 5.204551e-06, 6.580946e-06, 1.017314e-05, 
    8.887755e-06, 3.374944e-06, 1.699321e-06, 1.49128e-06, 5.742854e-07,
  2.409309e-05, 1.893252e-05, 1.237677e-05, 1.022907e-05, 1.100531e-05, 
    9.130623e-06, 8.341334e-06, 4.155506e-06, 6.438552e-06, 1.118064e-05, 
    1.187264e-05, 9.324905e-06, 4.979966e-06, 2.779455e-06, 2.247607e-06,
  1.624958e-05, 1.251341e-05, 1.176749e-05, 6.665174e-06, 4.967611e-06, 
    5.519866e-06, 6.29837e-06, 7.938393e-06, 8.115549e-06, 7.680006e-06, 
    9.873776e-06, 1.232066e-05, 9.883292e-06, 6.932671e-06, 5.175779e-06,
  2.127666e-06, 1.491698e-06, 2.210309e-06, 2.843156e-06, 6.470639e-07, 
    9.822237e-07, 1.016336e-06, 1.757282e-06, 1.75382e-06, 1.382677e-06, 
    1.654525e-06, 1.67525e-06, 1.407593e-06, 7.831504e-07, 1.222631e-06,
  2.642817e-07, 2.761549e-07, 2.826359e-06, 2.979736e-06, 1.33406e-06, 
    8.772185e-07, 4.699261e-07, 8.060669e-07, 9.248104e-07, 1.886758e-06, 
    2.00992e-06, 1.734768e-06, 1.885357e-06, 1.218886e-06, 1.357243e-06,
  4.73204e-06, 8.657358e-07, 5.139525e-07, 3.677617e-06, 3.289098e-06, 
    1.44594e-06, 2.820031e-07, 1.39488e-06, 1.631928e-06, 6.523464e-07, 
    9.726308e-07, 1.670331e-06, 2.001053e-06, 2.386467e-06, 2.102225e-06,
  2.12238e-05, 1.67713e-05, 1.022043e-05, 1.742943e-06, 6.915172e-06, 
    2.788783e-06, 6.314569e-07, 1.110657e-06, 2.766114e-06, 2.522109e-06, 
    1.727508e-06, 2.080569e-06, 2.069154e-06, 3.433987e-06, 3.37548e-06,
  2.402893e-05, 2.163293e-05, 1.920456e-05, 6.801034e-06, 5.57798e-06, 
    6.638588e-06, 5.302069e-06, 5.452933e-07, 3.248362e-07, 2.980783e-06, 
    2.728302e-06, 1.268828e-06, 1.875953e-06, 3.0271e-06, 4.594582e-06,
  2.652872e-05, 2.33165e-05, 2.283241e-05, 1.591398e-05, 1.449091e-05, 
    8.025558e-06, 8.986673e-06, 6.084706e-06, 5.256754e-06, 5.92576e-06, 
    2.9678e-06, 2.102873e-06, 1.012753e-06, 3.13785e-06, 5.594371e-06,
  2.974565e-05, 3.02163e-05, 2.779469e-05, 2.72184e-05, 2.318653e-05, 
    9.192082e-06, 8.604084e-06, 7.365986e-06, 7.034303e-06, 5.747999e-06, 
    3.169106e-06, 2.034967e-06, 1.021119e-06, 1.557656e-06, 6.302173e-06,
  3.209148e-05, 3.002474e-05, 2.987702e-05, 1.652072e-05, 1.598648e-05, 
    8.869193e-06, 8.450893e-06, 8.149206e-06, 7.734687e-06, 6.052152e-06, 
    4.9507e-06, 2.234332e-06, 1.995417e-06, 2.478942e-06, 6.015149e-06,
  2.918527e-05, 1.956466e-05, 1.07687e-05, 8.26741e-06, 6.998775e-06, 
    4.829887e-06, 5.968186e-06, 9.448709e-06, 9.775013e-06, 8.909926e-06, 
    6.791229e-06, 3.836899e-06, 1.871363e-06, 2.005161e-06, 4.848538e-06,
  1.984759e-05, 1.009382e-05, 4.556801e-06, 3.176567e-06, 2.211771e-06, 
    2.806811e-06, 3.845162e-06, 9.283475e-06, 8.329998e-06, 7.369511e-06, 
    6.215758e-06, 5.852249e-06, 3.965003e-06, 2.454553e-06, 2.897894e-06,
  2.213573e-06, 2.067568e-06, 7.204149e-07, 7.515467e-07, 1.173558e-06, 
    9.697495e-07, 8.014809e-07, 6.343073e-07, 8.986715e-07, 1.980124e-06, 
    2.580897e-06, 2.951725e-06, 2.730782e-06, 2.23495e-06, 1.295311e-06,
  6.789421e-07, 1.329427e-07, 8.17214e-07, 5.32371e-07, 7.086199e-07, 
    5.220808e-07, 4.453571e-07, 7.62159e-07, 5.99008e-07, 1.599047e-06, 
    2.36845e-06, 3.546369e-06, 3.4845e-06, 3.116416e-06, 1.511272e-06,
  3.332791e-06, 1.626436e-07, 1.920225e-06, 9.924978e-07, 1.073941e-06, 
    7.729652e-07, 2.111399e-07, 4.21218e-07, 4.010832e-07, 4.722034e-07, 
    1.235279e-06, 2.494958e-06, 2.830952e-06, 2.768413e-06, 2.315957e-06,
  1.37533e-05, 1.118841e-05, 4.426928e-06, 1.472192e-06, 5.606419e-06, 
    1.63128e-06, 1.718231e-07, 1.969219e-07, 2.68458e-07, 5.878442e-07, 
    1.45589e-06, 2.093212e-06, 2.410064e-06, 3.249468e-06, 3.168449e-06,
  1.790215e-05, 1.811551e-05, 1.406684e-05, 3.597919e-06, 2.426129e-06, 
    3.823049e-06, 2.79311e-06, 4.384274e-07, 3.251406e-07, 1.802535e-06, 
    2.903221e-06, 2.076898e-06, 1.985946e-06, 2.429749e-06, 3.879693e-06,
  1.528511e-05, 1.714566e-05, 1.131189e-05, 8.431703e-06, 6.019888e-06, 
    4.07928e-06, 5.078743e-06, 4.129086e-06, 2.852899e-06, 2.631132e-06, 
    1.730742e-06, 1.348245e-06, 8.213319e-07, 3.404058e-06, 3.49776e-06,
  1.308645e-05, 1.797787e-05, 1.691305e-05, 1.673264e-05, 1.575873e-05, 
    3.96159e-06, 3.626669e-06, 3.798298e-06, 3.539248e-06, 2.144847e-06, 
    8.586729e-07, 7.002837e-07, 6.573763e-07, 1.93639e-06, 3.182102e-06,
  1.573968e-05, 1.744213e-05, 1.98479e-05, 1.58414e-05, 1.053238e-05, 
    3.313136e-06, 2.623521e-06, 2.710925e-06, 2.702079e-06, 2.049739e-06, 
    1.172872e-06, 8.330847e-07, 7.907828e-07, 1.900642e-06, 3.283298e-06,
  1.296856e-05, 1.427695e-05, 1.187815e-05, 6.565706e-06, 2.129818e-06, 
    2.312142e-06, 3.551499e-06, 3.738761e-06, 3.007281e-06, 2.431161e-06, 
    1.841431e-06, 1.444264e-06, 1.264558e-06, 2.276696e-06, 3.675862e-06,
  9.192044e-06, 4.430045e-06, 1.561775e-06, 2.0613e-06, 4.168063e-06, 
    5.483426e-06, 7.551071e-06, 1.148819e-05, 6.720082e-06, 2.517126e-06, 
    1.491383e-06, 1.547162e-06, 1.688042e-06, 2.483654e-06, 3.787181e-06,
  1.208575e-07, 4.032256e-07, 7.988679e-07, 7.013358e-07, 3.990068e-07, 
    6.522548e-07, 6.60233e-07, 6.213457e-07, 3.188078e-07, 7.275413e-07, 
    3.616136e-06, 9.714195e-06, 1.820508e-05, 2.371835e-05, 2.849306e-05,
  1.008418e-09, 1.172534e-07, 6.482917e-08, 4.239405e-08, 1.445942e-07, 
    4.539877e-07, 6.013208e-07, 7.883549e-07, 8.201721e-07, 7.01423e-07, 
    7.20745e-07, 1.607078e-06, 3.38047e-06, 6.528724e-06, 1.310444e-05,
  7.822359e-07, 2.028556e-08, 2.686908e-07, 3.338853e-07, 3.159661e-07, 
    1.602955e-06, 7.586546e-07, 5.285083e-07, 6.543796e-07, 3.439291e-07, 
    5.315486e-07, 1.314691e-06, 2.232676e-06, 2.08331e-06, 3.556703e-06,
  7.393344e-06, 3.963489e-06, 2.401912e-06, 2.614953e-06, 4.498228e-06, 
    6.488928e-06, 9.601748e-06, 6.521206e-06, 4.61145e-06, 5.51766e-06, 
    5.036363e-06, 2.174571e-06, 1.087148e-06, 9.844539e-07, 1.472091e-06,
  7.949875e-06, 8.473869e-06, 1.601866e-05, 5.116159e-06, 8.759104e-06, 
    1.681481e-05, 2.223554e-05, 2.111947e-05, 1.031482e-05, 8.357851e-06, 
    1.660607e-05, 1.134877e-05, 4.227488e-06, 2.689186e-06, 2.737804e-06,
  1.573487e-05, 1.877009e-05, 2.032089e-05, 9.8597e-06, 1.294573e-05, 
    2.060454e-05, 3.405183e-05, 3.814528e-05, 2.69999e-05, 1.977953e-05, 
    1.644714e-05, 1.188854e-05, 7.94899e-06, 7.221995e-06, 5.336737e-06,
  3.760064e-05, 4.836873e-05, 2.696183e-05, 1.507105e-05, 2.364936e-05, 
    2.169555e-05, 2.951597e-05, 3.147883e-05, 2.681516e-05, 1.881533e-05, 
    1.478008e-05, 1.203901e-05, 1.205224e-05, 1.166489e-05, 8.845827e-06,
  6.268493e-05, 4.086014e-05, 2.924143e-05, 2.845631e-05, 3.054038e-05, 
    2.655625e-05, 2.481787e-05, 2.2607e-05, 1.916257e-05, 1.638137e-05, 
    1.514842e-05, 1.395273e-05, 1.336436e-05, 1.217759e-05, 9.338996e-06,
  5.115058e-05, 3.200006e-05, 3.089594e-05, 2.783715e-05, 2.20804e-05, 
    2.242987e-05, 2.325457e-05, 2.084364e-05, 1.810271e-05, 1.438095e-05, 
    1.253625e-05, 1.144619e-05, 1.268719e-05, 1.139237e-05, 8.40762e-06,
  2.467376e-05, 1.522089e-05, 1.551134e-05, 2.060487e-05, 2.097989e-05, 
    1.629154e-05, 1.594637e-05, 2.182606e-05, 1.980596e-05, 1.347328e-05, 
    1.289846e-05, 1.218126e-05, 1.075808e-05, 1.037779e-05, 8.041709e-06,
  1.248813e-07, 6.986331e-07, 1.692257e-06, 1.856714e-06, 9.959947e-07, 
    1.812949e-06, 8.020675e-07, 3.15631e-07, 2.486522e-07, 2.19038e-07, 
    1.402101e-07, 1.694663e-07, 2.945862e-07, 4.498586e-07, 4.236643e-07,
  1.217088e-08, 3.572632e-08, 7.24375e-07, 2.108116e-06, 1.010094e-06, 
    2.688542e-06, 1.135773e-06, 1.654247e-06, 1.367513e-06, 1.000646e-06, 
    8.906674e-07, 7.19136e-07, 3.997027e-07, 6.179675e-07, 4.564822e-07,
  5.187848e-07, 9.933014e-08, 1.346566e-06, 6.27906e-06, 8.008457e-06, 
    1.548221e-05, 4.106656e-06, 8.898815e-06, 1.320396e-05, 1.079847e-05, 
    8.503763e-06, 8.469654e-06, 7.710201e-06, 4.752413e-06, 4.251252e-06,
  1.599092e-07, 3.643712e-06, 4.133853e-06, 1.047465e-05, 1.179667e-05, 
    1.013913e-05, 1.166701e-05, 3.800349e-06, 5.795989e-06, 1.710112e-05, 
    1.798751e-05, 1.303011e-05, 1.171578e-05, 1.177518e-05, 1.106349e-05,
  1.50438e-06, 6.541744e-06, 3.775845e-05, 1.3656e-05, 6.511764e-06, 
    8.112595e-06, 1.075828e-05, 1.178481e-05, 5.601099e-06, 6.88696e-06, 
    9.326823e-06, 7.877062e-06, 9.849963e-06, 1.145472e-05, 1.279621e-05,
  8.580659e-06, 4.491996e-05, 2.003376e-05, 9.868859e-06, 3.484829e-06, 
    9.302657e-06, 2.521649e-05, 2.222795e-05, 1.375169e-05, 7.003605e-06, 
    2.549688e-06, 2.969858e-06, 3.450701e-06, 6.062195e-06, 1.160766e-05,
  7.296288e-05, 3.776253e-05, 1.945438e-05, 1.089955e-05, 1.742854e-05, 
    2.070434e-05, 2.082797e-05, 1.047325e-05, 4.663524e-06, 2.073678e-06, 
    5.822682e-07, 3.403713e-07, 1.03722e-06, 1.627765e-06, 4.55058e-06,
  5.147436e-05, 2.927658e-05, 2.130247e-05, 2.180288e-05, 2.458381e-05, 
    1.291947e-05, 2.483252e-06, 1.389254e-06, 2.148701e-06, 1.059223e-06, 
    1.049898e-06, 1.050521e-06, 2.185791e-06, 2.923127e-06, 4.235852e-06,
  3.031698e-05, 2.585314e-05, 2.930941e-05, 2.015456e-05, 1.285967e-05, 
    3.325459e-06, 1.372301e-06, 2.821933e-06, 2.971228e-06, 7.793284e-06, 
    2.385233e-06, 2.557913e-06, 3.799994e-06, 4.813322e-06, 4.612807e-06,
  2.023492e-05, 1.486777e-05, 1.601154e-05, 1.351638e-05, 2.520957e-06, 
    1.47461e-06, 4.007647e-06, 8.057581e-06, 8.667391e-06, 4.417219e-06, 
    4.317028e-06, 3.600794e-06, 2.937313e-06, 3.52487e-06, 4.701229e-06,
  1.80594e-07, 2.053463e-08, 7.284962e-10, 4.767139e-09, 1.271713e-06, 
    2.539312e-06, 3.866496e-06, 1.496927e-06, 2.540087e-06, 3.001475e-06, 
    1.942126e-06, 1.512177e-06, 1.524177e-06, 1.021611e-06, 9.43807e-07,
  7.177132e-08, 8.087165e-09, 9.271001e-09, 1.958687e-07, 1.22026e-06, 
    5.311316e-06, 4.343138e-06, 7.183871e-07, 1.259661e-06, 3.147119e-06, 
    2.999526e-06, 2.955589e-06, 2.688704e-06, 2.565107e-06, 1.731896e-06,
  2.195624e-09, 3.776736e-10, 6.065251e-08, 3.340673e-06, 1.079772e-05, 
    1.829059e-05, 2.368498e-06, 2.452187e-06, 3.269849e-06, 4.479722e-06, 
    5.131011e-06, 4.133414e-06, 5.233893e-06, 4.422926e-06, 3.229686e-06,
  2.224176e-10, 4.058815e-08, 4.009165e-06, 2.514197e-05, 2.546623e-05, 
    5.360716e-06, 4.366052e-06, 2.111572e-06, 7.597134e-06, 1.263041e-05, 
    1.047231e-05, 8.043347e-06, 7.755868e-06, 6.98678e-06, 7.067491e-06,
  2.916179e-08, 3.06054e-06, 3.147623e-05, 3.76061e-05, 1.08273e-05, 
    1.386404e-06, 1.275843e-06, 3.332001e-06, 3.606139e-06, 1.089086e-05, 
    1.43848e-05, 1.056448e-05, 1.008902e-05, 9.828463e-06, 1.031196e-05,
  2.240929e-06, 3.250428e-05, 3.524979e-05, 1.044008e-05, 1.08546e-06, 
    2.867964e-07, 2.967988e-07, 1.781188e-06, 2.601633e-06, 2.396661e-06, 
    3.780905e-06, 5.51287e-06, 5.937238e-06, 6.988422e-06, 1.013903e-05,
  5.070297e-05, 3.409633e-05, 1.588854e-05, 6.08382e-06, 9.946469e-06, 
    1.033721e-06, 5.075067e-07, 7.183899e-07, 5.487612e-07, 5.8805e-07, 
    6.427246e-07, 9.961443e-07, 9.964291e-07, 1.176553e-06, 1.412371e-06,
  3.713957e-05, 1.522254e-05, 6.739696e-06, 7.936998e-06, 9.245709e-06, 
    1.639172e-06, 9.058567e-07, 9.174428e-07, 9.435637e-07, 7.468592e-07, 
    6.563514e-07, 1.688224e-06, 1.064976e-06, 8.488569e-07, 1.834775e-06,
  2.202958e-05, 4.749607e-06, 9.295182e-06, 8.023248e-06, 4.478879e-06, 
    2.510673e-06, 2.332137e-06, 3.122876e-06, 4.269317e-06, 4.026739e-06, 
    3.46501e-07, 2.640098e-07, 2.896388e-06, 2.000829e-06, 1.905298e-06,
  1.056164e-05, 3.300258e-06, 7.077395e-06, 2.58608e-06, 1.599519e-06, 
    3.376234e-06, 4.31516e-06, 1.176594e-05, 9.217517e-06, 1.908047e-06, 
    2.820715e-06, 4.198562e-07, 7.956857e-07, 3.433741e-06, 1.989288e-06,
  2.685793e-06, 1.782934e-06, 1.078179e-06, 6.899973e-07, 5.420082e-07, 
    5.610473e-07, 8.058383e-07, 1.262516e-06, 8.478331e-07, 4.407702e-07, 
    7.256671e-07, 4.991812e-07, 5.21202e-07, 5.71717e-07, 9.812269e-07,
  3.411124e-06, 2.515136e-06, 1.770924e-06, 1.361233e-06, 1.092209e-06, 
    1.865516e-06, 2.916063e-06, 1.966137e-06, 8.563865e-07, 9.515333e-07, 
    7.026792e-07, 1.677631e-07, 3.573781e-07, 1.767726e-06, 1.667915e-06,
  3.313019e-06, 3.458553e-06, 2.688375e-06, 2.397775e-06, 2.818067e-06, 
    8.825654e-06, 4.124186e-06, 5.498396e-06, 2.498391e-06, 8.409432e-07, 
    2.823847e-07, 2.297231e-07, 7.480983e-07, 8.776882e-07, 1.438055e-06,
  1.02271e-05, 5.855537e-06, 4.348386e-06, 4.612282e-06, 8.828351e-06, 
    8.601313e-06, 6.580472e-06, 3.114558e-06, 2.093347e-06, 6.829973e-07, 
    4.170571e-07, 7.542821e-07, 7.925127e-07, 9.28395e-07, 1.547487e-06,
  1.261516e-05, 1.089884e-05, 1.291016e-05, 7.624131e-06, 1.125504e-05, 
    7.960832e-06, 2.874835e-06, 5.708402e-06, 1.1887e-06, 6.8548e-08, 
    1.590269e-06, 1.064126e-06, 7.63423e-07, 1.40419e-06, 2.883637e-06,
  8.940412e-06, 1.006738e-05, 1.039383e-05, 1.066602e-05, 7.987232e-06, 
    5.183768e-06, 3.795188e-06, 2.118858e-06, 6.893283e-07, 8.769333e-07, 
    1.058742e-06, 1.463893e-06, 1.80645e-06, 1.798488e-06, 1.906361e-06,
  4.057249e-06, 1.437272e-05, 2.005262e-05, 1.357086e-05, 7.203781e-06, 
    3.144851e-06, 3.947948e-06, 2.846255e-06, 1.710971e-06, 1.347973e-06, 
    1.324574e-06, 2.554018e-06, 2.406281e-06, 2.1652e-06, 1.909075e-06,
  1.785454e-05, 1.978271e-05, 1.615496e-05, 7.606292e-06, 8.691098e-06, 
    6.630974e-06, 4.232588e-06, 1.807252e-06, 1.78078e-06, 1.536439e-06, 
    1.452721e-06, 2.655294e-06, 1.950684e-06, 1.533247e-06, 1.798178e-06,
  3.098622e-05, 1.986832e-05, 9.374673e-06, 1.446184e-05, 1.685255e-05, 
    8.859904e-06, 2.721404e-06, 1.929062e-06, 3.288076e-06, 2.062718e-06, 
    1.045978e-06, 1.026179e-06, 1.371295e-06, 1.888801e-06, 1.182879e-06,
  1.78484e-05, 1.95914e-05, 3.10087e-05, 3.282864e-05, 1.745862e-05, 
    4.266079e-06, 1.980388e-06, 5.861489e-06, 7.066651e-06, 1.78932e-06, 
    2.016384e-06, 3.802206e-07, 8.17496e-07, 1.578522e-06, 1.577511e-06,
  2.229675e-05, 1.806293e-05, 1.238953e-05, 6.271703e-06, 2.414155e-06, 
    1.215607e-06, 1.07038e-06, 1.070831e-06, 9.894637e-07, 1.023375e-06, 
    8.722344e-07, 1.203922e-06, 1.573736e-06, 1.937693e-06, 1.784025e-06,
  1.593504e-05, 1.700456e-05, 1.183503e-05, 6.989644e-06, 3.564628e-06, 
    1.964827e-06, 1.578303e-06, 1.618991e-06, 1.58744e-06, 1.903233e-06, 
    2.667989e-06, 2.890205e-06, 2.679538e-06, 3.329167e-06, 2.602107e-06,
  1.229424e-05, 1.404041e-05, 1.097461e-05, 6.601852e-06, 3.607694e-06, 
    4.043823e-06, 2.57701e-06, 2.768309e-06, 3.152019e-06, 2.873457e-06, 
    2.98838e-06, 3.498994e-06, 3.080626e-06, 3.06775e-06, 4.393512e-06,
  1.454092e-05, 1.557934e-05, 1.416321e-05, 7.648295e-06, 3.940404e-06, 
    3.176742e-06, 4.730146e-06, 3.845633e-06, 4.263049e-06, 4.211444e-06, 
    4.472868e-06, 4.094562e-06, 4.190538e-06, 5.311122e-06, 8.777375e-06,
  1.631286e-05, 1.554409e-05, 1.518412e-05, 1.009629e-05, 5.518741e-06, 
    4.44222e-06, 4.045267e-06, 5.116954e-06, 4.377687e-06, 3.86019e-06, 
    6.011271e-06, 5.442946e-06, 4.904917e-06, 7.779627e-06, 1.116968e-05,
  1.189253e-05, 1.726224e-05, 1.808169e-05, 1.101739e-05, 8.386477e-06, 
    5.500256e-06, 5.701416e-06, 6.010598e-06, 4.035692e-06, 6.808547e-06, 
    8.33687e-06, 6.133911e-06, 6.921141e-06, 9.720386e-06, 9.776637e-06,
  1.046815e-05, 1.610478e-05, 1.827963e-05, 1.440013e-05, 1.301857e-05, 
    6.243121e-06, 6.887706e-06, 1.25474e-05, 1.614517e-05, 1.296065e-05, 
    9.048308e-06, 8.558403e-06, 9.478555e-06, 7.499088e-06, 3.911407e-06,
  1.423629e-05, 1.59529e-05, 1.4574e-05, 1.444978e-05, 1.587191e-05, 
    7.178458e-06, 1.222021e-05, 1.81579e-05, 1.884957e-05, 1.622518e-05, 
    1.403671e-05, 1.13627e-05, 5.666949e-06, 2.358719e-06, 1.707372e-06,
  1.430404e-05, 1.765369e-05, 1.775783e-05, 1.362731e-05, 7.727194e-06, 
    1.729421e-05, 2.664163e-05, 2.827206e-05, 2.213174e-05, 1.44398e-05, 
    7.155728e-06, 2.706602e-06, 1.742475e-06, 1.05106e-06, 9.786324e-07,
  1.563852e-05, 2.78672e-05, 1.482931e-05, 1.749023e-05, 2.996789e-05, 
    3.873275e-05, 3.277592e-05, 1.837437e-05, 8.47854e-06, 2.089538e-06, 
    7.046715e-07, 6.89121e-07, 4.383204e-07, 1.254055e-06, 2.499214e-06,
  2.357137e-06, 6.770687e-06, 1.370914e-05, 1.506099e-05, 1.296124e-05, 
    8.541745e-06, 6.485814e-06, 5.455179e-06, 5.57744e-06, 7.547234e-06, 
    7.594253e-06, 5.960915e-06, 4.120192e-06, 3.366984e-06, 3.070883e-06,
  4.835043e-06, 9.88687e-06, 1.887682e-05, 2.458689e-05, 2.43693e-05, 
    1.597134e-05, 1.089123e-05, 1.069841e-05, 9.57825e-06, 9.929677e-06, 
    8.408115e-06, 7.088377e-06, 4.733559e-06, 3.640385e-06, 2.942863e-06,
  1.066835e-05, 8.026489e-06, 1.969154e-05, 3.043207e-05, 3.190414e-05, 
    2.066354e-05, 1.748518e-05, 2.054906e-05, 1.741733e-05, 1.137003e-05, 
    7.815408e-06, 7.122303e-06, 5.950579e-06, 4.365609e-06, 3.560063e-06,
  1.931941e-05, 1.432774e-05, 2.687361e-05, 3.280207e-05, 3.607689e-05, 
    2.777914e-05, 2.170529e-05, 2.081443e-05, 1.706914e-05, 1.321958e-05, 
    1.002122e-05, 8.190933e-06, 7.639231e-06, 6.779766e-06, 5.593988e-06,
  1.693828e-05, 1.380663e-05, 2.400543e-05, 3.744852e-05, 3.632809e-05, 
    3.144824e-05, 2.190977e-05, 9.262796e-06, 7.929289e-06, 1.090261e-05, 
    1.35968e-05, 1.004323e-05, 8.728556e-06, 7.288558e-06, 6.666672e-06,
  1.911411e-05, 1.592975e-05, 1.958639e-05, 3.68096e-05, 3.65427e-05, 
    2.368558e-05, 1.69529e-05, 1.098328e-05, 8.438401e-06, 8.302274e-06, 
    7.861698e-06, 7.053489e-06, 6.733959e-06, 6.53976e-06, 7.843531e-06,
  2.694474e-05, 2.310234e-05, 2.768668e-05, 3.771338e-05, 3.644886e-05, 
    1.850991e-05, 8.997544e-06, 7.106433e-06, 5.698098e-06, 4.241961e-06, 
    4.022028e-06, 4.367607e-06, 4.871067e-06, 6.193531e-06, 9.545039e-06,
  4.272882e-05, 3.513519e-05, 3.481135e-05, 3.698807e-05, 3.168832e-05, 
    1.637493e-05, 7.011251e-06, 5.007201e-06, 3.77187e-06, 4.068133e-06, 
    4.554726e-06, 7.649685e-06, 1.042263e-05, 9.823353e-06, 7.897075e-06,
  4.091962e-05, 4.613561e-05, 3.594806e-05, 2.629157e-05, 1.842831e-05, 
    1.398514e-05, 1.124266e-05, 1.043277e-05, 9.877552e-06, 8.944126e-06, 
    5.487955e-06, 2.916468e-06, 1.955952e-06, 8.250584e-07, 5.364593e-07,
  2.980238e-05, 1.842049e-05, 1.249301e-05, 7.852163e-06, 9.556576e-06, 
    9.546022e-06, 5.661635e-06, 5.988201e-06, 4.011185e-06, 8.52552e-07, 
    4.43657e-07, 3.815752e-07, 2.537111e-07, 2.168471e-07, 4.061581e-07,
  4.909546e-06, 3.405466e-06, 6.015767e-06, 8.085258e-06, 8.685886e-06, 
    9.358845e-06, 8.947199e-06, 9.63804e-06, 1.445951e-05, 1.523138e-05, 
    7.9204e-06, 9.325228e-06, 1.209241e-05, 1.264227e-05, 1.66668e-05,
  2.380655e-06, 3.104394e-06, 5.204581e-06, 6.503514e-06, 9.207677e-06, 
    7.787364e-06, 8.654167e-06, 1.247453e-05, 1.569669e-05, 1.879325e-05, 
    1.550862e-05, 1.513965e-05, 1.35654e-05, 1.262273e-05, 1.35675e-05,
  9.179865e-06, 4.660564e-06, 5.891153e-06, 6.675009e-06, 9.398344e-06, 
    1.423284e-05, 7.58787e-06, 1.493324e-05, 1.395308e-05, 1.431522e-05, 
    1.421766e-05, 1.414393e-05, 1.451593e-05, 1.470729e-05, 1.598787e-05,
  2.016406e-05, 2.620385e-05, 2.245969e-05, 1.377953e-05, 1.329553e-05, 
    1.348808e-05, 1.250149e-05, 1.586084e-05, 1.556388e-05, 1.257019e-05, 
    1.229451e-05, 1.317211e-05, 1.423787e-05, 1.742431e-05, 1.666613e-05,
  2.934751e-05, 3.030226e-05, 3.026717e-05, 2.112452e-05, 1.472341e-05, 
    1.397412e-05, 1.09987e-05, 9.497604e-06, 9.903657e-06, 1.565081e-05, 
    1.690704e-05, 1.450632e-05, 1.499709e-05, 1.747352e-05, 1.827471e-05,
  3.515164e-05, 3.081218e-05, 2.85897e-05, 2.203028e-05, 1.357792e-05, 
    1.121986e-05, 1.175549e-05, 1.634201e-05, 2.465887e-05, 2.72171e-05, 
    2.526472e-05, 2.553394e-05, 2.464514e-05, 2.42728e-05, 2.552467e-05,
  3.461646e-05, 3.463996e-05, 3.246075e-05, 2.528125e-05, 1.483736e-05, 
    7.166952e-06, 6.97308e-06, 1.155051e-05, 1.882808e-05, 2.215541e-05, 
    2.526158e-05, 2.80041e-05, 2.667534e-05, 2.511445e-05, 2.501554e-05,
  3.051609e-05, 3.091655e-05, 2.685323e-05, 2.154522e-05, 1.481579e-05, 
    5.774513e-06, 4.531724e-06, 4.274327e-06, 5.097461e-06, 7.861648e-06, 
    1.061615e-05, 1.251236e-05, 1.230348e-05, 1.116292e-05, 1.051271e-05,
  3.174938e-05, 2.451474e-05, 1.765125e-05, 8.807538e-06, 3.215458e-06, 
    1.916248e-06, 2.410724e-06, 2.403719e-06, 2.077795e-06, 9.681193e-07, 
    4.131875e-07, 3.570376e-07, 4.725566e-07, 3.665193e-07, 3.696804e-07,
  2.688095e-05, 2.120903e-05, 1.416987e-05, 3.944517e-06, 1.418146e-06, 
    1.36502e-06, 1.287233e-06, 2.22265e-06, 1.750496e-06, 3.242727e-07, 
    4.325672e-07, 4.526933e-07, 3.60305e-07, 2.323158e-07, 2.141756e-07,
  3.998788e-07, 6.963038e-08, 3.674177e-08, 7.157196e-08, 4.111437e-07, 
    1.791936e-06, 4.139951e-06, 3.452632e-06, 4.090749e-06, 9.055969e-06, 
    9.816889e-06, 1.329898e-05, 1.777081e-05, 1.977997e-05, 1.711927e-05,
  9.722713e-08, 1.821511e-08, 7.167203e-09, 2.234615e-07, 1.993144e-07, 
    5.916309e-07, 1.316063e-06, 1.675597e-06, 8.682349e-07, 2.979599e-06, 
    8.977568e-06, 1.508627e-05, 1.906269e-05, 1.896363e-05, 1.432491e-05,
  6.114923e-06, 1.836594e-07, 1.005445e-07, 6.059562e-07, 7.142229e-07, 
    5.10889e-06, 1.484119e-06, 1.962736e-06, 3.465372e-06, 4.066663e-06, 
    6.659467e-06, 1.0625e-05, 1.328531e-05, 1.585407e-05, 1.839682e-05,
  1.459387e-05, 1.282071e-05, 1.021314e-05, 3.222748e-06, 3.795857e-06, 
    5.530244e-06, 4.571159e-06, 7.343016e-07, 1.820295e-06, 5.026159e-06, 
    4.634129e-06, 5.917308e-06, 7.830048e-06, 1.227274e-05, 1.60426e-05,
  1.752058e-05, 1.32018e-05, 1.569916e-05, 8.468629e-06, 1.298882e-05, 
    1.157688e-05, 7.281296e-06, 1.599018e-06, 3.484447e-06, 4.400486e-06, 
    4.839403e-06, 4.535521e-06, 5.033768e-06, 5.849617e-06, 8.930686e-06,
  2.543651e-05, 1.094763e-05, 1.285109e-05, 2.312789e-05, 2.763908e-05, 
    2.11858e-05, 7.515304e-06, 3.346433e-06, 4.466824e-06, 5.241063e-06, 
    3.899541e-06, 5.153176e-06, 7.060192e-06, 8.93894e-06, 1.092814e-05,
  4.561491e-05, 3.148537e-05, 3.468828e-05, 5.678512e-05, 5.499419e-05, 
    1.088827e-05, 2.169524e-06, 2.352457e-06, 2.571505e-06, 2.325852e-06, 
    2.514665e-06, 3.240747e-06, 4.603381e-06, 7.19585e-06, 1.133592e-05,
  5.905917e-05, 5.666031e-05, 7.610414e-05, 7.586123e-05, 1.467651e-05, 
    1.475074e-06, 7.118794e-07, 1.280352e-06, 1.743521e-06, 2.211792e-06, 
    2.095132e-06, 1.358917e-06, 1.19686e-06, 2.145927e-06, 4.392459e-06,
  5.352266e-05, 5.870904e-05, 6.717681e-05, 2.595508e-05, 2.798153e-06, 
    7.971179e-07, 1.185024e-06, 1.456019e-06, 2.444524e-06, 3.407905e-06, 
    2.549235e-06, 1.081782e-06, 3.476506e-07, 4.107979e-07, 6.976858e-07,
  4.646806e-05, 4.094244e-05, 3.413262e-05, 1.002089e-05, 7.991576e-07, 
    1.056546e-06, 1.642215e-06, 3.710451e-06, 3.53861e-06, 2.593778e-06, 
    2.390609e-06, 1.435535e-06, 5.153219e-07, 2.551616e-07, 2.958951e-07,
  4.115419e-06, 4.509863e-06, 5.264014e-06, 5.220728e-06, 4.370555e-06, 
    3.741314e-06, 4.624622e-06, 5.649318e-06, 5.107532e-06, 4.649345e-06, 
    3.665195e-06, 2.497364e-06, 2.286863e-06, 2.294823e-06, 4.340702e-06,
  1.779456e-06, 2.074192e-06, 2.971874e-06, 4.15516e-06, 3.461752e-06, 
    2.542168e-06, 3.589937e-06, 4.109815e-06, 4.082977e-06, 2.974092e-06, 
    2.968075e-06, 4.538788e-06, 5.462869e-06, 6.976812e-06, 7.425596e-06,
  9.410035e-07, 3.365367e-06, 2.053925e-06, 2.723077e-06, 9.002674e-07, 
    2.091205e-06, 1.628823e-06, 3.662745e-06, 3.114402e-06, 3.74337e-06, 
    5.782893e-06, 9.8747e-06, 1.369723e-05, 1.595266e-05, 1.631466e-05,
  4.985486e-06, 6.191286e-06, 5.860712e-06, 4.477513e-06, 6.626279e-07, 
    4.197716e-07, 5.465154e-06, 8.646e-06, 1.277626e-05, 1.720442e-05, 
    1.581655e-05, 1.260884e-05, 1.139258e-05, 1.108014e-05, 1.048636e-05,
  1.689815e-05, 1.693712e-05, 1.956372e-05, 5.099536e-06, 3.755324e-06, 
    8.820569e-06, 1.58333e-05, 2.923606e-05, 1.734128e-05, 1.243366e-05, 
    9.956118e-06, 5.895695e-06, 4.377902e-06, 4.007692e-06, 4.497198e-06,
  3.335627e-05, 3.202609e-05, 3.536393e-05, 2.90359e-05, 2.905321e-05, 
    3.839867e-05, 3.528488e-05, 1.291379e-05, 3.982007e-06, 2.198185e-06, 
    1.692195e-06, 2.212261e-06, 2.609171e-06, 2.868915e-06, 2.497096e-06,
  5.323295e-05, 4.951038e-05, 3.673269e-05, 3.272396e-05, 2.269534e-05, 
    1.293157e-05, 3.7264e-06, 2.217595e-06, 1.251857e-06, 1.283711e-06, 
    2.253322e-06, 2.652329e-06, 2.07234e-06, 2.14846e-06, 2.045121e-06,
  4.054676e-05, 3.503322e-05, 2.178072e-05, 9.740887e-06, 3.900291e-06, 
    1.539585e-06, 9.043328e-07, 4.236316e-07, 1.045431e-06, 1.413401e-06, 
    1.536086e-06, 1.379464e-06, 8.331945e-07, 1.07897e-06, 1.35625e-06,
  2.156424e-05, 2.009707e-05, 9.755225e-06, 6.817098e-06, 2.721866e-06, 
    1.024218e-06, 5.31224e-07, 5.287101e-07, 1.027831e-06, 9.018125e-07, 
    9.735803e-07, 1.466101e-06, 2.482745e-06, 2.850761e-06, 2.17753e-06,
  1.087821e-05, 8.922071e-06, 7.001562e-06, 1.6411e-06, 7.212939e-07, 
    5.097515e-07, 4.171369e-07, 1.525672e-06, 1.761364e-06, 1.292811e-06, 
    2.694502e-06, 4.727234e-06, 6.446136e-06, 5.088122e-06, 2.702967e-06,
  1.382932e-05, 2.62202e-05, 8.028926e-05, 0.0001393281, 0.0001429296, 
    0.0001290288, 0.0001057481, 7.795159e-05, 5.522622e-05, 4.731688e-05, 
    4.716304e-05, 4.923122e-05, 5.002783e-05, 4.408939e-05, 3.861147e-05,
  9.162965e-06, 1.124388e-05, 3.320499e-05, 0.0001045496, 0.0001427837, 
    0.0001336592, 0.0001171391, 8.987501e-05, 6.469672e-05, 5.146631e-05, 
    4.928187e-05, 5.14723e-05, 4.563592e-05, 4.023583e-05, 4.01132e-05,
  6.69046e-06, 4.52662e-06, 7.513324e-06, 2.211895e-05, 5.766088e-05, 
    9.645944e-05, 0.0001038359, 0.0001065164, 9.5966e-05, 7.804141e-05, 
    6.135907e-05, 5.086347e-05, 4.161417e-05, 3.185804e-05, 2.687448e-05,
  2.123619e-05, 1.495856e-05, 1.026701e-05, 4.30716e-06, 1.027787e-05, 
    2.891645e-05, 5.757955e-05, 6.262466e-05, 6.803749e-05, 6.847796e-05, 
    5.319432e-05, 3.927577e-05, 2.853585e-05, 1.957708e-05, 1.097696e-05,
  2.800252e-05, 2.124255e-05, 1.791507e-05, 2.855123e-06, 1.83136e-06, 
    6.509983e-06, 9.803878e-06, 1.843315e-05, 3.432885e-05, 3.256711e-05, 
    2.38208e-05, 1.663034e-05, 9.516535e-06, 4.738639e-06, 2.519299e-06,
  2.598838e-05, 2.255016e-05, 1.320579e-05, 3.813932e-06, 1.681987e-06, 
    2.653044e-06, 3.070676e-06, 4.636831e-06, 6.297482e-06, 5.770738e-06, 
    4.215714e-06, 2.479135e-06, 1.305673e-06, 5.92279e-07, 3.506735e-07,
  1.718816e-05, 9.16703e-06, 3.897636e-06, 1.276852e-08, 3.400267e-09, 
    2.225003e-07, 4.341221e-07, 2.029621e-06, 1.346267e-06, 9.380963e-07, 
    7.134956e-07, 4.75037e-07, 2.782302e-07, 1.407254e-07, 9.236664e-08,
  1.071745e-05, 1.247921e-05, 8.366643e-06, 3.850108e-06, 1.759572e-07, 
    8.101851e-08, 4.000256e-08, 6.097103e-08, 3.486591e-07, 3.660222e-07, 
    1.73065e-07, 2.330981e-07, 4.898197e-07, 9.50513e-07, 2.157175e-06,
  1.153235e-05, 9.988294e-06, 9.647932e-06, 6.287079e-06, 1.955942e-07, 
    6.950057e-08, 2.010743e-07, 4.93089e-07, 4.949882e-07, 5.585829e-07, 
    4.415905e-07, 4.723441e-07, 2.200445e-06, 6.007785e-06, 9.146805e-06,
  2.194183e-05, 1.5827e-05, 1.398104e-05, 3.401965e-06, 4.207266e-07, 
    5.498288e-08, 2.150613e-07, 8.987222e-07, 3.290286e-07, 6.604113e-07, 
    1.217465e-06, 1.942988e-06, 5.841284e-06, 1.151689e-05, 1.581442e-05,
  1.27105e-06, 6.418084e-06, 4.543457e-05, 9.93421e-05, 8.997634e-05, 
    6.460482e-05, 4.522901e-05, 2.847009e-05, 1.961976e-05, 9.082013e-06, 
    3.958487e-06, 4.069648e-06, 2.314717e-06, 5.998032e-06, 5.260761e-06,
  9.539234e-07, 1.528715e-06, 1.621191e-05, 8.46378e-05, 0.0001126973, 
    9.356533e-05, 7.920782e-05, 3.483188e-05, 1.806266e-05, 8.057896e-06, 
    2.619543e-06, 2.585358e-06, 1.202804e-06, 4.911942e-06, 3.23577e-06,
  6.658607e-06, 1.770935e-06, 4.092759e-06, 4.512348e-05, 0.0001046662, 
    0.0001017736, 8.26652e-05, 6.217987e-05, 2.190505e-05, 8.427603e-06, 
    3.487214e-06, 2.424922e-06, 2.326795e-06, 4.104957e-06, 6.88745e-06,
  9.169349e-06, 3.772298e-06, 2.476328e-06, 1.325308e-05, 7.146217e-05, 
    9.567245e-05, 8.426827e-05, 6.622593e-05, 4.025456e-05, 1.88659e-05, 
    1.274446e-05, 9.335682e-06, 1.170693e-05, 1.558151e-05, 1.930249e-05,
  9.803961e-06, 2.456559e-06, 3.738681e-07, 2.951748e-06, 2.647152e-05, 
    9.520617e-05, 8.060009e-05, 5.876657e-05, 7.822653e-05, 4.892761e-05, 
    3.440371e-05, 2.615372e-05, 2.616225e-05, 2.560151e-05, 2.813205e-05,
  3.909835e-06, 8.191795e-07, 2.884808e-09, 4.03501e-07, 4.182345e-06, 
    3.316128e-05, 0.0001071334, 9.217676e-05, 6.053752e-05, 4.83284e-05, 
    3.544313e-05, 2.956725e-05, 2.683557e-05, 2.471603e-05, 2.590719e-05,
  1.741254e-06, 5.193853e-07, 2.222914e-09, 8.366613e-08, 1.020116e-06, 
    3.777513e-06, 2.988616e-05, 7.797305e-05, 6.398784e-05, 3.50898e-05, 
    2.735727e-05, 2.632581e-05, 2.502395e-05, 2.257059e-05, 2.11457e-05,
  1.123855e-06, 1.52073e-06, 6.360384e-07, 5.596669e-07, 8.311298e-07, 
    4.394382e-07, 2.921525e-06, 1.637577e-05, 2.913807e-05, 3.182172e-05, 
    3.230324e-05, 3.074719e-05, 2.816907e-05, 2.726118e-05, 2.581952e-05,
  2.097509e-05, 1.695331e-05, 1.418526e-05, 1.135159e-05, 5.228318e-06, 
    8.849697e-07, 4.091885e-07, 2.094044e-06, 1.147909e-05, 2.019986e-05, 
    2.509717e-05, 2.817512e-05, 3.106585e-05, 3.463577e-05, 3.101984e-05,
  8.424965e-05, 9.195059e-05, 6.750884e-05, 4.836814e-05, 3.534351e-05, 
    1.494673e-05, 1.236816e-06, 1.849693e-07, 1.066521e-06, 5.516538e-06, 
    1.200099e-05, 2.2991e-05, 2.90035e-05, 3.017067e-05, 2.168488e-05,
  3.642578e-08, 5.593555e-09, 2.206906e-08, 2.239176e-06, 1.079628e-05, 
    2.581876e-05, 1.688167e-05, 3.123885e-06, 3.690692e-07, 3.541106e-06, 
    4.448807e-06, 4.836881e-06, 6.018652e-06, 1.021168e-05, 1.214272e-05,
  1.576469e-06, 1.563465e-07, 1.334255e-07, 4.902794e-06, 1.272386e-05, 
    2.229711e-05, 1.765728e-05, 5.156907e-06, 3.945821e-06, 3.615541e-06, 
    2.885761e-06, 3.649986e-06, 8.62764e-06, 1.62642e-05, 1.224378e-05,
  9.672151e-06, 3.191669e-06, 6.009247e-07, 6.632486e-06, 1.923448e-05, 
    2.748349e-05, 2.291134e-05, 1.696496e-05, 1.21012e-05, 6.053163e-06, 
    2.669027e-06, 6.081967e-06, 1.325308e-05, 1.600583e-05, 1.112037e-05,
  2.035674e-05, 1.27442e-05, 6.523913e-06, 5.500369e-06, 2.155213e-05, 
    3.032636e-05, 2.704067e-05, 2.346879e-05, 1.567385e-05, 8.154543e-06, 
    7.233792e-06, 1.321387e-05, 1.719178e-05, 1.267106e-05, 9.842167e-06,
  2.797102e-05, 2.177122e-05, 1.157515e-05, 3.3051e-06, 1.52937e-05, 
    3.54704e-05, 2.169382e-05, 2.738391e-05, 2.603352e-05, 8.507252e-06, 
    1.63359e-05, 2.212358e-05, 1.339393e-05, 7.230904e-06, 6.868157e-06,
  2.487049e-05, 2.374646e-05, 1.141959e-05, 2.822598e-06, 6.237781e-06, 
    2.002859e-05, 3.356009e-05, 9.175748e-06, 4.057615e-06, 7.936133e-06, 
    1.868164e-05, 1.615506e-05, 8.796331e-06, 5.612947e-06, 7.30815e-06,
  2.929017e-05, 2.394767e-05, 1.71588e-05, 4.264676e-06, 2.05871e-06, 
    9.905368e-06, 2.145599e-05, 1.607743e-05, 5.774696e-06, 8.744107e-06, 
    1.688987e-05, 1.141123e-05, 7.750362e-06, 6.710735e-06, 5.619077e-06,
  4.313924e-05, 3.035152e-05, 1.999962e-05, 9.383009e-06, 1.079418e-06, 
    4.647899e-06, 1.336936e-05, 2.046905e-05, 9.417749e-06, 8.883308e-06, 
    1.256715e-05, 1.026764e-05, 7.068888e-06, 6.47792e-06, 6.409043e-06,
  5.26428e-05, 3.810195e-05, 2.585025e-05, 1.443809e-05, 4.000138e-06, 
    2.14208e-06, 7.262773e-06, 1.268062e-05, 1.760943e-05, 1.037576e-05, 
    9.256534e-06, 8.796308e-06, 7.085468e-06, 9.493761e-06, 1.114797e-05,
  2.089038e-05, 2.081962e-05, 3.243902e-05, 2.66497e-05, 1.322971e-05, 
    5.491115e-06, 4.80583e-06, 6.843585e-06, 9.554927e-06, 1.034041e-05, 
    9.256945e-06, 9.017022e-06, 1.012425e-05, 1.659999e-05, 1.7259e-05,
  8.481023e-06, 6.53405e-06, 5.400012e-06, 7.007673e-06, 4.656521e-06, 
    2.01286e-06, 3.636959e-06, 3.722636e-06, 2.864392e-06, 5.077317e-06, 
    3.951695e-06, 3.776035e-06, 4.277756e-06, 4.780653e-06, 7.457878e-06,
  1.013628e-05, 9.264144e-06, 8.082746e-06, 7.761374e-06, 6.675528e-06, 
    3.878734e-06, 3.505148e-06, 3.397304e-06, 3.927722e-06, 1.479694e-06, 
    5.75172e-06, 5.597981e-06, 6.040478e-06, 6.242711e-06, 7.095908e-06,
  1.893335e-05, 1.309389e-05, 1.341858e-05, 1.198077e-05, 9.415575e-06, 
    9.447467e-06, 4.875717e-06, 3.385524e-06, 3.46035e-06, 3.995917e-06, 
    5.951469e-06, 5.195654e-06, 6.15457e-06, 5.419266e-06, 7.476406e-06,
  2.331684e-05, 3.800853e-05, 4.324695e-05, 1.575238e-05, 1.291972e-05, 
    1.368389e-05, 1.172765e-05, 5.943537e-06, 3.459609e-06, 7.962256e-06, 
    4.900692e-06, 6.288496e-06, 7.871667e-06, 6.723245e-06, 6.04847e-06,
  2.967002e-05, 3.017539e-05, 4.040391e-05, 1.511947e-05, 1.113899e-05, 
    1.123224e-05, 1.427566e-05, 1.764728e-05, 6.470272e-06, 3.354538e-06, 
    7.903473e-06, 9.856101e-06, 5.48155e-06, 4.346108e-06, 6.12227e-06,
  3.751572e-05, 3.572556e-05, 3.689205e-05, 1.3198e-05, 6.760674e-06, 
    3.060755e-06, 1.012052e-05, 5.972306e-06, 2.960349e-06, 6.008652e-06, 
    4.430103e-06, 5.27165e-06, 5.905492e-06, 8.341573e-06, 1.829272e-05,
  4.305034e-05, 4.725371e-05, 4.470745e-05, 2.509654e-05, 1.36527e-05, 
    3.307246e-06, 8.20689e-06, 3.146501e-06, 4.916117e-06, 9.283932e-06, 
    4.237649e-06, 5.103183e-06, 8.552883e-06, 1.65871e-05, 2.148382e-05,
  4.983707e-05, 5.708155e-05, 4.891448e-05, 3.134017e-05, 1.989397e-05, 
    4.721412e-06, 6.198904e-06, 6.116865e-06, 7.261492e-06, 1.148576e-05, 
    4.482326e-06, 5.697063e-06, 1.34636e-05, 1.799986e-05, 4.663428e-06,
  4.510094e-05, 4.597657e-05, 2.312474e-05, 2.219962e-05, 1.57358e-05, 
    6.86397e-06, 6.507978e-06, 7.596538e-06, 1.428982e-05, 1.207051e-05, 
    5.400243e-06, 9.764682e-06, 1.498271e-05, 5.202085e-06, 1.255411e-07,
  2.986728e-05, 1.103538e-05, 1.030925e-05, 1.193648e-05, 1.369841e-05, 
    1.085532e-05, 8.580066e-06, 8.937765e-06, 1.64112e-05, 1.041705e-05, 
    8.126878e-06, 1.224948e-05, 6.971083e-06, 6.116763e-07, 8.282745e-09,
  6.607635e-06, 2.125458e-07, 2.785012e-08, 7.492371e-08, 4.398102e-06, 
    2.066878e-05, 1.282213e-05, 5.245375e-06, 7.872985e-06, 7.268103e-06, 
    7.635869e-06, 5.66121e-06, 1.058756e-05, 2.362747e-05, 3.812885e-05,
  1.90378e-06, 3.708344e-07, 1.04083e-07, 3.391265e-07, 1.909752e-06, 
    1.373915e-05, 1.134152e-05, 4.403176e-06, 3.818216e-06, 4.122018e-06, 
    6.108969e-06, 7.867166e-06, 6.391823e-06, 1.126034e-05, 2.330612e-05,
  1.889085e-05, 3.994734e-06, 2.192639e-06, 1.180042e-06, 1.184242e-06, 
    1.557324e-05, 7.648276e-06, 6.401814e-06, 2.028099e-06, 3.113584e-06, 
    8.206164e-06, 1.004037e-05, 8.613671e-06, 9.121035e-06, 1.143439e-05,
  2.434197e-05, 2.999737e-05, 2.294804e-05, 2.148646e-06, 1.60997e-06, 
    7.410611e-06, 1.219802e-05, 5.060331e-06, 2.637071e-06, 6.730004e-06, 
    8.58821e-06, 1.118646e-05, 1.055054e-05, 1.2076e-05, 1.096156e-05,
  2.587703e-05, 3.021942e-05, 3.187018e-05, 2.859549e-06, 1.594139e-06, 
    2.406332e-06, 8.714184e-06, 3.446839e-06, 1.699565e-05, 8.363882e-06, 
    9.987151e-06, 1.383155e-05, 1.084549e-05, 7.119776e-06, 7.983376e-06,
  3.125373e-05, 3.334905e-05, 3.285695e-05, 9.025805e-06, 2.372536e-06, 
    2.422983e-06, 4.973431e-06, 5.214021e-06, 2.976991e-06, 1.179669e-05, 
    8.523619e-06, 1.05623e-05, 1.030235e-05, 4.359851e-06, 3.034301e-06,
  2.725951e-05, 4.327426e-05, 4.492772e-05, 1.350278e-05, 3.154659e-06, 
    2.265656e-06, 2.026268e-06, 2.471129e-06, 2.328946e-06, 4.54286e-06, 
    9.010092e-06, 1.038079e-05, 7.873236e-06, 2.130791e-06, 3.477297e-07,
  1.771883e-05, 2.341048e-05, 2.06271e-05, 1.472146e-05, 5.924024e-06, 
    3.005916e-06, 1.571931e-06, 1.99982e-06, 1.58743e-06, 4.259709e-06, 
    6.42828e-06, 6.715696e-06, 3.376934e-06, 2.406562e-07, 6.35125e-08,
  8.103398e-06, 1.308263e-05, 1.154724e-05, 1.414536e-05, 9.459099e-06, 
    4.535834e-06, 2.292271e-06, 2.808212e-06, 4.400434e-06, 4.75193e-06, 
    4.885818e-06, 3.100638e-06, 3.353226e-07, 1.185335e-07, 1.183013e-07,
  3.864111e-06, 3.660641e-06, 4.450253e-06, 4.324278e-06, 4.596581e-06, 
    5.834619e-06, 4.925723e-06, 3.659024e-06, 4.849994e-06, 4.143268e-06, 
    3.032139e-06, 3.781487e-07, 1.690023e-07, 1.938869e-07, 2.811093e-08,
  2.857191e-06, 5.346594e-07, 1.018487e-06, 3.544548e-06, 3.12978e-06, 
    4.81503e-06, 2.807589e-06, 7.934032e-06, 4.042604e-06, 4.73671e-06, 
    4.413885e-06, 7.094928e-06, 1.284469e-05, 1.618195e-05, 2.085001e-05,
  9.88438e-07, 4.376413e-07, 7.632441e-07, 2.576837e-06, 1.473213e-06, 
    1.277459e-06, 1.165012e-06, 5.494247e-06, 2.31569e-06, 3.299954e-06, 
    3.065879e-06, 7.529067e-06, 1.269657e-05, 1.160607e-05, 1.981632e-05,
  7.517819e-06, 2.262272e-06, 3.633168e-06, 4.092271e-06, 1.360018e-06, 
    4.11438e-06, 7.791501e-07, 6.342854e-06, 5.29449e-06, 3.549571e-06, 
    3.108519e-06, 3.975685e-06, 5.920167e-06, 1.093358e-05, 2.057857e-05,
  6.336073e-06, 1.269551e-05, 1.519842e-05, 6.266868e-06, 3.913744e-06, 
    1.283425e-06, 1.569684e-06, 1.237406e-06, 1.226707e-06, 4.308298e-06, 
    1.580506e-06, 1.403533e-06, 1.284495e-06, 1.874241e-06, 4.085938e-06,
  7.653063e-06, 1.011568e-05, 1.365362e-05, 2.694714e-06, 3.143737e-06, 
    3.32889e-06, 2.485794e-07, 7.563926e-07, 4.831329e-06, 3.421967e-06, 
    1.493111e-06, 6.539587e-07, 2.414693e-07, 2.475111e-07, 4.331943e-07,
  6.284085e-06, 8.299573e-06, 1.107776e-05, 5.578059e-06, 3.240955e-06, 
    2.519808e-06, 3.444077e-06, 2.977996e-06, 2.083112e-06, 2.298547e-06, 
    1.278447e-06, 4.85706e-07, 5.277755e-07, 3.209139e-07, 4.682665e-07,
  5.667449e-06, 9.084449e-06, 1.113338e-05, 1.023215e-05, 4.777486e-06, 
    3.118325e-06, 1.304222e-06, 9.321028e-07, 1.306599e-06, 2.005176e-06, 
    7.785719e-07, 7.175892e-07, 5.512348e-07, 4.537835e-07, 4.422032e-07,
  4.472454e-06, 6.322271e-06, 1.14048e-05, 1.159712e-05, 1.071348e-05, 
    7.451675e-06, 3.450014e-06, 1.143211e-06, 6.235186e-07, 4.78601e-07, 
    5.927112e-07, 5.075577e-07, 4.805089e-07, 4.390865e-07, 4.3637e-07,
  1.630206e-06, 3.181437e-06, 6.266865e-06, 1.486956e-05, 1.863558e-05, 
    1.418427e-05, 1.010827e-05, 4.587484e-06, 9.418278e-07, 2.991382e-07, 
    2.34524e-07, 3.202003e-07, 3.589327e-07, 3.916416e-07, 5.183081e-07,
  6.41131e-07, 1.683331e-06, 6.492434e-06, 2.12884e-05, 3.302706e-05, 
    2.687819e-05, 1.629229e-05, 1.139107e-05, 4.484291e-06, 9.588658e-07, 
    3.746926e-07, 3.49707e-07, 3.265016e-07, 1.595646e-07, 5.14249e-07,
  1.47573e-06, 4.681267e-06, 1.096231e-05, 1.867182e-05, 2.005293e-05, 
    2.12676e-05, 2.307491e-05, 1.911818e-05, 1.607486e-05, 1.444973e-05, 
    8.315509e-06, 6.12312e-06, 6.3127e-06, 7.124946e-06, 1.162888e-05,
  2.324768e-06, 5.893228e-06, 9.977083e-06, 1.795271e-05, 1.989312e-05, 
    1.618533e-05, 1.820699e-05, 2.225043e-05, 1.833913e-05, 1.678139e-05, 
    1.318427e-05, 6.906214e-06, 3.855583e-06, 5.020598e-06, 5.64721e-06,
  2.961664e-06, 4.809544e-06, 8.928617e-06, 1.824091e-05, 2.773656e-05, 
    2.330862e-05, 9.512338e-06, 1.372136e-05, 2.082867e-05, 2.164031e-05, 
    1.712713e-05, 1.144661e-05, 4.140995e-06, 7.719232e-07, 1.304104e-06,
  4.829899e-06, 6.863836e-06, 1.299045e-05, 2.016821e-05, 3.093778e-05, 
    3.403832e-05, 2.499657e-05, 9.493758e-06, 1.23764e-05, 1.914739e-05, 
    2.207797e-05, 1.517006e-05, 7.069396e-06, 1.623893e-06, 1.405448e-07,
  4.950021e-06, 8.538244e-06, 1.319024e-05, 2.05941e-05, 3.252845e-05, 
    3.424469e-05, 3.582356e-05, 2.98941e-05, 1.405257e-05, 1.020829e-05, 
    2.216998e-05, 1.734244e-05, 9.578234e-06, 1.949431e-06, 4.327527e-07,
  1.036081e-05, 9.171087e-06, 1.179108e-05, 1.898813e-05, 3.115443e-05, 
    3.548579e-05, 4.542008e-05, 4.144385e-05, 2.589331e-05, 2.081293e-05, 
    1.893556e-05, 1.516937e-05, 1.15919e-05, 3.001192e-06, 1.034431e-06,
  1.029333e-05, 1.029146e-05, 1.026155e-05, 1.598244e-05, 3.049712e-05, 
    3.306435e-05, 4.00658e-05, 4.503851e-05, 3.962109e-05, 2.78166e-05, 
    1.909394e-05, 1.582813e-05, 1.293234e-05, 3.302793e-06, 1.595655e-06,
  1.086769e-05, 7.851952e-06, 7.468249e-06, 1.392239e-05, 3.282418e-05, 
    3.330136e-05, 3.895648e-05, 4.494853e-05, 3.96005e-05, 3.265101e-05, 
    2.580519e-05, 1.954489e-05, 1.265498e-05, 2.905529e-06, 1.296804e-06,
  7.232183e-06, 4.765081e-06, 5.13095e-06, 1.060454e-05, 2.717554e-05, 
    2.785868e-05, 3.011778e-05, 3.958883e-05, 4.081932e-05, 3.512866e-05, 
    2.844026e-05, 2.151632e-05, 1.057615e-05, 2.788373e-06, 1.391776e-06,
  4.65598e-06, 2.958412e-06, 1.869267e-06, 3.818021e-06, 8.458086e-06, 
    1.030271e-05, 1.555328e-05, 2.550311e-05, 3.388518e-05, 3.088626e-05, 
    2.844049e-05, 2.07881e-05, 9.294458e-06, 3.4123e-06, 1.841372e-06,
  9.733226e-06, 1.875568e-05, 2.651564e-05, 2.304172e-05, 1.272898e-05, 
    9.729786e-06, 9.520051e-06, 7.494637e-06, 7.103237e-06, 1.037166e-05, 
    1.898014e-05, 2.832575e-05, 3.325667e-05, 3.550378e-05, 3.058705e-05,
  7.763367e-06, 1.213667e-05, 1.662779e-05, 1.153484e-05, 5.994943e-06, 
    3.006253e-06, 4.228052e-06, 6.557891e-06, 3.647682e-06, 4.179559e-06, 
    8.185476e-06, 2.009327e-05, 3.054514e-05, 2.855056e-05, 2.503689e-05,
  7.515002e-06, 1.28927e-05, 1.14329e-05, 7.15745e-06, 3.609601e-06, 
    6.09406e-06, 1.681594e-06, 4.555905e-06, 5.776456e-06, 3.290057e-06, 
    4.625274e-06, 1.239697e-05, 2.416136e-05, 2.497244e-05, 2.340945e-05,
  7.804935e-06, 1.288256e-05, 1.581812e-05, 8.004167e-06, 3.433952e-06, 
    5.514425e-06, 8.027847e-06, 2.483973e-06, 2.76999e-06, 3.255914e-06, 
    3.303554e-06, 8.285539e-06, 1.769989e-05, 2.529624e-05, 2.410843e-05,
  6.310185e-06, 9.406443e-06, 9.276744e-06, 3.511243e-06, 3.896857e-06, 
    6.158067e-06, 8.561957e-06, 1.516191e-05, 2.861026e-05, 8.464671e-06, 
    4.195615e-06, 6.184771e-06, 1.717815e-05, 2.349467e-05, 1.832574e-05,
  4.235699e-06, 5.524889e-06, 6.871463e-06, 4.358541e-06, 7.908058e-06, 
    1.264859e-05, 9.754162e-06, 1.193614e-05, 1.890591e-05, 1.093329e-05, 
    7.395244e-06, 5.494631e-06, 1.724666e-05, 1.391357e-05, 6.551376e-06,
  5.68476e-06, 3.668855e-06, 6.026113e-06, 9.007333e-06, 9.011469e-06, 
    7.040855e-06, 9.246983e-06, 9.58131e-06, 8.591444e-06, 6.703292e-06, 
    4.7662e-06, 4.726931e-06, 9.971376e-06, 6.376828e-06, 1.776155e-06,
  3.432311e-06, 2.191285e-06, 7.256084e-06, 7.374222e-06, 8.216655e-06, 
    4.075862e-06, 3.641343e-06, 5.203771e-06, 6.831413e-06, 7.614181e-06, 
    1.262799e-06, 4.38916e-06, 4.447214e-06, 2.453785e-06, 1.305363e-06,
  2.62367e-06, 2.521291e-06, 3.868792e-06, 4.745079e-06, 7.172675e-06, 
    3.788321e-06, 2.045917e-06, 1.754687e-06, 4.381861e-06, 4.971848e-06, 
    4.031809e-06, 3.25722e-06, 2.191298e-06, 1.574767e-06, 5.740289e-07,
  3.140642e-06, 2.410171e-06, 2.835434e-06, 4.17163e-06, 5.493984e-06, 
    6.114498e-06, 3.638081e-06, 2.885893e-06, 3.424661e-06, 3.027928e-06, 
    3.590222e-06, 2.712324e-06, 1.343521e-06, 1.057863e-06, 7.29107e-07,
  6.031657e-07, 1.94382e-06, 3.410537e-06, 4.938014e-06, 5.027573e-06, 
    5.831987e-06, 4.758986e-06, 2.792258e-06, 4.627833e-06, 5.826408e-06, 
    3.46825e-06, 4.841118e-06, 3.235692e-06, 5.692445e-07, 3.738388e-06,
  5.795418e-07, 1.629186e-06, 3.52746e-06, 5.99646e-06, 9.114502e-06, 
    9.48582e-06, 9.81892e-06, 7.166051e-06, 7.011585e-06, 4.677683e-06, 
    1.511134e-06, 3.331346e-06, 1.243811e-06, 2.872758e-06, 3.267209e-07,
  9.452701e-07, 2.546745e-06, 4.160592e-06, 6.845165e-06, 1.462973e-05, 
    2.779147e-05, 9.089025e-06, 1.166943e-05, 1.222739e-05, 7.492119e-06, 
    3.872279e-06, 2.206101e-06, 2.138923e-06, 5.066991e-06, 1.570892e-06,
  2.129821e-06, 5.353869e-06, 6.735141e-06, 9.347216e-06, 1.728749e-05, 
    2.363886e-05, 2.898831e-05, 1.047337e-05, 1.259775e-05, 1.164794e-05, 
    8.356772e-06, 3.753139e-06, 4.394614e-06, 3.573502e-06, 4.118218e-06,
  3.623582e-06, 5.799456e-06, 8.645906e-06, 1.21087e-05, 1.838479e-05, 
    2.239284e-05, 2.676448e-05, 3.112967e-05, 1.996907e-05, 1.212694e-05, 
    1.40082e-05, 6.826506e-06, 4.064396e-06, 2.444458e-06, 5.434849e-06,
  6.456984e-06, 9.351489e-06, 1.261726e-05, 1.383309e-05, 1.789056e-05, 
    2.250986e-05, 3.320343e-05, 2.49549e-05, 2.007926e-05, 2.543923e-05, 
    2.014254e-05, 1.082849e-05, 5.305354e-06, 2.66434e-06, 2.830016e-06,
  7.804975e-06, 8.765212e-06, 1.31097e-05, 1.553636e-05, 2.051566e-05, 
    2.574728e-05, 3.293706e-05, 3.804691e-05, 3.631381e-05, 3.400521e-05, 
    3.049661e-05, 1.93004e-05, 8.791612e-06, 3.469265e-06, 1.369635e-06,
  7.71608e-06, 7.050313e-06, 1.086156e-05, 1.428533e-05, 1.800622e-05, 
    2.426667e-05, 3.35074e-05, 3.668338e-05, 3.93657e-05, 4.757883e-05, 
    4.763911e-05, 2.974239e-05, 1.325197e-05, 4.295082e-06, 1.245787e-06,
  9.319819e-06, 1.00787e-05, 1.29644e-05, 1.550233e-05, 1.671849e-05, 
    2.183804e-05, 3.235508e-05, 4.351713e-05, 5.341333e-05, 5.798023e-05, 
    5.21623e-05, 3.524373e-05, 1.556818e-05, 4.215314e-06, 1.078931e-06,
  1.008973e-05, 1.493605e-05, 1.685692e-05, 1.725286e-05, 1.690627e-05, 
    1.81432e-05, 2.709248e-05, 4.661396e-05, 6.857825e-05, 7.167758e-05, 
    5.696597e-05, 3.455849e-05, 1.19796e-05, 2.402789e-06, 1.132654e-06,
  6.638101e-06, 1.301942e-05, 1.782543e-05, 2.534626e-05, 2.907985e-05, 
    3.178216e-05, 3.381485e-05, 3.40043e-05, 3.841773e-05, 3.806161e-05, 
    2.752172e-05, 2.280989e-05, 1.840255e-05, 7.980732e-06, 2.107726e-06,
  6.158331e-06, 9.597584e-06, 1.545364e-05, 2.167601e-05, 2.038195e-05, 
    1.895581e-05, 2.530723e-05, 2.447783e-05, 2.11715e-05, 2.53448e-05, 
    3.069444e-05, 3.189598e-05, 2.547427e-05, 1.704046e-05, 9.442443e-06,
  5.017254e-06, 8.856165e-06, 1.329597e-05, 1.968556e-05, 2.390478e-05, 
    3.343881e-05, 1.409842e-05, 2.202973e-05, 2.487752e-05, 2.165356e-05, 
    2.435174e-05, 2.882192e-05, 3.017202e-05, 2.44482e-05, 2.298088e-05,
  5.98784e-06, 9.637763e-06, 1.741905e-05, 1.720458e-05, 2.334792e-05, 
    2.606469e-05, 3.442667e-05, 9.60217e-06, 1.584214e-05, 2.589181e-05, 
    2.743678e-05, 2.668694e-05, 3.397054e-05, 3.953476e-05, 3.369067e-05,
  5.072397e-06, 5.444701e-06, 1.310047e-05, 1.128843e-05, 1.354665e-05, 
    1.884197e-05, 2.447491e-05, 4.525565e-05, 3.229326e-05, 1.54449e-05, 
    2.218269e-05, 2.665855e-05, 3.638975e-05, 4.991259e-05, 4.753424e-05,
  5.772853e-06, 5.985385e-06, 1.033504e-05, 8.9901e-06, 8.447533e-06, 
    1.106621e-05, 1.649515e-05, 2.615687e-05, 2.328879e-05, 2.098322e-05, 
    2.40832e-05, 3.449217e-05, 5.279537e-05, 6.314324e-05, 5.560234e-05,
  7.536327e-06, 9.849145e-06, 7.960937e-06, 8.109299e-06, 6.285924e-06, 
    5.2246e-06, 6.717226e-06, 1.129161e-05, 1.338691e-05, 1.873858e-05, 
    2.850707e-05, 4.820794e-05, 6.713028e-05, 7.130772e-05, 4.782142e-05,
  1.143997e-05, 1.257395e-05, 9.801111e-06, 8.646679e-06, 6.033489e-06, 
    7.181767e-06, 4.738357e-06, 5.243964e-06, 6.67086e-06, 1.598077e-05, 
    3.030236e-05, 5.653385e-05, 8.246356e-05, 6.431402e-05, 2.46858e-05,
  1.568762e-05, 2.093203e-05, 1.19412e-05, 6.450409e-06, 4.943589e-06, 
    3.751538e-06, 3.309372e-06, 2.665819e-06, 5.97453e-06, 1.256368e-05, 
    2.302296e-05, 5.474315e-05, 5.482605e-05, 2.258072e-05, 3.99523e-06,
  1.615375e-05, 2.131334e-05, 1.489193e-05, 6.682694e-06, 4.159382e-06, 
    3.944489e-06, 3.437529e-06, 2.347167e-06, 4.853558e-06, 1.155209e-05, 
    1.946909e-05, 2.767286e-05, 1.818673e-05, 2.763691e-06, 4.463305e-07,
  4.101512e-05, 3.133074e-05, 2.57897e-05, 1.857648e-05, 9.792497e-06, 
    4.089478e-06, 3.961394e-06, 1.963772e-06, 6.483915e-06, 1.018852e-05, 
    1.775774e-05, 3.282847e-05, 3.984452e-05, 2.646388e-05, 1.063493e-05,
  4.14328e-05, 2.873408e-05, 2.162288e-05, 1.692032e-05, 1.024103e-05, 
    3.806688e-06, 2.175893e-06, 9.934391e-07, 1.750088e-06, 3.924121e-06, 
    9.03964e-06, 2.035352e-05, 2.824403e-05, 2.290268e-05, 2.156869e-05,
  3.803498e-05, 3.216425e-05, 2.395353e-05, 1.707575e-05, 1.112399e-05, 
    7.389408e-06, 1.732106e-06, 1.260554e-06, 3.015616e-06, 5.387753e-06, 
    7.448266e-06, 1.120346e-05, 1.593324e-05, 2.278015e-05, 3.73276e-05,
  3.938888e-05, 3.486237e-05, 2.75401e-05, 2.239769e-05, 1.197531e-05, 
    4.690702e-06, 3.687309e-06, 4.944704e-07, 5.355678e-07, 2.80055e-06, 
    4.339315e-06, 5.797706e-06, 1.162503e-05, 1.856421e-05, 3.396555e-05,
  4.30659e-05, 3.924857e-05, 3.195913e-05, 2.603415e-05, 1.750872e-05, 
    6.323052e-06, 3.976286e-06, 3.716373e-06, 6.83831e-06, 2.884454e-06, 
    5.072425e-06, 6.368673e-06, 6.990531e-06, 1.10531e-05, 3.025123e-05,
  4.477098e-05, 4.128373e-05, 3.466855e-05, 3.092836e-05, 2.254233e-05, 
    9.554949e-06, 9.21378e-06, 3.886159e-06, 3.719564e-06, 3.547747e-06, 
    3.352349e-06, 5.740018e-06, 7.484824e-06, 1.35696e-05, 3.697495e-05,
  3.856458e-05, 4.085762e-05, 3.604017e-05, 3.031586e-05, 2.750986e-05, 
    1.406261e-05, 8.285342e-06, 5.242468e-06, 1.917005e-06, 9.820038e-07, 
    3.329853e-06, 5.168516e-06, 1.064854e-05, 2.363082e-05, 3.947963e-05,
  3.346894e-05, 4.297211e-05, 3.737487e-05, 2.776522e-05, 2.617969e-05, 
    1.721402e-05, 8.585906e-06, 5.213619e-06, 2.027785e-06, 1.252404e-06, 
    2.887381e-06, 1.354412e-06, 3.892639e-06, 9.236095e-06, 1.191479e-05,
  2.917784e-05, 3.858234e-05, 3.012253e-05, 2.325791e-05, 2.1916e-05, 
    1.889723e-05, 1.216116e-05, 6.770893e-06, 4.00053e-06, 2.555603e-06, 
    1.662173e-06, 1.523119e-06, 1.367869e-06, 1.157944e-06, 1.861623e-06,
  2.025328e-05, 2.366154e-05, 2.109369e-05, 2.015796e-05, 1.74276e-05, 
    1.704446e-05, 1.408262e-05, 9.34011e-06, 8.745174e-06, 1.104247e-05, 
    8.11157e-06, 3.61347e-06, 1.644223e-06, 1.041105e-06, 6.044559e-07,
  3.889613e-05, 4.117163e-05, 4.374503e-05, 3.295602e-05, 1.796316e-05, 
    8.894998e-06, 4.047855e-06, 4.508968e-06, 2.520714e-06, 3.133598e-06, 
    5.248157e-06, 4.943696e-06, 3.532622e-06, 6.722124e-06, 1.425048e-05,
  3.598855e-05, 3.733556e-05, 4.268298e-05, 3.206674e-05, 1.660696e-05, 
    5.61484e-06, 4.23752e-06, 3.602456e-06, 1.177572e-06, 3.418594e-07, 
    1.108947e-06, 3.577455e-06, 5.80003e-06, 6.092935e-06, 7.500123e-06,
  2.591107e-05, 3.39742e-05, 3.995591e-05, 3.338035e-05, 2.344384e-05, 
    1.678593e-05, 3.896346e-06, 5.369693e-06, 2.418677e-06, 7.122343e-07, 
    1.172658e-06, 2.306061e-06, 3.439695e-06, 3.581982e-06, 3.295255e-06,
  2.303939e-05, 2.741561e-05, 3.64737e-05, 3.621188e-05, 2.147714e-05, 
    1.876957e-05, 2.200099e-05, 3.607297e-06, 3.594878e-06, 1.795983e-06, 
    1.472443e-06, 1.384547e-06, 2.727595e-06, 3.715613e-06, 3.154121e-06,
  1.460509e-05, 2.108531e-05, 3.129655e-05, 3.04531e-05, 1.947203e-05, 
    1.428495e-05, 2.022769e-05, 2.776962e-05, 7.999642e-06, 1.798253e-06, 
    2.061307e-06, 1.857879e-06, 3.446252e-06, 5.965988e-06, 6.494792e-06,
  1.006728e-05, 1.258265e-05, 2.490653e-05, 2.407088e-05, 1.525813e-05, 
    1.068547e-05, 1.273063e-05, 1.194606e-05, 6.227807e-06, 6.395406e-06, 
    5.623945e-06, 4.213111e-06, 4.251625e-06, 4.853247e-06, 5.560096e-06,
  7.860331e-06, 1.352633e-05, 2.021242e-05, 1.922524e-05, 1.450123e-05, 
    9.149779e-06, 7.660852e-06, 9.469903e-06, 8.367711e-06, 5.869184e-06, 
    7.839971e-06, 9.727079e-06, 7.599115e-06, 7.589967e-06, 3.810824e-06,
  1.200404e-05, 1.341312e-05, 1.631941e-05, 1.468135e-05, 1.159511e-05, 
    8.448323e-06, 8.014434e-06, 7.353605e-06, 7.203326e-06, 9.405928e-06, 
    1.287964e-05, 1.288467e-05, 1.227618e-05, 1.078916e-05, 8.249416e-06,
  1.055901e-05, 1.295019e-05, 1.46495e-05, 8.415638e-06, 6.028593e-06, 
    6.719053e-06, 8.023253e-06, 7.712202e-06, 5.832712e-06, 9.469477e-06, 
    1.601327e-05, 1.90663e-05, 1.684608e-05, 1.286778e-05, 1.007646e-05,
  3.715172e-06, 9.530222e-06, 1.100721e-05, 6.094502e-06, 4.448116e-06, 
    5.125815e-06, 4.408828e-06, 5.145233e-06, 4.792059e-06, 7.750371e-06, 
    1.920909e-05, 2.666587e-05, 2.475762e-05, 1.927682e-05, 1.416791e-05,
  1.439743e-05, 1.192392e-05, 1.245272e-05, 9.383219e-06, 3.219293e-06, 
    4.963544e-06, 6.567281e-06, 6.815436e-06, 1.556924e-05, 1.71741e-05, 
    8.469676e-06, 3.56599e-06, 5.689407e-06, 4.914103e-06, 5.438765e-06,
  1.019714e-05, 1.05648e-05, 1.179964e-05, 7.093552e-06, 1.537817e-06, 
    2.009106e-06, 6.853895e-06, 7.140505e-06, 1.135985e-05, 1.909482e-05, 
    2.007678e-05, 1.17695e-05, 5.602792e-06, 6.108985e-06, 4.572797e-06,
  9.197968e-06, 1.050248e-05, 1.017436e-05, 5.201524e-06, 2.462209e-06, 
    8.972913e-06, 3.371903e-06, 1.009156e-05, 1.45952e-05, 2.250028e-05, 
    2.582111e-05, 2.325742e-05, 1.432057e-05, 6.51588e-06, 4.255116e-06,
  1.102068e-05, 1.261986e-05, 1.40299e-05, 7.50139e-06, 3.516194e-06, 
    7.932478e-06, 8.234923e-06, 3.980907e-06, 7.364662e-06, 1.412486e-05, 
    1.918843e-05, 2.466567e-05, 2.628754e-05, 1.815756e-05, 9.966549e-06,
  1.183686e-05, 1.099616e-05, 1.211055e-05, 7.232907e-06, 4.052902e-06, 
    4.564081e-06, 5.427207e-06, 9.233634e-06, 1.271872e-05, 9.297801e-06, 
    1.403614e-05, 1.957972e-05, 2.795052e-05, 2.849449e-05, 2.24433e-05,
  1.161815e-05, 1.016236e-05, 1.052998e-05, 8.818809e-06, 6.866701e-06, 
    3.930336e-06, 4.154159e-06, 9.433869e-06, 1.220731e-05, 9.187334e-06, 
    8.967043e-06, 1.198132e-05, 1.713449e-05, 2.53968e-05, 2.971306e-05,
  1.64255e-05, 1.471155e-05, 9.100119e-06, 8.152577e-06, 6.290172e-06, 
    4.756052e-06, 4.342132e-06, 2.696957e-06, 3.256094e-06, 3.327058e-06, 
    4.064829e-06, 5.303519e-06, 8.289448e-06, 1.503204e-05, 2.376429e-05,
  1.847534e-05, 1.780826e-05, 1.051144e-05, 6.323956e-06, 3.919811e-06, 
    3.470754e-06, 2.769641e-06, 3.105492e-06, 3.135676e-06, 2.599355e-06, 
    2.823292e-06, 3.322484e-06, 4.056401e-06, 6.919201e-06, 1.488002e-05,
  2.089241e-05, 1.916016e-05, 7.797305e-06, 3.713711e-06, 1.398799e-06, 
    3.352866e-06, 2.999853e-06, 1.828931e-06, 1.780411e-06, 2.347998e-06, 
    3.041642e-06, 2.834437e-06, 3.425802e-06, 5.319316e-06, 1.049865e-05,
  1.96816e-05, 1.166406e-05, 4.822872e-06, 2.600563e-06, 2.331818e-06, 
    2.684914e-06, 1.80937e-06, 4.229384e-06, 3.939029e-06, 1.533045e-06, 
    1.775857e-06, 1.92466e-06, 2.155235e-06, 3.326262e-06, 8.052419e-06,
  3.823036e-06, 1.722837e-06, 2.204176e-06, 2.273771e-06, 1.405613e-06, 
    2.315569e-06, 2.078667e-06, 2.647844e-06, 3.857057e-06, 1.059463e-05, 
    2.449346e-05, 3.355649e-05, 3.444398e-05, 1.858728e-05, 1.108764e-05,
  5.232086e-06, 2.482222e-06, 2.120563e-06, 9.907995e-07, 4.684273e-07, 
    2.670209e-07, 9.218193e-07, 1.665502e-06, 2.605895e-06, 4.361797e-06, 
    1.326324e-05, 2.732466e-05, 3.239726e-05, 2.653765e-05, 1.551077e-05,
  1.469253e-05, 1.40163e-05, 9.697645e-06, 2.069293e-06, 7.75413e-07, 
    2.253259e-06, 5.82697e-08, 2.958585e-07, 7.874264e-07, 1.629659e-06, 
    2.906928e-06, 1.164672e-05, 2.451922e-05, 3.267221e-05, 2.197865e-05,
  1.727625e-05, 1.787983e-05, 1.610623e-05, 2.155446e-06, 1.018584e-06, 
    1.060212e-06, 1.487366e-06, 8.257927e-08, 8.39409e-08, 1.500305e-06, 
    1.614224e-06, 3.215107e-06, 1.070458e-05, 2.531942e-05, 2.790932e-05,
  2.503722e-05, 1.91714e-05, 2.041499e-05, 2.967036e-06, 2.198851e-06, 
    1.826794e-06, 2.044904e-06, 2.151331e-06, 3.415986e-06, 2.049169e-06, 
    2.687041e-06, 1.864304e-06, 2.848835e-06, 1.544285e-05, 2.835187e-05,
  3.044366e-05, 2.771818e-05, 2.079203e-05, 6.830613e-06, 9.339456e-06, 
    1.881258e-06, 2.889221e-06, 3.549088e-06, 2.335091e-06, 1.35121e-06, 
    1.074721e-06, 1.068414e-06, 1.184083e-06, 4.810095e-06, 2.195123e-05,
  3.564577e-05, 3.625392e-05, 2.317411e-05, 1.352968e-05, 9.56525e-06, 
    2.860366e-06, 2.665161e-06, 3.26491e-06, 2.920588e-06, 1.656448e-06, 
    1.049178e-06, 1.191714e-06, 1.072693e-06, 1.542606e-06, 8.505226e-06,
  3.979902e-05, 4.084666e-05, 3.001386e-05, 9.130778e-06, 8.880575e-06, 
    4.07709e-06, 3.380457e-06, 3.002475e-06, 2.808185e-06, 1.848268e-06, 
    1.405174e-06, 1.070136e-06, 1.221202e-06, 8.560918e-07, 4.147924e-06,
  4.423504e-05, 4.132604e-05, 2.842616e-05, 2.443813e-06, 3.22052e-06, 
    6.298375e-06, 4.001747e-06, 4.490335e-06, 4.33632e-06, 3.725397e-06, 
    1.550007e-06, 1.142719e-06, 9.107201e-07, 9.147846e-07, 3.854056e-06,
  3.296093e-05, 2.239185e-05, 1.072381e-05, 8.602588e-07, 1.359883e-06, 
    4.440075e-06, 5.437851e-06, 9.599296e-06, 8.575014e-06, 3.751373e-06, 
    1.571621e-06, 7.843593e-07, 5.573798e-07, 8.179219e-07, 2.622607e-06,
  1.036346e-05, 1.360376e-05, 2.481936e-05, 1.585209e-05, 1.685585e-05, 
    1.81655e-05, 8.874928e-06, 1.084374e-06, 4.586457e-07, 7.286239e-07, 
    4.338559e-07, 3.284416e-07, 6.252796e-06, 1.510548e-05, 1.615662e-05,
  1.119172e-05, 9.357195e-06, 1.37781e-05, 1.758245e-05, 1.509957e-05, 
    2.341924e-05, 8.253883e-06, 3.759668e-07, 3.184863e-07, 5.120792e-07, 
    4.087873e-07, 3.89433e-07, 4.326457e-07, 3.312893e-06, 9.599643e-06,
  2.73434e-05, 2.76329e-05, 2.314893e-05, 1.005164e-05, 1.553409e-05, 
    2.752692e-05, 1.889557e-05, 1.38869e-06, 1.049718e-06, 4.142709e-07, 
    5.936309e-07, 5.095709e-07, 3.250611e-07, 8.352626e-07, 7.032056e-06,
  4.083438e-05, 4.346398e-05, 3.969638e-05, 1.491101e-05, 1.549417e-05, 
    2.102976e-05, 2.26428e-05, 5.385126e-06, 2.836296e-06, 1.285035e-06, 
    1.507062e-06, 6.126218e-07, 6.446154e-07, 5.317975e-07, 5.187976e-06,
  4.286005e-05, 3.804749e-05, 3.836197e-05, 4.25552e-06, 1.182079e-05, 
    2.357537e-05, 1.580712e-05, 8.805299e-06, 5.517543e-06, 5.925048e-07, 
    2.183015e-06, 6.358276e-07, 3.411167e-07, 3.716581e-07, 5.011133e-06,
  4.719413e-05, 3.620649e-05, 3.188103e-05, 1.500135e-05, 1.513138e-05, 
    1.395509e-05, 2.14386e-05, 8.585695e-06, 8.529556e-07, 2.062883e-07, 
    5.028103e-07, 5.299337e-07, 3.795314e-07, 2.961817e-07, 1.864357e-06,
  4.610274e-05, 4.705646e-05, 3.886412e-05, 2.32709e-05, 1.45475e-05, 
    5.466135e-06, 1.093817e-05, 1.077893e-05, 3.9524e-06, 1.245871e-06, 
    1.098131e-06, 1.041297e-06, 7.719915e-07, 2.390306e-07, 4.621059e-07,
  5.787944e-05, 5.332554e-05, 4.313867e-05, 2.293134e-05, 1.379623e-05, 
    6.400764e-06, 5.807088e-06, 4.203606e-06, 2.729658e-06, 2.172636e-06, 
    1.320552e-06, 1.497271e-06, 7.790243e-07, 2.273655e-07, 4.042923e-07,
  5.795346e-05, 5.514608e-05, 3.714349e-05, 1.305042e-05, 7.986494e-06, 
    5.546428e-06, 6.445732e-06, 6.040099e-06, 4.095583e-06, 2.31147e-06, 
    1.050234e-06, 1.416139e-06, 4.471771e-07, 2.420637e-07, 5.058898e-07,
  3.879571e-05, 2.271585e-05, 2.327551e-05, 1.447414e-05, 6.821438e-06, 
    6.990836e-06, 6.644602e-06, 6.919451e-06, 5.254493e-06, 2.16782e-06, 
    7.922299e-07, 1.209045e-06, 4.952789e-07, 2.184421e-07, 4.751644e-07,
  7.528243e-06, 1.446315e-06, 2.434826e-06, 2.262369e-06, 2.14769e-06, 
    3.616951e-06, 1.114268e-05, 1.523413e-05, 1.13557e-05, 5.034968e-06, 
    2.546715e-06, 1.195922e-06, 4.745231e-06, 1.49068e-05, 7.316783e-06,
  1.612865e-05, 5.285975e-06, 1.544466e-06, 4.129111e-06, 6.624329e-06, 
    1.567154e-05, 2.456007e-05, 1.935913e-05, 1.404894e-05, 6.90858e-06, 
    2.06976e-06, 4.734865e-07, 5.382559e-06, 1.561649e-05, 1.027983e-05,
  3.255886e-05, 3.482883e-05, 2.705075e-05, 8.844693e-06, 2.117623e-05, 
    2.549434e-05, 3.965773e-05, 3.366292e-05, 1.71038e-05, 4.894079e-06, 
    9.385685e-07, 6.146185e-07, 5.733202e-06, 1.871468e-05, 9.504618e-06,
  4.249178e-05, 4.442212e-05, 4.354524e-05, 1.545418e-05, 1.371496e-05, 
    1.383258e-05, 2.945132e-05, 3.001557e-05, 7.30953e-06, 2.535631e-06, 
    1.187597e-06, 7.591621e-07, 6.387875e-06, 1.52229e-05, 6.707423e-06,
  5.130782e-05, 4.902794e-05, 4.162485e-05, 7.452168e-06, 1.577248e-06, 
    7.344394e-06, 1.735911e-05, 1.096811e-05, 2.531563e-06, 1.161019e-06, 
    1.361019e-06, 9.949189e-07, 7.918285e-06, 1.171788e-05, 5.437718e-06,
  5.455736e-05, 5.70782e-05, 4.628299e-05, 1.621962e-05, 5.839102e-06, 
    2.34199e-06, 1.892278e-05, 9.405491e-06, 6.244283e-07, 8.754186e-07, 
    9.740389e-07, 1.506899e-06, 5.372193e-06, 6.859064e-06, 5.384763e-06,
  5.459883e-05, 6.420424e-05, 6.116135e-05, 3.364755e-05, 1.261837e-05, 
    2.751327e-06, 1.202968e-05, 1.459076e-05, 1.72946e-06, 1.265919e-06, 
    1.814428e-06, 2.113854e-06, 3.503101e-06, 5.650661e-06, 6.927757e-06,
  5.457462e-05, 6.151434e-05, 5.422429e-05, 3.39173e-05, 1.866792e-05, 
    1.137819e-05, 1.029524e-05, 5.164635e-06, 6.677683e-07, 2.411643e-06, 
    2.451962e-06, 3.694953e-06, 5.828005e-06, 7.242197e-06, 7.300567e-06,
  3.81868e-05, 4.593965e-05, 3.345068e-05, 1.938471e-05, 1.32838e-05, 
    1.129551e-05, 7.065895e-06, 1.463857e-06, 3.223007e-07, 1.818908e-06, 
    2.232792e-06, 4.461019e-06, 6.912608e-06, 6.498795e-06, 3.839779e-06,
  1.557918e-05, 1.257006e-05, 1.240801e-05, 1.092262e-05, 5.17454e-06, 
    2.648219e-06, 2.15417e-06, 2.020126e-06, 1.057492e-06, 1.542339e-06, 
    2.248254e-06, 3.781749e-06, 5.182141e-06, 4.588097e-06, 3.386362e-06,
  3.292527e-06, 5.734955e-08, 1.295232e-07, 4.857708e-08, 4.048519e-06, 
    9.66181e-06, 4.655707e-06, 6.025221e-07, 1.055885e-05, 5.452209e-05, 
    3.57853e-05, 1.541386e-05, 1.061291e-05, 5.460783e-06, 1.19437e-06,
  1.398212e-05, 1.995626e-06, 3.662454e-07, 8.472109e-07, 7.871649e-06, 
    1.457547e-05, 9.66577e-06, 4.810332e-06, 2.114518e-05, 3.879038e-05, 
    1.999221e-05, 9.277997e-06, 4.778016e-06, 1.723537e-06, 1.136958e-06,
  2.905924e-05, 2.161065e-05, 1.277884e-05, 2.657395e-06, 6.045068e-06, 
    1.604977e-05, 1.615227e-05, 1.762682e-05, 2.464797e-05, 2.484825e-05, 
    6.413655e-06, 3.556189e-06, 1.963622e-06, 4.906129e-07, 4.249999e-07,
  3.069475e-05, 2.692691e-05, 1.578927e-05, 4.813944e-06, 4.433013e-06, 
    1.151461e-05, 2.308534e-05, 2.71505e-05, 3.037892e-05, 2.154262e-05, 
    2.589233e-06, 7.534198e-07, 1.24184e-06, 7.932331e-07, 1.417205e-06,
  3.36261e-05, 2.104814e-05, 1.324541e-05, 2.321099e-06, 2.316746e-06, 
    9.134583e-06, 1.233277e-05, 4.76415e-06, 1.28316e-05, 9.238175e-06, 
    1.423202e-06, 3.864123e-07, 1.674765e-06, 2.289295e-06, 2.220255e-06,
  3.803916e-05, 2.679455e-05, 1.709909e-05, 7.768039e-06, 4.523618e-06, 
    2.01426e-06, 3.734376e-06, 2.652005e-06, 1.118229e-06, 1.641779e-06, 
    9.941945e-07, 1.318152e-06, 6.676422e-06, 6.72483e-06, 2.84363e-06,
  3.887402e-05, 3.898483e-05, 2.520305e-05, 1.005716e-05, 4.871879e-06, 
    1.7516e-06, 1.563863e-06, 1.951823e-06, 1.850995e-06, 8.076502e-07, 
    7.973737e-07, 3.836462e-06, 9.452622e-06, 7.071502e-06, 2.533354e-06,
  3.634424e-05, 4.086846e-05, 2.373827e-05, 1.00171e-05, 7.350951e-06, 
    2.432289e-06, 1.902244e-06, 1.25948e-06, 8.820438e-07, 1.217381e-06, 
    4.050309e-06, 9.4794e-06, 9.987806e-06, 6.120271e-06, 5.163393e-06,
  2.26961e-05, 2.465637e-05, 1.502509e-05, 8.206363e-06, 3.787861e-06, 
    3.544382e-06, 2.947006e-06, 2.878321e-06, 4.304604e-06, 9.443647e-06, 
    1.674718e-05, 1.775188e-05, 1.026903e-05, 5.180252e-06, 5.46927e-06,
  8.251242e-06, 7.844588e-06, 7.819345e-06, 6.827952e-06, 3.389176e-06, 
    4.48139e-06, 7.553874e-06, 1.301371e-05, 1.835902e-05, 2.525477e-05, 
    2.709822e-05, 1.88154e-05, 7.553695e-06, 5.883565e-06, 5.267404e-06,
  2.898717e-06, 1.357256e-07, 6.958245e-08, 1.498683e-06, 9.395266e-06, 
    2.625244e-05, 4.793517e-05, 4.216493e-05, 2.572031e-05, 2.124036e-05, 
    2.918977e-05, 7.369843e-05, 7.74613e-05, 3.925146e-05, 1.843908e-05,
  7.558808e-06, 1.718726e-07, 2.851523e-07, 2.631039e-06, 9.051459e-06, 
    2.2169e-05, 4.720248e-05, 4.903386e-05, 3.50634e-05, 3.856812e-05, 
    6.266893e-05, 7.064889e-05, 4.054882e-05, 2.24851e-05, 1.129477e-05,
  2.608262e-05, 1.055124e-05, 5.150415e-06, 2.695944e-06, 3.469645e-06, 
    9.905069e-06, 3.618771e-05, 6.261298e-05, 5.257616e-05, 3.955854e-05, 
    3.326119e-05, 3.008116e-05, 2.404346e-05, 1.745535e-05, 1.385699e-05,
  3.005619e-05, 1.721676e-05, 1.112396e-05, 2.949321e-06, 3.431205e-06, 
    8.475981e-06, 1.827267e-05, 1.671576e-05, 2.145009e-05, 2.374686e-05, 
    1.599407e-05, 8.070751e-06, 7.323173e-06, 1.226444e-05, 1.313567e-05,
  2.646152e-05, 2.123364e-05, 1.226498e-05, 1.728546e-06, 2.95703e-06, 
    9.203402e-06, 6.175153e-06, 2.395293e-06, 4.217765e-06, 2.557856e-06, 
    1.47339e-06, 4.541643e-07, 3.693925e-07, 2.158342e-06, 6.016266e-06,
  3.054748e-05, 2.623643e-05, 1.834208e-05, 7.762389e-06, 4.935257e-06, 
    4.009736e-06, 4.077767e-06, 3.141953e-06, 2.297615e-06, 2.329092e-06, 
    2.088267e-06, 1.210866e-06, 3.566193e-07, 4.22934e-07, 1.829853e-06,
  2.849091e-05, 2.739203e-05, 2.336584e-05, 1.194727e-05, 6.981873e-06, 
    4.693655e-06, 1.840367e-06, 3.268515e-06, 2.995027e-06, 1.88779e-06, 
    1.866536e-06, 2.009608e-06, 9.329672e-07, 1.421984e-07, 2.09325e-06,
  2.397311e-05, 2.581124e-05, 1.230213e-05, 1.134372e-05, 8.555475e-06, 
    5.064493e-06, 8.829943e-07, 2.140609e-06, 3.618506e-06, 3.328185e-06, 
    2.81244e-06, 2.153495e-06, 7.539465e-07, 9.696142e-07, 3.112848e-06,
  1.472081e-05, 1.406697e-05, 6.995674e-06, 6.233252e-06, 5.861046e-06, 
    3.408277e-06, 2.790145e-06, 1.436311e-06, 3.554064e-06, 4.574599e-06, 
    3.799669e-06, 2.988626e-06, 3.258891e-06, 3.187959e-06, 3.916128e-06,
  3.794487e-06, 2.22587e-06, 2.022351e-06, 2.389183e-06, 5.468324e-06, 
    1.046363e-05, 1.277559e-05, 1.568698e-05, 9.398338e-06, 5.462684e-06, 
    3.713042e-06, 4.550453e-06, 3.515921e-06, 5.01868e-06, 4.296347e-06,
  5.323516e-07, 1.277419e-07, 1.644544e-06, 2.779366e-06, 3.593812e-06, 
    2.2623e-06, 1.184345e-06, 1.184347e-06, 4.142381e-06, 9.64064e-06, 
    2.005407e-05, 1.024778e-05, 4.500026e-06, 4.953749e-06, 3.961036e-06,
  3.876926e-06, 6.246534e-07, 6.358787e-07, 2.020022e-06, 1.745354e-06, 
    7.481898e-07, 5.653611e-07, 6.476265e-07, 1.395245e-06, 8.743399e-06, 
    2.0474e-05, 2.585025e-05, 6.080733e-06, 4.775279e-06, 4.319269e-06,
  1.117965e-05, 1.07573e-05, 7.46861e-06, 2.036048e-06, 6.64049e-07, 
    1.064054e-06, 3.02207e-07, 6.397585e-07, 6.841312e-07, 2.103672e-06, 
    1.675206e-05, 4.346582e-05, 2.010099e-05, 2.783993e-06, 3.076174e-06,
  1.369987e-05, 1.615334e-05, 1.430994e-05, 2.385181e-06, 1.722708e-06, 
    2.877811e-06, 5.027799e-06, 6.570021e-07, 4.258827e-07, 1.088411e-06, 
    5.50501e-06, 3.0867e-05, 4.223803e-05, 2.087944e-05, 9.370398e-06,
  1.368079e-05, 1.485728e-05, 1.297178e-05, 1.336365e-06, 2.93399e-06, 
    6.847153e-06, 8.461397e-06, 1.280995e-05, 1.196139e-05, 1.991645e-06, 
    6.985001e-06, 1.433353e-05, 3.181936e-05, 2.604738e-05, 1.770886e-05,
  1.103966e-05, 1.318467e-05, 1.050242e-05, 7.093404e-06, 6.157145e-06, 
    7.542047e-06, 1.298965e-05, 1.047669e-05, 6.346706e-06, 5.749377e-06, 
    5.252555e-06, 7.565513e-06, 1.820781e-05, 2.153951e-05, 1.751746e-05,
  6.866665e-06, 1.193934e-05, 1.190734e-05, 1.331869e-05, 1.051227e-05, 
    6.707584e-06, 1.113318e-05, 1.121063e-05, 6.362132e-06, 3.704291e-06, 
    3.727654e-06, 5.603398e-06, 1.142532e-05, 1.596005e-05, 1.626657e-05,
  5.567697e-06, 1.29756e-05, 2.23788e-05, 2.66888e-05, 1.130455e-05, 
    4.56928e-06, 8.986112e-06, 1.202879e-05, 7.521045e-06, 5.151893e-06, 
    4.120964e-06, 3.658136e-06, 8.810186e-06, 1.170538e-05, 1.624058e-05,
  1.3009e-05, 2.256759e-05, 3.963885e-05, 2.78499e-05, 6.567406e-06, 
    2.491728e-06, 9.122941e-06, 1.287135e-05, 8.972473e-06, 6.291833e-06, 
    4.350223e-06, 3.868162e-06, 5.257569e-06, 7.575064e-06, 9.833291e-06,
  2.076958e-05, 2.294534e-05, 2.222091e-05, 8.940188e-06, 1.204208e-06, 
    1.691511e-06, 8.059924e-06, 1.453837e-05, 1.022704e-05, 5.22073e-06, 
    4.976749e-06, 4.303528e-06, 4.227956e-06, 6.664054e-06, 5.534073e-06,
  3.156184e-07, 1.807282e-06, 3.808477e-06, 2.495993e-06, 1.536956e-06, 
    5.40334e-06, 1.890624e-05, 1.560808e-05, 2.781654e-06, 4.877565e-06, 
    1.467418e-05, 9.73091e-06, 3.083955e-06, 3.649606e-06, 1.111391e-05,
  1.109473e-06, 2.385802e-06, 2.106078e-06, 1.473223e-06, 2.313792e-06, 
    1.075905e-05, 2.62326e-05, 1.251777e-05, 1.539587e-06, 6.058102e-06, 
    1.124377e-05, 9.292037e-06, 2.639526e-06, 9.103175e-07, 2.71025e-06,
  1.485218e-06, 2.916562e-06, 2.63963e-06, 3.619959e-06, 8.633775e-06, 
    2.50631e-05, 2.096622e-05, 1.084777e-05, 1.131901e-06, 6.215093e-06, 
    1.148469e-05, 9.11693e-06, 3.109155e-06, 4.740142e-07, 9.75034e-08,
  1.793386e-06, 3.264255e-06, 5.083843e-06, 6.068235e-06, 2.30153e-05, 
    3.382811e-05, 2.771163e-05, 3.728297e-06, 5.117324e-07, 5.346499e-06, 
    1.080153e-05, 1.092712e-05, 6.84836e-06, 2.687164e-06, 1.443574e-07,
  2.0328e-06, 3.284924e-06, 6.291843e-06, 1.031499e-05, 3.816497e-05, 
    3.892391e-05, 1.070317e-05, 2.735153e-06, 6.280241e-06, 5.040283e-06, 
    1.104317e-05, 9.732056e-06, 1.413611e-05, 9.937722e-06, 4.742109e-06,
  2.797538e-06, 4.239166e-06, 6.940984e-06, 2.478969e-05, 4.472362e-05, 
    2.620594e-05, 5.022292e-06, 2.088542e-06, 2.457344e-06, 5.733789e-06, 
    5.627317e-06, 7.49123e-06, 1.174361e-05, 1.94632e-05, 2.184172e-05,
  7.579746e-06, 6.419939e-06, 1.400986e-05, 4.066253e-05, 3.627884e-05, 
    6.666571e-06, 1.907922e-06, 3.543454e-06, 4.33141e-06, 5.16989e-06, 
    5.057566e-06, 5.865274e-06, 7.341663e-06, 1.611346e-05, 3.272553e-05,
  1.037792e-05, 1.147903e-05, 2.047236e-05, 3.02731e-05, 1.18384e-05, 
    3.225928e-07, 1.020043e-06, 4.704448e-06, 3.704356e-06, 4.49757e-06, 
    5.267837e-06, 5.125835e-06, 6.293076e-06, 9.224111e-06, 2.148271e-05,
  1.290395e-05, 1.217902e-05, 8.397769e-06, 5.692709e-06, 1.035192e-06, 
    9.06909e-08, 2.641946e-06, 5.693264e-06, 6.326152e-06, 5.144697e-06, 
    5.554875e-06, 4.600591e-06, 7.124866e-06, 7.713465e-06, 1.018028e-05,
  5.731024e-06, 5.556336e-06, 3.141272e-06, 1.402443e-06, 1.059724e-06, 
    1.429849e-07, 3.54666e-06, 7.389069e-06, 8.435556e-06, 4.354943e-06, 
    4.437004e-06, 3.443902e-06, 8.486231e-06, 7.837415e-06, 8.496941e-06,
  1.543435e-06, 2.992006e-06, 5.688071e-06, 7.348355e-06, 7.208627e-06, 
    1.062819e-05, 9.920059e-06, 7.316326e-06, 5.313528e-06, 1.480563e-06, 
    8.239836e-07, 4.082977e-06, 3.325903e-06, 5.521421e-07, 2.083148e-06,
  2.118912e-06, 5.076282e-06, 6.902759e-06, 5.965581e-06, 5.025163e-06, 
    6.528333e-06, 6.376831e-06, 3.224033e-06, 2.701555e-06, 8.132173e-07, 
    7.604668e-07, 4.780743e-06, 5.446217e-06, 4.082616e-06, 1.110587e-06,
  3.324517e-06, 4.685681e-06, 5.6463e-06, 4.135304e-06, 2.035418e-06, 
    5.215838e-06, 2.293768e-06, 2.947083e-06, 7.330193e-07, 3.80613e-07, 
    1.087998e-06, 4.415562e-06, 7.34359e-06, 8.922819e-06, 5.602761e-06,
  3.542878e-06, 5.473011e-06, 5.210865e-06, 2.051257e-06, 5.475555e-07, 
    7.967345e-07, 1.021923e-06, 1.095975e-06, 3.209103e-07, 6.213775e-07, 
    6.349459e-07, 3.836683e-06, 1.065308e-05, 1.251287e-05, 7.600436e-06,
  3.680271e-06, 3.480943e-06, 2.131875e-06, 6.486439e-07, 7.430297e-07, 
    1.303543e-06, 2.02777e-06, 2.455876e-06, 2.057217e-06, 1.147098e-06, 
    5.751916e-06, 4.154211e-06, 8.738986e-06, 1.305961e-05, 1.336543e-05,
  8.344194e-06, 4.390176e-06, 4.389308e-06, 2.498998e-06, 1.365588e-06, 
    2.101776e-06, 4.046542e-06, 4.479223e-06, 4.776629e-06, 2.696555e-06, 
    4.073824e-06, 1.861382e-06, 9.150152e-06, 1.297634e-05, 1.151874e-05,
  7.582512e-06, 8.601054e-06, 1.195515e-05, 7.924447e-06, 3.328704e-06, 
    2.349566e-06, 4.116174e-06, 5.963641e-06, 7.375565e-06, 6.737183e-06, 
    7.047554e-06, 2.648663e-06, 1.032465e-05, 1.149508e-05, 1.167878e-05,
  1.07683e-05, 1.150683e-05, 1.017349e-05, 1.220003e-05, 3.887095e-06, 
    1.515062e-06, 4.064539e-06, 5.93732e-06, 4.892334e-06, 7.734679e-06, 
    6.948925e-06, 5.350943e-06, 9.208563e-06, 9.549319e-06, 1.358778e-05,
  1.173609e-05, 1.43891e-05, 6.674452e-06, 1.264869e-05, 7.791195e-06, 
    1.095246e-06, 3.278209e-06, 7.646722e-06, 5.042938e-06, 6.55714e-06, 
    1.01525e-05, 8.209398e-06, 1.119622e-05, 1.298343e-05, 1.111334e-05,
  6.639925e-06, 6.761882e-06, 6.656212e-06, 1.10782e-05, 8.05979e-06, 
    7.406612e-07, 3.617925e-06, 1.002968e-05, 8.472523e-06, 7.362145e-06, 
    1.029738e-05, 9.979448e-06, 1.352283e-05, 1.19502e-05, 4.452745e-06,
  3.215561e-07, 2.049615e-07, 1.09823e-06, 4.217547e-06, 1.008369e-05, 
    7.587405e-06, 1.407202e-06, 2.149964e-06, 3.373489e-06, 5.395998e-06, 
    5.635868e-06, 5.075245e-06, 6.816713e-06, 5.009585e-06, 5.985041e-06,
  1.42725e-07, 8.464364e-07, 3.521363e-06, 1.386715e-05, 1.957349e-05, 
    1.212835e-05, 2.247518e-06, 5.933703e-07, 1.705629e-06, 3.798267e-06, 
    5.780422e-06, 7.845866e-06, 6.828348e-06, 6.862384e-06, 5.004872e-06,
  6.646462e-07, 3.289919e-06, 7.186494e-06, 1.754973e-05, 1.992434e-05, 
    1.637798e-05, 1.284353e-06, 8.500168e-07, 2.047139e-06, 2.119529e-06, 
    3.675501e-06, 9.123585e-06, 9.501859e-06, 8.948919e-06, 6.656277e-06,
  1.220261e-06, 3.689985e-06, 1.199091e-05, 2.12032e-05, 1.917678e-05, 
    9.321382e-06, 4.747669e-06, 5.176364e-07, 1.74738e-06, 5.477984e-06, 
    8.154086e-06, 8.883001e-06, 9.441746e-06, 5.856224e-06, 6.998355e-06,
  2.722694e-06, 5.738849e-06, 1.726977e-05, 2.401865e-05, 1.436975e-05, 
    4.76159e-06, 4.966053e-06, 7.16611e-06, 1.220599e-05, 7.358246e-06, 
    1.226996e-05, 7.429725e-06, 7.505235e-06, 3.451752e-06, 7.68579e-06,
  4.740108e-06, 6.953398e-06, 1.777113e-05, 1.980248e-05, 1.020475e-05, 
    3.285646e-06, 3.275134e-06, 6.449662e-06, 8.743288e-06, 8.059457e-06, 
    9.291128e-06, 8.199452e-06, 8.079075e-06, 8.303552e-06, 7.174278e-06,
  6.195709e-06, 5.925664e-06, 1.076247e-05, 1.418046e-05, 7.500093e-06, 
    2.659126e-06, 1.687099e-06, 5.864336e-06, 5.820405e-06, 8.107652e-06, 
    8.390381e-06, 8.26736e-06, 1.052028e-05, 1.122275e-05, 9.616949e-06,
  1.00384e-05, 5.380807e-06, 5.975739e-06, 4.954682e-06, 4.987147e-06, 
    1.16215e-06, 2.052053e-06, 4.981421e-06, 5.626207e-06, 9.050165e-06, 
    9.793655e-06, 1.337881e-05, 1.675383e-05, 1.600675e-05, 1.371636e-05,
  1.345146e-05, 5.611921e-06, 2.884998e-06, 3.506012e-06, 2.883068e-06, 
    7.580072e-07, 2.925286e-06, 4.460692e-06, 5.053355e-06, 7.386171e-06, 
    1.088366e-05, 1.693357e-05, 2.202123e-05, 2.303777e-05, 2.277378e-05,
  1.065421e-05, 7.786193e-06, 1.653294e-06, 3.117382e-06, 4.938846e-07, 
    8.283479e-07, 2.446548e-06, 6.464751e-06, 5.981298e-06, 5.231069e-06, 
    7.713187e-06, 1.46416e-05, 2.35733e-05, 2.920553e-05, 3.863197e-05,
  8.713056e-07, 3.954883e-06, 6.830134e-06, 7.684704e-06, 7.732163e-06, 
    9.361038e-06, 7.482475e-06, 3.003411e-06, 1.450124e-06, 2.861144e-06, 
    4.800856e-06, 5.6202e-06, 8.911518e-06, 7.826965e-06, 6.687508e-06,
  1.131194e-06, 3.136627e-06, 4.462481e-06, 4.778419e-06, 3.399985e-06, 
    4.025989e-06, 3.339464e-06, 8.293194e-07, 5.893386e-07, 1.085762e-06, 
    4.296339e-06, 8.350937e-06, 8.210082e-06, 1.242846e-05, 6.363053e-06,
  2.485856e-06, 2.826721e-06, 4.358097e-06, 2.771756e-06, 7.270388e-07, 
    2.617711e-06, 3.009385e-07, 1.251122e-06, 1.336609e-06, 4.956204e-06, 
    7.996295e-06, 1.013023e-05, 9.430782e-06, 1.084886e-05, 9.6763e-06,
  3.743073e-06, 2.305869e-06, 6.004716e-06, 1.76225e-06, 9.05417e-07, 
    1.503785e-06, 2.497504e-06, 3.455023e-07, 6.267672e-07, 1.646435e-06, 
    7.793597e-06, 1.14632e-05, 1.205789e-05, 1.196875e-05, 1.426607e-05,
  7.599352e-06, 3.445971e-06, 6.539876e-06, 1.476099e-06, 2.474324e-07, 
    2.402804e-06, 1.897871e-06, 5.197558e-06, 7.976014e-06, 1.832977e-06, 
    1.143505e-05, 1.004454e-05, 1.255554e-05, 1.242007e-05, 1.335429e-05,
  1.064481e-05, 3.519277e-06, 5.536758e-06, 2.249839e-06, 2.542722e-06, 
    1.607096e-06, 9.395628e-07, 9.723568e-07, 1.661518e-06, 4.196352e-06, 
    1.026087e-05, 1.202447e-05, 1.208792e-05, 1.364161e-05, 1.335686e-05,
  9.970053e-06, 3.715864e-06, 5.727615e-06, 2.113938e-06, 2.740554e-06, 
    9.714699e-07, 3.193143e-07, 8.108063e-07, 8.00518e-07, 2.142213e-06, 
    5.567463e-06, 1.194963e-05, 1.005626e-05, 1.189651e-05, 1.190699e-05,
  1.380317e-05, 3.951166e-06, 3.398557e-07, 2.76038e-06, 2.622786e-06, 
    1.413825e-06, 1.557217e-07, 2.661444e-07, 6.877062e-07, 1.360234e-06, 
    2.317289e-06, 1.045231e-05, 1.013445e-05, 1.301333e-05, 1.029672e-05,
  1.497143e-05, 4.21616e-06, 1.957247e-07, 1.077453e-06, 3.228658e-06, 
    9.361463e-07, 2.260387e-07, 2.467196e-07, 4.737921e-07, 7.546746e-07, 
    1.169522e-06, 6.708837e-06, 1.393417e-05, 1.487375e-05, 2.319506e-05,
  1.155281e-05, 5.454936e-06, 7.921876e-07, 9.157948e-07, 3.819666e-06, 
    2.826215e-06, 2.458816e-07, 4.678452e-07, 2.649e-07, 4.283511e-07, 
    8.023864e-07, 3.631927e-06, 1.367452e-05, 1.563034e-05, 2.782737e-05,
  1.755342e-07, 3.693575e-08, 1.885437e-07, 7.12518e-08, 7.839323e-08, 
    1.153617e-07, 3.756604e-07, 2.201743e-07, 1.646792e-07, 9.542601e-07, 
    1.534558e-06, 8.300324e-07, 4.097426e-06, 5.851371e-06, 5.770988e-06,
  6.078334e-07, 1.401939e-07, 8.603056e-08, 1.242806e-07, 1.170803e-07, 
    1.738134e-07, 1.628842e-07, 2.527306e-07, 1.302392e-07, 1.221857e-07, 
    4.17927e-07, 2.283653e-06, 1.709856e-06, 5.726914e-06, 4.167016e-06,
  1.34336e-06, 1.735068e-06, 1.811736e-06, 9.192192e-07, 3.916518e-07, 
    6.76639e-07, 5.152517e-07, 2.343245e-07, 1.70104e-07, 2.08597e-07, 
    3.414819e-07, 1.609587e-06, 4.333059e-06, 6.224974e-06, 5.628613e-06,
  1.486276e-06, 4.192633e-06, 8.552086e-06, 4.656338e-06, 2.678532e-06, 
    1.433068e-06, 2.069253e-06, 4.22362e-07, 9.788252e-08, 3.873157e-07, 
    7.073596e-07, 1.957204e-06, 3.780631e-06, 6.101679e-06, 9.189072e-06,
  1.090016e-06, 5.950302e-06, 1.074602e-05, 7.50811e-06, 5.407789e-06, 
    5.103831e-06, 6.57358e-06, 4.924271e-06, 7.018867e-07, 1.350637e-06, 
    3.61635e-06, 3.883139e-06, 4.395656e-06, 5.64284e-06, 8.020791e-06,
  8.601058e-07, 7.749246e-06, 1.138645e-05, 9.781375e-06, 9.76143e-06, 
    9.307299e-06, 8.4825e-06, 5.000875e-06, 3.578432e-06, 6.956227e-06, 
    9.028734e-06, 7.070536e-06, 7.912556e-06, 6.301764e-06, 6.286053e-06,
  3.720542e-06, 7.930032e-06, 9.092426e-06, 5.923579e-06, 6.152767e-06, 
    6.329199e-06, 7.385226e-06, 1.052425e-05, 1.24207e-05, 1.167609e-05, 
    1.272003e-05, 9.956096e-06, 7.487959e-06, 7.223181e-06, 8.114638e-06,
  9.478859e-06, 8.69725e-06, 6.604937e-06, 4.855015e-06, 5.722913e-06, 
    6.159935e-06, 9.909905e-06, 1.240159e-05, 1.459995e-05, 1.448463e-05, 
    1.400151e-05, 9.169143e-06, 6.72277e-06, 1.057852e-05, 1.131189e-05,
  5.943016e-06, 4.651089e-06, 7.436043e-06, 6.276094e-06, 5.703423e-06, 
    7.839858e-06, 1.199107e-05, 1.630815e-05, 1.76372e-05, 1.383997e-05, 
    9.00082e-06, 7.580625e-06, 7.730479e-06, 1.167245e-05, 1.867656e-05,
  2.588337e-06, 5.354013e-06, 6.7889e-06, 6.552552e-06, 6.995861e-06, 
    7.911104e-06, 1.170765e-05, 1.752873e-05, 1.537549e-05, 1.096089e-05, 
    8.005075e-06, 6.478224e-06, 4.577631e-06, 1.128874e-05, 1.930935e-05,
  3.781741e-07, 1.237963e-06, 5.5337e-06, 9.679648e-06, 1.058393e-05, 
    7.191661e-06, 2.328265e-06, 9.259577e-07, 7.80928e-07, 1.005733e-06, 
    1.394693e-06, 8.390703e-07, 1.392735e-06, 2.496672e-06, 1.073756e-06,
  6.936139e-07, 2.113649e-06, 6.35909e-06, 1.162598e-05, 8.834611e-06, 
    4.87803e-06, 2.151424e-06, 1.084619e-06, 8.616763e-07, 7.855396e-07, 
    6.258423e-07, 9.599573e-07, 2.264525e-06, 3.999279e-06, 1.839546e-06,
  1.850352e-07, 1.521264e-06, 6.811038e-06, 1.223476e-05, 1.069279e-05, 
    6.14494e-06, 1.14749e-06, 3.208836e-06, 4.374134e-06, 3.290597e-06, 
    2.217723e-06, 2.211757e-06, 3.538829e-06, 4.442336e-06, 3.524817e-06,
  1.694048e-07, 1.299836e-07, 3.713213e-06, 9.598549e-06, 9.461483e-06, 
    7.527732e-06, 1.79858e-05, 3.367695e-06, 3.23946e-06, 5.198206e-06, 
    4.276774e-06, 2.936624e-06, 4.064075e-06, 6.506683e-06, 7.591039e-06,
  1.52554e-07, 8.887751e-08, 2.168337e-06, 6.03025e-06, 7.514971e-06, 
    1.331357e-05, 2.049797e-05, 3.521379e-05, 1.578509e-05, 6.52827e-06, 
    1.206431e-05, 1.036293e-05, 1.163945e-05, 1.426775e-05, 1.852617e-05,
  9.501427e-08, 6.571656e-07, 3.393928e-06, 6.406227e-06, 5.064465e-06, 
    5.966905e-06, 1.42519e-05, 2.021734e-05, 2.37644e-05, 2.804364e-05, 
    2.054597e-05, 1.822551e-05, 2.106415e-05, 2.245636e-05, 2.640003e-05,
  1.365918e-06, 4.748534e-06, 7.796994e-06, 8.216205e-06, 7.757308e-06, 
    1.408096e-05, 2.75617e-05, 4.014324e-05, 2.618998e-05, 1.641056e-05, 
    1.529979e-05, 1.874015e-05, 2.512732e-05, 2.848938e-05, 2.984308e-05,
  2.876123e-06, 4.093572e-06, 6.365388e-06, 7.374272e-06, 1.250982e-05, 
    2.642126e-05, 2.666043e-05, 8.545364e-06, 8.934364e-06, 1.354417e-05, 
    1.51343e-05, 1.566887e-05, 1.532614e-05, 1.548521e-05, 1.512192e-05,
  2.995182e-06, 3.656126e-06, 8.103116e-06, 1.054137e-05, 1.932532e-05, 
    2.505996e-05, 5.20964e-06, 5.910249e-06, 1.246048e-05, 1.417072e-05, 
    6.100379e-06, 4.975809e-06, 6.591538e-06, 1.172803e-05, 1.399344e-05,
  7.077655e-06, 8.897893e-06, 8.415237e-06, 1.390506e-05, 1.871489e-05, 
    6.488202e-06, 4.928981e-06, 9.80918e-06, 1.600453e-05, 1.028984e-05, 
    4.527337e-06, 4.063413e-06, 7.961256e-06, 1.321169e-05, 1.408649e-05,
  4.878432e-06, 6.320469e-06, 6.645233e-06, 7.40355e-06, 1.143562e-05, 
    9.865056e-06, 9.7685e-06, 4.379702e-06, 6.862185e-06, 7.441257e-06, 
    5.191076e-06, 3.299039e-06, 5.713394e-06, 5.302712e-06, 5.915094e-06,
  3.775703e-06, 3.85386e-06, 3.991315e-06, 5.83247e-06, 6.89032e-06, 
    4.662371e-06, 4.420113e-06, 3.850755e-06, 5.443421e-06, 1.125489e-05, 
    1.485787e-05, 1.390562e-05, 9.914324e-06, 1.302014e-05, 7.436976e-06,
  1.654487e-06, 2.910497e-06, 2.908676e-06, 3.787831e-06, 6.819105e-06, 
    7.252257e-06, 1.306007e-06, 4.979522e-06, 8.458135e-06, 1.499947e-05, 
    2.029667e-05, 2.686299e-05, 2.723608e-05, 2.293644e-05, 1.785007e-05,
  2.480451e-06, 2.664902e-06, 3.16429e-06, 5.384321e-06, 4.033062e-06, 
    1.102181e-05, 1.598501e-05, 2.197985e-06, 1.291084e-05, 3.049559e-05, 
    3.208499e-05, 3.232689e-05, 3.648525e-05, 3.719882e-05, 3.418984e-05,
  4.738322e-06, 4.408664e-06, 3.481152e-06, 3.312801e-06, 8.127306e-06, 
    1.346566e-05, 1.876798e-05, 2.594959e-05, 2.752894e-05, 2.614243e-05, 
    3.204732e-05, 1.965209e-05, 1.063513e-05, 4.829596e-06, 6.84815e-06,
  6.965286e-06, 5.373375e-06, 3.910638e-06, 3.489382e-06, 8.140807e-06, 
    1.152998e-05, 2.087715e-05, 2.699587e-05, 2.297563e-05, 1.220204e-05, 
    4.237481e-06, 1.482675e-06, 5.825194e-07, 1.958806e-07, 8.853519e-07,
  9.606641e-06, 5.824074e-06, 3.878974e-06, 5.420557e-06, 3.859335e-06, 
    4.491857e-06, 5.924459e-06, 4.773492e-06, 2.766624e-06, 1.391779e-06, 
    8.925024e-07, 7.913793e-07, 9.695102e-07, 9.702567e-07, 7.744725e-07,
  8.102078e-06, 2.857011e-06, 3.44958e-06, 2.658855e-06, 1.004491e-06, 
    4.073128e-07, 2.236381e-07, 1.204115e-06, 2.519202e-06, 3.761427e-06, 
    4.252487e-06, 6.806961e-06, 7.697318e-06, 9.84108e-06, 1.06753e-05,
  8.264749e-06, 4.315871e-06, 1.116037e-06, 9.709373e-07, 1.512068e-06, 
    9.425627e-07, 8.31017e-07, 4.954389e-06, 6.418692e-06, 1.067037e-05, 
    6.201181e-06, 4.854137e-06, 8.075305e-06, 8.4648e-06, 7.691016e-06,
  7.241079e-06, 3.186321e-06, 4.590457e-07, 8.051169e-07, 6.424104e-07, 
    4.179838e-07, 2.989645e-06, 5.476466e-06, 1.440994e-05, 1.085338e-05, 
    6.913308e-06, 3.892073e-06, 6.791963e-06, 1.131631e-05, 1.012695e-05,
  2.514019e-06, 2.028581e-06, 1.528356e-06, 2.473746e-06, 4.108772e-06, 
    3.619026e-06, 1.791916e-06, 1.805208e-06, 2.437225e-06, 4.805061e-06, 
    1.284084e-05, 1.865854e-05, 2.011748e-05, 1.914101e-05, 1.981994e-05,
  2.952366e-06, 2.539735e-06, 3.709131e-07, 1.354706e-07, 1.019088e-06, 
    1.439373e-06, 1.046597e-06, 8.951375e-07, 1.736801e-06, 3.038384e-06, 
    3.29926e-06, 1.153653e-05, 1.765662e-05, 2.337819e-05, 2.366644e-05,
  5.653335e-06, 4.611266e-06, 3.360344e-06, 1.475835e-07, 5.041271e-08, 
    1.721783e-06, 6.882274e-08, 1.625781e-07, 2.367506e-06, 1.000242e-06, 
    5.540012e-07, 2.863908e-06, 6.952709e-06, 1.685214e-05, 1.707135e-05,
  7.899918e-06, 6.101635e-06, 5.828168e-06, 3.601881e-06, 1.891268e-06, 
    5.997113e-07, 3.138584e-06, 9.546986e-08, 5.538513e-07, 5.555424e-06, 
    1.409214e-06, 5.677595e-07, 5.549257e-07, 2.830157e-06, 7.967198e-06,
  7.188409e-06, 6.538898e-06, 7.197375e-06, 3.856665e-06, 3.385531e-06, 
    4.288583e-06, 3.652533e-06, 4.874527e-06, 1.343093e-05, 8.630304e-06, 
    4.783438e-06, 2.358521e-06, 2.724985e-07, 6.325507e-08, 8.04164e-07,
  9.371713e-06, 7.485931e-06, 7.000785e-06, 5.849617e-06, 4.692403e-06, 
    1.828198e-06, 4.389577e-06, 7.398023e-06, 9.798255e-06, 5.874771e-06, 
    1.371107e-06, 4.93573e-06, 3.773073e-06, 4.078771e-07, 1.45044e-07,
  7.95854e-06, 7.256165e-06, 9.175111e-06, 5.404362e-06, 5.576398e-06, 
    1.002513e-06, 3.653444e-06, 5.088924e-06, 3.545601e-06, 5.372989e-06, 
    4.72202e-06, 4.639247e-06, 8.307076e-06, 4.530646e-06, 4.183126e-07,
  7.298588e-06, 1.284558e-05, 1.08886e-05, 5.420007e-06, 5.971358e-06, 
    1.301265e-06, 5.836954e-06, 6.572974e-06, 3.421313e-06, 3.709273e-06, 
    4.334709e-06, 6.58624e-06, 6.579597e-06, 5.451142e-06, 6.063033e-06,
  1.207949e-05, 1.392345e-05, 9.280138e-06, 4.269275e-06, 8.605283e-06, 
    3.168313e-06, 5.617103e-06, 7.77081e-06, 8.829566e-06, 1.185977e-05, 
    5.445032e-06, 6.861902e-06, 4.158199e-06, 6.155454e-06, 8.272576e-06,
  1.022263e-05, 1.248589e-05, 6.898865e-06, 5.656462e-06, 1.140926e-05, 
    6.031389e-06, 6.604143e-06, 6.243949e-06, 9.002672e-06, 1.035217e-05, 
    6.630079e-06, 8.306211e-06, 1.363605e-06, 3.270536e-06, 3.502376e-06,
  3.862832e-06, 4.650759e-06, 3.768082e-06, 1.262223e-06, 3.919595e-06, 
    1.786157e-05, 2.678162e-05, 2.391565e-05, 1.413255e-05, 4.223184e-06, 
    1.083457e-06, 1.807675e-07, 9.319e-07, 4.10453e-06, 6.886479e-06,
  2.926439e-06, 3.492507e-06, 4.067575e-06, 2.95474e-06, 1.071337e-05, 
    2.066267e-05, 2.302523e-05, 2.457367e-05, 1.823842e-05, 7.629724e-06, 
    1.248147e-06, 1.711647e-07, 2.958026e-07, 2.482692e-06, 4.277709e-06,
  3.189126e-06, 3.656513e-06, 4.314562e-06, 7.878569e-06, 2.549024e-05, 
    4.898949e-05, 1.668707e-05, 3.013343e-05, 3.132698e-05, 1.508874e-05, 
    3.586172e-06, 4.282727e-07, 6.700711e-08, 8.950472e-07, 3.958863e-07,
  3.421615e-06, 4.504378e-06, 5.561319e-06, 1.621624e-05, 3.369983e-05, 
    4.639975e-05, 6.169933e-05, 2.987337e-05, 3.297358e-05, 2.503394e-05, 
    9.560295e-06, 1.013428e-06, 1.916907e-07, 1.242021e-06, 1.388064e-07,
  5.940767e-06, 5.06184e-06, 7.4186e-06, 2.084322e-05, 3.144327e-05, 
    4.736938e-05, 7.549708e-05, 8.74094e-05, 3.567924e-05, 1.914168e-05, 
    1.409155e-05, 2.182309e-06, 4.285555e-07, 1.911415e-06, 2.153766e-06,
  4.536085e-06, 3.883431e-06, 8.66048e-06, 1.754519e-05, 2.59201e-05, 
    4.882933e-05, 6.966646e-05, 6.261593e-05, 3.626464e-05, 2.218886e-05, 
    1.321459e-05, 2.073848e-06, 5.102925e-07, 7.965907e-07, 1.791912e-06,
  1.192388e-06, 3.564452e-06, 9.639432e-06, 1.623474e-05, 3.250649e-05, 
    4.036534e-05, 4.338711e-05, 4.458096e-05, 3.011992e-05, 1.476266e-05, 
    9.648266e-06, 2.889169e-06, 5.785329e-07, 8.928534e-07, 2.336401e-06,
  1.432983e-06, 4.782587e-06, 1.136311e-05, 2.373198e-05, 3.508971e-05, 
    3.306643e-05, 3.54153e-05, 3.117997e-05, 1.958219e-05, 1.016191e-05, 
    8.019207e-06, 2.931979e-06, 1.399179e-06, 3.096168e-06, 3.988133e-06,
  2.262047e-06, 5.272163e-06, 1.782321e-05, 3.132492e-05, 2.718845e-05, 
    2.433518e-05, 3.066314e-05, 2.989906e-05, 1.97521e-05, 8.996923e-06, 
    2.709129e-06, 2.213173e-06, 2.213236e-06, 2.26789e-06, 8.466697e-06,
  3.955232e-06, 1.286214e-05, 2.569641e-05, 2.970359e-05, 1.551822e-05, 
    1.776408e-05, 2.413248e-05, 2.524105e-05, 1.477588e-05, 4.193634e-06, 
    2.421665e-06, 2.968536e-06, 2.95919e-06, 2.031678e-06, 7.447518e-06,
  6.461377e-05, 6.507822e-05, 5.986479e-05, 5.402783e-05, 5.923898e-05, 
    7.78544e-05, 8.169987e-05, 7.956062e-05, 9.130304e-05, 8.39505e-05, 
    6.52397e-05, 4.943591e-05, 3.067562e-05, 9.44105e-06, 2.401593e-06,
  6.417975e-05, 2.838288e-05, 3.64703e-05, 4.607282e-05, 4.977719e-05, 
    5.512065e-05, 5.717625e-05, 5.027973e-05, 4.748543e-05, 4.472793e-05, 
    3.959297e-05, 4.082702e-05, 3.010405e-05, 1.767065e-05, 4.290698e-06,
  2.080155e-05, 1.996842e-05, 2.600208e-05, 3.275987e-05, 2.975375e-05, 
    1.682398e-05, 1.608102e-05, 3.28491e-05, 3.203885e-05, 2.561113e-05, 
    2.608112e-05, 3.18099e-05, 3.223883e-05, 1.796887e-05, 5.078018e-06,
  1.431001e-05, 1.810461e-05, 2.21465e-05, 1.681119e-05, 1.691286e-05, 
    1.393882e-05, 1.625338e-05, 6.685225e-06, 6.051623e-06, 2.285291e-05, 
    2.432314e-05, 3.395477e-05, 3.342493e-05, 1.672774e-05, 5.451942e-06,
  1.19985e-05, 1.25202e-05, 1.231426e-05, 7.662401e-06, 1.115774e-05, 
    2.306164e-05, 1.939345e-05, 1.745769e-05, 1.962989e-05, 1.309996e-05, 
    2.799822e-05, 3.817716e-05, 2.930619e-05, 1.189763e-05, 5.138241e-06,
  8.602404e-06, 7.569498e-06, 7.725691e-06, 6.356518e-06, 1.039707e-05, 
    1.316196e-05, 9.195706e-06, 9.53128e-06, 6.596741e-06, 6.205194e-06, 
    1.475851e-05, 2.616756e-05, 1.801352e-05, 8.004384e-06, 2.844504e-06,
  8.602453e-06, 7.850917e-06, 8.701125e-06, 8.911398e-06, 9.183531e-06, 
    4.35107e-06, 1.508443e-06, 4.442307e-06, 2.108636e-06, 6.207292e-07, 
    5.636314e-06, 9.130522e-06, 7.912977e-06, 5.510292e-06, 2.526419e-06,
  1.551147e-05, 1.147526e-05, 9.422093e-06, 7.659754e-06, 4.935473e-06, 
    5.208264e-06, 4.853966e-06, 5.614264e-06, 4.293328e-06, 1.399319e-06, 
    1.031833e-06, 2.490117e-06, 3.18157e-06, 3.472348e-06, 5.307211e-06,
  1.649235e-05, 9.016857e-06, 6.444661e-06, 4.607419e-06, 3.89109e-06, 
    4.377793e-06, 5.886901e-06, 7.247306e-06, 5.786321e-06, 4.678986e-06, 
    2.167106e-06, 1.601072e-06, 1.682475e-06, 2.816206e-06, 8.796897e-06,
  1.28925e-05, 8.043104e-06, 5.117885e-06, 3.741282e-06, 2.963866e-06, 
    3.137131e-06, 3.730607e-06, 5.464627e-06, 6.250188e-06, 2.74299e-06, 
    1.726156e-06, 1.451052e-06, 1.559048e-06, 3.297399e-06, 5.020292e-06,
  3.359725e-06, 6.03348e-06, 4.303819e-06, 2.324897e-06, 1.877393e-06, 
    2.273445e-06, 1.733497e-06, 2.760112e-06, 6.894362e-06, 1.721251e-05, 
    3.363118e-05, 5.572694e-05, 6.968444e-05, 5.985574e-05, 3.298965e-05,
  6.269426e-06, 5.953673e-06, 3.567141e-06, 3.205713e-06, 3.87944e-07, 
    6.184524e-07, 4.938087e-07, 1.706442e-06, 3.178325e-06, 6.164846e-06, 
    6.391213e-06, 2.096638e-05, 5.59963e-05, 6.087698e-05, 3.850452e-05,
  9.065649e-06, 1.111895e-05, 8.463851e-06, 1.475339e-06, 1.392365e-07, 
    1.356421e-06, 1.495328e-07, 1.165369e-06, 2.876144e-06, 7.954432e-06, 
    1.224587e-05, 1.298626e-05, 3.321913e-05, 6.280216e-05, 5.219805e-05,
  1.173317e-05, 1.175566e-05, 1.100042e-05, 5.118707e-06, 5.06315e-07, 
    3.477321e-07, 1.813039e-06, 1.245782e-07, 7.889429e-07, 8.33144e-06, 
    2.177875e-05, 3.236045e-05, 5.693999e-05, 7.879869e-05, 5.59507e-05,
  1.464674e-05, 1.238633e-05, 1.214291e-05, 7.160526e-06, 5.906104e-06, 
    5.965382e-06, 2.129646e-06, 5.020975e-06, 1.789345e-05, 1.041693e-05, 
    2.300761e-05, 3.717156e-05, 6.320227e-05, 6.656095e-05, 3.978308e-05,
  1.82848e-05, 1.203602e-05, 1.060639e-05, 8.487829e-06, 8.21758e-06, 
    6.613093e-06, 8.592815e-06, 8.112135e-06, 9.654927e-06, 6.554472e-06, 
    5.792043e-06, 1.707795e-05, 3.441784e-05, 3.448162e-05, 1.44177e-05,
  2.144331e-05, 1.282136e-05, 1.021438e-05, 9.254536e-06, 6.164056e-06, 
    6.230129e-06, 6.350104e-06, 8.05849e-06, 9.578451e-06, 3.372919e-06, 
    2.310569e-06, 7.019619e-06, 9.986312e-06, 9.721003e-06, 3.733622e-06,
  2.006228e-05, 1.214473e-05, 9.479532e-06, 7.323357e-06, 5.310974e-06, 
    7.037753e-06, 6.775839e-06, 7.315845e-06, 7.481306e-06, 2.933258e-06, 
    1.937417e-06, 3.005122e-06, 5.410015e-06, 5.495407e-06, 6.340781e-06,
  1.558215e-05, 1.144097e-05, 7.398492e-06, 5.335171e-06, 6.035847e-06, 
    6.778323e-06, 7.170054e-06, 9.161747e-06, 8.694434e-06, 6.543021e-06, 
    3.652082e-06, 2.354643e-06, 2.290107e-06, 2.292288e-06, 1.950452e-06,
  7.788136e-06, 8.656011e-06, 5.568119e-06, 4.62207e-06, 5.583302e-06, 
    6.06863e-06, 7.872999e-06, 1.208101e-05, 1.089694e-05, 3.422396e-06, 
    1.502841e-06, 1.160206e-06, 3.287708e-06, 1.901703e-06, 6.451165e-07,
  2.845214e-06, 5.396534e-06, 1.182744e-05, 1.489051e-05, 1.182591e-05, 
    6.380966e-06, 1.685761e-06, 1.418815e-07, 2.515129e-08, 6.231208e-06, 
    7.566636e-06, 4.726092e-06, 8.309521e-06, 5.814773e-06, 7.722375e-06,
  7.493979e-06, 4.923939e-06, 8.529282e-06, 1.007786e-05, 5.451554e-06, 
    2.708955e-06, 1.310354e-06, 1.139693e-06, 7.068342e-07, 1.77273e-06, 
    7.5666e-06, 7.090767e-06, 6.949012e-06, 1.405779e-05, 8.521966e-06,
  1.154778e-05, 1.51161e-05, 1.316927e-05, 8.123363e-06, 4.62918e-06, 
    7.193065e-06, 6.797027e-07, 3.443915e-06, 2.567739e-06, 4.539624e-06, 
    1.181261e-05, 1.470166e-05, 1.643124e-05, 1.324899e-05, 1.18981e-05,
  1.141203e-05, 2.03815e-05, 2.20015e-05, 8.394721e-06, 6.42352e-06, 
    4.948467e-06, 7.182133e-06, 1.374579e-06, 1.027474e-06, 4.633133e-06, 
    1.558213e-05, 2.54884e-05, 2.815473e-05, 2.215511e-05, 2.443428e-05,
  1.756067e-05, 1.807823e-05, 2.287497e-05, 1.179774e-05, 8.070798e-06, 
    8.225065e-06, 6.4192e-06, 8.882375e-06, 1.381452e-05, 7.287821e-06, 
    1.714361e-05, 3.233731e-05, 4.297637e-05, 4.162932e-05, 3.981017e-05,
  2.14276e-05, 2.287844e-05, 1.977942e-05, 1.505577e-05, 8.04585e-06, 
    8.874482e-06, 9.081114e-06, 4.928652e-06, 6.43767e-06, 1.076298e-05, 
    1.491195e-05, 2.751815e-05, 4.075731e-05, 4.945203e-05, 4.599309e-05,
  1.87864e-05, 1.914364e-05, 1.951267e-05, 1.264083e-05, 7.711642e-06, 
    8.659074e-06, 7.095453e-06, 6.069449e-06, 3.489412e-06, 4.612597e-06, 
    1.047411e-05, 2.019438e-05, 3.119526e-05, 3.620093e-05, 3.144771e-05,
  1.919834e-05, 1.925062e-05, 1.561718e-05, 1.04055e-05, 9.018997e-06, 
    8.798526e-06, 6.040141e-06, 3.940791e-06, 2.323787e-06, 4.173093e-06, 
    4.432208e-06, 9.502231e-06, 1.547135e-05, 1.90258e-05, 1.837428e-05,
  2.011809e-05, 1.865637e-05, 9.398602e-06, 7.82988e-06, 6.203267e-06, 
    6.613338e-06, 6.818678e-06, 8.016848e-06, 5.113476e-06, 5.978412e-06, 
    7.21035e-06, 6.778709e-06, 6.821499e-06, 1.452486e-05, 2.070841e-05,
  1.273336e-05, 1.072904e-05, 2.702808e-06, 4.456861e-06, 4.378082e-06, 
    7.166221e-06, 3.651907e-06, 1.132792e-05, 9.766618e-06, 4.985898e-06, 
    3.790623e-06, 3.759085e-06, 5.019163e-06, 7.89492e-06, 1.91533e-05,
  9.389407e-06, 4.923389e-06, 2.33367e-06, 4.257169e-06, 3.288059e-06, 
    3.417835e-06, 2.553482e-07, 3.314005e-07, 5.075444e-07, 3.560409e-06, 
    3.170666e-06, 1.799695e-06, 9.516944e-06, 3.764661e-05, 6.742976e-05,
  1.903616e-05, 4.682043e-06, 7.517605e-07, 3.709709e-06, 2.831196e-06, 
    1.754399e-06, 4.620528e-07, 1.246545e-06, 1.51343e-06, 1.349563e-06, 
    2.493294e-06, 5.077207e-06, 5.165042e-06, 1.661293e-05, 3.600595e-05,
  2.742939e-05, 4.106066e-06, 5.212498e-06, 2.359099e-06, 1.445039e-06, 
    5.325367e-06, 4.127486e-07, 5.768156e-06, 9.148152e-06, 3.978858e-06, 
    1.47957e-06, 6.947022e-06, 6.237659e-06, 8.77788e-06, 1.555931e-05,
  1.842362e-05, 4.711033e-06, 8.872401e-06, 6.503246e-06, 2.246325e-06, 
    7.116068e-07, 3.352368e-06, 2.419495e-06, 5.429523e-06, 1.107076e-05, 
    4.448295e-06, 6.391241e-06, 4.816054e-06, 3.907436e-06, 5.488695e-06,
  8.549784e-06, 6.228712e-06, 9.792414e-06, 7.274047e-06, 4.503674e-06, 
    3.079495e-06, 6.503979e-07, 6.919499e-06, 1.545094e-05, 1.870832e-05, 
    1.845104e-05, 8.897237e-06, 5.334015e-06, 5.608882e-06, 4.389419e-06,
  6.928535e-06, 6.734562e-06, 8.793344e-06, 7.602413e-06, 7.374924e-06, 
    5.326502e-06, 2.846697e-06, 4.340938e-06, 1.423411e-05, 2.739145e-05, 
    3.411393e-05, 2.248124e-05, 8.959225e-06, 2.819704e-06, 4.275845e-06,
  8.584811e-06, 8.952844e-06, 6.862953e-06, 6.645283e-06, 6.480727e-06, 
    5.409923e-06, 3.935086e-06, 4.481546e-06, 7.502397e-06, 1.95835e-05, 
    4.067889e-05, 4.866456e-05, 2.453122e-05, 1.034355e-05, 4.316948e-06,
  8.286435e-06, 1.043514e-05, 6.112895e-06, 6.029956e-06, 6.459568e-06, 
    5.812283e-06, 4.058685e-06, 4.127491e-06, 6.032338e-06, 1.231752e-05, 
    3.431906e-05, 5.859361e-05, 5.80564e-05, 2.705385e-05, 1.146482e-05,
  1.358285e-05, 5.995799e-06, 4.934856e-06, 4.691866e-06, 4.963572e-06, 
    6.269283e-06, 5.489763e-06, 6.080716e-06, 6.405039e-06, 1.056082e-05, 
    2.339522e-05, 5.37753e-05, 6.96634e-05, 5.706725e-05, 2.392282e-05,
  9.629186e-06, 4.804518e-06, 4.166627e-07, 5.699289e-06, 6.934064e-06, 
    6.763335e-06, 7.090568e-06, 1.041666e-05, 1.050823e-05, 9.015092e-06, 
    1.422628e-05, 3.322393e-05, 5.854638e-05, 6.618677e-05, 5.102866e-05,
  2.838961e-05, 4.293687e-05, 1.286352e-05, 1.923257e-07, 6.803951e-07, 
    4.265347e-07, 1.831827e-06, 3.788339e-06, 4.46395e-06, 2.998645e-06, 
    5.219167e-06, 5.09348e-06, 4.574867e-06, 2.367142e-05, 3.462048e-05,
  5.276811e-05, 4.2183e-05, 1.612191e-06, 1.562236e-08, 6.942684e-07, 
    2.055875e-07, 1.933013e-06, 4.497392e-06, 5.154453e-06, 1.362628e-06, 
    4.492301e-06, 5.068258e-06, 1.199078e-06, 9.91334e-06, 1.323074e-05,
  3.302747e-05, 8.940449e-06, 3.224037e-06, 1.143672e-06, 5.992043e-07, 
    2.544583e-06, 2.518903e-06, 2.019903e-05, 2.855547e-05, 1.228235e-05, 
    2.911834e-06, 4.834078e-06, 2.18011e-06, 1.621031e-06, 6.9292e-06,
  1.465577e-05, 8.114616e-06, 7.788531e-06, 5.097275e-06, 4.404361e-06, 
    9.917136e-07, 7.774606e-06, 1.228641e-05, 2.142596e-05, 2.506648e-05, 
    7.757378e-06, 6.512585e-06, 4.000954e-06, 3.504094e-07, 4.045992e-06,
  1.33218e-05, 1.086862e-05, 1.085247e-05, 6.340147e-06, 5.743324e-06, 
    8.077638e-06, 5.424725e-06, 1.576309e-05, 2.777896e-05, 2.954742e-05, 
    2.444868e-05, 8.265697e-06, 5.024435e-06, 6.606811e-07, 9.088951e-07,
  1.484656e-05, 9.999098e-06, 1.040249e-05, 8.48972e-06, 6.4598e-06, 
    7.052226e-06, 8.763221e-06, 1.432985e-05, 3.580184e-05, 5.419345e-05, 
    3.362312e-05, 9.54183e-06, 5.752278e-06, 2.711237e-06, 3.152865e-07,
  1.536469e-05, 1.150616e-05, 1.019974e-05, 8.377626e-06, 6.411725e-06, 
    8.383535e-06, 6.740983e-06, 8.230184e-06, 1.933781e-05, 3.111472e-05, 
    3.120402e-05, 1.597647e-05, 5.565149e-06, 5.318601e-06, 2.804229e-07,
  1.766537e-05, 1.277791e-05, 7.092728e-06, 7.165505e-06, 6.945709e-06, 
    7.831264e-06, 3.268345e-06, 2.962955e-06, 5.264912e-06, 1.278364e-05, 
    2.304449e-05, 1.729121e-05, 5.796038e-06, 2.614139e-06, 2.357514e-06,
  1.386916e-05, 8.690902e-06, 3.909901e-06, 6.233429e-06, 6.612791e-06, 
    1.767547e-06, 2.220731e-06, 5.502704e-06, 4.323792e-06, 8.566977e-06, 
    1.244704e-05, 1.878849e-05, 8.908642e-06, 2.703116e-06, 5.614037e-06,
  9.952251e-06, 7.690353e-06, 5.604056e-07, 5.931749e-06, 5.349448e-06, 
    5.528561e-07, 2.281944e-06, 6.77284e-06, 7.883456e-06, 3.596257e-06, 
    5.285882e-06, 1.168526e-05, 1.365869e-05, 8.34545e-06, 2.739745e-06,
  3.989811e-05, 2.413897e-05, 3.638578e-06, 1.412971e-07, 3.915336e-07, 
    6.779588e-07, 1.341254e-06, 1.513547e-06, 4.188093e-06, 1.050763e-05, 
    1.168858e-05, 5.694007e-06, 6.355109e-06, 7.173945e-06, 2.029438e-05,
  1.743335e-05, 8.551776e-06, 4.894281e-07, 6.508861e-07, 4.315931e-07, 
    2.564081e-07, 2.220632e-06, 2.979275e-06, 3.712224e-06, 5.289214e-06, 
    8.760476e-06, 7.598447e-06, 6.856458e-06, 6.52363e-06, 1.438404e-05,
  1.107205e-05, 1.115702e-05, 7.580691e-06, 1.912974e-06, 8.936844e-07, 
    3.027986e-06, 1.814738e-06, 1.071057e-05, 1.672846e-05, 1.359904e-05, 
    4.139702e-06, 5.128421e-06, 6.173279e-06, 3.129782e-06, 1.982566e-05,
  1.418445e-05, 1.376191e-05, 1.211515e-05, 4.69484e-06, 4.168801e-06, 
    3.490268e-06, 4.156155e-06, 5.271762e-06, 1.080165e-05, 1.153084e-05, 
    6.900013e-06, 6.217233e-06, 6.371837e-06, 2.524052e-06, 2.236203e-05,
  1.395991e-05, 1.29161e-05, 1.132093e-05, 7.142793e-06, 6.916533e-06, 
    5.377354e-06, 1.700053e-06, 1.158965e-05, 2.741596e-05, 1.307032e-05, 
    7.732603e-06, 1.040722e-05, 5.40429e-06, 6.424003e-06, 1.94738e-05,
  1.153432e-05, 1.00639e-05, 9.275299e-06, 8.227691e-06, 6.88167e-06, 
    4.941586e-06, 3.199269e-06, 5.904402e-06, 1.53815e-05, 2.094056e-05, 
    8.361374e-06, 9.122399e-06, 4.763739e-06, 5.732988e-06, 1.502902e-05,
  1.059946e-05, 9.333927e-06, 7.998836e-06, 5.684186e-06, 3.924346e-06, 
    4.906349e-06, 2.466575e-06, 2.240974e-06, 8.411208e-06, 1.114641e-05, 
    8.334076e-06, 5.215964e-06, 2.36861e-06, 5.020339e-06, 1.158219e-05,
  1.018485e-05, 6.658588e-06, 2.952958e-06, 2.154654e-06, 2.107293e-06, 
    5.886133e-06, 3.69111e-06, 1.086924e-06, 2.432814e-06, 4.880168e-06, 
    8.282212e-06, 5.362387e-06, 2.04608e-06, 4.981138e-06, 7.508297e-06,
  8.40073e-06, 8.193314e-06, 1.572888e-06, 1.034046e-06, 1.174002e-07, 
    3.282769e-06, 4.868092e-06, 7.330556e-06, 9.492485e-06, 7.399083e-06, 
    6.501946e-06, 6.270732e-06, 3.435731e-06, 2.527366e-06, 3.679643e-06,
  6.184221e-06, 4.218939e-06, 3.23161e-07, 1.341632e-06, 3.710132e-08, 
    1.931183e-06, 4.236612e-06, 1.11407e-05, 1.582171e-05, 6.908372e-06, 
    1.904617e-06, 5.834456e-06, 4.196407e-06, 1.977476e-06, 2.601492e-06,
  6.056479e-07, 2.13069e-06, 1.743898e-06, 1.623723e-06, 9.577798e-07, 
    1.132442e-06, 5.834523e-07, 3.110098e-06, 4.37123e-06, 8.45628e-06, 
    1.444106e-05, 1.066454e-05, 9.194448e-06, 1.036927e-05, 1.038049e-05,
  7.288066e-07, 9.081153e-07, 2.717202e-06, 3.832453e-06, 1.724363e-06, 
    5.163744e-07, 2.861252e-07, 2.156581e-06, 3.736128e-06, 7.83951e-06, 
    1.148922e-05, 1.038634e-05, 7.142264e-06, 1.380672e-05, 9.95038e-06,
  5.79082e-06, 8.380599e-06, 3.961726e-06, 4.848121e-06, 2.586926e-06, 
    5.379894e-06, 1.814268e-07, 2.282043e-06, 6.965292e-06, 8.364095e-06, 
    1.084264e-05, 9.994698e-06, 6.591789e-06, 7.377065e-06, 1.0306e-05,
  5.834726e-06, 1.02177e-05, 7.104295e-06, 5.410906e-06, 2.895097e-06, 
    1.199247e-06, 3.662365e-06, 7.290485e-07, 4.050084e-06, 8.606365e-06, 
    9.257197e-06, 1.191007e-05, 7.87401e-06, 4.936049e-06, 1.379013e-05,
  6.235086e-06, 8.206705e-06, 7.543603e-06, 7.477081e-06, 4.11795e-06, 
    7.256714e-06, 4.860563e-06, 1.149099e-05, 2.574859e-05, 1.045803e-05, 
    9.264287e-06, 9.072e-06, 8.422388e-06, 5.513799e-06, 1.442384e-05,
  8.136131e-06, 8.379619e-06, 6.21716e-06, 6.556558e-06, 5.108728e-06, 
    6.348198e-06, 6.423345e-06, 5.189011e-06, 6.839606e-06, 9.622095e-06, 
    8.187149e-06, 8.182608e-06, 7.771333e-06, 6.001315e-06, 1.583472e-05,
  9.020778e-06, 7.040358e-06, 2.418379e-06, 1.5075e-06, 5.519734e-06, 
    4.857622e-06, 6.885512e-06, 5.491183e-06, 4.1839e-06, 6.040667e-06, 
    8.361265e-06, 7.722088e-06, 7.352641e-06, 5.840513e-06, 1.239284e-05,
  1.056075e-05, 6.483214e-06, 2.589122e-07, 1.221089e-08, 3.927523e-06, 
    4.443479e-06, 6.89566e-06, 5.415431e-06, 4.619128e-06, 5.821777e-06, 
    7.364273e-06, 6.793421e-06, 5.745113e-06, 8.790387e-06, 1.270546e-05,
  1.00984e-05, 7.050213e-06, 3.247074e-07, 1.901261e-08, 1.323229e-06, 
    4.439068e-06, 3.230183e-06, 7.52968e-06, 1.206934e-05, 9.842935e-06, 
    7.104733e-06, 6.168612e-06, 7.793624e-06, 8.939269e-06, 1.105671e-05,
  7.285989e-06, 3.098031e-06, 2.002163e-07, 1.631011e-08, 1.977538e-06, 
    3.031299e-06, 1.109105e-06, 1.375479e-05, 1.530847e-05, 7.484025e-06, 
    8.941593e-06, 7.562183e-06, 7.559953e-06, 8.445249e-06, 8.70114e-06,
  2.611773e-07, 4.337942e-06, 4.208377e-06, 3.761073e-06, 3.420587e-06, 
    3.441579e-06, 2.771427e-06, 2.111887e-06, 8.020303e-07, 4.468932e-06, 
    8.306841e-06, 1.095987e-05, 1.570445e-05, 1.077637e-05, 1.271455e-05,
  3.698739e-06, 3.098672e-06, 3.782154e-06, 4.79585e-06, 4.257683e-06, 
    2.720651e-06, 2.047976e-06, 2.269103e-07, 3.93218e-07, 4.622375e-06, 
    7.306754e-06, 7.859457e-06, 1.648674e-05, 1.498587e-05, 1.137283e-05,
  5.801015e-06, 6.245021e-06, 3.814876e-06, 5.687535e-06, 4.479904e-06, 
    8.597227e-06, 3.61167e-07, 7.938921e-07, 2.622192e-06, 5.160054e-06, 
    5.881831e-06, 7.135762e-06, 9.404992e-06, 8.470261e-06, 9.900173e-06,
  4.196726e-06, 4.143412e-06, 7.819132e-06, 6.016027e-06, 6.031475e-06, 
    3.021594e-06, 7.449645e-06, 1.732298e-07, 1.020722e-06, 5.154212e-06, 
    7.434706e-06, 5.850917e-06, 9.010485e-06, 7.43258e-06, 9.410864e-06,
  3.742164e-06, 3.869968e-06, 6.211324e-06, 5.952541e-06, 6.554128e-06, 
    7.961448e-06, 5.141805e-06, 7.80449e-06, 1.604802e-05, 5.43488e-06, 
    8.053631e-06, 5.474173e-06, 8.599882e-06, 6.145081e-06, 7.185337e-06,
  4.679287e-06, 4.029462e-06, 4.657964e-06, 6.566689e-06, 4.325641e-06, 
    7.222531e-06, 7.503176e-06, 6.959099e-06, 6.732367e-06, 7.027473e-06, 
    8.380153e-06, 5.64817e-06, 5.447398e-06, 6.705685e-06, 5.579553e-06,
  8.35373e-06, 6.833466e-06, 4.918893e-06, 3.605372e-06, 4.410154e-06, 
    8.320009e-06, 7.291238e-06, 5.901411e-06, 5.807071e-06, 6.453925e-06, 
    6.545053e-06, 4.957339e-06, 6.123102e-06, 3.650779e-06, 6.252352e-06,
  9.46384e-06, 8.022608e-06, 1.785473e-06, 3.404444e-06, 5.111402e-06, 
    3.815979e-06, 6.557791e-06, 4.749054e-06, 3.556216e-06, 6.454394e-06, 
    3.640192e-06, 5.157017e-06, 4.744413e-06, 5.572864e-06, 8.861061e-06,
  6.687053e-06, 4.588681e-06, 8.367055e-07, 4.61829e-06, 6.218947e-06, 
    4.811147e-06, 5.28841e-06, 7.487231e-06, 8.95105e-06, 9.952866e-06, 
    8.176257e-06, 6.493965e-06, 5.119073e-06, 4.340986e-06, 5.971518e-06,
  2.835211e-06, 3.821602e-07, 1.310176e-06, 1.622634e-06, 4.511311e-06, 
    1.509542e-06, 4.347524e-06, 1.006876e-05, 1.247458e-05, 3.668493e-06, 
    6.761957e-06, 6.773733e-06, 8.315877e-06, 5.233764e-06, 6.16075e-06,
  2.095979e-06, 3.067616e-06, 4.874391e-06, 4.581895e-06, 4.768546e-06, 
    5.74298e-06, 5.780656e-06, 1.55817e-06, 2.282394e-07, 6.492478e-06, 
    9.642883e-06, 8.572297e-06, 7.311778e-06, 6.268122e-06, 7.689195e-06,
  1.884853e-06, 1.799058e-06, 4.161214e-06, 4.603378e-06, 5.485687e-06, 
    4.241877e-06, 5.149102e-06, 5.643259e-07, 8.69593e-08, 2.35404e-06, 
    6.779997e-06, 7.682668e-06, 5.645602e-06, 1.001784e-05, 1.511874e-05,
  4.578945e-06, 6.462405e-06, 3.282389e-06, 4.304963e-06, 6.035822e-06, 
    1.249601e-05, 3.871674e-06, 3.907481e-06, 1.130625e-06, 3.803997e-06, 
    5.747557e-06, 4.915524e-06, 4.7435e-06, 6.620992e-06, 1.034022e-05,
  6.652499e-06, 8.914006e-06, 7.015916e-06, 6.299372e-06, 9.344161e-06, 
    1.490736e-05, 1.909305e-05, 5.936425e-06, 3.092047e-06, 2.329433e-06, 
    5.575994e-06, 4.407123e-06, 4.990393e-06, 5.904996e-06, 9.93608e-06,
  1.199119e-05, 1.087057e-05, 1.282865e-05, 1.123883e-05, 1.225617e-05, 
    1.633364e-05, 2.244075e-05, 2.639715e-05, 1.253168e-05, 7.958913e-06, 
    8.494752e-06, 4.401197e-06, 5.165242e-06, 8.296392e-06, 3.761277e-06,
  2.163738e-05, 2.322283e-05, 1.749081e-05, 1.207661e-05, 1.397617e-05, 
    1.701125e-05, 2.309536e-05, 2.140637e-05, 1.334351e-05, 1.182065e-05, 
    7.856927e-06, 6.100754e-06, 4.734115e-06, 5.337135e-06, 4.400919e-06,
  2.735102e-05, 2.520279e-05, 1.821167e-05, 1.153253e-05, 1.695701e-05, 
    1.654068e-05, 1.796387e-05, 2.14131e-05, 2.268322e-05, 1.464193e-05, 
    6.17554e-06, 5.023048e-06, 6.000335e-06, 4.735313e-06, 5.857567e-06,
  2.422906e-05, 2.353912e-05, 1.569389e-05, 1.45913e-05, 1.707527e-05, 
    1.883429e-05, 1.906126e-05, 2.016446e-05, 1.960277e-05, 1.351131e-05, 
    8.141598e-06, 6.591441e-06, 7.015998e-06, 7.522758e-06, 7.467049e-06,
  2.085529e-05, 2.108236e-05, 8.984331e-06, 1.660191e-05, 1.680727e-05, 
    1.792167e-05, 1.928013e-05, 1.859755e-05, 1.064125e-05, 8.687392e-06, 
    4.589583e-06, 7.477478e-06, 7.65428e-06, 8.113688e-06, 6.657326e-06,
  1.721837e-05, 1.016369e-05, 8.952329e-06, 9.471502e-06, 1.12613e-05, 
    1.151969e-05, 1.411113e-05, 1.107e-05, 6.383593e-06, 5.563375e-06, 
    8.938476e-06, 1.105803e-05, 7.595227e-06, 7.015813e-06, 1.017228e-05,
  1.782578e-06, 3.22923e-06, 6.918455e-06, 6.804899e-06, 8.347937e-06, 
    9.176383e-06, 4.155751e-06, 2.951112e-06, 4.689839e-06, 8.074616e-06, 
    7.178495e-06, 6.392584e-06, 6.593618e-06, 6.771851e-06, 6.037263e-06,
  3.215257e-06, 5.725815e-06, 1.065847e-05, 1.301614e-05, 1.77361e-05, 
    1.406376e-05, 1.326245e-05, 1.195667e-05, 6.900247e-06, 4.924406e-06, 
    3.42282e-06, 4.218472e-06, 4.379473e-06, 5.771277e-06, 5.573941e-06,
  1.399526e-05, 1.933587e-05, 2.011687e-05, 2.685711e-05, 3.032076e-05, 
    2.903551e-05, 1.457189e-05, 2.40553e-05, 1.651247e-05, 6.410206e-06, 
    4.530044e-06, 4.219682e-06, 4.929037e-06, 4.007073e-06, 4.549105e-06,
  2.203258e-05, 2.631875e-05, 3.175759e-05, 2.86388e-05, 2.640731e-05, 
    2.479604e-05, 2.707212e-05, 1.199603e-05, 1.383608e-05, 1.257739e-05, 
    1.036582e-05, 6.99467e-06, 5.034933e-06, 5.500086e-06, 4.420331e-06,
  3.372532e-05, 2.374452e-05, 2.673326e-05, 1.659183e-05, 9.951003e-06, 
    9.550849e-06, 1.043408e-05, 2.519083e-05, 1.900613e-05, 1.433172e-05, 
    2.258677e-05, 1.111355e-05, 4.939542e-06, 4.883922e-06, 4.403716e-06,
  2.478356e-05, 2.00882e-05, 1.644239e-05, 1.038278e-05, 8.898221e-06, 
    1.088945e-05, 9.925691e-06, 7.520319e-06, 8.963007e-06, 9.258461e-06, 
    1.014453e-05, 8.676429e-06, 5.957372e-06, 2.675794e-06, 4.491417e-06,
  1.926636e-05, 1.917187e-05, 1.886822e-05, 8.165467e-06, 1.278935e-05, 
    1.452134e-05, 1.420452e-05, 9.85033e-06, 1.177458e-05, 5.927822e-06, 
    5.473451e-06, 1.045551e-05, 6.20706e-06, 5.628861e-07, 3.771422e-06,
  1.870147e-05, 2.218678e-05, 1.40896e-05, 8.274948e-06, 1.339558e-05, 
    1.589059e-05, 1.392011e-05, 1.453043e-05, 1.050091e-05, 4.643707e-06, 
    7.51995e-06, 9.942572e-06, 5.922609e-06, 4.098054e-06, 8.869508e-06,
  1.644109e-05, 1.476475e-05, 1.133932e-05, 5.876432e-06, 1.362282e-05, 
    1.591509e-05, 1.632928e-05, 1.792258e-05, 9.353378e-06, 4.506242e-06, 
    6.540481e-06, 8.380321e-06, 5.453115e-06, 6.010367e-06, 5.963785e-06,
  1.112557e-05, 1.159018e-05, 5.104506e-06, 7.193107e-06, 1.248466e-05, 
    1.642607e-05, 1.721589e-05, 1.790713e-05, 1.820265e-05, 8.182139e-06, 
    3.566142e-06, 1.141517e-05, 8.83361e-06, 6.150678e-06, 7.928998e-06,
  1.113531e-06, 1.029691e-07, 3.108016e-06, 1.897409e-06, 2.159002e-06, 
    2.839541e-06, 2.581419e-06, 3.057695e-06, 4.257372e-06, 7.50464e-06, 
    1.01566e-05, 1.02192e-05, 8.178878e-06, 6.02294e-06, 6.571536e-06,
  1.521334e-06, 8.371508e-07, 2.325548e-06, 1.84644e-06, 3.948257e-06, 
    5.237966e-06, 6.702269e-06, 4.989425e-06, 6.006117e-06, 9.835803e-06, 
    9.008456e-06, 8.456307e-06, 7.223276e-06, 5.353216e-06, 5.237839e-06,
  4.095622e-06, 3.728219e-06, 2.986538e-06, 3.954819e-06, 6.024413e-06, 
    1.435775e-05, 6.235713e-06, 4.19664e-06, 4.875905e-06, 7.704435e-06, 
    1.111856e-05, 9.777211e-06, 5.988908e-06, 3.489962e-06, 3.627544e-06,
  9.832254e-06, 1.293861e-05, 8.624815e-06, 7.881592e-06, 1.331988e-05, 
    1.86185e-05, 2.079032e-05, 6.284899e-06, 1.48224e-06, 5.849969e-06, 
    8.92803e-06, 9.904407e-06, 8.718639e-06, 4.275557e-06, 3.033398e-06,
  2.178335e-05, 1.008813e-05, 1.156358e-05, 8.417145e-06, 1.502638e-05, 
    2.31608e-05, 2.201376e-05, 2.019151e-05, 5.547063e-06, 1.378546e-06, 
    8.810755e-06, 8.739399e-06, 9.309953e-06, 3.948394e-06, 7.489896e-07,
  1.975764e-05, 1.515233e-05, 7.454674e-06, 1.13223e-05, 1.423967e-05, 
    1.882553e-05, 2.665962e-05, 1.46603e-05, 5.277146e-06, 1.327995e-06, 
    3.385115e-06, 9.459944e-06, 1.205812e-05, 1.853093e-06, 6.922648e-07,
  1.792643e-05, 1.59898e-05, 9.812662e-06, 1.120771e-05, 1.062295e-05, 
    1.16221e-05, 1.581112e-05, 1.861501e-05, 1.050499e-05, 6.7088e-07, 
    1.382568e-06, 1.31514e-05, 1.512929e-05, 4.767173e-07, 1.395008e-06,
  2.013841e-05, 2.21958e-05, 1.407341e-05, 1.055352e-05, 1.138855e-05, 
    1.334688e-05, 1.713566e-05, 1.063736e-05, 8.333321e-06, 1.531126e-06, 
    3.490821e-06, 1.265936e-05, 1.326678e-05, 3.75521e-07, 3.496927e-06,
  2.21475e-05, 2.183869e-05, 7.165751e-06, 7.188112e-06, 1.569237e-05, 
    1.194859e-05, 1.176899e-05, 1.409728e-05, 1.153341e-05, 8.197136e-06, 
    5.970841e-06, 1.259525e-05, 9.063008e-06, 4.314562e-07, 6.82112e-06,
  1.894101e-05, 1.562858e-05, 6.498307e-06, 6.224376e-06, 1.343714e-05, 
    1.492066e-05, 1.047722e-05, 1.300403e-05, 1.347983e-05, 9.206179e-06, 
    6.496903e-06, 1.193048e-05, 1.892327e-06, 4.85328e-07, 5.265168e-06,
  1.338008e-05, 1.322545e-05, 1.47536e-05, 1.365724e-05, 1.430145e-05, 
    5.741347e-06, 1.126747e-06, 2.276434e-06, 1.400954e-06, 1.378734e-06, 
    1.256712e-06, 1.556993e-06, 5.624585e-06, 5.090664e-06, 9.993593e-06,
  4.664325e-06, 4.018085e-06, 5.847404e-06, 9.652461e-06, 1.410705e-05, 
    1.326486e-05, 5.814594e-06, 4.912898e-06, 3.288699e-06, 2.685129e-06, 
    1.045434e-06, 8.029342e-07, 9.097098e-07, 5.326046e-06, 8.206428e-06,
  2.515197e-06, 4.940296e-06, 6.293445e-06, 9.243849e-06, 2.302832e-05, 
    4.502611e-05, 1.926744e-05, 1.75374e-05, 7.844334e-06, 5.628972e-06, 
    3.770931e-06, 1.310221e-06, 1.475646e-06, 1.876325e-06, 6.230901e-06,
  1.075402e-05, 9.283735e-06, 8.901518e-06, 6.498615e-06, 1.111579e-05, 
    2.053784e-05, 4.180365e-05, 2.619596e-05, 7.133768e-06, 8.335394e-06, 
    4.546348e-06, 1.642582e-06, 2.760889e-06, 1.668976e-06, 7.007174e-06,
  1.350217e-05, 7.549202e-06, 7.32409e-06, 2.160784e-06, 2.288017e-06, 
    1.252095e-05, 1.749264e-05, 2.820432e-05, 2.095336e-05, 2.7495e-06, 
    7.2868e-06, 1.714735e-06, 2.035854e-06, 2.498359e-06, 1.122495e-06,
  1.683163e-05, 1.454685e-05, 5.683569e-06, 5.295418e-06, 4.214345e-06, 
    1.862306e-06, 1.232847e-05, 8.709054e-06, 7.803201e-06, 3.674023e-06, 
    8.101571e-06, 4.045035e-06, 5.195822e-06, 6.994046e-07, 1.191702e-06,
  2.130992e-05, 1.880686e-05, 8.234084e-06, 4.410213e-06, 7.521577e-06, 
    9.892415e-07, 3.575002e-06, 1.011248e-05, 8.493947e-06, 2.957126e-06, 
    8.584131e-06, 4.713784e-06, 3.905498e-06, 7.184983e-07, 2.800818e-06,
  2.594156e-05, 2.084652e-05, 7.949171e-06, 4.117465e-06, 9.78106e-06, 
    4.241623e-06, 4.288946e-06, 5.524353e-06, 1.450774e-06, 3.113849e-06, 
    8.22205e-06, 4.757394e-06, 1.687705e-06, 2.973543e-06, 9.178653e-06,
  2.994456e-05, 2.574921e-05, 1.030277e-05, 9.29489e-06, 5.910275e-06, 
    1.002e-05, 1.216551e-05, 1.065707e-05, 4.779045e-06, 7.121593e-06, 
    4.790232e-06, 2.601917e-06, 6.130936e-07, 8.676553e-06, 9.026505e-06,
  2.561211e-05, 2.326172e-05, 5.299088e-06, 1.074412e-05, 8.677855e-06, 
    9.844896e-06, 1.181205e-05, 1.313489e-05, 6.024266e-06, 7.44326e-06, 
    4.555445e-06, 4.853513e-06, 4.866965e-07, 7.100963e-06, 7.215333e-06,
  3.167338e-06, 1.231235e-06, 2.935558e-07, 7.732265e-08, 7.340853e-07, 
    3.356865e-06, 5.017556e-06, 4.178977e-06, 3.261609e-06, 4.778559e-06, 
    2.022744e-06, 1.818585e-06, 2.473961e-06, 4.598301e-06, 2.020742e-05,
  1.047694e-06, 3.203615e-07, 7.57004e-08, 1.863919e-07, 5.584192e-06, 
    9.170856e-06, 8.432019e-06, 7.015666e-06, 3.304082e-06, 4.798489e-06, 
    2.82751e-06, 5.326272e-07, 8.717445e-07, 7.697642e-06, 2.603401e-05,
  2.9417e-07, 2.917097e-07, 2.075009e-07, 5.396617e-06, 9.323279e-06, 
    2.310076e-05, 1.240488e-05, 1.673812e-05, 1.000012e-05, 7.010097e-06, 
    2.775061e-06, 7.355273e-07, 1.253131e-06, 6.106121e-06, 2.098424e-05,
  1.08731e-05, 4.698024e-06, 4.478209e-06, 1.442063e-06, 7.1043e-06, 
    2.144379e-05, 2.985759e-05, 2.113099e-05, 1.188741e-05, 8.334438e-06, 
    3.420341e-06, 2.035585e-06, 1.718545e-06, 5.542941e-06, 1.477594e-05,
  1.424782e-05, 1.004057e-05, 1.371094e-05, 7.790535e-06, 2.956083e-06, 
    1.2277e-05, 1.247535e-05, 2.713626e-05, 2.111318e-05, 3.831128e-06, 
    5.221447e-06, 3.518086e-06, 1.894795e-06, 4.305618e-06, 8.801993e-06,
  1.849227e-05, 1.420247e-05, 8.19851e-06, 1.198515e-05, 6.29809e-06, 
    1.274391e-06, 1.055663e-05, 8.844759e-06, 7.445094e-06, 2.318687e-06, 
    4.904097e-06, 6.137117e-06, 4.143594e-06, 4.647893e-06, 7.835031e-06,
  1.876107e-05, 1.407945e-05, 5.750503e-06, 6.813788e-06, 1.321155e-05, 
    1.542098e-06, 4.045587e-06, 7.956153e-06, 8.024434e-06, 2.272338e-06, 
    6.652273e-06, 5.595378e-06, 7.387211e-06, 4.904846e-06, 7.982475e-06,
  2.183854e-05, 1.99401e-05, 5.50461e-06, 5.728175e-06, 9.841597e-06, 
    5.385994e-06, 3.528418e-06, 4.311667e-06, 3.07005e-06, 2.377793e-06, 
    6.136239e-06, 6.323168e-06, 2.954612e-06, 3.313041e-06, 7.894871e-06,
  2.798026e-05, 2.743454e-05, 8.273474e-06, 8.771637e-06, 4.894625e-06, 
    3.96203e-06, 4.938634e-06, 7.947272e-06, 7.534205e-06, 3.370069e-06, 
    8.410346e-06, 7.379105e-06, 1.594463e-06, 4.277339e-06, 7.113137e-06,
  3.022443e-05, 2.690999e-05, 9.369484e-06, 9.860248e-06, 5.533958e-06, 
    6.870958e-06, 1.049187e-05, 1.377318e-05, 8.839231e-06, 4.004863e-06, 
    1.322694e-05, 8.582563e-06, 1.488507e-06, 7.397462e-06, 6.212709e-06,
  2.705026e-06, 5.509025e-07, 5.167341e-07, 3.263452e-06, 2.21005e-06, 
    2.655246e-06, 3.336198e-06, 1.007403e-06, 3.306345e-06, 7.397969e-06, 
    6.833525e-06, 1.657771e-06, 2.648073e-06, 2.790493e-06, 1.337134e-05,
  2.217421e-06, 7.248319e-08, 6.554799e-07, 8.274841e-07, 6.919846e-06, 
    3.135047e-06, 3.367897e-06, 4.979512e-06, 4.940514e-06, 2.252444e-06, 
    5.297505e-06, 1.742022e-06, 1.13315e-06, 1.470647e-05, 3.466002e-05,
  1.020594e-06, 6.130541e-08, 8.123749e-08, 6.578584e-07, 1.246181e-06, 
    2.797118e-05, 3.054624e-06, 7.35909e-06, 3.530355e-06, 2.466744e-06, 
    4.595498e-06, 1.659958e-06, 3.396638e-06, 2.555001e-05, 4.20639e-05,
  7.854394e-07, 3.047339e-06, 1.012519e-05, 8.677314e-06, 5.468737e-06, 
    9.702086e-06, 3.119441e-05, 1.042654e-05, 3.41678e-06, 2.293918e-06, 
    8.789527e-07, 1.039416e-06, 1.427552e-05, 3.043073e-05, 2.813967e-05,
  9.612903e-06, 7.313115e-06, 8.749026e-06, 6.504634e-06, 4.751564e-06, 
    6.633546e-06, 8.340253e-06, 2.484023e-05, 6.669411e-06, 2.285504e-06, 
    2.546715e-06, 7.423231e-06, 3.143702e-05, 2.770609e-05, 1.010619e-05,
  1.456901e-05, 1.255861e-05, 4.216918e-06, 2.779554e-06, 3.996735e-06, 
    4.963079e-06, 9.385041e-06, 4.437075e-06, 5.877404e-06, 3.199579e-06, 
    8.614017e-06, 2.35326e-05, 3.714504e-05, 1.629694e-05, 4.179299e-06,
  1.401956e-05, 1.164742e-05, 4.646233e-06, 1.963739e-06, 5.081511e-06, 
    4.083122e-06, 6.245573e-06, 5.136423e-06, 5.23856e-06, 5.648236e-06, 
    2.179679e-05, 3.522647e-05, 2.858627e-05, 1.241017e-05, 3.893031e-06,
  1.771029e-05, 1.283893e-05, 5.842081e-06, 9.900863e-07, 9.405692e-06, 
    5.1204e-06, 9.029779e-06, 9.67828e-06, 8.319872e-06, 2.030364e-05, 
    3.698111e-05, 3.2961e-05, 2.152696e-05, 1.173722e-05, 5.940464e-06,
  1.981996e-05, 1.450448e-05, 4.332986e-06, 6.567584e-06, 1.076185e-05, 
    9.925618e-06, 1.082913e-05, 1.057583e-05, 1.429966e-05, 2.483502e-05, 
    3.033044e-05, 2.337012e-05, 1.629036e-05, 8.863473e-06, 4.115205e-06,
  1.598857e-05, 1.179625e-05, 5.821536e-06, 7.596353e-06, 7.219906e-06, 
    9.06383e-06, 9.440597e-06, 1.4108e-05, 1.440219e-05, 2.106159e-05, 
    2.274917e-05, 1.449874e-05, 8.004317e-06, 5.697449e-06, 3.120522e-06,
  9.83459e-05, 8.600657e-05, 6.056247e-05, 3.148778e-05, 2.166172e-05, 
    1.29587e-05, 8.394814e-06, 5.575288e-06, 7.284473e-06, 1.196236e-05, 
    8.232824e-06, 8.147053e-06, 1.213531e-05, 1.009125e-05, 6.123435e-06,
  8.887391e-05, 3.467713e-05, 1.065405e-05, 7.17457e-06, 1.904907e-06, 
    3.003553e-06, 4.047192e-06, 7.483589e-06, 1.086461e-05, 1.451018e-05, 
    9.743354e-06, 5.300002e-06, 4.947787e-06, 1.61653e-05, 5.748785e-06,
  1.407395e-05, 1.681872e-06, 2.181979e-07, 7.735151e-07, 1.884857e-06, 
    1.868234e-05, 4.09733e-06, 3.600416e-06, 5.920359e-06, 4.293547e-06, 
    7.639688e-06, 7.060587e-06, 7.494187e-06, 3.602851e-06, 4.136344e-06,
  6.341827e-08, 1.402778e-06, 2.272358e-06, 1.006471e-07, 5.158839e-08, 
    5.343267e-07, 2.011364e-05, 2.399097e-06, 2.090733e-06, 3.460385e-06, 
    2.596579e-06, 1.793696e-06, 1.81578e-06, 1.681128e-06, 4.335522e-06,
  4.66903e-06, 3.734839e-06, 8.434731e-06, 3.558075e-06, 1.760604e-07, 
    3.008622e-06, 7.421188e-06, 2.332532e-05, 8.932428e-06, 1.501242e-06, 
    1.273029e-06, 8.062237e-07, 8.524834e-07, 2.688192e-06, 8.200792e-06,
  6.57438e-06, 9.688406e-06, 3.516534e-06, 3.528587e-06, 4.612958e-06, 
    6.206918e-06, 7.058266e-06, 5.540864e-06, 4.017062e-06, 9.227006e-07, 
    6.222254e-07, 7.796302e-07, 5.217145e-06, 9.982228e-06, 1.120683e-05,
  7.400231e-06, 8.293876e-06, 6.52246e-06, 2.97463e-06, 5.832438e-06, 
    9.00729e-06, 8.350464e-06, 1.425896e-06, 1.442042e-06, 3.874963e-06, 
    5.196844e-06, 9.602774e-06, 1.309053e-05, 1.26223e-05, 1.091024e-05,
  1.057393e-05, 1.059877e-05, 8.606714e-06, 2.295533e-06, 7.039107e-06, 
    5.870631e-06, 3.770297e-06, 4.152185e-06, 4.658227e-06, 1.229055e-05, 
    1.566284e-05, 1.530758e-05, 1.224301e-05, 1.323733e-05, 1.394434e-05,
  1.403623e-05, 9.939935e-06, 4.946573e-06, 1.009161e-05, 1.093905e-05, 
    1.070393e-05, 1.003589e-05, 1.644451e-05, 2.626995e-05, 2.623618e-05, 
    1.888651e-05, 1.272741e-05, 1.189145e-05, 1.164125e-05, 1.240221e-05,
  9.686781e-06, 9.23746e-06, 6.624244e-06, 1.353198e-05, 1.476709e-05, 
    1.66987e-05, 2.241367e-05, 3.082293e-05, 3.159871e-05, 2.261946e-05, 
    1.551885e-05, 1.070955e-05, 1.031375e-05, 1.124889e-05, 1.057466e-05,
  9.587196e-06, 7.552876e-06, 8.060745e-06, 1.563116e-05, 3.096406e-05, 
    1.962835e-05, 1.054713e-05, 7.498156e-06, 9.033e-06, 1.492964e-05, 
    7.848799e-06, 7.153686e-06, 1.063166e-05, 1.05718e-05, 9.599272e-06,
  4.787671e-05, 4.5596e-05, 5.048017e-05, 7.78712e-05, 6.591436e-05, 
    2.93002e-05, 1.158016e-05, 8.017913e-06, 1.140831e-05, 2.368347e-05, 
    1.456639e-05, 5.079435e-06, 7.608837e-06, 1.565873e-05, 9.652244e-06,
  0.0001853494, 0.00016551, 0.0001502272, 0.0001159967, 5.652727e-05, 
    2.914749e-05, 4.248236e-06, 2.485376e-06, 1.627474e-06, 4.768667e-06, 
    7.763819e-06, 7.987446e-06, 7.131525e-06, 5.101707e-06, 7.447324e-06,
  0.0002372157, 0.0001987353, 0.0001318293, 6.254038e-05, 1.667865e-05, 
    1.059621e-05, 1.892553e-05, 7.003916e-07, 7.121612e-07, 1.33557e-06, 
    4.403883e-06, 8.592147e-06, 1.199303e-05, 9.347177e-06, 5.379097e-06,
  0.0001243226, 8.670025e-05, 3.908065e-05, 7.869057e-06, 1.625046e-06, 
    2.079536e-06, 7.328568e-06, 1.868432e-05, 9.860069e-06, 3.649432e-06, 
    6.584254e-06, 6.147208e-06, 1.105916e-05, 6.73159e-06, 4.271153e-06,
  2.90577e-05, 1.064268e-05, 2.239528e-06, 1.163224e-06, 4.35257e-07, 
    4.548715e-06, 1.014712e-05, 5.702609e-06, 7.510783e-06, 5.413701e-06, 
    4.983461e-06, 5.644318e-06, 4.255181e-06, 6.375798e-06, 5.979365e-06,
  2.712655e-06, 2.446426e-06, 8.506669e-07, 1.376108e-06, 3.403319e-06, 
    7.334986e-06, 9.281921e-06, 8.161323e-06, 6.348349e-06, 4.392113e-06, 
    6.185484e-06, 9.632561e-06, 6.703734e-06, 4.92425e-06, 4.696521e-06,
  1.601808e-06, 6.2657e-06, 6.814994e-07, 6.544915e-07, 7.74722e-06, 
    7.873925e-06, 5.020844e-06, 2.353286e-06, 3.670817e-07, 3.316751e-06, 
    3.98971e-06, 6.254033e-06, 5.571103e-06, 6.924374e-06, 7.148537e-06,
  4.063202e-06, 6.151064e-06, 2.297738e-07, 5.765382e-06, 1.065606e-05, 
    5.411837e-06, 5.915958e-07, 2.586339e-07, 3.134697e-06, 5.526545e-06, 
    5.06995e-06, 4.204615e-06, 7.259145e-06, 9.081195e-06, 9.414553e-06,
  5.901187e-06, 8.285924e-06, 4.514608e-06, 1.081144e-05, 8.690403e-06, 
    2.004875e-06, 8.480116e-07, 2.254305e-06, 6.559288e-06, 7.871101e-06, 
    4.699438e-06, 6.875561e-06, 9.454657e-06, 9.669971e-06, 1.058072e-05,
  3.568546e-06, 8.26111e-06, 7.987193e-06, 5.507056e-06, 1.029102e-05, 
    3.660446e-05, 4.707001e-05, 7.075619e-05, 0.0001199011, 0.0001488983, 
    0.0001396842, 0.0001218911, 9.484539e-05, 6.629421e-05, 3.387565e-05,
  9.218155e-06, 1.122503e-05, 8.58357e-06, 1.172148e-05, 5.635448e-05, 
    0.000117571, 0.0001281546, 0.0001654076, 0.0001716862, 0.0001481969, 
    0.0001162965, 0.0001010821, 7.325471e-05, 5.300889e-05, 2.157334e-05,
  7.979922e-06, 1.201097e-05, 3.699036e-05, 0.0001059424, 0.0001739289, 
    0.0002317273, 0.0001870005, 0.000178798, 0.0001394646, 0.0001187425, 
    8.892706e-05, 6.676853e-05, 4.681418e-05, 2.104954e-05, 9.243106e-06,
  1.313164e-05, 4.378114e-05, 0.0001020789, 0.0001571442, 0.0002049163, 
    0.0001436152, 0.0001850918, 0.0001433026, 0.0001022208, 6.103663e-05, 
    3.614201e-05, 2.312106e-05, 1.793017e-05, 1.146345e-05, 4.231832e-06,
  4.409558e-05, 9.722313e-05, 0.0001539169, 0.0001691248, 0.0001517255, 
    9.197403e-05, 3.633395e-05, 3.269333e-05, 3.605777e-05, 9.89392e-06, 
    3.678322e-06, 4.885484e-06, 6.630637e-06, 6.880437e-06, 2.511879e-06,
  0.0001301694, 0.0001481312, 0.000118559, 6.852249e-05, 3.725644e-05, 
    1.692784e-05, 3.445118e-06, 1.218507e-06, 6.219471e-07, 2.355329e-07, 
    5.869523e-07, 2.85412e-07, 5.501387e-06, 7.189607e-06, 3.425575e-06,
  8.625799e-05, 5.453044e-05, 2.686353e-05, 9.263142e-06, 2.068513e-06, 
    3.64856e-07, 7.599544e-08, 1.819801e-07, 2.970512e-06, 3.702066e-06, 
    3.290276e-06, 4.038485e-06, 7.204895e-06, 3.92659e-06, 2.951364e-06,
  2.715626e-05, 1.324635e-05, 4.85328e-06, 4.51887e-07, 1.082575e-07, 
    8.159549e-07, 3.794767e-07, 3.281727e-06, 3.918165e-06, 3.321026e-06, 
    3.285598e-06, 3.331346e-06, 5.760868e-06, 6.059668e-06, 3.821711e-06,
  1.852764e-05, 9.548067e-06, 7.036572e-07, 7.522431e-07, 2.167524e-06, 
    1.645066e-06, 2.102948e-06, 2.974133e-06, 4.606984e-06, 3.831485e-06, 
    3.69954e-06, 3.509846e-06, 4.55956e-06, 5.333847e-06, 3.835213e-06,
  1.516815e-05, 1.071506e-05, 2.989555e-06, 1.76292e-06, 4.043978e-06, 
    4.877214e-06, 4.463232e-06, 5.278631e-06, 6.226782e-06, 5.386793e-06, 
    4.844779e-06, 6.295631e-06, 5.611012e-06, 4.911853e-06, 3.764132e-06,
  1.864037e-07, 8.37636e-08, 1.599357e-07, 5.347224e-07, 2.953401e-06, 
    7.325123e-06, 1.068988e-05, 1.394263e-05, 1.424042e-05, 1.611154e-05, 
    8.798511e-06, 9.111786e-06, 2.437213e-05, 5.014108e-05, 7.534603e-05,
  2.617798e-07, 6.733438e-07, 1.474709e-06, 4.117542e-06, 9.890023e-06, 
    1.667921e-05, 2.531116e-05, 3.204885e-05, 2.937405e-05, 2.834685e-05, 
    2.594483e-05, 1.965735e-05, 2.641913e-05, 6.088919e-05, 7.129172e-05,
  2.798221e-06, 6.449861e-06, 7.264181e-06, 1.078117e-05, 1.81405e-05, 
    5.091878e-05, 5.046092e-05, 8.169937e-05, 6.424828e-05, 4.318147e-05, 
    2.64106e-05, 2.461978e-05, 2.901283e-05, 4.031639e-05, 5.393052e-05,
  1.135992e-05, 1.363341e-05, 1.860282e-05, 2.09661e-05, 3.361756e-05, 
    4.547169e-05, 0.0001173486, 6.715429e-05, 4.630395e-05, 2.932688e-05, 
    1.474123e-05, 1.814204e-05, 3.549201e-05, 5.625163e-05, 5.71764e-05,
  2.531081e-05, 3.406168e-05, 4.213412e-05, 3.773408e-05, 3.358505e-05, 
    4.177201e-05, 2.409408e-05, 2.530681e-05, 3.833271e-05, 1.024245e-05, 
    1.055454e-05, 1.711839e-05, 4.133104e-05, 5.993967e-05, 4.139381e-05,
  2.7548e-05, 3.872777e-05, 3.524408e-05, 2.264243e-05, 1.461882e-05, 
    7.99047e-06, 2.123951e-06, 9.295869e-07, 1.13813e-06, 4.557402e-06, 
    5.468539e-06, 1.521501e-05, 3.136032e-05, 3.207885e-05, 1.698028e-05,
  2.133838e-05, 1.930087e-05, 1.163292e-05, 2.234577e-06, 5.954727e-07, 
    1.102299e-07, 1.137677e-08, 2.403904e-08, 4.303616e-07, 4.587824e-06, 
    1.179572e-05, 1.624703e-05, 1.986742e-05, 1.108106e-05, 5.576657e-06,
  1.72904e-05, 1.15861e-05, 7.684321e-06, 2.703666e-06, 9.712857e-07, 
    2.835212e-08, 3.807921e-08, 4.06495e-07, 4.613568e-07, 3.12106e-06, 
    6.532793e-06, 1.161108e-05, 1.797538e-05, 1.143634e-05, 4.240003e-06,
  1.630093e-05, 7.662548e-06, 7.623943e-06, 8.552048e-06, 7.25488e-06, 
    4.582305e-06, 3.749743e-06, 5.196272e-06, 3.186084e-06, 3.828278e-06, 
    7.149869e-06, 1.037165e-05, 1.054104e-05, 7.119992e-06, 8.427669e-06,
  1.644615e-05, 6.85081e-06, 6.220307e-06, 7.975323e-06, 6.710323e-06, 
    6.573245e-06, 5.468386e-06, 4.064951e-06, 4.132105e-06, 7.01453e-06, 
    9.559807e-06, 8.450765e-06, 7.165743e-06, 8.042894e-06, 7.384329e-06,
  1.138042e-05, 5.56817e-06, 9.122266e-06, 1.259913e-05, 1.587942e-05, 
    1.093583e-05, 3.799849e-06, 2.725312e-06, 4.732253e-06, 6.760184e-06, 
    5.77969e-06, 5.993655e-06, 1.043235e-05, 1.251102e-05, 1.647177e-05,
  5.520193e-05, 4.585877e-05, 4.459174e-05, 4.559851e-05, 3.95675e-05, 
    1.494856e-05, 3.703307e-06, 2.575638e-06, 4.734699e-06, 6.640323e-06, 
    1.075846e-05, 1.641598e-05, 1.639021e-05, 2.196054e-05, 1.450328e-05,
  0.0001203476, 0.0001040955, 9.111509e-05, 8.665041e-05, 4.297456e-05, 
    1.443993e-05, 2.607836e-06, 5.319735e-07, 7.146675e-07, 4.294249e-06, 
    3.06062e-06, 1.119028e-05, 2.020544e-05, 2.567252e-05, 2.217399e-05,
  0.0001187038, 0.0001124142, 0.0001061657, 7.614818e-05, 2.477719e-05, 
    3.708239e-06, 6.569343e-06, 5.044822e-07, 1.005484e-06, 2.198793e-06, 
    1.584113e-06, 3.657867e-06, 1.013808e-05, 2.760497e-05, 2.723501e-05,
  0.0001274411, 0.0001006393, 6.049286e-05, 2.393078e-05, 5.639853e-06, 
    1.174086e-06, 3.488727e-06, 9.113613e-06, 2.408612e-05, 1.665473e-06, 
    4.380242e-06, 3.148002e-06, 1.422245e-05, 3.808331e-05, 2.867619e-05,
  5.028414e-05, 3.299211e-05, 1.547025e-05, 4.212407e-06, 9.473141e-07, 
    1.380151e-07, 1.735811e-06, 1.490275e-06, 3.240406e-06, 9.327697e-07, 
    2.860622e-06, 6.083909e-06, 4.6213e-05, 6.620164e-05, 3.849351e-05,
  1.159275e-05, 1.203413e-05, 8.346166e-06, 1.36876e-06, 1.470639e-07, 
    2.092012e-07, 2.201945e-07, 1.949113e-06, 2.965999e-06, 2.670553e-07, 
    1.07682e-06, 1.575524e-05, 8.036332e-05, 9.124381e-05, 5.506205e-05,
  1.273245e-05, 1.302441e-05, 7.2412e-06, 5.77144e-06, 4.905639e-06, 
    5.171725e-06, 9.495715e-07, 5.518639e-08, 6.09943e-07, 9.772101e-08, 
    5.497273e-06, 2.737289e-05, 8.357732e-05, 7.688565e-05, 3.494373e-05,
  1.206407e-05, 7.354665e-06, 5.443977e-06, 6.80084e-06, 6.856766e-06, 
    7.747631e-06, 1.463869e-06, 2.625012e-08, 1.09243e-08, 1.58931e-07, 
    4.910929e-06, 3.451258e-05, 5.872103e-05, 3.839674e-05, 1.211809e-05,
  5.882516e-06, 7.849143e-06, 6.485119e-06, 4.28168e-06, 6.507201e-06, 
    7.287822e-06, 6.516727e-06, 1.709023e-07, 2.2631e-07, 1.062591e-06, 
    8.218265e-06, 2.693375e-05, 3.365298e-05, 1.583197e-05, 8.364146e-06,
  3.165079e-06, 9.103375e-07, 1.778623e-06, 6.165657e-06, 1.296933e-05, 
    3.068023e-05, 5.340554e-05, 6.11197e-05, 6.574106e-05, 7.411036e-05, 
    7.790417e-05, 4.300072e-05, 7.438287e-06, 2.588432e-06, 2.573285e-06,
  1.555576e-06, 2.78019e-06, 4.934564e-06, 8.203964e-06, 3.371295e-05, 
    9.2473e-05, 9.031992e-05, 9.827138e-05, 0.0001055145, 0.0001079094, 
    7.776615e-05, 2.372867e-05, 1.878905e-06, 3.561999e-06, 3.598973e-06,
  8.654672e-06, 8.653822e-06, 7.228685e-06, 1.018748e-05, 7.341924e-05, 
    0.0001445106, 0.0001562903, 0.000160857, 0.0001596773, 0.0001164821, 
    5.0183e-05, 9.221146e-06, 9.728079e-07, 1.754583e-06, 5.441277e-06,
  1.431254e-05, 1.86754e-05, 2.723506e-05, 6.879943e-05, 0.0001357163, 
    0.0001210498, 0.0001803959, 0.0001454892, 0.0001158177, 6.750024e-05, 
    2.117848e-05, 3.731695e-06, 5.253112e-07, 1.668527e-06, 9.807277e-06,
  1.71817e-05, 3.765064e-05, 6.054178e-05, 7.858438e-05, 9.91546e-05, 
    0.0001133616, 6.728398e-05, 4.625862e-05, 4.578352e-05, 1.969e-05, 
    5.342338e-06, 6.035143e-07, 9.437338e-07, 9.976063e-06, 1.831993e-05,
  9.253498e-06, 1.594937e-05, 2.170591e-05, 1.6259e-05, 1.323536e-05, 
    2.004354e-05, 2.745365e-05, 2.102762e-05, 1.24109e-05, 7.710801e-06, 
    2.245131e-06, 1.254019e-06, 1.037574e-05, 3.387492e-05, 1.298145e-05,
  5.6515e-06, 9.607707e-06, 8.662123e-06, 3.029857e-06, 4.383302e-06, 
    4.376709e-06, 6.423893e-06, 6.916751e-06, 7.637287e-06, 2.375422e-06, 
    3.671796e-07, 4.668406e-06, 1.985412e-05, 4.19953e-05, 1.60545e-05,
  8.972059e-06, 8.867404e-06, 7.674685e-06, 6.392791e-06, 7.738647e-06, 
    7.191852e-06, 3.547688e-06, 1.364822e-07, 2.132106e-06, 2.088547e-07, 
    1.922016e-06, 7.29585e-06, 1.817667e-05, 3.060889e-05, 2.239872e-05,
  8.895318e-06, 7.689549e-06, 5.746804e-06, 6.300641e-06, 5.003569e-06, 
    3.057291e-06, 2.510306e-06, 8.021405e-09, 4.841145e-09, 6.602769e-07, 
    1.75323e-06, 1.089565e-05, 1.782961e-05, 1.59243e-05, 7.311705e-06,
  5.766032e-06, 4.245308e-06, 4.929521e-06, 8.834838e-06, 8.029647e-06, 
    3.854436e-07, 1.687786e-08, 9.082076e-09, 2.276306e-08, 2.474569e-06, 
    1.372589e-05, 2.143398e-05, 1.276969e-05, 8.5473e-06, 7.510165e-06,
  2.903832e-09, 1.121875e-08, 4.457436e-07, 2.067718e-06, 1.121298e-06, 
    2.192375e-06, 1.602448e-05, 1.655637e-05, 1.842863e-05, 2.113633e-05, 
    2.852695e-05, 8.767148e-05, 0.0001302964, 7.704629e-05, 3.321464e-05,
  1.166713e-08, 5.975383e-07, 2.124015e-06, 2.098652e-06, 2.203652e-06, 
    2.418948e-06, 9.62842e-06, 2.129607e-05, 3.012862e-05, 4.042138e-05, 
    7.555514e-05, 0.0001180948, 7.448291e-05, 2.064769e-05, 3.442895e-06,
  2.977203e-07, 5.391788e-06, 5.220139e-06, 2.035558e-06, 2.435185e-06, 
    9.052002e-06, 8.160486e-06, 3.758724e-05, 6.115388e-05, 8.499435e-05, 
    9.217262e-05, 6.04741e-05, 1.544273e-05, 1.320418e-06, 6.449993e-07,
  2.895787e-06, 7.217696e-06, 1.655169e-06, 4.277527e-06, 3.913024e-06, 
    3.550397e-06, 1.530105e-05, 2.543669e-05, 4.222675e-05, 5.877756e-05, 
    3.86987e-05, 1.551658e-05, 2.463847e-06, 1.535141e-06, 2.674687e-06,
  3.193757e-06, 1.468341e-06, 4.777386e-07, 4.856572e-06, 5.122322e-06, 
    5.362076e-06, 1.005824e-05, 2.02166e-05, 4.011705e-05, 3.041985e-05, 
    2.081619e-05, 8.720947e-06, 5.800341e-06, 4.419519e-06, 3.834399e-06,
  5.060083e-07, 3.929165e-07, 2.143159e-06, 4.052242e-06, 5.539242e-06, 
    6.741428e-06, 5.270555e-06, 1.367423e-05, 1.511672e-05, 1.828346e-05, 
    1.273983e-05, 6.910584e-06, 5.398105e-06, 2.827742e-06, 2.269231e-06,
  1.203553e-06, 4.877533e-06, 2.902673e-06, 4.291666e-06, 6.104857e-06, 
    5.26042e-06, 3.011865e-06, 6.068834e-06, 9.612725e-06, 9.377946e-06, 
    7.647634e-06, 5.643575e-06, 5.841728e-06, 3.655308e-06, 3.076326e-06,
  5.624937e-06, 1.130001e-05, 4.766551e-06, 8.482755e-06, 1.079171e-05, 
    7.256165e-06, 4.626218e-06, 1.332008e-06, 3.473209e-06, 5.515866e-06, 
    6.249429e-06, 4.023552e-06, 5.001848e-06, 4.047665e-06, 3.335817e-06,
  1.081226e-05, 7.262755e-06, 6.467155e-06, 8.285076e-06, 1.00601e-05, 
    5.872705e-06, 4.489558e-06, 2.947012e-07, 2.031667e-06, 6.23752e-06, 
    2.513091e-06, 2.585014e-06, 3.001436e-06, 1.965459e-06, 1.857058e-06,
  5.916047e-06, 3.533484e-06, 6.569253e-06, 1.109222e-05, 1.255683e-05, 
    7.930379e-06, 2.795286e-06, 6.694068e-08, 3.910816e-06, 5.728592e-06, 
    3.289668e-06, 8.888681e-07, 2.678575e-06, 2.658744e-06, 4.428422e-06,
  2.974041e-08, 3.68083e-08, 3.172809e-08, 9.861672e-08, 7.094177e-08, 
    1.776991e-09, 2.864215e-10, 3.234124e-08, 2.536833e-06, 9.624742e-06, 
    1.278282e-05, 6.134519e-06, 7.427691e-06, 6.724117e-06, 1.238212e-05,
  4.050195e-08, 3.280584e-08, 5.449377e-08, 2.968503e-07, 1.182564e-08, 
    7.598291e-10, 2.912559e-08, 1.901451e-07, 2.98879e-06, 9.879538e-06, 
    1.307344e-05, 7.545135e-06, 3.745638e-06, 1.469295e-05, 1.022714e-05,
  3.549271e-08, 2.382785e-06, 3.015217e-07, 2.929257e-08, 1.505426e-09, 
    1.322888e-07, 1.128732e-07, 6.301052e-07, 4.352828e-06, 1.442227e-05, 
    1.178161e-05, 7.877818e-06, 5.108652e-06, 3.65082e-06, 3.057509e-06,
  4.985417e-06, 2.771944e-07, 6.474336e-07, 5.387228e-07, 9.724633e-09, 
    3.723113e-08, 5.019743e-06, 7.631716e-07, 4.464975e-06, 1.382377e-05, 
    6.86362e-06, 8.742765e-06, 6.769612e-06, 2.182856e-06, 2.240045e-06,
  7.859078e-07, 2.149204e-07, 3.194183e-06, 1.144916e-06, 2.156149e-07, 
    1.140732e-06, 3.580804e-06, 9.803568e-06, 2.183076e-05, 1.236075e-05, 
    7.757168e-06, 6.694402e-06, 6.92234e-06, 4.160401e-06, 3.02334e-06,
  1.331102e-08, 6.866301e-07, 1.628712e-06, 5.103627e-06, 2.755854e-06, 
    4.572013e-06, 5.638502e-06, 7.382097e-06, 8.342445e-06, 1.272821e-05, 
    8.938806e-06, 7.632112e-06, 7.754479e-06, 6.922778e-06, 6.510779e-06,
  1.217519e-06, 1.339245e-06, 3.457626e-07, 4.4546e-06, 1.635169e-05, 
    1.629727e-05, 1.070615e-05, 6.838774e-06, 8.943667e-06, 1.121253e-05, 
    7.422752e-06, 5.528997e-06, 7.319448e-06, 9.26195e-06, 1.072221e-05,
  1.780451e-06, 2.458364e-06, 1.359701e-06, 1.437906e-06, 6.503934e-06, 
    1.200413e-05, 7.429603e-06, 2.36396e-06, 7.798483e-06, 9.185358e-06, 
    7.518042e-06, 5.506055e-06, 6.916037e-06, 8.910984e-06, 8.143639e-06,
  3.479413e-06, 5.038539e-06, 1.129347e-06, 1.113914e-06, 5.091847e-06, 
    7.018498e-06, 5.721068e-06, 7.043824e-07, 6.714306e-06, 8.573896e-06, 
    5.654773e-06, 5.668511e-06, 6.675195e-06, 8.856972e-06, 7.095488e-06,
  2.463273e-06, 3.524227e-06, 4.823236e-06, 1.581984e-06, 2.119675e-06, 
    1.009754e-05, 3.856446e-06, 1.611738e-06, 7.42797e-06, 6.395091e-06, 
    5.67213e-06, 6.344477e-06, 6.226019e-06, 8.091512e-06, 7.492257e-06,
  7.119082e-05, 8.905376e-06, 5.920327e-07, 8.754702e-08, 4.367596e-08, 
    3.857017e-09, 2.683423e-08, 1.001368e-08, 1.467445e-07, 6.129695e-06, 
    1.057695e-05, 1.439145e-05, 1.225828e-05, 5.3303e-06, 6.55154e-06,
  3.054627e-05, 2.725055e-06, 2.278875e-07, 3.384017e-08, 4.984615e-09, 
    2.213951e-09, 9.588241e-09, 9.715385e-08, 2.722456e-07, 7.264602e-06, 
    1.17639e-05, 1.754185e-05, 1.214942e-05, 1.159219e-05, 9.251931e-06,
  6.854327e-06, 7.924968e-07, 4.896701e-08, 7.084199e-09, 6.640707e-09, 
    1.896333e-07, 1.684528e-07, 1.27012e-06, 1.708495e-06, 7.628061e-06, 
    1.025227e-05, 1.850894e-05, 1.168471e-05, 9.991859e-06, 1.003144e-05,
  1.039388e-06, 8.907348e-08, 2.021918e-08, 9.728991e-09, 1.243943e-08, 
    2.18158e-07, 5.932581e-06, 8.476618e-07, 2.667183e-06, 6.997117e-06, 
    1.321667e-05, 1.843144e-05, 1.529798e-05, 1.065983e-05, 9.071809e-06,
  1.206672e-06, 2.547682e-06, 6.915589e-07, 1.433456e-07, 1.190273e-07, 
    1.305965e-06, 2.149003e-06, 1.992414e-05, 1.963278e-05, 4.739533e-06, 
    1.028828e-05, 1.546772e-05, 1.63235e-05, 1.272315e-05, 1.024776e-05,
  4.338297e-06, 3.25868e-06, 1.526686e-06, 1.828606e-06, 9.487197e-07, 
    2.252789e-06, 2.597748e-06, 5.999513e-06, 4.271722e-06, 8.007293e-06, 
    1.01784e-05, 1.205988e-05, 1.332345e-05, 1.203004e-05, 8.859324e-06,
  7.502979e-06, 6.636025e-06, 1.862689e-06, 2.764305e-06, 5.357752e-06, 
    4.576268e-06, 3.538135e-06, 6.588414e-06, 5.475801e-06, 7.460206e-06, 
    1.063341e-05, 1.102461e-05, 1.095012e-05, 8.604708e-06, 7.12066e-06,
  6.576747e-06, 8.754219e-06, 6.871791e-06, 1.725251e-06, 5.427681e-06, 
    3.536813e-06, 3.692096e-06, 2.24785e-06, 6.732589e-06, 8.810019e-06, 
    1.013685e-05, 1.098335e-05, 9.831836e-06, 5.909075e-06, 6.525857e-06,
  8.303829e-06, 8.286767e-06, 3.957961e-06, 2.192751e-06, 5.002963e-06, 
    6.075485e-06, 3.244034e-06, 2.841919e-06, 4.401137e-06, 1.000227e-05, 
    1.080557e-05, 1.262173e-05, 9.431063e-06, 6.514853e-06, 8.047046e-06,
  8.393482e-06, 8.227054e-06, 7.522347e-06, 5.793265e-06, 3.458457e-06, 
    4.638498e-06, 5.046668e-06, 5.661121e-06, 6.473749e-06, 7.538718e-06, 
    1.114515e-05, 1.204353e-05, 1.003626e-05, 8.914363e-06, 1.147573e-05,
  8.106539e-07, 1.374883e-07, 2.925999e-08, 2.613039e-08, 2.079881e-07, 
    4.079815e-07, 7.607626e-07, 1.192991e-06, 1.007046e-06, 9.792086e-06, 
    1.086052e-05, 1.582801e-05, 1.85313e-05, 1.061585e-05, 1.044649e-05,
  2.889866e-07, 3.899455e-07, 5.592565e-07, 7.378401e-07, 1.433504e-06, 
    1.357173e-06, 1.379249e-06, 1.805432e-06, 9.758523e-07, 6.595121e-06, 
    1.166942e-05, 1.83661e-05, 1.623835e-05, 2.313665e-05, 1.912296e-05,
  8.286104e-07, 1.28145e-06, 3.063568e-06, 3.763254e-06, 2.13561e-06, 
    8.434077e-06, 8.916714e-07, 1.097831e-06, 3.543963e-06, 8.950007e-06, 
    9.60748e-06, 1.928566e-05, 1.602209e-05, 1.521196e-05, 1.578794e-05,
  1.458616e-06, 2.116213e-06, 4.362954e-06, 5.694791e-06, 5.230723e-06, 
    5.566933e-06, 7.879244e-06, 9.867703e-07, 3.006491e-06, 1.158566e-05, 
    1.060288e-05, 1.786712e-05, 1.624469e-05, 1.882386e-05, 1.902209e-05,
  1.651747e-06, 6.531037e-06, 6.3391e-06, 4.41987e-06, 4.687502e-06, 
    8.058456e-06, 9.704611e-06, 1.353548e-05, 1.969906e-05, 8.701732e-06, 
    1.508783e-05, 1.460381e-05, 1.765224e-05, 1.690563e-05, 2.287203e-05,
  6.17275e-06, 1.030234e-05, 5.224456e-06, 5.26519e-06, 6.914531e-06, 
    6.675074e-06, 8.243162e-06, 5.809993e-06, 8.391604e-06, 1.381293e-05, 
    1.629746e-05, 1.511163e-05, 1.71242e-05, 1.781108e-05, 2.208649e-05,
  9.866297e-06, 1.094008e-05, 7.197146e-06, 5.424665e-06, 7.312194e-06, 
    7.515446e-06, 6.741453e-06, 7.836456e-06, 9.326747e-06, 9.874485e-06, 
    1.332607e-05, 1.726854e-05, 1.65146e-05, 1.6652e-05, 2.087971e-05,
  1.094817e-05, 9.507081e-06, 5.971923e-06, 7.463601e-06, 7.648416e-06, 
    8.464328e-06, 7.696109e-06, 5.291489e-06, 5.261831e-06, 7.959212e-06, 
    1.303238e-05, 1.718324e-05, 1.677066e-05, 1.563942e-05, 1.356164e-05,
  9.496885e-06, 8.500595e-06, 4.235576e-06, 7.103009e-06, 7.944004e-06, 
    7.988041e-06, 6.667972e-06, 5.170024e-06, 4.051111e-06, 5.913769e-06, 
    1.028561e-05, 1.210516e-05, 1.464839e-05, 1.49274e-05, 1.212624e-05,
  8.867564e-06, 4.716073e-06, 3.80421e-06, 6.288325e-06, 6.724388e-06, 
    6.82839e-06, 9.51919e-06, 8.411502e-06, 4.402285e-06, 7.073937e-06, 
    6.779591e-06, 8.357351e-06, 1.01213e-05, 1.416344e-05, 1.136958e-05,
  3.912873e-07, 1.171671e-06, 1.111175e-06, 1.526e-06, 5.021704e-06, 
    5.751e-06, 6.948166e-06, 5.204474e-06, 4.848241e-06, 4.844692e-06, 
    7.080685e-06, 1.209478e-05, 1.654732e-05, 2.10431e-05, 2.444634e-05,
  1.535228e-06, 2.439141e-06, 3.332889e-06, 4.791045e-06, 6.134288e-06, 
    3.600889e-06, 5.730121e-06, 3.004018e-06, 3.525233e-06, 2.396465e-06, 
    6.986557e-06, 1.303162e-05, 1.655154e-05, 2.401093e-05, 2.156987e-05,
  1.896278e-06, 5.493565e-06, 6.52044e-06, 6.19809e-06, 3.534597e-06, 
    1.174894e-05, 2.303367e-06, 5.810264e-06, 4.719802e-06, 4.045287e-06, 
    6.559704e-06, 1.423777e-05, 1.602781e-05, 1.707578e-05, 1.597914e-05,
  3.977482e-06, 5.262842e-06, 6.322818e-06, 7.232093e-06, 5.284339e-06, 
    6.988974e-06, 1.078588e-05, 2.561141e-06, 3.323439e-06, 3.475985e-06, 
    9.856089e-06, 1.542322e-05, 1.482621e-05, 1.270772e-05, 1.211266e-05,
  3.14157e-06, 5.334869e-06, 6.443129e-06, 7.425245e-06, 7.408913e-06, 
    7.228713e-06, 8.17782e-06, 1.438875e-05, 1.677509e-05, 2.973055e-06, 
    1.282762e-05, 1.541071e-05, 1.355551e-05, 1.023695e-05, 1.120836e-05,
  6.315623e-06, 5.696588e-06, 8.008595e-06, 6.818971e-06, 7.334378e-06, 
    8.7322e-06, 9.742149e-06, 6.930032e-06, 7.168044e-06, 8.713221e-06, 
    1.253782e-05, 1.245592e-05, 1.117562e-05, 1.143769e-05, 1.163867e-05,
  6.454849e-06, 6.386203e-06, 8.579429e-06, 5.07842e-06, 6.818642e-06, 
    8.461419e-06, 5.75271e-06, 5.910701e-06, 6.802131e-06, 5.858045e-06, 
    1.133857e-05, 1.155081e-05, 8.400769e-06, 1.260441e-05, 1.31947e-05,
  6.296748e-06, 7.659074e-06, 7.918297e-06, 6.61858e-06, 7.419943e-06, 
    8.911768e-06, 7.209273e-06, 8.658054e-06, 7.376535e-06, 7.677558e-06, 
    1.221704e-05, 1.170561e-05, 9.650424e-06, 1.149941e-05, 1.336686e-05,
  6.744105e-06, 8.329905e-06, 4.294168e-06, 5.116076e-06, 6.959245e-06, 
    1.119035e-05, 1.20066e-05, 1.401614e-05, 1.389451e-05, 1.208746e-05, 
    1.273605e-05, 1.290032e-05, 1.116189e-05, 8.994254e-06, 8.072378e-06,
  7.01052e-06, 3.746104e-06, 3.229645e-06, 3.985587e-06, 7.679111e-06, 
    1.270544e-05, 1.716967e-05, 1.856431e-05, 1.925597e-05, 2.169897e-05, 
    1.968951e-05, 1.726751e-05, 1.104212e-05, 6.849974e-06, 6.187303e-06,
  4.523477e-07, 2.84189e-06, 2.51169e-06, 3.757545e-06, 4.665817e-06, 
    6.13571e-06, 4.631884e-06, 2.764237e-06, 3.269653e-06, 4.122027e-06, 
    5.208252e-06, 7.667778e-06, 9.380826e-06, 9.772461e-06, 8.578445e-06,
  2.086102e-06, 2.096025e-06, 3.624623e-06, 5.422108e-06, 6.990754e-06, 
    3.184972e-06, 4.832053e-06, 6.425947e-06, 3.440166e-06, 3.737045e-06, 
    5.100059e-06, 6.117238e-06, 9.949886e-06, 1.270385e-05, 8.210641e-06,
  2.463082e-06, 4.246502e-06, 5.082849e-06, 6.531872e-06, 8.10859e-06, 
    1.231325e-05, 2.580346e-06, 1.208483e-05, 1.098918e-05, 6.339234e-06, 
    3.673509e-06, 5.991854e-06, 8.970118e-06, 1.04633e-05, 1.021045e-05,
  3.302465e-06, 2.751296e-06, 7.338667e-06, 8.42078e-06, 8.907754e-06, 
    1.11565e-05, 1.91425e-05, 4.459042e-06, 7.998513e-06, 9.878951e-06, 
    7.950905e-06, 6.808222e-06, 5.420949e-06, 6.892879e-06, 1.018967e-05,
  3.605105e-06, 5.478448e-06, 8.982902e-06, 7.908493e-06, 1.074535e-05, 
    1.402369e-05, 2.538685e-05, 4.375432e-05, 2.688821e-05, 8.590778e-06, 
    1.375939e-05, 9.935065e-06, 7.519395e-06, 7.45953e-06, 1.013786e-05,
  1.532759e-06, 5.983879e-06, 9.266151e-06, 5.265761e-06, 9.648394e-06, 
    1.849179e-05, 3.069185e-05, 3.63882e-05, 2.61169e-05, 2.432897e-05, 
    1.86536e-05, 1.543636e-05, 1.254694e-05, 1.174609e-05, 1.148457e-05,
  3.951091e-06, 8.851625e-06, 5.340657e-06, 5.72618e-06, 7.905971e-06, 
    1.734627e-05, 2.330589e-05, 2.787258e-05, 2.408738e-05, 1.859874e-05, 
    1.763818e-05, 2.001421e-05, 1.919391e-05, 1.702827e-05, 1.392543e-05,
  5.790321e-06, 7.530508e-06, 4.276504e-06, 5.803855e-06, 8.476391e-06, 
    1.46066e-05, 1.709709e-05, 1.760535e-05, 1.768725e-05, 1.742369e-05, 
    1.889086e-05, 1.806882e-05, 1.863872e-05, 2.002047e-05, 1.307769e-05,
  5.659839e-06, 5.389864e-06, 2.75608e-06, 3.517599e-06, 9.146994e-06, 
    1.070963e-05, 1.177676e-05, 1.223795e-05, 1.201516e-05, 1.397621e-05, 
    1.513878e-05, 1.51312e-05, 1.585053e-05, 1.385959e-05, 1.068861e-05,
  3.276266e-06, 2.714169e-06, 1.074057e-06, 1.996846e-06, 4.898937e-06, 
    7.563874e-06, 5.799611e-06, 5.19466e-06, 7.460085e-06, 1.189172e-05, 
    1.480914e-05, 1.381238e-05, 1.405627e-05, 9.950767e-06, 1.084933e-05,
  2.646972e-08, 1.061404e-06, 2.919e-06, 4.583988e-06, 6.103596e-06, 
    6.246332e-06, 4.773686e-06, 6.214832e-06, 9.048165e-06, 1.442293e-05, 
    1.413381e-05, 1.381076e-05, 9.702833e-06, 6.784684e-06, 3.246774e-06,
  6.515451e-07, 2.189315e-06, 3.955533e-06, 5.581296e-06, 7.777316e-06, 
    4.746705e-06, 5.126178e-06, 4.722572e-06, 3.747979e-06, 6.41795e-06, 
    1.32377e-05, 1.582521e-05, 1.027565e-05, 7.3985e-06, 6.26906e-06,
  3.027919e-06, 4.880542e-06, 6.570615e-06, 6.159803e-06, 7.226404e-06, 
    1.431837e-05, 7.940042e-06, 9.692099e-06, 7.314312e-06, 3.775854e-06, 
    6.21242e-06, 1.213979e-05, 1.216251e-05, 4.896308e-06, 3.8792e-06,
  1.680103e-06, 6.837982e-06, 1.018513e-05, 6.23325e-06, 7.525481e-06, 
    1.305957e-05, 2.876801e-05, 1.136175e-05, 1.19985e-05, 6.721481e-06, 
    5.372247e-06, 8.741787e-06, 1.060633e-05, 5.507269e-06, 3.65145e-06,
  4.869759e-06, 8.259743e-06, 1.11789e-05, 4.98807e-06, 7.562994e-06, 
    2.06478e-05, 2.851612e-05, 4.32679e-05, 3.050583e-05, 1.07311e-05, 
    8.622578e-06, 9.523055e-06, 6.619201e-06, 4.35488e-06, 4.570147e-06,
  5.921286e-06, 7.172615e-06, 6.075949e-06, 3.919019e-06, 1.092046e-05, 
    2.632668e-05, 3.88147e-05, 3.465027e-05, 2.011893e-05, 1.222433e-05, 
    1.233974e-05, 8.803908e-06, 8.815192e-06, 6.138552e-06, 4.599481e-06,
  5.786156e-06, 4.835401e-06, 4.483507e-06, 4.470488e-06, 1.124583e-05, 
    2.029341e-05, 3.101377e-05, 3.291586e-05, 2.02127e-05, 1.061858e-05, 
    1.478368e-05, 1.494552e-05, 8.866962e-06, 6.291075e-06, 6.007328e-06,
  4.916373e-06, 8.098643e-06, 5.766863e-06, 2.625685e-06, 1.211312e-05, 
    1.823273e-05, 2.686824e-05, 2.666355e-05, 2.127695e-05, 1.070201e-05, 
    1.120486e-05, 1.55472e-05, 7.082154e-06, 7.264041e-06, 7.199342e-06,
  2.431976e-06, 4.370297e-06, 3.051223e-06, 1.331932e-06, 9.992367e-06, 
    1.863971e-05, 2.102923e-05, 2.756272e-05, 2.385457e-05, 1.109142e-05, 
    1.127476e-05, 1.037486e-05, 5.079833e-06, 5.482505e-06, 8.635976e-06,
  2.84333e-06, 2.152823e-06, 8.249049e-07, 1.29915e-06, 9.165445e-06, 
    1.983229e-05, 2.129568e-05, 2.145857e-05, 2.654881e-05, 2.044459e-05, 
    1.422445e-05, 1.005362e-05, 4.689422e-06, 4.823833e-06, 7.665792e-06,
  5.926337e-07, 2.80349e-06, 4.26311e-06, 2.075071e-06, 1.933895e-06, 
    3.801155e-06, 4.863788e-06, 7.03756e-06, 1.403466e-05, 1.704586e-05, 
    2.218143e-05, 1.275767e-05, 6.374897e-06, 1.320499e-06, 3.151797e-06,
  3.46861e-06, 2.468169e-06, 2.774525e-06, 9.420359e-07, 3.666332e-06, 
    3.100691e-06, 7.05311e-06, 8.890293e-06, 9.244167e-06, 1.639747e-05, 
    1.474127e-05, 1.043121e-05, 7.06135e-06, 4.58399e-06, 4.106098e-06,
  3.852278e-06, 5.926252e-06, 8.000427e-06, 2.300517e-06, 5.589896e-06, 
    2.09324e-05, 7.665009e-06, 1.628302e-05, 1.289808e-05, 1.737995e-05, 
    1.317476e-05, 5.920121e-06, 8.545002e-06, 7.935485e-07, 2.159346e-06,
  5.32653e-06, 7.183799e-06, 8.877419e-06, 3.375422e-06, 6.404915e-06, 
    1.994819e-05, 3.700584e-05, 1.923286e-05, 1.693431e-05, 1.655151e-05, 
    1.458063e-05, 7.905443e-06, 7.058634e-06, 1.870239e-06, 9.40198e-07,
  6.019833e-06, 9.035482e-06, 8.037658e-06, 4.96048e-06, 5.688147e-06, 
    1.519657e-05, 2.343924e-05, 3.60018e-05, 3.060348e-05, 1.054324e-05, 
    1.042496e-05, 6.258771e-06, 3.99692e-06, 1.585641e-06, 9.085427e-07,
  6.739318e-06, 8.608006e-06, 7.546485e-06, 7.023743e-06, 5.516451e-06, 
    9.364065e-06, 1.169902e-05, 1.37007e-05, 1.109931e-05, 6.91497e-06, 
    5.751187e-06, 3.447561e-06, 2.867047e-06, 1.674084e-06, 9.574596e-07,
  8.55896e-06, 1.00457e-05, 6.099426e-06, 6.154239e-06, 3.518101e-06, 
    3.135999e-06, 4.126988e-06, 9.019202e-06, 1.20296e-05, 5.84552e-06, 
    4.642452e-06, 3.550003e-06, 2.69675e-06, 1.814982e-06, 1.047844e-06,
  9.630337e-06, 1.188102e-05, 6.228116e-06, 6.609655e-06, 5.531047e-06, 
    1.428935e-06, 2.902945e-06, 3.575277e-06, 5.204328e-06, 6.037715e-06, 
    4.579042e-06, 5.421771e-06, 2.507439e-06, 1.870058e-06, 8.969197e-07,
  1.045207e-05, 1.037252e-05, 5.965482e-06, 5.570539e-06, 4.767401e-06, 
    9.077019e-07, 1.991374e-06, 5.844438e-06, 5.476812e-06, 4.941832e-06, 
    3.098008e-06, 4.953462e-06, 2.583526e-06, 1.759212e-06, 9.265092e-07,
  9.226315e-06, 6.563863e-06, 4.310464e-06, 3.625379e-06, 4.264242e-06, 
    2.929684e-06, 2.312097e-06, 1.987934e-06, 3.457274e-06, 3.34678e-06, 
    2.940559e-06, 3.680355e-06, 1.963259e-06, 1.762059e-06, 7.340411e-07,
  7.344276e-06, 6.389371e-06, 4.672474e-06, 5.138068e-06, 8.298674e-07, 
    1.335935e-06, 2.795095e-06, 3.885406e-06, 6.941541e-06, 9.71084e-06, 
    9.675191e-06, 3.818655e-06, 1.044008e-06, 1.013216e-07, 7.132709e-06,
  1.180529e-05, 5.146307e-06, 5.083079e-06, 5.396095e-06, 2.13254e-06, 
    1.313664e-06, 2.342632e-06, 3.948339e-06, 6.899731e-06, 9.692156e-06, 
    1.037452e-05, 4.906086e-06, 6.718473e-07, 4.401666e-06, 1.922995e-05,
  1.136784e-05, 6.483189e-06, 6.982447e-06, 7.078588e-06, 9.662381e-07, 
    1.195043e-05, 9.30196e-06, 6.409212e-06, 6.782447e-06, 1.324186e-05, 
    1.041392e-05, 4.968296e-06, 7.135702e-07, 7.795095e-06, 2.90856e-05,
  8.623593e-06, 7.195693e-06, 6.398568e-06, 6.458414e-06, 1.636325e-06, 
    6.006665e-06, 2.700777e-05, 1.524917e-05, 7.555918e-06, 1.790037e-05, 
    1.171647e-05, 5.802456e-06, 2.587439e-06, 1.552161e-05, 2.917876e-05,
  9.550244e-06, 6.896942e-06, 7.344362e-06, 4.90222e-06, 1.902663e-06, 
    3.371019e-06, 3.430805e-06, 2.117881e-05, 3.096764e-05, 1.405821e-05, 
    1.068054e-05, 4.752599e-06, 8.375962e-06, 2.973047e-05, 3.180407e-05,
  9.570016e-06, 8.584212e-06, 6.988756e-06, 3.508608e-06, 1.921092e-06, 
    3.923961e-07, 2.318787e-06, 6.187534e-06, 6.559841e-06, 8.436266e-06, 
    7.462107e-06, 4.78924e-06, 2.391591e-05, 4.501179e-05, 1.805565e-05,
  1.090533e-05, 8.029598e-06, 5.552262e-06, 2.70247e-06, 2.095837e-06, 
    2.839586e-06, 2.45448e-06, 6.28713e-06, 1.549179e-05, 1.031383e-05, 
    8.507224e-06, 2.189135e-05, 4.764558e-05, 4.418943e-05, 2.007477e-05,
  1.003507e-05, 9.480201e-06, 1.93476e-06, 1.60456e-06, 4.725126e-06, 
    3.748888e-06, 4.75888e-06, 1.012375e-05, 1.278897e-05, 1.460423e-05, 
    2.497565e-05, 4.044253e-05, 4.487316e-05, 2.450953e-05, 1.328316e-05,
  1.176642e-05, 5.682937e-06, 1.472846e-06, 3.464019e-06, 3.825111e-06, 
    5.340075e-06, 9.388621e-06, 1.391331e-05, 1.749319e-05, 2.164264e-05, 
    2.487938e-05, 2.607317e-05, 1.955969e-05, 9.470165e-06, 6.618184e-06,
  8.996812e-06, 7.258453e-06, 1.932129e-06, 3.060662e-06, 4.913995e-06, 
    6.73109e-06, 9.8066e-06, 9.060047e-06, 1.025783e-05, 1.556542e-05, 
    1.652353e-05, 1.485053e-05, 1.21573e-05, 7.876954e-06, 6.023457e-06,
  7.895542e-06, 6.709738e-06, 5.401867e-06, 5.575598e-06, 8.00717e-06, 
    8.026652e-06, 2.689595e-06, 2.497016e-06, 2.38503e-06, 1.380975e-06, 
    1.128247e-06, 5.439954e-07, 2.62303e-06, 3.840762e-08, 1.629724e-06,
  2.453137e-05, 1.273342e-05, 1.026212e-05, 9.885386e-06, 6.544662e-06, 
    2.963733e-06, 2.094437e-06, 2.277457e-06, 1.178645e-06, 1.63694e-06, 
    3.158834e-06, 4.099679e-06, 7.278701e-09, 7.264836e-07, 7.548731e-06,
  8.264324e-05, 4.1757e-05, 1.573469e-05, 7.023224e-06, 3.821232e-06, 
    3.178838e-06, 3.61398e-06, 1.32324e-06, 1.471225e-06, 1.572186e-06, 
    1.686653e-06, 2.155909e-06, 2.599735e-08, 5.876609e-07, 1.868363e-05,
  8.311804e-05, 3.066171e-05, 6.643072e-06, 3.492285e-06, 4.084097e-06, 
    3.614534e-06, 1.298233e-05, 1.317068e-05, 3.10366e-06, 1.608414e-06, 
    1.06663e-06, 6.310058e-07, 5.874281e-08, 1.742092e-06, 2.041106e-05,
  2.395574e-05, 7.261128e-06, 4.782446e-06, 3.944346e-06, 4.055746e-06, 
    4.958363e-06, 1.307482e-06, 2.746211e-05, 1.555009e-05, 2.020484e-06, 
    1.400563e-06, 8.305323e-07, 4.429626e-07, 6.453301e-06, 1.713445e-05,
  8.760189e-06, 9.93956e-06, 6.474291e-06, 4.599454e-06, 5.151265e-07, 
    1.642915e-06, 3.171521e-06, 1.69121e-06, 1.218961e-06, 6.620139e-07, 
    1.741478e-07, 3.663247e-07, 4.079476e-06, 1.769048e-05, 3.901438e-06,
  1.009894e-05, 1.024832e-05, 5.47468e-06, 5.393103e-06, 8.270485e-07, 
    9.919642e-07, 1.575261e-06, 1.249824e-06, 8.45049e-07, 1.880355e-07, 
    9.258957e-07, 6.734335e-06, 2.158974e-05, 1.20755e-05, 2.825924e-06,
  8.058072e-06, 9.066483e-06, 1.663057e-06, 1.73959e-06, 3.263511e-06, 
    5.948525e-06, 4.11133e-06, 3.915728e-06, 3.173073e-06, 4.676894e-06, 
    1.269204e-05, 2.482642e-05, 2.466742e-05, 3.751073e-06, 2.531953e-06,
  1.233086e-05, 4.98117e-06, 2.887424e-06, 4.876227e-06, 7.051634e-06, 
    1.052188e-05, 9.958942e-06, 1.129246e-05, 1.051033e-05, 2.301504e-05, 
    3.443976e-05, 3.04055e-05, 1.020596e-05, 3.812564e-06, 2.357185e-06,
  8.773099e-06, 9.077756e-06, 4.043794e-06, 6.867982e-06, 1.322332e-05, 
    1.555212e-05, 1.774566e-05, 1.708184e-05, 2.881955e-05, 4.523864e-05, 
    3.946312e-05, 1.621033e-05, 6.161652e-06, 4.186171e-06, 3.278574e-06,
  4.338736e-05, 9.652389e-06, 1.676138e-06, 8.531437e-09, 1.733245e-07, 
    6.455188e-07, 8.424939e-07, 7.555849e-07, 1.127039e-06, 2.590594e-06, 
    2.310843e-06, 3.232198e-07, 1.154162e-08, 7.019412e-07, 1.481848e-06,
  4.298279e-05, 1.069826e-05, 5.85825e-07, 7.755375e-07, 1.878989e-06, 
    1.967865e-06, 1.315584e-06, 1.274746e-06, 8.466635e-07, 1.293043e-07, 
    3.335504e-07, 1.582101e-07, 3.355454e-08, 1.978448e-06, 7.507722e-06,
  4.634236e-05, 8.830412e-06, 4.024019e-06, 4.107579e-06, 2.11275e-06, 
    4.575499e-06, 4.29191e-06, 2.768255e-06, 7.950787e-07, 4.90163e-07, 
    2.059679e-06, 4.695813e-07, 6.750079e-07, 2.996056e-06, 3.442677e-05,
  8.351645e-05, 4.738573e-05, 2.139416e-05, 1.517785e-05, 1.449024e-05, 
    2.187422e-06, 9.322008e-06, 2.783185e-06, 1.472708e-06, 7.138196e-07, 
    2.13731e-07, 1.977024e-07, 1.78261e-06, 1.149165e-05, 4.335975e-05,
  8.47785e-05, 5.10553e-05, 3.351742e-05, 2.523362e-05, 1.979493e-05, 
    9.243931e-06, 8.218272e-07, 5.464954e-06, 3.823761e-06, 3.990832e-07, 
    7.124697e-07, 1.237665e-06, 3.923798e-06, 2.252767e-05, 2.805983e-05,
  2.648435e-05, 2.697423e-05, 2.349529e-05, 1.800237e-05, 8.798283e-06, 
    4.924282e-06, 2.023671e-06, 3.659367e-07, 2.20592e-07, 8.963985e-08, 
    9.125463e-08, 1.567766e-06, 1.279836e-05, 1.975784e-05, 7.883454e-06,
  9.255647e-06, 1.009504e-05, 6.629948e-06, 4.409793e-06, 3.879672e-06, 
    3.170102e-06, 2.429147e-06, 1.76054e-07, 9.678103e-07, 3.2867e-06, 
    1.095783e-06, 6.061148e-06, 2.590096e-05, 5.498563e-06, 3.366831e-06,
  8.169873e-06, 6.452491e-06, 2.749292e-07, 2.028877e-06, 3.658773e-06, 
    2.926256e-06, 1.31694e-06, 2.122061e-07, 3.050658e-08, 5.861215e-07, 
    2.090727e-06, 2.099842e-05, 1.587204e-05, 3.760456e-06, 3.22399e-06,
  7.622808e-06, 4.409098e-06, 1.608644e-06, 2.482359e-06, 2.859235e-06, 
    1.388927e-06, 1.132063e-06, 7.64462e-07, 7.85692e-07, 1.73918e-06, 
    6.437728e-06, 2.377122e-05, 1.032071e-05, 5.833641e-06, 4.279034e-06,
  6.951736e-06, 5.874231e-06, 4.137132e-06, 4.551218e-06, 2.884079e-06, 
    6.601549e-07, 2.207081e-06, 4.440734e-07, 3.854245e-07, 3.566779e-06, 
    1.779001e-05, 1.83241e-05, 1.374272e-05, 1.168039e-05, 7.061196e-06,
  3.121014e-05, 1.350647e-06, 3.937793e-06, 1.216645e-05, 1.187108e-05, 
    3.420775e-06, 1.574205e-06, 7.805852e-08, 1.559472e-07, 5.704311e-07, 
    1.416022e-06, 8.733524e-07, 9.574451e-07, 2.052045e-06, 3.652099e-06,
  4.340641e-06, 6.136947e-06, 1.158773e-05, 2.311699e-05, 2.78405e-05, 
    7.72867e-06, 1.714813e-06, 4.937287e-07, 2.789099e-07, 9.806179e-07, 
    1.320379e-06, 1.301117e-06, 1.809396e-06, 4.929678e-06, 5.833524e-06,
  1.783823e-05, 2.767351e-05, 3.166177e-05, 3.92641e-05, 2.20303e-05, 
    1.965396e-05, 2.202906e-06, 1.211239e-06, 1.379448e-06, 1.342161e-06, 
    1.1482e-06, 1.157802e-06, 2.912061e-06, 5.942347e-06, 8.838418e-06,
  4.902093e-05, 5.37404e-05, 5.239122e-05, 4.392569e-05, 3.781723e-05, 
    2.636676e-06, 1.191288e-05, 4.043151e-06, 1.522286e-06, 5.654209e-07, 
    8.042263e-08, 2.098472e-06, 4.673119e-06, 4.011887e-06, 1.105087e-05,
  7.186081e-05, 6.428784e-05, 7.044246e-05, 4.223268e-05, 4.616623e-05, 
    7.446478e-06, 6.481993e-07, 1.805258e-06, 2.426912e-06, 1.052925e-07, 
    1.129096e-07, 1.825519e-06, 6.742845e-06, 1.434762e-05, 1.937298e-05,
  9.334298e-05, 6.406202e-05, 7.052271e-05, 3.888652e-05, 2.334073e-05, 
    5.939933e-06, 8.320415e-07, 1.995717e-07, 8.152585e-08, 9.206747e-08, 
    2.841307e-06, 3.679169e-06, 1.161034e-05, 1.874448e-05, 1.550687e-05,
  9.313328e-05, 7.941599e-05, 7.397558e-05, 3.465098e-05, 1.351281e-05, 
    2.145395e-06, 3.989206e-07, 3.212188e-07, 2.040576e-06, 2.311828e-06, 
    4.182796e-06, 8.732144e-06, 1.255106e-05, 1.580167e-05, 1.188699e-05,
  8.111116e-05, 8.233149e-05, 5.38003e-05, 2.573213e-05, 8.614518e-06, 
    1.808565e-06, 2.907703e-07, 2.70523e-07, 2.1296e-07, 2.426401e-07, 
    3.19413e-06, 9.716211e-06, 9.44778e-06, 1.201859e-05, 1.390734e-05,
  6.593615e-05, 4.521498e-05, 3.348492e-05, 2.127185e-05, 9.145507e-06, 
    3.429547e-06, 4.078375e-07, 1.956933e-08, 2.82637e-07, 1.23111e-06, 
    2.569246e-06, 7.107279e-06, 2.786697e-06, 4.643927e-06, 1.445775e-05,
  4.417586e-05, 2.812409e-05, 2.459428e-05, 1.635117e-05, 8.949819e-06, 
    4.047391e-06, 1.326214e-06, 4.656348e-09, 3.098256e-08, 8.091889e-07, 
    6.275515e-06, 6.906662e-06, 3.496206e-06, 9.555836e-06, 2.71675e-05,
  0.0002113222, 0.0001145875, 3.003439e-05, 2.609931e-05, 8.583514e-05, 
    7.893132e-05, 4.049469e-05, 3.39929e-05, 1.94006e-05, 6.343992e-06, 
    1.223202e-06, 1.464819e-07, 4.5976e-07, 7.91421e-07, 8.123135e-07,
  0.0002139223, 8.386411e-05, 3.052607e-05, 4.303544e-05, 7.994242e-05, 
    6.182535e-05, 4.798458e-05, 4.282839e-05, 2.2181e-05, 4.45474e-06, 
    1.399935e-06, 6.640398e-07, 7.22814e-07, 7.913197e-07, 7.848607e-07,
  0.0001130912, 7.127326e-05, 4.000849e-05, 5.054593e-05, 4.131992e-05, 
    7.82345e-05, 5.635581e-05, 5.163649e-05, 2.317318e-05, 3.403051e-06, 
    1.189264e-06, 7.310713e-07, 4.825101e-07, 7.829873e-07, 2.549943e-06,
  0.0001049201, 6.664647e-05, 3.136679e-05, 3.709766e-05, 3.360808e-05, 
    3.427682e-06, 6.743347e-05, 3.325725e-05, 1.039933e-05, 1.453668e-06, 
    7.356713e-07, 8.029025e-07, 6.256373e-07, 5.080493e-07, 4.714198e-06,
  8.645145e-05, 4.712394e-05, 1.482407e-05, 2.189291e-05, 3.809252e-05, 
    2.115236e-05, 9.2825e-07, 2.444664e-06, 5.641452e-06, 1.465608e-06, 
    7.282003e-07, 3.627026e-07, 4.054804e-06, 5.751867e-06, 1.116721e-05,
  3.843896e-05, 1.17567e-05, 4.442732e-06, 1.041467e-05, 1.555528e-05, 
    1.06603e-05, 1.220463e-06, 8.113168e-08, 9.215588e-08, 4.230787e-07, 
    1.26016e-06, 9.21188e-07, 9.525153e-06, 1.22102e-05, 1.266241e-05,
  2.106689e-05, 9.944149e-06, 1.233575e-05, 9.504382e-06, 5.826416e-06, 
    2.337511e-06, 9.389067e-07, 1.061066e-06, 1.127842e-06, 2.803858e-06, 
    1.742747e-06, 7.158165e-06, 1.2435e-05, 6.790042e-06, 5.069112e-06,
  2.365056e-05, 2.421536e-05, 2.213557e-05, 3.632741e-06, 2.839994e-06, 
    1.038214e-06, 5.763507e-07, 7.631073e-07, 1.435176e-06, 2.148287e-06, 
    1.007068e-05, 5.503626e-06, 7.778077e-06, 9.640227e-06, 1.15372e-05,
  4.180657e-05, 4.460938e-05, 1.430006e-05, 3.733556e-06, 3.013039e-06, 
    2.487383e-06, 2.69529e-06, 3.631697e-06, 2.964999e-06, 6.265465e-06, 
    6.079433e-06, 4.846755e-06, 6.642627e-06, 1.225938e-05, 1.898379e-05,
  6.938841e-05, 2.688162e-05, 4.730759e-06, 3.369776e-06, 2.956067e-06, 
    2.497551e-06, 3.52892e-06, 5.131539e-06, 5.528585e-06, 4.583209e-06, 
    3.423335e-06, 3.818571e-06, 6.942985e-06, 1.242567e-05, 1.337194e-05,
  1.31786e-06, 8.630015e-07, 2.020291e-06, 0.0001004908, 8.379132e-05, 
    8.287871e-06, 7.602714e-06, 3.116684e-05, 0.000115177, 0.0001267818, 
    1.9862e-05, 2.965577e-07, 1.940224e-07, 3.494416e-06, 5.768429e-06,
  5.448451e-05, 1.529499e-05, 2.313657e-06, 1.924741e-05, 1.315856e-06, 
    1.151377e-06, 6.446797e-06, 2.858551e-05, 8.983369e-05, 0.0001562026, 
    4.696885e-05, 4.680359e-06, 1.017868e-07, 1.267496e-06, 3.110017e-06,
  4.450688e-05, 9.872416e-06, 2.770097e-06, 2.530272e-06, 7.4485e-07, 
    2.30474e-06, 2.770083e-06, 3.421729e-05, 0.0001035505, 0.0001715561, 
    0.0001093117, 1.753107e-05, 3.900607e-06, 2.032632e-07, 1.7829e-06,
  1.157105e-05, 3.771173e-06, 3.273548e-06, 2.293609e-06, 1.28769e-06, 
    6.985413e-07, 2.741573e-05, 5.588908e-05, 9.963413e-05, 0.0001135662, 
    0.0001144716, 4.515129e-05, 9.150951e-06, 4.276225e-07, 1.332105e-06,
  1.09915e-05, 6.554352e-06, 7.350328e-06, 6.874904e-06, 8.742698e-06, 
    1.86186e-05, 1.163365e-05, 4.975027e-05, 8.76562e-05, 4.47849e-05, 
    7.636067e-05, 7.341934e-05, 2.384125e-05, 7.476158e-06, 2.747016e-06,
  1.536372e-05, 1.515523e-05, 1.154854e-05, 1.035507e-05, 9.283849e-06, 
    2.112604e-05, 2.424164e-05, 7.396187e-06, 1.457153e-05, 6.474983e-05, 
    4.182907e-05, 6.928142e-05, 6.403251e-05, 3.095257e-05, 8.055739e-06,
  8.802214e-06, 1.269607e-05, 1.643112e-05, 1.908315e-05, 1.878765e-05, 
    2.966009e-05, 6.071846e-05, 0.0001104034, 0.0001051587, 6.082495e-05, 
    4.421376e-05, 4.507462e-05, 3.987291e-05, 1.911724e-05, 6.644385e-06,
  5.939214e-06, 1.034955e-05, 1.771901e-05, 2.393526e-05, 2.824839e-05, 
    2.88267e-05, 2.25266e-05, 2.286982e-05, 2.188398e-05, 1.654145e-05, 
    1.16318e-05, 9.204033e-06, 7.371837e-06, 5.887997e-06, 3.694526e-06,
  6.744292e-06, 6.976892e-06, 7.919195e-06, 8.654553e-06, 6.259821e-06, 
    3.943785e-06, 3.593305e-06, 4.072404e-06, 3.614938e-06, 3.328968e-06, 
    2.433589e-06, 3.144558e-06, 4.543335e-06, 5.836301e-06, 3.825598e-06,
  2.114916e-06, 3.572456e-06, 4.460374e-06, 4.089978e-06, 4.019782e-06, 
    3.94021e-06, 3.45161e-06, 3.362335e-06, 2.661293e-06, 3.103098e-06, 
    3.780812e-06, 7.474986e-06, 5.023797e-06, 4.682877e-06, 5.787593e-06,
  8.970062e-06, 8.024747e-06, 6.715713e-06, 7.846768e-05, 0.0001478834, 
    6.235861e-05, 1.07843e-05, 2.765415e-06, 4.353412e-06, 1.82245e-05, 
    2.81722e-06, 1.308699e-06, 3.119668e-07, 2.014489e-06, 1.718482e-06,
  5.667334e-06, 5.697173e-06, 2.658954e-05, 0.00014446, 0.0001447652, 
    6.939075e-05, 3.481226e-05, 7.932595e-06, 7.956173e-06, 1.626835e-05, 
    5.959112e-06, 6.050012e-07, 3.932473e-07, 3.243607e-06, 4.291542e-06,
  7.611137e-06, 2.849901e-05, 9.448864e-05, 0.0001526904, 0.0001175295, 
    9.114653e-05, 3.647436e-05, 2.492966e-05, 2.039342e-05, 2.365303e-05, 
    6.848669e-06, 2.162995e-06, 3.412455e-07, 1.926227e-06, 3.335604e-06,
  8.050841e-06, 1.663684e-05, 5.118054e-05, 0.0001393521, 0.0001250141, 
    6.419563e-05, 6.187573e-05, 2.421743e-05, 3.000011e-05, 4.341259e-05, 
    1.101433e-05, 1.996903e-06, 1.104118e-06, 5.174729e-06, 3.341695e-06,
  5.085238e-06, 5.751572e-06, 2.042528e-05, 8.580886e-05, 8.798151e-05, 
    6.389927e-05, 9.170407e-06, 1.182843e-05, 5.902087e-05, 5.144083e-05, 
    3.161605e-05, 1.084999e-05, 3.776793e-06, 5.607359e-06, 4.167421e-06,
  7.996578e-06, 9.408252e-06, 1.401796e-05, 2.966215e-05, 4.563672e-05, 
    3.197346e-05, 9.135611e-06, 2.694302e-06, 2.035619e-06, 3.710618e-05, 
    5.930583e-05, 4.184111e-05, 2.663478e-05, 7.568274e-06, 6.530605e-06,
  8.366725e-06, 1.13026e-05, 1.281126e-05, 1.943487e-05, 3.908251e-05, 
    3.03168e-05, 1.210928e-05, 6.926763e-06, 1.42544e-05, 4.369254e-05, 
    6.418446e-05, 7.585368e-05, 5.67967e-05, 3.594166e-05, 9.981125e-06,
  8.455397e-06, 8.210334e-06, 1.362451e-05, 1.895524e-05, 3.071647e-05, 
    4.377947e-05, 2.398986e-05, 1.352184e-05, 1.910232e-05, 5.167384e-05, 
    6.519025e-05, 6.839605e-05, 9.221478e-05, 7.937625e-05, 4.971685e-05,
  6.072714e-06, 4.329478e-06, 7.604378e-06, 8.232397e-06, 1.304136e-05, 
    2.24878e-05, 2.732184e-05, 2.349389e-05, 2.164824e-05, 4.313601e-05, 
    4.641791e-05, 5.001905e-05, 6.706622e-05, 6.504409e-05, 5.856044e-05,
  2.866576e-06, 2.58372e-06, 2.793606e-06, 2.827046e-06, 3.303822e-06, 
    5.099478e-06, 8.175732e-06, 1.087401e-05, 1.112991e-05, 1.797708e-05, 
    2.167056e-05, 2.261678e-05, 2.714252e-05, 2.724957e-05, 2.862432e-05,
  8.290558e-06, 7.822549e-06, 7.262534e-06, 9.317696e-06, 6.432711e-06, 
    2.236152e-06, 4.834541e-07, 6.045839e-08, 1.269181e-08, 5.517218e-07, 
    1.523903e-06, 1.716643e-05, 5.589139e-06, 3.388943e-06, 7.732552e-07,
  1.01655e-05, 9.990745e-06, 1.078138e-05, 1.159371e-05, 8.405423e-06, 
    9.35401e-06, 8.721107e-07, 6.959448e-08, 2.49697e-08, 1.032198e-06, 
    8.459922e-07, 1.547759e-05, 5.492011e-06, 4.218291e-06, 1.077756e-06,
  8.598439e-06, 1.104004e-05, 2.572215e-05, 2.201596e-05, 1.486453e-05, 
    1.933037e-05, 3.948659e-06, 1.079047e-06, 4.39583e-07, 6.978651e-07, 
    2.637287e-07, 9.950127e-06, 3.753661e-06, 1.294217e-06, 8.661851e-08,
  9.958285e-06, 1.150108e-05, 3.725536e-05, 4.787864e-05, 3.274052e-05, 
    8.021841e-06, 1.715147e-05, 5.511195e-06, 2.010594e-06, 3.019829e-07, 
    5.265642e-07, 9.708701e-06, 3.348729e-06, 1.860299e-06, 2.013154e-07,
  8.84516e-06, 1.053314e-05, 3.724795e-05, 6.75449e-05, 5.837076e-05, 
    2.129399e-05, 2.13129e-06, 2.323383e-05, 1.222441e-05, 1.155495e-07, 
    5.880081e-07, 6.712001e-06, 5.131983e-06, 2.539621e-06, 1.221226e-06,
  1.080438e-05, 1.613595e-05, 2.919837e-05, 4.394999e-05, 4.269119e-05, 
    2.158594e-05, 2.807358e-06, 2.212151e-07, 5.185376e-07, 1.227409e-07, 
    2.920928e-07, 4.38641e-06, 4.144098e-06, 3.884815e-06, 2.497266e-06,
  1.368521e-05, 1.951996e-05, 3.343062e-05, 3.945988e-05, 3.734825e-05, 
    2.381297e-05, 3.41346e-06, 6.309243e-07, 6.228528e-07, 1.720766e-07, 
    9.258977e-07, 5.127358e-06, 4.784124e-06, 6.754755e-06, 3.977434e-06,
  1.492074e-05, 2.179316e-05, 4.268641e-05, 5.011417e-05, 5.773428e-05, 
    4.288991e-05, 7.256131e-06, 1.437733e-06, 7.093695e-07, 9.144026e-07, 
    2.006112e-06, 6.137424e-06, 6.343017e-06, 8.595436e-06, 8.472906e-06,
  1.483766e-05, 2.714774e-05, 4.799396e-05, 6.832034e-05, 7.963824e-05, 
    6.203664e-05, 2.609861e-05, 8.16008e-06, 5.035623e-06, 1.470606e-05, 
    2.020996e-05, 6.487334e-06, 7.191812e-06, 9.797674e-06, 1.212546e-05,
  1.192534e-05, 2.530381e-05, 4.822528e-05, 6.268195e-05, 6.778711e-05, 
    6.354198e-05, 4.083433e-05, 1.911271e-05, 1.73753e-05, 3.213361e-05, 
    3.173972e-05, 1.144127e-05, 1.044275e-05, 1.180327e-05, 1.328066e-05,
  3.472713e-07, 1.159877e-06, 7.81355e-07, 3.761231e-06, 3.316383e-06, 
    1.956326e-06, 2.551845e-06, 3.468517e-06, 3.896267e-06, 1.327e-06, 
    3.07475e-07, 2.83625e-06, 2.158117e-05, 4.949829e-05, 6.396668e-05,
  1.496799e-07, 3.333101e-07, 2.359845e-06, 4.618273e-06, 7.471235e-06, 
    3.022918e-06, 1.816052e-06, 2.600732e-06, 2.449357e-06, 1.589368e-06, 
    3.331382e-07, 7.35161e-06, 3.358743e-05, 7.301837e-05, 7.617828e-05,
  2.532328e-06, 1.65361e-06, 3.787832e-06, 4.096613e-06, 6.146458e-06, 
    1.623433e-05, 2.04173e-06, 1.503026e-06, 1.439246e-06, 9.929064e-07, 
    1.176186e-06, 2.491709e-05, 5.416349e-05, 7.921879e-05, 8.091572e-05,
  2.783071e-06, 2.986276e-06, 4.690554e-06, 6.321613e-06, 9.783455e-06, 
    1.279147e-05, 1.327661e-05, 3.257519e-06, 2.431606e-06, 3.695016e-07, 
    4.760427e-06, 4.736019e-05, 6.784906e-05, 9.270412e-05, 6.997376e-05,
  4.771518e-06, 1.007536e-05, 6.350603e-06, 4.786916e-06, 6.492722e-06, 
    1.59086e-05, 7.585353e-06, 1.227576e-05, 8.496408e-06, 7.447668e-07, 
    1.772965e-05, 6.807232e-05, 7.138098e-05, 5.640325e-05, 2.577782e-05,
  1.684173e-05, 1.731847e-05, 1.302306e-05, 9.070111e-06, 6.129214e-06, 
    9.442996e-06, 7.915005e-06, 9.337988e-07, 2.93471e-07, 1.605929e-07, 
    3.221192e-05, 7.436339e-05, 5.422825e-05, 1.798088e-05, 2.445913e-06,
  1.928926e-05, 2.372843e-05, 1.903972e-05, 1.089759e-05, 5.731958e-06, 
    7.846432e-06, 6.294898e-06, 2.559454e-06, 2.180143e-06, 1.575763e-06, 
    5.225163e-05, 6.141272e-05, 2.08588e-05, 3.868197e-06, 2.207006e-06,
  1.834382e-05, 2.417997e-05, 1.962677e-05, 8.190964e-06, 7.725798e-06, 
    1.095513e-05, 5.936305e-06, 1.41802e-06, 8.222893e-07, 1.935909e-05, 
    5.904615e-05, 2.738099e-05, 5.294511e-06, 3.655412e-06, 4.608925e-06,
  1.537749e-05, 2.355642e-05, 2.623865e-05, 1.765342e-05, 1.639454e-05, 
    1.446516e-05, 6.768009e-06, 6.319514e-07, 5.191992e-06, 3.104529e-05, 
    4.58089e-05, 7.71481e-06, 4.447608e-06, 4.602469e-06, 7.274705e-06,
  1.090825e-05, 1.952959e-05, 3.000567e-05, 2.809484e-05, 2.320253e-05, 
    1.299441e-05, 3.670598e-06, 1.135965e-06, 4.962305e-06, 1.73732e-05, 
    2.369461e-05, 5.823147e-06, 4.98175e-06, 7.493432e-06, 8.751144e-06,
  3.908692e-06, 3.778584e-06, 3.958631e-06, 3.051723e-06, 2.360186e-06, 
    2.089355e-06, 1.455399e-06, 1.633656e-06, 2.40714e-06, 4.932377e-06, 
    4.24995e-06, 3.187641e-06, 3.700365e-06, 2.177717e-06, 4.574229e-06,
  7.589335e-07, 4.138884e-07, 5.077612e-07, 1.206531e-06, 2.266883e-06, 
    1.882712e-06, 1.339251e-06, 2.363679e-06, 3.596122e-06, 3.646161e-06, 
    1.989688e-06, 1.228086e-06, 1.549484e-06, 5.119702e-06, 4.192392e-06,
  1.261664e-07, 3.274246e-08, 8.063184e-07, 1.968847e-06, 2.956954e-06, 
    5.864394e-06, 5.03765e-07, 1.06446e-06, 1.500865e-06, 1.029421e-06, 
    7.993705e-07, 6.635937e-07, 3.256222e-06, 2.184649e-06, 6.092805e-06,
  1.073137e-07, 6.254319e-07, 2.154371e-06, 3.035072e-06, 4.741313e-06, 
    4.64601e-06, 1.1117e-05, 9.096759e-07, 3.66387e-07, 2.530349e-07, 
    3.348684e-07, 2.512429e-06, 1.304443e-05, 8.594911e-06, 1.660594e-05,
  7.109643e-07, 4.041649e-06, 7.534967e-06, 8.916758e-06, 1.084274e-05, 
    1.966459e-05, 1.197095e-05, 3.506378e-05, 5.638339e-06, 7.616785e-07, 
    7.38054e-07, 1.385304e-05, 3.773831e-05, 2.072387e-05, 3.560722e-05,
  4.081059e-06, 1.130967e-05, 1.370579e-05, 1.212152e-05, 8.642119e-06, 
    7.658015e-06, 1.041002e-05, 1.787697e-06, 9.161816e-07, 8.571641e-07, 
    2.340752e-06, 4.197969e-05, 5.470482e-05, 2.622007e-05, 1.994801e-05,
  7.825077e-06, 1.077143e-05, 9.777444e-06, 1.102959e-05, 8.610867e-06, 
    5.45971e-06, 5.50994e-06, 6.194572e-06, 4.841583e-06, 2.014178e-06, 
    2.244983e-05, 7.103716e-05, 4.855235e-05, 1.397276e-05, 1.259776e-05,
  1.068892e-05, 1.109107e-05, 4.726063e-06, 4.18728e-06, 4.942785e-06, 
    4.661038e-06, 3.319984e-06, 4.896723e-06, 3.45338e-06, 8.315069e-06, 
    7.371239e-05, 6.673652e-05, 2.164971e-05, 1.009179e-05, 9.085303e-06,
  1.156579e-05, 5.550651e-06, 4.156227e-06, 3.661475e-06, 4.206776e-06, 
    3.759696e-06, 4.571931e-06, 4.601665e-06, 1.055532e-05, 5.209296e-05, 
    7.992285e-05, 3.466556e-05, 8.042593e-06, 8.160477e-06, 3.079128e-06,
  6.000434e-06, 7.445579e-06, 5.125473e-06, 3.235878e-06, 3.14443e-06, 
    4.389287e-06, 5.970431e-06, 1.126657e-05, 4.585152e-05, 9.094828e-05, 
    4.721541e-05, 9.79133e-06, 7.553771e-06, 4.570599e-06, 3.789345e-07,
  0.0001081594, 7.650707e-05, 5.391962e-05, 3.164092e-05, 2.149284e-05, 
    6.002922e-06, 4.05526e-06, 2.975958e-06, 4.269033e-06, 1.005071e-06, 
    1.429176e-06, 1.793098e-06, 1.431754e-06, 6.103737e-07, 4.350245e-06,
  0.0001555561, 8.088604e-05, 5.561955e-05, 3.776797e-05, 1.737194e-05, 
    4.956497e-06, 1.248297e-06, 2.885675e-06, 3.582628e-06, 1.042864e-06, 
    8.442415e-07, 4.655374e-07, 9.516254e-07, 4.074163e-06, 2.220686e-05,
  0.0002435826, 9.811465e-05, 2.877013e-05, 2.750908e-05, 1.805144e-05, 
    1.992673e-05, 2.866127e-06, 8.391329e-07, 1.072269e-06, 6.516879e-07, 
    9.930444e-07, 3.556431e-08, 2.376008e-06, 5.47039e-06, 6.874976e-05,
  0.0002311492, 0.0001540563, 3.964918e-05, 1.127577e-05, 1.113391e-05, 
    9.380189e-07, 2.20334e-05, 4.29776e-07, 8.620593e-08, 1.750201e-08, 
    2.677238e-09, 4.832201e-09, 3.599806e-06, 6.752647e-06, 9.735669e-05,
  6.465123e-05, 7.827678e-05, 4.148381e-05, 1.001558e-05, 6.528474e-06, 
    7.50089e-06, 2.503431e-06, 1.42165e-05, 2.806888e-06, 1.977354e-08, 
    2.827901e-08, 1.112465e-07, 1.939793e-06, 6.793946e-06, 6.325773e-05,
  6.960008e-07, 4.177937e-06, 5.093906e-06, 3.734901e-06, 3.068282e-06, 
    4.224704e-06, 6.152459e-06, 1.965678e-06, 2.381435e-07, 1.023895e-07, 
    1.316101e-07, 3.27988e-06, 3.089769e-06, 6.488798e-06, 1.630041e-05,
  2.429915e-06, 3.74408e-06, 4.423493e-06, 4.482871e-06, 4.626642e-06, 
    3.894159e-06, 5.145163e-06, 8.660514e-06, 3.876296e-06, 5.143983e-07, 
    2.524543e-07, 9.290566e-07, 3.325821e-06, 8.335894e-06, 1.01929e-05,
  1.013725e-06, 5.015831e-06, 3.463879e-06, 4.627167e-06, 4.277888e-06, 
    4.656695e-06, 4.634829e-06, 4.466349e-06, 3.39724e-06, 6.420412e-07, 
    1.622815e-06, 1.530081e-06, 5.97588e-06, 8.89488e-06, 7.558565e-06,
  2.964614e-06, 8.805739e-06, 1.111722e-05, 1.147567e-05, 1.211668e-05, 
    9.442761e-06, 6.219278e-06, 4.280007e-06, 3.058806e-06, 1.520031e-06, 
    7.998305e-07, 2.867912e-06, 5.535902e-06, 8.395293e-06, 5.632386e-06,
  5.840627e-06, 2.401578e-05, 2.638901e-05, 2.313442e-05, 2.023618e-05, 
    1.58146e-05, 7.28923e-06, 3.980022e-06, 4.866596e-06, 1.761644e-06, 
    8.792509e-07, 3.933916e-06, 5.855939e-06, 1.014388e-05, 2.510395e-06,
  3.340001e-05, 3.226859e-05, 4.847837e-05, 0.00014287, 0.0001312251, 
    9.749053e-05, 7.897235e-05, 5.728327e-05, 2.17409e-05, 6.309074e-06, 
    4.348211e-07, 1.882424e-08, 1.43743e-07, 3.303874e-06, 6.174172e-06,
  7.606853e-05, 3.338964e-05, 5.494629e-05, 9.89523e-05, 8.434065e-05, 
    8.309961e-05, 5.378892e-05, 2.225498e-05, 7.599494e-06, 3.779239e-06, 
    9.285998e-08, 8.235298e-07, 1.773178e-06, 5.973086e-06, 6.379086e-06,
  0.0001437772, 6.610037e-05, 6.981823e-05, 8.38466e-05, 3.726858e-05, 
    5.589697e-05, 1.886732e-05, 7.873966e-06, 4.408619e-06, 1.008208e-06, 
    1.030895e-06, 1.794554e-06, 1.802053e-06, 5.210684e-06, 2.356081e-06,
  0.0001944586, 0.0001593125, 0.0001103443, 7.627908e-05, 4.724378e-05, 
    6.314529e-06, 3.344057e-05, 1.144985e-05, 2.140102e-06, 9.365223e-07, 
    1.850003e-06, 2.097742e-06, 2.850266e-06, 6.037331e-06, 4.979602e-06,
  0.0001435317, 0.0002556331, 0.0001942703, 8.980372e-05, 5.171655e-05, 
    2.505156e-05, 2.743892e-06, 1.129633e-05, 6.23597e-06, 2.396444e-06, 
    1.544003e-06, 3.028772e-06, 4.885042e-06, 5.907547e-06, 6.78019e-06,
  2.51026e-05, 0.0002254853, 0.0002379092, 9.650859e-05, 4.208794e-05, 
    3.493145e-05, 2.309319e-05, 4.233603e-06, 8.482265e-07, 1.201391e-06, 
    1.51049e-06, 2.008898e-06, 4.935785e-06, 7.132558e-06, 6.488201e-06,
  4.1317e-06, 0.0001188884, 0.000234859, 0.0001062806, 2.565285e-05, 
    1.485951e-05, 2.969966e-05, 1.010451e-05, 2.772539e-06, 1.365584e-06, 
    1.68233e-06, 4.107156e-06, 6.214811e-06, 9.315527e-06, 7.828132e-06,
  4.370704e-07, 3.216999e-05, 0.0001939245, 0.0001397285, 2.226021e-05, 
    9.247733e-06, 4.799681e-06, 1.239574e-06, 9.306313e-07, 7.889881e-07, 
    1.99165e-06, 3.009506e-06, 7.531637e-06, 8.776196e-06, 7.215312e-06,
  2.392124e-06, 8.093954e-06, 0.0001213035, 0.0001409431, 3.239936e-05, 
    8.765348e-06, 3.784539e-06, 1.663552e-06, 1.724382e-06, 1.580014e-06, 
    5.648639e-07, 7.60144e-06, 9.532007e-06, 9.076497e-06, 5.391629e-06,
  3.977326e-06, 3.68691e-06, 4.252683e-05, 9.418633e-05, 5.057058e-05, 
    1.609822e-05, 5.669522e-06, 4.571248e-06, 3.663108e-06, 3.283747e-06, 
    8.955937e-07, 8.953618e-06, 9.267427e-06, 8.30625e-06, 6.133222e-06,
  2.709407e-08, 5.707263e-06, 1.996823e-05, 4.304051e-05, 1.581247e-05, 
    6.148317e-06, 1.792555e-05, 7.524552e-05, 0.0001175657, 7.458196e-05, 
    3.626676e-05, 9.09651e-06, 2.668482e-07, 4.194442e-07, 9.577374e-07,
  2.672546e-08, 7.388853e-06, 2.158389e-05, 3.94638e-05, 1.909203e-05, 
    2.608634e-05, 5.631389e-05, 9.750679e-05, 9.739656e-05, 4.461916e-05, 
    4.473131e-06, 2.568505e-07, 3.361181e-07, 2.610563e-06, 2.749923e-06,
  4.456937e-06, 6.488205e-06, 2.101943e-05, 3.895192e-05, 1.905128e-05, 
    6.253172e-05, 5.472432e-05, 8.132857e-05, 5.836913e-05, 4.611938e-06, 
    2.665099e-06, 2.719208e-06, 2.279485e-06, 1.832857e-06, 3.182735e-06,
  3.041193e-05, 6.161588e-06, 2.09732e-05, 1.300168e-05, 1.98526e-05, 
    3.394877e-06, 6.910937e-05, 1.647119e-05, 7.409469e-06, 5.596525e-06, 
    4.891426e-06, 3.260811e-06, 4.157535e-06, 3.975068e-06, 2.278987e-06,
  2.726382e-05, 2.711719e-06, 3.930186e-05, 4.549335e-06, 7.098208e-06, 
    9.903423e-06, 5.286007e-07, 1.0193e-06, 8.339989e-06, 4.339629e-06, 
    6.064787e-06, 4.680501e-06, 4.380373e-06, 2.080521e-06, 1.70863e-06,
  9.539825e-06, 2.176303e-06, 4.548305e-05, 7.467915e-06, 1.147061e-06, 
    4.782435e-06, 1.745004e-06, 1.36864e-06, 3.439388e-07, 4.712746e-06, 
    4.601749e-06, 4.439773e-06, 4.071372e-06, 3.316056e-06, 3.312366e-06,
  3.410795e-06, 1.854827e-06, 5.005777e-05, 1.551557e-05, 2.653333e-06, 
    4.656818e-06, 8.030849e-07, 2.609175e-06, 3.559623e-06, 3.777202e-06, 
    3.559202e-06, 3.556532e-06, 3.686333e-06, 3.284482e-06, 4.713856e-06,
  2.884949e-06, 1.641682e-06, 6.546518e-05, 3.10784e-05, 1.326998e-05, 
    1.060352e-05, 1.860985e-06, 1.751783e-06, 2.725848e-06, 3.587703e-06, 
    2.929371e-06, 4.772606e-06, 5.790781e-06, 5.438678e-06, 5.993681e-06,
  2.377726e-06, 1.704202e-06, 7.466268e-05, 7.051629e-05, 3.358272e-05, 
    2.185132e-05, 4.951018e-06, 3.502187e-06, 3.376852e-06, 4.797446e-06, 
    3.834832e-06, 4.255941e-06, 6.173607e-06, 5.98583e-06, 5.320979e-06,
  2.31764e-06, 3.414581e-06, 7.942537e-05, 0.0001106023, 5.585309e-05, 
    3.464794e-05, 1.268793e-05, 3.516681e-06, 2.928283e-06, 5.200527e-06, 
    7.004304e-06, 5.638472e-06, 5.620592e-06, 6.285713e-06, 6.598602e-06,
  6.173373e-06, 4.783639e-06, 3.440523e-05, 3.610761e-05, 1.320031e-05, 
    6.059841e-06, 6.831408e-06, 9.384058e-06, 5.944439e-06, 3.112352e-06, 
    2.995144e-06, 2.082507e-06, 1.976699e-06, 2.497237e-06, 1.5054e-06,
  2.470741e-05, 2.725163e-05, 5.102103e-05, 4.495131e-05, 1.57972e-05, 
    7.915215e-06, 6.724986e-06, 5.322236e-06, 1.353809e-06, 2.706013e-06, 
    3.294711e-06, 1.604045e-06, 6.37682e-07, 1.039368e-06, 2.255576e-06,
  0.0001047949, 6.132588e-05, 5.034842e-05, 4.112595e-05, 1.694267e-05, 
    2.837889e-05, 1.192108e-05, 5.38664e-06, 4.062617e-06, 2.505079e-06, 
    1.173095e-06, 5.937964e-07, 1.057231e-06, 1.087775e-06, 1.395005e-06,
  0.0001311233, 7.074752e-05, 4.866217e-05, 3.515026e-05, 3.117603e-05, 
    7.168722e-06, 3.41303e-05, 9.676643e-06, 6.962214e-06, 4.4345e-06, 
    2.881885e-06, 2.145651e-06, 1.101977e-06, 1.221791e-06, 2.599689e-06,
  0.0001101728, 8.204015e-05, 6.319572e-05, 4.154263e-05, 3.827765e-05, 
    3.558964e-05, 8.708283e-06, 6.788286e-06, 6.060187e-06, 3.847761e-06, 
    5.937317e-06, 2.549769e-06, 3.863887e-06, 4.980689e-06, 3.949971e-06,
  8.439962e-05, 7.352493e-05, 6.005052e-05, 4.678681e-05, 4.276112e-05, 
    4.661302e-05, 2.934239e-05, 8.302558e-07, 6.631209e-07, 6.550931e-06, 
    4.548865e-06, 4.344083e-06, 3.993498e-06, 4.181179e-06, 5.459651e-06,
  8.239935e-05, 7.791026e-05, 7.254394e-05, 7.205083e-05, 6.876957e-05, 
    5.914621e-05, 4.182504e-05, 1.136193e-05, 4.679386e-06, 7.162048e-06, 
    4.309424e-06, 4.535932e-06, 3.049297e-06, 2.809288e-06, 5.099508e-06,
  0.0001013861, 0.0001090557, 0.0001181682, 0.0001203567, 0.0001038697, 
    7.91382e-05, 3.660339e-05, 9.959997e-06, 6.632161e-06, 7.267229e-06, 
    4.015164e-06, 4.193443e-06, 4.174119e-06, 5.92457e-06, 5.085889e-06,
  9.183311e-05, 0.0001057912, 0.0001512452, 0.0001770577, 0.0001404901, 
    7.414663e-05, 2.701628e-05, 7.992846e-06, 9.044874e-06, 7.279265e-06, 
    4.295306e-06, 3.785088e-06, 5.678671e-06, 5.542453e-06, 4.072953e-06,
  7.738436e-05, 9.58516e-05, 0.0001657027, 0.000198335, 0.0001450121, 
    6.062534e-05, 1.773434e-05, 8.040258e-06, 1.004507e-05, 5.919314e-06, 
    5.182443e-06, 5.548916e-06, 6.262648e-06, 6.344531e-06, 7.938707e-06,
  8.106342e-05, 5.043065e-05, 4.762126e-05, 4.889701e-05, 2.846042e-05, 
    1.698882e-05, 1.079923e-05, 1.159384e-05, 1.398122e-05, 1.090507e-05, 
    6.347475e-06, 5.484216e-06, 7.784164e-06, 8.300276e-06, 5.333437e-06,
  0.0001323275, 0.0001068078, 9.989813e-05, 7.896017e-05, 4.07296e-05, 
    1.110437e-05, 1.371413e-05, 1.137611e-05, 1.32332e-05, 2.079007e-05, 
    1.724176e-05, 7.743224e-06, 5.440074e-06, 2.367651e-06, 3.583237e-06,
  0.0001069144, 7.972173e-05, 5.628862e-05, 3.11604e-05, 1.273031e-05, 
    1.500079e-05, 1.111029e-05, 3.458604e-05, 2.356902e-05, 2.380088e-05, 
    2.022942e-05, 1.410325e-05, 5.348613e-06, 3.59162e-06, 4.022064e-06,
  4.724999e-05, 1.422996e-05, 5.81683e-06, 4.001076e-06, 4.894605e-06, 
    7.297007e-06, 3.035312e-05, 3.862141e-05, 3.204144e-05, 3.261615e-05, 
    3.069348e-05, 2.195755e-05, 1.069742e-05, 5.234617e-06, 3.602605e-06,
  2.037526e-06, 1.656096e-06, 1.39468e-06, 2.123004e-06, 3.508791e-06, 
    1.112393e-05, 1.948985e-05, 4.791009e-05, 2.986778e-05, 3.957266e-05, 
    4.489045e-05, 2.813027e-05, 1.237552e-05, 6.852018e-06, 5.812761e-06,
  3.340918e-07, 2.381915e-07, 1.280915e-07, 3.597199e-07, 1.233044e-06, 
    6.469271e-06, 2.454398e-05, 2.909916e-05, 2.306407e-05, 4.987634e-05, 
    3.63613e-05, 2.824672e-05, 1.654923e-05, 9.312451e-06, 5.160993e-06,
  1.689221e-07, 5.395545e-09, 1.811449e-07, 7.676675e-07, 3.974877e-06, 
    7.866285e-06, 2.578349e-05, 5.946639e-05, 5.49094e-05, 4.170472e-05, 
    3.264385e-05, 3.199396e-05, 1.617818e-05, 8.352903e-06, 5.157142e-06,
  3.193998e-07, 2.281513e-07, 8.374851e-07, 4.564908e-06, 7.520713e-06, 
    1.202709e-05, 3.085612e-05, 4.565046e-05, 3.524598e-05, 3.504802e-05, 
    3.708022e-05, 3.505298e-05, 1.493833e-05, 6.992681e-06, 5.032644e-06,
  1.632532e-06, 8.298836e-07, 5.394475e-06, 7.944098e-06, 1.220594e-05, 
    3.063892e-05, 4.549322e-05, 5.287751e-05, 4.500811e-05, 4.129663e-05, 
    3.706639e-05, 2.693567e-05, 1.1716e-05, 6.350873e-06, 4.365369e-06,
  1.884061e-07, 2.105094e-06, 4.225267e-05, 5.717297e-05, 4.785026e-05, 
    5.49584e-05, 5.49488e-05, 4.993537e-05, 4.047313e-05, 3.477364e-05, 
    2.877654e-05, 1.681646e-05, 6.564568e-06, 2.596992e-06, 1.371531e-06,
  4.946742e-05, 2.748588e-05, 1.891292e-05, 4.088505e-05, 8.894761e-05, 
    0.0001303004, 0.0001605006, 0.0001865876, 0.0001918969, 0.0001737485, 
    0.0001485556, 0.0001281684, 0.0001067343, 6.9815e-05, 1.889831e-05,
  0.0002939305, 0.0002468555, 0.0002007448, 0.000199407, 0.0001882382, 
    0.0001713263, 0.0001091593, 5.560452e-05, 2.90376e-05, 2.966675e-05, 
    2.672828e-05, 3.191287e-05, 3.908796e-05, 3.97701e-05, 1.366501e-05,
  0.0003382408, 0.0002966511, 0.0002558414, 0.0002040488, 0.0001144879, 
    5.244252e-05, 1.403227e-05, 6.608504e-06, 3.926149e-06, 4.063079e-06, 
    4.430528e-06, 8.607247e-06, 1.741773e-05, 2.130755e-05, 1.637181e-05,
  0.0002105539, 0.0001900147, 0.0001446507, 8.237961e-05, 2.372291e-05, 
    2.97477e-06, 2.30912e-06, 2.438522e-06, 8.420415e-07, 3.945929e-06, 
    4.095562e-06, 8.401155e-06, 1.678075e-05, 2.039959e-05, 2.165539e-05,
  2.771424e-05, 2.097184e-05, 1.297812e-05, 6.760443e-06, 4.352262e-06, 
    5.440804e-06, 3.848804e-06, 3.180863e-06, 1.568267e-06, 3.66239e-07, 
    2.972267e-06, 9.260754e-06, 2.034335e-05, 2.047599e-05, 2.284881e-05,
  4.650096e-06, 4.467095e-06, 2.860265e-06, 2.688545e-06, 4.26875e-06, 
    5.584617e-06, 8.420006e-06, 3.370052e-06, 1.870766e-06, 2.701039e-06, 
    4.065597e-06, 8.243637e-06, 1.969788e-05, 2.087834e-05, 1.952924e-05,
  3.57055e-06, 5.032567e-06, 4.577975e-06, 3.041315e-06, 4.087425e-06, 
    4.952666e-06, 5.531354e-06, 8.532677e-06, 1.09883e-05, 6.644395e-06, 
    4.141948e-06, 7.411052e-06, 1.649797e-05, 1.895092e-05, 1.200176e-05,
  4.422766e-06, 5.81235e-06, 6.502257e-06, 5.447669e-06, 2.744794e-06, 
    3.045798e-06, 8.937664e-06, 2.534161e-05, 2.868591e-05, 2.920906e-05, 
    2.074456e-05, 1.069106e-05, 1.925584e-05, 1.988547e-05, 1.105813e-05,
  5.618391e-06, 3.152634e-06, 2.613845e-06, 2.245689e-06, 5.747503e-06, 
    5.847646e-06, 1.835533e-05, 3.09588e-05, 3.663174e-05, 4.171679e-05, 
    3.467384e-05, 2.072148e-05, 2.577609e-05, 2.528816e-05, 1.086984e-05,
  3.765324e-06, 3.762976e-06, 2.103256e-06, 3.669016e-06, 4.913247e-06, 
    4.992665e-06, 9.695449e-06, 1.24199e-05, 1.775689e-05, 2.013382e-05, 
    1.8748e-05, 2.085981e-05, 2.467438e-05, 1.911841e-05, 1.431613e-05,
  4.137768e-07, 8.603013e-07, 6.479875e-07, 2.842469e-06, 2.630467e-06, 
    2.494636e-06, 5.618427e-06, 1.231248e-05, 2.664713e-05, 2.348684e-05, 
    2.159283e-05, 2.035031e-05, 1.875299e-05, 3.340933e-05, 6.477744e-05,
  1.113073e-05, 6.463021e-06, 6.236363e-06, 1.152875e-05, 3.675618e-05, 
    6.250764e-05, 7.996574e-05, 9.458941e-05, 0.0001018119, 9.912252e-05, 
    9.374091e-05, 9.641955e-05, 8.282917e-05, 8.981829e-05, 9.578004e-05,
  9.844197e-05, 8.950161e-05, 6.913004e-05, 8.058715e-05, 0.0001324312, 
    0.0001778564, 0.0001754605, 0.0001615509, 0.000157529, 0.000159734, 
    0.0001478783, 0.0001301626, 0.0001173198, 0.0001018688, 0.0001205608,
  0.0001459567, 0.0001951866, 0.0001909095, 0.0001836673, 0.0001914191, 
    0.0001436942, 0.0001805015, 0.0001676433, 0.00013523, 0.0001156476, 
    9.799752e-05, 7.459956e-05, 6.833801e-05, 7.365737e-05, 8.411792e-05,
  6.549548e-05, 0.0001078801, 0.0001222138, 0.0001003681, 9.47441e-05, 
    0.000104617, 5.898853e-05, 7.02547e-05, 0.0001399298, 0.0001204871, 
    8.83414e-05, 6.334551e-05, 4.012885e-05, 3.370461e-05, 3.893817e-05,
  1.275258e-05, 1.919025e-05, 2.44829e-05, 2.578673e-05, 2.040225e-05, 
    1.930484e-05, 1.928208e-05, 4.127424e-05, 5.066923e-05, 3.635948e-05, 
    2.62764e-05, 1.43103e-05, 8.887157e-06, 9.695143e-06, 1.365529e-05,
  6.569357e-06, 9.221552e-06, 4.806639e-06, 4.967509e-06, 4.702216e-06, 
    4.841904e-06, 4.015899e-06, 6.92914e-06, 1.169126e-05, 1.070982e-05, 
    8.034664e-06, 5.810272e-06, 5.381275e-06, 6.288982e-06, 1.128975e-05,
  6.152326e-06, 5.715471e-06, 3.206276e-06, 3.18522e-06, 2.053019e-06, 
    4.976106e-06, 4.646276e-06, 3.756636e-06, 3.487228e-06, 5.428966e-06, 
    6.919101e-06, 5.48077e-06, 5.077287e-06, 9.093308e-06, 1.023026e-05,
  7.833988e-06, 2.013917e-06, 2.255937e-06, 4.750069e-06, 3.646955e-06, 
    3.434919e-06, 4.63988e-06, 5.654545e-06, 5.117258e-06, 4.497586e-06, 
    5.708629e-06, 7.209864e-06, 5.879091e-06, 1.128349e-05, 7.950074e-06,
  6.786358e-06, 1.536359e-06, 1.198545e-06, 4.406839e-06, 4.703102e-06, 
    3.796576e-06, 5.767257e-06, 8.438149e-06, 7.712628e-06, 4.77482e-06, 
    5.531161e-06, 5.586976e-06, 5.512582e-06, 4.880228e-06, 4.723136e-06,
  0.000384161, 0.0001901183, 6.929762e-05, 3.406258e-05, 1.776729e-05, 
    1.019573e-05, 1.399835e-06, 1.900097e-08, 1.308973e-07, 9.681722e-07, 
    2.520936e-06, 2.728149e-06, 5.863787e-06, 1.886106e-05, 1.229915e-05,
  0.0003003632, 0.0002811599, 0.0001777928, 9.287971e-05, 2.983528e-05, 
    6.899572e-06, 1.62108e-07, 1.28451e-08, 1.153254e-07, 3.119427e-07, 
    1.211596e-06, 4.279444e-06, 1.098475e-05, 3.655463e-05, 2.010872e-05,
  0.0001262678, 0.000141637, 9.957921e-05, 4.86391e-05, 1.154197e-05, 
    5.994822e-06, 7.602474e-07, 7.666343e-08, 5.104543e-07, 7.957319e-07, 
    1.75128e-06, 6.795833e-06, 1.253357e-05, 2.071067e-05, 2.483386e-05,
  6.82537e-06, 9.864296e-06, 9.450957e-06, 4.849647e-06, 1.4395e-06, 
    1.831993e-06, 1.549016e-05, 4.465361e-07, 7.968052e-07, 3.306748e-06, 
    6.057935e-06, 7.421292e-06, 8.161213e-06, 1.1893e-05, 2.055197e-05,
  2.576198e-06, 3.353693e-06, 3.661235e-06, 2.636621e-06, 2.661968e-06, 
    1.782414e-06, 2.43734e-06, 8.692353e-06, 1.472236e-05, 9.136469e-06, 
    1.731411e-05, 1.724035e-05, 1.335489e-05, 1.613071e-05, 3.25145e-05,
  3.805676e-06, 3.247841e-06, 3.713739e-06, 2.117585e-06, 1.551752e-06, 
    2.051031e-06, 3.609546e-06, 4.549301e-06, 5.479133e-06, 7.405362e-06, 
    2.006565e-05, 3.382065e-05, 4.397351e-05, 5.186226e-05, 6.175668e-05,
  5.527605e-06, 3.710242e-06, 2.586114e-06, 2.85858e-06, 4.194448e-06, 
    4.462929e-06, 5.780243e-06, 4.704702e-06, 5.295444e-06, 8.391251e-06, 
    1.640815e-05, 2.156228e-05, 4.204553e-05, 5.391487e-05, 3.800068e-05,
  6.34721e-06, 2.863738e-06, 2.211409e-06, 5.369318e-06, 4.816938e-06, 
    4.95099e-06, 3.495485e-06, 4.033541e-06, 6.494188e-06, 8.726352e-06, 
    1.611563e-05, 1.404014e-05, 2.238565e-05, 2.351768e-05, 1.736638e-05,
  6.080586e-06, 1.747996e-06, 2.117109e-06, 7.026777e-06, 4.537689e-06, 
    6.014006e-06, 3.918153e-06, 2.768318e-06, 3.099628e-06, 4.148657e-06, 
    1.146003e-05, 1.391573e-05, 1.233312e-05, 1.280622e-05, 7.653259e-06,
  2.300719e-06, 2.434293e-06, 3.74928e-06, 3.279286e-06, 3.233303e-06, 
    3.03204e-06, 3.158003e-06, 2.307919e-06, 3.501487e-06, 1.447525e-06, 
    9.054722e-06, 1.154502e-05, 5.964357e-06, 6.118541e-06, 5.991289e-06,
  1.18644e-05, 4.500873e-06, 2.115623e-06, 5.630082e-06, 9.209676e-07, 
    3.38927e-06, 1.239014e-05, 1.024726e-05, 6.752086e-06, 5.091524e-06, 
    5.514629e-06, 5.080251e-06, 5.249619e-06, 3.013818e-06, 3.958578e-06,
  9.541825e-05, 8.549583e-05, 6.264204e-05, 5.441114e-05, 3.680338e-05, 
    3.4434e-05, 2.834329e-05, 2.306508e-05, 2.142669e-05, 2.267187e-05, 
    1.904234e-05, 1.364263e-05, 5.415781e-06, 5.842224e-06, 5.800077e-06,
  0.0001752641, 0.0001970042, 0.0002001279, 0.0001888102, 0.0001288289, 
    0.0001392783, 9.410972e-05, 5.654791e-05, 4.051752e-05, 3.434722e-05, 
    2.213718e-05, 1.253016e-05, 3.928658e-06, 4.341863e-06, 5.466675e-06,
  0.0001052766, 0.0001752743, 0.0001966651, 0.0001883942, 0.0001725992, 
    9.804912e-05, 0.0001377881, 0.000106635, 7.420794e-05, 4.721642e-05, 
    3.601947e-05, 1.529277e-05, 7.233553e-06, 3.023192e-06, 5.952856e-06,
  2.138256e-05, 5.332571e-05, 8.498751e-05, 8.84553e-05, 0.0001039815, 
    0.0001169445, 4.857585e-05, 8.674481e-05, 9.254582e-05, 4.249943e-05, 
    3.414778e-05, 8.379499e-06, 4.85093e-06, 3.960371e-06, 9.287319e-06,
  4.916831e-06, 9.943153e-06, 2.265314e-05, 3.637608e-05, 3.984183e-05, 
    5.578074e-05, 6.009778e-05, 1.81637e-05, 1.036329e-05, 1.553456e-05, 
    8.131494e-06, 2.45567e-06, 2.804434e-06, 9.160167e-06, 1.661879e-05,
  6.019722e-06, 3.073661e-06, 4.340307e-06, 9.103918e-06, 1.386751e-05, 
    1.686234e-05, 2.493563e-05, 3.19419e-05, 1.944754e-05, 8.76488e-06, 
    5.364449e-06, 4.097878e-07, 1.60991e-06, 1.192919e-05, 1.828211e-05,
  5.063775e-06, 3.45053e-06, 1.226641e-06, 2.932715e-06, 4.916266e-06, 
    5.961322e-06, 5.790323e-06, 6.055016e-06, 5.895786e-06, 4.461036e-06, 
    3.177753e-06, 2.114682e-06, 1.383295e-06, 1.092883e-05, 1.37237e-05,
  7.977015e-06, 1.713918e-06, 1.764497e-06, 2.872031e-06, 2.381674e-06, 
    2.639339e-06, 3.558544e-06, 4.355642e-06, 3.865506e-06, 4.147666e-06, 
    3.555106e-06, 3.167919e-06, 1.637408e-06, 1.020444e-05, 1.376132e-05,
  1.973403e-06, 2.024517e-06, 2.373569e-06, 1.623738e-06, 2.144936e-06, 
    1.59362e-06, 4.500351e-06, 3.460634e-06, 3.308527e-07, 4.296347e-06, 
    3.84631e-06, 4.420938e-06, 6.859859e-06, 1.328109e-05, 1.110465e-05,
  2.752676e-06, 1.917036e-06, 1.506785e-05, 7.631961e-05, 1.61785e-05, 
    2.885268e-07, 7.065025e-06, 3.366434e-06, 8.688731e-06, 8.600147e-08, 
    5.165208e-08, 1.101368e-07, 2.118275e-07, 1.240865e-06, 9.677915e-07,
  5.275477e-06, 4.872217e-06, 2.587371e-06, 1.582906e-05, 2.627115e-05, 
    1.302849e-06, 2.606661e-06, 3.075169e-06, 2.808893e-06, 7.070432e-06, 
    1.333611e-07, 7.847387e-07, 1.683622e-06, 3.551018e-06, 1.042632e-06,
  5.297663e-06, 5.2241e-06, 3.960506e-06, 4.457403e-06, 4.291802e-06, 
    7.301289e-06, 2.901123e-06, 9.852087e-07, 3.252471e-06, 6.49703e-06, 
    9.164423e-06, 2.532432e-06, 8.049217e-06, 1.891574e-06, 5.696456e-06,
  4.377638e-06, 6.726222e-06, 7.338283e-06, 4.816916e-06, 8.95845e-06, 
    2.978046e-06, 9.049431e-06, 4.76029e-06, 2.627898e-06, 2.388377e-06, 
    5.218104e-06, 9.300384e-06, 9.731486e-06, 3.253531e-06, 1.457612e-05,
  6.136221e-06, 8.13306e-06, 9.86964e-06, 1.438785e-05, 1.121553e-05, 
    6.913699e-06, 5.0876e-06, 2.639229e-05, 2.710314e-05, 1.076152e-05, 
    2.439907e-05, 1.723778e-05, 1.328058e-05, 1.884859e-05, 4.646628e-05,
  6.70829e-06, 5.427326e-06, 9.168781e-06, 1.779031e-05, 1.81136e-05, 
    2.183073e-05, 3.581342e-05, 7.987302e-06, 6.410161e-06, 6.783618e-05, 
    6.572807e-05, 4.295797e-05, 6.420945e-05, 7.404913e-05, 8.637822e-05,
  9.410211e-06, 4.816217e-06, 3.695424e-06, 1.999555e-05, 1.97123e-05, 
    2.168477e-05, 3.716182e-05, 9.265346e-05, 0.0001439404, 0.0001222752, 
    9.450957e-05, 9.362733e-05, 0.000105168, 0.0001014653, 6.460346e-05,
  8.527129e-06, 4.711717e-06, 3.497023e-06, 6.231729e-06, 1.468894e-05, 
    2.019077e-05, 2.406631e-05, 4.432288e-05, 9.046667e-05, 9.787574e-05, 
    8.942954e-05, 8.081026e-05, 7.993801e-05, 6.536092e-05, 2.083464e-05,
  2.830758e-06, 2.9612e-06, 3.677819e-06, 3.842774e-06, 1.250806e-05, 
    2.505797e-05, 5.080365e-05, 8.305164e-05, 0.0001056214, 0.0001019166, 
    7.643614e-05, 5.929258e-05, 5.039621e-05, 2.692704e-05, 5.136287e-06,
  2.14831e-06, 2.231518e-06, 4.330397e-06, 4.228681e-06, 1.304368e-05, 
    3.836955e-05, 6.440593e-05, 8.91584e-05, 9.022309e-05, 7.287315e-05, 
    6.034249e-05, 4.731334e-05, 3.119857e-05, 1.212358e-05, 5.012777e-06,
  5.918642e-05, 8.614919e-05, 9.851828e-05, 6.610613e-05, 7.146527e-06, 
    1.737335e-06, 7.460935e-06, 8.957199e-06, 1.15206e-05, 1.422903e-07, 
    2.802864e-07, 4.959377e-09, 1.741172e-08, 9.210027e-08, 5.160717e-07,
  2.878695e-05, 2.075289e-05, 2.278368e-05, 7.003683e-05, 5.767717e-05, 
    1.372465e-06, 3.191523e-06, 5.020219e-06, 6.405707e-06, 1.020191e-05, 
    4.566939e-07, 1.170736e-06, 1.49224e-06, 9.069252e-08, 1.749162e-06,
  6.398904e-06, 8.096235e-06, 4.363558e-06, 9.780828e-06, 5.328346e-05, 
    5.936528e-05, 6.598023e-07, 5.5015e-06, 6.22895e-06, 1.076447e-05, 
    1.279941e-05, 8.361322e-06, 8.516244e-06, 1.002128e-06, 1.061028e-07,
  4.308263e-06, 4.682963e-06, 2.379824e-06, 2.963473e-06, 2.481427e-06, 
    3.02626e-05, 3.688321e-05, 1.759583e-06, 2.928952e-06, 8.395467e-06, 
    1.20118e-05, 1.337296e-05, 5.966037e-06, 3.699069e-06, 9.797969e-08,
  1.700078e-06, 5.318815e-06, 2.732038e-06, 1.581243e-06, 2.857618e-06, 
    1.887031e-06, 1.459132e-05, 1.911064e-05, 1.106923e-05, 3.380178e-06, 
    6.311506e-06, 9.736894e-06, 1.187874e-05, 4.049289e-06, 1.315153e-06,
  1.174463e-06, 5.423818e-06, 3.104041e-06, 1.403106e-06, 3.338268e-06, 
    2.7401e-06, 2.363208e-06, 2.891863e-06, 1.627768e-06, 8.178349e-07, 
    3.047774e-06, 7.124852e-06, 7.174e-06, 6.541105e-06, 4.564696e-06,
  2.033298e-06, 3.992001e-06, 4.232915e-06, 1.155657e-06, 2.507601e-06, 
    3.661428e-06, 2.310895e-06, 1.406115e-06, 2.951982e-06, 2.29098e-06, 
    1.560806e-06, 1.303401e-06, 2.830177e-06, 4.164892e-06, 2.106685e-05,
  1.678019e-06, 2.569211e-06, 4.624319e-06, 1.532989e-06, 3.048266e-06, 
    3.639355e-06, 2.079136e-06, 2.048776e-06, 1.498535e-06, 1.234602e-06, 
    2.254108e-06, 2.764638e-06, 3.569952e-06, 1.195628e-05, 4.436642e-05,
  2.623695e-06, 2.362427e-06, 5.4351e-06, 9.540685e-07, 2.848915e-06, 
    3.866e-06, 2.783515e-06, 3.863993e-06, 7.318364e-06, 3.932028e-06, 
    3.614686e-06, 4.500136e-06, 1.383594e-05, 4.079557e-05, 4.997733e-05,
  2.11246e-06, 2.184241e-06, 3.201791e-06, 2.239081e-06, 2.956437e-06, 
    3.262216e-06, 6.042126e-06, 8.276013e-06, 1.160978e-05, 8.011248e-06, 
    9.663162e-06, 1.736636e-05, 3.627808e-05, 5.494072e-05, 5.372731e-05,
  0.0005030062, 0.0001558666, 5.775887e-05, 6.341383e-06, 5.583871e-06, 
    4.38295e-06, 6.374818e-06, 4.484948e-06, 5.57471e-06, 1.547525e-07, 
    2.630606e-08, 2.747471e-09, 3.700864e-07, 1.894648e-08, 2.665784e-07,
  0.0004493719, 0.00025492, 0.0001351986, 7.365417e-05, 1.000751e-05, 
    3.18993e-06, 3.799345e-06, 3.348254e-06, 9.396372e-06, 1.604937e-05, 
    1.481096e-06, 1.420596e-05, 1.483858e-05, 5.879825e-07, 1.982397e-07,
  0.0002491354, 0.0003036468, 0.0001753387, 0.000133376, 3.976267e-05, 
    1.974126e-05, 5.917193e-06, 8.364481e-06, 7.003922e-06, 1.239781e-05, 
    1.4027e-05, 1.080457e-05, 1.317407e-05, 9.714905e-06, 2.932764e-07,
  7.047668e-05, 0.0001709874, 0.0002070343, 0.0001429371, 0.0001091089, 
    2.248178e-05, 3.305396e-05, 6.61881e-06, 5.348347e-06, 9.172345e-06, 
    6.634879e-06, 9.672035e-06, 9.818003e-06, 1.36906e-05, 1.321491e-05,
  8.353342e-06, 4.539646e-05, 0.0001201523, 0.0001429017, 0.0001271873, 
    0.000117857, 1.185888e-05, 1.776133e-05, 1.972553e-05, 4.659362e-06, 
    4.835405e-06, 5.761331e-06, 8.051049e-06, 9.992542e-06, 1.626352e-05,
  8.055529e-07, 6.446124e-06, 2.824721e-05, 7.930391e-05, 0.0001163647, 
    0.0001216886, 0.0001158023, 3.694814e-06, 9.695235e-07, 1.038541e-06, 
    1.432517e-06, 2.049062e-06, 4.635258e-06, 6.905907e-06, 1.028011e-05,
  1.022065e-07, 8.119676e-07, 4.326796e-06, 1.60264e-05, 5.325566e-05, 
    8.76809e-05, 0.0001068124, 0.0001109356, 4.167564e-05, 4.378237e-06, 
    1.680563e-06, 4.535127e-07, 7.748412e-07, 4.268693e-06, 5.766542e-06,
  3.376393e-07, 6.828632e-08, 4.871071e-07, 4.433698e-06, 1.253026e-05, 
    4.281037e-05, 7.014209e-05, 5.848556e-05, 3.93087e-05, 2.40214e-05, 
    9.709534e-06, 1.01229e-06, 1.914175e-07, 2.766826e-07, 1.11813e-06,
  1.862482e-06, 2.118187e-08, 2.778557e-06, 3.037838e-06, 4.317501e-06, 
    7.581244e-06, 1.911152e-05, 4.287743e-05, 4.814212e-05, 3.213134e-05, 
    1.097476e-05, 1.215158e-06, 7.406776e-07, 4.237284e-07, 4.72889e-07,
  2.279471e-07, 8.902628e-08, 2.292859e-07, 3.238455e-06, 2.732606e-06, 
    4.144564e-06, 4.583095e-06, 5.953108e-06, 1.24029e-05, 1.513995e-05, 
    9.794424e-06, 3.800723e-06, 1.701842e-06, 1.23723e-06, 1.098469e-06,
  5.315629e-05, 1.778166e-05, 1.324532e-06, 1.179163e-08, 6.36063e-09, 
    1.635117e-05, 4.699533e-05, 1.100923e-05, 1.165822e-05, 1.787551e-07, 
    5.648144e-08, 7.116004e-11, 3.420546e-08, 1.240077e-08, 3.890361e-10,
  8.622507e-05, 2.014183e-05, 3.177331e-06, 2.624371e-08, 5.578366e-08, 
    1.295059e-05, 4.805432e-05, 1.80147e-05, 3.717415e-06, 2.073072e-05, 
    2.167061e-07, 1.016231e-05, 2.047964e-06, 1.913458e-08, 8.355717e-09,
  0.0001685021, 6.546926e-05, 7.914487e-06, 1.923991e-07, 1.002157e-07, 
    3.054795e-05, 5.475919e-05, 3.640288e-05, 2.678906e-06, 7.765671e-06, 
    1.565345e-05, 2.35146e-06, 2.72435e-06, 8.976797e-06, 1.660945e-08,
  0.0001896875, 0.0001524061, 5.028877e-05, 1.687033e-06, 2.732199e-07, 
    9.276078e-06, 6.957883e-05, 5.769591e-05, 3.533307e-06, 1.025557e-05, 
    5.951209e-06, 6.229978e-06, 5.902653e-06, 7.470656e-06, 1.402716e-05,
  8.116505e-05, 0.0001750793, 0.0001377715, 4.924429e-05, 1.272972e-05, 
    4.665556e-05, 1.033753e-05, 7.252801e-05, 2.05009e-05, 5.65872e-06, 
    1.311672e-05, 8.840202e-06, 6.221465e-06, 1.173791e-05, 1.605813e-05,
  2.342481e-05, 0.0001016399, 0.0001505653, 0.0001275743, 9.64938e-05, 
    5.405631e-05, 2.437443e-05, 2.000268e-05, 1.896261e-06, 4.661332e-06, 
    6.753272e-06, 6.264058e-06, 6.320614e-06, 6.255615e-06, 1.007467e-05,
  5.057602e-07, 2.184147e-05, 8.199342e-05, 0.0001445798, 0.0001565742, 
    8.962808e-05, 2.716684e-05, 6.36297e-05, 1.839108e-05, 4.79889e-06, 
    6.126572e-06, 5.11755e-06, 4.263494e-06, 5.268809e-06, 5.94133e-06,
  1.216105e-06, 5.777878e-06, 2.045435e-05, 7.869246e-05, 0.0001439636, 
    0.0001525985, 6.221713e-05, 2.239099e-05, 1.519092e-05, 5.917581e-06, 
    4.037255e-06, 4.553749e-06, 3.455888e-06, 4.475103e-06, 5.124519e-06,
  1.631368e-06, 9.947665e-07, 5.432198e-06, 1.973142e-05, 7.635118e-05, 
    0.0001446078, 0.0001624199, 0.0001102682, 5.798394e-05, 2.474498e-05, 
    1.785689e-05, 9.093082e-06, 4.017948e-06, 3.232326e-06, 4.59913e-06,
  7.578137e-07, 2.19984e-07, 1.600646e-06, 4.513123e-06, 1.693958e-05, 
    7.812857e-05, 0.0001318391, 0.0001398519, 0.0001123476, 7.780647e-05, 
    4.195979e-05, 1.4858e-05, 6.406699e-06, 3.874874e-06, 2.855839e-06,
  8.068814e-05, 2.963968e-05, 1.820964e-06, 5.70356e-07, 2.045339e-08, 
    8.76278e-08, 1.229898e-05, 0.0001326726, 2.002453e-05, 6.19449e-06, 
    1.092543e-08, 2.052598e-25, 3.010437e-12, 1.507175e-11, 7.119658e-11,
  8.162703e-05, 3.0103e-05, 7.165615e-06, 1.037402e-06, 2.323887e-07, 
    4.030123e-08, 1.5166e-05, 0.0001191901, 8.294125e-06, 1.287781e-05, 
    1.708833e-08, 2.766468e-10, 1.03674e-13, 6.998988e-12, 3.205724e-11,
  7.883955e-05, 3.80027e-05, 1.294483e-05, 2.342473e-06, 6.228877e-07, 
    2.474731e-07, 2.236015e-05, 0.0001248187, 5.313088e-06, 1.227313e-05, 
    1.972305e-06, 8.778837e-09, 9.282866e-07, 1.341207e-05, 9.66413e-11,
  5.04971e-05, 5.122949e-05, 1.452738e-05, 5.788771e-06, 3.582131e-07, 
    3.680166e-08, 3.989632e-05, 8.215888e-05, 5.845768e-06, 7.975137e-06, 
    2.333134e-06, 1.502779e-06, 4.964587e-06, 8.244678e-06, 4.879592e-06,
  3.182319e-05, 7.35093e-05, 2.741939e-05, 7.632856e-06, 1.326191e-06, 
    8.487547e-07, 2.538579e-05, 6.642153e-05, 1.755342e-05, 5.814923e-06, 
    5.185285e-06, 2.095352e-06, 3.853183e-06, 9.281107e-06, 1.343942e-05,
  1.830383e-05, 4.978305e-05, 4.872248e-05, 1.883002e-05, 2.050396e-05, 
    6.151563e-06, 1.133316e-05, 2.220876e-05, 8.828348e-07, 5.99643e-06, 
    7.000584e-06, 2.047917e-06, 5.36843e-06, 2.780647e-06, 5.299942e-06,
  2.882669e-06, 2.407962e-05, 4.559908e-05, 4.365638e-05, 8.079599e-05, 
    5.08943e-05, 1.211001e-05, 1.350057e-05, 2.373962e-06, 5.897387e-06, 
    9.509585e-06, 1.371807e-06, 3.307807e-06, 1.744955e-06, 3.090053e-06,
  6.587253e-07, 1.125467e-05, 1.483797e-05, 4.902978e-05, 0.0001250223, 
    0.0001283348, 2.77338e-05, 3.672043e-06, 2.302375e-06, 2.098782e-06, 
    5.761357e-06, 2.029296e-06, 2.11799e-06, 3.253412e-06, 2.920803e-06,
  9.37107e-07, 1.912092e-06, 4.949651e-06, 1.255686e-05, 0.0001015194, 
    0.0001558507, 8.439616e-05, 4.383929e-06, 3.863826e-06, 2.859053e-06, 
    1.864213e-06, 4.669436e-06, 5.926095e-06, 2.833095e-06, 1.341465e-06,
  1.219691e-06, 6.473096e-07, 7.813104e-07, 3.598291e-06, 4.246258e-05, 
    0.0001639377, 0.0001240859, 5.409143e-05, 1.305388e-05, 4.919177e-06, 
    2.462655e-06, 3.495879e-06, 4.910356e-06, 3.308768e-06, 2.832701e-06,
  7.947369e-06, 4.405259e-06, 6.423565e-06, 4.526877e-06, 4.411527e-06, 
    2.724794e-06, 1.065876e-06, 3.223993e-06, 2.342774e-05, 4.507113e-06, 
    3.442319e-06, 1.179401e-07, 3.88072e-09, 3.250308e-09, 1.675692e-09,
  3.273921e-06, 3.509487e-06, 3.882529e-06, 5.166414e-06, 6.345642e-06, 
    4.100568e-06, 1.227776e-06, 8.535409e-06, 1.410916e-05, 7.139808e-06, 
    3.031824e-06, 1.481075e-07, 4.434132e-08, 1.354031e-06, 1.009753e-06,
  5.702151e-06, 6.142648e-06, 3.977022e-06, 4.934268e-06, 4.074514e-06, 
    8.007838e-06, 1.055482e-06, 2.418185e-05, 1.48488e-05, 9.110924e-06, 
    1.388936e-06, 2.157836e-07, 1.468243e-06, 1.265424e-05, 1.243068e-07,
  8.191632e-06, 1.156613e-05, 8.413035e-06, 8.623075e-06, 3.730313e-06, 
    2.272983e-06, 1.806548e-05, 3.841209e-05, 1.35112e-05, 6.599854e-06, 
    5.589148e-06, 1.527636e-06, 8.488384e-06, 1.18255e-05, 7.660522e-08,
  8.580339e-06, 1.780142e-05, 1.262389e-05, 6.893963e-06, 5.309301e-06, 
    4.612375e-06, 3.976746e-05, 5.190476e-05, 1.565012e-05, 7.515059e-06, 
    9.652387e-06, 4.139248e-06, 6.012268e-06, 1.150448e-05, 1.296629e-05,
  6.738239e-06, 1.622464e-05, 2.083663e-05, 7.129526e-06, 6.44651e-06, 
    9.293573e-06, 6.714836e-05, 4.862268e-05, 1.595576e-06, 9.814918e-06, 
    8.139425e-06, 6.003373e-06, 8.483759e-06, 8.463433e-06, 8.802011e-06,
  5.042069e-06, 1.066963e-05, 2.637637e-05, 1.406313e-05, 8.117722e-06, 
    9.590418e-06, 6.864582e-05, 9.69582e-05, 9.301815e-06, 1.514316e-05, 
    9.206085e-06, 6.85917e-06, 1.073191e-05, 9.867138e-06, 9.94261e-06,
  3.04571e-06, 1.121406e-05, 2.553615e-05, 2.792297e-05, 7.652616e-06, 
    1.238162e-05, 6.588375e-05, 6.108329e-05, 6.444955e-06, 1.375494e-05, 
    6.99149e-06, 5.333548e-06, 1.051123e-05, 8.087361e-06, 9.100104e-06,
  1.479104e-06, 1.039318e-05, 2.265863e-05, 4.15268e-05, 2.005401e-05, 
    2.494932e-05, 5.914433e-05, 6.015715e-05, 9.455612e-06, 1.213074e-05, 
    8.025627e-06, 8.192392e-06, 9.001926e-06, 9.710556e-06, 7.572178e-06,
  1.482705e-06, 4.9099e-06, 1.606293e-05, 5.049585e-05, 5.247984e-05, 
    5.327123e-05, 6.071269e-05, 5.376215e-05, 1.056967e-05, 8.913834e-06, 
    4.666862e-06, 8.125743e-06, 7.035312e-06, 6.050684e-06, 5.780911e-06,
  5.132506e-07, 2.047324e-07, 1.900865e-06, 2.621426e-06, 3.496478e-06, 
    3.415145e-06, 4.100834e-06, 3.600638e-06, 2.428525e-07, 3.620529e-07, 
    7.880131e-06, 5.551718e-06, 1.207358e-05, 3.623887e-06, 5.536934e-07,
  4.49316e-09, 1.751149e-07, 5.905045e-07, 2.96311e-06, 5.637949e-06, 
    1.735262e-06, 1.361547e-06, 9.281378e-07, 1.000309e-07, 1.029857e-06, 
    2.520606e-06, 6.83809e-06, 2.238723e-06, 6.874802e-06, 1.23216e-06,
  1.960552e-07, 1.569406e-07, 1.302025e-06, 3.735731e-06, 7.963295e-06, 
    9.733858e-06, 3.60275e-07, 1.208467e-06, 8.375141e-08, 3.814941e-06, 
    5.489115e-06, 4.626103e-06, 2.219782e-06, 2.200762e-06, 2.429799e-07,
  2.277577e-08, 5.328938e-07, 3.628842e-06, 4.668108e-06, 4.138758e-06, 
    9.67055e-06, 8.210268e-06, 1.210342e-07, 9.02286e-08, 7.215547e-06, 
    1.329602e-05, 1.093197e-05, 4.026867e-06, 2.132093e-06, 3.592665e-08,
  7.808097e-08, 5.985646e-07, 3.434517e-06, 5.121937e-06, 4.815425e-06, 
    5.313701e-06, 5.969575e-06, 1.054464e-05, 2.344109e-06, 3.51703e-06, 
    1.738971e-05, 1.634729e-05, 4.541886e-06, 3.73595e-06, 2.589311e-06,
  7.371389e-07, 4.352218e-07, 2.3752e-06, 2.502064e-06, 2.820359e-06, 
    3.636486e-06, 4.460229e-06, 3.313147e-06, 6.417713e-06, 3.757165e-06, 
    1.130701e-05, 1.881647e-05, 7.204673e-06, 1.466913e-06, 2.238158e-06,
  2.289828e-06, 2.359888e-06, 4.195808e-06, 2.123959e-06, 1.586173e-06, 
    1.748687e-06, 4.458313e-06, 4.563777e-06, 4.595629e-06, 3.733014e-06, 
    7.176203e-06, 1.560568e-05, 1.101439e-05, 1.963749e-06, 2.863261e-06,
  4.106101e-06, 5.12097e-06, 9.528677e-06, 9.730598e-06, 4.541092e-06, 
    2.440082e-06, 3.305631e-06, 2.176491e-06, 3.182518e-06, 5.04321e-06, 
    5.937639e-06, 1.168603e-05, 1.69531e-05, 3.869014e-06, 2.747339e-06,
  8.759085e-06, 9.409358e-06, 1.5124e-05, 1.516767e-05, 5.098119e-06, 
    2.755855e-06, 4.689511e-06, 1.406426e-06, 2.450965e-06, 4.265859e-06, 
    5.006654e-06, 9.862553e-06, 2.06763e-05, 8.494744e-06, 7.596824e-06,
  8.291918e-06, 8.729433e-06, 1.546256e-05, 2.330941e-05, 1.512681e-05, 
    5.9212e-06, 5.012377e-06, 2.990155e-06, 4.304609e-06, 4.302113e-06, 
    4.535686e-06, 6.726454e-06, 1.755487e-05, 9.045098e-06, 7.838393e-06,
  4.31121e-09, 3.516037e-08, 4.952718e-07, 1.883714e-06, 3.765735e-06, 
    2.766744e-06, 2.369893e-06, 4.637514e-06, 3.713476e-06, 6.332411e-06, 
    3.439291e-06, 1.870285e-06, 4.48181e-07, 6.652729e-08, 7.361859e-08,
  2.164003e-08, 3.085102e-08, 1.879883e-08, 4.179065e-07, 4.000275e-06, 
    6.107191e-07, 6.466792e-07, 1.257575e-06, 3.881923e-06, 1.065642e-05, 
    4.60424e-06, 2.014811e-06, 1.639836e-06, 2.676942e-06, 5.311339e-06,
  1.783442e-07, 2.274084e-08, 9.389782e-08, 3.157288e-07, 9.11025e-07, 
    7.063614e-06, 1.985206e-07, 1.690855e-06, 1.311166e-06, 1.931627e-05, 
    5.716719e-06, 9.51559e-07, 5.067443e-06, 7.922281e-06, 4.563819e-07,
  6.320097e-07, 2.423662e-07, 1.117632e-06, 2.815509e-07, 1.191767e-06, 
    1.870248e-06, 5.198242e-06, 5.437837e-08, 1.480592e-07, 8.71796e-06, 
    9.503712e-06, 2.838931e-06, 7.554742e-06, 1.087679e-05, 1.281537e-07,
  9.060742e-09, 1.972817e-08, 7.068929e-07, 1.265563e-06, 1.169998e-06, 
    1.115628e-06, 3.464067e-06, 2.479568e-06, 3.795855e-06, 1.145582e-06, 
    8.100205e-06, 1.176885e-05, 6.114071e-06, 8.011136e-06, 3.813829e-06,
  3.51737e-07, 5.067248e-07, 1.292138e-06, 8.703175e-07, 1.083539e-07, 
    9.585376e-07, 1.060566e-06, 2.353572e-06, 5.935485e-06, 1.257698e-06, 
    5.953702e-07, 1.204511e-05, 5.141228e-06, 8.695578e-06, 4.652111e-06,
  3.017029e-06, 3.582433e-06, 3.940171e-06, 4.815094e-06, 4.717233e-06, 
    1.944431e-06, 1.236397e-06, 1.613786e-06, 2.1069e-06, 1.911864e-06, 
    1.341584e-06, 2.364174e-06, 9.312658e-06, 8.525692e-06, 3.59332e-06,
  4.987256e-06, 3.565184e-06, 4.530831e-06, 6.387419e-06, 4.498636e-06, 
    4.616617e-06, 3.40939e-06, 3.128582e-06, 1.613143e-06, 1.806191e-06, 
    1.746757e-06, 1.040848e-06, 6.796685e-06, 7.251197e-06, 4.336337e-06,
  9.114415e-06, 6.036812e-06, 5.219517e-06, 3.903279e-06, 5.001434e-06, 
    2.886504e-06, 3.825489e-06, 3.620652e-06, 2.336184e-06, 1.894108e-06, 
    2.062875e-06, 1.091066e-06, 4.376878e-06, 8.398772e-06, 8.507018e-06,
  7.697294e-06, 7.683064e-06, 5.335255e-06, 4.780029e-06, 3.518667e-06, 
    3.438246e-06, 4.61609e-06, 4.266741e-06, 4.424621e-06, 3.04527e-06, 
    2.498964e-06, 2.668529e-06, 3.7478e-06, 3.356839e-06, 1.112358e-05 ;

 prw =
  2.036014, 2.124499, 2.119642, 2.054166, 1.88181, 1.658246, 1.541344, 
    1.476863, 1.429647, 1.29525, 1.309881, 1.31477, 1.256765, 1.265899, 
    1.246869,
  2.042166, 2.0126, 2.021447, 2.007962, 1.868574, 1.587368, 1.474908, 
    1.37251, 1.350663, 1.283472, 1.193976, 1.243345, 1.241907, 1.149893, 
    1.176628,
  2.111785, 1.939402, 1.901277, 1.880857, 1.723977, 1.397114, 1.33706, 
    1.23978, 1.196588, 1.177276, 1.123363, 1.149438, 1.18258, 1.193347, 
    1.167726,
  2.366038, 1.938049, 1.779327, 1.693885, 1.628971, 1.438841, 1.048375, 
    1.075261, 1.088357, 1.050704, 1.028553, 1.038929, 1.083523, 1.140173, 
    1.139975,
  2.521959, 2.035335, 1.714991, 1.580541, 1.46528, 1.343131, 1.196122, 
    0.8293736, 0.8102834, 0.9567543, 0.9609662, 0.9658884, 1.002234, 1.06713, 
    1.142902,
  2.423422, 2.059092, 1.734291, 1.55157, 1.427177, 1.278052, 1.17375, 
    1.147495, 1.029498, 0.9568139, 0.92349, 0.9333751, 0.9622366, 1.019358, 
    1.132788,
  2.278565, 1.997543, 1.748291, 1.54159, 1.411964, 1.281725, 1.175069, 
    1.103963, 1.058935, 1.009219, 0.963406, 0.9363506, 0.9692344, 1.012931, 
    1.111831,
  2.153393, 1.98274, 1.749464, 1.569473, 1.422637, 1.273878, 1.182859, 
    1.135532, 1.086018, 1.038717, 0.9962353, 0.9741663, 0.996155, 1.046058, 
    1.132185,
  2.146832, 1.971833, 1.769265, 1.607337, 1.481247, 1.340947, 1.242999, 
    1.179098, 1.137094, 1.076594, 1.050018, 1.031432, 1.057579, 1.126636, 
    1.200978,
  2.201155, 2.031859, 1.86018, 1.702352, 1.564635, 1.43773, 1.347416, 
    1.275562, 1.191596, 1.120213, 1.102757, 1.101996, 1.122254, 1.181631, 
    1.255197,
  2.004152, 2.126981, 1.890525, 1.620552, 1.451821, 1.465685, 1.598991, 
    1.890474, 2.18169, 2.480823, 2.872702, 3.336399, 3.620271, 3.398443, 
    3.112815,
  1.885042, 1.947541, 1.942041, 1.710487, 1.455901, 1.410084, 1.531172, 
    1.716163, 1.980952, 2.244127, 2.603157, 3.030496, 3.313485, 3.059313, 
    2.881178,
  1.650874, 1.645519, 1.68719, 1.635924, 1.436052, 1.241271, 1.439304, 
    1.570002, 1.776262, 2.014865, 2.358258, 2.733421, 2.994879, 2.901547, 
    2.727514,
  1.53552, 1.440826, 1.374271, 1.328929, 1.319849, 1.320294, 1.179388, 
    1.435496, 1.594495, 1.767254, 2.101635, 2.435312, 2.670916, 2.614287, 
    2.523355,
  1.526935, 1.389305, 1.284342, 1.226875, 1.195105, 1.233054, 1.283976, 
    1.03657, 1.180679, 1.506597, 1.805086, 2.116553, 2.362056, 2.359786, 
    2.342415,
  1.636703, 1.458461, 1.307388, 1.210311, 1.148375, 1.114625, 1.148372, 
    1.222117, 1.274301, 1.409709, 1.606081, 1.835571, 2.063927, 2.139172, 
    2.149809,
  1.800845, 1.588599, 1.414718, 1.279848, 1.191923, 1.127294, 1.104859, 
    1.121944, 1.189152, 1.311523, 1.425297, 1.569036, 1.767177, 1.879873, 
    1.918632,
  1.971695, 1.759978, 1.563292, 1.392803, 1.278133, 1.174655, 1.110591, 
    1.102988, 1.125024, 1.203999, 1.258848, 1.354046, 1.503906, 1.618963, 
    1.677801,
  2.092687, 1.93839, 1.750866, 1.57128, 1.39423, 1.276314, 1.190911, 
    1.153596, 1.124337, 1.131094, 1.161449, 1.208133, 1.319413, 1.412319, 
    1.47046,
  2.200639, 2.06552, 1.934187, 1.775814, 1.593537, 1.43521, 1.271584, 
    1.168868, 1.113114, 1.105379, 1.130383, 1.159069, 1.233285, 1.300463, 
    1.354373,
  2.179666, 1.778112, 1.549966, 1.534384, 1.590414, 1.666282, 1.860751, 
    2.025964, 2.209512, 2.406099, 2.428964, 2.244107, 2.245626, 2.491726, 
    2.897235,
  1.905409, 1.562365, 1.497655, 1.535461, 1.646383, 1.784971, 2.015992, 
    2.080303, 2.362989, 2.527198, 2.481583, 2.322342, 2.483794, 2.700888, 
    3.108073,
  1.860934, 1.529795, 1.466675, 1.523592, 1.727452, 1.815641, 2.123094, 
    2.089706, 2.480499, 2.567486, 2.501175, 2.467051, 2.721347, 3.151836, 
    3.224109,
  1.887523, 1.572408, 1.469836, 1.509385, 1.658801, 2.023458, 1.972108, 
    2.188642, 2.41761, 2.480923, 2.535369, 2.661442, 3.003722, 3.33148, 
    3.180763,
  1.922536, 1.620063, 1.504481, 1.480565, 1.62598, 1.942108, 2.339976, 
    2.006105, 2.101439, 2.50307, 2.652372, 2.882663, 3.262797, 3.367057, 
    3.092994,
  1.9878, 1.663803, 1.524991, 1.485403, 1.603973, 1.875471, 2.259758, 
    2.40341, 2.51059, 2.610121, 2.801283, 3.097477, 3.395849, 3.370767, 
    3.001431,
  2.046041, 1.716222, 1.543113, 1.517755, 1.625227, 1.86321, 2.243011, 
    2.477299, 2.651349, 2.803682, 2.956397, 3.261099, 3.460223, 3.334376, 
    3.010609,
  2.157556, 1.831843, 1.594471, 1.540834, 1.634796, 1.840795, 2.168701, 
    2.424442, 2.675078, 2.908178, 3.062994, 3.33493, 3.474738, 3.330117, 
    3.097743,
  2.246712, 1.98288, 1.717635, 1.596406, 1.632608, 1.846367, 2.111862, 
    2.368623, 2.662617, 2.933372, 3.086429, 3.326493, 3.443136, 3.298564, 
    3.148275,
  2.309666, 2.0866, 1.869021, 1.723249, 1.688545, 1.814174, 2.029509, 
    2.267485, 2.559783, 2.792291, 3.028033, 3.273871, 3.344669, 3.23086, 
    3.203682,
  3.055305, 2.832185, 2.498091, 2.394161, 2.256492, 2.356336, 2.298321, 
    1.926842, 1.758348, 1.809908, 1.981845, 1.727213, 1.437757, 1.498875, 
    1.793046,
  3.040552, 2.70498, 2.38677, 2.284971, 2.124019, 2.198784, 2.429556, 
    2.265481, 2.03222, 2.058096, 2.013394, 1.664677, 1.50411, 1.573719, 
    1.983335,
  2.993245, 2.593576, 2.243449, 2.199288, 2.077471, 2.072085, 2.555586, 
    2.457112, 2.303948, 2.153418, 1.972339, 1.601554, 1.580096, 1.853224, 
    2.256481,
  2.898877, 2.459719, 2.1849, 2.190542, 2.312569, 2.568421, 2.281396, 
    2.445759, 2.290865, 2.082767, 1.839483, 1.597921, 1.709783, 2.113593, 
    2.390258,
  2.758655, 2.301917, 2.176519, 2.208518, 2.344545, 2.670683, 2.71104, 
    2.018789, 1.788242, 1.948546, 1.736548, 1.67664, 1.97015, 2.336439, 
    2.402447,
  2.602104, 2.226301, 2.219943, 2.280401, 2.435264, 2.714382, 2.9465, 
    2.546546, 2.089772, 1.904676, 1.740081, 1.893097, 2.234831, 2.437163, 
    2.211511,
  2.456368, 2.196976, 2.267575, 2.407389, 2.561468, 2.849991, 2.858751, 
    2.595422, 2.283296, 2.090522, 1.922557, 2.161715, 2.407193, 2.280069, 
    1.959964,
  2.294868, 2.186431, 2.348787, 2.562814, 2.736404, 2.935253, 2.790833, 
    2.536685, 2.321634, 2.228704, 2.18641, 2.378649, 2.337547, 2.025958, 
    1.695443,
  2.161565, 2.208914, 2.474759, 2.766481, 2.897798, 2.965155, 2.730681, 
    2.594974, 2.496928, 2.523389, 2.412759, 2.401991, 2.102689, 1.768477, 
    1.608011,
  2.114661, 2.296285, 2.686898, 2.88703, 2.976065, 2.949556, 2.753205, 
    2.718222, 2.644098, 2.541462, 2.467788, 2.229278, 1.861447, 1.641367, 
    1.74873,
  2.636564, 2.952397, 3.245565, 3.374597, 3.31058, 3.133308, 2.380275, 
    1.466518, 1.238105, 1.272677, 1.462177, 1.430792, 1.58998, 1.882865, 
    2.063908,
  2.984625, 3.31957, 3.622252, 3.568614, 3.274271, 2.636302, 1.871027, 
    1.368608, 1.307054, 1.454117, 1.499045, 1.529367, 1.764666, 1.916283, 
    2.112662,
  3.189699, 3.515224, 3.721495, 3.510464, 3.034897, 2.014801, 1.89371, 
    1.540183, 1.495031, 1.564011, 1.558415, 1.630996, 1.872533, 2.105292, 
    2.220788,
  3.41937, 3.664707, 3.681489, 3.436942, 3.105665, 2.150332, 1.746749, 
    1.617179, 1.606107, 1.62027, 1.594191, 1.725515, 1.946937, 2.14664, 
    2.254221,
  3.60609, 3.727909, 3.566683, 3.298806, 3.071157, 2.552563, 2.118461, 
    1.468475, 1.377522, 1.635572, 1.646116, 1.802162, 2.009746, 2.187564, 
    2.320002,
  3.685462, 3.672386, 3.380851, 3.142237, 3.027331, 2.933054, 2.669308, 
    2.055202, 1.718687, 1.697269, 1.706842, 1.861355, 2.045607, 2.211203, 
    2.291915,
  3.714015, 3.542948, 3.19671, 3.014542, 2.97216, 3.062452, 2.823719, 
    2.369753, 2.024556, 1.937291, 1.811673, 1.899188, 2.092017, 2.219777, 
    2.233577,
  3.70303, 3.359107, 2.998073, 2.925783, 2.961287, 3.197894, 2.830941, 
    2.328519, 2.149297, 2.035228, 1.855125, 1.955347, 2.158235, 2.201646, 
    2.185401,
  3.581423, 3.131249, 2.889327, 2.909638, 3.045817, 3.27546, 2.786404, 
    2.355305, 2.260454, 2.164586, 1.926237, 2.046354, 2.206815, 2.149949, 
    2.211332,
  3.361123, 2.969145, 2.902673, 2.989866, 3.15127, 3.292745, 2.684651, 
    2.384241, 2.23958, 2.079775, 2.011202, 2.156992, 2.20347, 2.110844, 
    2.401335,
  2.029093, 2.070578, 1.900426, 2.279298, 2.486137, 2.504626, 2.197853, 
    1.653492, 1.327998, 1.517983, 1.8339, 2.105449, 2.340276, 2.321133, 
    2.154482,
  2.3162, 2.323905, 2.31908, 2.685727, 2.741594, 2.472214, 1.854014, 1.44593, 
    1.304171, 1.570916, 1.885877, 2.247623, 2.562917, 2.467433, 2.281672,
  2.409742, 2.484149, 2.597338, 3.054617, 2.98578, 2.198492, 1.674196, 
    1.351496, 1.323036, 1.599188, 1.958963, 2.391023, 2.740638, 2.754759, 
    2.481947,
  2.466971, 2.608061, 2.82176, 3.321146, 3.330787, 2.676784, 1.582087, 
    1.238673, 1.293441, 1.608985, 1.998054, 2.504348, 2.906297, 2.952834, 
    2.733997,
  2.582218, 2.740689, 3.022678, 3.534821, 3.586303, 3.096498, 2.125746, 
    1.041833, 1.005094, 1.531074, 2.008482, 2.575075, 3.03228, 3.183835, 
    3.168472,
  2.729201, 2.969946, 3.230791, 3.687889, 3.714531, 3.360904, 2.787886, 
    1.721773, 1.27844, 1.570544, 2.013122, 2.639032, 3.045661, 3.274385, 
    3.430741,
  2.884246, 3.143709, 3.436603, 3.801435, 3.796213, 3.46112, 3.017962, 
    2.240917, 1.663899, 1.782495, 2.108341, 2.677844, 3.025493, 3.237813, 
    3.484311,
  3.100317, 3.363107, 3.634044, 3.889158, 3.815321, 3.480026, 3.046467, 
    2.381171, 1.919402, 1.951916, 2.143658, 2.67626, 2.984223, 3.133328, 
    3.39172,
  3.348587, 3.617025, 3.811892, 3.953739, 3.85122, 3.487466, 2.981958, 
    2.437589, 2.103189, 2.123482, 2.200256, 2.656098, 2.900518, 3.033858, 
    3.223168,
  3.629613, 3.847722, 3.892586, 3.992592, 3.865472, 3.504563, 2.921439, 
    2.416131, 2.149781, 2.128368, 2.216006, 2.606405, 2.832075, 2.960068, 
    3.127487,
  2.068769, 2.270184, 1.85374, 1.68072, 1.426476, 1.775929, 1.724522, 
    1.796935, 2.009498, 2.11329, 2.125411, 2.106428, 1.95533, 1.86379, 
    1.899571,
  2.445396, 2.551626, 2.325598, 1.999605, 1.481363, 1.772464, 1.669405, 
    1.752058, 2.0086, 2.23891, 2.281306, 2.248903, 2.060352, 1.794443, 
    1.865601,
  2.853595, 2.751977, 2.637017, 2.324984, 1.636889, 1.473558, 1.596685, 
    1.705081, 2.001976, 2.291899, 2.452512, 2.456524, 2.263733, 2.010987, 
    1.876579,
  3.087267, 2.981964, 2.809227, 2.551567, 2.106863, 1.731829, 1.305034, 
    1.574085, 1.92228, 2.353174, 2.670208, 2.854345, 2.702724, 2.391875, 
    2.04643,
  3.284592, 3.158846, 2.997234, 2.753203, 2.406346, 2.099216, 1.589801, 
    1.218477, 1.523305, 2.317833, 2.867229, 3.200538, 3.272377, 3.053697, 
    2.719347,
  3.59439, 3.375852, 3.16476, 2.949343, 2.64342, 2.312614, 2.001225, 
    1.788009, 1.935735, 2.459678, 2.927417, 3.267545, 3.367324, 3.309404, 
    3.054943,
  3.633703, 3.561556, 3.306607, 3.124031, 2.919977, 2.581909, 2.2999, 
    2.131229, 2.113906, 2.613807, 2.913512, 3.170758, 3.253057, 3.224634, 
    3.009701,
  3.662924, 3.654692, 3.44018, 3.251019, 3.119098, 2.832411, 2.708303, 
    2.581969, 2.311673, 2.572051, 2.756918, 3.063631, 3.146313, 3.082778, 
    2.880514,
  3.794517, 3.745155, 3.543237, 3.375056, 3.25477, 2.993234, 3.046126, 
    3.148309, 2.69378, 2.597599, 2.565747, 2.942183, 3.119227, 3.094164, 
    2.841695,
  3.960176, 3.83367, 3.64694, 3.466425, 3.337625, 3.125607, 3.277212, 
    3.536569, 3.035135, 2.508945, 2.360167, 2.733297, 3.051332, 3.156456, 
    2.935086,
  3.498902, 2.986935, 1.780671, 1.472756, 1.603001, 1.977785, 2.156056, 
    2.160396, 2.021456, 1.793517, 1.631391, 1.546786, 1.50706, 1.551636, 
    1.672018,
  3.724712, 3.359482, 2.394797, 1.825707, 1.496348, 1.878047, 2.147497, 
    2.258929, 2.190226, 1.999613, 1.819354, 1.739411, 1.711336, 1.658665, 
    1.753168,
  3.946648, 3.690036, 2.920411, 2.22658, 1.465366, 1.525148, 2.093026, 
    2.333557, 2.388777, 2.233015, 2.023976, 1.919064, 1.891768, 1.921329, 
    1.941488,
  4.047876, 3.79924, 3.238379, 2.603445, 1.828426, 1.791251, 1.804091, 
    2.337181, 2.540094, 2.493731, 2.281815, 2.088667, 1.996094, 2.01979, 
    2.039189,
  4.076694, 3.85322, 3.346349, 2.776972, 2.095326, 2.201416, 2.184368, 
    2.053341, 2.365332, 2.777049, 2.65276, 2.373302, 2.207377, 2.111074, 
    2.061503,
  4.205072, 3.924536, 3.423395, 2.937152, 2.324927, 2.263412, 2.339975, 
    2.781718, 2.987675, 3.070634, 2.890739, 2.576121, 2.374906, 2.233407, 
    2.108237,
  4.065059, 3.952965, 3.561502, 3.154026, 2.655923, 2.432075, 2.342172, 
    2.853351, 3.266142, 3.250901, 2.937237, 2.671041, 2.451057, 2.265646, 
    2.042701,
  3.744573, 3.935295, 3.725135, 3.442694, 2.997086, 2.730621, 2.433354, 
    2.848526, 3.327921, 3.309344, 2.914073, 2.683259, 2.432379, 2.160757, 
    1.909375,
  4.049784, 3.874349, 3.881394, 3.763298, 3.370235, 2.965776, 2.620248, 
    2.765836, 3.302165, 3.320935, 2.878342, 2.696459, 2.390613, 2.093171, 
    1.944506,
  4.950273, 4.182684, 3.943411, 3.941289, 3.65343, 3.320408, 2.807671, 
    2.677579, 3.181018, 3.220834, 2.893994, 2.752202, 2.495273, 2.291713, 
    2.238907,
  3.121949, 3.289534, 2.374338, 1.811442, 1.767101, 1.698251, 1.53624, 
    1.460846, 1.456758, 1.450177, 1.481246, 1.558079, 1.641439, 1.714987, 
    1.74812,
  3.377173, 3.544241, 2.817282, 2.113654, 1.812752, 1.755073, 1.604507, 
    1.462948, 1.404616, 1.399307, 1.421201, 1.560357, 1.691079, 1.713117, 
    1.791978,
  3.549693, 3.72425, 3.179663, 2.42826, 1.892353, 1.658906, 1.698474, 
    1.564009, 1.435812, 1.371993, 1.396851, 1.55253, 1.747873, 1.871566, 
    1.924353,
  3.690898, 3.80282, 3.437869, 2.729718, 2.194995, 1.992837, 1.62353, 
    1.61402, 1.481098, 1.398058, 1.391554, 1.5553, 1.806904, 1.93357, 1.993272,
  3.962279, 3.936142, 3.549721, 2.900745, 2.458964, 2.474242, 2.0206, 
    1.473309, 1.300308, 1.451228, 1.456298, 1.624865, 1.859082, 1.961645, 
    1.980752,
  4.113629, 4.002833, 3.604032, 2.9816, 2.543774, 2.706835, 2.544171, 
    2.180973, 1.835645, 1.674973, 1.582888, 1.732738, 1.918124, 1.999372, 
    1.971245,
  4.20523, 4.066583, 3.612828, 2.995519, 2.689019, 2.895671, 2.820703, 
    2.743864, 2.43139, 2.011544, 1.783603, 1.878698, 1.996511, 2.035771, 
    1.988349,
  4.235242, 4.005407, 3.594332, 2.971605, 2.712082, 2.995926, 3.066309, 
    3.089973, 2.845423, 2.463378, 2.061274, 2.051979, 2.092944, 2.094266, 
    1.965887,
  3.978405, 3.998395, 3.509651, 3.003152, 2.792056, 3.035217, 3.210876, 
    3.396326, 3.31057, 2.889519, 2.36881, 2.232107, 2.196302, 2.127816, 
    1.930187,
  3.741729, 3.775847, 3.517568, 3.169472, 2.894895, 3.042743, 3.218366, 
    3.542372, 3.575256, 3.136307, 2.620222, 2.397691, 2.285071, 2.141229, 
    1.945048,
  2.127622, 1.837365, 1.654583, 1.744614, 1.695448, 1.717326, 1.741324, 
    1.766205, 1.794763, 1.80573, 1.862584, 1.983651, 2.014842, 1.987241, 
    1.949545,
  2.419106, 2.191926, 1.972175, 1.934128, 1.672118, 1.661086, 1.653975, 
    1.647455, 1.692044, 1.801283, 1.902269, 2.050317, 2.133486, 2.050418, 
    2.084641,
  2.71611, 2.531603, 2.212805, 2.12225, 1.627883, 1.381736, 1.484702, 
    1.492728, 1.539628, 1.661928, 1.866464, 2.056856, 2.184756, 2.276778, 
    2.311969,
  2.989405, 2.781846, 2.481274, 2.280217, 1.870183, 1.560875, 1.252778, 
    1.369538, 1.366469, 1.50084, 1.766773, 2.043175, 2.233188, 2.365772, 
    2.449116,
  3.294242, 3.014099, 2.633203, 2.413348, 2.113608, 1.973158, 1.622376, 
    1.138513, 1.093043, 1.378584, 1.670694, 2.000529, 2.237009, 2.395895, 
    2.550989,
  3.540985, 3.263879, 2.857458, 2.684299, 2.377542, 2.217084, 2.03537, 
    1.826023, 1.598672, 1.455716, 1.600207, 1.950673, 2.218713, 2.410392, 
    2.609895,
  3.756959, 3.539422, 3.103742, 2.940172, 2.779784, 2.656692, 2.36512, 
    2.161801, 1.905295, 1.595242, 1.561483, 1.869304, 2.148883, 2.344786, 
    2.573555,
  3.910519, 3.713587, 3.353457, 3.133581, 3.028595, 3.006728, 2.865995, 
    2.512108, 2.262485, 1.886724, 1.552791, 1.818411, 2.026071, 2.181938, 
    2.363441,
  4.01757, 4.010929, 3.623053, 3.38509, 3.246238, 3.244989, 3.176155, 
    3.000918, 2.577671, 2.18992, 1.641593, 1.787414, 1.951435, 2.052254, 
    2.165608,
  4.281896, 4.027165, 3.876555, 3.652115, 3.351372, 3.338269, 3.379333, 
    3.269706, 2.970045, 2.355074, 1.779415, 1.822892, 1.918343, 2.00588, 
    2.08139,
  1.667185, 1.766818, 1.663821, 1.675908, 1.573807, 1.600885, 1.738894, 
    2.039551, 2.322076, 2.444556, 2.445686, 2.43994, 2.321203, 2.200185, 
    2.100434,
  2.009794, 2.074583, 1.966324, 1.848928, 1.609919, 1.559807, 1.677613, 
    1.950188, 2.317331, 2.567246, 2.615038, 2.602126, 2.535265, 2.330307, 
    2.288795,
  2.316624, 2.347208, 2.222157, 2.036803, 1.778367, 1.510679, 1.653426, 
    1.909398, 2.286856, 2.604597, 2.754809, 2.774049, 2.71652, 2.653704, 
    2.610008,
  2.516417, 2.515703, 2.37815, 2.192611, 2.055464, 1.983807, 1.647306, 
    1.781565, 2.130215, 2.575575, 2.786146, 2.877316, 2.90252, 2.866826, 
    2.829654,
  2.732226, 2.702835, 2.570869, 2.383247, 2.275909, 2.242463, 2.206604, 
    1.524394, 1.660828, 2.436072, 2.738717, 2.888947, 2.957297, 2.96197, 
    2.914971,
  2.838867, 2.791279, 2.688986, 2.601363, 2.501572, 2.460761, 2.414809, 
    2.304841, 2.061104, 2.373421, 2.639389, 2.808543, 2.884188, 2.910182, 
    2.893063,
  3.319404, 3.142812, 2.971356, 2.939042, 2.934447, 2.830654, 2.632175, 
    2.609819, 2.254394, 2.216393, 2.52135, 2.604022, 2.636028, 2.657279, 
    2.648688,
  4.353325, 4.036014, 3.665583, 3.38899, 3.271721, 3.210565, 3.178779, 
    2.962901, 2.604523, 2.115102, 2.251747, 2.387556, 2.4185, 2.390099, 
    2.369084,
  6.389129, 5.706524, 5.087755, 4.415614, 3.8218, 3.476792, 3.3938, 3.326745, 
    2.984276, 2.117991, 2.018188, 2.207556, 2.23397, 2.237861, 2.229782,
  7.288489, 6.575529, 6.002488, 5.422728, 4.555577, 3.781194, 3.434939, 
    3.391373, 3.228623, 2.193716, 1.87344, 2.012796, 2.116738, 2.16215, 
    2.131247,
  1.400323, 1.730625, 2.117574, 2.291899, 2.275359, 2.287167, 2.495184, 
    2.720048, 2.76547, 2.664253, 2.601047, 2.616827, 2.541899, 2.419134, 
    2.355755,
  1.749776, 2.098265, 2.313213, 2.389693, 2.513746, 2.334982, 2.40832, 
    2.676003, 2.735876, 2.70615, 2.651021, 2.649761, 2.585211, 2.405694, 
    2.460246,
  2.182157, 2.271046, 2.461575, 2.573303, 2.779896, 2.346617, 2.308613, 
    2.595216, 2.712044, 2.648891, 2.611166, 2.574788, 2.51515, 2.490819, 
    2.567189,
  2.467262, 2.526014, 2.617263, 2.774518, 2.887807, 2.894917, 2.137717, 
    2.291146, 2.501173, 2.536559, 2.500491, 2.465774, 2.435802, 2.420916, 
    2.514434,
  2.653947, 2.833338, 2.871559, 2.96455, 3.015277, 3.003153, 2.726584, 
    1.756847, 1.894112, 2.409941, 2.378106, 2.333007, 2.290593, 2.29066, 
    2.387384,
  2.833658, 3.010636, 3.193214, 3.274357, 3.284261, 3.073033, 3.052756, 
    2.432973, 2.228229, 2.311323, 2.275749, 2.23158, 2.19379, 2.193914, 
    2.281785,
  4.129415, 3.730178, 3.508546, 3.498678, 3.653688, 3.534758, 3.159447, 
    2.581563, 2.229589, 2.156673, 2.205199, 2.158719, 2.124457, 2.104147, 
    2.160765,
  6.385473, 5.78515, 5.160148, 4.432234, 4.069162, 3.772116, 3.338543, 
    3.131433, 2.605034, 2.12402, 2.117266, 2.1277, 2.090041, 2.044969, 
    2.060504,
  5.966174, 6.103193, 6.124759, 5.91453, 5.433851, 4.796654, 3.719249, 
    3.506775, 3.341224, 2.373942, 2.050401, 2.089931, 2.053518, 1.971772, 
    1.957863,
  4.528097, 4.744389, 5.038771, 5.685344, 5.91063, 5.635309, 4.553733, 
    3.80936, 3.596003, 2.704048, 2.17428, 2.01981, 2.018018, 1.902067, 
    1.812714,
  1.650702, 2.111407, 2.516941, 2.814054, 2.712037, 2.413544, 2.292126, 
    2.282833, 2.163863, 2.040204, 2.047503, 2.309074, 2.495913, 2.4972, 
    2.409636,
  1.921387, 2.467329, 3.0076, 3.097864, 3.030648, 2.625363, 2.320456, 
    2.195474, 2.076271, 2.017202, 1.996037, 2.186076, 2.473504, 2.49735, 
    2.493755,
  2.165298, 2.451748, 2.838827, 3.180566, 3.396414, 2.653873, 2.393722, 
    2.219075, 2.05845, 1.973924, 1.927918, 2.016995, 2.32938, 2.659257, 
    2.713442,
  2.313118, 2.49394, 2.695608, 3.208403, 3.516371, 3.481467, 2.397811, 
    2.02864, 1.866188, 1.930427, 1.875932, 1.904103, 2.110013, 2.608805, 
    2.817006,
  2.433379, 2.622483, 2.808761, 3.139391, 3.445731, 3.825061, 3.302769, 
    1.763724, 1.466474, 1.876028, 1.912066, 1.877347, 1.910031, 2.342689, 
    2.813297,
  2.504434, 2.709647, 2.914109, 3.165135, 3.475769, 3.71047, 3.632783, 
    2.778735, 2.0938, 1.966562, 1.98662, 1.952827, 1.836271, 1.999652, 
    2.589877,
  2.857234, 2.945949, 3.036823, 3.159348, 3.377784, 3.676866, 3.777973, 
    3.2343, 2.673441, 2.236225, 2.161971, 2.117227, 1.917515, 1.795218, 
    2.161172,
  3.675585, 3.461751, 3.35418, 3.28324, 3.378829, 3.569419, 3.765607, 
    3.603162, 3.355394, 2.92976, 2.635807, 2.40779, 2.124393, 1.845095, 
    1.806859,
  4.632875, 4.226145, 4.097587, 3.927501, 3.772861, 3.810055, 3.95944, 
    3.966561, 3.853273, 3.527953, 3.207003, 2.858323, 2.450976, 2.067674, 
    1.797786,
  5.483633, 5.004962, 4.734599, 4.526692, 4.352557, 4.328135, 4.369364, 
    4.319125, 4.223039, 4.025676, 3.78822, 3.406561, 2.929601, 2.471906, 
    2.061916,
  2.544695, 2.382713, 2.093151, 1.934916, 1.949822, 1.975195, 1.891132, 
    1.798187, 1.733385, 1.738238, 1.884179, 2.169235, 2.432997, 2.54756, 
    2.463691,
  2.540132, 2.50329, 2.344604, 2.217757, 2.148247, 2.130145, 2.113183, 
    1.79924, 1.651479, 1.731298, 1.906205, 2.12488, 2.364062, 2.481788, 
    2.562687,
  2.622039, 2.671159, 2.64706, 2.604091, 2.412178, 2.057935, 2.299196, 
    2.022267, 1.870064, 1.778867, 1.941087, 2.148379, 2.356146, 2.654316, 
    2.755744,
  2.639979, 2.752367, 2.818612, 2.935945, 3.035872, 2.872438, 2.24379, 
    2.444687, 2.228805, 1.985659, 2.068812, 2.291048, 2.514923, 2.699893, 
    2.833959,
  2.653968, 2.778413, 2.875449, 3.060232, 3.350735, 3.605624, 3.455905, 
    2.625127, 2.378925, 2.41919, 2.424757, 2.597986, 2.816967, 2.869673, 
    2.865945,
  2.701621, 2.792488, 2.901178, 3.053065, 3.250175, 3.394952, 3.631588, 
    3.710983, 3.550462, 3.143145, 2.905076, 3.020446, 3.207443, 3.206751, 
    2.979721,
  2.718997, 2.82464, 2.916604, 3.031856, 3.139115, 3.223326, 3.310008, 
    3.477008, 3.691908, 3.684327, 3.516322, 3.499745, 3.569155, 3.549495, 
    3.249436,
  2.742696, 2.863936, 2.954508, 3.039724, 3.141601, 3.21433, 3.305202, 
    3.410219, 3.594052, 3.767052, 3.80311, 3.808882, 3.849303, 3.853233, 
    3.672065,
  2.825693, 2.95649, 3.075451, 3.141229, 3.234274, 3.316412, 3.3949, 
    3.473401, 3.646242, 3.780327, 3.852113, 3.944274, 4.10308, 4.140076, 
    4.11505,
  3.238691, 3.215699, 3.283986, 3.375599, 3.458706, 3.543562, 3.632037, 
    3.779545, 3.907182, 3.93602, 4.045988, 4.189956, 4.387928, 4.533351, 
    4.597218,
  3.344943, 3.549598, 3.30993, 2.960667, 2.132197, 1.746347, 1.678046, 
    1.617644, 1.560811, 1.717795, 2.077971, 2.638738, 3.186612, 3.097048, 
    2.547077,
  3.517906, 3.795904, 3.543648, 2.97864, 2.064389, 1.718651, 1.693641, 
    1.647916, 1.643669, 2.010383, 2.313966, 2.927213, 3.492604, 3.186521, 
    2.517973,
  3.686439, 3.961074, 3.72469, 3.079492, 2.060401, 1.55978, 1.725234, 
    1.725243, 2.24371, 2.388963, 2.615165, 3.189012, 3.780629, 3.678622, 
    2.651867,
  3.696496, 3.933552, 3.758122, 3.215384, 2.340805, 1.763075, 1.625522, 
    2.2677, 2.72212, 2.729613, 2.956568, 3.402737, 3.96039, 4.014263, 2.796983,
  3.588005, 3.781101, 3.653419, 3.260054, 2.620446, 2.259567, 2.06244, 
    2.047233, 2.268015, 3.012784, 3.255661, 3.538774, 3.990668, 4.318762, 
    3.271669,
  3.547033, 3.684081, 3.562818, 3.253729, 2.839025, 2.63721, 2.693283, 
    2.937668, 3.136899, 3.223521, 3.355816, 3.560446, 3.910879, 4.436273, 
    3.984598,
  3.533966, 3.600508, 3.50284, 3.32342, 3.061181, 2.916446, 2.943302, 
    3.211159, 3.319096, 3.392653, 3.390242, 3.532219, 3.811015, 4.349061, 
    4.503071,
  3.492007, 3.512006, 3.420944, 3.32479, 3.201219, 3.108995, 3.115772, 
    3.264912, 3.391344, 3.493871, 3.488697, 3.557603, 3.802853, 4.252605, 
    4.794655,
  3.40289, 3.39347, 3.32475, 3.306649, 3.255496, 3.230092, 3.25013, 3.315263, 
    3.458993, 3.535339, 3.496064, 3.567729, 3.86567, 4.273613, 5.015484,
  3.223151, 3.232614, 3.237096, 3.255456, 3.266817, 3.282911, 3.324101, 
    3.387585, 3.51062, 3.591095, 3.735194, 3.96268, 4.280613, 4.69076, 5.35817,
  3.019217, 2.344692, 1.991827, 1.852636, 1.707218, 1.630126, 1.682741, 
    1.990626, 2.491732, 2.960884, 3.19013, 3.040555, 2.372927, 2.008596, 
    1.928156,
  3.090875, 2.576397, 2.288003, 1.984298, 1.735759, 1.623255, 1.651516, 
    1.921199, 2.452171, 2.994497, 3.312814, 3.467066, 3.061417, 2.40194, 
    2.301049,
  3.294712, 2.962778, 2.747076, 2.329041, 1.858383, 1.488158, 1.595977, 
    1.857437, 2.443778, 2.923589, 3.333726, 3.56449, 3.662759, 3.247829, 
    2.860515,
  3.528604, 3.340685, 3.196438, 2.79246, 2.287841, 1.775267, 1.44147, 
    1.809013, 2.49497, 2.854282, 3.21546, 3.452803, 3.862778, 3.932309, 
    3.431793,
  3.658885, 3.608049, 3.569518, 3.288776, 2.796718, 2.317421, 1.805036, 
    1.562286, 1.913852, 2.771426, 3.106448, 3.282131, 3.743652, 4.171597, 
    4.014177,
  3.706658, 3.782535, 3.830714, 3.726712, 3.233495, 2.769533, 2.381788, 
    2.053228, 2.376018, 2.768091, 3.012554, 3.181931, 3.528994, 4.09493, 
    4.39877,
  3.779833, 3.902972, 4.00761, 4.010237, 3.701541, 3.182784, 2.772092, 
    2.609084, 2.708144, 2.82993, 3.016484, 3.125766, 3.408356, 3.893445, 
    4.465868,
  3.857013, 4.031548, 4.161604, 4.155557, 3.966625, 3.555729, 3.133798, 
    2.867496, 2.78843, 2.892281, 3.061681, 3.20096, 3.384481, 3.770376, 
    4.355263,
  4.010852, 4.115012, 4.219223, 4.210567, 4.09202, 3.831273, 3.478299, 
    3.197492, 3.090057, 3.12581, 3.133659, 3.191939, 3.389931, 3.743971, 
    4.200869,
  4.272057, 4.283057, 4.278655, 4.236792, 4.112764, 3.925345, 3.68045, 
    3.441264, 3.338375, 3.202742, 3.166489, 3.199191, 3.45541, 3.789682, 
    4.153955,
  1.572467, 1.478335, 1.535112, 1.719053, 1.91271, 2.111352, 2.263701, 
    2.408319, 2.511331, 2.595132, 2.727825, 3.294891, 3.690323, 3.295213, 
    2.562439,
  1.801494, 1.670119, 1.692262, 1.69087, 1.777974, 1.942286, 2.159927, 
    2.211745, 2.318739, 2.555285, 2.649358, 3.138438, 3.650645, 3.224768, 
    2.580719,
  2.126593, 1.987249, 1.99431, 1.878712, 1.686792, 1.505153, 1.767306, 
    2.007597, 2.176003, 2.442255, 2.55037, 2.931799, 3.547993, 3.412619, 
    2.697005,
  2.480856, 2.296509, 2.286561, 2.220249, 2.090183, 1.875923, 1.559711, 
    1.75697, 2.085341, 2.373446, 2.448717, 2.722939, 3.408537, 3.454471, 
    2.774662,
  2.80134, 2.600507, 2.568313, 2.540291, 2.532562, 2.473628, 2.348938, 
    1.776901, 1.734953, 2.273446, 2.40919, 2.563774, 3.251082, 3.479078, 
    2.91647,
  3.137358, 2.908484, 2.868037, 2.894375, 2.941865, 3.019201, 3.035542, 
    2.848592, 2.666826, 2.560937, 2.41085, 2.462928, 3.074095, 3.49878, 
    3.113906,
  3.551164, 3.362088, 3.334489, 3.380599, 3.464505, 3.501899, 3.522244, 
    3.484625, 3.33276, 3.034595, 2.724584, 2.474662, 2.927628, 3.516007, 
    3.369787,
  3.959987, 3.831544, 3.794205, 3.773197, 3.835508, 3.881647, 3.851048, 
    3.754623, 3.633971, 3.411661, 3.025142, 2.585619, 2.809241, 3.434248, 
    3.634101,
  4.436715, 4.330461, 4.278201, 4.284812, 4.27276, 4.20963, 4.165701, 
    4.058781, 3.888721, 3.699086, 3.304067, 2.823959, 2.76028, 3.196957, 
    3.744568,
  4.47938, 4.505273, 4.535535, 4.550434, 4.556727, 4.569515, 4.508738, 
    4.442185, 4.308876, 4.054236, 3.723084, 3.128004, 2.800482, 2.947349, 
    3.521004,
  1.659538, 1.926338, 2.059, 2.125743, 2.157456, 2.255749, 2.340507, 
    2.406772, 2.277987, 2.051631, 1.854766, 1.499804, 1.104731, 0.9722319, 
    0.9742713,
  1.935301, 2.046978, 2.121532, 2.062838, 2.110074, 2.201164, 2.499349, 
    2.644014, 2.506173, 2.138796, 1.946563, 1.56009, 1.128179, 0.9450114, 
    0.9851353,
  2.131236, 2.175725, 2.206913, 2.172686, 2.157042, 1.989984, 2.565119, 
    3.037067, 3.018088, 2.359994, 2.050266, 1.641257, 1.172461, 1.02347, 
    1.050219,
  2.324811, 2.333905, 2.386307, 2.444928, 2.543334, 2.747498, 2.581202, 
    3.278915, 3.373021, 2.842326, 2.155782, 1.835577, 1.27096, 1.047083, 
    1.089183,
  2.463434, 2.448563, 2.485214, 2.603874, 2.801177, 3.203521, 3.450718, 
    3.044195, 3.029691, 3.416199, 2.416678, 2.071129, 1.452336, 1.103588, 
    1.158852,
  2.644527, 2.674563, 2.691453, 2.818912, 3.090833, 3.464718, 3.786433, 
    3.962227, 3.995702, 3.873599, 2.708179, 2.348673, 1.770355, 1.217235, 
    1.222013,
  2.7742, 2.897454, 3.071947, 3.287759, 3.572761, 3.914255, 4.104847, 
    4.191792, 4.113323, 4.021512, 3.28511, 2.507272, 2.243791, 1.487079, 
    1.299656,
  2.9603, 3.143952, 3.372414, 3.710886, 4.036468, 4.208531, 4.275872, 
    4.20662, 4.065174, 4.045587, 3.739653, 2.688047, 2.695817, 1.953406, 
    1.457166,
  3.443969, 3.667094, 3.968747, 4.217564, 4.359908, 4.313402, 4.278698, 
    4.254638, 4.137568, 4.07407, 3.982979, 2.949026, 2.79788, 2.651939, 
    1.928271,
  4.229989, 4.377867, 4.493926, 4.532587, 4.455677, 4.401487, 4.440388, 
    4.444228, 4.538065, 4.435203, 4.304012, 3.657137, 2.779077, 2.985966, 
    2.838384,
  2.069746, 2.186058, 2.337677, 2.616, 2.95532, 3.300351, 3.664669, 3.32357, 
    2.213366, 1.367082, 1.00811, 1.05637, 1.189363, 1.309356, 1.423681,
  2.150945, 2.195672, 2.356202, 2.465039, 2.907889, 3.36867, 3.928558, 
    3.837675, 3.033148, 1.923353, 1.23868, 1.089689, 1.227656, 1.311745, 
    1.460508,
  2.295333, 2.287171, 2.306558, 2.565538, 3.043077, 3.274679, 4.003442, 
    4.125255, 3.572496, 2.606322, 1.569763, 1.175244, 1.231937, 1.412657, 
    1.544267,
  2.486362, 2.451311, 2.431497, 2.732278, 3.439203, 3.962591, 3.946958, 
    4.097351, 3.751468, 3.111992, 2.037281, 1.324397, 1.222874, 1.430516, 
    1.587652,
  2.673372, 2.611817, 2.634438, 3.009174, 3.604654, 4.20105, 4.421587, 
    3.488046, 2.985772, 3.241489, 2.475444, 1.464242, 1.237993, 1.445218, 
    1.616581,
  2.887482, 2.870275, 2.954133, 3.377462, 3.742908, 4.240174, 4.37234, 
    4.21369, 3.958184, 3.613152, 2.627354, 1.650447, 1.368713, 1.487003, 
    1.632473,
  3.048421, 3.245897, 3.410056, 3.570213, 3.845242, 4.253043, 4.334596, 
    4.265017, 4.119966, 3.698653, 2.924335, 2.115604, 1.786516, 1.611733, 
    1.638042,
  2.959234, 3.219552, 3.396498, 3.566722, 3.954953, 4.280416, 4.302022, 
    4.258995, 4.064438, 3.899601, 3.470592, 2.740367, 2.314943, 1.83417, 
    1.677846,
  2.83345, 3.079778, 3.339185, 3.696443, 4.12039, 4.264022, 4.324671, 
    4.427054, 4.318248, 4.126709, 3.85012, 3.253455, 2.711325, 2.141707, 
    1.786718,
  2.927206, 3.18546, 3.49436, 3.874859, 4.131302, 4.21236, 4.427234, 
    4.463505, 4.318713, 4.172891, 4.145761, 3.855678, 3.088802, 2.597581, 
    2.096621,
  1.743189, 2.043083, 2.319583, 2.366215, 2.581135, 3.512663, 4.172647, 
    4.029018, 3.708008, 3.367285, 3.037547, 2.46793, 1.995484, 1.732327, 
    1.58159,
  2.020586, 2.171924, 2.385766, 2.385731, 2.715181, 3.480363, 4.058763, 
    3.990699, 3.699764, 3.56498, 3.278614, 2.688831, 2.15384, 1.785104, 
    1.611359,
  2.340162, 2.34533, 2.470915, 2.576958, 2.967976, 3.250968, 3.902441, 
    4.039618, 3.830565, 3.734537, 3.443856, 2.85134, 2.298301, 1.974968, 
    1.72245,
  2.620609, 2.538657, 2.574327, 2.69097, 3.209321, 3.735841, 3.711897, 
    3.758912, 3.676998, 3.88748, 3.616019, 3.001888, 2.481864, 2.067292, 
    1.764706,
  2.781378, 2.80207, 2.806696, 2.925579, 3.34585, 3.795279, 4.060781, 
    3.28882, 3.175838, 3.947906, 3.801807, 3.199254, 2.687743, 2.170277, 
    1.811531,
  2.821498, 2.923802, 3.034391, 3.232369, 3.504504, 3.737009, 3.956388, 
    4.03187, 4.104485, 4.194167, 3.941278, 3.419298, 2.907686, 2.26715, 
    1.850436,
  2.699134, 2.963304, 3.185854, 3.350286, 3.521234, 3.665224, 3.799732, 
    3.983072, 4.187767, 4.236513, 4.016136, 3.567942, 3.072672, 2.363814, 
    1.891818,
  2.638029, 2.866041, 3.096566, 3.300318, 3.41665, 3.550564, 3.684489, 
    3.842133, 4.078042, 4.156939, 3.926365, 3.55564, 3.159752, 2.448157, 
    1.940323,
  2.776414, 2.921826, 3.09517, 3.277068, 3.365396, 3.492792, 3.645785, 
    3.95891, 4.179295, 4.146881, 3.82438, 3.435593, 3.19504, 2.549724, 
    1.998298,
  3.137426, 3.195504, 3.254344, 3.301067, 3.393402, 3.640136, 3.969961, 
    4.239477, 4.441546, 4.228542, 3.760588, 3.245758, 3.18379, 2.744165, 
    2.086249,
  2.088138, 1.931079, 2.018244, 2.173636, 2.163029, 2.100361, 2.152435, 
    2.468494, 2.879695, 3.286702, 3.544952, 3.632874, 3.543287, 3.048601, 
    2.221083,
  2.63659, 2.350502, 2.266014, 2.209863, 2.113672, 2.093099, 2.264324, 
    2.715869, 3.12709, 3.421031, 3.590083, 3.666491, 3.612311, 3.01234, 
    2.155706,
  3.142243, 2.939168, 2.794341, 2.741968, 2.699827, 2.41288, 2.654197, 
    3.059837, 3.295074, 3.407917, 3.560732, 3.680799, 3.661286, 3.178267, 
    2.205401,
  3.218814, 3.095123, 2.976001, 2.921886, 3.010157, 3.098497, 2.895137, 
    3.104508, 3.181508, 3.3421, 3.579237, 3.691583, 3.722761, 3.199862, 
    2.19422,
  3.098976, 3.068238, 3.041893, 3.101082, 3.241229, 3.418489, 3.577298, 
    3.123744, 2.911176, 3.386396, 3.686112, 3.773095, 3.783426, 3.250785, 
    2.241421,
  2.839848, 2.984565, 3.226616, 3.461474, 3.683274, 3.858915, 3.958985, 
    3.97314, 3.951885, 3.994442, 4.035449, 4.035453, 3.914082, 3.28839, 
    2.250171,
  3.319444, 3.671548, 3.944398, 4.196621, 4.358674, 4.4708, 4.491699, 
    4.477716, 4.43236, 4.329222, 4.323081, 4.279749, 4.040996, 3.280462, 
    2.212004,
  4.441336, 4.611253, 4.800241, 4.962861, 5.056736, 5.080181, 4.97655, 
    4.661514, 4.388048, 4.3501, 4.435767, 4.448283, 4.157408, 3.240051, 
    2.167603,
  5.251266, 5.314081, 5.403155, 5.497388, 5.574198, 5.470351, 5.051029, 
    4.45095, 4.240962, 4.333437, 4.473963, 4.529471, 4.201729, 3.155827, 
    2.145133,
  5.453005, 5.56733, 5.755095, 5.918138, 5.908617, 5.534344, 4.702491, 
    4.126965, 4.170285, 4.312754, 4.495556, 4.547011, 4.170025, 3.064012, 
    2.118908,
  1.810007, 1.771371, 1.777444, 1.887495, 1.985746, 2.053648, 2.080755, 
    2.1089, 2.154991, 2.254985, 2.655968, 3.298265, 3.607436, 3.61532, 
    3.272688,
  2.083441, 2.021428, 2.024522, 2.005206, 1.958576, 1.997325, 2.108883, 
    2.275538, 2.543197, 3.026623, 3.664865, 4.159272, 4.168699, 3.826427, 
    3.317219,
  2.525334, 2.485961, 2.520678, 2.561569, 2.547343, 2.242736, 2.570037, 
    3.079482, 3.508201, 3.987773, 4.583456, 4.829535, 4.532962, 4.199662, 
    3.427938,
  3.241634, 2.812129, 2.746476, 2.822899, 2.975441, 3.086775, 2.987109, 
    3.530612, 3.961445, 4.843575, 5.417083, 5.255138, 4.48983, 4.187422, 
    3.281169,
  4.205723, 3.532644, 3.073945, 3.049538, 3.30474, 3.735713, 4.172151, 
    3.806801, 4.041322, 5.507208, 5.779248, 4.920279, 4.23932, 4.122637, 
    3.276824,
  5.362722, 4.586002, 3.93714, 3.688522, 3.856793, 4.3536, 4.783912, 
    5.164809, 5.571721, 5.887417, 5.250687, 4.296909, 4.014673, 4.088217, 
    3.194032,
  6.352824, 5.863862, 5.275298, 4.80044, 4.626497, 4.799838, 5.172287, 
    5.585792, 5.847158, 5.309427, 4.42954, 3.86389, 3.866889, 3.912281, 
    3.032622,
  7.096664, 6.886362, 6.431458, 5.871194, 5.460636, 5.297284, 5.437103, 
    5.653255, 5.322565, 4.639537, 4.072979, 3.702606, 3.867161, 3.690552, 
    2.78564,
  7.808833, 7.603997, 7.235746, 6.654061, 6.074246, 5.719695, 5.651188, 
    5.53459, 5.024933, 4.478083, 3.963429, 3.758563, 3.857259, 3.417336, 
    2.50529,
  8.717179, 8.537355, 8.125257, 7.477561, 6.777167, 6.249618, 5.889047, 
    5.35878, 4.810339, 4.289214, 3.983199, 3.771577, 3.650726, 3.150608, 
    2.281805,
  3.62075, 2.627389, 1.819557, 1.40671, 1.195545, 1.056693, 1.001308, 
    1.025987, 1.100109, 1.171248, 1.308954, 1.574072, 2.172743, 2.908593, 
    3.4383,
  4.934602, 3.779659, 2.566194, 1.75125, 1.357743, 1.193944, 1.135048, 
    1.092285, 1.11132, 1.239864, 1.435422, 1.918838, 2.648563, 3.189314, 
    3.373745,
  6.933646, 5.691297, 4.459338, 3.045791, 1.885109, 1.264775, 1.281833, 
    1.314688, 1.345678, 1.466835, 1.736814, 2.350817, 3.051722, 3.505545, 
    3.114793,
  8.131297, 7.257216, 6.183366, 5.094098, 3.91371, 2.653301, 1.735413, 
    1.615763, 1.664121, 1.787551, 2.132524, 2.743889, 3.350646, 3.492805, 
    2.778164,
  8.658787, 7.914532, 7.230507, 6.436078, 5.541102, 4.608807, 3.658006, 
    2.395279, 1.874094, 2.10771, 2.515413, 3.044676, 3.513877, 3.420542, 
    2.632226,
  8.627933, 7.979042, 7.536982, 7.193607, 6.622987, 5.905724, 5.018671, 
    4.274391, 3.558837, 3.145075, 2.9448, 3.250206, 3.611374, 3.191415, 
    2.408446,
  8.092876, 7.522339, 7.316613, 7.309878, 7.231703, 6.838679, 6.194789, 
    5.482537, 4.760839, 3.987875, 3.466366, 3.462028, 3.59452, 2.964835, 
    2.213465,
  7.257357, 6.616862, 6.520074, 6.724125, 6.933199, 6.995768, 6.715082, 
    6.174625, 5.620133, 4.821074, 4.171319, 3.772216, 3.552155, 2.782374, 
    2.090858,
  5.250083, 4.709209, 5.019265, 5.727783, 6.392821, 6.7709, 6.788949, 
    6.519369, 6.139256, 5.495547, 4.79798, 4.172719, 3.583462, 2.662041, 
    1.948691,
  4.233907, 4.184747, 4.891122, 6.029036, 6.99765, 7.584465, 7.535536, 
    7.074533, 6.533185, 5.950325, 5.238084, 4.496523, 3.583186, 2.592152, 
    1.858629,
  6.440376, 5.209987, 3.654431, 2.363938, 2.163949, 1.868531, 1.505754, 
    1.196659, 1.059922, 1.025839, 1.120063, 1.188159, 1.116553, 1.121856, 
    1.417928,
  7.147505, 6.306877, 4.881848, 2.882809, 2.066034, 1.89104, 1.658849, 
    1.27614, 1.038181, 0.9738326, 1.010497, 1.06569, 1.064211, 1.141526, 
    1.476147,
  7.724419, 7.112007, 6.075565, 4.16822, 2.27239, 1.682316, 1.710513, 
    1.483274, 1.189811, 1.013457, 0.9929052, 1.036182, 1.093556, 1.279996, 
    1.620386,
  8.571683, 7.631632, 6.821801, 5.532739, 3.318877, 2.078441, 1.699214, 
    1.569579, 1.365609, 1.174747, 1.072211, 1.062708, 1.136315, 1.382492, 
    1.674603,
  9.125089, 8.143505, 7.146725, 6.254291, 4.660822, 3.079095, 2.311915, 
    1.549772, 1.262933, 1.431035, 1.402375, 1.31234, 1.305473, 1.528858, 
    1.72094,
  7.410616, 7.985404, 7.154473, 6.441028, 5.601406, 4.279726, 3.344156, 
    2.662282, 2.249014, 2.227301, 2.029333, 1.725752, 1.525777, 1.699968, 
    1.775673,
  5.78, 6.857364, 6.71341, 6.341802, 5.844105, 5.27246, 4.441796, 3.842979, 
    3.487399, 3.108819, 2.901951, 2.465843, 1.852441, 1.875592, 1.795699,
  4.708716, 5.450994, 6.263652, 6.385596, 6.132143, 5.892812, 5.517201, 
    4.967257, 4.423421, 3.977951, 3.716815, 3.242349, 2.285748, 2.044538, 
    1.82212,
  3.824823, 4.257717, 4.749404, 5.28217, 5.494783, 5.573618, 5.671115, 
    5.630496, 5.380859, 4.908406, 4.451158, 3.951508, 2.803354, 2.233681, 
    1.860859,
  3.069049, 3.207719, 3.392486, 3.832226, 4.382112, 4.895625, 5.275731, 
    5.497499, 5.692514, 5.55476, 5.130406, 4.588766, 3.392591, 2.445721, 
    1.919528,
  4.412238, 3.740005, 3.209656, 2.660863, 2.402913, 2.15349, 1.971351, 
    1.794467, 1.663426, 1.524412, 1.549342, 1.522856, 1.360313, 1.214811, 
    1.304572,
  4.877134, 4.10305, 3.484071, 2.758187, 2.407928, 2.206834, 2.033737, 
    1.831096, 1.669707, 1.533388, 1.543528, 1.517915, 1.317795, 1.106708, 
    1.202418,
  5.449555, 4.637691, 3.879401, 2.923632, 2.433972, 2.011188, 2.040609, 
    1.917216, 1.76336, 1.549862, 1.518135, 1.478857, 1.274651, 1.120759, 
    1.150201,
  5.944845, 5.154608, 4.284942, 3.302493, 2.659743, 2.234712, 1.841524, 
    1.872473, 1.78862, 1.579582, 1.462641, 1.431241, 1.263045, 1.122434, 
    1.089308,
  6.249093, 5.53708, 4.675217, 3.774558, 2.959873, 2.589957, 2.13547, 
    1.566573, 1.455149, 1.574658, 1.460874, 1.380418, 1.311042, 1.176711, 
    1.105558,
  6.296103, 5.682518, 4.933122, 4.218417, 3.353117, 2.868008, 2.552957, 
    2.069702, 1.780105, 1.686021, 1.529954, 1.388436, 1.346424, 1.272605, 
    1.161197,
  6.163689, 5.875724, 5.246302, 4.648065, 3.866446, 3.191501, 2.844862, 
    2.636497, 2.372206, 1.947912, 1.677673, 1.476009, 1.40439, 1.392125, 
    1.237159,
  5.793097, 5.742467, 5.379933, 4.948008, 4.347842, 3.749384, 3.239897, 
    2.907566, 2.689488, 2.272583, 1.910042, 1.678763, 1.520242, 1.493484, 
    1.318089,
  5.2442, 5.539894, 5.485685, 5.21886, 4.713498, 4.221811, 3.72884, 3.338206, 
    2.991336, 2.637231, 2.227404, 1.939901, 1.714996, 1.615069, 1.391972,
  3.88668, 4.493695, 4.87051, 5.100056, 4.979118, 4.705266, 4.316068, 
    3.930587, 3.530564, 3.050763, 2.564792, 2.17856, 1.888284, 1.743941, 
    1.47067,
  2.62174, 1.904145, 1.553918, 1.421419, 1.350087, 1.339221, 1.372733, 
    1.383332, 1.466703, 1.489291, 1.543062, 1.616749, 1.647114, 1.635991, 
    1.641872,
  2.394923, 1.897759, 1.631556, 1.444683, 1.368794, 1.381498, 1.398379, 
    1.417192, 1.478695, 1.519621, 1.545165, 1.593839, 1.597027, 1.520707, 
    1.546144,
  2.517398, 2.139463, 1.858999, 1.548776, 1.40435, 1.254353, 1.413326, 
    1.475958, 1.524322, 1.543446, 1.529347, 1.509332, 1.522179, 1.519753, 
    1.508405,
  2.855246, 2.536198, 2.228464, 1.880143, 1.665743, 1.380531, 1.264563, 
    1.436219, 1.487389, 1.509807, 1.487341, 1.42065, 1.405261, 1.419191, 
    1.451574,
  3.256002, 2.964213, 2.634629, 2.279908, 2.021703, 1.704909, 1.430511, 
    1.142293, 1.161278, 1.449985, 1.44934, 1.373058, 1.306249, 1.293228, 
    1.34505,
  3.737888, 3.403799, 3.008659, 2.64439, 2.344338, 2.035483, 1.80472, 
    1.464339, 1.336571, 1.438024, 1.424567, 1.390896, 1.308924, 1.232524, 
    1.237579,
  4.206481, 3.83894, 3.336025, 2.954654, 2.651467, 2.334179, 2.101954, 
    1.911662, 1.72025, 1.512917, 1.425177, 1.440259, 1.423664, 1.363987, 
    1.24764,
  4.677312, 4.199065, 3.615238, 3.216698, 2.911359, 2.623705, 2.36366, 
    2.195692, 1.985324, 1.610419, 1.458822, 1.459924, 1.49424, 1.497004, 
    1.403181,
  5.054821, 4.518651, 3.921464, 3.465204, 3.135049, 2.875937, 2.660493, 
    2.485684, 2.284491, 1.809362, 1.5623, 1.497497, 1.490348, 1.522593, 
    1.515608,
  5.393035, 4.846113, 4.244586, 3.74104, 3.319893, 3.092509, 2.903841, 
    2.745993, 2.529319, 2.146438, 1.816353, 1.641841, 1.560946, 1.562144, 
    1.581211,
  3.113069, 2.573945, 1.778866, 1.520357, 1.474479, 1.546514, 1.68935, 
    1.796004, 1.914352, 2.00835, 2.127013, 2.272918, 2.393567, 2.537, 2.673486,
  3.062209, 2.390116, 1.717509, 1.466933, 1.434307, 1.533392, 1.682094, 
    1.753618, 1.833546, 1.964482, 2.081407, 2.258039, 2.443284, 2.556559, 
    2.802029,
  2.971888, 2.226848, 1.73501, 1.445203, 1.441334, 1.43084, 1.669618, 
    1.720564, 1.772276, 1.868136, 1.999686, 2.170398, 2.384262, 2.630475, 
    2.889993,
  2.811818, 2.23028, 1.862785, 1.608185, 1.650915, 1.597014, 1.552132, 
    1.654427, 1.665504, 1.75419, 1.914583, 2.114699, 2.374714, 2.69032, 
    3.040377,
  2.708483, 2.280126, 1.999163, 1.857118, 1.888977, 1.886575, 1.763466, 
    1.368806, 1.330699, 1.635476, 1.790344, 2.02651, 2.342856, 2.715444, 
    3.177701,
  2.589547, 2.301372, 2.145853, 2.065375, 2.10512, 2.14135, 2.070087, 
    1.728367, 1.559289, 1.55532, 1.63575, 1.897307, 2.270955, 2.710949, 
    3.245146,
  2.49027, 2.29957, 2.220927, 2.254376, 2.319673, 2.334724, 2.267373, 
    2.037791, 1.790028, 1.535218, 1.524019, 1.759559, 2.152474, 2.626073, 
    3.198037,
  2.534882, 2.434395, 2.364644, 2.431943, 2.478258, 2.480786, 2.365846, 
    2.107312, 1.73868, 1.47822, 1.493531, 1.639947, 1.993599, 2.509829, 
    3.118617,
  2.671109, 2.567976, 2.556794, 2.597299, 2.619664, 2.556811, 2.400748, 
    2.172484, 1.752756, 1.398624, 1.43779, 1.553589, 1.850268, 2.368828, 
    3.018521,
  2.8392, 2.754788, 2.743848, 2.732239, 2.676175, 2.547374, 2.347479, 
    2.095195, 1.581665, 1.331488, 1.446702, 1.561891, 1.768026, 2.196926, 
    2.842606,
  2.191988, 1.826762, 1.899053, 2.068522, 2.215396, 2.365858, 2.513344, 
    2.643212, 2.700854, 2.670622, 2.710514, 2.777165, 2.844355, 2.933959, 
    2.974912,
  2.448979, 1.994811, 2.019738, 2.114648, 2.285291, 2.463037, 2.690722, 
    2.875419, 2.994828, 3.101283, 3.175944, 3.263387, 3.350589, 3.375391, 
    3.429675,
  2.759189, 2.161852, 2.139642, 2.153956, 2.333302, 2.357358, 2.762495, 
    3.046543, 3.277072, 3.454927, 3.595194, 3.696987, 3.779251, 3.871939, 
    3.889314,
  3.055787, 2.447312, 2.372242, 2.376945, 2.589208, 2.612461, 2.699042, 
    3.246815, 3.526274, 3.759005, 3.990922, 4.146934, 4.271425, 4.371921, 
    4.331103,
  3.273289, 2.672632, 2.574904, 2.632137, 2.760605, 2.842844, 2.959164, 
    2.766469, 3.092453, 3.851897, 4.148805, 4.405353, 4.570686, 4.693851, 
    4.610757,
  3.438453, 2.871588, 2.701896, 2.722982, 2.798972, 2.858279, 2.989393, 
    3.099806, 3.362558, 3.741676, 4.126576, 4.462887, 4.690965, 4.831612, 
    4.80708,
  3.587149, 3.054321, 2.822703, 2.750813, 2.797496, 2.842658, 2.886015, 
    2.972376, 3.125406, 3.410263, 3.859645, 4.301685, 4.616182, 4.81215, 
    4.900963,
  3.666447, 3.172917, 2.921077, 2.784414, 2.726333, 2.699943, 2.67983, 
    2.62657, 2.610293, 2.855208, 3.339759, 3.864261, 4.305709, 4.622119, 
    4.843228,
  3.65828, 3.23251, 3.018371, 2.878811, 2.734227, 2.596246, 2.450141, 
    2.331565, 2.277222, 2.41829, 2.776479, 3.20095, 3.653706, 4.056886, 
    4.398104,
  3.637316, 3.308014, 3.123933, 2.969293, 2.799484, 2.543613, 2.280192, 
    2.105198, 1.999023, 2.277735, 2.508298, 2.681149, 2.983137, 3.259125, 
    3.541384,
  2.359887, 2.504012, 2.502416, 2.394704, 2.313561, 2.280273, 2.262632, 
    2.285653, 2.361228, 2.440593, 2.632575, 2.901278, 3.200481, 3.544931, 
    3.898865,
  2.614945, 2.707106, 2.69048, 2.610825, 2.579733, 2.557548, 2.596598, 
    2.622408, 2.635077, 2.669734, 2.767966, 3.00386, 3.322792, 3.568811, 
    3.976249,
  2.903183, 2.957365, 3.086139, 3.073945, 3.136021, 2.986397, 3.14986, 
    3.038851, 3.019254, 3.030494, 3.051923, 3.170428, 3.429387, 3.766691, 
    4.046581,
  3.229138, 3.497204, 3.705619, 3.745124, 3.841548, 3.755402, 3.426568, 
    3.483742, 3.367476, 3.267588, 3.26152, 3.325668, 3.517068, 3.79463, 
    4.075505,
  3.509341, 3.796072, 4.064156, 4.230657, 4.238424, 4.211638, 4.112155, 
    3.409219, 3.185481, 3.560854, 3.513974, 3.521667, 3.666832, 3.884469, 
    4.114587,
  3.678489, 3.99477, 4.24223, 4.435629, 4.481044, 4.419476, 4.32578, 
    4.158386, 3.940531, 3.863191, 3.76415, 3.716614, 3.760212, 3.886371, 
    4.068177,
  3.864173, 4.135283, 4.277676, 4.402246, 4.459279, 4.476558, 4.401984, 
    4.269484, 4.110611, 3.969502, 3.885567, 3.807304, 3.725362, 3.7919, 
    4.012993,
  3.981368, 4.092041, 4.157434, 4.235077, 4.258143, 4.283865, 4.235883, 
    4.127958, 3.996569, 3.992168, 3.958865, 3.888633, 3.860662, 3.975408, 
    4.254228,
  4.062729, 4.035809, 3.971967, 3.912183, 3.896892, 3.902715, 3.903088, 
    3.835229, 3.786329, 3.837748, 3.920385, 3.989186, 4.066322, 4.121011, 
    4.10623,
  4.106324, 3.920707, 3.704149, 3.477287, 3.349727, 3.35156, 3.417311, 
    3.458808, 3.446293, 3.518598, 3.579972, 3.696788, 3.75523, 3.590346, 
    3.207673,
  2.044543, 1.957575, 1.983227, 2.22317, 2.476595, 2.737609, 2.970032, 
    3.17518, 3.361462, 3.491801, 3.711186, 4.039424, 4.209085, 4.203324, 
    4.013913,
  2.2227, 2.111456, 2.156163, 2.353408, 2.570585, 2.828642, 3.097358, 
    3.397517, 3.641807, 3.908127, 4.187582, 4.343782, 4.328886, 4.00631, 
    3.710009,
  2.533373, 2.360219, 2.423017, 2.468443, 2.640736, 2.737558, 3.180426, 
    3.438767, 3.808549, 4.134095, 4.350921, 4.432306, 4.337733, 4.067686, 
    3.692737,
  3.06098, 2.92524, 2.88373, 2.788712, 2.893011, 2.990839, 3.054457, 
    3.589128, 3.876258, 4.125386, 4.364372, 4.38256, 4.267578, 4.009261, 
    3.620907,
  3.596164, 3.444573, 3.340592, 3.25385, 3.271147, 3.302064, 3.402672, 
    3.16615, 3.344218, 4.123346, 4.287518, 4.313176, 4.200467, 3.90182, 
    3.471612,
  4.123393, 3.983253, 3.869571, 3.679045, 3.597305, 3.528507, 3.57091, 
    3.62204, 3.781383, 4.110532, 4.208237, 4.230185, 4.054082, 3.716081, 
    3.262857,
  4.579695, 4.524399, 4.265182, 4.029646, 3.926513, 3.76781, 3.658028, 
    3.723582, 3.875702, 4.071033, 4.188256, 4.122888, 3.869286, 3.521679, 
    3.046368,
  4.886582, 4.74644, 4.544802, 4.294386, 4.114523, 3.938783, 3.798494, 
    3.793788, 3.778435, 4.046427, 4.160519, 4.027031, 3.780926, 3.414341, 
    2.850062,
  4.929243, 4.666463, 4.504583, 4.373504, 4.252604, 4.061386, 3.860741, 
    3.798781, 3.770943, 4.040143, 4.147546, 4.010513, 3.692923, 3.174815, 
    2.40778,
  4.780481, 4.482925, 4.335034, 4.26517, 4.25612, 4.103128, 3.885878, 
    3.745654, 3.693519, 3.950914, 4.107846, 3.989113, 3.453816, 2.570478, 
    2.065439,
  1.795863, 1.809474, 2.057577, 2.362318, 2.544184, 2.655875, 2.730718, 
    2.844359, 3.073253, 3.228063, 3.324944, 3.22471, 2.890492, 2.504372, 
    2.100505,
  1.92502, 2.04675, 2.381491, 2.550523, 2.661743, 2.707604, 2.750143, 
    2.896303, 3.160999, 3.378475, 3.348994, 2.966593, 2.489326, 1.958825, 
    1.665201,
  2.272502, 2.548461, 2.791082, 2.770571, 2.759079, 2.530784, 2.745615, 
    2.945914, 3.301949, 3.550724, 3.249011, 2.705346, 2.225218, 1.860501, 
    1.636082,
  2.810586, 3.114202, 3.203971, 3.105223, 3.021137, 2.867502, 2.611616, 
    3.061007, 3.546649, 3.540617, 3.071275, 2.466549, 2.067045, 1.805348, 
    1.684721,
  3.208054, 3.398233, 3.471903, 3.495023, 3.413263, 3.229917, 3.159601, 
    2.950795, 3.27203, 3.481967, 2.857691, 2.330456, 1.987701, 1.771908, 
    1.716261,
  3.448737, 3.566477, 3.708815, 3.819722, 3.771587, 3.609395, 3.582074, 
    3.786345, 3.891832, 3.453059, 2.738164, 2.271358, 1.91809, 1.752014, 
    1.699519,
  3.729513, 3.785554, 3.965466, 4.085588, 4.059296, 3.921046, 3.871627, 
    4.105748, 4.054372, 3.402323, 2.703245, 2.231226, 1.8869, 1.729016, 
    1.651031,
  4.043009, 3.975061, 4.048615, 4.195384, 4.191502, 4.131752, 4.165029, 
    4.30806, 4.01036, 3.388463, 2.704994, 2.22035, 1.894005, 1.703917, 1.60974,
  4.35857, 4.246112, 4.18021, 4.236284, 4.280087, 4.256407, 4.282763, 
    4.298241, 3.996482, 3.43891, 2.751675, 2.256824, 1.924949, 1.68248, 
    1.594877,
  4.636502, 4.447911, 4.261693, 4.19131, 4.217913, 4.267322, 4.2483, 
    4.183838, 3.922422, 3.529042, 2.89066, 2.361338, 2.020228, 1.731121, 
    1.627735,
  1.708901, 1.841151, 2.20236, 2.532205, 2.750969, 2.948871, 3.026086, 
    2.859594, 2.647577, 2.422371, 2.320961, 2.227055, 2.235485, 2.376145, 
    2.280338,
  1.70368, 1.785209, 2.069283, 2.506341, 2.78024, 2.873608, 2.854272, 
    2.572001, 2.345531, 2.337991, 2.347736, 2.258847, 2.229739, 2.104263, 
    1.883625,
  2.006398, 1.963049, 2.169999, 2.595361, 2.840645, 2.70643, 2.7299, 
    2.298256, 2.123632, 2.249924, 2.325992, 2.224176, 2.116202, 1.987138, 
    1.715312,
  2.334712, 2.31408, 2.484935, 2.75514, 3.029771, 2.998735, 2.465986, 
    2.23834, 1.973184, 2.099942, 2.224004, 2.144445, 1.993487, 1.846117, 
    1.706988,
  2.648652, 2.706021, 2.796489, 2.92071, 3.189815, 3.318612, 2.87088, 
    1.940632, 1.635347, 1.952366, 2.108749, 2.050967, 1.923512, 1.824251, 
    1.821847,
  2.9685, 3.036604, 3.010468, 3.05867, 3.215269, 3.475396, 3.270153, 2.64847, 
    2.03051, 1.900644, 1.990465, 1.961917, 1.894206, 1.869609, 1.942624,
  3.254988, 3.396111, 3.348846, 3.312761, 3.377921, 3.502052, 3.571567, 
    2.950338, 2.245998, 1.84082, 1.875382, 1.880094, 1.861324, 1.901525, 
    2.030507,
  3.558786, 3.743093, 3.750889, 3.653094, 3.546272, 3.507695, 3.657946, 
    3.358208, 2.41171, 1.851759, 1.790794, 1.800915, 1.83594, 1.912639, 
    2.062059,
  3.863669, 4.078916, 4.156399, 3.999318, 3.782154, 3.570141, 3.682093, 
    3.783226, 2.772586, 1.950381, 1.765391, 1.758352, 1.815913, 1.903358, 
    2.038621,
  4.176558, 4.340549, 4.42201, 4.27941, 3.99251, 3.646909, 3.647321, 4.01444, 
    3.237811, 2.229167, 1.801137, 1.740336, 1.791608, 1.875159, 1.979812,
  1.81217, 1.917431, 2.451449, 2.720746, 2.688049, 2.568426, 2.282227, 
    1.933945, 1.769931, 1.787897, 1.904285, 2.037081, 2.093211, 2.071906, 
    2.000934,
  1.836148, 1.761678, 2.198472, 2.763445, 2.716581, 2.451586, 2.339042, 
    2.118356, 1.879959, 1.822872, 1.840998, 1.918585, 2.056974, 2.041833, 
    2.033856,
  2.195479, 1.948328, 2.128477, 2.711756, 2.971925, 2.422772, 2.123052, 
    2.169327, 2.048953, 1.863493, 1.790606, 1.78775, 1.987126, 2.199979, 
    2.126342,
  2.694539, 2.348447, 2.317129, 2.646713, 3.332891, 3.161383, 2.083535, 
    2.082241, 2.152858, 1.989617, 1.788708, 1.675817, 1.880498, 2.1927, 
    2.144601,
  3.116824, 2.687385, 2.570835, 2.692968, 3.156504, 3.963407, 3.059973, 
    1.694465, 1.829245, 2.142623, 1.935464, 1.667259, 1.758675, 2.141065, 
    2.159799,
  3.530999, 3.048202, 2.799717, 2.794606, 3.061367, 3.712661, 3.804441, 
    2.798527, 2.251482, 2.38623, 2.17015, 1.820625, 1.748912, 2.014978, 
    2.103356,
  3.812478, 3.33182, 3.04734, 2.975907, 3.081399, 3.435118, 3.902744, 
    3.520446, 2.568064, 2.470553, 2.403711, 2.09003, 1.837254, 1.880285, 
    2.000426,
  3.968668, 3.539329, 3.262656, 3.184007, 3.204937, 3.383394, 3.744761, 
    3.750725, 2.910728, 2.468565, 2.514713, 2.340102, 1.978451, 1.862157, 
    1.879731,
  4.046474, 3.690166, 3.472984, 3.423055, 3.438361, 3.514033, 3.753606, 
    3.962806, 3.334584, 2.633783, 2.488669, 2.447289, 2.182769, 1.910924, 
    1.829645,
  4.097671, 3.79458, 3.711806, 3.678072, 3.704421, 3.734061, 3.854322, 
    4.051369, 3.556877, 2.745482, 2.378078, 2.376276, 2.276489, 2.065119, 
    1.878335,
  3.683974, 3.102919, 2.632848, 2.15988, 1.794443, 1.613935, 1.646164, 
    1.813704, 1.89833, 1.898086, 2.058512, 2.112047, 1.937326, 1.844285, 
    1.791181,
  3.810511, 3.23566, 2.747777, 2.344372, 1.905726, 1.644973, 1.591349, 
    1.696604, 1.820936, 1.873244, 2.051778, 2.14572, 2.003392, 1.847714, 
    1.828867,
  4.126482, 3.481237, 2.916723, 2.475009, 2.049285, 1.603498, 1.58595, 
    1.608013, 1.72711, 1.863143, 2.019712, 2.175366, 2.101512, 2.023772, 
    1.943839,
  4.573232, 3.907857, 3.263579, 2.72409, 2.270575, 1.8855, 1.560694, 
    1.571041, 1.636831, 1.787331, 1.977836, 2.135609, 2.128502, 2.093156, 
    2.02448,
  4.796628, 4.34809, 3.667565, 3.082837, 2.6135, 2.343427, 2.038941, 1.47291, 
    1.37986, 1.630795, 1.843917, 2.039829, 2.113011, 2.12619, 2.125097,
  4.798264, 4.591825, 4.00628, 3.387022, 2.892824, 2.656549, 2.55917, 
    2.215196, 1.996694, 1.807556, 1.744323, 1.879337, 1.991892, 2.076526, 
    2.192587,
  4.79836, 4.714086, 4.285177, 3.646173, 3.128266, 2.858093, 2.875197, 
    2.857787, 2.699096, 2.236449, 1.870838, 1.791697, 1.83249, 1.911808, 
    2.073739,
  4.827458, 4.78299, 4.445781, 3.876532, 3.329238, 2.987574, 2.990537, 
    3.09142, 3.103477, 2.862835, 2.363072, 1.925096, 1.783684, 1.75446, 
    1.843543,
  4.820624, 4.796874, 4.571938, 4.112782, 3.516187, 3.141464, 3.101474, 
    3.196136, 3.372639, 3.412113, 3.085963, 2.504677, 2.019198, 1.772254, 
    1.707541,
  4.848789, 4.838666, 4.688388, 4.351267, 3.777157, 3.353229, 3.224044, 
    3.274628, 3.414433, 3.560075, 3.503486, 3.133216, 2.677624, 2.187687, 
    1.818885,
  4.521499, 4.161002, 3.634007, 3.059983, 2.332924, 1.74568, 1.739771, 
    1.953121, 1.984333, 1.961195, 1.845775, 1.69349, 1.55863, 1.469424, 
    1.433405,
  4.869389, 4.344817, 3.754072, 3.139951, 2.410112, 1.74234, 1.722994, 
    1.917294, 1.953777, 1.970895, 1.898541, 1.736451, 1.604598, 1.502782, 
    1.495162,
  5.302622, 4.731591, 3.899826, 3.253905, 2.573526, 1.655567, 1.664548, 
    1.871838, 1.941015, 1.934103, 1.928503, 1.809732, 1.68865, 1.641205, 
    1.589921,
  5.475699, 5.171091, 4.243711, 3.436619, 2.848589, 1.86778, 1.511695, 
    1.7793, 1.914742, 1.904049, 1.908912, 1.887886, 1.78405, 1.717166, 1.65774,
  5.483415, 5.412207, 4.598015, 3.695566, 3.140708, 2.176226, 1.693837, 
    1.492962, 1.534028, 1.850465, 1.876614, 1.920603, 1.877669, 1.807349, 
    1.744478,
  5.426174, 5.41278, 4.904999, 3.963918, 3.453565, 2.580997, 1.941061, 
    1.771871, 1.800364, 1.871822, 1.822204, 1.911439, 1.943587, 1.898142, 
    1.829546,
  5.266388, 5.313758, 5.055744, 4.217366, 3.680512, 2.938678, 2.167306, 
    1.966074, 1.915738, 1.854085, 1.778799, 1.861763, 1.953224, 1.957927, 
    1.923783,
  5.117031, 5.200859, 5.037066, 4.409512, 3.79661, 3.216942, 2.469012, 
    2.151118, 1.945192, 1.813959, 1.743157, 1.762846, 1.897739, 1.954112, 
    1.957308,
  4.841054, 5.036423, 4.950941, 4.556508, 3.965998, 3.33691, 2.674224, 
    2.325751, 2.08572, 1.864268, 1.752754, 1.697472, 1.79733, 1.877996, 
    1.910684,
  4.579772, 4.897096, 4.913361, 4.655373, 4.134663, 3.448898, 2.803189, 
    2.474163, 2.156616, 1.930022, 1.848443, 1.77674, 1.763441, 1.821856, 
    1.853835,
  4.525552, 4.784342, 4.882761, 4.402286, 3.589037, 2.99851, 2.293939, 
    1.880058, 1.793973, 1.782416, 1.737706, 1.613153, 1.469524, 1.399533, 
    1.410896,
  4.7949, 5.092517, 5.107729, 4.446153, 3.490238, 2.901319, 2.136222, 
    1.78705, 1.765597, 1.804777, 1.728259, 1.589132, 1.441625, 1.329489, 
    1.361419,
  4.930585, 5.297724, 5.270796, 4.446949, 3.527709, 2.737555, 2.033285, 
    1.713185, 1.736373, 1.77534, 1.706128, 1.559537, 1.420386, 1.382237, 
    1.37601,
  5.068439, 5.368017, 5.45251, 4.599356, 3.636243, 2.985393, 1.850673, 
    1.637684, 1.717747, 1.726881, 1.6519, 1.528418, 1.422935, 1.395663, 
    1.383251,
  5.16363, 5.275987, 5.455807, 4.799193, 3.833809, 3.105321, 2.084588, 
    1.409562, 1.435982, 1.725556, 1.640155, 1.528949, 1.461347, 1.438922, 
    1.427299,
  5.210386, 5.08974, 5.363454, 4.958488, 4.047402, 3.331952, 2.334267, 
    1.724945, 1.761728, 1.802562, 1.643741, 1.553893, 1.502762, 1.500014, 
    1.480285,
  5.059486, 4.883413, 5.178283, 5.067508, 4.177773, 3.544818, 2.497801, 
    1.876903, 1.866493, 1.832354, 1.693796, 1.593014, 1.550416, 1.555725, 
    1.540412,
  4.451146, 4.540268, 5.004434, 5.082018, 4.235119, 3.581556, 2.671959, 
    1.988452, 1.889741, 1.842604, 1.725403, 1.64526, 1.613097, 1.611174, 
    1.595932,
  4.136501, 4.363962, 4.907134, 5.083199, 4.273622, 3.546145, 2.669537, 
    2.149611, 1.930629, 1.858824, 1.751614, 1.708134, 1.691912, 1.681397, 
    1.660811,
  4.131753, 4.538002, 5.087013, 5.064405, 4.194277, 3.513819, 2.697013, 
    2.220173, 1.925554, 1.856421, 1.774122, 1.743747, 1.754425, 1.755487, 
    1.745547,
  4.64857, 4.378712, 4.207864, 4.107648, 4.07368, 3.847112, 3.515404, 
    3.109461, 2.552317, 2.036128, 1.774069, 1.643846, 1.58716, 1.543659, 
    1.558736,
  4.981187, 4.675282, 4.418983, 4.289014, 4.030888, 3.663199, 3.299248, 
    2.908719, 2.409459, 2.000656, 1.794865, 1.682178, 1.617772, 1.49245, 
    1.488022,
  5.403461, 5.144409, 4.779935, 4.459298, 4.036578, 3.267812, 3.05035, 
    2.604001, 2.174192, 1.884901, 1.785224, 1.709307, 1.626632, 1.556001, 
    1.489345,
  5.57177, 5.361402, 5.116442, 4.800616, 4.221442, 3.582551, 2.887313, 
    2.528821, 2.123183, 1.807415, 1.731462, 1.687942, 1.6137, 1.517795, 
    1.457599,
  5.789573, 5.688546, 5.448214, 5.12655, 4.472645, 3.729465, 3.223058, 
    2.317985, 1.812979, 1.753551, 1.697455, 1.652045, 1.579672, 1.496659, 
    1.43394,
  5.659152, 5.746325, 5.600898, 5.344661, 4.723233, 3.939357, 3.366598, 
    2.667461, 2.054586, 1.762027, 1.660935, 1.62638, 1.535231, 1.462505, 
    1.40495,
  4.786129, 5.329621, 5.490013, 5.337231, 4.803764, 4.051486, 3.497148, 
    2.668058, 2.038986, 1.730512, 1.655946, 1.593033, 1.49107, 1.424629, 
    1.384998,
  4.580173, 5.053392, 5.305294, 5.128204, 4.681612, 4.042532, 3.496279, 
    2.575389, 1.875947, 1.681964, 1.629615, 1.534323, 1.4426, 1.393473, 
    1.372195,
  4.268027, 4.634512, 4.836019, 4.851488, 4.480917, 3.890699, 3.260732, 
    2.379282, 1.747218, 1.645434, 1.582384, 1.472643, 1.401025, 1.372492, 
    1.369777,
  4.23612, 4.479296, 4.678986, 4.719479, 4.210669, 3.597051, 2.849382, 
    2.016826, 1.648708, 1.618528, 1.541021, 1.436307, 1.393162, 1.382883, 
    1.383362,
  5.528044, 5.245844, 5.028286, 4.758188, 4.469923, 4.212589, 4.030357, 
    3.843134, 3.599078, 3.24798, 2.881789, 2.390356, 1.988232, 1.691985, 
    1.557335,
  5.740099, 5.43191, 5.062346, 4.718165, 4.312395, 4.019938, 3.85326, 
    3.67785, 3.466588, 3.171166, 2.82316, 2.357501, 1.985679, 1.596596, 
    1.492664,
  5.752593, 5.583603, 5.215931, 4.753405, 4.265551, 3.603693, 3.631934, 
    3.359938, 3.183552, 2.978954, 2.695652, 2.289227, 1.915538, 1.657595, 
    1.48307,
  5.372627, 5.319482, 5.205024, 4.814943, 4.277617, 3.79941, 3.113296, 
    3.079044, 2.973603, 2.731019, 2.525446, 2.180466, 1.827488, 1.617604, 
    1.440836,
  5.098987, 5.22093, 5.089585, 4.833339, 4.279698, 3.727194, 3.327636, 
    2.660903, 2.55483, 2.644753, 2.414691, 2.102489, 1.768028, 1.604325, 
    1.414223,
  4.713169, 4.976498, 5.180631, 4.863329, 4.225089, 3.692261, 3.425874, 
    3.131325, 2.988402, 2.644462, 2.315553, 2.007397, 1.725643, 1.590626, 
    1.386857,
  4.521641, 4.727492, 5.170196, 4.971595, 4.205411, 3.690332, 3.337668, 
    3.163477, 2.940929, 2.530876, 2.182086, 1.902212, 1.688733, 1.565894, 
    1.373133,
  4.805034, 4.951599, 5.220437, 4.768292, 4.224569, 3.681341, 3.332182, 
    3.094912, 2.778603, 2.391265, 2.055842, 1.798023, 1.654203, 1.535488, 
    1.366145,
  4.882858, 4.896246, 4.798244, 4.53573, 4.077374, 3.658636, 3.441742, 
    3.114496, 2.560825, 2.152794, 1.880057, 1.708153, 1.61007, 1.499419, 
    1.362598,
  4.297719, 4.501082, 4.413497, 4.211579, 3.877959, 3.602323, 3.333656, 
    2.587211, 2.106064, 1.885065, 1.742776, 1.626587, 1.565453, 1.46193, 
    1.3544,
  4.887339, 4.734329, 4.6323, 4.476873, 4.325252, 4.153572, 4.000087, 
    3.899827, 3.839363, 3.773678, 3.792028, 3.746608, 3.495224, 3.163703, 
    2.760149,
  5.346019, 5.235638, 5.098322, 4.924997, 4.65775, 4.494824, 4.432621, 
    4.239624, 4.10286, 3.988375, 3.843011, 3.637241, 3.331842, 2.949488, 
    2.589027,
  5.323614, 5.492297, 5.531773, 5.401736, 4.972276, 4.305323, 4.429929, 
    4.222595, 4.006103, 3.842153, 3.639657, 3.393782, 3.110332, 2.856266, 
    2.468216,
  4.919829, 5.13846, 5.391294, 5.649536, 5.342371, 4.724898, 3.950394, 
    3.840281, 3.766633, 3.58891, 3.378705, 3.142011, 2.886275, 2.641544, 
    2.31131,
  4.46144, 4.754405, 4.929075, 5.202793, 5.524415, 4.99697, 4.267519, 
    3.139627, 2.888139, 3.189279, 3.06398, 2.909757, 2.701927, 2.474459, 
    2.147114,
  4.135324, 4.589265, 4.82653, 5.170429, 5.386999, 4.848954, 4.109844, 
    3.548088, 3.255514, 3.065, 2.886736, 2.768565, 2.523547, 2.30566, 1.948812,
  3.774305, 4.229119, 4.992829, 5.316667, 5.145739, 4.263243, 3.596684, 
    3.216491, 3.065542, 2.901616, 2.774852, 2.610918, 2.347235, 2.123513, 
    1.740887,
  3.570791, 3.655191, 3.904514, 4.106555, 3.843789, 3.462675, 3.191814, 
    2.944126, 2.773054, 2.711441, 2.565135, 2.39222, 2.162428, 1.92497, 
    1.563588,
  3.459413, 3.408722, 3.434366, 3.435649, 3.348487, 3.082867, 2.887486, 
    2.679507, 2.579672, 2.535402, 2.379378, 2.211361, 1.969181, 1.729638, 
    1.457936,
  3.405388, 3.33797, 3.326807, 3.343951, 3.334947, 3.171639, 2.867373, 
    2.500935, 2.425847, 2.37025, 2.204026, 2.014014, 1.804555, 1.591224, 
    1.43421,
  4.27066, 4.262416, 4.255798, 4.190647, 4.054972, 3.733029, 3.395129, 
    3.059568, 2.773463, 2.527392, 2.428483, 2.421973, 2.463505, 2.571786, 
    2.688191,
  4.232012, 4.230173, 4.310639, 4.357398, 4.193788, 3.977561, 3.823086, 
    3.506314, 3.146389, 2.838018, 2.628018, 2.605089, 2.650426, 2.651648, 
    2.736982,
  4.02194, 4.103236, 4.360877, 4.568481, 4.470432, 3.821227, 4.030507, 
    3.81482, 3.534405, 3.248798, 2.9879, 2.865853, 2.830429, 2.843779, 
    2.765651,
  3.754267, 3.884959, 4.154918, 4.576334, 4.75801, 4.493512, 3.808777, 
    3.777677, 3.697858, 3.546919, 3.317209, 3.124275, 2.9806, 2.870455, 
    2.728467,
  3.578577, 3.701007, 4.000485, 4.412419, 4.905484, 4.957658, 4.403597, 
    3.425022, 3.278837, 3.711875, 3.511623, 3.302559, 3.065351, 2.899693, 
    2.727787,
  3.382594, 3.426964, 3.718512, 4.098424, 4.652957, 4.899287, 4.354213, 
    4.147607, 4.048808, 3.965934, 3.648143, 3.399078, 3.114989, 2.899999, 
    2.669657,
  3.25507, 3.078469, 3.183307, 3.414454, 3.636147, 3.946404, 3.872973, 
    3.887794, 3.811821, 3.825385, 3.551656, 3.289125, 3.029582, 2.803205, 
    2.540856,
  3.179433, 2.899691, 2.735165, 2.740706, 2.797927, 2.896521, 3.027374, 
    3.095929, 3.256198, 3.387264, 3.23485, 3.033508, 2.852143, 2.644343, 
    2.364008,
  3.145671, 2.864869, 2.657268, 2.569632, 2.569027, 2.623928, 2.575178, 
    2.575116, 2.709468, 2.885429, 2.837247, 2.737468, 2.605138, 2.428534, 
    2.131909,
  3.173738, 2.943611, 2.597624, 2.309626, 2.19662, 2.375522, 2.369845, 
    2.236044, 2.293797, 2.457588, 2.518293, 2.451718, 2.361676, 2.19868, 
    1.893221,
  3.795857, 3.592428, 3.434844, 3.431823, 3.52, 3.673919, 3.759638, 3.667109, 
    3.356124, 3.148537, 3.166561, 3.133118, 3.009529, 2.905876, 2.837885,
  3.75261, 3.349895, 3.205983, 3.29538, 3.441088, 3.677687, 3.92036, 
    3.757898, 3.506591, 3.24112, 3.156176, 3.115603, 2.985325, 2.719023, 
    2.635597,
  3.570767, 3.223995, 3.094257, 3.170673, 3.320564, 3.163023, 3.722723, 
    3.839781, 3.640146, 3.462959, 3.248959, 3.128722, 2.982719, 2.777843, 
    2.592351,
  3.615546, 3.071173, 3.067108, 3.122989, 3.25441, 3.376594, 2.928416, 
    3.242747, 3.360332, 3.495957, 3.358739, 3.192545, 2.967888, 2.703759, 
    2.500847,
  3.583847, 3.028976, 3.087355, 3.102653, 3.110445, 3.255442, 3.15304, 
    2.505844, 2.617204, 3.483205, 3.386174, 3.174564, 2.90742, 2.670647, 
    2.460198,
  3.464289, 3.153081, 3.246153, 3.290884, 3.156802, 3.053187, 2.873859, 
    2.804309, 3.090416, 3.490281, 3.471881, 3.206422, 2.838395, 2.61173, 
    2.426646,
  3.332463, 3.32374, 3.527655, 3.602556, 3.389853, 3.123157, 2.850856, 
    2.555168, 2.70943, 3.223005, 3.350437, 3.102291, 2.788458, 2.572035, 
    2.413588,
  3.27594, 3.465862, 3.936756, 3.946704, 3.577249, 3.266658, 2.940564, 
    2.479461, 2.444365, 2.848581, 3.103779, 2.949922, 2.742892, 2.546471, 
    2.367687,
  3.354987, 3.814299, 4.312762, 4.238518, 3.729039, 3.296462, 2.988486, 
    2.468553, 2.216289, 2.548786, 2.885978, 2.806, 2.687092, 2.491775, 
    2.278345,
  3.844996, 4.452731, 4.70664, 4.403151, 3.812288, 3.329388, 2.990074, 
    2.463611, 2.079384, 2.254006, 2.704703, 2.669733, 2.596589, 2.414025, 
    2.190136,
  2.736415, 2.830964, 3.004344, 3.049299, 3.212472, 3.399187, 3.532938, 
    3.625079, 3.723223, 3.551794, 3.220431, 2.96369, 2.73361, 2.613723, 
    2.50203,
  2.782033, 2.879762, 3.028728, 3.213945, 3.378365, 3.469151, 3.635412, 
    3.764258, 3.793402, 3.675399, 3.331605, 3.033712, 2.829153, 2.590097, 
    2.512663,
  3.023624, 3.007282, 3.321536, 3.523751, 3.796134, 3.780841, 4.110814, 
    4.230995, 4.022933, 3.728851, 3.334533, 3.043358, 2.860055, 2.726168, 
    2.584824,
  3.419456, 3.354272, 3.691622, 4.073738, 4.521393, 4.837092, 4.508602, 
    4.414213, 3.997355, 3.630449, 3.209904, 2.911331, 2.809898, 2.707399, 
    2.56201,
  3.855003, 3.815952, 4.195246, 4.64123, 5.135583, 5.426343, 5.192701, 
    3.896363, 3.253844, 3.260894, 2.961773, 2.738391, 2.747609, 2.686542, 
    2.531752,
  3.891258, 4.28959, 4.745486, 5.188329, 5.506899, 5.36119, 4.964831, 
    4.467289, 3.818587, 3.100965, 2.62285, 2.572711, 2.687686, 2.687433, 
    2.5139,
  4.267162, 4.930391, 5.429746, 5.60076, 5.508776, 4.97333, 4.354538, 
    3.88405, 3.618057, 2.90794, 2.425733, 2.436748, 2.59663, 2.593257, 
    2.434142,
  5.036967, 5.663421, 6.018705, 5.683088, 5.258733, 4.484602, 3.558616, 
    3.447969, 3.409104, 2.71875, 2.284992, 2.356305, 2.477424, 2.417627, 
    2.298174,
  5.885721, 6.437386, 6.342959, 5.499072, 4.979043, 3.935501, 2.997927, 
    3.124786, 3.102779, 2.481572, 2.192421, 2.273014, 2.346735, 2.254172, 
    2.151079,
  6.634229, 6.851945, 6.383711, 5.282698, 4.690689, 3.523858, 2.583278, 
    2.738132, 2.787259, 2.346691, 2.138467, 2.200893, 2.251216, 2.108496, 
    2.026877,
  2.04451, 2.713982, 3.497098, 3.833365, 3.7425, 3.398872, 3.254761, 
    3.384336, 3.629431, 3.854897, 4.099056, 4.334648, 4.239892, 3.853402, 
    3.473069,
  2.962347, 3.912694, 4.38133, 4.449698, 4.152509, 3.645855, 3.461779, 
    3.462576, 3.558327, 3.842003, 4.239518, 4.49194, 4.341331, 3.717918, 
    3.313793,
  4.370255, 5.042226, 5.389349, 5.208729, 4.61956, 3.454976, 3.154586, 
    3.132128, 3.246342, 3.627883, 4.045679, 4.149666, 3.908523, 3.42229, 
    2.976398,
  5.426885, 5.940609, 5.930327, 5.493429, 4.761976, 3.596579, 2.419807, 
    2.428507, 2.720069, 3.231806, 3.397132, 3.24623, 2.881519, 2.59232, 
    2.43601,
  6.144226, 6.372095, 5.97424, 5.478157, 4.838246, 3.645009, 2.571569, 
    1.889767, 2.016931, 2.525308, 2.613576, 2.519355, 2.364251, 2.261986, 
    2.249726,
  6.613986, 6.495787, 6.014808, 5.502478, 5.022298, 3.927962, 2.981172, 
    2.542249, 2.420862, 2.258492, 2.179378, 2.175864, 2.237822, 2.269738, 
    2.254509,
  6.67774, 6.370508, 5.976454, 5.668782, 5.287899, 4.415727, 3.472265, 
    2.877124, 2.563402, 2.141437, 1.984422, 2.087821, 2.174764, 2.293273, 
    2.220922,
  6.389153, 6.119469, 5.833632, 5.689239, 5.413386, 4.805974, 3.988211, 
    3.301634, 2.807002, 2.229231, 1.921853, 2.05148, 2.206369, 2.255799, 
    2.175986,
  6.055979, 5.854376, 5.628391, 5.575171, 5.497488, 5.076264, 4.520589, 
    3.831748, 3.268566, 2.535743, 2.009332, 1.973598, 2.086096, 2.142931, 
    2.072369,
  5.747773, 5.539015, 5.354067, 5.363799, 5.434149, 5.319563, 4.923282, 
    4.359054, 3.803235, 2.948604, 2.273238, 1.976647, 1.965838, 2.022547, 
    2.023149,
  3.083823, 2.983557, 3.017925, 3.355186, 3.589029, 3.767349, 4.010459, 
    3.954238, 3.344509, 2.330862, 1.925735, 2.307038, 2.86849, 3.040132, 
    2.796067,
  3.356334, 3.263705, 3.680746, 4.078942, 4.195507, 4.212711, 4.434217, 
    4.368593, 3.747204, 2.671778, 1.900443, 2.019855, 2.541352, 2.880324, 
    2.889988,
  3.814914, 4.178786, 4.704768, 4.852725, 4.751363, 4.292853, 4.678019, 
    4.894486, 4.394277, 3.244824, 2.095948, 1.841346, 2.006215, 2.627074, 
    2.809684,
  4.564494, 5.057589, 5.306047, 5.454934, 5.30549, 5.180134, 4.594281, 
    4.920154, 4.823125, 4.053501, 2.600819, 1.895799, 1.82238, 2.004732, 
    2.436879,
  4.85438, 5.20578, 5.331381, 5.319778, 5.331044, 5.451581, 5.407171, 
    4.401888, 4.321147, 4.83711, 3.355431, 2.164118, 1.869168, 1.800367, 
    1.958765,
  5.225626, 5.437982, 5.256311, 5.045784, 4.977851, 5.226171, 5.47911, 
    5.588774, 5.638952, 5.363334, 4.037151, 2.735894, 2.057119, 1.849598, 
    1.865834,
  5.25377, 5.133553, 5.013772, 4.912285, 4.715758, 4.852046, 5.148393, 
    5.536162, 5.798296, 5.790118, 4.792615, 3.495618, 2.359829, 1.965109, 
    1.825539,
  5.246682, 4.977178, 4.644659, 4.648111, 4.51085, 4.588384, 4.793557, 
    5.187246, 5.635542, 5.879761, 5.340922, 4.13196, 2.930486, 2.126976, 
    1.85247,
  5.291718, 4.859084, 4.43157, 4.44116, 4.397732, 4.37178, 4.551995, 4.95139, 
    5.474386, 5.815437, 5.559721, 4.580888, 3.465349, 2.50049, 1.919537,
  5.066193, 4.574836, 4.301958, 4.245258, 4.229156, 4.227399, 4.405152, 
    4.7564, 5.317232, 5.769854, 5.639225, 4.792958, 3.799039, 2.920217, 
    2.191461,
  3.713856, 3.151053, 3.987281, 3.899028, 3.849325, 4.130472, 4.423466, 
    4.603493, 3.903011, 2.702111, 2.097468, 1.942233, 1.914149, 1.871643, 
    1.855618,
  3.336135, 3.630045, 4.083676, 3.786873, 3.697912, 3.85028, 4.228422, 
    4.59086, 4.561651, 3.53168, 2.525236, 2.066779, 1.923653, 1.759178, 
    1.742943,
  3.470296, 4.12324, 4.050531, 3.711261, 3.551913, 3.20467, 3.907758, 
    4.513314, 4.804511, 4.41454, 3.294286, 2.38732, 1.998851, 1.855991, 
    1.759551,
  3.967988, 4.408451, 4.06439, 3.752099, 3.724645, 3.618879, 3.289892, 
    3.883472, 4.409256, 4.813604, 4.152995, 3.115324, 2.303682, 1.948018, 
    1.771509,
  4.483611, 4.50423, 4.112099, 3.905533, 3.910121, 4.021386, 3.910671, 
    3.133761, 3.370722, 4.612019, 4.593187, 3.947203, 2.990889, 2.240206, 
    1.884528,
  4.690982, 4.591971, 4.102718, 4.024456, 4.023264, 4.06778, 4.14361, 
    4.164496, 4.304642, 4.555366, 4.60715, 4.407977, 3.799702, 2.911462, 
    2.244818,
  4.89987, 4.750076, 4.213514, 4.160532, 4.131018, 4.235003, 4.229884, 
    4.326857, 4.42742, 4.500655, 4.544247, 4.415417, 4.17407, 3.560903, 
    2.820143,
  5.042724, 4.936444, 4.583458, 4.455819, 4.420928, 4.48829, 4.434524, 
    4.416887, 4.431806, 4.507104, 4.534455, 4.406209, 4.210647, 3.93284, 
    3.34312,
  5.270839, 5.272729, 5.170011, 4.953173, 4.895093, 4.777849, 4.64238, 
    4.596183, 4.609558, 4.60036, 4.611984, 4.505519, 4.184517, 3.991824, 
    3.672948,
  5.311493, 5.364504, 5.288306, 5.127612, 4.96934, 4.839574, 4.779903, 
    4.744056, 4.725828, 4.703823, 4.754266, 4.69091, 4.270759, 3.932166, 
    3.727994,
  5.559754, 3.3078, 3.012749, 3.157317, 3.330345, 3.514612, 3.603626, 
    3.728756, 3.625567, 3.283427, 2.966391, 2.56897, 2.226244, 1.983634, 
    1.861498,
  4.399729, 3.162359, 3.072172, 3.243367, 3.341671, 3.510347, 3.658494, 
    3.687994, 3.749485, 3.789304, 3.663287, 3.272482, 2.853132, 2.374454, 
    2.203829,
  3.627982, 3.135522, 3.158517, 3.210752, 3.215644, 2.771914, 3.268953, 
    3.661471, 3.956369, 4.045588, 4.156587, 3.968183, 3.61205, 3.276248, 
    2.922104,
  3.315627, 3.120562, 3.117261, 3.071038, 3.146008, 3.242316, 3.01252, 
    3.575468, 3.999747, 4.387131, 4.603121, 4.62493, 4.455505, 4.150748, 
    3.741874,
  3.275675, 3.135478, 3.133454, 3.142135, 3.337187, 3.723586, 4.10201, 
    3.717632, 3.882689, 4.840007, 5.21364, 5.305782, 5.279354, 5.059187, 
    4.677324,
  3.318208, 3.226206, 3.235356, 3.388077, 3.748033, 4.418985, 5.121386, 
    5.592104, 5.900028, 6.254828, 6.292105, 6.222023, 6.094228, 5.857819, 
    5.522586,
  3.673414, 3.716758, 3.864946, 4.193789, 4.903391, 5.790216, 6.473702, 
    6.901308, 7.149176, 7.303684, 7.273504, 7.108212, 6.851109, 6.5163, 
    6.174111,
  4.080423, 4.373256, 4.827997, 5.731261, 6.690418, 7.398878, 7.868924, 
    8.122927, 8.279251, 8.317642, 8.20334, 7.942629, 7.589462, 7.153646, 
    6.728615,
  4.594279, 5.395119, 6.616138, 7.638729, 8.331982, 8.783899, 9.047191, 
    9.161665, 9.153598, 9.05999, 8.893471, 8.609389, 8.166223, 7.596354, 
    7.009057,
  6.540873, 7.772036, 8.743342, 9.337576, 9.670608, 9.872321, 9.938328, 
    9.890908, 9.79205, 9.638295, 9.389328, 8.973196, 8.387412, 7.652432, 
    6.777925,
  5.097998, 3.914584, 2.689798, 2.217457, 2.148535, 2.388498, 2.658282, 
    3.183065, 3.783031, 4.505714, 5.475461, 6.740159, 7.480626, 7.580586, 
    7.409992,
  4.810546, 3.802149, 2.892451, 2.476914, 2.317166, 2.489228, 2.753241, 
    3.310561, 3.987805, 5.085411, 6.625026, 7.931365, 8.395107, 7.871041, 
    7.510259,
  4.548337, 3.682806, 3.024923, 2.633204, 2.463544, 2.28159, 2.620727, 
    3.537996, 4.537196, 6.24305, 8.086846, 8.946004, 8.877808, 8.336595, 
    7.772752,
  4.398565, 3.722742, 3.304142, 2.993309, 2.767808, 2.768227, 2.89129, 
    3.968784, 5.149147, 7.844388, 9.274776, 9.411018, 8.723991, 8.018349, 
    7.471778,
  4.338193, 3.77659, 3.490468, 3.301303, 3.265932, 3.483883, 4.077614, 
    4.396906, 5.978549, 9.031935, 9.72122, 9.014407, 7.999499, 7.351927, 
    6.927733,
  4.279672, 3.843416, 3.589783, 3.455548, 3.498632, 3.917748, 4.911637, 
    6.636294, 8.714529, 9.714646, 9.313575, 7.931938, 7.079092, 6.579397, 
    6.254851,
  4.322184, 3.936245, 3.743702, 3.676732, 3.9356, 4.740199, 6.466166, 
    8.851675, 10.00534, 9.673103, 7.97175, 6.747988, 6.109734, 5.761037, 
    5.606012,
  4.353605, 4.10382, 3.982032, 4.118698, 4.854979, 6.508889, 8.720287, 
    9.778175, 9.637251, 7.811699, 6.320961, 5.528695, 5.128856, 4.965803, 
    5.000391,
  4.266148, 4.244913, 4.513381, 5.265203, 6.907878, 8.835044, 9.7705, 
    9.737714, 7.893451, 6.098412, 5.086552, 4.528053, 4.299236, 4.316566, 
    4.48181,
  4.452566, 4.88673, 5.915639, 7.478728, 8.999819, 9.761307, 9.656394, 
    7.831623, 5.956699, 4.696225, 3.993634, 3.637471, 3.624745, 3.800206, 
    4.037615,
  6.543622, 5.923394, 4.965102, 3.880348, 2.981554, 2.322423, 1.934334, 
    1.863478, 1.928918, 2.012449, 2.640596, 3.985361, 4.774733, 4.587357, 
    3.965768,
  6.869175, 6.509265, 5.645144, 4.549574, 3.508941, 2.673627, 2.181754, 
    1.931746, 1.877846, 2.04244, 2.878074, 4.026171, 4.516771, 3.964421, 
    3.580426,
  6.882507, 6.735772, 6.223009, 5.316919, 4.176412, 3.050029, 2.664305, 
    2.402411, 2.235069, 2.399885, 3.268533, 4.115371, 4.293418, 3.912352, 
    3.577349,
  6.783719, 6.655993, 6.412994, 5.979884, 5.127976, 4.124205, 3.159807, 
    2.880941, 2.679177, 3.026625, 3.876072, 4.405927, 4.33582, 4.00142, 
    3.66847,
  6.524669, 6.498244, 6.341258, 6.097038, 5.72438, 5.224326, 4.46141, 
    3.268058, 2.877834, 3.654819, 4.59513, 4.851158, 4.631417, 4.258963, 
    3.831345,
  6.104496, 6.207087, 6.12994, 5.988297, 5.753663, 5.508546, 5.175869, 
    4.640909, 4.424415, 4.853394, 5.245153, 5.221072, 4.902544, 4.434458, 
    3.903691,
  5.699457, 5.821143, 5.826228, 5.712727, 5.536161, 5.346607, 5.117544, 
    4.979807, 4.93384, 5.170893, 5.371892, 5.257593, 4.906146, 4.393277, 
    3.846302,
  5.216744, 5.31773, 5.356766, 5.290329, 5.194353, 5.02856, 4.828059, 
    4.718219, 4.892655, 5.256947, 5.383842, 5.209919, 4.818576, 4.302369, 
    3.823864,
  5.165815, 5.142116, 5.136963, 5.120988, 5.016389, 4.831224, 4.712808, 
    4.862409, 5.255255, 5.507985, 5.485386, 5.218078, 4.815463, 4.384313, 
    3.971661,
  5.396215, 5.198876, 5.098543, 4.976322, 4.790765, 4.749579, 4.860894, 
    5.151303, 5.461016, 5.525695, 5.489451, 5.28412, 4.907378, 4.370533, 
    3.790828,
  4.82194, 4.690736, 4.926147, 5.278934, 5.563002, 5.77025, 5.819945, 5.5734, 
    5.162547, 4.598377, 4.110873, 3.6352, 3.13123, 2.740694, 2.57989,
  4.252348, 4.492095, 5.047249, 5.552595, 5.84864, 5.988791, 6.102662, 
    5.805789, 5.36652, 4.929992, 4.473081, 4.006107, 3.634853, 3.31176, 
    3.072404,
  4.351115, 4.881764, 5.463831, 5.956769, 6.141671, 5.650795, 6.065678, 
    5.947238, 5.585594, 5.285566, 5.013164, 4.762712, 4.547759, 4.016771, 
    3.453586,
  4.835914, 5.363734, 5.830015, 6.245858, 6.409525, 6.305477, 5.632074, 
    5.815242, 5.712417, 5.745558, 5.658171, 5.424119, 4.831592, 4.050888, 
    3.27266,
  5.447654, 5.884704, 6.219235, 6.485665, 6.596837, 6.566957, 6.254086, 
    4.992027, 4.889236, 5.762846, 5.685014, 5.136997, 4.248663, 3.238172, 
    2.757402,
  6.201349, 6.463098, 6.623313, 6.646461, 6.544914, 6.408811, 6.29189, 
    6.041527, 5.9146, 5.761964, 5.333737, 4.516078, 3.335416, 2.65565, 
    2.355226,
  6.840149, 6.83324, 6.772384, 6.550977, 6.384284, 6.148426, 5.970605, 
    5.872787, 5.749022, 5.532421, 4.887552, 3.648844, 2.753423, 2.253605, 
    1.975065,
  7.099051, 6.901833, 6.618137, 6.29, 6.041293, 5.76124, 5.589357, 5.47931, 
    5.405546, 4.82147, 3.70041, 2.801739, 2.21017, 1.830255, 1.634552,
  7.141587, 6.845467, 6.357128, 5.924464, 5.609967, 5.347904, 5.229154, 
    5.263348, 4.91275, 3.800843, 2.991377, 2.327744, 1.873526, 1.590268, 
    1.460154,
  7.157784, 6.736472, 6.104851, 5.451207, 5.031217, 4.8669, 5.025916, 
    4.771803, 3.918581, 3.161376, 2.706449, 2.259664, 1.86944, 1.581905, 
    1.374539,
  4.564432, 4.540592, 5.3153, 6.018901, 6.47956, 6.743817, 6.77281, 6.569669, 
    6.230556, 5.822865, 5.398033, 5.125192, 4.81364, 4.557201, 4.290481,
  4.713554, 5.137384, 6.133391, 6.670547, 6.947762, 6.86982, 6.848512, 
    6.528722, 6.094428, 5.754458, 5.373805, 5.145485, 4.890574, 4.477664, 
    4.307067,
  5.149794, 6.184126, 6.812186, 7.212432, 7.29075, 6.452995, 6.635927, 
    6.525606, 6.148968, 5.713291, 5.373283, 5.177062, 4.96603, 4.774935, 
    4.445347,
  6.074249, 6.878973, 7.275542, 7.514921, 7.48742, 7.183383, 6.060719, 
    6.043313, 5.719576, 5.673297, 5.489041, 5.223672, 5.015026, 4.852605, 
    4.443217,
  6.861699, 7.281833, 7.61451, 7.607469, 7.376355, 7.097871, 6.783235, 
    5.19712, 4.799904, 5.684722, 5.622054, 5.257758, 5.025724, 4.802997, 
    4.31098,
  7.214756, 7.545286, 7.711848, 7.488711, 7.083134, 6.795038, 6.584219, 
    6.35463, 6.172163, 6.047036, 5.679691, 5.280918, 5.11877, 4.814079, 
    3.95228,
  7.536763, 7.703909, 7.595053, 7.241059, 6.856253, 6.516082, 6.353308, 
    6.394168, 6.364405, 6.05114, 5.663146, 5.411775, 5.201857, 4.471214, 
    3.161101,
  7.738714, 7.631446, 7.396339, 7.029884, 6.677802, 6.414483, 6.334958, 
    6.385554, 6.333087, 6.060157, 5.838093, 5.577487, 4.899899, 3.433375, 
    2.393153,
  7.605064, 7.460984, 7.237514, 6.889665, 6.559622, 6.445138, 6.495823, 
    6.58601, 6.51694, 6.352585, 6.109649, 5.276246, 3.688518, 2.330417, 
    1.866696,
  7.242235, 7.06461, 6.904234, 6.729468, 6.630962, 6.683042, 6.794945, 
    6.919722, 6.876537, 6.627269, 5.723454, 3.954727, 2.321604, 1.696346, 
    1.52724,
  2.288861, 2.71122, 3.212473, 3.6426, 4.358759, 4.849752, 4.948586, 
    5.103117, 5.255121, 5.424476, 5.657144, 5.919544, 6.015646, 5.913454, 
    5.863404,
  2.550856, 2.901799, 3.271232, 3.645295, 4.214787, 4.41741, 4.646165, 
    4.901392, 4.978701, 5.291297, 5.661945, 5.999887, 6.205244, 5.996519, 
    5.968494,
  2.843173, 3.189733, 3.4263, 3.802203, 4.270299, 3.961355, 4.347747, 
    4.808161, 5.031778, 5.335604, 5.763722, 6.152486, 6.437975, 6.586234, 
    6.332426,
  3.078422, 3.420658, 3.705147, 4.109356, 4.615678, 4.795407, 4.378125, 
    4.584639, 4.69123, 5.323485, 6.045961, 6.421776, 6.75326, 6.832841, 
    6.287227,
  3.519325, 3.84362, 4.175779, 4.646849, 5.127306, 5.493149, 5.527477, 
    4.374145, 4.258182, 5.620875, 6.442733, 6.707942, 6.984461, 6.889423, 
    6.088853,
  4.427685, 4.793218, 5.137952, 5.530352, 5.725717, 5.836425, 5.934409, 
    5.851313, 5.981356, 6.43413, 6.691588, 6.874148, 7.106693, 6.809032, 
    5.730103,
  5.436039, 5.744611, 6.005338, 6.15907, 6.202915, 6.171582, 6.123216, 
    6.200536, 6.344871, 6.542277, 6.708213, 6.992466, 7.154169, 6.462652, 
    5.030549,
  6.496987, 6.623427, 6.636988, 6.621688, 6.536956, 6.441738, 6.336697, 
    6.252226, 6.354701, 6.590213, 6.8213, 7.152886, 6.994187, 5.74518, 
    3.960642,
  7.0309, 6.99328, 6.908564, 6.834877, 6.723651, 6.547678, 6.37583, 6.363068, 
    6.546174, 6.779795, 7.04018, 7.240156, 6.443818, 4.612416, 2.779444,
  7.279115, 7.092278, 6.953277, 6.783028, 6.618738, 6.427487, 6.308573, 
    6.373062, 6.639979, 6.935071, 7.230309, 6.948561, 5.35748, 3.386439, 
    1.978899,
  2.944956, 2.936996, 2.964303, 3.027021, 3.137367, 3.237336, 3.271822, 
    3.27907, 3.388711, 3.637146, 4.098254, 4.722582, 5.260712, 5.607224, 
    5.976892,
  3.335102, 3.422847, 3.518597, 3.652286, 3.761868, 3.664166, 3.719023, 
    3.88354, 4.13121, 4.565296, 5.019499, 5.46805, 5.876733, 5.830024, 
    6.132226,
  4.082127, 4.268767, 4.364917, 4.44662, 4.424898, 3.875334, 4.121636, 
    4.698605, 5.097621, 5.44579, 5.694561, 5.999257, 6.272686, 6.468881, 
    6.584811,
  4.673826, 4.811355, 4.859915, 4.875787, 4.918365, 4.849952, 4.409787, 
    4.94271, 5.350649, 5.902118, 6.199097, 6.347323, 6.556075, 6.692309, 
    6.726801,
  5.024539, 5.050215, 5.034611, 5.010979, 5.091165, 5.319659, 5.557806, 
    4.612638, 4.529063, 5.847629, 6.461204, 6.575193, 6.720369, 6.762844, 
    6.80171,
  5.057623, 5.145631, 5.184874, 5.234683, 5.419852, 5.695582, 5.999353, 
    6.122834, 6.249148, 6.520441, 6.661422, 6.734444, 6.799518, 6.853961, 
    6.83626,
  5.149322, 5.315792, 5.432775, 5.614095, 5.857996, 6.080928, 6.285934, 
    6.515651, 6.638584, 6.683582, 6.774459, 6.857811, 6.909635, 6.954645, 
    6.711984,
  5.541094, 5.786471, 6.017544, 6.204575, 6.369379, 6.522864, 6.662047, 
    6.745187, 6.797951, 6.885313, 6.979374, 7.027102, 7.064749, 7.01879, 
    6.469038,
  6.657916, 6.826922, 6.940319, 7.00705, 7.041629, 7.015293, 7.028172, 
    7.085088, 7.162371, 7.235014, 7.272919, 7.258709, 7.244226, 6.992596, 
    6.187354,
  7.752478, 7.729572, 7.682735, 7.602525, 7.494473, 7.394616, 7.339579, 
    7.331366, 7.420403, 7.539233, 7.541951, 7.446705, 7.336329, 6.851138, 
    5.811662,
  1.737541, 1.722019, 1.732738, 1.771093, 1.84115, 1.999427, 2.255993, 
    2.580834, 2.933596, 3.240308, 3.57497, 3.936819, 4.223848, 4.400268, 
    4.648497,
  2.189817, 2.102363, 2.039105, 2.055708, 2.182635, 2.429288, 2.784718, 
    3.139875, 3.463241, 3.78915, 4.142372, 4.476066, 4.774019, 4.701842, 
    4.935938,
  3.029831, 3.038446, 2.967345, 2.950364, 3.047447, 2.996848, 3.43147, 
    3.89959, 4.265731, 4.5307, 4.750573, 4.992116, 5.205491, 5.322107, 
    5.419495,
  4.195873, 4.278383, 4.375084, 4.547287, 4.683177, 4.64583, 4.307142, 
    4.707929, 4.961585, 5.2065, 5.339712, 5.378099, 5.449463, 5.474706, 
    5.526127,
  5.516164, 5.586661, 5.651837, 5.696205, 5.760607, 5.805361, 5.736901, 
    4.724051, 4.452266, 5.322911, 5.577883, 5.504866, 5.533392, 5.543075, 
    5.65317,
  5.584229, 5.665474, 5.695168, 5.679581, 5.649391, 5.659091, 5.680055, 
    5.664192, 5.6494, 5.768085, 5.729419, 5.662009, 5.679623, 5.7246, 5.861261,
  5.213956, 5.309218, 5.334626, 5.369776, 5.359392, 5.349615, 5.368968, 
    5.490129, 5.645815, 5.677126, 5.731544, 5.792492, 5.829538, 5.924535, 
    6.098144,
  4.874389, 4.992208, 5.072848, 5.229224, 5.360495, 5.384701, 5.374713, 
    5.371039, 5.437495, 5.578542, 5.747889, 5.858692, 5.966691, 6.100622, 
    6.2802,
  4.991755, 5.091367, 5.255723, 5.535305, 5.89592, 6.174648, 6.257218, 
    6.208351, 6.134407, 6.109544, 6.152895, 6.220006, 6.349892, 6.49598, 
    6.615129,
  4.358741, 4.428253, 4.613317, 5.012167, 5.50032, 6.037916, 6.516255, 
    6.779764, 6.854425, 6.8753, 6.872062, 6.883344, 6.927369, 6.930995, 
    6.898457,
  2.497932, 2.444649, 2.504144, 2.635791, 2.727331, 2.733894, 2.683745, 
    2.580959, 2.435743, 2.247809, 2.105604, 2.028362, 2.007841, 2.050686, 
    2.220962,
  2.742392, 2.466575, 2.300963, 2.244852, 2.239716, 2.299905, 2.380099, 
    2.349086, 2.266104, 2.200638, 2.157058, 2.179204, 2.275725, 2.336972, 
    2.649319,
  3.714927, 3.340694, 2.922129, 2.597587, 2.320071, 2.005975, 2.165873, 
    2.287168, 2.280094, 2.268549, 2.352051, 2.534308, 2.785568, 3.095683, 
    3.505652,
  4.605692, 4.532687, 4.311107, 4.04516, 3.678231, 3.130851, 2.694137, 
    2.920235, 3.05004, 3.158552, 3.327927, 3.499584, 3.779606, 4.11905, 
    4.381349,
  4.826478, 5.110899, 5.232081, 5.161623, 5.047563, 4.87559, 4.476286, 
    3.529684, 3.297631, 4.023502, 4.494327, 4.554348, 4.723368, 4.886041, 
    5.011653,
  4.027363, 4.344891, 4.738288, 5.098549, 5.299098, 5.430134, 5.440308, 
    5.224347, 5.095391, 5.25815, 5.268236, 5.211351, 5.228313, 5.195863, 
    5.116974,
  3.228566, 3.246002, 3.272353, 3.373086, 3.563278, 3.855954, 4.202698, 
    4.634122, 4.923009, 5.07544, 5.204984, 5.302404, 5.325379, 5.255915, 
    5.127759,
  2.885157, 2.812878, 2.749558, 2.690635, 2.721019, 2.929301, 3.33189, 
    3.792693, 4.101442, 4.351336, 4.554356, 4.683278, 4.764018, 4.807579, 
    4.849703,
  2.711071, 2.552251, 2.437184, 2.343456, 2.324324, 2.456253, 2.841953, 
    3.313877, 3.653702, 3.873094, 4.089134, 4.311354, 4.474827, 4.657374, 
    4.89202,
  2.599497, 2.405565, 2.2925, 2.199797, 2.127119, 2.139613, 2.221676, 
    2.572885, 3.261153, 3.830271, 4.243752, 4.610195, 4.97367, 5.298624, 
    5.453845,
  3.351484, 3.324034, 3.317766, 3.313849, 3.346342, 3.370953, 3.399065, 
    3.408825, 3.394103, 3.304773, 3.241091, 3.22227, 3.134929, 2.976034, 
    2.892229,
  3.526655, 3.486847, 3.494261, 3.436917, 3.32115, 3.32003, 3.341158, 
    3.366249, 3.365051, 3.370582, 3.354423, 3.337433, 3.258167, 3.019855, 
    2.981145,
  4.050552, 4.188807, 4.132556, 3.92588, 3.52651, 3.095993, 3.349635, 
    3.434987, 3.367864, 3.281401, 3.255839, 3.257308, 3.22494, 3.160577, 
    3.080992,
  3.796627, 3.970981, 4.227851, 4.487032, 4.370866, 3.773178, 3.241335, 
    3.414072, 3.398921, 3.337706, 3.214048, 3.105736, 3.032195, 2.974406, 
    2.886635,
  3.443455, 3.495065, 3.67842, 3.912963, 4.222859, 4.430419, 3.922255, 
    3.032319, 2.819826, 3.316082, 3.395837, 3.286137, 3.188467, 3.09126, 
    3.044552,
  3.246655, 3.149493, 3.16899, 3.359086, 3.623993, 4.040213, 4.215322, 
    3.991236, 3.869272, 3.877722, 3.839182, 3.84571, 3.883463, 3.879391, 
    3.861387,
  3.156067, 3.019014, 2.944682, 2.912147, 2.934999, 3.041372, 3.346123, 
    3.585829, 3.77865, 3.715865, 3.598878, 3.582287, 3.618077, 3.707177, 
    3.80397,
  3.217053, 2.962395, 2.783756, 2.683901, 2.656662, 2.642557, 2.584033, 
    2.564058, 2.614595, 2.602941, 2.574358, 2.517784, 2.465682, 2.4345, 
    2.48156,
  3.27862, 2.96693, 2.684355, 2.534432, 2.420448, 2.355299, 2.305445, 
    2.238791, 2.189347, 2.153633, 2.248035, 2.295308, 2.301346, 2.297561, 
    2.30884,
  3.336713, 2.873811, 2.548827, 2.472989, 2.351278, 2.220094, 1.997714, 
    1.932203, 1.980528, 2.054746, 2.179359, 2.240506, 2.292253, 2.375162, 
    2.581676,
  3.011969, 2.983482, 2.996247, 2.976754, 2.997951, 3.038524, 3.076871, 
    3.152994, 3.187706, 3.133394, 3.097147, 3.077209, 2.990159, 2.861576, 
    2.767696,
  3.478575, 3.374259, 3.248376, 3.158717, 3.016937, 3.023095, 3.05043, 
    3.064027, 3.081286, 3.097193, 3.091818, 3.073761, 3.025919, 2.884157, 
    2.875618,
  4.258898, 4.292642, 4.127709, 3.902926, 3.420372, 2.871255, 3.163258, 
    3.195693, 3.140887, 3.101373, 3.088244, 3.063356, 3.004654, 2.956691, 
    2.910845,
  4.387245, 4.134823, 3.982316, 3.978689, 4.051847, 3.666887, 3.180543, 
    3.421649, 3.494847, 3.51423, 3.419107, 3.302291, 3.181462, 3.046452, 
    2.899747,
  4.253808, 4.056625, 3.859525, 3.621191, 3.601877, 3.91737, 3.660317, 
    2.764651, 2.584987, 3.077009, 3.342946, 3.352273, 3.320164, 3.213175, 
    3.079631,
  3.958777, 3.810285, 3.717396, 3.59633, 3.369951, 3.274471, 3.352295, 
    3.462981, 3.481693, 3.554541, 3.508576, 3.455213, 3.406477, 3.317036, 
    3.236724,
  3.544793, 3.473639, 3.37901, 3.18056, 3.053132, 3.002922, 2.952378, 
    2.99195, 3.085894, 3.13343, 3.25329, 3.321764, 3.315119, 3.268175, 
    3.222744,
  3.201616, 3.087088, 2.909168, 2.720804, 2.554869, 2.516357, 2.423276, 
    2.373397, 2.315655, 2.290929, 2.38766, 2.49221, 2.611418, 2.697509, 
    2.734934,
  2.788101, 2.633733, 2.485489, 2.298637, 2.122225, 1.989953, 1.897684, 
    1.820041, 1.755729, 1.754223, 1.886382, 2.007585, 2.114419, 2.188217, 
    2.251835,
  2.463654, 2.217625, 2.112121, 1.919416, 1.71855, 1.626383, 1.561558, 
    1.53887, 1.539309, 1.552354, 1.586973, 1.61355, 1.692266, 1.793197, 
    1.917863,
  3.410725, 3.194935, 2.979239, 2.77136, 2.69725, 2.761494, 2.871233, 
    2.979843, 3.005019, 2.89067, 2.795325, 2.679922, 2.541533, 2.460566, 
    2.426652,
  3.827935, 3.621762, 3.372484, 3.076975, 2.800134, 2.613041, 2.622825, 
    2.715408, 2.839294, 2.903412, 2.901449, 2.867094, 2.766561, 2.565025, 
    2.56016,
  4.005075, 4.14265, 4.217665, 4.070086, 3.564313, 2.779209, 2.864789, 
    2.84036, 2.754465, 2.738364, 2.802497, 2.851201, 2.81129, 2.750615, 
    2.676242,
  3.638643, 3.664461, 3.906222, 4.318347, 4.378847, 3.842211, 3.172423, 
    3.20794, 3.045918, 2.891614, 2.828967, 2.827886, 2.839678, 2.795679, 
    2.684257,
  3.365579, 3.291891, 3.309943, 3.55871, 4.021036, 4.164228, 3.731918, 
    2.974221, 2.686186, 3.032307, 2.991284, 2.861872, 2.841217, 2.80776, 
    2.723498,
  3.332524, 3.016197, 2.739587, 2.843377, 3.081598, 3.43349, 3.573404, 
    3.510617, 3.45792, 3.442222, 3.322463, 3.080645, 2.998105, 2.928735, 
    2.846038,
  3.277198, 2.803821, 2.385655, 2.222974, 2.263013, 2.363423, 2.564573, 
    2.904625, 3.07204, 3.183713, 3.278701, 3.235076, 3.139697, 3.05095, 
    2.986779,
  3.123694, 2.665032, 2.24646, 2.015399, 1.880851, 1.808457, 1.76612, 
    1.745418, 1.80115, 2.103054, 2.570998, 2.797835, 2.932509, 2.961365, 
    2.960498,
  3.075182, 2.612887, 2.229543, 1.964111, 1.749773, 1.630352, 1.548474, 
    1.483967, 1.468732, 1.525248, 1.778952, 1.988984, 2.240497, 2.45273, 
    2.632771,
  3.351388, 2.618037, 2.136061, 1.809344, 1.622897, 1.459661, 1.36047, 
    1.333912, 1.356675, 1.444418, 1.494219, 1.560115, 1.658916, 1.803726, 
    2.051528,
  4.152782, 3.869488, 3.660498, 3.488593, 3.363526, 3.157639, 2.964657, 
    2.838525, 2.727901, 2.58023, 2.514036, 2.459523, 2.381575, 2.335935, 
    2.270777,
  4.424258, 4.055778, 3.818137, 3.65234, 3.426943, 3.300939, 3.17101, 
    2.975749, 2.788609, 2.681631, 2.595407, 2.502914, 2.41454, 2.276943, 
    2.303852,
  4.823235, 4.36881, 4.083692, 3.900001, 3.635388, 3.047878, 3.259628, 
    3.211464, 2.986654, 2.768521, 2.675848, 2.582751, 2.466444, 2.390906, 
    2.369749,
  5.143134, 4.562955, 4.063838, 3.748088, 3.734089, 3.486148, 2.966569, 
    3.130156, 3.124646, 2.988011, 2.799211, 2.68765, 2.593135, 2.463848, 
    2.386498,
  4.948802, 3.754199, 2.970972, 2.658657, 2.871326, 3.278367, 3.249309, 
    2.550946, 2.481463, 2.957628, 2.918163, 2.758504, 2.677656, 2.565477, 
    2.435109,
  3.891393, 2.907511, 2.370867, 2.237403, 2.447146, 2.65765, 2.890763, 
    2.86087, 2.722541, 2.786807, 2.884607, 2.840337, 2.709775, 2.617731, 
    2.490263,
  3.658982, 2.972508, 2.595369, 2.34675, 2.192948, 2.091057, 2.071761, 
    1.992959, 1.79912, 1.876968, 2.318274, 2.679288, 2.751983, 2.632913, 
    2.520186,
  3.754321, 3.328807, 2.853099, 2.518348, 2.277064, 2.103886, 1.92286, 
    1.710154, 1.46751, 1.450552, 1.696879, 2.186047, 2.586707, 2.654804, 
    2.535058,
  3.553924, 3.07762, 2.531468, 2.218637, 2.179541, 2.05227, 1.828455, 
    1.60184, 1.427028, 1.332605, 1.421298, 1.750944, 2.329253, 2.602074, 
    2.569001,
  2.55354, 2.176107, 1.912086, 1.734135, 1.592152, 1.447355, 1.321248, 
    1.247343, 1.228169, 1.257884, 1.285199, 1.494183, 2.025695, 2.474137, 
    2.557838,
  4.102125, 4.219934, 4.140201, 3.897689, 3.576816, 3.276733, 3.065558, 
    2.881897, 2.753715, 2.544688, 2.426083, 2.343003, 2.251794, 2.222773, 
    2.292784,
  3.847037, 4.022149, 4.022267, 3.86034, 3.545558, 3.290762, 3.132912, 
    2.98149, 2.85503, 2.727144, 2.590307, 2.475073, 2.357721, 2.125962, 
    2.130038,
  3.887361, 4.081895, 3.992821, 3.824706, 3.516258, 3.016669, 3.15791, 
    3.063561, 2.941423, 2.86322, 2.77744, 2.648827, 2.49035, 2.333725, 
    2.205275,
  4.083957, 4.183601, 4.094968, 3.8999, 3.625699, 3.278816, 2.886139, 
    2.991934, 2.976373, 2.944513, 2.901477, 2.819334, 2.667998, 2.507444, 
    2.317087,
  4.310367, 4.131438, 3.830679, 3.527684, 3.411547, 3.249496, 3.072663, 
    2.490751, 2.400228, 2.896988, 2.948892, 2.893279, 2.799779, 2.664397, 
    2.500196,
  3.924044, 3.377093, 3.012022, 2.764758, 2.716519, 2.841769, 3.053513, 
    2.953861, 2.84366, 2.905452, 2.897785, 2.889874, 2.845849, 2.755126, 
    2.646206,
  3.437963, 3.069771, 2.888886, 2.772609, 2.714339, 2.581043, 2.655329, 
    2.769348, 2.548074, 2.364071, 2.379343, 2.487569, 2.639166, 2.703561, 
    2.663415,
  3.671435, 3.313497, 3.015185, 2.686133, 2.274574, 2.085675, 2.131998, 
    2.365931, 2.329961, 2.034539, 1.809036, 1.776189, 1.851348, 2.112824, 
    2.402863,
  3.349905, 2.944844, 2.359149, 1.808538, 1.477052, 1.501043, 2.013378, 
    2.285083, 2.251925, 2.058139, 1.78278, 1.567968, 1.433708, 1.485526, 
    1.736558,
  2.195942, 1.808922, 1.504767, 1.188264, 1.096391, 1.162866, 1.502441, 
    1.859228, 1.858605, 1.745605, 1.555534, 1.382656, 1.26766, 1.255153, 
    1.38853,
  2.559627, 3.046424, 3.459731, 3.900415, 4.327384, 4.487566, 4.410347, 
    4.139423, 3.775071, 3.317206, 2.907952, 2.564612, 2.30938, 2.285623, 
    2.43242,
  2.447379, 2.643162, 2.992472, 3.387501, 3.74534, 4.084911, 4.229139, 
    4.068477, 3.751863, 3.349658, 2.933699, 2.562339, 2.315676, 2.078854, 
    2.296559,
  2.673239, 2.955006, 3.142699, 3.307989, 3.431977, 3.261643, 3.883358, 
    3.870646, 3.610471, 3.256332, 2.935941, 2.582571, 2.314692, 2.193534, 
    2.237426,
  3.501585, 3.547734, 3.55918, 3.576592, 3.569178, 3.42182, 3.216361, 
    3.442178, 3.3177, 3.061918, 2.826467, 2.581831, 2.358809, 2.209208, 
    2.149524,
  3.518275, 3.48369, 3.523154, 3.516245, 3.477737, 3.447818, 3.289941, 
    2.654222, 2.470244, 2.841421, 2.735954, 2.55331, 2.406939, 2.255189, 
    2.120914,
  3.215732, 3.12489, 3.038422, 3.013495, 3.05267, 3.147238, 3.247345, 
    3.027553, 2.809539, 2.77051, 2.680659, 2.574974, 2.465735, 2.339117, 
    2.190444,
  3.015709, 2.947202, 2.864438, 2.764163, 2.643183, 2.587053, 2.653578, 
    2.759554, 2.899637, 2.810316, 2.665786, 2.601621, 2.522898, 2.423956, 
    2.285209,
  2.527034, 2.371949, 2.235388, 2.038093, 1.794757, 1.642991, 1.564654, 
    1.676361, 2.072558, 2.710474, 2.740729, 2.632318, 2.561413, 2.495937, 
    2.386234,
  1.969079, 1.766723, 1.582315, 1.410041, 1.201538, 1.098326, 1.06982, 
    1.080529, 1.191785, 1.692863, 2.52061, 2.639638, 2.582665, 2.515245, 
    2.423447,
  1.532239, 1.425124, 1.32196, 1.130552, 1.058083, 1.023108, 1.015253, 
    1.092424, 1.228176, 1.485226, 1.938941, 2.483387, 2.526993, 2.443354, 
    2.325523,
  2.640986, 2.782962, 2.816889, 2.871123, 3.098684, 3.487725, 3.871498, 
    3.954915, 3.854898, 3.662309, 3.535959, 3.444049, 3.325594, 3.184212, 
    3.060155,
  2.728161, 2.71545, 2.837961, 2.934962, 3.017753, 3.222098, 3.620775, 
    3.964809, 4.005007, 3.951555, 3.819443, 3.698545, 3.519726, 3.193594, 
    3.080916,
  3.230111, 3.124644, 2.954696, 2.883903, 2.950663, 2.786287, 3.330011, 
    3.798161, 4.047525, 4.085305, 4.061361, 3.929171, 3.71988, 3.50219, 
    3.293689,
  3.257814, 3.333782, 3.387235, 3.278371, 3.052939, 2.996872, 2.899859, 
    3.475124, 3.876068, 4.057443, 4.147246, 4.076686, 3.870344, 3.616017, 
    3.353789,
  2.755835, 2.819278, 3.07565, 3.370173, 3.332246, 3.240315, 3.237165, 
    2.752916, 2.824587, 3.764524, 4.055507, 4.05249, 3.876287, 3.627175, 
    3.381231,
  2.24879, 2.21489, 2.497968, 3.079325, 3.306947, 3.347404, 3.465032, 
    3.408338, 3.332254, 3.677382, 3.882061, 3.927996, 3.754751, 3.53685, 
    3.28969,
  1.961815, 1.900413, 1.914891, 2.215289, 2.670021, 3.013542, 3.293875, 
    3.401477, 3.458081, 3.533292, 3.669519, 3.732887, 3.569899, 3.356624, 
    3.099898,
  1.716631, 1.607221, 1.536729, 1.434802, 1.428236, 1.609728, 2.290737, 
    2.907799, 3.186968, 3.394993, 3.470965, 3.484485, 3.351127, 3.146705, 
    2.898116,
  1.704857, 1.548811, 1.473212, 1.308087, 1.119716, 1.045794, 1.210551, 
    1.877712, 2.579965, 3.058124, 3.257454, 3.238855, 3.09968, 2.912924, 
    2.686782,
  1.798753, 1.512919, 1.347692, 1.165294, 1.032699, 0.9566881, 0.9903604, 
    1.301825, 1.831279, 2.416856, 2.869399, 2.953559, 2.868106, 2.723666, 
    2.517958,
  2.576997, 2.676694, 2.588656, 2.817073, 3.07064, 3.142004, 3.167388, 
    3.246325, 3.386451, 3.451677, 3.689911, 3.877402, 3.982665, 3.995785, 
    3.780584,
  2.690562, 2.691834, 2.48247, 2.68703, 3.005469, 3.119343, 3.146731, 
    3.253147, 3.384149, 3.501604, 3.745899, 3.874354, 3.952761, 3.754711, 
    3.503651,
  2.905558, 3.277749, 2.69416, 2.508575, 2.822309, 2.778764, 3.133036, 
    3.203061, 3.401395, 3.53852, 3.717015, 3.798515, 3.833336, 3.674086, 
    3.275241,
  2.378155, 3.014162, 3.318175, 2.824265, 2.705199, 2.906438, 2.82539, 
    3.238801, 3.336802, 3.482155, 3.666018, 3.692096, 3.657496, 3.443112, 
    2.951751,
  1.916509, 2.417268, 3.040878, 3.213427, 2.821478, 2.939121, 2.94685, 
    2.634492, 2.758235, 3.424002, 3.615335, 3.633158, 3.541956, 3.221389, 
    2.763366,
  1.847153, 1.870271, 2.633673, 3.192727, 3.096454, 3.043258, 3.068497, 
    3.057969, 3.145138, 3.390033, 3.529065, 3.577449, 3.450349, 3.097827, 
    2.797792,
  1.827607, 1.685616, 1.927634, 2.652194, 3.090459, 3.106454, 3.162961, 
    3.237147, 3.203441, 3.283135, 3.37055, 3.460001, 3.333669, 3.088126, 
    2.929462,
  1.731026, 1.636, 1.581843, 1.878991, 2.490928, 2.770956, 3.065243, 
    3.184304, 3.149395, 3.162281, 3.207538, 3.290171, 3.253152, 3.173242, 
    3.110366,
  1.63602, 1.571194, 1.475205, 1.454785, 1.691154, 2.052142, 2.454069, 
    2.937194, 3.188054, 3.155481, 3.136797, 3.169895, 3.238207, 3.261116, 
    3.243402,
  1.551136, 1.420981, 1.306503, 1.15054, 1.241418, 1.461394, 1.763405, 
    2.457603, 2.97811, 3.123664, 3.106887, 3.127066, 3.237503, 3.333315, 
    3.333124,
  2.654989, 3.072129, 2.963388, 3.088963, 3.090735, 2.945055, 2.717162, 
    2.652936, 2.616624, 2.463994, 2.426462, 2.473751, 2.51619, 2.57648, 
    2.69773,
  2.60595, 3.140285, 3.077645, 3.208791, 3.130528, 2.811917, 2.581924, 
    2.594228, 2.557433, 2.514284, 2.543352, 2.626553, 2.684188, 2.625852, 
    2.826343,
  2.392829, 3.118623, 3.22566, 3.242774, 2.912932, 2.398451, 2.463454, 
    2.447618, 2.508788, 2.562824, 2.686316, 2.778476, 2.862248, 2.989999, 
    3.161332,
  2.234922, 2.907805, 3.229302, 3.268118, 2.93353, 2.578315, 2.289621, 
    2.401186, 2.482903, 2.653856, 2.883106, 2.964118, 3.11535, 3.297706, 
    3.457041,
  2.19639, 2.834046, 3.240186, 3.339859, 3.1445, 2.827346, 2.679422, 
    2.261313, 2.252629, 2.879795, 3.104029, 3.240477, 3.447133, 3.619687, 
    3.602804,
  2.171765, 2.751537, 3.193961, 3.396256, 3.36691, 3.164222, 3.02923, 
    3.00277, 3.01718, 3.266981, 3.459516, 3.636129, 3.783915, 3.749932, 
    3.393183,
  2.109957, 2.563194, 3.148807, 3.440859, 3.498391, 3.458738, 3.378705, 
    3.374698, 3.492692, 3.687561, 3.856398, 3.976004, 3.877558, 3.429931, 
    2.846252,
  2.088821, 2.449076, 2.940926, 3.410169, 3.567621, 3.697397, 3.72749, 
    3.807584, 3.918833, 4.031242, 4.07006, 3.976677, 3.466585, 2.767305, 
    2.291503,
  1.930151, 2.2957, 2.711761, 3.090947, 3.374547, 3.634154, 3.777952, 
    3.922831, 4.031366, 4.042335, 3.948935, 3.521655, 2.768366, 2.255825, 
    2.114613,
  1.568943, 1.901674, 2.285334, 2.704751, 3.102178, 3.448151, 3.67656, 
    3.795248, 3.853245, 3.846827, 3.554419, 2.914276, 2.362498, 2.155565, 
    2.110488,
  3.301705, 3.424446, 3.380431, 3.12036, 3.11144, 3.286918, 3.075727, 
    2.511474, 2.142438, 2.196923, 2.233975, 2.279165, 2.298226, 2.28679, 
    2.248942,
  3.26327, 3.202632, 2.891728, 2.431162, 2.403483, 2.991841, 2.978045, 
    2.544606, 2.19698, 2.205744, 2.178741, 2.168109, 2.1527, 2.008584, 
    2.034619,
  3.134234, 3.117567, 2.735567, 2.287424, 2.307364, 2.466429, 2.730497, 
    2.411561, 2.261165, 2.213348, 2.155346, 2.106159, 2.08366, 2.073946, 
    2.074204,
  3.092939, 2.942849, 2.722636, 2.407109, 2.400731, 2.486481, 2.231607, 
    2.218914, 2.169253, 2.183185, 2.154274, 2.091125, 2.075354, 2.090982, 
    2.066646,
  3.113048, 2.950501, 2.772356, 2.518677, 2.402067, 2.411592, 2.208198, 
    1.747675, 1.709552, 2.123668, 2.143793, 2.081381, 2.061489, 2.0422, 
    2.053347,
  3.179851, 2.99035, 2.795239, 2.602279, 2.42792, 2.34703, 2.218302, 
    2.039403, 1.992538, 2.100097, 2.068448, 2.025989, 2.038441, 2.056959, 
    2.13166,
  3.310815, 3.078827, 2.863361, 2.6769, 2.476611, 2.300073, 2.214794, 
    2.132061, 2.095268, 2.055972, 2.027165, 2.065524, 2.154726, 2.281495, 
    2.407438,
  3.535772, 3.296424, 3.050283, 2.835855, 2.613224, 2.42239, 2.258384, 
    2.126657, 2.08686, 2.130655, 2.219998, 2.370555, 2.506231, 2.59334, 
    2.59537,
  3.706218, 3.470701, 3.226065, 2.963588, 2.777728, 2.594169, 2.465512, 
    2.382958, 2.384259, 2.471821, 2.598379, 2.704077, 2.678122, 2.569508, 
    2.42808,
  3.335447, 3.44956, 3.275069, 3.042424, 2.912871, 2.774383, 2.675301, 
    2.612543, 2.62467, 2.705439, 2.699482, 2.568511, 2.347978, 2.130765, 
    1.758435,
  2.602285, 2.535604, 2.662213, 2.716288, 2.481537, 2.279589, 2.300446, 
    2.389756, 2.379632, 2.372946, 2.378955, 2.365041, 2.296921, 2.804338, 
    4.026101,
  2.658303, 2.528714, 2.507041, 2.551129, 2.577372, 2.591768, 2.672551, 
    2.608439, 2.355829, 2.408337, 2.486266, 2.493883, 2.420532, 2.336033, 
    3.213828,
  2.658708, 2.659269, 2.649041, 2.696026, 2.729091, 2.478029, 2.497045, 
    2.315446, 2.258705, 2.377628, 2.416308, 2.503222, 2.510223, 2.393246, 
    2.76082,
  2.429959, 2.559017, 2.662323, 2.635403, 2.608824, 2.328426, 1.949306, 
    2.018665, 2.031295, 2.163563, 2.341861, 2.462849, 2.48632, 2.38307, 
    2.455627,
  2.350542, 2.304978, 2.274744, 2.207061, 2.108678, 2.039159, 1.851517, 
    1.470358, 1.491564, 2.04784, 2.246478, 2.36727, 2.442715, 2.381467, 
    2.330301,
  2.507517, 2.363151, 2.264719, 2.159434, 2.043299, 1.948592, 1.896637, 
    1.853504, 1.79448, 1.889672, 2.07899, 2.205038, 2.320027, 2.294005, 
    2.212489,
  2.724792, 2.546647, 2.394626, 2.296849, 2.150354, 2.009223, 1.934347, 
    1.798241, 1.755319, 1.768723, 1.872778, 2.012582, 2.128468, 2.141615, 
    2.104903,
  2.895565, 2.707936, 2.565622, 2.481903, 2.373703, 2.248206, 2.043912, 
    1.812747, 1.709214, 1.703928, 1.746799, 1.842528, 1.940068, 1.976475, 
    2.00242,
  3.143039, 2.75949, 2.52767, 2.295517, 2.304696, 2.275258, 2.208357, 
    2.08559, 1.988432, 1.887682, 1.834315, 1.851267, 1.891498, 1.930338, 
    1.961209,
  3.269247, 2.652305, 2.213566, 2.013745, 2.128578, 2.212106, 2.296785, 
    2.340418, 2.345576, 2.254467, 2.155577, 2.074947, 2.030419, 2.004705, 
    1.996002,
  2.219727, 2.049856, 1.874993, 1.656075, 1.534662, 1.546639, 1.597669, 
    1.733321, 2.00604, 2.409196, 2.927117, 3.56405, 4.023077, 4.111809, 
    3.894635,
  2.182843, 2.006208, 1.828434, 1.696509, 1.687925, 1.791174, 1.914182, 
    1.927979, 1.969386, 2.1729, 2.595315, 3.172796, 3.717917, 3.853438, 
    3.902936,
  2.449855, 2.281697, 2.178483, 2.147329, 2.114338, 1.897536, 1.946985, 
    1.88762, 1.813842, 1.922062, 2.265667, 2.790916, 3.33531, 3.809942, 
    4.055464,
  2.337218, 2.358551, 2.320433, 2.180102, 2.122661, 1.935059, 1.570912, 
    1.635317, 1.64065, 1.857225, 2.047439, 2.476959, 2.95282, 3.496398, 
    3.919436,
  2.366163, 2.153105, 2.033166, 1.893285, 1.732427, 1.730833, 1.680188, 
    1.323442, 1.340559, 1.837031, 1.956171, 2.228052, 2.644602, 3.163025, 
    3.659582,
  2.707591, 2.5112, 2.271055, 2.034113, 1.874292, 1.685587, 1.653106, 
    1.711664, 1.803476, 1.88464, 1.941367, 2.045908, 2.386804, 2.826903, 
    3.314636,
  3.166316, 2.90598, 2.626151, 2.423055, 2.123477, 1.860936, 1.63448, 
    1.550692, 1.712878, 1.85474, 1.933508, 2.035954, 2.248274, 2.588812, 
    3.050803,
  3.369167, 3.11175, 2.874799, 2.774013, 2.512877, 2.031336, 1.701484, 
    1.485309, 1.512371, 1.707187, 1.915131, 2.03455, 2.150604, 2.33566, 
    2.77551,
  3.750268, 3.253866, 2.708164, 2.446521, 2.381948, 2.225699, 1.946568, 
    1.658758, 1.509461, 1.560452, 1.797336, 1.991302, 2.058052, 2.113123, 
    2.455183,
  3.88364, 3.303044, 2.744222, 2.261674, 2.19423, 2.241384, 2.224256, 
    2.093575, 1.80696, 1.577779, 1.644821, 1.869439, 1.979489, 1.988425, 
    2.165588,
  1.573063, 1.609697, 1.630317, 1.656404, 1.645123, 1.604234, 1.72174, 
    2.062022, 2.506408, 2.764242, 2.89948, 2.87231, 2.612549, 2.412219, 
    2.499957,
  1.806614, 1.69458, 1.661888, 1.663228, 1.663246, 1.542472, 1.684101, 
    1.994795, 2.462575, 2.8106, 3.071866, 3.026823, 2.781424, 2.408276, 
    2.385541,
  2.106014, 1.913282, 1.776537, 1.679119, 1.605395, 1.408134, 1.634243, 
    1.977897, 2.345962, 2.777407, 3.124331, 3.110275, 2.868449, 2.581417, 
    2.433218,
  2.314264, 1.993336, 1.854055, 1.686569, 1.653688, 1.603391, 1.49166, 
    1.815597, 2.189515, 2.675034, 3.03106, 3.103861, 2.880173, 2.644433, 
    2.476339,
  2.767825, 2.338519, 2.10339, 1.926522, 1.795542, 1.698321, 1.614325, 
    1.519179, 1.783929, 2.438267, 2.874742, 3.045105, 2.903477, 2.68066, 
    2.552103,
  3.756686, 3.360266, 2.890405, 2.433425, 2.136261, 1.832438, 1.602828, 
    1.723103, 1.948644, 2.299385, 2.700152, 2.940387, 2.894226, 2.731356, 
    2.638933,
  4.624542, 4.292852, 3.833743, 3.34052, 2.805073, 2.132053, 1.691163, 
    1.657876, 1.92175, 2.175389, 2.497296, 2.757754, 2.856017, 2.79281, 
    2.717645,
  5.232853, 4.86757, 4.300916, 3.611088, 3.228853, 2.41946, 1.772839, 
    1.584661, 1.743082, 1.999302, 2.265886, 2.545405, 2.777676, 2.878776, 
    2.840895,
  5.958511, 5.560679, 4.833351, 3.661468, 2.975925, 2.451033, 1.961928, 
    1.671878, 1.655205, 1.826955, 2.081092, 2.329739, 2.635023, 2.957182, 
    3.035838,
  6.754212, 6.145454, 5.520443, 4.284199, 3.070348, 2.433423, 2.068092, 
    1.831505, 1.703975, 1.693689, 1.914389, 2.178107, 2.431999, 2.837313, 
    3.200204,
  1.74406, 1.617667, 1.637876, 1.680769, 1.805156, 2.076456, 2.232334, 
    2.330396, 2.323823, 2.162403, 2.049411, 2.160843, 2.344429, 2.578085, 
    2.760217,
  2.238409, 1.899457, 1.859699, 1.855695, 2.123042, 2.359422, 2.570369, 
    2.524796, 2.405908, 2.270564, 2.117383, 2.178061, 2.302411, 2.347955, 
    2.631883,
  2.628488, 2.361441, 2.28309, 2.392189, 2.788004, 2.701558, 2.749109, 
    2.522414, 2.318781, 2.273379, 2.184322, 2.202054, 2.296849, 2.445293, 
    2.685841,
  2.732774, 2.709225, 2.839098, 3.137867, 3.373915, 3.164492, 2.318136, 
    2.279937, 2.243936, 2.291312, 2.266186, 2.256533, 2.290221, 2.435652, 
    2.690298,
  2.978134, 3.017783, 3.236603, 3.617579, 3.448076, 2.702533, 2.245927, 
    2.034965, 1.960962, 2.312014, 2.332006, 2.278866, 2.295979, 2.420774, 
    2.700519,
  3.40947, 3.28869, 3.602581, 3.649806, 3.212551, 2.444709, 2.280077, 
    2.276476, 2.297108, 2.371432, 2.328388, 2.265731, 2.281032, 2.426454, 
    2.682954,
  3.875713, 3.606937, 3.706532, 3.463199, 2.890538, 2.379506, 2.338391, 
    2.322225, 2.35529, 2.353846, 2.268676, 2.218649, 2.26774, 2.445901, 
    2.610694,
  4.123889, 3.892859, 3.689898, 3.106004, 2.532668, 2.278248, 2.280523, 
    2.272511, 2.267483, 2.237884, 2.17591, 2.1681, 2.271731, 2.429237, 
    2.462787,
  4.298273, 4.039387, 3.452468, 2.621531, 2.14104, 2.053617, 2.114775, 
    2.176913, 2.15408, 2.110916, 2.091008, 2.149606, 2.255891, 2.330669, 
    2.293571,
  4.417773, 3.888492, 2.962399, 2.204489, 1.958999, 1.945181, 2.009702, 
    2.065866, 2.064611, 2.03416, 2.04507, 2.119794, 2.181822, 2.199815, 
    2.198293,
  3.175913, 2.86436, 2.492883, 2.079733, 1.727486, 1.557727, 1.533887, 
    1.6027, 1.770583, 1.927063, 2.031044, 2.124578, 2.213733, 2.191101, 
    2.116437,
  2.684364, 2.599368, 2.468149, 2.251562, 1.990563, 1.814736, 1.807529, 
    1.939729, 2.110318, 2.295183, 2.352184, 2.321103, 2.3874, 2.246313, 
    2.184132,
  2.431969, 2.306206, 2.228942, 2.174903, 2.139752, 1.909537, 2.098163, 
    2.28091, 2.435272, 2.608078, 2.485136, 2.325128, 2.420205, 2.434353, 
    2.33414,
  2.715966, 2.540087, 2.596606, 2.598276, 2.564182, 2.477005, 2.241294, 
    2.421038, 2.66965, 2.616852, 2.236993, 2.302958, 2.475862, 2.454179, 
    2.394288,
  3.103133, 3.155726, 2.986819, 2.88683, 2.492897, 2.337069, 2.46184, 
    2.107666, 2.002381, 2.157345, 2.149696, 2.454365, 2.509584, 2.51929, 
    2.489101,
  2.818273, 2.748388, 2.655749, 2.624647, 2.547669, 2.448733, 2.544102, 
    2.439009, 2.150803, 2.170272, 2.363698, 2.512815, 2.524848, 2.518353, 
    2.480184,
  2.567894, 2.532825, 2.539053, 2.503925, 2.46128, 2.409581, 2.319611, 
    2.211514, 2.207609, 2.322062, 2.437819, 2.484152, 2.469058, 2.411313, 
    2.354849,
  2.459725, 2.422223, 2.39688, 2.381908, 2.351451, 2.297098, 2.240086, 
    2.15659, 2.289553, 2.376098, 2.414167, 2.419672, 2.362196, 2.262268, 
    2.170022,
  2.357816, 2.33875, 2.301082, 2.246152, 2.202196, 2.174734, 2.177979, 
    2.239125, 2.324012, 2.333852, 2.357467, 2.342819, 2.28883, 2.207016, 
    2.169776,
  2.211822, 2.145183, 2.032815, 1.947394, 2.018525, 2.09185, 2.127126, 
    2.17313, 2.231541, 2.238887, 2.26777, 2.265038, 2.221414, 2.19732, 
    2.220562,
  2.989013, 3.204481, 3.152929, 2.793715, 2.158915, 1.753133, 1.558537, 
    1.362465, 1.231207, 1.150756, 1.177785, 1.247426, 1.326151, 1.429689, 
    1.545218,
  2.435733, 2.540384, 2.964402, 2.916924, 2.436663, 1.93998, 1.646504, 
    1.41091, 1.266132, 1.203544, 1.218168, 1.331887, 1.516089, 1.592982, 
    1.74009,
  2.529107, 2.290589, 2.544963, 2.777924, 2.560512, 1.965476, 1.757952, 
    1.569621, 1.3964, 1.307466, 1.370077, 1.603149, 1.840507, 2.065421, 
    2.166846,
  2.407412, 2.33996, 2.4503, 2.600854, 2.546023, 2.233087, 1.71513, 1.578874, 
    1.474294, 1.573528, 1.752578, 1.961274, 2.199912, 2.303377, 2.277974,
  2.382034, 2.325996, 2.404135, 2.556248, 2.437279, 2.315973, 1.90124, 
    1.426146, 1.312094, 1.71214, 1.964072, 2.240801, 2.316665, 2.290413, 
    2.27282,
  2.420426, 2.337055, 2.356577, 2.424278, 2.354279, 2.226003, 2.031769, 
    1.883896, 1.851253, 2.138854, 2.353817, 2.345261, 2.293789, 2.293992, 
    2.302763,
  2.468014, 2.379843, 2.378381, 2.366079, 2.346465, 2.244102, 2.102155, 
    2.116806, 2.280631, 2.321642, 2.278229, 2.279495, 2.259342, 2.259088, 
    2.289415,
  2.477084, 2.417418, 2.368174, 2.36499, 2.376928, 2.394283, 2.318604, 
    2.270279, 2.283398, 2.250812, 2.272656, 2.273484, 2.268826, 2.243309, 
    2.21374,
  2.648253, 2.55927, 2.56628, 2.524482, 2.452814, 2.399786, 2.299122, 
    2.246865, 2.224998, 2.235147, 2.270956, 2.319104, 2.359351, 2.406751, 
    2.371936,
  2.70701, 2.569558, 2.419074, 2.286696, 2.257346, 2.18162, 2.146924, 
    2.098006, 2.093389, 2.095811, 2.115026, 2.175201, 2.289498, 2.432972, 
    2.525658,
  2.700207, 2.760291, 2.82603, 2.908219, 2.961178, 2.844587, 2.639227, 
    2.144341, 1.708541, 1.31307, 1.11152, 1.083749, 1.088703, 1.12357, 
    1.239361,
  2.68568, 2.676069, 2.780803, 2.889011, 2.802588, 2.659895, 2.349954, 
    1.819761, 1.409698, 1.150129, 1.067313, 1.085836, 1.15436, 1.210182, 
    1.439455,
  3.005494, 2.641675, 2.807207, 2.83209, 2.761612, 2.32783, 2.037868, 
    1.557375, 1.294015, 1.158475, 1.11856, 1.192934, 1.366407, 1.69692, 
    1.960052,
  2.984963, 2.843989, 2.890613, 2.855757, 2.74672, 2.268672, 1.546987, 
    1.35575, 1.258282, 1.258015, 1.285909, 1.427477, 1.795833, 2.124316, 
    2.15783,
  2.906706, 2.928572, 2.950037, 2.914728, 2.607424, 2.156986, 1.542144, 
    1.143442, 1.063792, 1.349067, 1.469583, 1.847235, 2.210237, 2.227609, 
    2.177799,
  2.904584, 2.951061, 2.959871, 2.834384, 2.421365, 2.048785, 1.714022, 
    1.568716, 1.456665, 1.580082, 2.00998, 2.352035, 2.28975, 2.198679, 
    2.188769,
  2.946853, 2.926195, 2.857923, 2.707735, 2.482406, 2.220597, 1.823703, 
    1.750177, 1.754778, 2.13127, 2.354871, 2.339519, 2.266914, 2.191285, 
    2.186102,
  2.829802, 2.79178, 2.712481, 2.602948, 2.436714, 2.277701, 1.979715, 
    1.862038, 2.097987, 2.286974, 2.360034, 2.41016, 2.382052, 2.235748, 
    2.185976,
  2.801018, 2.679689, 2.6205, 2.534883, 2.377937, 2.267126, 2.115029, 
    2.108236, 2.244539, 2.303376, 2.341808, 2.42109, 2.444108, 2.3505, 
    2.202059,
  2.844322, 2.713576, 2.523867, 2.309283, 2.251676, 2.206033, 2.124472, 
    2.107277, 2.095349, 2.085049, 2.078876, 2.249503, 2.419888, 2.442345, 
    2.329409,
  2.684062, 2.551772, 2.530371, 2.603245, 2.607792, 2.566161, 2.748787, 
    2.879609, 2.85932, 2.868949, 2.714651, 2.328144, 1.920823, 1.572871, 
    1.389475,
  2.725095, 2.631297, 2.64227, 2.641137, 2.492104, 2.536421, 2.719781, 
    2.798523, 2.777146, 2.614834, 2.163335, 1.604022, 1.276158, 1.169821, 
    1.460046,
  3.267834, 2.888979, 2.623827, 2.573409, 2.500204, 2.418243, 2.555953, 
    2.489523, 2.206254, 1.700233, 1.256395, 1.138368, 1.287656, 1.793992, 
    2.107051,
  3.036485, 2.771526, 2.646839, 2.547123, 2.61342, 2.544578, 2.070981, 
    1.740166, 1.305058, 1.128169, 1.149414, 1.41537, 1.983722, 2.221464, 
    2.227017,
  2.907151, 2.753416, 2.720259, 2.622475, 2.516835, 2.229352, 1.512641, 
    0.9404567, 0.854208, 1.198003, 1.461582, 1.983513, 2.254116, 2.226274, 
    2.20718,
  2.883831, 2.695959, 2.586057, 2.405967, 1.985978, 1.582527, 1.280757, 
    1.149546, 1.154503, 1.526993, 1.980029, 2.252419, 2.211344, 2.210279, 
    2.226759,
  2.864821, 2.596461, 2.357441, 2.135499, 1.91073, 1.642115, 1.369693, 
    1.444326, 1.69966, 2.120363, 2.2445, 2.201213, 2.172813, 2.212228, 2.25204,
  2.984492, 2.724068, 2.491698, 2.319643, 2.136845, 1.936766, 1.689833, 
    1.803001, 2.141173, 2.271751, 2.25273, 2.216327, 2.202812, 2.245876, 
    2.271557,
  3.215137, 2.973449, 2.72789, 2.492773, 2.291536, 2.067318, 1.976479, 
    2.176938, 2.312529, 2.286494, 2.262874, 2.252569, 2.239559, 2.281247, 
    2.313852,
  3.358688, 3.115876, 2.88322, 2.521775, 2.295714, 2.17044, 2.146558, 
    2.240552, 2.27706, 2.259452, 2.278054, 2.308851, 2.308863, 2.326972, 
    2.364478,
  2.303159, 2.162802, 2.152658, 2.177819, 2.121254, 2.111328, 2.183786, 
    2.264794, 2.30053, 2.273231, 2.336259, 2.371493, 2.286266, 2.203269, 
    2.085899,
  2.267727, 2.23118, 2.129828, 2.029909, 1.945853, 1.97083, 2.087312, 
    2.160125, 2.193463, 2.18439, 2.079381, 1.954041, 1.845415, 1.644963, 
    1.656259,
  2.500868, 2.220187, 2.019889, 1.875922, 1.685868, 1.555578, 1.792927, 
    1.872559, 1.888316, 1.876661, 1.872762, 1.906082, 1.981259, 2.00973, 
    1.983442,
  2.77737, 2.483604, 2.173327, 1.80778, 1.618025, 1.56289, 1.522432, 
    1.758742, 1.863243, 1.973759, 2.05433, 2.031679, 1.958709, 1.862213, 
    1.775535,
  2.914234, 2.545797, 2.334467, 1.860288, 1.526248, 1.648096, 1.750618, 
    1.538846, 1.699642, 2.0653, 2.063783, 1.98284, 1.869868, 1.719072, 
    1.574264,
  2.957535, 2.59639, 2.255374, 1.868158, 1.675113, 1.686247, 1.876729, 
    2.034837, 2.111773, 2.141574, 2.104913, 2.030744, 1.903964, 1.740439, 
    1.584497,
  2.944948, 2.600441, 2.232299, 2.031882, 2.077046, 2.04696, 2.01678, 
    2.155802, 2.199193, 2.191818, 2.163668, 2.119529, 2.020088, 1.874358, 
    1.733066,
  2.864099, 2.520735, 2.34037, 2.29156, 2.255319, 2.310719, 2.273251, 
    2.215263, 2.216238, 2.226043, 2.222721, 2.195361, 2.137382, 2.048613, 
    1.929637,
  2.826956, 2.632818, 2.511468, 2.432172, 2.320213, 2.28532, 2.246411, 
    2.239591, 2.247564, 2.268617, 2.279668, 2.267473, 2.231558, 2.184163, 
    2.127958,
  2.911349, 2.842443, 2.41495, 2.128459, 2.202296, 2.248258, 2.264809, 
    2.265373, 2.271208, 2.274816, 2.278727, 2.277921, 2.271818, 2.261752, 
    2.245006,
  2.105629, 1.985597, 1.824655, 1.723884, 1.712563, 1.827187, 1.876855, 
    1.915979, 1.918597, 1.800559, 1.707644, 1.63598, 1.554713, 1.538163, 
    1.625622,
  1.838094, 1.693905, 1.565022, 1.573303, 1.732786, 1.877608, 1.926309, 
    1.886871, 1.844849, 1.774726, 1.662413, 1.538152, 1.450845, 1.356144, 
    1.496178,
  1.731255, 1.454039, 1.438817, 1.647244, 1.876804, 1.811467, 1.970355, 
    1.93798, 1.870371, 1.770993, 1.612294, 1.461728, 1.383139, 1.356898, 
    1.51012,
  2.022357, 1.848234, 1.769434, 1.839122, 2.130703, 2.225102, 1.854367, 
    1.966968, 1.889422, 1.784027, 1.601852, 1.462618, 1.402931, 1.364221, 
    1.481054,
  2.363222, 2.088567, 2.127219, 2.190487, 2.271885, 2.282354, 2.290649, 
    1.765488, 1.674191, 1.807628, 1.664857, 1.526573, 1.466083, 1.47114, 
    1.539973,
  2.668677, 2.261891, 2.289898, 2.367324, 2.343664, 2.246978, 2.243913, 
    2.179101, 2.047651, 1.857795, 1.72755, 1.592021, 1.550953, 1.565133, 
    1.598251,
  2.836402, 2.519582, 2.479068, 2.553384, 2.570925, 2.410759, 2.231647, 
    2.163398, 2.075633, 1.969851, 1.814368, 1.680287, 1.605742, 1.598983, 
    1.608219,
  2.875291, 2.717704, 2.727226, 2.677266, 2.638166, 2.527939, 2.346782, 
    2.183999, 2.101251, 2.02171, 1.897456, 1.758792, 1.650059, 1.567683, 
    1.524781,
  2.905288, 2.867994, 2.846883, 2.676772, 2.521419, 2.416037, 2.312814, 
    2.188921, 2.096953, 2.040247, 1.985723, 1.897653, 1.789028, 1.687036, 
    1.596941,
  3.051282, 2.974192, 2.493542, 2.283006, 2.301129, 2.345566, 2.338315, 
    2.246936, 2.110936, 2.03844, 1.996122, 1.972264, 1.945339, 1.923568, 
    1.900971,
  2.595185, 2.712906, 2.851665, 2.954879, 2.967734, 2.900172, 2.774905, 
    2.554646, 2.286526, 2.018117, 1.847356, 1.681268, 1.536016, 1.402672, 
    1.31251,
  2.043161, 2.039968, 2.07581, 2.104101, 2.105133, 2.055756, 1.991554, 
    1.903823, 1.834988, 1.755637, 1.637951, 1.49289, 1.425894, 1.250673, 
    1.22377,
  1.966199, 1.860458, 1.854294, 1.837676, 1.782415, 1.605766, 1.753816, 
    1.76437, 1.756931, 1.665829, 1.473813, 1.380077, 1.358374, 1.348836, 
    1.321726,
  2.336009, 2.229057, 2.068032, 1.935226, 1.911335, 1.847852, 1.596157, 
    1.778893, 1.666367, 1.524549, 1.419213, 1.420344, 1.444921, 1.498018, 
    1.579064,
  2.556377, 2.479702, 2.376612, 2.189179, 2.130343, 2.07116, 2.006041, 
    1.480792, 1.336646, 1.501168, 1.511103, 1.547586, 1.642943, 1.671226, 
    1.667061,
  2.702318, 2.593615, 2.47538, 2.371109, 2.217339, 2.136965, 2.024801, 
    1.878963, 1.673137, 1.579344, 1.59438, 1.615321, 1.64598, 1.616688, 
    1.515419,
  2.83153, 2.82416, 2.740935, 2.654417, 2.558941, 2.269583, 1.98595, 
    1.817157, 1.668321, 1.609067, 1.601591, 1.597694, 1.55593, 1.492686, 
    1.430917,
  2.993896, 3.018326, 2.90837, 2.817538, 2.710412, 2.484629, 2.054145, 
    1.801707, 1.65148, 1.579503, 1.54844, 1.533832, 1.492847, 1.450722, 
    1.443248,
  3.135148, 3.210375, 3.086301, 2.820135, 2.649068, 2.472567, 2.051202, 
    1.800205, 1.681876, 1.5849, 1.524776, 1.526935, 1.594212, 1.709126, 
    1.835157,
  3.362487, 3.15734, 2.806175, 2.539102, 2.478908, 2.34316, 2.035467, 
    1.814843, 1.687961, 1.661583, 1.733507, 1.890557, 2.102594, 2.347251, 
    2.607333,
  2.857137, 3.224768, 3.64806, 4.08859, 4.498582, 4.824485, 5.087849, 
    5.229372, 5.266478, 5.161638, 5.012353, 4.815612, 4.532474, 4.165972, 
    3.758109,
  2.400416, 2.795482, 3.215021, 3.526956, 3.808609, 3.948966, 4.101376, 
    4.25341, 4.23143, 4.14575, 3.974028, 3.770502, 3.541715, 3.109029, 
    2.824366,
  2.212227, 2.141183, 2.342475, 2.590461, 2.794483, 2.743019, 2.963364, 
    2.946066, 2.959189, 2.874711, 2.766037, 2.613836, 2.434013, 2.212575, 
    1.958756,
  2.369517, 2.20024, 1.990933, 1.910729, 2.020419, 2.091543, 2.052542, 
    2.178554, 2.042656, 1.928407, 1.860816, 1.744992, 1.655036, 1.567242, 
    1.44151,
  2.496405, 2.285997, 2.103166, 1.842112, 1.740466, 1.822032, 1.747501, 
    1.389168, 1.319599, 1.539818, 1.509064, 1.518286, 1.504409, 1.466229, 
    1.468344,
  2.620572, 2.401913, 2.220422, 1.966981, 1.732745, 1.642024, 1.642349, 
    1.563369, 1.401125, 1.407191, 1.394134, 1.397722, 1.407474, 1.406703, 
    1.455416,
  2.992959, 2.553411, 2.47865, 2.272967, 2.002839, 1.679922, 1.438243, 
    1.368478, 1.34164, 1.338707, 1.340973, 1.35352, 1.352531, 1.337188, 
    1.34615,
  3.917292, 3.269644, 3.131489, 2.85474, 2.339637, 1.845994, 1.54849, 
    1.438949, 1.423487, 1.454211, 1.467257, 1.486878, 1.508192, 1.481287, 
    1.400951,
  4.041552, 3.765485, 3.689809, 3.271013, 2.629102, 2.108927, 1.906895, 
    1.968621, 2.092021, 2.19993, 2.254734, 2.256961, 2.187285, 2.068968, 
    1.804421,
  4.038087, 3.842913, 3.695229, 2.92493, 2.31459, 2.287912, 2.420656, 
    2.654142, 2.864843, 2.995243, 3.059171, 3.067699, 3.01403, 2.838178, 
    2.575694,
  2.503378, 3.208885, 3.955026, 4.459637, 5.009972, 5.691623, 6.378085, 
    6.839779, 7.066282, 7.194243, 7.37847, 7.432809, 7.329151, 7.179989, 
    7.032523,
  2.356916, 2.659539, 3.366771, 4.091595, 4.782711, 5.325657, 5.811289, 
    6.438375, 6.729591, 6.951837, 6.991695, 7.005958, 6.923004, 6.58211, 
    6.497849,
  2.485778, 2.420231, 2.673613, 3.114705, 3.767481, 4.211597, 4.830159, 
    5.219991, 5.778687, 6.13982, 6.354415, 6.389342, 6.333065, 6.095051, 
    5.803114,
  2.681593, 2.537733, 2.538246, 2.530493, 2.731024, 3.110682, 3.303508, 
    4.097166, 4.490998, 4.785321, 5.254565, 5.415439, 5.297952, 4.970802, 
    4.645643,
  3.044434, 2.67548, 2.664902, 2.600424, 2.333314, 2.457196, 2.46541, 
    2.296023, 2.519175, 3.099865, 3.709372, 4.001231, 3.96233, 3.729908, 
    3.395936,
  3.59116, 3.101102, 2.94141, 2.906429, 2.487595, 2.278659, 2.202413, 
    1.910616, 1.732546, 1.762917, 2.002594, 2.399447, 2.641969, 2.599623, 
    2.431504,
  4.23234, 3.669245, 3.439556, 3.177694, 2.910003, 2.688342, 2.409253, 
    2.159664, 1.814921, 1.420702, 1.239292, 1.276802, 1.410308, 1.573805, 
    1.66383,
  4.470465, 4.13292, 3.874866, 3.516061, 3.411753, 3.499199, 3.453732, 
    3.338497, 3.097388, 2.767287, 2.219502, 1.653884, 1.37633, 1.308975, 
    1.341063,
  4.158926, 4.090651, 4.291153, 3.953518, 3.939755, 3.930734, 3.828376, 
    3.722779, 3.568023, 3.321867, 3.056813, 2.619443, 2.014801, 1.591352, 
    1.448745,
  3.565573, 3.591564, 3.663426, 3.775076, 3.995217, 3.954425, 3.879111, 
    3.738866, 3.554225, 3.22493, 3.010498, 2.867627, 2.60684, 2.120011, 
    1.714468,
  3.23536, 3.584335, 3.827004, 4.014127, 4.655273, 5.122819, 5.726336, 
    6.084725, 6.083846, 5.918895, 5.785577, 5.51843, 5.180199, 5.046474, 
    5.166288,
  3.19981, 3.522109, 3.819443, 3.688123, 4.111733, 4.640361, 5.30478, 6.0505, 
    6.493455, 6.61698, 6.592305, 6.369689, 5.992766, 5.245276, 5.180672,
  3.302979, 3.595976, 3.988952, 3.645691, 3.526571, 3.639191, 4.238079, 
    4.798883, 5.507759, 6.057228, 6.477801, 6.585441, 6.492052, 6.200182, 
    5.882754,
  3.478788, 3.79203, 4.164839, 3.891791, 3.531593, 3.516773, 3.230204, 
    3.929447, 4.424637, 4.869664, 5.56883, 6.0213, 6.233781, 6.183374, 
    6.083885,
  3.684944, 3.924686, 4.192854, 4.153917, 3.83675, 3.638644, 3.111683, 
    2.478684, 2.528584, 3.134244, 3.859185, 4.763534, 5.425458, 5.770604, 
    5.873772,
  3.970315, 4.119133, 4.207747, 3.994456, 3.995077, 4.008524, 3.552236, 
    2.95179, 2.50934, 2.192614, 2.129853, 2.574347, 3.663227, 4.764097, 
    5.288465,
  4.148643, 4.240555, 4.177129, 3.871408, 3.985429, 4.196594, 3.793515, 
    3.537221, 3.209019, 2.697006, 1.997456, 1.68762, 1.841775, 2.695267, 
    3.909652,
  4.072381, 4.192387, 4.132463, 3.855751, 4.143263, 4.095012, 3.667872, 
    3.401182, 3.201933, 3.012075, 2.83636, 2.293931, 1.830283, 1.764634, 
    2.187565,
  3.949336, 4.054927, 4.207775, 4.204428, 4.054839, 3.83587, 3.526292, 
    3.317129, 3.189454, 3.023767, 2.787102, 2.517551, 2.047766, 1.756538, 
    1.626561,
  3.790302, 4.087138, 4.301732, 4.055789, 3.690545, 3.445541, 3.338345, 
    3.232794, 3.170294, 3.070687, 2.823626, 2.572924, 2.266701, 1.887602, 
    1.644051,
  3.759861, 3.53235, 3.770328, 3.673223, 3.276344, 3.190621, 4.18399, 
    5.223636, 5.588305, 5.415029, 5.091154, 4.667791, 4.753746, 4.98771, 
    5.147355,
  3.991481, 3.57803, 3.579973, 3.800206, 3.480694, 3.084638, 3.444741, 
    4.236523, 4.957581, 5.546768, 5.667401, 5.399114, 4.95854, 4.293939, 
    4.26199,
  4.241625, 3.722664, 3.487681, 3.723517, 3.690734, 3.138555, 3.154359, 
    3.359924, 3.732805, 4.305474, 5.066781, 5.414394, 5.447914, 5.294012, 
    5.036603,
  4.459887, 4.124694, 3.792244, 3.766545, 3.769296, 3.813485, 3.147332, 
    3.1522, 3.112369, 3.038463, 3.261327, 3.691314, 4.15912, 4.525817, 4.80024,
  4.568007, 4.363423, 4.129536, 3.936335, 3.852663, 3.990376, 3.862914, 
    2.969549, 2.651851, 2.566397, 2.250098, 2.228774, 2.545312, 3.097644, 
    3.689508,
  4.583089, 4.514028, 4.335338, 4.083166, 3.913632, 4.02305, 3.975458, 
    3.781781, 3.389599, 2.68568, 2.097631, 1.895782, 1.937614, 2.143766, 
    2.582189,
  4.604996, 4.594443, 4.468983, 4.242836, 4.126545, 4.228108, 4.00045, 
    3.664225, 3.299172, 2.893082, 2.312596, 2.070849, 2.023092, 1.836871, 
    1.86633,
  4.661915, 4.691793, 4.56325, 4.30623, 4.151777, 4.241806, 3.954604, 
    3.558255, 3.190159, 2.887206, 2.66129, 2.491409, 2.192026, 1.749977, 
    1.590441,
  4.748299, 4.751111, 4.605668, 4.416256, 4.244461, 4.223026, 3.864554, 
    3.448621, 3.079973, 2.834801, 2.803052, 2.791499, 2.260576, 1.729332, 
    1.570504,
  4.811379, 4.762827, 4.680954, 4.347826, 4.100862, 3.999176, 3.687927, 
    3.32552, 2.967337, 2.864635, 3.098063, 2.813399, 2.197472, 1.734627, 
    1.563886,
  4.414967, 4.245558, 4.285539, 4.283919, 4.012506, 3.307632, 3.026098, 
    3.495044, 4.192091, 4.583123, 4.663161, 4.582639, 4.57551, 4.435743, 
    4.401582,
  4.516161, 4.188236, 4.120398, 4.140047, 3.921227, 3.331203, 2.912615, 
    3.08831, 3.512074, 4.049805, 4.543633, 4.598105, 4.441675, 3.722807, 
    3.848525,
  4.625569, 4.321041, 4.047609, 4.039734, 3.925052, 3.129137, 3.168905, 
    2.896484, 3.048125, 3.175032, 3.593318, 3.598597, 3.025132, 2.837373, 
    3.0039,
  4.723565, 4.576776, 4.294813, 4.019278, 3.95665, 3.615541, 3.031278, 
    3.152301, 3.042416, 2.908989, 2.695403, 2.30009, 2.029528, 1.975778, 
    2.011995,
  4.87901, 4.691761, 4.544859, 4.224253, 3.968802, 3.834494, 3.658921, 
    2.807674, 2.850649, 3.00001, 2.534514, 2.126721, 2.044159, 1.979672, 
    1.85764,
  5.113337, 4.785267, 4.674979, 4.463229, 4.063819, 3.875198, 3.836566, 
    3.813633, 3.893507, 3.450371, 2.608101, 2.142285, 2.287817, 1.993064, 
    1.742166,
  5.18858, 4.916624, 4.715245, 4.598172, 4.285007, 4.020572, 3.896863, 
    3.870733, 3.659534, 3.378274, 2.654564, 2.330904, 2.337015, 1.787763, 
    1.70561,
  5.098687, 4.954908, 4.825487, 4.725836, 4.450336, 4.167477, 4.02104, 
    3.824595, 3.473926, 3.20758, 2.668751, 2.617899, 2.161348, 1.655714, 
    1.856305,
  4.953884, 4.911141, 4.882492, 4.870154, 4.625636, 4.331089, 4.090789, 
    3.759681, 3.33004, 3.051789, 2.694434, 2.736895, 1.762322, 1.666511, 
    2.048252,
  4.818166, 4.864913, 4.9547, 4.868351, 4.59973, 4.35433, 4.084484, 3.620577, 
    3.203837, 2.916997, 2.705067, 2.504984, 1.664377, 1.70743, 2.133906,
  5.6736, 4.8322, 4.09879, 3.735924, 3.761302, 3.808583, 3.95094, 4.126518, 
    4.320654, 4.409081, 4.530981, 4.381005, 4.221494, 3.804918, 3.705235,
  5.406042, 4.579321, 3.936615, 3.602873, 3.497998, 3.542281, 3.656673, 
    3.969458, 4.190757, 4.311966, 4.450965, 4.289163, 4.199808, 3.413573, 
    3.164793,
  5.165172, 4.534675, 3.806608, 3.542209, 3.396995, 2.997395, 3.331899, 
    3.553061, 3.911349, 4.089089, 4.247153, 4.040288, 3.484251, 2.803531, 
    2.463559,
  5.031785, 4.793203, 3.862227, 3.546145, 3.432588, 3.178956, 2.877356, 
    3.328128, 3.487261, 3.557319, 3.62248, 3.217436, 2.634983, 2.332423, 
    2.159322,
  4.887925, 4.961313, 3.983897, 3.707255, 3.500331, 3.242826, 3.104896, 
    2.752953, 2.757424, 3.108808, 2.961485, 2.642151, 2.416716, 2.271652, 
    2.266014,
  4.892609, 5.013134, 4.042079, 3.836771, 3.570464, 3.305173, 3.308405, 
    3.335117, 3.27935, 2.952898, 2.675306, 2.49768, 2.451561, 2.25436, 
    2.239486,
  5.055473, 4.901707, 4.185092, 4.01281, 3.803034, 3.573863, 3.503103, 
    3.582222, 3.323057, 2.950925, 2.646239, 2.460527, 2.432201, 2.160652, 
    2.270133,
  4.967281, 4.733292, 4.166725, 4.005882, 3.949874, 3.781265, 3.682922, 
    3.555652, 3.207311, 2.893041, 2.609589, 2.392647, 2.156059, 2.160277, 
    2.445982,
  4.983539, 4.790454, 4.301978, 4.028386, 4.018953, 3.930573, 3.724279, 
    3.511492, 3.105239, 2.820275, 2.571913, 2.405677, 1.982997, 2.253572, 
    2.508862,
  5.101469, 5.110323, 4.878252, 4.283519, 4.072145, 4.044328, 3.745172, 
    3.424295, 2.977711, 2.799271, 2.548256, 2.333367, 1.971895, 2.324802, 
    2.515325,
  5.578668, 5.700188, 5.49145, 4.846353, 4.03737, 3.409755, 3.304986, 
    3.527232, 3.730039, 3.87436, 4.046166, 4.238466, 4.247188, 3.941377, 
    3.63971,
  5.917355, 5.890029, 5.454083, 4.683604, 3.820315, 3.202346, 3.248356, 
    3.513533, 3.751759, 3.89466, 4.034509, 4.204752, 4.216075, 3.78777, 
    3.614526,
  6.167646, 5.923012, 5.229564, 4.383102, 3.568341, 2.70642, 3.094521, 
    3.410461, 3.71866, 3.849672, 4.001051, 4.143622, 4.130078, 3.91375, 
    3.666054,
  6.200689, 5.886169, 4.983715, 3.919598, 3.316943, 2.895566, 2.688074, 
    3.357868, 3.492447, 3.638675, 3.844729, 3.836329, 3.762557, 3.556139, 
    3.228072,
  6.123568, 5.75247, 4.632145, 3.508815, 3.079876, 2.909718, 3.06797, 
    2.876505, 2.916433, 3.350062, 3.32525, 3.218046, 3.210931, 3.012809, 
    2.799908,
  5.89535, 5.317086, 4.018509, 3.161405, 3.023418, 3.017085, 3.155224, 
    3.317487, 3.221817, 3.036239, 2.879379, 2.849613, 2.818059, 2.699452, 
    2.640376,
  5.423081, 4.699914, 3.461983, 3.215678, 3.301774, 3.246232, 3.138378, 
    3.015323, 2.86555, 2.755977, 2.669616, 2.66261, 2.617245, 2.568761, 
    2.565292,
  4.875417, 4.038808, 3.252717, 3.398293, 3.489477, 3.413893, 2.970086, 
    2.782963, 2.63767, 2.564069, 2.485185, 2.450767, 2.466121, 2.496407, 
    2.476894,
  4.236475, 3.557708, 3.239318, 3.472724, 3.615205, 3.223904, 2.814824, 
    2.64146, 2.506804, 2.429291, 2.36347, 2.334056, 2.383562, 2.485775, 
    2.531207,
  3.858091, 3.420936, 3.227978, 3.25424, 3.305098, 3.047801, 2.726119, 
    2.562827, 2.433318, 2.364078, 2.285831, 2.308423, 2.383764, 2.564965, 
    2.681748,
  6.566571, 6.394082, 6.221983, 6.083345, 5.92871, 5.727954, 5.329839, 
    4.882394, 4.39377, 3.980031, 3.805095, 3.737827, 3.717755, 3.740147, 
    3.736966,
  6.025455, 5.842585, 5.625525, 5.47738, 5.376709, 4.924475, 4.593893, 
    4.208993, 3.871921, 3.689896, 3.596832, 3.556458, 3.637998, 3.640441, 
    3.696462,
  5.619944, 5.23291, 4.972184, 4.858625, 4.629445, 3.853374, 3.97498, 
    3.702619, 3.519953, 3.432996, 3.406855, 3.479838, 3.584831, 3.75371, 
    3.752453,
  5.040122, 4.677696, 4.40824, 4.246851, 4.104469, 3.800057, 3.090053, 
    3.225787, 3.191686, 3.169546, 3.271096, 3.445558, 3.563534, 3.686462, 
    3.720522,
  4.382185, 4.176211, 3.975249, 3.701823, 3.372146, 3.1174, 2.96325, 
    2.422934, 2.495063, 2.970649, 3.144762, 3.409532, 3.541765, 3.653697, 
    3.635198,
  3.881597, 3.631793, 3.378858, 3.095346, 2.873553, 2.837304, 2.907876, 
    2.91888, 2.927742, 2.861904, 3.08581, 3.322628, 3.419713, 3.479536, 
    3.444937,
  3.489106, 3.233834, 3.036936, 2.955863, 2.902519, 2.850552, 2.824828, 
    2.761693, 2.718133, 2.789423, 3.009743, 3.158478, 3.249354, 3.262301, 
    3.160626,
  3.304432, 3.154606, 3.026441, 3.023003, 2.930138, 2.783443, 2.628417, 
    2.601584, 2.61611, 2.723729, 2.887239, 3.001466, 3.045335, 2.970647, 
    2.788564,
  3.451565, 3.289695, 3.108138, 2.909621, 2.759414, 2.541281, 2.437578, 
    2.462587, 2.522467, 2.641692, 2.757663, 2.822492, 2.798246, 2.674992, 
    2.5122,
  3.655856, 3.415322, 3.049843, 2.620046, 2.472304, 2.391181, 2.335299, 
    2.375347, 2.445888, 2.542122, 2.627212, 2.647234, 2.594083, 2.532649, 
    2.463595,
  3.52476, 3.260545, 2.982584, 2.76727, 2.813019, 2.915798, 2.970438, 
    3.051914, 3.274152, 3.374674, 3.489874, 3.607292, 3.70074, 3.74901, 
    3.821548,
  3.569757, 3.197821, 2.90956, 2.685239, 2.705106, 2.730148, 2.854319, 
    2.906057, 3.121275, 3.280648, 3.412292, 3.490592, 3.576244, 3.461438, 
    3.548976,
  3.856027, 3.321713, 3.010742, 2.763719, 2.667698, 2.46411, 2.692753, 
    2.748455, 2.869939, 3.023514, 3.174401, 3.299659, 3.343775, 3.400768, 
    3.449331,
  3.978801, 3.406958, 3.080614, 2.811256, 2.678703, 2.604814, 2.4096, 
    2.590033, 2.681628, 2.846693, 3.006834, 3.183663, 3.195076, 3.260994, 
    3.325349,
  3.994869, 3.417119, 3.017407, 2.828505, 2.71642, 2.582376, 2.575509, 
    2.204797, 2.225474, 2.726057, 2.897777, 3.089916, 3.168605, 3.201529, 
    3.222541,
  4.051609, 3.466769, 2.961959, 2.783466, 2.724686, 2.585469, 2.53874, 
    2.535919, 2.611018, 2.800527, 2.986622, 3.115205, 3.161571, 3.191586, 
    3.207307,
  4.131752, 3.553211, 2.95605, 2.703845, 2.717156, 2.61382, 2.571231, 
    2.589235, 2.705567, 2.896123, 3.010824, 3.094533, 3.1652, 3.213937, 
    3.302652,
  4.226844, 3.652373, 3.01931, 2.596182, 2.610683, 2.621669, 2.584391, 
    2.634647, 2.683481, 2.826039, 2.974296, 3.084124, 3.167696, 3.216861, 
    3.272968,
  4.338632, 3.756764, 3.125925, 2.507779, 2.365034, 2.445173, 2.543603, 
    2.646354, 2.689242, 2.769266, 2.875472, 2.979288, 3.056154, 3.091675, 
    3.034945,
  4.511607, 3.908036, 3.241445, 2.450047, 2.165372, 2.290308, 2.457994, 
    2.616735, 2.702, 2.757297, 2.807566, 2.873109, 2.921968, 2.926346, 
    2.942821,
  4.880228, 4.061924, 3.250276, 2.879734, 2.808273, 2.588785, 2.491156, 
    2.448638, 2.5301, 2.61546, 2.651269, 2.704204, 2.738046, 2.752957, 
    2.790883,
  5.388565, 4.336475, 3.327461, 2.842534, 2.767249, 2.596524, 2.527971, 
    2.454487, 2.578045, 2.730847, 2.807197, 2.893487, 2.898207, 2.796845, 
    2.891287,
  5.957193, 4.802399, 3.62321, 2.855274, 2.70134, 2.434325, 2.537684, 
    2.517222, 2.617072, 2.778411, 2.896821, 2.99633, 3.009549, 3.062157, 
    3.157583,
  6.63689, 5.561844, 4.151696, 2.953891, 2.683599, 2.618904, 2.387594, 
    2.553355, 2.618728, 2.806813, 2.939528, 3.059396, 3.125435, 3.189662, 
    3.250767,
  7.495402, 6.382266, 4.811173, 3.259557, 2.653665, 2.653653, 2.625298, 
    2.212265, 2.216083, 2.795746, 2.981572, 3.092749, 3.199535, 3.263013, 
    3.289651,
  8.4103, 7.349167, 5.697266, 3.867262, 2.594417, 2.574501, 2.6803, 2.667006, 
    2.741254, 2.841615, 3.021846, 3.110632, 3.208551, 3.262067, 3.25928,
  9.288527, 8.330306, 6.822595, 4.748635, 2.797737, 2.472472, 2.684034, 
    2.758147, 2.866153, 2.965612, 3.045752, 3.12224, 3.18886, 3.224818, 
    3.191996,
  10.00479, 9.307317, 7.932907, 5.852784, 3.366228, 2.353397, 2.568934, 
    2.734813, 2.828465, 2.964168, 3.057409, 3.126645, 3.150371, 3.121669, 
    3.020566,
  10.44412, 10.06073, 8.931305, 7.086571, 4.557563, 2.251903, 2.398862, 
    2.701685, 2.817322, 2.908893, 2.985504, 3.027937, 3.020497, 2.963704, 
    2.853981,
  10.70363, 10.47701, 9.716398, 8.171358, 5.811597, 2.626175, 2.193741, 
    2.56512, 2.751893, 2.849892, 2.91501, 2.950022, 2.947766, 2.917998, 
    2.862457,
  8.829076, 8.522467, 6.619843, 3.478814, 2.336532, 2.43772, 2.436054, 
    2.482452, 2.570319, 2.546747, 2.506133, 2.452698, 2.225626, 2.152548, 
    2.135924,
  8.82708, 8.561148, 6.44213, 3.370943, 2.319877, 2.434659, 2.500803, 
    2.536109, 2.625987, 2.65125, 2.634334, 2.571521, 2.39464, 2.151715, 
    2.133327,
  8.732321, 8.516495, 6.411767, 3.539211, 2.336123, 2.246545, 2.507646, 
    2.587589, 2.634421, 2.651504, 2.614925, 2.519241, 2.413035, 2.321375, 
    2.330253,
  8.555111, 8.387134, 6.429745, 3.801525, 2.456189, 2.481005, 2.365744, 
    2.636358, 2.648111, 2.701851, 2.720182, 2.641488, 2.596171, 2.631057, 
    2.714754,
  8.237911, 8.104054, 6.53535, 4.115181, 2.518781, 2.605692, 2.655588, 
    2.253817, 2.303957, 2.813128, 2.951024, 2.960482, 2.963809, 3.009112, 
    3.076338,
  7.741168, 7.643981, 6.648442, 4.409588, 2.607176, 2.601309, 2.775859, 
    2.81887, 2.848945, 2.915422, 3.018896, 3.048766, 3.051908, 3.064706, 
    3.060853,
  7.162722, 7.042535, 6.726081, 4.632854, 2.857345, 2.597953, 2.726518, 
    2.801547, 2.870635, 2.904655, 2.935031, 2.969415, 2.989161, 3.013506, 
    3.054167,
  6.635352, 6.44396, 6.601757, 4.716166, 3.060752, 2.602897, 2.635028, 
    2.692919, 2.729913, 2.775643, 2.807064, 2.844414, 2.898032, 2.975948, 
    3.083313,
  6.219466, 5.923695, 6.314904, 4.813567, 3.259052, 2.474113, 2.540073, 
    2.601394, 2.627559, 2.650989, 2.692029, 2.761119, 2.858243, 2.984349, 
    3.141331,
  5.956964, 5.638827, 5.885926, 4.788693, 3.27936, 2.382991, 2.460022, 
    2.516754, 2.559596, 2.62448, 2.695318, 2.773008, 2.884063, 3.035313, 
    3.221332,
  3.769207, 3.010783, 2.435681, 2.3113, 2.347379, 2.313058, 2.245164, 
    2.259884, 2.245535, 2.187663, 2.179, 2.110739, 2.044801, 2.000051, 
    1.994117,
  3.448986, 2.833715, 2.528011, 2.54518, 2.561914, 2.46416, 2.390204, 
    2.294704, 2.253304, 2.246685, 2.203553, 2.139053, 2.043957, 1.89423, 
    1.938874,
  3.313766, 2.815188, 2.663935, 2.742287, 2.760252, 2.487127, 2.572355, 
    2.503, 2.408482, 2.341049, 2.215662, 2.106463, 2.019144, 2.000819, 
    1.995216,
  3.387639, 3.015616, 2.848655, 2.870998, 2.929149, 2.874936, 2.603025, 
    2.657244, 2.584975, 2.591049, 2.532078, 2.351456, 2.18548, 2.076627, 
    2.02902,
  3.428515, 3.161292, 3.072189, 2.959124, 3.003769, 3.001245, 2.942407, 
    2.476342, 2.401444, 2.694059, 2.702592, 2.656812, 2.520684, 2.339561, 
    2.214261,
  3.386173, 3.205769, 3.111996, 3.055039, 3.037946, 3.029613, 3.02663, 
    2.928463, 2.814015, 2.845805, 2.852671, 2.790308, 2.732647, 2.610397, 
    2.447706,
  3.433589, 3.308647, 3.199578, 3.13027, 3.105227, 3.005423, 3.05438, 
    3.09415, 3.129179, 3.157641, 3.108537, 3.020395, 2.92643, 2.845757, 
    2.744349,
  3.432881, 3.350151, 3.24193, 3.149458, 3.077819, 2.982639, 3.009167, 
    3.11003, 3.2036, 3.281452, 3.326939, 3.285578, 3.171824, 3.062088, 
    2.971752,
  3.408216, 3.301356, 3.135415, 3.033203, 2.971058, 2.930531, 2.993231, 
    3.071983, 3.159569, 3.292459, 3.398565, 3.505725, 3.485301, 3.370403, 
    3.269415,
  3.230593, 3.075054, 2.88378, 2.789258, 2.843711, 2.957877, 3.026604, 
    3.024158, 3.040415, 3.122929, 3.306726, 3.494341, 3.648538, 3.663981, 
    3.573052,
  3.110829, 3.124996, 3.082316, 3.026596, 2.956512, 2.736509, 2.57082, 
    2.418769, 2.319696, 2.111153, 2.050189, 2.112633, 2.246897, 2.455003, 
    2.840005,
  3.326763, 3.261224, 3.165091, 3.089528, 2.993697, 2.774766, 2.629182, 
    2.421319, 2.309417, 2.188158, 2.033633, 2.054104, 2.154019, 2.18776, 
    2.53102,
  3.50878, 3.408894, 3.278797, 3.109878, 2.995192, 2.66005, 2.692295, 
    2.535909, 2.379632, 2.308799, 2.066683, 1.979145, 2.042005, 2.154443, 
    2.385636,
  3.567247, 3.493462, 3.358724, 3.096745, 2.996511, 2.852952, 2.562161, 
    2.617999, 2.468917, 2.377861, 2.204569, 1.994933, 1.970636, 2.039939, 
    2.198588,
  3.599338, 3.51632, 3.379548, 3.10142, 2.918633, 2.840181, 2.776306, 
    2.358419, 2.233269, 2.504625, 2.253693, 2.087522, 1.955859, 1.96356, 
    2.07249,
  3.584497, 3.528516, 3.322725, 3.065435, 2.86184, 2.725006, 2.728231, 
    2.731059, 2.702751, 2.6853, 2.438711, 2.201853, 2.011493, 1.954312, 
    1.962367,
  3.551021, 3.405365, 3.268064, 3.013203, 2.81654, 2.601059, 2.638374, 
    2.762546, 2.842315, 2.905492, 2.762199, 2.37037, 2.147954, 2.011114, 
    1.945638,
  3.406328, 3.254358, 3.018402, 2.830195, 2.635802, 2.447572, 2.487075, 
    2.643857, 2.80375, 2.868329, 2.925482, 2.712742, 2.36283, 2.149333, 
    2.012757,
  3.220894, 3.019503, 2.717193, 2.453267, 2.247628, 2.213274, 2.345506, 
    2.529446, 2.678129, 2.816826, 2.882972, 2.930212, 2.669406, 2.369013, 
    2.167147,
  2.972429, 2.666237, 2.314812, 2.01875, 1.930109, 1.968033, 2.133614, 
    2.370121, 2.52512, 2.696371, 2.799011, 2.923142, 2.948766, 2.667836, 
    2.388793,
  2.846477, 2.759174, 2.640351, 2.502876, 2.395095, 2.210621, 2.130596, 
    2.090662, 2.110445, 2.071746, 2.040877, 2.019826, 1.988874, 1.999921, 
    2.05494,
  2.982183, 2.724228, 2.477839, 2.28416, 2.173656, 2.001037, 2.000643, 
    2.010682, 2.114316, 2.182004, 2.121616, 2.06439, 2.010911, 1.884276, 
    1.955582,
  3.232942, 2.721133, 2.346227, 2.076553, 1.955758, 1.708745, 1.863816, 
    2.037545, 2.19801, 2.314792, 2.241054, 2.118373, 2.017739, 1.977366, 
    2.029522,
  3.087285, 2.728932, 2.268313, 1.936105, 1.81941, 1.8148, 1.681619, 1.99846, 
    2.209213, 2.337719, 2.27144, 2.110063, 2.001844, 1.958975, 2.035665,
  2.943214, 2.571918, 2.188862, 1.875028, 1.798964, 1.830879, 1.89813, 
    1.747708, 1.905576, 2.283992, 2.242412, 2.097089, 1.979593, 1.937582, 
    2.052426,
  2.737466, 2.412143, 2.067032, 1.859682, 1.807087, 1.856395, 1.951075, 
    2.04918, 2.179014, 2.277509, 2.259531, 2.072081, 1.974901, 1.922315, 
    2.020906,
  2.57669, 2.299641, 2.062486, 1.875569, 1.863455, 1.891137, 2.014532, 
    2.117981, 2.227136, 2.366571, 2.34381, 2.057253, 1.93281, 1.887803, 
    1.951528,
  2.398163, 2.183104, 1.979277, 1.887526, 1.784628, 1.828946, 2.016291, 
    2.126958, 2.205227, 2.317598, 2.312735, 2.137713, 1.940842, 1.836005, 
    1.882163,
  2.266284, 2.049253, 1.838294, 1.625739, 1.547366, 1.650446, 1.882907, 
    2.092, 2.17552, 2.268677, 2.325882, 2.2423, 1.996346, 1.87944, 1.843564,
  2.029052, 1.736221, 1.529386, 1.38771, 1.42614, 1.494093, 1.649043, 
    1.921302, 2.107294, 2.191011, 2.301972, 2.318972, 2.142768, 1.947407, 
    1.868753,
  2.076421, 1.998398, 1.94734, 1.881371, 1.825163, 1.773653, 1.767228, 
    1.759212, 1.776778, 1.80317, 1.844281, 1.871463, 1.852174, 1.837133, 
    1.843576,
  1.85624, 1.755584, 1.706241, 1.694783, 1.686303, 1.607976, 1.6695, 
    1.652128, 1.678094, 1.731114, 1.786015, 1.837021, 1.862915, 1.773596, 
    1.808663,
  2.017216, 1.763986, 1.646494, 1.603018, 1.644269, 1.51706, 1.722607, 
    1.792399, 1.826356, 1.906797, 1.996935, 2.036763, 2.024253, 1.986026, 
    1.944438,
  2.263001, 2.018357, 1.833748, 1.613231, 1.661356, 1.749636, 1.668098, 
    1.887123, 1.971912, 2.110363, 2.170865, 2.186749, 2.15946, 2.091252, 
    1.997201,
  2.298739, 2.117794, 1.971173, 1.730795, 1.689718, 1.766279, 1.864036, 
    1.653082, 1.716928, 2.083221, 2.137702, 2.152522, 2.103267, 2.036233, 
    1.961098,
  2.385991, 2.19095, 2.049792, 1.839733, 1.724446, 1.67304, 1.777577, 
    1.860675, 1.935546, 2.052967, 2.120887, 2.103969, 2.072977, 1.960136, 
    1.88141,
  2.449023, 2.296716, 2.117816, 1.945772, 1.799524, 1.62769, 1.704942, 
    1.808863, 1.887429, 2.007162, 2.058381, 2.020459, 1.977486, 1.898849, 
    1.809708,
  2.449764, 2.301458, 2.141231, 2.034668, 1.857993, 1.6355, 1.614063, 
    1.697627, 1.748279, 1.826685, 1.870888, 1.91092, 1.90813, 1.859981, 
    1.798488,
  2.516356, 2.298128, 2.187455, 2.03077, 1.836428, 1.710447, 1.637564, 
    1.653637, 1.677107, 1.719584, 1.761242, 1.808556, 1.819249, 1.813208, 
    1.787113,
  2.458666, 2.308625, 2.143175, 2.039037, 1.995348, 1.885159, 1.76299, 
    1.722137, 1.650207, 1.621682, 1.646061, 1.704975, 1.754914, 1.769215, 
    1.765567,
  1.420703, 1.353775, 1.32543, 1.299149, 1.286863, 1.281124, 1.308308, 
    1.345733, 1.418541, 1.505525, 1.773857, 2.171446, 2.506041, 2.776565, 
    3.03194,
  1.489696, 1.491012, 1.492002, 1.480168, 1.466771, 1.398054, 1.43246, 
    1.412297, 1.412752, 1.458634, 1.523265, 1.635356, 1.80482, 1.959493, 
    2.244585,
  2.312932, 2.287694, 2.218882, 2.119734, 2.020513, 1.729312, 1.807248, 
    1.834582, 1.761836, 1.697099, 1.671289, 1.665632, 1.657225, 1.706604, 
    1.820893,
  2.984789, 3.09348, 3.170905, 2.964852, 2.802545, 2.591587, 2.190241, 
    2.221341, 2.192952, 2.189632, 2.111871, 2.012828, 1.918792, 1.838224, 
    1.773772,
  3.228428, 3.517589, 3.670171, 3.520744, 3.362681, 3.134801, 2.878339, 
    2.263198, 2.084151, 2.35991, 2.309689, 2.207591, 2.11491, 2.012287, 
    1.904261,
  3.604748, 4.009013, 4.010974, 3.81466, 3.608803, 3.301901, 2.958404, 
    2.637395, 2.435998, 2.303071, 2.198479, 2.14606, 2.120923, 2.069363, 
    1.98345,
  4.180996, 4.304989, 4.151465, 3.854073, 3.573845, 3.190729, 2.792316, 
    2.447033, 2.17118, 1.972822, 1.86706, 1.862778, 1.918977, 1.978665, 
    1.961115,
  4.524554, 4.421459, 4.019697, 3.669724, 3.340418, 2.905283, 2.450804, 
    2.095869, 1.859344, 1.707279, 1.625009, 1.602427, 1.660802, 1.781711, 
    1.859268,
  4.646818, 4.291821, 3.872576, 3.501789, 3.068916, 2.539515, 2.061903, 
    1.802211, 1.634458, 1.524523, 1.4707, 1.464097, 1.512606, 1.613001, 
    1.716207,
  4.582055, 4.201317, 3.744541, 3.27928, 2.799306, 2.175695, 1.733701, 
    1.524693, 1.420178, 1.372605, 1.364154, 1.38444, 1.44099, 1.524399, 
    1.595708,
  2.556095, 2.657556, 2.896948, 3.438415, 3.519482, 3.221019, 2.71454, 
    2.2149, 1.921678, 1.672787, 1.491373, 1.400603, 1.344443, 1.301999, 
    1.318503,
  2.782409, 2.945051, 3.45862, 4.386598, 4.550415, 4.274088, 4.067047, 
    3.623225, 3.182746, 2.846799, 2.566788, 2.311371, 2.056621, 1.723405, 
    1.503854,
  2.907382, 3.292214, 4.380324, 5.356662, 5.342598, 4.650587, 4.590822, 
    4.069533, 3.527228, 3.192793, 2.976145, 2.785742, 2.603262, 2.430816, 
    2.242567,
  3.049744, 4.227799, 5.405537, 5.732276, 5.584029, 5.010503, 3.682801, 
    3.279019, 2.968798, 2.79049, 2.672503, 2.592587, 2.540253, 2.495643, 
    2.413271,
  3.95765, 5.384482, 5.797081, 5.707027, 4.962571, 4.097747, 3.429935, 
    2.464427, 2.124611, 2.221017, 2.11019, 2.030499, 2.037008, 2.088742, 
    2.174095,
  5.397937, 5.824794, 5.820663, 5.08432, 4.285778, 3.739866, 3.200961, 
    2.658117, 2.24409, 1.913854, 1.665141, 1.531103, 1.517061, 1.615103, 
    1.781338,
  5.801974, 5.772429, 5.21175, 4.436633, 3.895373, 3.286866, 2.620435, 
    2.022883, 1.632309, 1.438587, 1.373342, 1.341714, 1.316523, 1.334649, 
    1.460963,
  5.772514, 5.278223, 4.624073, 3.926656, 3.256294, 2.3665, 1.665128, 
    1.429521, 1.399367, 1.384073, 1.362227, 1.324566, 1.271652, 1.22972, 
    1.284407,
  5.355798, 4.800439, 4.050297, 3.26394, 2.405552, 1.601116, 1.381286, 
    1.412254, 1.456406, 1.401641, 1.350849, 1.275458, 1.190238, 1.113062, 
    1.135731,
  4.952781, 4.175662, 3.42356, 2.531712, 1.734504, 1.374139, 1.395324, 
    1.483148, 1.459595, 1.387315, 1.298667, 1.198604, 1.093858, 1.002226, 
    1.029505,
  2.441555, 1.990762, 1.827558, 2.486516, 3.979226, 5.141922, 5.387837, 
    4.987765, 4.114708, 3.367419, 2.951994, 2.712827, 2.500415, 2.326627, 
    2.365986,
  1.920681, 1.819652, 2.087126, 3.448901, 4.95458, 5.485059, 5.391809, 
    4.490245, 3.719285, 3.336783, 3.121652, 3.00179, 2.899051, 2.698376, 
    2.718704,
  1.961599, 2.126989, 3.044084, 4.877547, 5.657837, 5.0377, 4.281178, 
    3.53372, 3.108821, 2.834859, 2.697453, 2.633745, 2.552809, 2.507519, 
    2.482375,
  2.067237, 2.968849, 4.883065, 5.888017, 5.629153, 4.350983, 2.835558, 
    2.451467, 2.401713, 2.375511, 2.335623, 2.296413, 2.276663, 2.253982, 
    2.225638,
  2.69413, 4.868754, 6.04656, 5.651599, 4.139098, 2.618182, 2.116895, 
    1.564419, 1.555082, 1.933993, 1.993035, 2.006733, 2.042443, 2.072263, 
    2.10038,
  5.144758, 6.226798, 5.94558, 4.303243, 2.733946, 1.798383, 1.561481, 
    1.569488, 1.609196, 1.635727, 1.649391, 1.665805, 1.689448, 1.729373, 
    1.768419,
  6.253769, 6.075163, 4.609441, 2.910388, 2.019016, 1.586165, 1.522894, 
    1.561906, 1.561165, 1.524949, 1.480495, 1.458638, 1.458843, 1.464043, 
    1.472226,
  6.146481, 4.719361, 3.152196, 2.176661, 1.744357, 1.573883, 1.613206, 
    1.621745, 1.577871, 1.503938, 1.480352, 1.46769, 1.46435, 1.45126, 
    1.431306,
  5.220062, 3.511931, 2.31134, 1.711178, 1.564558, 1.664666, 1.692898, 
    1.645878, 1.527149, 1.485401, 1.481173, 1.474006, 1.437443, 1.414235, 
    1.374328,
  4.204216, 2.485511, 1.739759, 1.535974, 1.678232, 1.738003, 1.713733, 
    1.567918, 1.48786, 1.462012, 1.44554, 1.451871, 1.446566, 1.388752, 
    1.285201,
  3.125657, 2.875783, 2.855021, 2.792567, 2.726227, 2.828443, 3.32281, 
    3.874795, 3.999868, 3.457875, 2.699031, 2.068245, 1.665916, 1.519485, 
    1.571855,
  3.413287, 3.080347, 2.882623, 2.728346, 2.796348, 3.176252, 3.852625, 
    4.017146, 3.578466, 2.829041, 2.138147, 1.739688, 1.578122, 1.446977, 
    1.466278,
  3.778055, 3.326323, 2.89758, 2.834867, 3.332708, 3.493816, 4.008098, 
    3.722039, 2.953863, 2.237406, 1.80457, 1.659171, 1.599808, 1.549998, 
    1.486013,
  3.747867, 3.606776, 3.471741, 3.804992, 4.225631, 4.3119, 3.536796, 
    3.003539, 2.422595, 2.031354, 1.770616, 1.658575, 1.602008, 1.530496, 
    1.45578,
  3.387079, 3.462805, 4.010755, 4.482351, 4.498254, 4.064336, 3.384737, 
    2.24673, 1.804011, 1.873159, 1.726601, 1.616544, 1.525204, 1.450308, 
    1.422984,
  3.152855, 3.846363, 4.531938, 4.755168, 4.405908, 3.789533, 3.098554, 
    2.459226, 1.978121, 1.699599, 1.590123, 1.50945, 1.454319, 1.427505, 
    1.419155,
  3.646114, 4.495758, 4.967306, 4.690514, 4.158626, 3.418138, 2.686435, 
    2.104417, 1.769825, 1.642321, 1.552088, 1.469141, 1.435001, 1.420221, 
    1.413929,
  4.948198, 5.220511, 5.015974, 4.423413, 3.743658, 2.779031, 2.139204, 
    1.799207, 1.655634, 1.546221, 1.479763, 1.437928, 1.425357, 1.424932, 
    1.410421,
  6.360097, 5.949055, 5.050315, 4.010471, 3.043747, 2.292472, 1.874036, 
    1.702215, 1.575073, 1.498431, 1.451175, 1.42506, 1.433933, 1.412395, 
    1.383479,
  5.904776, 5.638301, 4.501854, 3.275488, 2.415523, 1.932119, 1.725145, 
    1.594455, 1.485816, 1.424103, 1.39959, 1.422099, 1.419599, 1.389737, 
    1.341172,
  5.168321, 4.817051, 4.481972, 4.167191, 3.736692, 3.361758, 3.16499, 
    3.054331, 2.969736, 2.977846, 3.118592, 3.263062, 3.197662, 2.963208, 
    2.775669,
  4.863168, 4.607527, 4.173654, 3.817303, 3.485397, 3.245363, 3.130176, 
    3.046452, 3.029975, 3.142521, 3.224994, 3.214293, 3.050578, 2.768167, 
    2.68215,
  4.507042, 4.448635, 4.003628, 3.578405, 3.216963, 2.733297, 2.970574, 
    3.112635, 3.204816, 3.251652, 3.243315, 3.121494, 2.965618, 2.843199, 
    2.6959,
  4.191165, 4.437346, 4.123668, 3.591479, 3.190908, 2.87754, 2.663109, 
    2.99472, 3.216565, 3.340365, 3.291511, 3.12301, 2.957256, 2.773854, 
    2.544175,
  3.897717, 4.391799, 4.461515, 3.998701, 3.450433, 3.170244, 2.993263, 
    2.572272, 2.586475, 3.138443, 3.203408, 3.017689, 2.819775, 2.592502, 
    2.357423,
  3.729333, 4.193415, 4.543295, 4.425178, 3.942323, 3.510928, 3.336613, 
    3.197483, 3.228848, 3.239036, 3.055108, 2.858047, 2.652899, 2.400061, 
    2.10672,
  3.727055, 4.126706, 4.469781, 4.568121, 4.365191, 4.043424, 3.852109, 
    3.745034, 3.521849, 3.194991, 2.939916, 2.67498, 2.351029, 1.997527, 
    1.712812,
  3.732136, 4.09547, 4.331801, 4.484864, 4.471096, 4.435165, 4.30754, 
    4.032444, 3.619797, 3.192614, 2.723557, 2.252337, 1.854811, 1.561607, 
    1.416125,
  4.39115, 4.445485, 4.463216, 4.528487, 4.642192, 4.711847, 4.469737, 
    3.949628, 3.346714, 2.721841, 2.139559, 1.667788, 1.41187, 1.341276, 
    1.344826,
  4.894297, 5.446766, 5.449596, 5.230968, 4.982625, 4.52052, 3.865992, 
    3.177341, 2.452089, 1.813657, 1.42274, 1.266946, 1.29019, 1.35331, 
    1.383783,
  3.763159, 4.066358, 4.323495, 4.515206, 4.681759, 4.757617, 4.806371, 
    4.834226, 4.823691, 4.62716, 4.295579, 3.799523, 3.150341, 2.664243, 
    2.410929,
  4.120901, 4.379006, 4.575004, 4.739347, 4.787203, 4.832919, 4.860508, 
    4.816553, 4.691329, 4.536241, 4.310521, 3.981466, 3.450163, 2.776039, 
    2.492051,
  4.390147, 4.456025, 4.671365, 4.862614, 4.90824, 4.457896, 4.748772, 
    4.68233, 4.550351, 4.389715, 4.222331, 4.005437, 3.67807, 3.170812, 
    2.770506,
  4.28099, 4.168594, 4.659686, 4.915593, 4.91349, 4.685968, 4.090189, 
    4.327584, 4.298345, 4.179272, 4.067008, 3.911374, 3.705392, 3.446139, 
    3.147988,
  4.059531, 4.008488, 4.682423, 4.855521, 4.750979, 4.61612, 4.24584, 
    3.486601, 3.360416, 3.912529, 3.892141, 3.768223, 3.615056, 3.416986, 
    3.26923,
  4.040253, 4.03474, 4.537928, 4.716491, 4.632745, 4.482243, 4.219835, 
    3.765679, 3.663936, 3.714953, 3.608074, 3.504822, 3.415647, 3.328675, 
    3.309894,
  4.097121, 4.239345, 4.441892, 4.622873, 4.484035, 4.276056, 3.923113, 
    3.646496, 3.459456, 3.267703, 3.170903, 3.147891, 3.178165, 3.222758, 
    3.215952,
  4.262802, 4.332946, 4.458386, 4.485265, 4.33369, 4.06626, 3.804883, 
    3.511234, 3.292163, 3.240011, 3.243615, 3.24236, 3.130532, 2.934258, 
    2.695883,
  4.407277, 4.27818, 4.292481, 4.242537, 4.090609, 3.91223, 3.724061, 
    3.532632, 3.388159, 3.177269, 2.977142, 2.623266, 2.156792, 1.812069, 
    1.611999,
  4.2537, 4.149518, 3.909172, 3.705539, 3.510824, 3.276522, 2.993136, 
    2.665421, 2.341967, 1.996677, 1.656106, 1.459364, 1.410735, 1.400434, 
    1.385034,
  4.582625, 4.537945, 4.459937, 4.344291, 4.292338, 4.235503, 4.134548, 
    3.985388, 3.827355, 3.667198, 3.752208, 4.031096, 4.234683, 4.243951, 
    4.393033,
  4.508286, 4.429366, 4.3007, 4.233129, 4.219345, 4.159282, 4.162744, 
    4.055068, 3.891069, 3.776588, 3.788456, 3.955165, 4.154433, 4.054345, 
    4.023181,
  4.262607, 4.1361, 4.047577, 3.99014, 4.030555, 3.681954, 3.928684, 3.95666, 
    3.862521, 3.790733, 3.778681, 3.883493, 4.048066, 4.198951, 4.112059,
  3.93993, 3.883201, 3.834888, 3.715624, 3.808176, 3.901461, 3.495225, 
    3.623025, 3.627804, 3.625225, 3.647299, 3.734085, 3.909628, 4.130099, 
    4.180693,
  3.723007, 3.672268, 3.557185, 3.402337, 3.510572, 3.702385, 3.729735, 
    3.069475, 2.988606, 3.559487, 3.606655, 3.646336, 3.798063, 3.977606, 
    4.144678,
  3.49135, 3.448149, 3.28808, 3.139749, 3.2279, 3.412003, 3.569619, 3.543015, 
    3.450726, 3.46836, 3.521413, 3.572208, 3.613893, 3.737867, 3.843696,
  3.291741, 3.198928, 3.031772, 2.839041, 2.847923, 2.912408, 3.063421, 
    3.178418, 3.227898, 3.244405, 3.233448, 3.235919, 3.258704, 3.312301, 
    3.382384,
  3.17201, 2.982378, 2.747434, 2.508388, 2.394092, 2.457709, 2.566898, 
    2.608723, 2.673464, 2.700805, 2.682453, 2.659291, 2.648, 2.66895, 2.729785,
  3.136897, 2.871837, 2.505146, 2.053057, 1.789423, 1.860275, 1.997856, 
    2.056608, 2.025125, 1.92849, 1.799732, 1.710942, 1.632236, 1.562481, 
    1.519657,
  3.264364, 2.921113, 2.478157, 1.914283, 1.574698, 1.444906, 1.48975, 
    1.506949, 1.468158, 1.411397, 1.334562, 1.285054, 1.266586, 1.278486, 
    1.284826,
  3.463579, 3.280653, 3.194951, 3.118724, 3.081979, 3.049367, 2.96253, 
    2.857233, 2.925427, 3.067434, 3.271471, 3.468799, 3.53483, 3.492618, 
    3.437011,
  3.288643, 3.199677, 3.174181, 3.085023, 2.99934, 2.850084, 2.792027, 
    2.664815, 2.746684, 2.98534, 3.216537, 3.378711, 3.462488, 3.295506, 
    3.300053,
  3.267629, 3.247201, 3.234632, 3.09758, 2.926214, 2.481366, 2.512413, 
    2.547056, 2.634884, 2.798263, 2.962851, 3.063161, 3.142516, 3.209182, 
    3.241966,
  3.37411, 3.395882, 3.442416, 3.235406, 2.951078, 2.618943, 2.215847, 
    2.287322, 2.355663, 2.453692, 2.556033, 2.613159, 2.707016, 2.798765, 
    2.887311,
  3.820287, 3.691689, 3.619812, 3.347472, 2.918151, 2.544782, 2.285371, 
    1.806506, 1.744205, 2.087563, 2.188375, 2.21375, 2.26963, 2.35509, 
    2.491706,
  4.388008, 4.116472, 3.895108, 3.614598, 2.929141, 2.326619, 1.996693, 
    1.897059, 1.817607, 1.812227, 1.875388, 1.916544, 1.972713, 2.052089, 
    2.19442,
  4.963189, 4.743766, 4.569963, 4.151511, 2.767774, 1.907633, 1.68333, 
    1.639721, 1.6125, 1.580809, 1.586835, 1.630733, 1.687488, 1.763379, 
    1.909094,
  5.23208, 5.237783, 5.172671, 3.999026, 2.251223, 1.498665, 1.509237, 
    1.457776, 1.410951, 1.383471, 1.389145, 1.435327, 1.464489, 1.486025, 
    1.566325,
  5.326402, 5.252702, 4.757375, 3.313448, 1.698218, 1.389645, 1.451217, 
    1.44011, 1.369883, 1.311556, 1.291569, 1.307631, 1.307714, 1.295569, 
    1.325701,
  4.974945, 4.594935, 3.975355, 2.57353, 1.587396, 1.370354, 1.40705, 
    1.390373, 1.319901, 1.265059, 1.22466, 1.193246, 1.1671, 1.130488, 1.13964,
  5.209971, 5.191075, 4.991117, 4.669372, 4.387869, 4.250992, 4.18965, 
    4.040911, 3.7259, 3.325316, 3.019767, 2.784122, 2.517431, 2.312912, 
    2.212768,
  4.211773, 4.730039, 4.784328, 4.570959, 4.261535, 4.014761, 3.958888, 
    3.847826, 3.584133, 3.322363, 3.081559, 2.879859, 2.649971, 2.319629, 
    2.181489,
  3.347034, 3.686962, 4.060645, 4.065914, 3.765645, 3.012247, 3.302559, 
    3.333231, 3.209174, 3.055653, 2.889526, 2.695604, 2.480784, 2.260233, 2.06,
  3.867169, 3.620638, 3.590192, 3.447243, 3.255411, 3.030537, 2.839547, 
    3.22749, 3.244277, 2.961369, 2.607136, 2.28606, 2.038443, 1.858533, 
    1.730654,
  4.618832, 4.242656, 4.117545, 3.894231, 3.775012, 3.916531, 3.90499, 
    2.843127, 2.273666, 2.034468, 1.693755, 1.487626, 1.400744, 1.364318, 
    1.358211,
  5.169518, 4.848168, 4.480595, 4.027264, 3.646996, 3.328207, 2.632135, 
    1.98244, 1.492396, 1.241535, 1.147377, 1.134308, 1.143898, 1.140839, 
    1.138159,
  4.490018, 4.065812, 3.380275, 2.688323, 2.040157, 1.605227, 1.240401, 
    1.089595, 1.064728, 1.060011, 1.069848, 1.06964, 1.058052, 0.9981198, 
    0.9639659,
  3.423694, 2.931065, 2.370043, 1.75601, 1.298744, 1.057997, 1.045731, 
    1.053096, 1.062606, 1.058314, 1.033004, 0.9999486, 0.9387261, 0.8755738, 
    0.8522716,
  2.427488, 2.041675, 1.672317, 1.336043, 1.123401, 1.116266, 1.111388, 
    1.108041, 1.095294, 1.071307, 1.032477, 0.9766001, 0.8967516, 0.8200499, 
    0.7766007,
  1.835746, 1.586965, 1.307075, 1.150169, 1.148537, 1.15038, 1.163673, 
    1.190304, 1.184809, 1.154112, 1.120064, 1.044962, 0.9356646, 0.830372, 
    0.756759,
  4.85899, 4.995584, 5.754312, 6.849527, 8.05136, 8.718051, 9.050338, 
    9.210615, 9.095597, 8.640331, 8.225248, 7.767088, 7.127757, 6.424788, 
    5.769371,
  4.685395, 4.743443, 5.16466, 5.862791, 6.58152, 7.204175, 7.707061, 
    8.038175, 8.145944, 8.020989, 7.749405, 7.420928, 6.907535, 6.000842, 
    5.459371,
  4.28351, 4.329667, 4.446549, 4.908632, 5.368392, 5.410052, 6.175375, 
    6.495432, 6.736487, 6.788753, 6.630639, 6.337442, 5.923739, 5.390963, 
    4.870706,
  3.926262, 3.869085, 3.795167, 3.771776, 3.983291, 4.139647, 4.104611, 
    4.830731, 4.887048, 4.914227, 4.829578, 4.604054, 4.228906, 3.794625, 
    3.326645,
  3.782562, 3.648348, 3.472153, 3.277526, 3.337713, 3.611979, 3.579975, 
    3.005352, 3.019072, 3.378108, 3.112404, 2.778081, 2.479717, 2.219335, 
    1.996887,
  3.189826, 3.071246, 2.854862, 2.517003, 2.314188, 2.356545, 2.61056, 
    2.556443, 2.322202, 1.990936, 1.733255, 1.583053, 1.468704, 1.412715, 
    1.349567,
  2.400585, 2.037685, 1.60104, 1.194191, 1.069434, 1.032634, 1.206529, 
    1.405023, 1.442328, 1.318211, 1.246101, 1.211725, 1.209012, 1.221626, 
    1.220624,
  2.614167, 2.293391, 2.034833, 1.773186, 1.44244, 1.180829, 1.180718, 
    1.211566, 1.246187, 1.263725, 1.271925, 1.287835, 1.311527, 1.337386, 
    1.354746,
  3.067219, 2.816547, 2.551878, 2.233801, 1.882716, 1.621117, 1.487236, 
    1.450665, 1.454342, 1.464668, 1.490301, 1.545624, 1.610962, 1.641634, 
    1.63297,
  3.658109, 3.371086, 3.029705, 2.560996, 2.189166, 2.009431, 1.938988, 
    1.899911, 1.869777, 1.83514, 1.857691, 1.9173, 1.948482, 1.935779, 
    1.854681,
  2.880343, 2.980473, 4.452437, 6.141675, 7.174526, 7.537774, 7.737728, 
    7.580461, 7.478529, 6.895574, 6.517358, 6.308734, 6.235462, 6.255989, 
    6.512051,
  2.802484, 2.649548, 3.924561, 5.832668, 6.931388, 7.824819, 8.134223, 
    8.009085, 7.596774, 6.89116, 6.46834, 6.249038, 6.21417, 5.987315, 
    6.403121,
  2.767845, 2.475387, 3.205205, 5.107605, 6.418568, 6.775819, 8.000493, 
    8.098373, 7.83745, 7.117929, 6.65395, 6.460875, 6.498897, 6.518589, 
    6.853773,
  2.692441, 2.410956, 2.747028, 3.949174, 5.79049, 6.765838, 6.787068, 
    7.690803, 7.675312, 7.365343, 7.102341, 6.917765, 6.910341, 6.91919, 
    7.167068,
  2.736143, 2.34724, 2.42227, 2.804399, 4.485392, 6.16001, 7.047057, 
    6.450584, 6.17669, 7.336764, 7.352697, 7.207138, 7.186746, 7.146554, 
    7.226553,
  2.882349, 2.527169, 2.455679, 2.375423, 2.928101, 4.569502, 6.060201, 
    6.702974, 6.887534, 7.165472, 7.151788, 7.126665, 7.116592, 7.059425, 
    6.854154,
  3.161272, 3.087829, 3.01447, 2.690786, 2.368173, 2.690667, 4.300435, 
    5.438426, 6.02347, 6.390869, 6.536343, 6.5751, 6.542778, 6.412807, 
    6.018038,
  3.498317, 3.585151, 3.719743, 3.813822, 3.117202, 2.065238, 2.310022, 
    3.717569, 4.691904, 5.264359, 5.576929, 5.708292, 5.687683, 5.508803, 
    5.04185,
  5.229099, 5.016211, 4.958512, 4.855851, 4.195187, 3.074119, 1.904404, 
    2.08639, 3.310408, 4.043128, 4.50019, 4.705191, 4.697924, 4.476276, 
    4.042296,
  6.332351, 6.27915, 6.162302, 5.881585, 5.456924, 4.328606, 2.677276, 
    1.674448, 2.156405, 3.044221, 3.517579, 3.731004, 3.716105, 3.539917, 
    3.206039,
  2.842209, 2.693594, 2.932964, 3.799031, 4.753502, 5.550584, 5.480368, 
    4.970708, 4.521391, 4.535578, 4.564947, 4.607347, 4.777975, 5.126349, 
    5.334717,
  3.875503, 3.370011, 3.459572, 4.261598, 4.959548, 5.657185, 5.450038, 
    4.858182, 4.735571, 4.785574, 4.665401, 4.769891, 5.170102, 5.276451, 
    5.516256,
  5.043345, 4.163461, 3.896659, 4.468479, 4.934148, 5.245346, 5.74575, 
    5.093059, 5.196861, 4.942849, 4.820559, 5.029574, 5.60161, 5.813528, 
    5.849651,
  5.407547, 4.64459, 4.187932, 4.446526, 4.832409, 5.523158, 5.139606, 
    5.371671, 5.26873, 5.066802, 5.083308, 5.473843, 5.851995, 5.935638, 
    6.18678,
  5.411853, 4.753894, 4.16021, 4.255702, 4.613512, 5.410459, 6.009761, 
    4.332826, 4.031295, 5.136641, 5.462096, 5.822658, 5.9783, 6.178277, 
    6.522039,
  4.868446, 4.490327, 4.04001, 3.952034, 4.264253, 5.109797, 5.869142, 
    5.168165, 4.760504, 5.22024, 5.626949, 5.900253, 6.034413, 6.376591, 
    6.527607,
  4.352332, 4.237411, 4.060153, 3.745079, 3.974472, 4.741427, 5.334013, 
    5.40908, 5.131669, 5.257598, 5.579911, 5.807872, 6.034515, 6.394638, 
    6.316137,
  4.280465, 4.229859, 4.192111, 4.008036, 3.978081, 4.342584, 4.985434, 
    5.382263, 5.215186, 5.364009, 5.526875, 5.706125, 5.978271, 6.261285, 
    5.989937,
  3.558317, 3.952133, 4.444713, 4.699707, 4.514793, 4.2692, 4.497172, 
    4.866295, 5.330228, 5.49758, 5.585335, 5.719444, 5.947673, 6.131499, 
    5.688922,
  2.296356, 2.582596, 3.535672, 4.724465, 5.157981, 4.835092, 4.396014, 
    4.198744, 5.198036, 5.553686, 5.673635, 5.830175, 6.033183, 6.063713, 
    5.544768,
  3.989848, 3.767631, 3.543747, 3.425541, 3.762631, 4.214483, 4.655097, 
    4.487042, 4.099543, 3.724952, 3.829626, 4.018326, 4.173112, 4.255723, 
    4.252446,
  3.776891, 3.785675, 3.761022, 3.660015, 4.036957, 4.294849, 4.806066, 
    4.196604, 3.696601, 3.665781, 3.62066, 3.843347, 4.016279, 3.93999, 
    4.049774,
  3.292086, 3.471569, 3.711678, 3.79788, 4.074711, 3.986922, 4.804647, 
    4.279834, 3.840243, 3.824947, 3.763091, 3.932591, 4.064262, 4.109886, 
    4.072978,
  2.734951, 2.917531, 3.469774, 3.721985, 4.004649, 4.460896, 4.200715, 
    4.550302, 4.170873, 3.961046, 4.094315, 4.128934, 4.120413, 4.064328, 
    4.043396,
  2.348217, 2.373394, 2.974496, 3.478438, 3.918372, 4.462808, 4.952353, 
    3.766846, 3.431001, 4.371184, 4.290861, 4.145262, 4.071382, 4.120478, 
    4.328499,
  2.102083, 1.933816, 2.401816, 3.056519, 3.64625, 4.276187, 5.051755, 
    4.781556, 4.417113, 4.721992, 4.432386, 4.174769, 4.248012, 4.527312, 
    4.918026,
  1.909567, 1.709554, 2.024058, 2.701716, 3.538997, 4.236028, 4.97447, 
    4.811882, 4.839747, 4.953069, 4.485791, 4.386406, 4.712715, 5.060243, 
    4.573309,
  1.751852, 1.595729, 1.872601, 2.584684, 3.789539, 4.398172, 5.010797, 
    4.803939, 5.078112, 5.036078, 4.639452, 4.806743, 5.178425, 4.672956, 
    3.106908,
  1.650129, 1.536036, 1.854415, 2.531846, 3.983759, 4.481713, 4.997337, 
    4.956159, 5.26625, 5.076952, 4.908373, 5.237398, 5.023798, 3.668142, 
    2.013397,
  1.572091, 1.409035, 1.678261, 2.489161, 4.04623, 4.556324, 5.006568, 
    5.042336, 5.266893, 5.157669, 5.231643, 5.353079, 4.401003, 2.739663, 
    1.731375,
  3.152741, 2.67493, 2.352203, 2.326431, 3.253319, 4.000698, 3.925527, 
    3.650451, 3.41356, 3.325089, 3.908326, 4.55624, 4.726718, 5.105676, 
    5.384404,
  3.236982, 2.805451, 2.485139, 2.484077, 3.365157, 4.047717, 4.019491, 
    3.652844, 3.466125, 3.305052, 3.474097, 4.036963, 4.269582, 4.249718, 
    4.534097,
  3.253012, 3.060625, 2.78334, 2.673657, 3.305277, 3.746269, 4.047632, 
    3.799907, 3.62161, 3.450997, 3.365864, 3.662967, 3.858253, 3.954947, 
    3.975285,
  3.230795, 3.201615, 3.131143, 2.918174, 3.336794, 4.026429, 3.726373, 
    3.784885, 3.500015, 3.525448, 3.525597, 3.536599, 3.607055, 3.590181, 
    3.515561,
  3.204145, 3.364191, 3.399517, 3.309447, 3.50434, 4.048776, 4.210865, 
    3.221734, 2.95514, 3.632204, 3.597862, 3.52586, 3.475894, 3.294895, 
    3.031646,
  3.113039, 3.461216, 3.70133, 3.825231, 3.871891, 4.054489, 4.206594, 
    4.058611, 3.769031, 3.695156, 3.653964, 3.477869, 3.249101, 2.925847, 
    2.487256,
  3.02576, 3.460017, 3.858174, 4.219009, 4.337049, 4.212338, 4.115528, 
    3.924215, 3.767757, 3.655356, 3.474433, 3.206799, 2.828926, 2.336837, 
    1.798757,
  2.896186, 3.383269, 3.865371, 4.343687, 4.609694, 4.347563, 4.030185, 
    3.719474, 3.512802, 3.34216, 3.049109, 2.654881, 2.15177, 1.702334, 
    1.493816,
  2.68729, 3.025867, 3.658717, 4.128526, 4.637852, 4.547298, 4.041896, 
    3.637363, 3.266467, 2.90567, 2.527024, 2.07141, 1.641024, 1.488396, 
    1.556695,
  2.564432, 2.447702, 3.158037, 3.710584, 4.412451, 4.736488, 4.258338, 
    3.584665, 3.0693, 2.588381, 2.154094, 1.675997, 1.435338, 1.498609, 
    1.622901,
  4.530949, 4.015162, 3.480858, 3.260346, 3.324287, 3.232089, 3.097164, 
    2.968708, 3.031175, 3.081416, 3.380271, 3.785471, 4.119775, 4.39464, 
    4.395212,
  4.666055, 4.221044, 3.555295, 3.162927, 3.108064, 2.980007, 2.908325, 
    2.771805, 2.749919, 2.788121, 2.952118, 3.414078, 3.927468, 4.15744, 
    4.319673,
  4.767997, 4.464066, 3.771263, 3.135352, 2.84808, 2.533081, 2.68922, 
    2.61353, 2.519, 2.433543, 2.436604, 2.61809, 3.079074, 3.632783, 3.949922,
  4.823618, 4.604214, 4.06298, 3.259818, 2.774046, 2.64416, 2.347292, 
    2.389529, 2.274925, 2.173398, 2.064066, 2.002428, 2.128346, 2.423166, 
    2.786891,
  4.980796, 4.73685, 4.332125, 3.662225, 2.827981, 2.533274, 2.426709, 
    1.888304, 1.82401, 2.032856, 1.879847, 1.696178, 1.621639, 1.608704, 
    1.652273,
  5.320511, 4.933294, 4.586428, 4.13404, 3.163338, 2.453605, 2.287863, 
    2.189328, 2.069984, 1.958663, 1.800894, 1.671277, 1.598834, 1.562139, 
    1.554238,
  5.748749, 5.077768, 4.869545, 4.568914, 3.839456, 2.685399, 2.112119, 
    1.971126, 1.912359, 1.820328, 1.759901, 1.724983, 1.694559, 1.659864, 
    1.630544,
  6.238425, 5.419972, 5.042031, 4.900532, 4.444712, 3.207993, 2.296686, 
    1.812312, 1.686306, 1.723851, 1.764485, 1.777743, 1.750013, 1.687733, 
    1.619032,
  6.798841, 5.843877, 5.337416, 4.935885, 4.664607, 3.99708, 2.776737, 
    1.992273, 1.644175, 1.634733, 1.752816, 1.803347, 1.77408, 1.67954, 
    1.588859,
  7.261636, 6.326945, 5.54692, 5.013553, 4.692529, 4.377725, 3.400143, 
    2.390939, 1.812614, 1.598161, 1.699025, 1.787225, 1.763278, 1.650284, 
    1.537937,
  7.325967, 6.855352, 6.31161, 5.688713, 5.017247, 4.286711, 3.681671, 
    3.184739, 2.757354, 2.367013, 2.21594, 2.408749, 2.754597, 3.130848, 
    3.36059,
  7.823298, 7.387142, 6.9673, 6.211422, 5.328627, 4.447277, 3.828233, 
    3.268951, 2.851064, 2.506495, 2.169285, 2.054064, 2.212057, 2.562371, 
    3.109579,
  8.242303, 7.847683, 7.455872, 6.551111, 5.429419, 4.135106, 3.667857, 
    3.189569, 2.806602, 2.484695, 2.187511, 1.913924, 1.754174, 1.920014, 
    2.438029,
  8.583893, 8.134821, 7.686901, 6.695713, 5.462612, 4.370785, 3.257237, 
    2.895887, 2.612975, 2.393206, 2.177396, 1.915389, 1.663995, 1.516888, 
    1.622039,
  8.845233, 8.258772, 7.59228, 6.451839, 5.23795, 4.180446, 3.410966, 
    2.404262, 2.041707, 2.255035, 2.164947, 1.961659, 1.694183, 1.448871, 
    1.438399,
  8.858706, 8.197088, 7.26159, 5.958924, 4.827975, 3.953078, 3.294512, 
    2.817241, 2.544633, 2.403706, 2.230205, 2.084712, 1.814345, 1.483222, 
    1.375173,
  8.659113, 7.886675, 6.693724, 5.325706, 4.306888, 3.663259, 3.265412, 
    2.918061, 2.616868, 2.396129, 2.26177, 2.186695, 1.967556, 1.609279, 
    1.386593,
  8.299469, 7.299924, 5.915369, 4.575546, 3.720959, 3.276059, 3.120589, 
    2.981866, 2.716533, 2.513861, 2.396214, 2.325147, 2.106475, 1.757356, 
    1.482819,
  7.939481, 6.534264, 5.008509, 3.705906, 3.058935, 2.82642, 2.843286, 
    2.890709, 2.777591, 2.648175, 2.590479, 2.478732, 2.214942, 1.875724, 
    1.631584,
  7.573672, 5.705915, 3.991034, 2.800445, 2.365408, 2.321173, 2.521175, 
    2.680733, 2.710653, 2.784381, 2.789739, 2.582603, 2.27515, 1.974388, 
    1.780701,
  5.990871, 5.420949, 4.770039, 4.030708, 3.37818, 2.914764, 2.701458, 
    2.541263, 2.463379, 2.46901, 2.575183, 2.649743, 2.626408, 2.622011, 
    2.670231,
  5.927097, 5.066359, 4.236558, 3.406641, 2.801244, 2.413457, 2.319085, 
    2.188177, 2.072657, 2.123238, 2.260912, 2.405395, 2.481812, 2.407641, 
    2.521737,
  5.921959, 4.76965, 3.797347, 2.937047, 2.432996, 2.027877, 2.129619, 
    2.167481, 2.080065, 2.058542, 2.0603, 2.174603, 2.356679, 2.464438, 
    2.540328,
  5.924091, 4.527116, 3.42482, 2.57592, 2.272482, 2.161448, 1.961714, 
    2.04473, 2.016983, 2.112522, 2.052494, 2.072169, 2.344825, 2.534724, 
    2.5252,
  6.022285, 4.397053, 3.180154, 2.389739, 2.235965, 2.250257, 2.210811, 
    1.781348, 1.670113, 2.111878, 2.116831, 2.160687, 2.522449, 2.655721, 
    2.454348,
  6.304735, 4.461998, 3.147582, 2.443994, 2.258277, 2.291396, 2.317623, 
    2.245443, 2.132444, 2.084442, 2.032302, 2.191521, 2.519897, 2.569552, 
    2.255248,
  6.67805, 4.683342, 3.369312, 2.716417, 2.389789, 2.301831, 2.350821, 
    2.337252, 2.219083, 2.055993, 1.972186, 2.089316, 2.297593, 2.233335, 
    1.943663,
  7.154835, 5.026504, 3.666634, 3.014992, 2.617163, 2.348064, 2.33194, 
    2.306239, 2.221155, 2.089863, 2.000596, 2.01125, 2.040158, 1.83172, 
    1.605445,
  7.562532, 5.440672, 4.056085, 3.250036, 2.878429, 2.515457, 2.340113, 
    2.325505, 2.284696, 2.22022, 2.151973, 2.065073, 1.952684, 1.666278, 
    1.433676,
  7.739046, 5.691365, 4.339107, 3.607538, 3.260447, 2.819548, 2.439703, 
    2.297567, 2.261639, 2.248911, 2.262279, 2.243552, 2.120707, 1.844254, 
    1.666508,
  6.111668, 5.679065, 5.097778, 4.530505, 4.033367, 3.539135, 3.154528, 
    2.806798, 2.536169, 2.351293, 2.279048, 2.152122, 2.079837, 2.038969, 
    2.061763,
  6.793546, 6.396019, 5.850847, 5.253456, 4.671209, 4.04314, 3.632232, 
    3.171391, 2.765962, 2.54537, 2.407386, 2.348467, 2.304309, 2.103138, 
    2.233206,
  7.489258, 7.075628, 6.604461, 5.979928, 5.315013, 4.303375, 4.092969, 
    3.665186, 3.164286, 2.794647, 2.529986, 2.439566, 2.405911, 2.432724, 
    2.553766,
  7.939807, 7.587979, 7.260186, 6.642092, 6.006068, 5.284532, 4.217343, 
    3.903455, 3.427089, 3.073653, 2.703547, 2.5025, 2.447626, 2.512365, 
    2.625912,
  8.299005, 8.050761, 7.763774, 7.203993, 6.584386, 5.918476, 5.159967, 
    3.807441, 3.346108, 3.428046, 2.9523, 2.544505, 2.394072, 2.379208, 
    2.490805,
  8.589693, 8.421563, 8.119189, 7.671114, 7.083718, 6.472326, 5.799258, 
    5.129817, 4.569621, 3.966049, 3.274777, 2.699296, 2.335592, 2.185435, 
    2.203225,
  8.743141, 8.597648, 8.295109, 7.929202, 7.480951, 6.956925, 6.387175, 
    5.814638, 5.172394, 4.464344, 3.684553, 2.985615, 2.474821, 2.180722, 
    2.042422,
  8.625211, 8.528567, 8.274516, 7.986099, 7.741352, 7.44863, 7.018749, 
    6.494545, 5.879335, 5.122853, 4.165174, 3.323427, 2.738189, 2.363776, 
    2.145818,
  8.282629, 8.231145, 8.11587, 7.941936, 7.822908, 7.74075, 7.534361, 
    7.149673, 6.527285, 5.652615, 4.546751, 3.542205, 2.898699, 2.507206, 
    2.319633,
  8.000219, 7.94959, 7.865576, 7.803851, 7.828434, 7.947626, 7.924758, 
    7.691671, 7.063043, 5.983007, 4.661269, 3.54187, 2.834967, 2.423382, 
    2.315637,
  7.60612, 7.81096, 8.207613, 8.521, 8.623829, 8.559502, 8.356553, 8.057966, 
    7.577387, 6.7956, 6.060929, 5.346844, 4.587476, 3.862378, 3.227666,
  7.367345, 7.515843, 7.923736, 8.350999, 8.477024, 8.343275, 8.41492, 
    8.19179, 7.876175, 7.390232, 6.696952, 5.916563, 5.109261, 4.222094, 
    3.651687,
  7.09854, 7.177381, 7.479711, 7.953096, 8.134372, 7.257461, 7.895354, 
    8.162504, 8.012968, 7.728634, 7.217318, 6.493237, 5.632297, 4.820558, 
    4.081011,
  6.84504, 6.817052, 6.998906, 7.395133, 7.727854, 7.726075, 6.864544, 
    7.42464, 7.618498, 7.806073, 7.524751, 6.932052, 6.10728, 5.139278, 
    4.256885,
  6.690215, 6.500786, 6.530815, 6.809023, 7.11934, 7.280737, 7.306108, 
    5.955792, 5.918492, 7.360216, 7.566185, 7.238135, 6.545895, 5.488195, 
    4.422957,
  6.606663, 6.269505, 6.090234, 6.229962, 6.415985, 6.550897, 6.716837, 
    6.859081, 7.050842, 7.415926, 7.539018, 7.373569, 6.756913, 5.6577, 
    4.415009,
  6.548616, 6.12279, 5.781674, 5.708186, 5.793103, 5.889762, 6.052062, 
    6.307394, 6.620762, 6.967875, 7.369603, 7.390039, 6.727244, 5.485428, 
    4.161627,
  6.5491, 6.084515, 5.603932, 5.280103, 5.215547, 5.267531, 5.403662, 
    5.550408, 5.812059, 6.35253, 6.916888, 6.949185, 6.047728, 4.691703, 
    3.670419,
  6.663761, 6.168548, 5.612597, 5.0356, 4.823233, 4.835423, 4.86722, 4.97327, 
    5.188738, 5.55781, 5.908551, 5.615217, 4.622052, 3.77801, 3.096632,
  6.842505, 6.291894, 5.644656, 4.993578, 4.595422, 4.467555, 4.416164, 
    4.406569, 4.492802, 4.577518, 4.514894, 4.044805, 3.463411, 2.91964, 
    2.27087,
  8.513837, 7.944526, 7.432318, 6.732757, 5.941603, 5.01576, 4.761534, 
    5.000237, 5.510416, 5.879306, 6.388119, 6.815612, 6.611206, 6.125069, 
    5.562473,
  8.998938, 8.297954, 7.663272, 6.882493, 5.910048, 4.638807, 4.279148, 
    4.262162, 4.587, 5.125633, 5.674108, 6.274784, 6.559511, 6.095191, 
    5.899978,
  9.5465, 8.703901, 8.014966, 7.210747, 6.097146, 4.429133, 3.8941, 3.928745, 
    4.131893, 4.440211, 4.96931, 5.69437, 6.274251, 6.440468, 6.172865,
  10.12925, 9.221289, 8.44635, 7.568935, 6.497611, 5.201779, 3.810127, 
    3.364443, 3.241275, 3.645022, 4.296573, 5.196465, 5.843472, 6.423974, 
    6.356822,
  10.5975, 9.738723, 8.85507, 7.919378, 6.892717, 5.729125, 4.653543, 
    3.244086, 2.733594, 3.249867, 3.905464, 4.808295, 5.622796, 6.202579, 
    6.44732,
  10.8574, 10.1314, 9.21021, 8.231205, 7.286629, 6.233813, 5.218288, 4.23245, 
    3.474863, 3.23151, 3.629226, 4.586052, 5.614941, 6.347838, 6.647988,
  10.88125, 10.27431, 9.443561, 8.50057, 7.620767, 6.693768, 5.719378, 
    4.802936, 3.927797, 3.338108, 3.291272, 4.003715, 5.178638, 6.018792, 
    5.912082,
  10.73062, 10.15806, 9.431022, 8.52554, 7.776574, 7.009819, 6.181186, 
    5.304677, 4.367595, 3.550026, 3.068122, 3.073252, 3.467907, 4.033159, 
    4.182919,
  10.43453, 9.881347, 9.141741, 8.300474, 7.76598, 7.241093, 6.596448, 
    5.822063, 4.928659, 4.017744, 3.280343, 2.868127, 2.687963, 2.633435, 
    2.519779,
  10.05585, 9.438891, 8.548856, 7.866091, 7.620677, 7.374695, 6.971637, 
    6.360987, 5.585664, 4.639149, 3.715099, 3.028218, 2.605498, 2.331719, 
    2.105798,
  9.582353, 9.249124, 9.347436, 9.769984, 9.491488, 8.582866, 7.393013, 
    6.083983, 4.861266, 3.847884, 3.384543, 3.440269, 3.877161, 4.664512, 
    5.263951,
  9.676685, 9.178324, 9.066001, 9.461491, 9.484057, 8.506057, 7.550257, 
    6.304546, 5.117249, 4.192827, 3.702318, 3.625715, 3.773305, 3.945634, 
    4.729197,
  9.657285, 9.198349, 8.8583, 8.989437, 9.183612, 7.640131, 7.622178, 
    6.711692, 5.60135, 4.621475, 3.953027, 3.750266, 3.78985, 4.024253, 
    4.546735,
  9.426965, 9.195604, 8.667191, 8.512291, 8.60268, 8.367999, 6.941072, 
    6.784792, 6.021437, 5.169592, 4.4301, 3.961621, 4.060268, 4.115557, 
    4.435039,
  9.14299, 9.086828, 8.462416, 8.091322, 7.830335, 7.684643, 7.50582, 
    5.642972, 5.150509, 5.729048, 5.181454, 4.443213, 4.308397, 4.356082, 
    4.529519,
  8.956667, 8.932019, 8.2104, 7.615618, 7.028758, 6.633527, 6.737008, 
    6.778304, 6.759799, 6.434334, 5.684899, 4.887474, 4.387047, 4.527463, 
    4.759449,
  8.83711, 8.726739, 7.973371, 7.090952, 6.21829, 5.793158, 5.940699, 
    6.319358, 6.57009, 6.536983, 6.078768, 5.386703, 4.706815, 4.57028, 
    4.899075,
  8.743425, 8.507912, 7.666651, 6.544174, 5.506983, 5.057573, 5.225665, 
    5.586634, 6.068942, 6.324464, 6.12724, 5.672739, 5.026517, 4.505733, 
    4.461388,
  8.57382, 8.248722, 7.33282, 6.066632, 5.071623, 4.50667, 4.592743, 
    4.940868, 5.376393, 5.586042, 5.51765, 5.286849, 4.923806, 4.473892, 
    4.068587,
  8.306756, 7.921785, 6.953909, 5.670521, 4.708972, 4.045765, 4.007372, 
    4.162869, 4.430986, 4.663077, 4.756469, 4.724737, 4.544703, 4.256732, 
    3.861443,
  8.019798, 7.145213, 6.598032, 6.097983, 5.994214, 6.150275, 6.563037, 
    7.000345, 7.070463, 6.341021, 5.212844, 4.369862, 3.903636, 3.74034, 
    3.810846,
  7.927999, 7.105817, 6.48687, 5.648983, 5.142137, 5.212721, 5.992762, 
    6.588723, 6.907987, 6.704432, 6.018454, 5.136569, 4.405558, 3.866603, 
    3.801108,
  7.773227, 6.968877, 6.382776, 5.426532, 4.510266, 3.989118, 4.92992, 
    5.957162, 6.36874, 6.368981, 6.182506, 5.798406, 5.136806, 4.494975, 
    4.110928,
  7.567249, 6.751995, 6.189417, 5.171385, 4.232962, 3.845719, 3.647242, 
    4.421848, 5.120361, 5.624772, 5.864594, 5.988565, 5.778203, 5.117535, 
    4.547856,
  7.309482, 6.440701, 5.871444, 4.880713, 3.898369, 3.529905, 3.509085, 
    2.947022, 3.124565, 4.422435, 5.067977, 5.578613, 5.966277, 5.754511, 
    5.198511,
  7.036446, 6.084363, 5.440097, 4.521108, 3.527798, 3.038768, 2.928547, 
    3.013509, 3.22144, 3.620855, 4.093831, 4.598403, 5.177783, 5.601701, 
    5.439557,
  6.666532, 5.679205, 4.974642, 4.069891, 3.173483, 2.646543, 2.453175, 
    2.421191, 2.563859, 2.797443, 3.05048, 3.455687, 4.025347, 4.705187, 
    5.269723,
  6.228957, 5.233988, 4.409181, 3.493507, 2.800054, 2.360166, 2.136018, 
    2.042744, 2.059196, 2.150563, 2.263716, 2.48978, 2.914998, 3.628472, 
    4.484847,
  5.691214, 4.801511, 3.928695, 2.955892, 2.444365, 2.137082, 1.952002, 
    1.854159, 1.828437, 1.868981, 1.928353, 2.047374, 2.257541, 2.716689, 
    3.461599,
  5.143183, 4.317367, 3.45525, 2.582783, 2.185315, 1.932308, 1.801414, 
    1.690472, 1.638377, 1.636443, 1.67916, 1.780024, 1.933213, 2.269741, 
    2.824316,
  3.769109, 2.939578, 2.462189, 2.215723, 2.197262, 2.135827, 2.084687, 
    2.1684, 2.591995, 3.194387, 4.011068, 4.914688, 5.029478, 4.667917, 
    4.25001,
  3.872506, 3.049498, 2.463341, 2.083217, 1.919248, 1.777549, 1.773216, 
    1.745679, 1.8997, 2.291166, 2.904683, 3.86157, 4.592413, 4.532933, 
    4.269999,
  3.847454, 3.136478, 2.607233, 2.120066, 1.86293, 1.52177, 1.545481, 
    1.564292, 1.565003, 1.620336, 1.919328, 2.639516, 3.568505, 4.298147, 
    4.509211,
  3.810828, 3.12462, 2.658334, 2.196708, 1.946514, 1.687204, 1.41824, 
    1.423338, 1.412689, 1.460363, 1.504281, 1.803439, 2.54633, 3.562495, 
    4.350646,
  3.786628, 3.131386, 2.686887, 2.284253, 2.041505, 1.798043, 1.642511, 
    1.29229, 1.22128, 1.421711, 1.408658, 1.428539, 1.769581, 2.743511, 
    3.901125,
  3.707685, 3.136702, 2.749124, 2.399574, 2.080578, 1.860101, 1.745682, 
    1.635185, 1.54055, 1.455679, 1.362104, 1.317002, 1.402129, 1.923368, 
    3.273971,
  3.575052, 3.100358, 2.768368, 2.410151, 2.092405, 1.922128, 1.825953, 
    1.735945, 1.626965, 1.486357, 1.354373, 1.256318, 1.271455, 1.516489, 
    2.56515,
  3.414002, 3.023933, 2.678634, 2.342391, 2.097594, 1.984164, 1.868955, 
    1.732145, 1.613569, 1.468285, 1.332678, 1.21614, 1.172201, 1.345723, 
    2.027724,
  3.267876, 2.94205, 2.582495, 2.245959, 2.127575, 2.005112, 1.85873, 
    1.694622, 1.573528, 1.419428, 1.297018, 1.181984, 1.109339, 1.216606, 
    1.883525,
  3.208295, 2.868111, 2.488598, 2.182267, 2.124245, 2.006307, 1.83227, 
    1.646906, 1.512541, 1.356119, 1.247633, 1.134344, 1.073512, 1.162644, 
    1.7976,
  4.536267, 4.1075, 3.805464, 3.677664, 3.719415, 3.409947, 2.762282, 
    2.062934, 1.626594, 1.491021, 1.313963, 1.530066, 3.029126, 4.227766, 
    4.813191,
  4.369241, 3.931174, 3.735861, 3.675129, 3.704293, 3.42501, 2.781728, 
    2.043318, 1.715231, 1.628276, 1.461497, 1.31245, 1.771453, 3.424371, 
    4.228174,
  3.998107, 3.654248, 3.575037, 3.543298, 3.530908, 2.929744, 2.774211, 
    2.264641, 1.896569, 1.725343, 1.649552, 1.403838, 1.316643, 2.234024, 
    3.852108,
  3.65104, 3.371601, 3.305238, 3.241618, 3.258797, 3.006374, 2.396686, 
    2.264121, 2.016956, 1.88579, 1.785051, 1.592459, 1.302472, 1.597885, 
    3.238964,
  3.323222, 3.114964, 3.047288, 3.012445, 2.913188, 2.892218, 2.584704, 
    1.917903, 1.66073, 1.930348, 1.89412, 1.726904, 1.402707, 1.368175, 
    2.498948,
  3.014462, 2.795365, 2.689163, 2.628078, 2.537979, 2.501832, 2.465235, 
    2.249787, 2.087581, 2.022979, 1.925523, 1.773542, 1.490897, 1.268733, 
    1.838897,
  2.722565, 2.459794, 2.287281, 2.198738, 2.068592, 2.014548, 2.089446, 
    2.03735, 1.954092, 1.940516, 1.914443, 1.793841, 1.552978, 1.246707, 
    1.466654,
  2.478042, 2.17813, 1.95896, 1.810403, 1.740245, 1.689956, 1.704992, 
    1.716157, 1.732989, 1.786479, 1.843251, 1.757955, 1.553614, 1.246341, 
    1.300442,
  2.354763, 2.008877, 1.745743, 1.601473, 1.557802, 1.5131, 1.522247, 
    1.55723, 1.587888, 1.646278, 1.738035, 1.690862, 1.506562, 1.222493, 
    1.229116,
  2.33116, 1.934345, 1.610672, 1.479798, 1.450746, 1.412218, 1.417094, 
    1.458552, 1.503439, 1.575206, 1.641823, 1.57774, 1.416765, 1.163081, 
    1.227992,
  3.15406, 2.905914, 2.693771, 2.541442, 2.519788, 2.826859, 3.204702, 
    3.396247, 3.109417, 2.572958, 2.093934, 1.821955, 2.490219, 3.488021, 
    4.586332,
  2.866443, 2.482595, 2.34057, 2.348196, 2.637012, 2.954729, 3.227617, 
    3.123157, 2.638121, 2.210353, 1.837693, 1.6393, 2.561898, 3.630217, 
    4.687994,
  2.421679, 2.049052, 1.994582, 2.208102, 2.663042, 2.397131, 2.822583, 
    2.648932, 2.158399, 1.826356, 1.618073, 1.512414, 2.473291, 3.903946, 
    4.971684,
  2.104327, 1.78173, 1.685473, 1.884246, 2.225315, 2.233244, 2.1319, 
    2.232756, 1.823661, 1.610183, 1.542084, 1.558325, 2.506053, 3.910938, 
    4.876163,
  1.878848, 1.601269, 1.500181, 1.529814, 1.801868, 2.002655, 2.215879, 
    1.867601, 1.447564, 1.605196, 1.619559, 1.670784, 2.510219, 3.768125, 
    4.736114,
  1.771057, 1.541195, 1.440375, 1.405123, 1.487169, 1.747647, 2.217613, 
    2.179204, 1.831471, 1.738648, 1.664211, 1.811844, 2.521975, 3.723763, 
    4.643833,
  1.722548, 1.559416, 1.515022, 1.532151, 1.62121, 1.870149, 2.30979, 
    2.282957, 1.976766, 1.774538, 1.725706, 1.923415, 2.572605, 3.611644, 
    4.485449,
  1.700495, 1.567119, 1.597502, 1.717481, 1.922209, 2.12496, 2.284757, 
    2.164126, 1.86151, 1.764301, 1.771911, 2.01001, 2.633698, 3.488863, 
    4.303257,
  1.732643, 1.523437, 1.519162, 1.702275, 1.959994, 2.084751, 2.105012, 
    1.966859, 1.785299, 1.766032, 1.807983, 2.050354, 2.605609, 3.347805, 
    4.117383,
  1.867072, 1.464745, 1.406947, 1.508201, 1.730555, 1.858871, 1.83519, 
    1.743814, 1.712906, 1.74737, 1.816828, 2.040767, 2.516214, 3.176467, 
    3.904764,
  2.411643, 2.164235, 1.981412, 1.825649, 2.082315, 2.196702, 2.045867, 
    1.741954, 2.194217, 3.286546, 3.60222, 3.37747, 3.201809, 2.939264, 
    2.709907,
  2.444198, 2.218212, 1.982644, 1.852035, 2.240699, 2.308425, 2.185968, 
    1.945933, 2.474958, 3.343773, 3.516072, 3.099657, 2.85287, 2.497269, 
    2.431468,
  2.389061, 2.187843, 2.018406, 1.851535, 2.176651, 2.185774, 2.330828, 
    2.367974, 2.846097, 3.331195, 3.224883, 2.736628, 2.545969, 2.415595, 
    2.42878,
  2.39871, 2.221126, 2.013129, 1.794183, 1.987014, 2.244708, 2.210894, 
    2.533186, 2.862989, 3.026896, 2.893695, 2.450206, 2.438728, 2.46039, 
    2.616019,
  2.417789, 2.309348, 2.045214, 1.77336, 1.797318, 1.968489, 2.225978, 
    2.073772, 2.093573, 2.577748, 2.532826, 2.297062, 2.602968, 2.764282, 
    2.972631,
  2.410807, 2.376847, 2.116833, 1.842827, 1.73066, 1.679141, 1.791264, 
    1.953914, 1.9827, 2.072559, 2.151103, 2.433065, 2.95521, 3.182327, 
    3.391471,
  2.3642, 2.328416, 2.198581, 1.925594, 1.772266, 1.655833, 1.612963, 
    1.68827, 1.768188, 1.8447, 2.247415, 2.946349, 3.489279, 3.634793, 
    3.829413,
  2.265363, 2.194674, 2.172286, 1.963321, 1.780094, 1.719429, 1.708549, 
    1.743212, 1.85408, 2.235138, 2.967615, 3.693604, 4.02868, 4.073915, 
    4.208518,
  2.160152, 1.971751, 1.924664, 1.936962, 1.837134, 1.766887, 1.874365, 
    2.093693, 2.431752, 2.99547, 3.70629, 4.212778, 4.395319, 4.420779, 
    4.52803,
  2.14248, 1.684593, 1.675236, 1.792032, 1.878468, 1.876631, 2.049428, 
    2.387505, 2.850558, 3.426763, 3.999462, 4.39463, 4.551628, 4.615529, 
    4.747889,
  3.499617, 2.722585, 2.051421, 1.932951, 2.558417, 2.922597, 3.167916, 
    3.31092, 3.369139, 3.223552, 3.387476, 3.89917, 4.080697, 3.89532, 
    3.591871,
  3.502519, 2.678802, 2.099275, 2.055174, 2.653282, 2.974746, 3.269577, 
    3.539887, 3.725445, 4.020655, 4.456006, 4.741135, 4.542035, 3.956384, 
    3.783752,
  3.226085, 2.665977, 2.196113, 2.090098, 2.57708, 2.74953, 3.122208, 
    3.398784, 3.604973, 3.829982, 4.107096, 4.300121, 4.283542, 4.107526, 
    3.982704,
  2.970419, 2.521852, 2.16479, 2.024146, 2.400759, 2.718449, 2.69633, 
    2.979332, 3.058571, 3.19086, 3.296524, 3.45876, 3.641802, 3.734059, 
    3.789937,
  2.713591, 2.455775, 2.120607, 1.945318, 2.195893, 2.48549, 2.555209, 
    2.091541, 2.134897, 2.593947, 2.633286, 2.598114, 2.76011, 3.015881, 
    3.310606,
  2.612645, 2.464987, 2.1329, 1.904138, 1.992888, 2.266583, 2.475016, 
    2.404246, 2.245494, 2.194064, 2.155559, 2.129079, 2.175689, 2.374182, 
    2.776566,
  2.59017, 2.542966, 2.330591, 2.054457, 1.920103, 1.974091, 2.123394, 
    2.220895, 2.14609, 1.983198, 1.943783, 1.947041, 1.946559, 2.027643, 
    2.392745,
  2.468713, 2.553684, 2.494981, 2.357512, 2.295097, 2.302902, 2.32888, 
    2.229841, 2.054839, 1.926285, 1.996235, 2.037472, 2.01649, 2.031497, 
    2.387814,
  2.278137, 2.359988, 2.387501, 2.477473, 2.676967, 2.90721, 3.11808, 
    3.226806, 3.156934, 2.853803, 2.588821, 2.423685, 2.266024, 2.222948, 
    2.636337,
  2.153186, 1.934063, 2.182054, 2.372834, 2.612033, 2.952683, 3.471967, 
    3.773368, 3.82539, 3.367615, 3.064547, 2.87625, 2.736865, 2.722194, 
    3.250064,
  2.983653, 3.087065, 3.070965, 2.850899, 2.648502, 2.410697, 2.344407, 
    2.480111, 2.909543, 3.256648, 3.324338, 2.547094, 1.788833, 1.925781, 
    2.096894,
  3.221552, 3.169874, 3.065052, 2.78472, 2.609705, 2.314236, 2.289453, 
    2.26175, 2.51339, 3.01686, 3.446888, 3.33045, 1.975819, 1.647293, 1.895318,
  3.323973, 3.232251, 3.061242, 2.718894, 2.553512, 2.210336, 2.267544, 
    2.277803, 2.275843, 2.533075, 3.159735, 3.707462, 3.069208, 2.039406, 
    1.903848,
  3.503249, 3.316522, 3.039274, 2.704776, 2.600042, 2.460929, 2.200347, 
    2.179606, 2.191279, 2.272087, 2.490753, 3.601891, 3.852657, 2.867699, 
    2.261142,
  3.686526, 3.447513, 3.137437, 2.804288, 2.670139, 2.576196, 2.545848, 
    2.019721, 1.941531, 2.309743, 2.121419, 2.984063, 3.947845, 3.722543, 
    3.049148,
  3.751791, 3.62179, 3.424654, 3.054268, 2.806206, 2.703575, 2.733234, 
    2.705329, 2.701415, 2.494325, 2.085754, 2.513022, 3.721604, 4.253849, 
    3.982718,
  3.905722, 3.929025, 3.806765, 3.415146, 3.061207, 2.87246, 2.963444, 
    3.009074, 3.030289, 2.70048, 2.190412, 2.326635, 3.343984, 4.315184, 
    4.615224,
  4.437584, 4.507526, 4.247693, 3.706094, 3.267431, 2.996235, 3.136557, 
    3.201927, 3.12257, 2.884858, 2.296323, 2.297559, 3.137633, 4.222907, 
    4.83084,
  5.623108, 5.348842, 4.73459, 3.947483, 3.337218, 2.944453, 3.153364, 
    3.350461, 3.195108, 3.039224, 2.435931, 2.304379, 3.070525, 4.159372, 
    4.878017,
  6.610403, 5.935197, 5.066625, 4.034491, 3.38537, 2.833153, 3.148825, 
    3.523294, 3.380194, 3.279673, 2.643945, 2.443153, 3.132267, 3.993731, 
    4.605543,
  4.557564, 4.791428, 4.95899, 4.681499, 4.296062, 4.218097, 4.255728, 
    3.838643, 3.166243, 3.139289, 2.899043, 2.403603, 1.969989, 2.314613, 
    2.640026,
  5.568845, 5.645477, 5.489126, 4.978655, 4.729512, 4.66319, 4.645331, 
    3.912897, 2.975162, 3.197607, 3.087128, 2.606234, 2.030283, 2.030647, 
    2.415592,
  6.368697, 6.213539, 5.751673, 5.361815, 5.296244, 4.834259, 4.747727, 
    3.793142, 2.81881, 3.232063, 3.320928, 2.956716, 2.315037, 2.017087, 
    2.141748,
  6.891578, 6.498988, 6.056515, 5.91925, 5.946109, 5.536232, 4.182575, 
    3.202742, 2.486424, 3.20617, 3.531276, 3.460044, 2.851543, 2.244046, 
    1.942619,
  7.38123, 6.727386, 6.429513, 6.460271, 6.156067, 5.341203, 3.905515, 
    2.498777, 1.964527, 3.066499, 3.62728, 3.910299, 3.63008, 3.014755, 
    2.436659,
  7.678977, 6.878423, 6.762096, 6.617901, 5.80089, 4.458975, 3.357278, 
    2.967176, 2.463767, 3.066922, 3.645983, 4.127822, 4.34306, 4.003935, 
    3.574688,
  7.851191, 7.049575, 6.939361, 6.378782, 5.112241, 3.477194, 3.241225, 
    3.105904, 2.516663, 3.029304, 3.515603, 4.194358, 4.624767, 4.691849, 
    4.525694,
  7.962706, 7.008347, 6.697079, 5.743005, 4.254813, 2.995071, 3.292023, 
    3.264719, 2.637813, 2.982671, 3.3281, 4.169497, 4.691402, 4.918298, 
    4.998994,
  7.870068, 6.634446, 6.146092, 5.093441, 3.832717, 2.832086, 3.315401, 
    3.423364, 2.854652, 2.828449, 3.137145, 4.073994, 4.759041, 5.028742, 
    5.151587,
  7.755088, 6.21642, 5.608957, 4.915828, 3.874058, 2.768068, 3.28879, 
    3.491171, 2.928774, 2.679589, 3.011765, 3.945305, 4.617472, 4.970911, 
    5.200715,
  7.209538, 7.254179, 7.02319, 6.64797, 6.27569, 6.010928, 5.866068, 
    5.466526, 4.834076, 3.512074, 3.338849, 3.672656, 3.67696, 3.221041, 
    3.067741,
  7.973291, 7.223732, 6.453267, 5.897141, 5.356953, 5.011526, 5.052474, 
    4.636077, 3.975995, 3.165289, 3.316692, 3.686141, 3.807479, 3.380313, 
    3.194874,
  8.087541, 6.674561, 5.825536, 5.228349, 4.526318, 3.578635, 4.009686, 
    3.941784, 3.357499, 2.958343, 3.150669, 3.551273, 3.816599, 3.903892, 
    3.664088,
  7.958426, 6.097031, 5.396305, 4.646915, 3.897831, 3.16182, 2.954016, 
    3.267595, 2.904658, 2.792337, 2.980856, 3.40336, 3.838939, 4.183229, 
    4.234686,
  7.835892, 5.82304, 5.149856, 4.383593, 3.586442, 2.788858, 3.042184, 
    2.636258, 2.283144, 2.643818, 2.869894, 3.383733, 3.901964, 4.366015, 
    4.621754,
  7.92003, 6.026717, 5.272566, 4.57075, 3.704987, 2.798908, 3.0323, 3.094627, 
    2.700342, 2.645845, 2.868876, 3.549366, 4.108202, 4.639934, 4.76426,
  8.056192, 6.562974, 5.84664, 5.009724, 3.987897, 2.89057, 3.026597, 
    3.161156, 2.850897, 2.79368, 3.088765, 3.849743, 4.497312, 4.826194, 
    4.75402,
  8.239469, 6.929266, 6.331998, 5.49061, 4.387389, 2.974763, 3.011258, 
    3.224801, 3.056551, 3.132137, 3.609109, 4.268995, 4.748509, 4.725841, 
    4.431614,
  8.369341, 7.351572, 6.589904, 5.914669, 4.678504, 3.004132, 2.987907, 
    3.366812, 3.36131, 3.547513, 4.081276, 4.559145, 4.628126, 4.253536, 
    3.857911,
  8.403455, 7.496348, 6.504117, 6.082783, 4.744597, 2.889343, 2.956067, 
    3.551405, 3.732574, 4.057195, 4.501506, 4.586694, 4.304857, 3.817433, 
    3.421602,
  6.293682, 5.428345, 5.32763, 5.072456, 4.548679, 3.472104, 3.089758, 
    3.088285, 3.198637, 3.220043, 3.195978, 3.171095, 3.104976, 3.076177, 
    3.136707,
  6.85218, 6.211093, 6.104483, 5.687582, 4.978448, 3.637371, 3.199186, 
    3.067528, 3.021036, 3.08744, 3.124286, 3.062515, 2.938617, 2.696341, 
    2.805709,
  7.280802, 7.041902, 6.856785, 6.173888, 5.282218, 3.473056, 3.174244, 
    3.187564, 3.136798, 3.228454, 3.271253, 3.222955, 3.116578, 3.179366, 
    3.36767,
  7.712852, 7.771276, 7.192163, 6.419303, 5.527432, 3.956396, 2.89543, 
    3.122161, 3.132908, 3.463544, 3.450401, 3.396644, 3.463445, 3.693292, 
    3.944455,
  8.2792, 8.244146, 7.212874, 6.568806, 5.591188, 4.087189, 3.297952, 
    2.769493, 2.759277, 3.585373, 3.549633, 3.487183, 3.483338, 3.524214, 
    3.532099,
  8.584555, 8.322996, 7.009855, 6.553939, 5.311927, 3.86762, 3.40652, 
    3.612133, 3.705238, 3.730592, 3.566783, 3.415786, 3.301656, 3.202378, 
    3.080674,
  8.620288, 8.070131, 6.562823, 6.290575, 4.866275, 3.550688, 3.558096, 
    3.765872, 3.831231, 3.70156, 3.484458, 3.292678, 3.14881, 3.169714, 
    3.154573,
  8.696455, 7.7811, 6.078976, 5.780819, 4.382883, 3.355908, 3.678395, 
    3.812224, 3.706637, 3.515254, 3.249784, 3.065049, 3.058991, 3.237072, 
    3.51458,
  8.695939, 7.630133, 5.788574, 5.229248, 3.781351, 3.254816, 3.826428, 
    3.857267, 3.611631, 3.297841, 2.97787, 2.902338, 3.113047, 3.412519, 
    3.7015,
  8.842023, 7.621782, 5.641138, 4.814659, 3.437655, 3.230013, 3.93778, 
    3.851342, 3.47382, 3.037254, 2.738965, 2.842078, 3.184585, 3.532647, 
    3.715823,
  6.654067, 7.416696, 7.671727, 6.750713, 5.27905, 4.379641, 3.8397, 
    3.428758, 3.333867, 3.456208, 3.548582, 3.575531, 3.480793, 3.29105, 
    3.175265,
  6.969968, 7.616425, 7.155265, 5.883026, 4.519498, 3.753013, 3.447439, 
    3.193373, 3.23579, 3.489512, 3.584736, 3.565717, 3.516615, 3.239524, 
    3.153322,
  7.447556, 7.614348, 6.572721, 5.159626, 3.801921, 2.919963, 3.071366, 
    3.158817, 3.214425, 3.421263, 3.445616, 3.443725, 3.398508, 3.334971, 
    3.306785,
  7.898911, 7.473766, 6.110063, 4.674467, 3.487794, 3.005955, 2.712054, 
    2.836778, 2.839649, 3.210677, 3.340852, 3.421202, 3.423479, 3.308456, 
    3.159357,
  8.276887, 7.326263, 5.828386, 4.349104, 3.286091, 3.054174, 2.944444, 
    2.361815, 2.337984, 3.045074, 3.343888, 3.534223, 3.647156, 3.560654, 
    3.324588,
  8.445845, 7.262885, 5.443128, 4.07661, 3.200236, 2.998349, 2.889374, 
    2.770776, 2.767639, 3.040771, 3.328365, 3.571512, 3.749479, 3.690703, 
    3.558584,
  8.592295, 7.205807, 5.018118, 3.889879, 3.243426, 3.010605, 2.692489, 
    2.67503, 2.735747, 2.898777, 3.194007, 3.466459, 3.656273, 3.632537, 
    3.452358,
  8.683373, 7.174921, 4.72156, 3.69364, 3.287718, 3.047639, 2.625286, 
    2.611311, 2.602797, 2.644559, 2.952937, 3.318614, 3.582505, 3.558244, 
    3.269605,
  8.818949, 7.35876, 4.690948, 3.65196, 3.317644, 3.118548, 2.669379, 
    2.645614, 2.549183, 2.460636, 2.656395, 3.144411, 3.534575, 3.634521, 
    3.220217,
  9.134672, 7.727361, 5.225503, 4.003109, 3.496824, 3.273197, 2.812458, 
    2.668115, 2.526073, 2.335699, 2.402152, 2.903871, 3.501468, 3.782116, 
    3.455901,
  6.267277, 5.38967, 4.122583, 3.075052, 2.643148, 2.61491, 2.5234, 2.541498, 
    2.60708, 2.713355, 2.827997, 2.896755, 2.944935, 3.028527, 3.163675,
  6.878769, 5.910535, 4.421914, 3.334965, 2.782611, 2.585108, 2.513308, 
    2.48876, 2.512913, 2.65404, 2.789406, 2.831569, 2.848107, 2.858712, 
    3.104759,
  7.76629, 6.776951, 5.279746, 3.888868, 3.150906, 2.468816, 2.543403, 
    2.600649, 2.599161, 2.742325, 2.816427, 2.823302, 2.808643, 2.96357, 
    3.216549,
  8.447409, 7.630986, 6.232863, 4.820366, 3.949048, 3.278011, 2.666593, 
    2.647185, 2.659385, 2.935404, 2.977797, 2.874072, 2.834172, 2.992055, 
    3.276508,
  8.92794, 8.353858, 7.047129, 5.786854, 4.82423, 4.068209, 3.517159, 
    2.625541, 2.576953, 3.220239, 3.264222, 3.022444, 2.883407, 3.036249, 
    3.364985,
  9.256662, 8.847778, 7.614021, 6.517859, 5.497707, 4.72356, 4.147725, 
    3.888714, 3.889632, 3.884087, 3.605391, 3.215132, 2.979491, 3.141366, 
    3.440402,
  9.69609, 9.261462, 8.020361, 6.974189, 6.03206, 5.328271, 4.950701, 
    4.819713, 4.662007, 4.402325, 3.956778, 3.410848, 3.116222, 3.255923, 
    3.470357,
  9.741774, 9.055382, 8.06637, 7.170731, 6.434175, 6.001569, 5.775923, 
    5.6134, 5.317965, 4.884771, 4.243186, 3.539583, 3.209622, 3.327228, 
    3.469884,
  9.318039, 8.680649, 8.172744, 7.586935, 7.074222, 6.760844, 6.537755, 
    6.25378, 5.749541, 5.137803, 4.381271, 3.581087, 3.265701, 3.362716, 
    3.453315,
  8.783124, 8.350867, 8.299927, 8.174428, 7.843135, 7.504353, 7.085124, 
    6.548901, 5.830253, 5.143632, 4.335726, 3.511354, 3.268041, 3.374387, 
    3.475027,
  8.85058, 9.226281, 9.221837, 8.657557, 7.775813, 6.822361, 5.786491, 
    4.866254, 4.490345, 4.321977, 4.332764, 4.34304, 4.067374, 3.675359, 
    3.113275,
  9.396871, 9.632346, 9.679029, 9.107429, 8.159036, 7.157727, 6.262831, 
    5.453461, 5.122083, 5.104277, 5.130974, 5.12098, 4.846115, 4.25899, 
    3.962982,
  9.550809, 9.889986, 9.866782, 9.281326, 8.268544, 6.842995, 6.653253, 
    6.344786, 6.172187, 6.112078, 6.029701, 5.968645, 5.745527, 5.339065, 
    4.851357,
  9.730026, 9.984319, 9.852345, 9.176452, 8.294284, 7.527454, 6.289605, 
    6.603657, 6.704593, 6.904984, 6.885777, 6.746643, 6.600075, 6.241902, 
    5.611917,
  9.922293, 10.00671, 9.68747, 9.016795, 8.284453, 7.737276, 7.467423, 
    6.067121, 6.004193, 7.419163, 7.570933, 7.349676, 7.115969, 6.772894, 
    6.218899,
  10.27588, 10.19715, 9.620399, 8.793287, 7.982997, 7.728567, 7.962442, 
    8.080276, 8.055662, 7.946735, 7.605737, 7.227837, 6.946789, 6.724551, 
    6.409473,
  10.71333, 10.36035, 9.491461, 8.418624, 7.900054, 8.102244, 8.384191, 
    8.335675, 7.827921, 7.081195, 6.59944, 6.387161, 6.285495, 6.160093, 
    6.00105,
  10.99513, 10.34578, 9.185271, 8.322007, 8.373759, 8.557677, 8.170141, 
    7.10098, 6.076751, 5.702322, 5.566389, 5.419391, 5.292042, 5.175341, 
    5.073308,
  11.09916, 10.04041, 8.85006, 8.489003, 8.495212, 7.836075, 6.461823, 
    5.269623, 4.909168, 4.68871, 4.370581, 4.217099, 4.20229, 4.146053, 
    4.107328,
  10.7998, 9.29021, 8.54826, 8.219111, 7.472632, 5.860778, 4.602911, 
    4.239028, 3.945697, 3.577632, 3.432049, 3.489847, 3.653716, 3.692054, 
    3.672468,
  10.76664, 10.52019, 10.55394, 10.61697, 10.25702, 9.313604, 8.470913, 
    7.715759, 6.927315, 6.216393, 5.976269, 6.096914, 6.268078, 6.177689, 
    6.041402,
  11.03305, 10.74892, 10.56515, 10.2733, 9.5359, 8.529042, 8.022726, 
    7.249798, 6.666927, 6.443257, 6.498727, 6.642282, 6.779911, 6.418138, 
    6.343586,
  10.778, 10.3616, 10.00322, 9.419996, 8.624924, 7.118848, 7.110012, 
    6.801836, 6.4748, 6.406756, 6.732176, 7.166802, 7.398701, 7.470784, 
    7.23982,
  10.42928, 9.83266, 9.109961, 8.356993, 7.934232, 7.07467, 5.566063, 
    5.692984, 5.797881, 6.101326, 6.387788, 6.713271, 6.992796, 7.138652, 
    7.196589,
  9.907288, 9.042927, 8.087173, 7.410185, 6.903185, 6.177038, 5.598679, 
    4.31191, 4.254658, 5.183249, 5.148353, 5.053649, 4.914062, 4.822609, 
    5.148086,
  9.179021, 8.075456, 7.12179, 6.426383, 5.743294, 5.037995, 4.651291, 
    4.539508, 4.451907, 4.06652, 3.744229, 3.495705, 3.326992, 3.21685, 
    3.232673,
  8.384148, 7.147874, 6.19138, 5.355512, 4.660345, 3.912553, 3.662837, 
    3.529296, 3.334952, 3.137414, 3.064641, 3.052295, 3.060934, 3.049845, 
    3.006008,
  7.680834, 6.270087, 5.146869, 4.382438, 3.64653, 3.038038, 2.996172, 
    3.010675, 3.03793, 3.008433, 3.050913, 3.095134, 3.127287, 3.114507, 
    3.056467,
  6.810222, 5.324772, 4.328925, 3.70101, 3.107615, 2.758437, 2.946965, 
    3.061856, 3.078398, 3.039018, 3.095463, 3.180629, 3.198543, 3.163159, 
    3.138822,
  5.970464, 4.596522, 3.873557, 3.480948, 3.02126, 2.781555, 3.043936, 
    3.126798, 3.088036, 3.066294, 3.107001, 3.181471, 3.187995, 3.146198, 
    3.120985,
  5.463943, 5.029842, 4.813928, 4.526978, 4.11249, 3.624468, 3.333274, 
    3.152622, 3.151715, 3.319501, 3.765445, 4.399313, 5.046099, 5.430715, 
    5.929385,
  5.172504, 4.490908, 4.121485, 3.930184, 3.554338, 3.070813, 2.907197, 
    2.76504, 2.768969, 2.902863, 3.211713, 3.732486, 4.523732, 4.926115, 
    5.525696,
  5.115424, 4.432615, 4.0086, 3.720655, 3.221225, 2.539096, 2.663334, 
    2.716339, 2.716554, 2.79564, 2.868831, 3.072874, 3.577985, 4.342608, 
    5.355569,
  5.298311, 4.604178, 4.221787, 3.850687, 3.32851, 2.760931, 2.442729, 
    2.549297, 2.565604, 2.77583, 2.8419, 2.861239, 3.016, 3.395089, 4.373087,
  5.743183, 4.995321, 4.572604, 4.116173, 3.477882, 2.899261, 2.798012, 
    2.204927, 2.139892, 2.768271, 2.839128, 2.804303, 2.899174, 3.000872, 
    3.290478,
  6.245255, 5.606478, 5.01426, 4.453892, 3.674314, 3.009749, 2.910751, 
    2.731631, 2.740515, 2.856979, 2.837739, 2.769518, 2.849031, 2.950528, 
    3.02642,
  6.872692, 6.289749, 5.517069, 4.780639, 3.889224, 3.175567, 3.004574, 
    2.82172, 2.847146, 2.896012, 2.828379, 2.757865, 2.819245, 2.891248, 
    3.01384,
  7.680988, 7.033404, 6.003826, 5.09022, 4.170074, 3.379894, 3.126625, 
    2.860132, 2.848122, 2.92895, 2.883335, 2.771353, 2.84232, 2.890123, 
    2.894142,
  8.486995, 7.688282, 6.458491, 5.571928, 4.556363, 3.662788, 3.307631, 
    2.994596, 2.932901, 2.966855, 2.939917, 2.820636, 2.835219, 2.904518, 
    2.933754,
  9.194354, 8.175853, 6.968814, 6.137554, 5.057213, 4.040121, 3.493856, 
    3.114326, 3.029386, 3.025489, 2.98042, 2.857137, 2.831261, 2.91769, 
    3.005715,
  7.045609, 6.569025, 6.170732, 5.905391, 5.794209, 5.569685, 5.122843, 
    4.41304, 3.747571, 3.17279, 2.84027, 2.679986, 2.704805, 3.178903, 
    4.075509,
  8.179524, 7.774349, 7.332254, 6.918001, 6.682171, 6.213165, 5.771207, 
    4.955486, 4.122656, 3.48633, 2.990872, 2.751672, 2.678679, 2.685604, 
    3.306127,
  9.159645, 8.734533, 8.311255, 7.921947, 7.547009, 6.366226, 6.224566, 
    5.496604, 4.536515, 3.744521, 3.132354, 2.845334, 2.752671, 2.688766, 
    2.988478,
  10.2074, 9.669072, 9.215437, 8.815309, 8.366987, 7.632214, 6.212741, 
    5.669998, 4.682748, 3.884167, 3.253049, 2.917571, 2.827582, 2.778262, 
    2.83354,
  11.09914, 10.40641, 9.916208, 9.478476, 9.007859, 8.304241, 7.243289, 
    5.139644, 4.151531, 4.022151, 3.411862, 3.007001, 2.894509, 2.825892, 
    2.814635,
  11.41244, 10.64705, 10.20854, 9.842825, 9.392253, 8.782264, 7.605326, 
    6.295743, 5.090904, 4.05763, 3.399667, 3.089553, 2.947623, 2.917498, 
    2.867538,
  11.06246, 10.47144, 10.2905, 10.02499, 9.700668, 8.976203, 7.570206, 
    6.2224, 4.736881, 3.812334, 3.370627, 3.181767, 3.032396, 2.966881, 
    2.886277,
  10.32509, 10.33652, 10.23693, 10.13812, 9.822941, 8.64498, 7.062391, 
    5.802555, 4.50318, 3.72433, 3.399537, 3.278613, 3.138141, 2.979936, 
    2.901738,
  10.16449, 10.33029, 10.18655, 10.16898, 9.484523, 7.712993, 6.506192, 
    5.409941, 4.27702, 3.643284, 3.385866, 3.296844, 3.17369, 2.994457, 
    2.847829,
  10.23451, 10.26163, 10.19668, 9.796324, 8.32756, 6.643465, 5.883527, 
    4.859286, 4.022707, 3.441894, 3.251856, 3.22424, 3.131345, 2.967885, 
    2.8142,
  14.18543, 13.5569, 12.73491, 11.87405, 11.07983, 10.38189, 9.768774, 
    9.344796, 8.856325, 8.112348, 7.234334, 6.248704, 5.123682, 3.895703, 
    2.880206,
  14.03906, 13.17919, 12.36962, 11.61609, 10.92364, 10.09231, 9.34963, 
    8.71602, 8.347219, 7.743145, 6.966982, 6.090709, 5.064558, 3.744072, 
    2.797523,
  13.57949, 12.51559, 11.78996, 10.94327, 9.981718, 8.240983, 8.062984, 
    7.546301, 6.875381, 6.079256, 5.635139, 5.28419, 4.625492, 3.699389, 
    2.850917,
  12.73877, 11.77883, 10.90338, 9.650856, 8.525114, 7.83366, 6.220677, 
    5.799187, 5.084248, 4.909005, 4.904626, 4.693609, 4.008946, 3.426654, 
    2.814178,
  11.92585, 10.85893, 9.672392, 8.25574, 7.308388, 6.600255, 5.656422, 
    3.768526, 3.336413, 4.234587, 4.329541, 3.992834, 3.522971, 3.203915, 
    2.845244,
  11.04632, 9.836801, 8.467513, 7.156545, 6.184958, 5.406956, 4.422915, 
    3.811089, 3.530524, 3.681994, 3.794293, 3.507472, 3.252291, 3.095807, 
    2.939279,
  10.21677, 8.996398, 7.628671, 6.245496, 5.247989, 4.321784, 3.610562, 
    3.397528, 3.314247, 3.33857, 3.364679, 3.245533, 3.142921, 3.083522, 
    3.027138,
  9.539071, 8.381443, 6.872789, 5.402499, 4.314101, 3.576802, 3.297981, 
    3.176, 3.186312, 3.221328, 3.237206, 3.197407, 3.193785, 3.17114, 3.085145,
  8.837901, 7.734121, 6.029738, 4.502728, 3.534803, 3.234166, 3.158798, 
    3.176, 3.227818, 3.243941, 3.239756, 3.228018, 3.190483, 3.185936, 
    3.039505,
  7.921786, 6.683078, 5.079771, 3.723272, 3.19792, 3.041039, 3.022671, 
    3.123523, 3.19601, 3.222903, 3.222173, 3.165977, 3.096612, 3.060966, 
    2.977906,
  5.892379, 5.009682, 4.392601, 4.211637, 3.983777, 3.599501, 3.399666, 
    3.42232, 3.680033, 4.133722, 4.851659, 5.731632, 6.103586, 6.392211, 
    6.380581,
  5.829034, 4.748981, 3.844049, 3.523578, 3.479873, 3.038227, 2.869786, 
    2.806178, 2.928677, 3.276571, 3.889992, 5.502242, 6.142882, 6.087595, 
    6.153087,
  5.748185, 4.598561, 3.558036, 3.088164, 2.963502, 2.579417, 2.671686, 
    2.730986, 2.794021, 3.060625, 3.445437, 4.210445, 5.920677, 6.032088, 
    5.857402,
  5.59837, 4.456343, 3.462892, 2.945196, 2.883201, 2.77233, 2.501907, 
    2.626981, 2.643039, 3.059616, 3.567781, 4.480979, 5.259212, 5.391499, 
    5.24451,
  5.415699, 4.313585, 3.45939, 2.97773, 2.932792, 2.934221, 2.870577, 
    2.326331, 2.289191, 2.987948, 3.320851, 3.832345, 4.421042, 4.678993, 
    4.773734,
  5.246943, 4.205981, 3.425029, 3.068, 3.000215, 3.018672, 3.033963, 
    2.989794, 2.928755, 3.007342, 3.147685, 3.423115, 3.779218, 3.994614, 
    3.99504,
  4.957024, 4.072452, 3.359761, 3.067152, 3.057974, 3.093873, 3.105323, 
    3.10513, 3.071731, 3.062741, 3.041126, 3.050044, 3.170765, 3.288404, 
    3.238453,
  4.512768, 3.851314, 3.215624, 3.069969, 3.098194, 3.138977, 3.177653, 
    3.162795, 3.112839, 3.111746, 3.090914, 3.055667, 2.978062, 2.912637, 
    2.838336,
  4.161303, 3.607565, 3.152175, 3.111004, 3.141785, 3.188162, 3.22245, 
    3.232113, 3.184228, 3.143195, 3.127604, 3.089555, 3.088202, 3.030011, 
    2.882259,
  3.703666, 3.383552, 3.206918, 3.169111, 3.17628, 3.211337, 3.248387, 
    3.249673, 3.201288, 3.16734, 3.192826, 3.161044, 3.027592, 3.018349, 
    3.013378,
  3.985511, 4.227221, 4.230577, 4.020228, 3.773885, 3.405806, 3.099493, 
    2.915393, 2.833059, 2.973823, 3.111104, 3.359109, 3.418058, 3.536018, 
    4.019014,
  4.337959, 4.541856, 4.371753, 4.043313, 3.765853, 3.331985, 3.090594, 
    2.916447, 2.817488, 3.10697, 3.319368, 3.626865, 3.701414, 3.451321, 
    3.662135,
  4.595344, 4.681103, 4.417688, 3.980273, 3.642334, 2.999025, 3.005172, 
    2.969352, 2.862635, 3.146253, 3.380323, 3.861221, 4.331372, 4.20361, 
    4.056159,
  4.785011, 4.762186, 4.359654, 3.869963, 3.549342, 3.235064, 2.77019, 
    2.854778, 2.722833, 3.070046, 3.282116, 3.852713, 4.582411, 4.68797, 
    4.48752,
  4.937435, 4.797616, 4.303345, 3.740504, 3.431587, 3.193539, 3.052465, 
    2.451422, 2.324183, 2.983249, 3.163333, 3.531717, 4.307925, 4.73169, 
    4.768223,
  5.019601, 4.829304, 4.244674, 3.642472, 3.316709, 3.146338, 3.069159, 
    3.034457, 2.917322, 2.963959, 3.1294, 3.30579, 3.657881, 4.207175, 
    4.529918,
  5.051663, 4.842809, 4.224565, 3.581525, 3.238136, 3.095406, 3.076197, 
    3.075033, 3.001448, 2.989743, 3.067723, 3.241222, 3.48811, 3.743306, 
    4.024806,
  5.072817, 4.819535, 4.217023, 3.564268, 3.167601, 3.020747, 3.026413, 
    3.035835, 2.954719, 2.925712, 2.969047, 3.055119, 3.247798, 3.457934, 
    3.580349,
  5.081898, 4.786375, 4.258551, 3.615716, 3.156576, 2.96368, 2.975163, 
    3.000161, 2.957304, 2.91418, 2.905661, 2.987212, 3.11499, 3.355955, 
    3.656809,
  5.086109, 4.719002, 4.316095, 3.715358, 3.170925, 2.917274, 2.903375, 
    2.928158, 2.918882, 2.911131, 2.913474, 2.925345, 3.018318, 3.33543, 
    3.791674,
  6.644754, 5.423779, 3.550655, 2.783544, 2.92422, 3.041261, 3.021804, 
    2.998224, 2.953147, 2.901919, 2.791601, 3.080317, 4.158951, 6.143224, 
    7.909285,
  6.905027, 5.099455, 3.354306, 2.654331, 2.756675, 2.872023, 2.979901, 
    2.968838, 2.980468, 3.108582, 3.027285, 3.01464, 3.611794, 4.809115, 
    6.517363,
  6.915849, 4.798855, 3.296916, 2.611594, 2.632788, 2.586519, 2.87696, 
    3.049021, 3.110345, 3.30222, 3.280678, 3.187842, 3.416404, 4.254824, 
    5.488406,
  6.581875, 4.49825, 3.26118, 2.584388, 2.619659, 2.797373, 2.655943, 
    2.896965, 3.061983, 3.385011, 3.493916, 3.427888, 3.41546, 4.017297, 
    4.700324,
  5.939834, 4.26915, 3.221918, 2.608145, 2.566927, 2.82085, 2.899627, 
    2.529669, 2.65819, 3.442392, 3.703838, 3.743537, 3.515305, 3.611672, 
    4.280304,
  5.443855, 4.252469, 3.19783, 2.649152, 2.490418, 2.676136, 2.924595, 
    3.000393, 3.172886, 3.547699, 3.94022, 4.151004, 3.929991, 3.423805, 
    3.712392,
  5.329051, 4.291383, 3.255826, 2.627599, 2.473739, 2.592916, 2.803555, 
    3.017307, 3.233854, 3.64925, 4.142776, 4.573569, 4.728231, 4.037848, 
    3.357547,
  5.348481, 4.28704, 3.283462, 2.659445, 2.463777, 2.541398, 2.676178, 
    2.884328, 3.133376, 3.607434, 4.276472, 4.926177, 5.358703, 5.077865, 
    4.031385,
  5.324184, 4.309698, 3.395927, 2.779561, 2.54064, 2.532774, 2.605325, 
    2.766968, 3.050172, 3.539179, 4.313266, 5.158752, 5.937226, 6.25639, 
    5.479428,
  5.248086, 4.310118, 3.697031, 2.96205, 2.613735, 2.565857, 2.573399, 
    2.653434, 2.915497, 3.407134, 4.167152, 5.181341, 6.15246, 6.888286, 
    7.046852,
  8.82457, 7.83271, 5.375149, 2.750547, 2.3787, 2.75746, 3.427728, 4.019059, 
    4.08758, 3.707071, 3.470421, 3.966929, 5.438085, 7.38829, 8.522181,
  8.719102, 6.875017, 3.420242, 2.356157, 2.32156, 2.908264, 3.700983, 
    4.221347, 4.296171, 4.128306, 3.647555, 3.724689, 4.658536, 6.293486, 
    8.07297,
  6.768447, 4.182883, 2.749778, 2.31911, 2.349488, 2.871315, 3.812479, 
    4.427012, 4.595894, 4.625468, 4.188391, 3.812716, 4.088717, 5.666996, 
    7.943676,
  4.598904, 3.263204, 2.682703, 2.344065, 2.580417, 3.256469, 3.681463, 
    4.480714, 4.79798, 5.103074, 5.023545, 4.095044, 3.779275, 4.829471, 
    7.364823,
  3.79999, 3.152031, 2.705509, 2.438466, 2.674974, 3.32763, 3.959683, 
    4.058691, 4.434918, 5.417962, 5.66346, 5.026763, 3.8974, 3.973474, 
    6.358493,
  3.696028, 3.147691, 2.655031, 2.481473, 2.677408, 3.274318, 3.886217, 
    4.500121, 5.121153, 5.706736, 6.165517, 5.633776, 4.387786, 3.533802, 
    5.261613,
  3.778836, 3.157418, 2.639052, 2.4364, 2.676336, 3.18018, 3.777841, 
    4.427625, 5.214302, 5.98966, 6.469923, 6.189132, 4.875529, 3.625152, 
    4.222855,
  3.912805, 3.138038, 2.54085, 2.360011, 2.580991, 3.03179, 3.593094, 
    4.166026, 4.869706, 5.815976, 6.512106, 6.756327, 5.661013, 3.842893, 
    3.567004,
  4.250782, 3.202864, 2.419354, 2.263978, 2.456391, 2.772592, 3.26143, 
    3.907244, 4.502256, 5.278383, 6.26334, 6.809597, 6.855027, 5.197858, 
    3.448346,
  4.570018, 3.375631, 2.521736, 2.225953, 2.315838, 2.557047, 2.927801, 
    3.5077, 4.125992, 4.766135, 5.59295, 6.556297, 6.994155, 6.831508, 
    5.023937,
  6.350302, 5.72562, 4.567909, 3.057617, 3.199033, 4.400226, 5.124045, 
    5.341657, 5.457307, 5.369331, 4.80918, 4.440909, 4.344868, 4.533328, 
    5.210587,
  4.973193, 4.192032, 3.114161, 3.04476, 3.874737, 4.714897, 5.229075, 
    5.393322, 5.583764, 5.709289, 5.080814, 4.496292, 4.235508, 4.099822, 
    5.542073,
  3.160149, 3.043683, 3.095636, 3.547371, 4.158083, 4.327519, 5.065696, 
    5.47828, 5.718697, 5.82546, 5.267461, 4.430523, 4.084139, 4.356663, 
    6.681802,
  3.136312, 3.24025, 3.409273, 3.696568, 4.089119, 4.339642, 4.478139, 
    5.258616, 5.596698, 5.926742, 5.342263, 4.249402, 3.945065, 4.830597, 
    7.375652,
  3.247619, 3.298428, 3.445845, 3.622361, 3.841468, 4.036067, 4.474403, 
    4.326298, 4.769092, 5.865235, 5.521691, 4.238805, 4.012156, 5.187053, 
    7.497765,
  3.148905, 3.217304, 3.199059, 3.404653, 3.563971, 3.653656, 4.145589, 
    4.764382, 5.46772, 5.939923, 5.856909, 4.486434, 3.988962, 5.097822, 
    7.331429,
  3.027417, 2.986433, 2.877722, 3.005196, 3.326825, 3.351944, 3.687102, 
    4.416773, 5.287983, 5.984889, 6.067017, 5.280947, 4.240752, 4.812168, 
    6.763542,
  3.484714, 2.904515, 2.554263, 2.595331, 3.000307, 3.082877, 3.347943, 
    3.889396, 4.626634, 5.630136, 6.079435, 5.895865, 4.843365, 4.528142, 
    6.230238,
  4.562276, 3.481507, 2.454605, 2.362693, 2.86063, 2.976278, 3.158226, 
    3.577785, 4.13092, 5.074824, 5.869604, 6.237959, 5.693004, 4.794134, 
    5.290415,
  5.337339, 4.341003, 2.924016, 2.474495, 2.878481, 3.030117, 3.136792, 
    3.361887, 3.693266, 4.390425, 5.339103, 6.138981, 6.244041, 5.511278, 
    4.831258,
  3.723861, 3.862599, 3.808548, 3.862782, 4.132409, 4.348326, 4.637301, 
    4.9793, 5.39051, 5.443401, 5.300668, 4.876699, 4.533432, 4.338349, 
    4.300478,
  3.820432, 3.933875, 3.758938, 3.649965, 3.742074, 3.88575, 4.333476, 
    4.740706, 5.230805, 5.472516, 5.270621, 4.722455, 4.407562, 3.942297, 
    3.990998,
  3.83909, 3.942585, 3.676576, 3.364746, 3.338852, 3.246246, 3.8956, 
    4.602273, 5.141907, 5.493045, 5.245322, 4.805157, 4.584448, 4.614549, 
    5.331467,
  3.774119, 3.671292, 3.443508, 3.130291, 3.175876, 3.294768, 3.393244, 
    4.178302, 4.774431, 5.436822, 5.330017, 5.106404, 4.939578, 5.341556, 
    6.196619,
  3.755534, 3.368829, 3.150214, 2.951604, 3.130647, 3.272747, 3.602834, 
    3.481642, 4.01655, 5.300421, 5.49718, 5.390389, 5.274856, 5.86565, 6.7096,
  3.935062, 3.267094, 2.866745, 2.841465, 3.161704, 3.305551, 3.622177, 
    4.029039, 4.644864, 5.293329, 5.573329, 5.58738, 5.606602, 6.25662, 
    6.917272,
  4.280797, 3.389571, 2.899544, 2.87579, 3.291631, 3.406836, 3.588976, 
    3.92581, 4.525057, 5.186847, 5.535639, 5.721312, 5.818935, 6.315932, 
    6.800651,
  4.589187, 3.773701, 3.244163, 3.002822, 3.478827, 3.553595, 3.607819, 
    3.689394, 3.969851, 4.752922, 5.398486, 5.756766, 5.905364, 6.160538, 
    6.531294,
  5.25848, 4.706454, 3.877631, 3.272702, 3.695086, 3.765875, 3.726037, 
    3.598398, 3.650437, 4.204259, 5.077169, 5.762227, 5.949746, 6.007783, 
    6.105289,
  5.510703, 5.100885, 4.462836, 3.616229, 3.900724, 4.022763, 3.903547, 
    3.552798, 3.424816, 3.648348, 4.56239, 5.567086, 5.964149, 5.893229, 
    5.630362,
  3.515729, 3.25887, 3.102432, 3.059436, 3.211041, 3.411878, 3.743125, 
    4.073208, 4.471073, 4.810862, 4.94919, 5.177694, 5.068556, 4.88563, 
    4.726756,
  3.732205, 3.274203, 3.114689, 3.090453, 3.284049, 3.417507, 3.739858, 
    3.91199, 4.188426, 4.661874, 4.868846, 5.15728, 5.207987, 4.954566, 
    4.917164,
  4.277629, 3.364885, 3.274544, 3.240288, 3.375644, 3.134811, 3.548086, 
    3.807502, 3.98641, 4.38414, 4.688457, 5.08346, 5.355931, 5.452112, 
    5.426034,
  4.718477, 3.350368, 3.455396, 3.459748, 3.631712, 3.546824, 3.146874, 
    3.397091, 3.481552, 4.069399, 4.498735, 4.959774, 5.376658, 5.500025, 
    5.499713,
  4.757939, 3.420001, 3.718678, 3.736843, 3.84478, 3.715595, 3.427455, 
    2.773153, 2.758204, 3.745333, 4.340508, 4.84997, 5.315141, 5.429391, 
    5.589932,
  4.290867, 3.653575, 3.982241, 3.954586, 4.054982, 3.878931, 3.473472, 
    3.213261, 3.17261, 3.552911, 4.214148, 4.810838, 5.176023, 5.208537, 
    5.422831,
  4.11245, 4.059583, 4.370005, 4.125602, 4.240799, 4.11605, 3.561053, 
    3.173044, 3.104141, 3.398776, 4.131972, 4.769953, 5.047933, 4.941909, 
    5.108086,
  4.28515, 4.472439, 4.790903, 4.352495, 4.382009, 4.370584, 3.776546, 
    3.168025, 2.981417, 3.246324, 4.060116, 4.717999, 4.881959, 4.550092, 
    4.700723,
  4.884003, 5.093466, 5.274498, 4.736913, 4.668046, 4.587744, 4.058814, 
    3.319362, 3.007473, 3.158207, 3.978078, 4.667572, 4.707645, 4.30073, 
    4.187574,
  5.338248, 5.714281, 5.830571, 5.351211, 5.047744, 4.793498, 4.311518, 
    3.487074, 3.089225, 3.130893, 3.890235, 4.636199, 4.587263, 4.221615, 
    3.971613,
  3.260335, 3.600207, 3.876246, 3.966507, 4.006679, 3.887808, 3.614661, 
    3.372159, 3.263116, 3.214326, 3.346262, 3.616633, 3.973162, 4.337355, 
    4.671113,
  3.665048, 4.034414, 4.319392, 4.400639, 4.38052, 4.101155, 3.770457, 
    3.412883, 3.148922, 3.212449, 3.311289, 3.514286, 3.889128, 3.993467, 
    4.384483,
  4.095064, 4.469721, 4.827999, 4.889021, 4.798652, 4.073195, 3.970737, 
    3.715029, 3.40271, 3.270767, 3.280509, 3.461918, 3.78806, 4.121643, 
    4.430967,
  4.44193, 4.948828, 5.31534, 5.336332, 5.265059, 4.92484, 3.991894, 
    3.864523, 3.505958, 3.434685, 3.40166, 3.487845, 3.773338, 4.042381, 
    4.297602,
  5.01015, 5.628889, 5.893338, 5.805709, 5.635029, 5.358533, 4.857839, 
    3.590969, 3.169784, 3.578531, 3.615969, 3.664919, 3.852125, 3.97226, 
    4.177942,
  5.678376, 6.199644, 6.302214, 6.063426, 5.693528, 5.354315, 5.045112, 
    4.656531, 4.300896, 4.019504, 3.856061, 3.831855, 3.942735, 4.021016, 
    4.065767,
  6.219377, 6.408194, 6.18927, 5.815124, 5.341372, 5.075509, 5.008593, 
    4.95377, 4.621851, 4.212658, 3.977906, 3.948317, 4.017429, 4.036192, 
    4.011262,
  6.346081, 6.089041, 5.738266, 5.417017, 5.055758, 4.914949, 5.027441, 
    5.068181, 4.798757, 4.340941, 3.990038, 3.953712, 3.997936, 3.972698, 
    3.971011,
  6.130648, 5.625319, 5.303728, 5.044803, 4.812641, 4.784123, 4.922358, 
    4.910172, 4.543625, 4.059396, 3.879295, 3.99451, 4.013956, 3.983623, 
    3.94085,
  5.865272, 5.176413, 4.838305, 4.60112, 4.436862, 4.462263, 4.587355, 
    4.518293, 4.22046, 3.976176, 3.929609, 4.158832, 4.073737, 4.000705, 
    4.031787,
  5.645579, 5.341863, 5.162006, 5.050932, 5.057148, 5.090675, 5.114978, 
    5.133607, 5.086522, 4.793546, 4.342838, 3.749768, 3.330108, 3.244886, 
    3.740754,
  5.743076, 5.527085, 5.481627, 5.562502, 5.654428, 5.671617, 5.749223, 
    5.658506, 5.490042, 5.275295, 4.899801, 4.278833, 3.545024, 3.044071, 
    3.386955,
  5.805978, 5.746578, 5.770576, 5.756599, 5.804108, 5.265975, 5.786347, 
    6.039828, 5.948762, 5.705729, 5.312792, 4.766472, 3.903595, 3.367682, 
    3.340101,
  5.904741, 5.740623, 5.514417, 5.264025, 5.180243, 5.151676, 4.602461, 
    5.126908, 5.587344, 5.84271, 5.624556, 5.170143, 4.389188, 3.601645, 
    3.366311,
  5.62276, 5.3639, 4.956474, 4.619962, 4.440424, 4.272322, 4.233459, 
    3.392412, 3.458329, 4.913641, 5.400998, 5.221714, 4.674643, 3.823371, 
    3.471255,
  5.214697, 4.859095, 4.431343, 4.172096, 4.011231, 3.885393, 3.78741, 
    3.71606, 3.830062, 4.277866, 4.999647, 5.124363, 4.785045, 4.013859, 
    3.629922,
  4.833889, 4.549791, 4.311646, 4.330655, 4.274099, 4.204374, 4.11994, 
    4.154055, 4.124629, 4.189389, 4.560622, 4.932455, 4.713439, 4.152057, 
    3.786437,
  4.666982, 4.571093, 4.495732, 4.648551, 4.619423, 4.601491, 4.625227, 
    4.541663, 4.511611, 4.507591, 4.617045, 4.80301, 4.619507, 4.132971, 
    3.833056,
  4.62216, 4.631789, 4.668494, 4.874087, 4.850365, 4.887334, 4.898212, 
    4.757218, 4.413251, 4.393976, 4.589824, 4.663985, 4.486282, 4.053871, 
    3.873875,
  4.524087, 4.617547, 4.729641, 4.914301, 4.950911, 5.036834, 5.108912, 
    5.129434, 4.701734, 4.285835, 4.433927, 4.486424, 4.300532, 3.973318, 
    3.885531,
  4.904961, 4.96518, 4.988471, 4.949974, 4.905694, 4.879106, 4.857978, 
    4.885207, 4.823367, 4.719929, 4.757766, 4.721573, 4.278291, 3.67346, 
    3.474303,
  5.334442, 5.374065, 5.375272, 5.307581, 5.143581, 4.883903, 4.823239, 
    4.87604, 4.953413, 4.89465, 4.855731, 4.932199, 4.615148, 3.63171, 
    3.340104,
  5.887897, 5.939816, 5.886685, 5.72801, 5.488479, 4.604633, 4.624527, 
    4.544629, 4.695958, 4.969909, 5.028634, 5.108093, 4.997837, 4.05968, 
    3.471101,
  6.283679, 6.151695, 6.033305, 5.856833, 5.62458, 5.264723, 4.299045, 
    4.202639, 4.105065, 4.606179, 5.121023, 5.31674, 5.280275, 4.341761, 
    3.500173,
  6.253937, 6.018162, 5.825492, 5.570728, 5.247132, 5.081073, 4.807581, 
    3.730586, 3.255375, 3.816442, 4.867839, 5.422654, 5.481702, 4.588939, 
    3.623611,
  5.94484, 5.603034, 5.435987, 5.010907, 4.73472, 4.720449, 4.706877, 
    4.557039, 4.187572, 3.908217, 4.539734, 5.44937, 5.610875, 4.608809, 
    3.783116,
  5.438511, 5.253666, 4.957055, 4.687739, 4.626975, 4.644791, 4.730006, 
    4.801519, 4.685439, 4.027876, 4.249475, 5.427367, 5.586824, 4.525873, 
    4.007368,
  5.083523, 4.897691, 4.676817, 4.667237, 4.658234, 4.706506, 4.692973, 
    4.773508, 4.738634, 4.099674, 4.22014, 5.437355, 5.445556, 4.377789, 
    4.034353,
  4.816869, 4.699262, 4.679294, 4.750573, 4.763626, 4.788539, 4.705624, 
    4.828766, 4.693625, 4.048247, 4.341983, 5.392386, 5.169812, 4.176078, 
    3.92328,
  4.661254, 4.586048, 4.677097, 4.772995, 4.777868, 4.785809, 4.77491, 
    4.833738, 4.369337, 4.027867, 4.656433, 5.285141, 4.831546, 4.001218, 
    3.84088,
  7.365091, 6.757993, 6.600976, 6.527381, 6.201225, 5.74603, 5.326058, 
    5.078353, 5.14316, 4.962692, 4.810902, 4.75011, 4.505614, 4.407472, 
    4.486797,
  6.613076, 6.152416, 6.165214, 6.385278, 6.351649, 6.166819, 5.927188, 
    5.408929, 5.189913, 5.13938, 4.963457, 4.739398, 4.445029, 4.124263, 
    4.26354,
  6.427453, 6.170388, 6.1847, 6.3809, 6.395211, 5.557898, 6.00842, 5.786137, 
    5.253263, 5.126643, 4.982383, 4.731596, 4.466168, 4.2753, 4.190828,
  6.223752, 5.944758, 5.818277, 5.822319, 5.940353, 5.907414, 5.302417, 
    5.56259, 5.218753, 5.018541, 4.967547, 4.723448, 4.486187, 4.219774, 
    3.967954,
  5.651186, 5.310864, 5.156356, 4.956841, 4.66438, 4.809893, 5.33762, 
    4.502073, 4.025147, 4.781906, 4.884277, 4.7256, 4.550387, 4.166806, 
    3.872601,
  5.101122, 4.933659, 4.905094, 4.591056, 4.206134, 4.16229, 4.739466, 
    5.038569, 4.717037, 4.721127, 4.714568, 4.701592, 4.591221, 4.123535, 
    3.924387,
  4.743028, 4.673593, 4.553111, 4.646507, 4.482783, 4.241437, 4.502053, 
    4.991091, 4.715879, 4.601959, 4.617946, 4.708406, 4.570684, 4.127833, 
    4.293896,
  4.462336, 4.390492, 4.347994, 4.593939, 4.63694, 4.466556, 4.624622, 
    4.769295, 4.572564, 4.513674, 4.606329, 4.751549, 4.534109, 4.28196, 
    4.520133,
  4.23211, 4.213715, 4.292699, 4.467487, 4.645226, 4.530768, 4.575742, 
    4.633207, 4.569987, 4.49176, 4.675977, 4.809297, 4.519726, 4.349548, 
    4.580296,
  4.12027, 4.157318, 4.325047, 4.43898, 4.526987, 4.515809, 4.538509, 
    4.581897, 4.558224, 4.566977, 4.809955, 4.818799, 4.479299, 4.369402, 
    4.773652,
  7.737146, 6.529377, 5.984783, 5.709911, 5.766935, 5.808616, 5.703575, 
    5.386406, 5.230023, 5.09997, 4.541944, 4.625045, 5.16672, 5.378985, 
    6.529498,
  6.771561, 6.259799, 5.922708, 5.69232, 5.662364, 5.740369, 5.731805, 
    5.362831, 5.163367, 5.208485, 4.798387, 4.666283, 4.974457, 5.196705, 
    6.230307,
  6.070923, 5.802882, 5.536706, 5.229709, 5.320487, 4.873766, 5.660914, 
    5.583327, 5.345354, 5.302098, 4.887243, 4.609983, 4.861804, 5.407516, 
    6.127517,
  5.353127, 5.129279, 4.966989, 4.880117, 5.11136, 5.450459, 5.056768, 
    5.570153, 5.430125, 5.311273, 4.969409, 4.521237, 4.743463, 5.213262, 
    5.758957,
  4.96611, 4.780544, 4.694907, 4.816522, 4.987415, 5.189332, 5.672471, 
    4.623959, 4.35796, 5.276621, 5.015587, 4.553001, 4.65533, 4.980824, 
    5.410345,
  4.474443, 4.444588, 4.445178, 4.546022, 4.727551, 4.420051, 5.176431, 
    5.458263, 5.249008, 5.301681, 4.915933, 4.542407, 4.568287, 4.826317, 
    5.216648,
  4.2979, 4.271456, 4.099177, 4.316322, 4.633866, 4.134239, 4.338233, 
    5.47186, 5.461203, 5.201215, 4.803629, 4.470585, 4.449139, 4.661764, 
    5.018309,
  4.146197, 4.08303, 4.067307, 4.181546, 4.525417, 4.109324, 4.387781, 
    5.242989, 5.316694, 5.076937, 4.71204, 4.409579, 4.356817, 4.448301, 
    4.694037,
  4.095007, 4.154604, 4.255568, 4.315868, 4.421647, 4.300401, 4.67797, 
    5.223461, 5.249936, 4.93914, 4.537024, 4.297607, 4.235783, 4.297802, 
    4.399486,
  4.138333, 4.247146, 4.411246, 4.407332, 4.459051, 4.530012, 4.883239, 
    5.111829, 5.025206, 4.688035, 4.324116, 4.17315, 4.140559, 4.148382, 
    4.266022,
  6.454898, 6.133728, 5.988581, 5.763577, 5.563638, 5.353765, 5.151044, 
    5.112419, 5.131438, 5.075381, 4.787569, 4.568731, 4.232384, 4.649711, 
    6.380251,
  6.112068, 5.816357, 5.73906, 5.689065, 5.451842, 5.204311, 5.227968, 
    5.21128, 5.121281, 5.147334, 4.842844, 4.485516, 4.474018, 5.469603, 
    7.293863,
  5.703559, 5.524366, 5.459242, 5.40651, 5.255918, 4.515402, 5.053722, 
    5.333293, 5.071553, 5.015274, 4.600283, 4.381247, 5.082631, 6.854538, 
    8.14941,
  5.207517, 5.186015, 5.129498, 5.06672, 5.007881, 5.07704, 4.342777, 
    5.011696, 5.039913, 5.070506, 4.667897, 4.693065, 6.105479, 7.604679, 
    8.041313,
  4.982486, 4.915493, 4.867216, 4.774, 4.748719, 4.848441, 4.956756, 
    3.859943, 3.832769, 4.938858, 4.750786, 5.457305, 6.998991, 7.707048, 
    7.340201,
  4.743904, 4.632926, 4.585577, 4.406107, 4.558769, 4.678853, 4.992074, 
    4.959479, 5.00368, 4.976371, 5.177407, 6.414291, 7.2258, 7.385285, 
    6.573813,
  4.54472, 4.422526, 4.251813, 4.232496, 4.614414, 4.543532, 5.081217, 
    5.365733, 5.037811, 5.183541, 5.935826, 6.708457, 7.120233, 6.894979, 
    6.390262,
  4.40116, 4.260923, 4.117637, 4.436627, 4.550867, 4.739592, 5.314936, 
    5.288487, 5.099141, 5.491738, 6.054403, 6.572533, 6.71263, 6.546977, 
    6.288923,
  4.308788, 4.309851, 4.25326, 4.455868, 4.678823, 4.959595, 5.328736, 
    5.222025, 5.151235, 5.490984, 5.925474, 6.22959, 6.264941, 6.248329, 
    6.121205,
  4.29006, 4.311852, 4.381712, 4.507974, 4.726516, 4.992727, 5.175085, 
    5.051923, 5.062601, 5.313941, 5.641682, 5.877026, 5.93412, 5.945551, 
    5.872939,
  9.91676, 8.681334, 7.570251, 7.057368, 6.662328, 6.259919, 5.837415, 
    5.633996, 5.37397, 5.011986, 4.908548, 4.9737, 5.044823, 4.737542, 
    4.361891,
  8.007552, 7.094957, 6.335136, 6.067854, 5.849843, 5.648045, 5.621027, 
    5.518122, 5.439791, 5.387284, 5.304078, 5.186845, 5.040203, 4.446685, 
    4.305575,
  6.391769, 5.471362, 5.153695, 5.216238, 5.077105, 4.403244, 4.846238, 
    5.134021, 5.136679, 5.163553, 5.195993, 5.131356, 4.917668, 4.670752, 
    4.611365,
  5.139633, 5.087931, 5.115446, 5.095452, 4.973137, 4.821455, 4.13129, 
    4.545197, 4.835531, 5.011731, 5.082733, 5.000282, 4.784405, 4.725583, 
    5.105031,
  5.443956, 5.363492, 5.137588, 4.80406, 4.468796, 4.297644, 4.312502, 
    3.437676, 3.392908, 4.362968, 4.753006, 4.721605, 4.732525, 5.139842, 
    5.771992,
  5.530918, 5.080518, 4.743664, 4.352135, 4.159997, 4.179133, 4.298861, 
    4.29824, 4.467036, 4.680048, 4.759135, 4.860395, 5.270569, 5.820667, 
    6.27603,
  4.973516, 4.658693, 4.169661, 4.191694, 4.34237, 4.396708, 4.480956, 
    4.673331, 4.708027, 4.771197, 5.158909, 5.615027, 6.073687, 6.370062, 
    6.246532,
  4.576488, 4.345528, 4.149171, 4.550009, 4.593574, 4.789037, 4.890808, 
    4.898081, 5.096138, 5.634343, 6.053996, 6.385904, 6.485511, 6.077157, 
    5.599658,
  4.347379, 4.390892, 4.577147, 4.818981, 4.919194, 4.986563, 5.16348, 
    5.581879, 6.191033, 6.515849, 6.620044, 6.435991, 5.913018, 5.513733, 
    5.412901,
  4.346294, 4.562497, 4.777995, 4.885877, 5.046092, 5.38453, 5.834748, 
    6.323254, 6.632944, 6.652816, 6.298483, 5.852717, 5.534607, 5.566853, 
    5.955554,
  14.25839, 12.0587, 10.19456, 8.81566, 7.465001, 6.51498, 5.978764, 
    5.683898, 5.411996, 5.166315, 5.117714, 5.065052, 5.211934, 5.062954, 
    4.623506,
  13.5517, 11.4843, 9.831657, 8.543782, 7.201745, 6.235527, 5.794151, 
    5.400924, 5.162457, 5.061801, 5.241858, 5.37996, 5.277854, 4.815022, 
    4.753751,
  13.02184, 11.18564, 9.557681, 8.14857, 6.815971, 5.223881, 5.039282, 
    4.833417, 4.60472, 4.624196, 4.962154, 5.374606, 5.49115, 5.286669, 
    5.047768,
  11.76427, 10.14912, 8.585298, 7.207009, 6.087895, 5.054202, 3.902477, 
    4.106472, 4.075791, 4.249837, 4.552721, 5.056479, 5.377128, 5.323848, 
    5.103245,
  10.082, 8.857173, 7.514538, 5.963575, 4.94653, 4.512905, 4.348728, 
    3.417743, 3.207625, 3.999749, 4.427582, 4.883243, 5.193317, 5.202284, 
    5.03586,
  8.545545, 7.177582, 5.762927, 4.783533, 4.455729, 4.588031, 4.591221, 
    4.469538, 4.305488, 4.321416, 4.575871, 4.845863, 5.074514, 5.009318, 
    4.760628,
  6.385391, 5.198792, 4.539752, 4.356009, 4.725857, 4.846497, 4.794483, 
    4.623126, 4.416979, 4.324417, 4.467766, 4.582718, 4.69702, 4.695924, 
    4.5835,
  4.724068, 4.290424, 4.294516, 4.865283, 4.982933, 4.847928, 4.672143, 
    4.489811, 4.354525, 4.201954, 4.255902, 4.307055, 4.472601, 4.632967, 
    4.81926,
  4.088384, 4.343897, 4.944896, 5.135736, 5.01209, 4.683917, 4.350206, 
    4.283563, 4.215791, 4.121438, 4.292933, 4.569987, 4.83741, 5.017484, 
    5.225212,
  4.342873, 4.943076, 5.238365, 5.276264, 5.10355, 4.775677, 4.567297, 
    4.591781, 4.627245, 4.749668, 5.099713, 5.299963, 5.44556, 5.577622, 
    5.777683,
  14.92711, 15.56124, 15.94728, 16.08604, 16.2338, 16.21742, 15.88408, 
    15.2681, 14.16973, 12.70134, 11.11051, 9.565188, 8.214218, 6.968133, 
    5.896882,
  15.26112, 15.7982, 16.17705, 16.453, 16.29861, 15.78514, 15.24884, 
    14.23203, 12.96213, 11.5138, 9.781942, 8.188803, 7.168466, 6.009943, 
    5.399935,
  15.2691, 15.82137, 16.31325, 16.4332, 15.91051, 13.8019, 13.57785, 
    12.31722, 10.90788, 9.466555, 7.988022, 6.633594, 6.077169, 5.748258, 
    5.195291,
  14.98912, 15.69788, 16.10773, 15.92182, 15.00657, 13.48691, 10.39107, 
    9.668763, 8.621585, 7.411311, 6.24148, 5.289453, 5.092775, 5.214893, 
    5.009505,
  13.7308, 14.46736, 14.50619, 13.9038, 12.47086, 10.57706, 8.507162, 
    6.08104, 4.994293, 5.431067, 4.648853, 4.281864, 4.372118, 4.802164, 
    4.87442,
  12.23363, 12.48937, 11.92989, 10.60993, 8.849778, 6.898891, 5.195059, 
    4.330599, 4.158777, 4.128959, 3.904293, 4.073164, 4.409044, 4.773659, 
    4.841393,
  9.805511, 9.220256, 8.033762, 6.478859, 4.901488, 4.031652, 3.873914, 
    3.886722, 3.742202, 3.699906, 3.84608, 4.196628, 4.666749, 4.889272, 
    4.808403,
  6.955925, 6.078982, 5.080926, 4.240249, 3.810723, 3.64126, 3.553493, 
    3.522224, 3.582758, 3.812558, 4.147591, 4.568031, 4.833432, 4.883451, 
    4.605137,
  5.589452, 5.004654, 4.384403, 3.955256, 3.6868, 3.662923, 3.679143, 
    3.650305, 3.59613, 3.792216, 4.127898, 4.385868, 4.535621, 4.444816, 
    4.095449,
  5.207161, 4.74313, 4.248806, 3.770014, 3.663226, 3.808493, 3.985449, 
    4.031107, 3.909292, 3.905911, 4.024631, 4.118791, 4.130126, 4.026196, 
    4.18175,
  6.406841, 6.502863, 7.297863, 8.50077, 9.342686, 9.788377, 10.07452, 
    10.4408, 10.88995, 11.15791, 11.52492, 12.0178, 12.39925, 12.49783, 
    12.35966,
  6.327606, 6.910822, 8.251599, 9.554957, 10.41565, 10.88872, 11.65674, 
    12.15791, 12.52954, 12.7978, 12.97083, 13.15335, 13.173, 12.32384, 
    12.01575,
  6.54783, 7.589495, 8.919974, 10.14889, 11.07008, 10.6256, 12.10405, 
    11.9083, 12.22012, 12.31334, 12.59216, 12.73688, 12.68415, 12.39269, 
    11.73122,
  6.877821, 7.947773, 9.054444, 9.972845, 11.22336, 11.40896, 9.365358, 
    9.725252, 10.14659, 10.54768, 10.80825, 11.17812, 11.5934, 11.32414, 
    10.56003,
  6.944764, 7.848419, 8.566441, 8.901286, 9.01792, 8.697894, 8.102155, 
    6.670927, 6.017432, 7.225636, 7.851842, 8.78935, 9.475686, 9.528082, 
    8.980897,
  6.526364, 6.769727, 6.837582, 6.812466, 6.271908, 5.432793, 4.711087, 
    4.330375, 4.310472, 4.764688, 5.291905, 6.049708, 6.944332, 7.447816, 
    7.173189,
  5.756582, 5.455112, 5.024112, 4.417832, 3.748029, 3.362339, 3.330996, 
    3.503883, 3.834767, 4.193734, 4.474915, 4.832458, 5.31206, 5.715576, 
    5.594507,
  4.960908, 4.323965, 3.957264, 3.90351, 3.769643, 3.64238, 3.560959, 
    3.565536, 3.852767, 4.167441, 4.360111, 4.490434, 4.640176, 4.797982, 
    4.749737,
  4.479569, 3.852681, 3.729327, 3.973881, 4.042306, 3.950278, 3.916146, 
    3.935318, 4.164358, 4.341557, 4.418484, 4.427548, 4.390243, 4.400733, 
    4.502315,
  4.183875, 3.702713, 3.810911, 4.107583, 4.235698, 4.155559, 3.977592, 
    3.912816, 4.143863, 4.334997, 4.36992, 4.331061, 4.258773, 4.313108, 
    4.879168,
  11.87718, 10.84641, 9.415943, 8.105849, 7.726443, 7.451804, 6.663894, 
    6.14194, 5.851572, 5.809385, 6.110537, 6.545533, 6.938434, 7.250404, 
    7.528633,
  10.67969, 9.78655, 8.765121, 7.688109, 7.061717, 6.481697, 5.821086, 
    5.385719, 5.220702, 5.486007, 6.069254, 6.903296, 7.717189, 7.985627, 
    8.422994,
  9.630642, 8.69885, 7.809747, 6.806912, 5.969285, 4.8864, 4.797205, 
    4.558881, 4.402559, 4.689988, 5.313138, 6.449, 7.994613, 9.292412, 
    9.770539,
  9.050932, 7.902633, 6.859334, 5.870042, 5.055161, 4.313527, 3.668785, 
    3.966835, 3.794995, 4.16129, 4.542437, 5.89594, 8.116668, 10.24394, 
    10.6792,
  7.883391, 6.713309, 5.761917, 4.913359, 4.374357, 4.206329, 4.055738, 
    3.215897, 3.092017, 3.825855, 4.022261, 5.461868, 8.270976, 10.94708, 
    11.14855,
  6.169166, 5.27736, 4.60196, 4.307763, 4.230525, 4.295691, 4.441974, 
    4.344877, 4.10399, 3.804363, 3.883984, 5.352706, 8.381677, 10.55691, 
    11.01026,
  4.672012, 4.210062, 3.973295, 4.121174, 4.256137, 4.355152, 4.445066, 
    4.479923, 4.232611, 3.856136, 3.973088, 5.60334, 8.088505, 9.705275, 
    10.28239,
  4.495276, 4.025907, 3.769669, 3.899469, 4.182022, 4.357625, 4.416538, 
    4.363548, 4.12494, 3.871874, 4.232677, 5.857615, 7.621554, 8.695663, 
    9.040557,
  4.916933, 4.171326, 3.710753, 4.099985, 4.575397, 4.684451, 4.487733, 
    4.280056, 4.065333, 3.972042, 4.516943, 6.00314, 7.319695, 7.983075, 
    7.843089,
  4.984563, 3.959607, 4.063638, 4.790043, 5.041988, 4.924786, 4.493426, 
    4.143205, 3.94471, 4.076817, 4.855137, 6.028255, 6.937554, 7.280705, 
    7.073916,
  5.645211, 6.22536, 7.316525, 8.706092, 9.876219, 10.24849, 10.15101, 
    9.810396, 9.325989, 8.687154, 7.786312, 6.540882, 5.334816, 4.459507, 
    4.192348,
  6.1373, 6.519025, 7.295702, 8.45642, 9.588531, 9.796331, 9.953561, 9.49263, 
    8.858642, 8.160971, 7.100102, 5.790068, 4.748821, 3.940357, 3.945763,
  6.352936, 6.71165, 7.364269, 8.347695, 9.382658, 8.732018, 9.460976, 
    8.781923, 7.958169, 7.169524, 6.125195, 5.00477, 4.23031, 3.924736, 
    4.881356,
  6.185966, 6.479761, 7.188025, 7.953534, 8.781305, 8.829353, 7.395727, 
    7.476087, 6.860694, 6.137423, 5.223866, 4.354841, 3.863335, 4.644472, 
    7.145609,
  5.650807, 5.713009, 6.117877, 6.655562, 7.163571, 7.344553, 6.838038, 
    5.639966, 5.037206, 5.212156, 4.460094, 3.793242, 4.335318, 7.089856, 
    9.169235,
  5.20575, 4.926644, 4.890823, 5.101312, 5.389118, 5.643286, 5.730948, 
    5.420663, 4.969615, 4.500037, 3.81045, 3.912547, 6.046873, 8.81863, 
    9.144388,
  5.090919, 4.479067, 4.108217, 4.087193, 4.129742, 4.213086, 4.377671, 
    4.518314, 4.399242, 3.876523, 3.712515, 5.043984, 7.337705, 9.098948, 
    9.322627,
  5.349814, 4.740298, 4.201581, 4.204046, 4.21511, 4.210343, 4.181389, 
    4.172451, 3.964236, 3.466438, 4.372652, 6.510089, 7.975109, 8.912865, 
    9.403912,
  5.744631, 5.313735, 4.848169, 4.931746, 5.007771, 4.940822, 4.731026, 
    4.370461, 3.685256, 3.750806, 5.910151, 7.483013, 8.183906, 8.58112, 
    8.414654,
  6.034657, 5.812436, 5.65065, 5.624492, 5.474593, 5.260741, 5.034436, 
    4.467406, 3.577926, 4.845999, 6.997901, 7.656367, 7.777878, 7.477937, 
    6.979175,
  7.951498, 7.513463, 6.911177, 5.953385, 5.234849, 5.648501, 6.590209, 
    7.184837, 7.874704, 8.056597, 8.35977, 8.978299, 9.324762, 8.723623, 
    7.671206,
  8.304208, 7.943293, 7.066955, 5.611001, 4.835987, 5.326079, 6.404516, 
    6.922851, 7.615361, 8.178694, 8.456458, 8.632527, 8.280547, 6.862574, 
    5.657233,
  9.232435, 8.361935, 6.971067, 4.929842, 4.54726, 4.701662, 5.924069, 
    6.586136, 7.210093, 7.703035, 7.705317, 7.381028, 6.287932, 5.209817, 
    4.509595,
  9.069743, 8.030821, 6.276868, 4.619741, 4.494102, 4.827186, 5.168734, 
    5.966688, 6.471679, 7.028198, 6.784283, 6.071615, 5.35619, 4.889267, 
    5.53784,
  7.976321, 7.061646, 5.80267, 4.73097, 4.559778, 4.649159, 5.125392, 
    4.938761, 5.259436, 6.67892, 6.651831, 6.161251, 5.94315, 6.613822, 
    7.614305,
  6.768383, 6.46911, 6.014529, 5.435952, 4.917388, 4.517385, 4.595988, 
    4.99872, 5.412334, 6.343759, 6.533993, 6.44992, 6.81232, 7.443212, 7.40584,
  6.491027, 6.706947, 6.670849, 6.263195, 5.639882, 4.939798, 4.404051, 
    4.546126, 4.909741, 5.861611, 6.496101, 6.751183, 7.317802, 7.666093, 
    7.51304,
  6.618378, 6.892859, 6.851322, 6.608001, 6.186615, 5.502665, 4.687781, 
    4.147897, 4.350819, 5.592326, 6.384091, 7.027702, 7.965723, 8.354622, 
    8.193735,
  6.60008, 6.561589, 6.431935, 6.371294, 6.272141, 5.766974, 5.160736, 
    4.364795, 4.203849, 5.506183, 6.219014, 6.998195, 7.843205, 8.270588, 
    8.248079,
  6.232543, 5.930829, 5.867024, 6.111548, 6.402027, 6.146202, 5.463527, 
    4.559544, 4.246175, 5.484103, 6.218317, 6.917245, 7.384332, 7.668101, 
    7.805079,
  11.21254, 10.18999, 9.652748, 8.690535, 7.025981, 5.140681, 4.142202, 
    4.681502, 5.855949, 6.790552, 6.967844, 6.704207, 6.683014, 6.542524, 
    6.88438,
  11.17183, 10.69549, 9.550282, 7.792159, 5.944557, 4.603718, 4.210313, 
    4.63163, 5.876821, 7.205347, 7.216067, 6.954609, 6.877038, 6.484887, 
    6.699941,
  12.00931, 11.048, 8.167379, 6.648224, 5.208882, 4.100545, 4.296981, 
    4.66292, 5.911308, 7.455583, 7.433627, 7.318239, 7.206492, 7.258617, 
    7.319241,
  12.33084, 8.612917, 6.716826, 5.879368, 4.984366, 4.607142, 4.053739, 
    4.31954, 5.516463, 7.347721, 7.51455, 7.526742, 7.345644, 7.322522, 
    7.34995,
  9.122158, 6.764294, 6.484012, 5.901103, 5.446709, 5.156208, 4.983652, 
    3.862548, 4.583096, 7.165763, 7.537755, 7.71453, 7.567082, 7.326039, 
    7.287356,
  6.751281, 6.072107, 6.404784, 6.4235, 6.302247, 5.891492, 5.655112, 
    5.107037, 5.265532, 7.091814, 7.501257, 7.880183, 7.895698, 7.764506, 
    7.59742,
  6.090818, 6.025572, 5.971192, 6.286772, 6.752335, 6.700509, 6.395645, 
    5.504986, 5.222978, 6.768857, 7.348418, 7.922085, 8.121777, 8.1679, 
    8.199862,
  5.980147, 5.683405, 5.155097, 5.290477, 5.882596, 6.524509, 6.48078, 
    5.334206, 5.000345, 6.351574, 7.152566, 7.768795, 8.154455, 8.37015, 
    8.526421,
  5.716526, 5.050273, 4.833363, 5.092774, 5.441423, 6.316943, 6.072194, 
    5.056571, 4.992439, 6.126202, 7.08566, 7.70435, 8.1616, 8.469276, 8.704692,
  5.710029, 4.891521, 4.983863, 5.591165, 5.874074, 6.222013, 5.740697, 
    4.992871, 5.178543, 6.250868, 7.273233, 7.835442, 8.240041, 8.557151, 
    8.834479,
  20.79451, 15.37659, 10.38903, 6.970646, 5.49087, 4.733488, 4.316225, 
    4.481107, 5.320235, 6.731403, 7.235433, 7.490223, 7.360777, 7.056675, 
    7.157313,
  16.88919, 11.1945, 7.110333, 5.443195, 4.906168, 4.457899, 4.550391, 
    4.780876, 5.628062, 7.060798, 7.557646, 7.863528, 7.663202, 7.00438, 
    7.121074,
  12.3781, 7.82091, 5.367177, 4.828961, 4.626075, 4.116652, 4.848151, 
    5.296195, 6.100849, 7.34007, 7.888921, 8.285617, 8.096183, 7.789761, 
    7.634924,
  8.7475, 5.646367, 4.661766, 4.582142, 4.664365, 4.644083, 4.61381, 
    5.449522, 6.140476, 7.51286, 8.160366, 8.61409, 8.565245, 8.306074, 
    8.086879,
  6.322541, 4.984122, 4.802955, 4.944048, 5.126644, 5.174501, 5.494435, 
    4.765505, 5.403254, 7.584103, 8.359239, 8.790294, 8.80966, 8.595158, 
    8.445714,
  5.44234, 4.865499, 4.868658, 5.121235, 5.604916, 5.605086, 5.866358, 
    6.197369, 6.833826, 7.885839, 8.557582, 8.885058, 8.880329, 8.665383, 
    8.544341,
  4.969607, 4.596859, 4.595294, 4.920719, 5.346857, 5.744303, 6.070282, 
    6.501028, 7.279092, 8.19098, 8.728001, 8.960433, 8.879791, 8.647281, 
    8.496541,
  4.846715, 4.489848, 4.580245, 4.986428, 5.241496, 5.684112, 6.146392, 
    6.846705, 7.710664, 8.432068, 8.849007, 9.020169, 8.87867, 8.600479, 
    8.412495,
  4.992311, 4.701379, 4.809817, 5.186926, 5.488195, 5.987385, 6.512586, 
    7.29664, 8.122619, 8.633157, 8.972378, 9.105022, 8.909689, 8.577149, 
    8.41651,
  5.223642, 4.806061, 4.796886, 5.176994, 5.588261, 6.266007, 6.919027, 
    7.658834, 8.307208, 8.749331, 9.084118, 9.225747, 8.980615, 8.633263, 
    8.518336,
  8.901625, 6.280758, 5.012523, 4.54322, 4.58328, 5.081033, 5.754296, 
    6.807908, 7.75067, 8.231141, 8.607704, 8.747169, 8.437998, 7.906092, 
    7.705615,
  7.839013, 5.773455, 4.746264, 4.387567, 4.571618, 5.128136, 5.996129, 
    7.046153, 7.865123, 8.423932, 8.740044, 8.785095, 8.403084, 7.563278, 
    7.511995,
  7.362391, 5.521627, 4.559674, 4.331389, 4.652195, 4.788958, 6.264094, 
    7.574373, 8.152235, 8.504476, 8.740373, 8.731754, 8.259433, 7.888075, 
    7.742461,
  6.950035, 5.175382, 4.506569, 4.519342, 5.102665, 5.872084, 6.093966, 
    7.665784, 8.130848, 8.549626, 8.699936, 8.621137, 8.171977, 7.896464, 
    7.847654,
  6.101727, 4.677606, 4.609361, 4.821906, 5.520239, 6.467723, 7.35764, 
    6.844442, 6.997819, 8.435668, 8.661749, 8.539585, 8.146626, 7.947586, 
    7.916438,
  5.037933, 4.461665, 4.640505, 5.217859, 6.061316, 6.9965, 7.769122, 
    8.300303, 8.414065, 8.549982, 8.684397, 8.52818, 8.202316, 8.003149, 
    7.902654,
  4.645627, 4.439081, 4.714848, 5.694064, 6.614119, 7.36055, 7.999432, 
    8.418526, 8.532223, 8.623588, 8.665451, 8.59315, 8.329848, 8.084992, 
    7.854404,
  4.578594, 4.398092, 4.869008, 6.093895, 6.983819, 7.574853, 8.097153, 
    8.38714, 8.478628, 8.565551, 8.678905, 8.736038, 8.551351, 8.283578, 
    7.994193,
  4.63128, 4.373046, 4.941544, 6.282487, 7.209681, 7.634396, 8.105759, 
    8.389924, 8.475291, 8.534037, 8.722226, 8.895736, 8.845812, 8.614042, 
    8.307601,
  4.732073, 4.380177, 4.807125, 6.181642, 7.22507, 7.617026, 8.07965, 
    8.413275, 8.474657, 8.521771, 8.753743, 8.987856, 9.05595, 8.937724, 
    8.706043,
  8.750816, 6.554, 5.152008, 4.685387, 4.991026, 5.665877, 6.416026, 
    7.404755, 7.906817, 8.033364, 8.006537, 7.994047, 7.908805, 7.661142, 
    7.496197,
  7.943386, 5.745392, 4.73993, 4.877424, 5.56841, 6.268767, 7.259295, 
    7.85638, 7.867751, 7.928304, 7.949532, 8.055895, 8.04146, 7.483315, 
    7.385118,
  6.76731, 4.936741, 4.709517, 5.371459, 6.131378, 6.288974, 7.613353, 
    7.981883, 7.7523, 7.771194, 8.011998, 8.268647, 8.216577, 8.054449, 
    7.754943,
  5.504275, 4.595582, 4.896726, 5.75658, 6.659871, 7.322092, 7.160746, 
    7.713319, 7.345947, 7.77157, 8.215401, 8.511453, 8.383269, 8.15681, 
    7.867924,
  4.677254, 4.511967, 5.035873, 6.058106, 7.036881, 7.627298, 7.908986, 
    6.639389, 6.246916, 7.79085, 8.411843, 8.639058, 8.453894, 8.173026, 
    7.998325,
  4.415639, 4.610238, 5.069729, 6.286215, 7.291309, 7.820016, 7.995822, 
    7.801025, 7.621345, 7.998217, 8.593103, 8.709345, 8.488501, 8.264803, 
    8.27588,
  4.516429, 4.741838, 5.139556, 6.507192, 7.54945, 7.989509, 8.167657, 
    8.054463, 7.926069, 8.244856, 8.647081, 8.671278, 8.493377, 8.366457, 
    8.490965,
  4.799869, 4.83926, 5.290655, 6.755543, 7.755351, 8.159489, 8.307885, 
    8.188595, 8.092487, 8.298169, 8.628609, 8.649222, 8.520951, 8.371423, 
    8.494102,
  5.000318, 5.064464, 5.698795, 7.09052, 8.009466, 8.386382, 8.574369, 
    8.462717, 8.337302, 8.48002, 8.694361, 8.734012, 8.583425, 8.348636, 
    8.368415,
  5.286648, 5.612872, 6.22387, 7.377277, 8.237932, 8.649895, 8.885566, 
    8.704051, 8.582907, 8.65948, 8.786345, 8.775846, 8.674512, 8.367174, 
    8.170189,
  4.840213, 4.300356, 4.470174, 5.010213, 6.130949, 7.16425, 7.803757, 
    7.943141, 7.731341, 7.513824, 7.473201, 7.821309, 7.998015, 8.044427, 
    8.121047,
  4.536325, 4.316646, 4.615436, 5.307121, 6.550829, 7.427148, 8.038128, 
    7.950766, 7.72303, 7.661046, 7.744743, 7.975108, 8.152325, 7.896633, 
    8.064974,
  4.366117, 4.477331, 4.959516, 5.86488, 7.062694, 7.144786, 8.019784, 
    8.100835, 7.927036, 7.723871, 7.854432, 7.977167, 8.097128, 8.22373, 
    8.306803,
  4.320742, 4.757911, 5.454323, 6.567672, 7.661934, 8.075935, 7.412395, 
    7.921312, 7.806339, 7.765512, 7.812449, 7.850685, 7.883544, 7.941721, 
    8.106407,
  4.461497, 5.224181, 6.295795, 7.371392, 8.135021, 8.382433, 8.267281, 
    6.780396, 6.554841, 7.780149, 7.88309, 7.80594, 7.836408, 7.840151, 
    7.954325,
  4.921549, 6.164867, 7.183359, 8.104373, 8.433802, 8.579097, 8.512277, 
    8.345788, 8.270303, 8.194683, 8.074393, 7.963049, 7.975875, 7.963416, 
    7.973928,
  5.731123, 7.087089, 7.982433, 8.534364, 8.623423, 8.723964, 8.72693, 
    8.669856, 8.53051, 8.35676, 8.292459, 8.188532, 8.15852, 8.184744, 8.14153,
  6.600141, 7.836315, 8.502016, 8.743834, 8.690906, 8.819137, 8.780136, 
    8.665447, 8.509717, 8.40809, 8.364996, 8.27473, 8.247774, 8.232541, 
    8.214351,
  7.262403, 8.379124, 8.869057, 8.847259, 8.704367, 8.793108, 8.729146, 
    8.637899, 8.500708, 8.44037, 8.408876, 8.383067, 8.392705, 8.329165, 
    8.219748,
  7.66162, 8.720184, 9.046493, 8.751584, 8.574229, 8.622604, 8.585787, 
    8.501839, 8.45774, 8.472602, 8.46655, 8.383736, 8.274733, 8.272435, 
    8.245391,
  5.187421, 4.486176, 5.386443, 6.912899, 8.057065, 8.411882, 8.326539, 
    8.216886, 8.169356, 8.066003, 8.069956, 7.874512, 7.65637, 7.408896, 
    7.542846,
  4.760683, 5.148792, 6.766276, 7.977601, 8.456261, 8.260503, 8.183236, 
    8.107355, 8.069856, 8.176769, 8.235369, 8.061718, 7.762105, 7.236134, 
    7.452247,
  5.11916, 6.455931, 7.842295, 8.46281, 8.381864, 7.395889, 7.895999, 
    8.07913, 8.007897, 8.027563, 8.107359, 8.1589, 7.868862, 7.665108, 
    7.707361,
  6.005344, 7.62322, 8.368285, 8.460715, 8.285329, 8.178974, 7.221774, 
    7.627183, 7.680525, 7.937523, 7.956721, 8.020147, 7.930284, 7.747699, 
    7.712173,
  7.109574, 8.302891, 8.409761, 8.331448, 8.313665, 8.356694, 8.140606, 
    6.557811, 6.32397, 7.729505, 7.946994, 7.898687, 7.912974, 7.773067, 
    7.665342,
  7.993965, 8.493989, 8.306816, 8.318116, 8.430954, 8.415507, 8.193215, 
    7.980344, 7.817626, 7.898694, 7.973284, 7.917518, 7.82649, 7.804097, 
    7.639951,
  8.189279, 8.468148, 8.305448, 8.478057, 8.586145, 8.456054, 8.241933, 
    8.131537, 8.004913, 7.925828, 8.104259, 8.060206, 7.815812, 7.776046, 
    7.64881,
  8.112718, 8.393941, 8.455173, 8.643102, 8.683296, 8.447026, 8.256893, 
    8.134052, 8.036176, 7.935485, 8.205399, 8.144233, 7.790879, 7.714501, 
    7.686869,
  8.028339, 8.457975, 8.688695, 8.861382, 8.856575, 8.525221, 8.334869, 
    8.251073, 8.226544, 8.127745, 8.299371, 8.31371, 7.995513, 7.766344, 
    7.713444,
  7.900581, 8.550908, 8.837299, 9.004695, 9.023638, 8.641643, 8.398547, 
    8.349608, 8.337667, 8.36051, 8.425892, 8.539454, 8.008303, 7.82011, 
    7.723857,
  5.860821, 6.820814, 7.801905, 7.986106, 7.946323, 7.799107, 7.664507, 
    7.691016, 7.77796, 7.774197, 7.815989, 7.75293, 7.358444, 6.810498, 
    6.685718,
  6.746802, 7.84404, 8.265152, 8.084988, 7.862044, 7.619413, 7.693607, 
    7.549892, 7.561364, 7.728022, 7.897138, 7.821138, 7.403366, 6.573681, 
    6.739357,
  7.642652, 8.455559, 8.340892, 8.004463, 7.768015, 6.860323, 7.569952, 
    7.573524, 7.451818, 7.576588, 7.800532, 7.889598, 7.456985, 7.043154, 
    7.088934,
  8.246367, 8.72449, 8.289422, 7.870897, 7.765004, 7.706987, 6.784382, 
    7.455029, 7.352024, 7.44085, 7.712764, 7.808574, 7.474184, 7.174065, 
    7.255661,
  8.690756, 8.761854, 8.125179, 7.728565, 7.66079, 7.782507, 7.865145, 
    6.159949, 5.8902, 7.435772, 7.714986, 7.681857, 7.487887, 7.20311, 
    7.282047,
  8.919509, 8.720912, 7.940634, 7.606867, 7.500807, 7.665452, 7.880173, 
    7.670488, 7.248968, 7.580786, 7.64767, 7.660425, 7.498013, 7.271107, 
    7.270211,
  8.965483, 8.627881, 7.833326, 7.486317, 7.435302, 7.621243, 7.753687, 
    7.84369, 7.641134, 7.530204, 7.623429, 7.662212, 7.518305, 7.307312, 
    7.277203,
  8.94434, 8.517235, 7.759647, 7.429811, 7.389055, 7.618199, 7.720232, 
    7.719755, 7.550667, 7.513198, 7.715295, 7.717186, 7.540168, 7.301377, 
    7.248275,
  8.875854, 8.487089, 7.784737, 7.496454, 7.468418, 7.590126, 7.623024, 
    7.622814, 7.578849, 7.67045, 7.85595, 7.726437, 7.523938, 7.271837, 
    7.184548,
  8.896629, 8.565101, 7.82203, 7.520863, 7.590753, 7.747289, 7.789733, 
    7.760098, 7.793835, 7.915633, 7.952894, 7.731022, 7.510241, 7.291475, 
    7.086231,
  9.690311, 9.627851, 8.788217, 7.405969, 6.789168, 6.774873, 6.984068, 
    6.966542, 6.847202, 6.995724, 7.266374, 7.507817, 7.078789, 6.701924, 
    10.59906,
  10.08815, 9.473365, 7.643043, 6.759028, 6.551363, 6.78352, 7.304765, 
    7.313622, 7.102247, 7.116429, 7.285014, 7.458132, 6.879104, 7.275959, 
    11.45341,
  10.03333, 8.451392, 6.823979, 6.461691, 6.683118, 6.215815, 7.644713, 
    7.460279, 7.147384, 7.256913, 7.369275, 7.345324, 6.887357, 8.935247, 
    12.30789,
  9.229448, 7.335937, 6.462806, 6.49784, 6.961573, 7.175309, 6.265441, 
    7.334574, 7.049489, 7.242134, 7.404908, 7.244576, 7.338381, 10.18449, 
    12.73658,
  8.156559, 6.731424, 6.426486, 6.618399, 6.970211, 7.398899, 7.194723, 
    5.672458, 5.452878, 7.227417, 7.420088, 7.332409, 8.518406, 11.04154, 
    13.08719,
  7.318725, 6.539383, 6.475072, 6.75571, 6.995002, 7.142433, 7.141909, 
    6.772615, 6.816204, 7.343669, 7.450216, 7.900047, 9.546025, 11.61782, 
    13.24144,
  6.857347, 6.520542, 6.587409, 6.908654, 7.081798, 7.167446, 7.133593, 
    7.180543, 7.269398, 7.507535, 7.838664, 8.853652, 10.28042, 11.94753, 
    13.08723,
  6.671527, 6.567016, 6.734117, 7.037998, 7.157868, 7.306572, 7.307117, 
    7.348511, 7.52811, 7.887859, 8.434896, 9.293634, 10.50647, 11.7678, 
    12.60269,
  6.71508, 6.755166, 6.930843, 7.123724, 7.219146, 7.331962, 7.41123, 
    7.57836, 7.79119, 8.088375, 8.549792, 9.226676, 10.12747, 11.00424, 
    11.73799,
  6.916975, 7.075245, 7.248939, 7.330939, 7.398808, 7.47144, 7.547958, 
    7.661247, 7.8203, 8.047292, 8.4374, 8.977753, 9.689393, 10.51325, 11.21692,
  16.3471, 15.06024, 13.78762, 12.0584, 10.26986, 8.753033, 7.565101, 
    6.761458, 6.124114, 6.085975, 6.701086, 6.769813, 6.823546, 6.550947, 
    9.766303,
  16.21801, 14.48748, 12.44452, 10.25566, 8.407814, 7.338682, 6.718338, 
    6.42551, 6.346431, 6.195708, 6.456947, 6.498941, 6.719894, 6.640139, 
    11.02519,
  15.23531, 13.14459, 10.3314, 8.231943, 6.93877, 5.629883, 7.102087, 
    6.729986, 6.482436, 6.337376, 6.455581, 6.468637, 6.615551, 7.759399, 
    12.62755,
  13.50648, 10.60458, 7.828278, 6.499754, 6.270201, 6.217205, 5.718689, 
    6.805924, 6.474819, 6.463946, 6.478984, 6.510171, 6.921309, 9.758589, 
    13.44564,
  10.3533, 7.238367, 6.083738, 5.889291, 6.12388, 6.668803, 6.614043, 
    5.274077, 4.989779, 6.317566, 6.524652, 6.741141, 8.095767, 11.96631, 
    14.23464,
  6.722586, 5.769119, 5.710915, 5.971829, 6.408427, 6.635896, 6.651865, 
    6.441097, 6.333313, 6.298043, 6.612573, 7.643045, 10.59225, 13.74839, 
    14.33309,
  5.843826, 5.766736, 5.973767, 6.318439, 6.591688, 6.565687, 6.372969, 
    6.289342, 6.377488, 6.435288, 7.454901, 9.827301, 12.95717, 14.26962, 
    13.38685,
  6.008677, 6.151432, 6.466839, 6.68604, 6.660369, 6.554801, 6.564278, 
    6.695314, 7.064935, 7.832421, 9.770194, 12.32049, 13.97095, 13.82395, 
    12.5021,
  6.323866, 6.583755, 6.85641, 6.996146, 7.07283, 7.1722, 7.368559, 7.622409, 
    8.394282, 9.993939, 12.18148, 13.63367, 13.92867, 12.99088, 12.47788,
  6.683291, 6.895072, 7.117823, 7.246051, 7.328657, 7.549247, 7.937912, 
    8.721953, 10.2997, 11.96304, 13.25282, 13.71789, 13.30824, 12.8409, 
    12.66199,
  19.67376, 17.94203, 15.94765, 13.95473, 12.9315, 12.3501, 11.93429, 
    11.40181, 9.828848, 7.830849, 6.482734, 5.858842, 5.623236, 5.470647, 
    7.10904,
  19.0626, 17.41881, 15.49089, 13.99167, 12.96844, 12.35885, 11.57162, 
    10.08229, 7.970351, 6.47765, 5.485056, 5.169205, 5.239451, 5.389895, 
    9.037321,
  18.51624, 17.03753, 15.30003, 14.08204, 12.98225, 10.80824, 10.51695, 
    8.697764, 6.879096, 5.756926, 5.142122, 5.155941, 5.396092, 7.309165, 
    12.20464,
  17.48298, 16.29496, 14.84795, 13.22661, 11.85544, 10.25056, 7.935041, 
    7.20533, 5.914505, 5.403914, 5.076687, 5.216016, 6.150467, 10.76237, 
    13.51633,
  15.38282, 14.03724, 12.45589, 11.03079, 9.798973, 8.783461, 7.4255, 
    5.088201, 4.296246, 5.135916, 5.171457, 5.625691, 8.724238, 12.73641, 
    14.09971,
  10.85079, 9.815653, 9.051292, 8.31769, 7.669269, 7.033227, 6.666437, 
    5.844014, 5.436131, 5.339143, 5.252937, 7.208296, 11.50259, 13.61258, 
    14.19459,
  6.903677, 6.718506, 6.550668, 6.458795, 6.519726, 6.226235, 6.224424, 
    5.997543, 5.548295, 5.125531, 6.005429, 10.0106, 13.04228, 13.79914, 
    14.02367,
  6.001774, 5.912986, 5.926667, 6.092052, 6.134049, 6.007184, 6.072279, 
    5.702537, 5.375964, 5.418921, 7.946751, 12.30085, 13.7256, 13.90802, 
    14.46614,
  6.249598, 6.400612, 6.426848, 6.359578, 6.366004, 6.2007, 6.120042, 
    5.617725, 5.578349, 6.941382, 11.05913, 13.41623, 13.9405, 14.22771, 
    15.04761,
  6.955944, 7.014346, 6.905422, 6.601909, 6.496072, 6.31837, 6.142055, 
    5.851148, 6.919814, 10.0017, 13.01444, 13.82206, 13.98935, 14.43605, 
    15.03565,
  19.26182, 18.93426, 19.4641, 19.76961, 19.36402, 17.78765, 15.24284, 
    12.69557, 11.99851, 11.69223, 9.601343, 6.778757, 5.041954, 4.59479, 
    4.633518,
  19.31655, 19.06728, 19.30123, 18.85481, 17.94381, 16.27025, 13.74049, 
    11.90102, 11.12694, 9.814721, 6.96571, 4.72896, 4.4303, 4.640965, 5.41003,
  19.46118, 19.24606, 18.83951, 17.76393, 16.65394, 13.49831, 12.41344, 
    10.81437, 9.792034, 7.560151, 5.158773, 4.530408, 5.565047, 7.601006, 
    8.933578,
  19.27611, 19.00786, 18.08805, 16.7636, 15.83613, 13.24251, 10.51073, 
    9.888384, 8.350696, 5.98931, 4.585978, 4.990383, 7.526949, 10.94497, 
    11.9513,
  18.77223, 18.38648, 17.35849, 16.08998, 14.75678, 12.70526, 10.4642, 
    7.93685, 5.589288, 4.654745, 4.522938, 7.260203, 11.66336, 13.62577, 
    14.07369,
  17.94218, 17.70165, 16.7116, 15.41806, 13.67584, 11.7684, 9.610641, 
    7.324113, 5.321502, 4.695965, 5.537889, 10.22253, 13.62951, 14.9925, 
    15.27006,
  16.70226, 16.63275, 15.67432, 14.25905, 12.62969, 10.56965, 8.151523, 
    6.131187, 4.83473, 4.52421, 7.835752, 12.77118, 14.538, 15.61608, 15.64629,
  14.57226, 14.59165, 13.80902, 12.58368, 11.27134, 9.172369, 6.802425, 
    5.281684, 4.47752, 4.943357, 9.430799, 13.79734, 15.01163, 15.49465, 
    15.68645,
  12.25096, 12.11882, 11.51472, 10.87227, 10.04085, 8.180675, 6.266888, 
    4.966286, 4.439005, 5.7795, 11.18357, 13.86661, 14.65371, 15.15852, 
    15.96287,
  10.44864, 10.26085, 9.973392, 9.681552, 9.011911, 7.475598, 5.874601, 
    4.681273, 4.62166, 7.904321, 12.55504, 13.75981, 14.50307, 15.39269, 
    16.02746,
  21.36833, 21.55908, 21.10266, 21.22701, 21.31153, 20.77676, 20.96805, 
    20.87685, 19.40141, 16.47364, 14.17884, 11.44058, 8.72119, 6.216761, 
    4.944338,
  21.62936, 21.80722, 21.42285, 21.59609, 20.90082, 20.22079, 20.6399, 
    19.99472, 17.98671, 15.53452, 13.00159, 9.946436, 7.459599, 6.104974, 
    6.082425,
  21.60697, 21.71659, 21.64502, 21.30637, 20.25898, 17.9438, 19.53538, 
    18.29402, 16.21269, 13.81692, 10.90288, 8.328595, 7.464386, 8.373396, 
    8.902364,
  21.48176, 21.63937, 21.26167, 20.45132, 19.83719, 18.15591, 16.14648, 
    15.86414, 14.02685, 11.74967, 8.879194, 7.246374, 8.233356, 9.73017, 
    10.51441,
  21.0225, 20.87559, 20.06509, 18.95659, 18.2646, 17.40461, 15.99293, 
    12.32926, 10.6792, 9.481541, 7.041527, 7.807046, 10.55307, 12.24546, 
    12.47128,
  20.2236, 19.49544, 18.08273, 17.0484, 16.27876, 15.44676, 13.96165, 
    11.78394, 9.874113, 7.115321, 7.100728, 10.63042, 12.85807, 13.51437, 
    13.27156,
  19.32998, 18.20495, 16.83663, 15.95782, 15.11821, 13.16832, 11.13733, 
    9.270543, 7.264003, 7.090916, 11.00757, 13.14882, 13.81493, 13.65757, 
    13.05633,
  18.61566, 17.29094, 16.02581, 14.49806, 12.18961, 9.643648, 8.127743, 
    7.090981, 7.277334, 10.7561, 13.1527, 14.06124, 14.14501, 13.91939, 
    13.54319,
  17.90923, 16.46134, 14.64423, 11.61583, 9.360712, 7.892857, 7.196799, 
    7.309912, 9.64447, 12.22693, 13.62989, 14.18229, 14.52189, 14.42048, 
    14.29771,
  16.98476, 15.08662, 11.55215, 8.857434, 7.746617, 6.967992, 6.785424, 
    7.812837, 10.0416, 11.95362, 12.82195, 13.66848, 14.51854, 14.52449, 
    14.04587,
  10.60232, 9.613351, 10.49529, 13.02127, 14.56097, 14.17772, 14.60164, 
    17.48459, 22.65298, 24.85431, 22.42822, 18.04557, 14.0081, 11.07604, 
    8.790551,
  13.41321, 11.72858, 11.46929, 12.48134, 12.91626, 12.0361, 12.8981, 
    15.60626, 20.30369, 23.93988, 22.54744, 18.68799, 15.49832, 12.36621, 
    9.346265,
  15.29656, 13.42664, 12.6125, 12.30312, 11.80293, 10.28393, 12.17592, 
    14.61005, 18.3019, 22.48666, 22.19096, 19.24485, 16.24737, 13.68201, 
    10.7953,
  16.06697, 14.5007, 13.45725, 12.44057, 11.9323, 11.63995, 11.64388, 
    14.40511, 16.49379, 20.24187, 21.16523, 19.49817, 16.40097, 13.76184, 
    11.57974,
  16.51, 15.25278, 14.19453, 13.27885, 13.0038, 13.52505, 14.26254, 12.80904, 
    13.01418, 18.07826, 19.49026, 18.32522, 15.7378, 13.44252, 11.90989,
  16.44722, 15.58643, 14.81765, 14.32975, 14.2731, 15.01434, 16.17753, 
    16.96077, 16.79992, 17.18177, 16.84891, 15.76355, 14.36853, 13.1603, 
    12.24006,
  16.12878, 15.70009, 15.52895, 15.8229, 16.34905, 16.96921, 17.30075, 
    17.4189, 16.53915, 15.03998, 14.0997, 13.71774, 13.32949, 12.84499, 
    12.29521,
  15.58127, 15.58019, 15.67286, 16.01758, 16.22016, 16.1861, 15.52996, 
    14.2437, 13.08812, 12.4812, 12.45228, 12.52144, 12.41675, 12.13843, 
    11.97792,
  13.82351, 13.8377, 13.79928, 13.61014, 12.99888, 11.89234, 10.81405, 
    10.60536, 10.99495, 11.43031, 11.92664, 12.26041, 12.35973, 11.76893, 
    11.76746,
  11.77672, 11.23792, 10.73689, 10.17915, 9.590722, 9.371308, 9.804784, 
    10.47557, 11.04814, 11.60274, 12.37306, 12.74449, 12.14711, 10.78261, 
    11.3475,
  11.807, 11.34931, 11.48521, 13.1815, 13.98035, 13.92812, 13.33383, 
    13.60932, 14.97188, 19.8112, 21.55492, 15.92748, 11.06479, 10.09808, 
    12.16935,
  11.32667, 11.84389, 13.14455, 13.87816, 14.08796, 14.23392, 14.30947, 
    14.67435, 15.67397, 20.0022, 21.15957, 15.97901, 11.236, 9.62829, 11.72643,
  11.76884, 12.89466, 13.89432, 13.84344, 13.84876, 12.93315, 14.39311, 
    15.40287, 16.83738, 20.25142, 20.90045, 16.02292, 11.55348, 10.49527, 
    11.97857,
  11.78387, 12.49417, 13.21926, 13.20137, 13.50596, 13.53436, 12.5115, 
    15.13627, 17.41107, 20.54564, 20.90732, 16.21175, 12.01678, 11.41331, 
    12.3303,
  11.13569, 11.20617, 11.56017, 12.00801, 12.62772, 13.12382, 13.0421, 
    11.98787, 14.23464, 20.75189, 21.27229, 16.91633, 12.85226, 12.44548, 
    13.04046,
  10.88325, 10.5395, 10.32894, 10.92913, 11.60288, 11.97711, 12.95087, 
    14.17354, 16.40582, 20.56267, 21.47969, 17.95969, 14.3812, 14.05814, 
    14.23742,
  10.92562, 10.89436, 10.77371, 11.2676, 12.25658, 13.04282, 13.67039, 
    15.17513, 16.98393, 19.84463, 20.77301, 18.23179, 15.96462, 15.68823, 
    15.44909,
  12.6791, 12.93387, 13.20703, 13.64497, 14.28144, 15.05171, 15.65352, 
    16.34838, 17.30626, 18.82547, 19.25806, 17.88861, 16.80474, 16.39631, 
    15.8699,
  14.49448, 14.56691, 14.77209, 14.97404, 15.12382, 15.3479, 15.75663, 
    16.17137, 16.43571, 16.80991, 17.01358, 16.69744, 16.10858, 15.54816, 
    14.75307,
  12.15579, 11.41619, 11.16608, 11.41324, 11.93334, 12.59106, 13.15867, 
    13.63252, 13.9555, 14.27591, 14.51308, 14.49258, 14.19974, 13.49418, 
    12.78052,
  11.99556, 12.03716, 12.35233, 12.67543, 13.47875, 14.33587, 15.03773, 
    14.90218, 13.98332, 12.44932, 16.02434, 17.73386, 15.98067, 14.8557, 
    15.01384,
  11.84417, 12.16998, 12.75744, 12.81586, 12.77899, 13.36189, 14.38881, 
    14.69742, 14.05022, 12.65693, 15.30352, 17.66359, 15.83947, 14.08438, 
    14.93081,
  11.65084, 12.3427, 13.47516, 13.62175, 13.02233, 11.59583, 13.43787, 
    14.32311, 14.0762, 12.80813, 14.4559, 17.15479, 15.71728, 14.62119, 
    15.62466,
  11.73173, 12.80401, 14.11707, 14.23934, 13.69764, 12.44238, 11.57582, 
    13.35089, 13.55293, 12.73749, 13.7985, 16.4334, 15.65337, 14.60208, 
    15.99963,
  12.2557, 13.43752, 14.40717, 14.55014, 13.95815, 12.95793, 12.12216, 
    10.69268, 10.76488, 12.25714, 13.21992, 15.61731, 15.65309, 14.47154, 
    15.92981,
  12.82645, 13.69598, 13.87809, 13.64664, 13.31671, 12.67759, 12.13158, 
    11.78308, 12.02104, 12.1691, 12.65296, 15.07366, 15.57766, 14.31414, 
    15.34751,
  12.83393, 13.39493, 13.13243, 12.49992, 12.64201, 12.24494, 11.68667, 
    11.85698, 12.27621, 12.11049, 12.55915, 15.01396, 15.368, 13.98889, 
    14.41578,
  12.20497, 12.92762, 12.81416, 12.6425, 12.67751, 12.33972, 11.75125, 
    11.86695, 12.25575, 12.5291, 13.16961, 15.1733, 15.20248, 13.64459, 
    13.54245,
  11.18269, 12.13547, 12.66791, 12.80004, 12.8565, 12.74874, 12.39919, 
    12.5293, 12.93256, 13.27811, 13.90713, 15.28955, 15.33501, 13.72707, 
    13.39338,
  9.937451, 11.02024, 11.86806, 12.55162, 12.90219, 12.99515, 12.98689, 
    13.16091, 13.50787, 13.83297, 14.51673, 15.68828, 15.67422, 14.28809, 
    13.79971,
  11.21246, 10.6146, 10.59667, 10.75886, 11.06289, 11.24911, 11.79701, 
    12.87452, 13.94275, 13.76719, 13.94336, 15.49156, 17.16528, 18.51172, 
    18.90356,
  10.5389, 10.31157, 10.37933, 10.74612, 11.14669, 11.30837, 11.6899, 
    12.5708, 13.62999, 13.76893, 14.20547, 16.22549, 17.88403, 18.29, 18.85392,
  10.2711, 10.62045, 10.94503, 11.26248, 11.49301, 10.72357, 11.58046, 
    12.44558, 13.49935, 13.59099, 14.41263, 16.99029, 18.48966, 19.32702, 
    19.17625,
  10.94721, 11.52506, 11.72556, 11.79966, 11.92344, 11.95899, 11.04015, 
    11.97235, 13.14899, 13.36188, 14.94776, 17.79476, 18.89507, 19.20568, 
    18.45369,
  11.64366, 11.84669, 11.7816, 11.77644, 11.91971, 12.23801, 12.13867, 
    10.46144, 10.48949, 12.7183, 15.51953, 18.3379, 19.08136, 18.4357, 
    17.27173,
  11.8001, 11.86082, 11.5613, 11.38048, 11.56541, 12.11496, 12.42561, 
    12.09137, 12.14976, 13.01212, 16.40826, 18.66677, 18.7035, 17.34603, 
    16.04172,
  11.88344, 11.95329, 11.71647, 11.24336, 11.30434, 12.01838, 12.43699, 
    12.30294, 12.79077, 13.5601, 17.02304, 18.47479, 17.87515, 16.1334, 
    15.70541,
  12.03939, 12.09902, 11.87649, 11.31481, 11.26048, 12.17917, 12.51883, 
    12.29179, 12.9243, 14.28074, 17.04457, 17.92183, 16.91771, 15.36465, 
    16.10884,
  12.10819, 12.19943, 11.98784, 11.67089, 11.832, 12.508, 12.63636, 12.66339, 
    13.3964, 14.59056, 16.56018, 17.12873, 15.96555, 15.49251, 16.48336,
  12.18184, 12.39307, 12.4209, 12.35805, 12.5176, 12.82599, 12.82608, 
    13.07538, 13.51807, 14.45099, 15.77019, 16.34839, 15.6198, 15.89921, 
    16.47443,
  15.72064, 14.92427, 14.18628, 13.3621, 12.55346, 11.88091, 11.32336, 
    11.01929, 10.91088, 10.64288, 10.83142, 11.46134, 12.04494, 12.32011, 
    12.79818,
  13.88597, 12.86493, 12.10199, 11.51379, 11.10668, 10.79556, 10.72734, 
    10.6293, 10.5924, 10.79843, 11.11175, 11.65282, 12.38844, 12.15277, 
    12.59575,
  10.99436, 10.4743, 10.30104, 10.32067, 10.38976, 9.624619, 10.32078, 
    10.72381, 10.69684, 10.7872, 11.03343, 11.59106, 12.40977, 12.9651, 
    13.34175,
  9.62243, 10.0967, 10.6377, 11.04142, 11.22135, 11.11909, 10.08378, 
    10.72349, 10.78762, 10.98598, 11.10882, 11.72407, 12.66452, 13.28555, 
    14.06817,
  10.91499, 11.77385, 12.13992, 12.14657, 12.04673, 11.7965, 11.42742, 
    9.343152, 9.064783, 10.86881, 11.42206, 12.38063, 13.23185, 13.80178, 
    14.98894,
  12.27589, 12.44131, 12.32902, 12.06124, 11.87528, 11.74208, 11.56163, 
    11.26019, 10.96648, 10.99144, 11.62152, 13.08074, 13.85835, 14.43931, 
    16.06561,
  12.54472, 12.40124, 11.74698, 11.42457, 11.39199, 11.38233, 11.28371, 
    11.36454, 11.09001, 10.96306, 12.83181, 14.24825, 14.75746, 15.30369, 
    16.07537,
  12.60199, 11.8414, 11.19605, 11.16054, 11.24298, 11.27518, 11.13378, 
    11.0387, 10.8734, 12.23973, 14.52816, 15.32626, 15.62823, 15.4398, 
    14.66969,
  12.47889, 11.62868, 11.08468, 11.07065, 11.17034, 11.1512, 10.98247, 
    10.9621, 11.85095, 14.53551, 15.83791, 16.10578, 15.62221, 14.61777, 
    12.63104,
  12.51025, 11.92079, 11.45342, 11.12125, 11.02144, 10.99542, 11.02924, 
    11.88814, 14.44163, 16.21304, 16.64516, 16.14786, 14.87255, 13.32136, 
    10.72783,
  22.91823, 22.13336, 21.69902, 20.98606, 20.16925, 19.54135, 18.86466, 
    18.17251, 17.13464, 15.7155, 13.46377, 10.62617, 9.274355, 9.138274, 
    10.66851,
  22.26204, 21.48071, 20.75546, 19.97268, 18.85309, 17.91436, 17.00237, 
    15.55546, 14.01365, 12.31976, 9.707758, 8.905135, 8.890784, 9.213311, 
    11.90497,
  20.26182, 19.46343, 18.49427, 17.80602, 16.91588, 14.41829, 14.86481, 
    13.68706, 12.03333, 10.20614, 8.88474, 8.913045, 9.110258, 10.54972, 
    13.87721,
  15.99664, 15.53718, 14.80874, 14.28215, 14.02304, 13.34212, 11.53012, 
    11.68579, 10.84424, 9.891729, 9.412979, 9.347104, 9.336912, 11.45671, 
    14.17795,
  11.36343, 12.07454, 12.33412, 12.24178, 12.2392, 12.29621, 11.69918, 
    9.398839, 8.608295, 9.757036, 9.706703, 9.526368, 9.613876, 12.01585, 
    12.70744,
  10.14138, 11.18936, 11.4852, 11.50414, 11.39499, 11.4225, 11.43629, 
    11.14907, 10.95372, 10.88435, 10.44158, 9.799985, 9.957029, 12.01855, 
    10.72952,
  11.35116, 11.61997, 11.57512, 11.3946, 11.27054, 11.20848, 11.25384, 
    11.353, 11.38943, 11.12801, 10.68894, 9.932803, 10.48409, 11.65676, 
    9.450728,
  11.70283, 11.89865, 11.84379, 11.64588, 11.46605, 11.31484, 11.24098, 
    11.20572, 11.1691, 11.10665, 10.73545, 10.00035, 10.87334, 11.0444, 
    8.435983,
  11.94182, 12.30309, 12.34663, 12.09841, 11.79437, 11.5247, 11.27045, 
    11.23537, 11.17944, 11.04535, 10.57913, 10.1468, 11.32139, 10.48592, 
    7.640438,
  12.08936, 12.95236, 12.98174, 12.40578, 11.63656, 11.22351, 11.06472, 
    10.98021, 10.93114, 10.82248, 10.43354, 10.53827, 11.67131, 9.760134, 
    6.952003,
  18.28478, 19.1622, 22.23342, 22.95694, 22.28155, 21.46605, 20.60613, 
    18.54587, 17.23651, 16.8019, 16.57766, 12.69796, 7.701912, 8.110134, 
    8.818724,
  19.27293, 20.07767, 22.19359, 22.56062, 21.80018, 20.62646, 19.38929, 
    17.87825, 17.27013, 16.85274, 14.24173, 8.814995, 7.202436, 7.908612, 
    8.190592,
  18.82613, 20.97065, 22.21622, 22.05802, 20.59426, 18.01949, 18.60634, 
    17.90016, 17.30425, 15.28845, 10.93366, 7.560099, 7.592659, 8.363091, 
    7.816685,
  17.58626, 20.90684, 22.05925, 21.48814, 19.88997, 18.37729, 16.54371, 
    17.38876, 16.35276, 13.45216, 9.17537, 7.85199, 7.981781, 8.155996, 
    7.322534,
  15.84387, 19.94069, 21.49883, 20.94957, 19.37623, 18.80504, 17.63128, 
    14.7002, 12.8871, 12.10093, 9.038307, 8.314142, 8.367245, 7.865679, 
    6.84489,
  12.76384, 18.14288, 20.10116, 20.01921, 18.64189, 18.32953, 17.90895, 
    16.45889, 14.12193, 11.52527, 9.264902, 8.574466, 8.468791, 7.479535, 
    6.688687,
  9.772075, 15.43995, 17.65347, 18.07458, 17.19048, 16.96224, 16.57589, 
    15.61316, 13.45781, 10.8963, 9.330712, 8.684098, 8.175124, 6.784187, 
    6.299907,
  9.673799, 12.64054, 15.16277, 15.91927, 15.57305, 15.52758, 15.00223, 
    13.63977, 11.71067, 10.2486, 9.386643, 8.825377, 7.955536, 6.576559, 
    6.156943,
  9.892729, 10.5392, 13.11048, 14.191, 14.37715, 14.36819, 13.86876, 
    12.67634, 11.1375, 10.14537, 9.650212, 8.991515, 7.857704, 6.502102, 
    5.869038,
  9.934582, 9.924302, 11.65575, 12.90469, 13.39858, 13.52527, 13.11583, 
    12.05358, 10.93358, 10.30363, 9.906206, 9.143471, 7.621955, 6.208087, 
    5.437527,
  9.727895, 13.09125, 17.76545, 18.75033, 18.32919, 17.93672, 18.53299, 
    20.06275, 19.61601, 19.31802, 19.04726, 16.91729, 11.62171, 8.405669, 
    7.964124,
  10.1019, 13.06528, 17.11996, 18.38532, 18.73733, 18.46778, 19.13805, 
    19.27388, 18.9535, 18.58344, 16.3181, 11.33339, 7.980973, 7.478792, 
    7.863215,
  10.6245, 12.74862, 16.56855, 17.38712, 18.17306, 16.77919, 18.17388, 
    18.1062, 17.55419, 15.12765, 10.62517, 7.880718, 7.660736, 7.681979, 
    7.601299,
  11.19497, 12.16237, 16.30298, 16.41138, 17.33136, 17.00209, 15.62738, 
    16.60513, 13.75454, 10.36318, 8.064266, 7.51787, 7.416947, 7.080672, 
    6.856368,
  11.37378, 11.43658, 16.00285, 15.89025, 16.31418, 16.63543, 14.93098, 
    11.56453, 8.938104, 8.662133, 7.761056, 7.366202, 6.578233, 6.009168, 
    5.801711,
  11.13001, 10.79015, 15.18043, 16.12312, 15.94888, 16.20093, 14.78661, 
    12.40543, 9.878896, 8.467919, 7.57033, 6.733121, 5.959327, 5.68583, 
    5.572539,
  10.56125, 10.41187, 14.08465, 16.35815, 16.32683, 16.30831, 14.52478, 
    12.5239, 10.2194, 8.528946, 7.291983, 6.158029, 5.622274, 5.417386, 
    5.400674,
  10.14592, 10.2161, 13.54046, 16.40168, 16.6374, 16.60678, 14.76582, 
    12.54477, 10.15139, 8.211206, 6.751862, 5.917784, 5.534167, 5.345983, 
    5.480686,
  10.13317, 9.81645, 13.22782, 16.24681, 16.85026, 16.76674, 14.95885, 
    12.6576, 9.965367, 7.926661, 6.67614, 5.947948, 5.552733, 5.466555, 
    6.248948,
  10.08065, 9.405106, 12.80984, 16.01954, 16.87155, 16.68439, 14.8262, 
    12.15225, 9.372896, 7.799098, 6.75658, 5.953224, 5.557716, 5.952252, 
    7.424871,
  27.71215, 26.02995, 24.96843, 22.78558, 20.11719, 19.59516, 18.90868, 
    18.02409, 18.19193, 17.50088, 15.12031, 11.94024, 9.859615, 8.721091, 
    8.153025,
  27.58954, 25.36319, 24.17687, 22.55916, 20.42942, 19.55928, 19.03212, 
    17.85349, 15.75621, 13.20411, 10.13237, 8.488246, 7.876667, 6.994647, 
    6.755535,
  22.89374, 21.72849, 21.27922, 20.73721, 19.68663, 17.25252, 18.1529, 
    16.33318, 13.00286, 9.630128, 7.953686, 7.417724, 7.011656, 6.506291, 
    6.107273,
  18.89437, 18.94609, 19.08333, 19.07148, 18.83025, 18.0429, 15.79732, 
    15.25192, 11.13865, 8.420966, 7.49516, 6.814208, 6.327603, 5.893529, 
    5.702439,
  16.92066, 17.34527, 17.4761, 17.59617, 17.53409, 17.53656, 16.17492, 
    12.20502, 8.144002, 7.960611, 7.124673, 6.252804, 5.71465, 5.429623, 
    5.861771,
  15.70636, 16.14163, 16.37816, 16.67579, 16.6939, 16.77507, 15.49278, 
    12.92101, 9.247994, 7.670941, 6.728334, 5.778232, 5.373778, 5.305434, 
    6.674505,
  15.16024, 15.57485, 15.88477, 16.1902, 16.26209, 16.24062, 14.58139, 
    12.03441, 9.033762, 7.281729, 6.266656, 5.438322, 5.006234, 5.916887, 
    8.423721,
  13.88625, 14.59625, 15.39083, 15.9917, 16.05655, 15.83872, 13.94963, 
    10.93288, 8.235812, 6.878309, 5.813262, 5.067345, 5.335649, 8.221654, 
    10.39866,
  12.99309, 13.69159, 14.35089, 15.19601, 15.573, 15.47778, 13.34346, 
    10.19133, 7.783617, 6.529865, 5.530193, 5.083833, 7.352757, 10.38766, 
    11.34077,
  12.34043, 12.84836, 13.21442, 13.83123, 14.68366, 14.89348, 12.69572, 
    9.536469, 7.525722, 6.117483, 5.151215, 6.015259, 9.502643, 10.97687, 
    10.9228,
  29.43139, 28.07939, 26.31157, 24.12653, 22.21614, 20.43427, 18.90639, 
    18.10553, 17.95577, 17.53517, 15.89514, 12.8458, 10.27365, 7.799921, 
    6.66742,
  25.32143, 22.91864, 19.74911, 16.74196, 15.13454, 14.6404, 15.02179, 
    15.70826, 16.4134, 16.45801, 14.7176, 11.92912, 9.268848, 6.645578, 
    6.048936,
  17.61731, 14.85534, 12.56812, 10.84376, 10.09709, 9.470624, 12.01735, 
    14.10229, 15.21768, 15.12697, 13.97844, 11.64924, 9.254333, 7.061949, 
    6.418223,
  12.00459, 10.00842, 8.675421, 8.025702, 7.940436, 8.811453, 9.313824, 
    12.03432, 14.02666, 14.40697, 13.55558, 11.60648, 9.232666, 7.395287, 
    6.868089,
  8.497072, 8.08089, 7.935196, 7.835486, 7.852678, 8.343977, 9.501844, 
    9.086398, 9.950169, 12.47278, 12.67931, 11.27617, 9.322632, 7.653017, 
    7.237579,
  8.664366, 8.541953, 8.24869, 7.968034, 7.852746, 8.106825, 9.063948, 
    10.27271, 11.43446, 11.71956, 11.41682, 10.54513, 9.192694, 7.608225, 
    7.685288,
  8.782378, 8.363455, 7.993177, 7.989675, 8.220836, 8.544554, 9.298658, 
    10.46013, 11.19728, 11.09055, 10.52752, 9.852201, 8.605197, 7.553944, 
    8.536304,
  8.526834, 8.268168, 8.343288, 8.894055, 9.503599, 9.781401, 10.14555, 
    10.80299, 11.01469, 10.60692, 9.879838, 9.002126, 7.999274, 8.303411, 
    9.597794,
  8.399248, 8.583541, 9.583527, 11.25378, 11.74132, 11.55894, 11.3718, 
    11.46645, 10.89613, 10.03524, 9.135501, 8.058693, 8.410859, 9.565495, 
    9.781285,
  8.49008, 9.925098, 11.72101, 13.00663, 13.23434, 12.54102, 11.86446, 
    11.40814, 10.32636, 9.305221, 8.116959, 8.088367, 9.277595, 9.237387, 
    9.163756,
  31.7895, 32.59174, 33.32624, 33.20451, 32.32535, 31.07198, 29.86718, 
    28.48605, 26.66275, 24.69075, 23.42371, 22.4725, 20.69626, 17.30694, 
    13.55501,
  28.32463, 28.28871, 28.34297, 27.57535, 26.26678, 24.81796, 23.87154, 
    22.13361, 20.51877, 19.32651, 18.82302, 18.95608, 18.71206, 15.89893, 
    13.1601,
  23.28852, 23.31083, 23.18922, 22.56167, 21.68128, 18.67338, 17.17989, 
    15.48474, 14.20338, 13.23121, 13.26395, 14.36813, 15.79922, 15.62846, 
    13.43715,
  19.66601, 19.14466, 17.95311, 16.28331, 14.47676, 12.90783, 10.10365, 
    9.760795, 9.208505, 9.178531, 9.720569, 10.90724, 12.52731, 13.46391, 
    12.59121,
  12.74722, 11.6897, 10.83298, 10.012, 9.250056, 8.742682, 8.150685, 
    6.362209, 5.990973, 7.36983, 7.84815, 9.118866, 10.88478, 11.98164, 
    11.71374,
  10.16632, 10.1071, 9.840775, 9.425303, 8.927055, 8.623515, 8.518847, 
    8.240629, 8.079941, 7.953475, 7.672533, 8.264424, 9.786052, 11.13556, 
    11.06563,
  10.35618, 9.924415, 9.19049, 8.674294, 8.667046, 8.878844, 9.036979, 
    9.132435, 9.107952, 8.859777, 8.502879, 8.421487, 9.242231, 10.30019, 
    10.41915,
  10.05322, 8.940406, 8.467208, 9.042999, 9.672853, 9.725388, 9.759286, 
    9.866219, 9.90424, 9.806798, 9.424562, 9.135739, 9.434347, 9.994549, 
    9.821022,
  8.626373, 8.295588, 9.50588, 10.36937, 9.989404, 9.431385, 9.4946, 
    9.924555, 10.14113, 9.903727, 9.532236, 9.315149, 9.613267, 9.770258, 
    9.605345,
  7.926195, 9.383184, 10.911, 10.35485, 9.005519, 8.713422, 9.375478, 
    10.23265, 10.31936, 9.804113, 9.416164, 9.40432, 9.692964, 9.632891, 
    9.572826,
  13.94739, 12.83355, 12.52167, 13.25688, 15.12249, 17.25922, 19.22919, 
    21.12579, 22.82963, 24.21607, 25.52568, 26.95086, 27.97671, 28.49316, 
    28.38187,
  14.30993, 13.6995, 13.52404, 14.28287, 16.04593, 18.03226, 20.13408, 
    21.67527, 22.74934, 23.35226, 23.70751, 24.08185, 24.88041, 24.62511, 
    25.3959,
  15.03226, 15.66989, 16.09849, 16.98782, 18.2946, 18.13312, 20.30464, 
    21.54948, 21.72102, 21.48462, 20.8636, 20.42664, 21.10746, 23.02717, 
    23.82151,
  13.91599, 14.95272, 16.20884, 17.43703, 18.53648, 19.47581, 18.06854, 
    18.96517, 19.15956, 18.72745, 17.93294, 17.16178, 16.89592, 17.94898, 
    19.55582,
  12.47046, 13.24336, 14.24653, 15.34795, 16.14956, 17.02766, 17.94184, 
    15.34994, 14.13391, 15.62176, 15.08848, 14.31343, 13.64758, 13.48923, 
    14.65267,
  10.86139, 11.17549, 11.60899, 11.97104, 12.28614, 12.83985, 13.74306, 
    14.09604, 13.53878, 12.75082, 11.94644, 11.10201, 10.51486, 10.61531, 
    11.52996,
  10.25116, 10.00733, 9.852929, 9.847524, 9.686238, 9.513801, 9.550582, 
    9.922639, 10.17038, 9.939618, 9.764295, 9.319119, 8.977516, 9.293625, 
    10.32793,
  9.947601, 9.793206, 9.319679, 8.943273, 8.490321, 8.0147, 7.726658, 
    7.571316, 7.6605, 7.88133, 8.397923, 8.754727, 8.865768, 9.181555, 
    10.13754,
  9.362836, 9.602841, 9.244495, 8.757053, 8.273976, 7.873767, 7.834569, 
    8.004966, 8.247281, 8.379782, 8.767745, 9.079998, 9.01283, 9.239394, 
    9.736491,
  9.106971, 9.485866, 9.037044, 8.439243, 7.95928, 7.930194, 8.266771, 
    8.543849, 8.880593, 9.275893, 9.444046, 9.384531, 9.152089, 9.317182, 
    9.494945,
  23.2146, 22.09434, 20.24925, 18.36459, 16.61683, 14.88393, 13.15587, 
    12.00872, 11.47844, 11.45907, 11.54824, 11.67101, 11.92235, 12.50953, 
    13.82041,
  19.4928, 18.99821, 17.70965, 16.22319, 14.61567, 12.89855, 11.83634, 
    11.57665, 11.67974, 12.03285, 12.2046, 12.47092, 13.1367, 13.30464, 
    14.10595,
  15.73872, 15.56707, 14.80389, 13.63439, 12.22103, 10.27542, 10.52276, 
    11.33136, 11.68535, 11.86799, 12.23791, 13.30557, 14.42211, 14.83656, 
    14.78756,
  11.77581, 11.87545, 11.50981, 10.80641, 10.05344, 9.480603, 8.718288, 
    10.1068, 10.59653, 11.23592, 12.7011, 14.62744, 15.49306, 15.58111, 
    15.23794,
  10.04403, 10.04214, 9.674687, 9.094797, 8.735958, 8.653517, 8.768576, 
    7.892628, 8.138078, 10.69028, 13.82394, 16.07693, 17.03105, 16.95031, 
    16.52609,
  9.75269, 9.515727, 8.952172, 8.547244, 8.444699, 8.423766, 8.39822, 
    8.622985, 9.290972, 10.43419, 13.7942, 16.31163, 17.64391, 18.36557, 
    17.93382,
  9.834674, 9.673909, 8.98936, 8.776731, 8.762244, 8.614841, 8.316049, 
    8.218482, 8.387332, 9.52444, 12.41097, 14.65265, 16.07278, 17.09476, 
    16.90297,
  9.8725, 9.470725, 8.898908, 8.763115, 8.718404, 8.565289, 8.325461, 
    8.144928, 8.143557, 8.843444, 10.2939, 11.88096, 13.23427, 13.76502, 
    13.16381,
  9.913646, 9.137703, 8.830211, 8.677243, 8.530439, 8.432868, 8.38382, 
    8.386885, 8.442211, 8.796964, 9.633841, 10.52178, 11.22676, 11.5003, 
    10.79904,
  9.636091, 8.9249, 8.842243, 8.633652, 8.523127, 8.534357, 8.516934, 
    8.517404, 8.59562, 8.833216, 9.263773, 9.831616, 10.07977, 10.32709, 
    9.909306,
  21.1559, 24.7736, 29.69938, 31.07525, 29.18625, 26.29606, 25.65495, 
    25.82683, 25.53125, 24.10063, 21.5918, 18.84611, 16.25638, 13.24305, 
    11.81811,
  20.18417, 22.76697, 26.16987, 29.40413, 29.7809, 27.86164, 26.25274, 
    24.97839, 23.78055, 22.2163, 19.79279, 17.30776, 14.70895, 11.87552, 
    11.78898,
  18.34176, 20.6528, 23.02939, 25.89602, 28.34627, 25.92608, 25.58922, 
    24.33154, 22.30568, 20.03021, 17.72445, 15.72819, 13.1918, 11.91123, 
    13.26129,
  16.49754, 18.09179, 19.93264, 21.82399, 23.81541, 24.5742, 21.5588, 
    20.98056, 19.6692, 17.76799, 16.01778, 14.13687, 11.81239, 12.04974, 
    14.50838,
  12.94325, 14.89525, 16.26555, 17.55196, 18.61516, 19.43698, 19.32992, 
    16.08875, 14.36977, 14.9439, 14.10922, 12.19419, 10.67167, 12.43073, 
    14.99113,
  9.597247, 11.01235, 12.32676, 13.40615, 14.30543, 14.97807, 15.20473, 
    14.70058, 13.55814, 12.61782, 12.13041, 10.55474, 10.27729, 12.5176, 
    14.7149,
  8.381977, 8.704504, 9.391, 10.26636, 11.06333, 11.53665, 11.75867, 11.7171, 
    11.27657, 11.06992, 10.94335, 9.751892, 10.14793, 12.27424, 13.94669,
  8.201084, 7.875609, 8.009806, 8.546621, 9.071587, 9.427311, 9.559116, 
    9.563473, 9.383512, 9.803818, 10.02539, 9.240803, 10.08755, 11.91499, 
    12.87656,
  8.267974, 7.956005, 8.170056, 8.229901, 8.32292, 8.400862, 8.481796, 
    8.501556, 8.427972, 8.92804, 9.217566, 8.908124, 10.16002, 11.90623, 
    12.42608,
  8.310481, 8.490709, 8.683267, 8.49879, 8.303118, 8.183683, 8.06119, 
    7.957604, 8.098245, 8.424688, 8.620414, 8.895761, 10.40521, 12.09119, 
    12.20263,
  16.83034, 18.43744, 23.11362, 27.7919, 29.07096, 27.2042, 24.1519, 
    21.97546, 22.45787, 24.73031, 26.95315, 27.54509, 25.67101, 23.21343, 
    21.75717,
  14.91395, 16.33952, 18.82784, 23.65392, 27.69119, 28.18721, 25.85145, 
    23.26067, 22.18937, 23.64755, 25.45602, 25.72484, 24.58524, 22.41631, 
    21.16735,
  13.06666, 14.42034, 16.49101, 19.65799, 24.37141, 25.3012, 26.696, 
    25.20879, 23.44082, 23.31995, 24.31577, 24.39528, 24.02381, 22.53099, 
    20.71341,
  12.04076, 13.14322, 14.97967, 17.71401, 21.40538, 24.74139, 24.77757, 
    25.84595, 24.89339, 24.06468, 24.10801, 24.18749, 23.66121, 21.35223, 
    19.56172,
  10.32086, 12.39533, 14.01294, 16.36156, 19.35313, 23.15071, 25.78043, 
    23.65209, 22.58425, 24.95625, 24.65563, 23.91639, 22.45605, 20.0766, 
    18.83885,
  8.500211, 10.87452, 13.22771, 15.26739, 17.75152, 20.95036, 24.14996, 
    26.39062, 27.06645, 26.28094, 24.73309, 23.23169, 21.204, 19.14876, 
    17.60772,
  7.662735, 8.77973, 11.74562, 14.57983, 16.56092, 18.97183, 21.95537, 
    24.27195, 26.03669, 25.6431, 24.1395, 22.09559, 19.77689, 17.61433, 
    15.48372,
  7.673236, 7.676712, 9.240571, 12.83762, 15.28891, 17.31958, 19.88855, 
    21.93242, 23.24041, 23.46213, 22.22193, 19.99086, 17.57451, 15.22433, 
    13.21827,
  7.961403, 7.683903, 7.904226, 10.18821, 13.25514, 15.26279, 17.29071, 
    18.8965, 19.92464, 20.04293, 18.92086, 16.93625, 14.77974, 12.96852, 
    12.24384,
  8.310343, 8.073271, 7.825768, 8.637675, 11.11888, 12.91632, 14.58244, 
    15.86064, 16.57696, 16.39767, 15.42351, 13.94139, 12.39681, 11.76711, 
    12.0237,
  18.62289, 21.91095, 25.27011, 27.86908, 29.42913, 29.20437, 28.03601, 
    26.17803, 23.69945, 24.07109, 25.49592, 27.32497, 27.81591, 26.97907, 
    24.8518,
  16.36034, 18.79462, 21.18595, 24.72588, 28.24817, 28.83505, 27.90445, 
    26.6754, 24.95261, 23.99022, 24.55713, 25.60169, 26.51849, 25.43647, 
    23.83576,
  13.10483, 15.42644, 17.6845, 19.863, 24.44555, 25.77116, 27.86825, 
    27.28372, 25.81892, 24.52375, 24.18757, 24.39591, 24.85769, 25.08725, 
    23.46918,
  9.68684, 11.3482, 13.97797, 16.01488, 18.65811, 22.75501, 24.9317, 
    27.54336, 27.05979, 25.76097, 24.62221, 24.29585, 24.54057, 24.76411, 
    23.40421,
  8.004177, 8.453995, 10.13162, 12.52921, 14.53873, 17.39674, 21.55138, 
    22.97515, 23.86168, 26.88761, 26.34531, 25.23063, 24.99246, 24.99438, 
    24.36623,
  7.974698, 7.628908, 7.81183, 9.531205, 11.40484, 13.31414, 16.26412, 
    19.37752, 22.62608, 25.82399, 26.84804, 26.41795, 26.00394, 25.70483, 
    25.32058,
  8.414824, 7.779929, 7.262484, 8.112849, 9.530959, 10.8326, 12.4532, 
    15.03089, 17.97255, 21.99444, 24.79708, 26.12247, 26.34661, 26.30126, 
    26.12789,
  8.922688, 8.123279, 7.406725, 7.852055, 8.836123, 9.729213, 10.69781, 
    12.21334, 14.47414, 17.54234, 21.30968, 24.27979, 25.56412, 26.12751, 
    26.04078,
  9.360091, 8.519067, 7.764781, 8.010258, 8.688075, 9.307614, 10.413, 
    11.67826, 13.17799, 15.51104, 18.52308, 21.51982, 23.87742, 24.92854, 
    24.68804,
  9.449499, 8.704049, 8.136049, 8.275272, 8.963667, 9.383555, 10.34703, 
    11.80948, 13.04758, 14.64988, 16.8512, 19.36144, 21.68274, 23.05633, 
    22.83835,
  24.65837, 26.5208, 26.21061, 26.21325, 26.53215, 26.85048, 26.20654, 
    25.42053, 25.16948, 25.29569, 25.19392, 25.35004, 25.50684, 24.8657, 
    24.27082,
  21.36302, 24.9164, 26.66667, 27.79173, 27.92317, 27.62631, 27.0458, 
    26.41814, 25.66319, 25.58675, 25.47361, 25.24315, 25.41333, 24.76037, 
    25.48739,
  17.3136, 21.68128, 24.85029, 27.32768, 28.60247, 26.29582, 27.62159, 
    27.33386, 26.79624, 26.27274, 25.93728, 25.46631, 25.36798, 25.95995, 
    27.03841,
  13.11659, 17.12792, 21.18848, 24.16665, 26.65083, 27.44812, 25.49966, 
    26.80661, 26.58474, 26.28732, 26.35659, 25.6816, 25.48768, 25.96575, 
    27.21079,
  10.18027, 12.59218, 16.30369, 20.30134, 23.03094, 25.2995, 26.71177, 
    23.75165, 22.87965, 25.59169, 26.37582, 26.02642, 25.71882, 25.66777, 
    26.62181,
  9.074833, 9.948637, 11.79954, 15.11935, 18.77352, 21.0163, 23.22317, 
    23.85572, 23.51437, 24.70717, 25.47446, 25.80246, 25.93773, 25.7546, 
    26.14298,
  8.873498, 8.928505, 9.447758, 11.02423, 13.93901, 16.68367, 18.6458, 
    19.83451, 20.43021, 21.21617, 22.47001, 23.91026, 25.03793, 25.73517, 
    26.43803,
  8.809943, 8.653973, 8.709722, 8.840936, 10.17951, 12.4575, 14.62996, 
    16.08266, 16.8992, 17.31058, 17.59987, 18.76179, 20.94071, 23.18233, 
    25.30271,
  8.457077, 8.369405, 8.298972, 8.17076, 8.305818, 9.218387, 10.80513, 
    12.28609, 13.39087, 13.99477, 14.0368, 14.05058, 14.89338, 17.14758, 
    20.17272,
  8.333945, 8.229517, 8.239014, 8.006861, 7.805157, 7.830093, 8.243883, 
    9.05373, 9.90432, 10.55098, 10.97373, 11.21407, 11.54003, 12.61055, 
    14.76206,
  15.89364, 15.96443, 13.07082, 12.99878, 18.66432, 26.13869, 29.25068, 
    29.33269, 28.41077, 24.58931, 23.50142, 23.18311, 22.45406, 21.98748, 
    21.60167,
  15.95635, 16.01425, 13.76335, 13.45492, 19.21393, 26.03696, 29.22773, 
    29.56287, 28.20477, 24.43558, 23.7566, 23.27365, 22.777, 21.98102, 
    22.31257,
  16.42538, 16.34451, 15.06741, 14.50226, 20.24325, 24.15286, 29.26254, 
    30.02714, 28.71345, 24.93123, 23.77597, 23.41741, 23.16892, 23.18633, 
    23.8198,
  16.2265, 16.9615, 16.53275, 16.35884, 22.00327, 26.38925, 27.16336, 
    29.92456, 28.78165, 25.54815, 24.26684, 23.63788, 23.59849, 23.96905, 
    24.66821,
  14.89283, 16.91535, 17.31465, 18.19909, 23.49259, 27.38016, 29.30141, 
    26.12815, 24.82378, 26.00991, 24.79726, 23.99446, 24.12228, 24.23696, 
    24.95854,
  12.17243, 15.62573, 17.50961, 19.02619, 23.75813, 27.03585, 29.65821, 
    29.71126, 28.41855, 27.34525, 25.61792, 24.60294, 24.73956, 24.86048, 
    25.10615,
  9.508683, 12.57224, 16.10934, 18.39138, 22.19157, 25.76192, 27.97513, 
    29.47529, 29.55541, 28.06768, 26.40375, 25.41143, 25.30497, 25.39365, 
    25.48453,
  8.059027, 9.401535, 12.76684, 16.39322, 19.68792, 23.27914, 26.20523, 
    27.86416, 28.1663, 27.42931, 26.65659, 25.85427, 25.38448, 25.28105, 
    25.26446,
  7.694977, 7.788277, 9.342004, 12.82384, 16.55544, 19.87788, 23.10805, 
    25.64283, 26.63862, 26.47124, 26.06869, 25.37641, 24.74047, 24.2238, 
    23.58016,
  7.838104, 7.552251, 7.700302, 9.335602, 12.68129, 16.22786, 19.31567, 
    22.08399, 23.8779, 24.62551, 24.62006, 24.10548, 23.42302, 22.71664, 
    21.73604,
  12.67472, 11.41633, 10.94265, 10.43629, 10.46702, 13.65997, 20.60576, 
    27.45696, 31.67653, 26.23177, 20.36061, 18.9045, 18.43421, 17.40475, 
    16.6246,
  12.83874, 11.29392, 11.05514, 10.44541, 10.43603, 13.6516, 20.82647, 
    26.91015, 30.50403, 26.01678, 20.32753, 18.87399, 18.57586, 17.89944, 
    18.30247,
  13.02777, 11.49501, 11.37807, 10.57315, 10.58222, 12.73277, 20.68116, 
    26.28288, 29.59612, 25.92903, 20.31519, 18.96258, 19.15236, 19.84696, 
    20.81637,
  13.08117, 12.18432, 11.22881, 10.87102, 11.0996, 14.08075, 19.07069, 
    25.9532, 28.91173, 25.41374, 20.67326, 19.12727, 19.55452, 20.68597, 
    21.7989,
  12.43627, 13.02664, 11.31446, 11.61755, 11.96189, 14.86348, 19.84233, 
    22.538, 24.4087, 25.27966, 21.31878, 19.43794, 19.70394, 20.41652, 
    21.67859,
  11.52712, 13.53256, 12.64555, 12.84798, 13.4104, 15.27679, 19.53663, 
    23.75667, 26.18265, 26.08444, 22.19923, 19.86249, 19.72544, 20.28538, 
    21.32511,
  10.12172, 12.68938, 13.72184, 14.30085, 15.46772, 16.26234, 18.82311, 
    23.27305, 26.18308, 26.80007, 23.42071, 20.76012, 19.87601, 20.14841, 
    20.88891,
  8.723917, 10.90507, 13.58379, 15.62401, 16.85527, 17.80191, 18.60493, 
    21.94777, 25.03655, 26.93332, 25.33991, 22.40298, 20.70709, 20.43203, 
    20.93925,
  8.397679, 8.63463, 11.42505, 15.03014, 17.5013, 19.16244, 19.32742, 
    20.99524, 24.07643, 26.44106, 27.02312, 24.80456, 22.41305, 21.42645, 
    21.5093,
  9.26048, 7.487309, 8.895594, 12.19496, 15.89468, 18.76068, 20.2854, 
    20.71408, 22.61744, 25.45657, 27.19968, 26.78003, 24.79695, 23.15795, 
    22.61774,
  11.20247, 10.68931, 10.38487, 10.11582, 9.849, 9.458875, 8.966724, 
    11.62458, 20.8364, 23.08335, 18.79443, 12.17869, 11.98668, 14.73133, 
    16.15866,
  11.32435, 10.80885, 10.48042, 10.22654, 9.847001, 9.328644, 9.379965, 
    12.41451, 19.51622, 21.64757, 16.82394, 10.99097, 11.75879, 13.45546, 
    14.48389,
  11.46175, 10.93464, 10.69311, 10.39, 9.984202, 8.569096, 10.05729, 13.7164, 
    19.51984, 20.66251, 14.72224, 11.08429, 12.24721, 14.68293, 17.04153,
  11.51979, 10.9406, 10.57606, 10.49741, 10.14313, 9.783349, 10.66742, 
    15.19839, 20.27543, 19.93004, 13.60169, 11.76301, 14.94263, 18.7249, 
    20.3604,
  11.5288, 10.89605, 10.58491, 10.66562, 10.29828, 10.86839, 13.42612, 
    15.08566, 18.0726, 19.40067, 13.55322, 13.52183, 18.52708, 21.62661, 
    22.03551,
  11.48553, 10.89786, 10.85606, 10.83564, 10.65218, 12.0909, 14.94046, 
    18.26154, 21.36585, 19.32971, 14.05002, 15.55996, 20.81448, 22.75369, 
    22.59914,
  11.26197, 10.84499, 11.21401, 10.86897, 11.00143, 13.25341, 16.18679, 
    19.82207, 23.02895, 19.11222, 14.69399, 17.0305, 21.65114, 22.84739, 
    23.03535,
  10.92125, 10.67937, 11.60607, 11.40165, 11.34426, 14.0436, 17.17238, 
    21.14727, 23.61312, 19.16516, 15.5323, 17.85402, 21.66007, 22.59587, 
    22.89856,
  10.82208, 10.15823, 11.44373, 12.33182, 12.42796, 14.89384, 17.78052, 
    21.97952, 24.2557, 19.50076, 16.60298, 18.32576, 21.23969, 21.96373, 
    22.3369,
  11.06631, 9.69854, 10.51106, 12.48145, 13.64318, 15.67704, 18.02698, 
    22.15834, 24.24379, 19.82893, 17.72895, 18.81837, 20.90178, 21.34943, 
    21.57139,
  11.13735, 10.26799, 9.699212, 9.46277, 9.46792, 9.440113, 9.344968, 
    9.648307, 12.64376, 17.89386, 17.31909, 19.44823, 21.81295, 19.06979, 
    17.35382,
  11.81064, 10.7866, 10.03258, 9.387238, 9.083305, 8.871445, 9.042868, 
    9.064712, 10.71726, 15.37783, 16.48537, 19.17399, 21.10839, 18.0887, 
    17.57075,
  11.67673, 10.88754, 10.45942, 9.823381, 8.949547, 7.652989, 8.394547, 
    8.843665, 9.632282, 13.59541, 15.70421, 18.98775, 20.57474, 18.46588, 
    18.08023,
  11.07798, 10.86705, 10.53874, 9.949553, 9.096061, 8.454979, 7.366805, 
    8.112137, 8.797331, 12.7186, 15.35799, 18.53137, 20.03369, 18.18899, 
    18.08044,
  11.17259, 10.98443, 10.3937, 9.817137, 9.278927, 8.696294, 8.301533, 
    6.502922, 6.678372, 12.09838, 14.63768, 18.42837, 19.64738, 17.47506, 
    17.71361,
  11.38857, 10.85313, 10.49714, 10.32462, 9.935654, 9.250162, 8.630021, 
    8.101003, 8.338975, 11.50357, 13.49116, 18.57388, 19.59853, 17.15844, 
    17.14721,
  11.12622, 11.03152, 11.41644, 11.60403, 11.34251, 10.52009, 9.330441, 
    8.551211, 8.324738, 10.98557, 12.60411, 18.75923, 19.97716, 17.13947, 
    16.65823,
  11.13818, 11.52751, 11.97011, 12.03227, 11.64839, 11.0446, 10.01476, 
    8.803171, 8.28686, 10.91377, 12.14941, 18.85956, 20.54295, 17.54243, 
    16.60297,
  11.33925, 11.67413, 11.98322, 12.04321, 11.69722, 11.08986, 10.34636, 
    9.180167, 8.671561, 11.20339, 11.94005, 18.96926, 20.92333, 18.29048, 
    16.95523,
  11.27893, 11.5263, 11.68995, 12.06055, 11.86002, 11.27843, 10.52814, 
    9.488717, 9.225771, 11.50312, 11.92086, 19.18975, 21.20851, 19.20739, 
    17.82002,
  11.88032, 10.95629, 9.42725, 8.410071, 8.020554, 8.088154, 9.23082, 
    11.29215, 14.58329, 18.25983, 19.80056, 20.14539, 18.93166, 18.13992, 
    17.20402,
  13.31017, 12.88827, 11.33711, 9.993632, 8.907856, 7.736219, 7.75653, 
    9.266178, 12.56286, 17.24113, 19.26846, 19.30388, 17.68852, 16.58831, 
    16.19072,
  13.6098, 13.16387, 11.92852, 10.65074, 9.83091, 7.682129, 7.600666, 
    7.842877, 9.844829, 15.42832, 18.3882, 19.05527, 17.7766, 17.48988, 
    16.44328,
  14.24943, 13.19792, 11.8209, 10.61616, 9.875998, 9.318376, 7.361887, 
    7.523442, 7.889496, 12.94628, 17.871, 18.47854, 18.41692, 18.29128, 
    16.77604,
  12.49876, 12.08397, 11.28568, 10.46229, 9.715335, 9.171323, 8.811816, 
    6.434441, 5.87449, 8.793468, 15.9683, 18.04452, 18.48977, 18.7523, 
    17.19903,
  10.22332, 10.43161, 10.5673, 10.46912, 10.136, 9.646504, 9.077819, 
    8.472917, 8.128862, 8.077406, 12.39929, 17.6983, 18.28114, 19.33956, 
    17.8677,
  10.38595, 10.5005, 10.54661, 10.60856, 10.61191, 10.47002, 9.951379, 
    9.261171, 8.593949, 8.123197, 9.515455, 16.16344, 17.69606, 19.64831, 
    18.72997,
  10.23493, 10.17066, 10.08752, 10.12573, 10.29413, 10.52049, 10.4909, 
    9.845833, 9.090178, 8.451334, 8.752976, 13.96021, 16.89555, 19.50107, 
    19.70638,
  9.752234, 9.762872, 9.892447, 10.04044, 10.10661, 10.22674, 10.39636, 
    10.24295, 9.529579, 8.755832, 8.566665, 11.97406, 15.8673, 18.57882, 
    20.38929,
  9.686715, 10.0583, 10.74483, 11.09531, 11.07567, 10.77788, 10.48991, 
    10.33948, 9.793509, 9.018047, 8.60404, 10.72566, 14.66346, 17.39311, 
    20.45876 ;

 ps =
  101029.5, 100948.3, 101092.3, 101193.2, 101319.1, 101478.1, 101571.2, 
    101658.9, 101803.2, 101718.2, 101906.6, 102368.2, 102403.8, 102097.4, 
    102104.7,
  101050.6, 100974.8, 101005.8, 101039.6, 101224.7, 101266.9, 101544, 101637, 
    101711.9, 101941, 102128.6, 102298.6, 102470.6, 100668.1, 101518.5,
  101144.6, 101084.1, 101087.9, 101113.8, 101200.6, 97804.13, 101447, 
    101733.2, 101750.6, 101895.3, 102059.5, 102186, 102370, 102558, 102746.2,
  101119.9, 101170.1, 101196.4, 101235.1, 101367.2, 101346.1, 97669.09, 
    101535.7, 101818.3, 101942.3, 102061.7, 102136.3, 102298.3, 102513.6, 
    102752,
  101040.1, 101213.3, 101286.8, 101356, 101451.6, 101592.3, 101607, 95427.53, 
    94772.33, 101866.3, 102112.1, 102154.3, 102279, 102411.6, 102697.5,
  101068.9, 101231.6, 101349.8, 101432.3, 101497, 101609.6, 101769.8, 
    101826.5, 101807.8, 102130, 102174.2, 102194.7, 102303.8, 102432.7, 
    102643.9,
  101223.7, 101368, 101468, 101569.1, 101634, 101724, 101804.4, 101969.2, 
    102088.8, 102146, 102213.2, 102282.1, 102358.3, 102474.1, 102640.2,
  101497.7, 101573.7, 101626.4, 101702.4, 101753.8, 101851.1, 101945.8, 
    102033.4, 102116.4, 102222.7, 102307, 102381.8, 102442.9, 102540.2, 
    102662.9,
  101740, 101796.8, 101838, 101902.6, 101967.5, 102036.3, 102110, 102210.9, 
    102286.9, 102354.2, 102437.2, 102513.5, 102573.9, 102677.8, 102795.5,
  101975.2, 101993.4, 102023.2, 102064.9, 102105.7, 102191, 102283.9, 
    102374.7, 102478.8, 102547.5, 102613, 102688.4, 102752.8, 102828, 102883.5,
  100537.1, 100555.7, 100697.4, 100621.5, 100624.3, 100432.4, 100179.9, 
    99936.51, 99790.98, 99442.31, 99576.24, 100075.7, 100235.7, 100245, 100561,
  100556.9, 100481.4, 100575, 100650.8, 100717.6, 100402.3, 100424.5, 
    100181.8, 100008.1, 100028.6, 100096.5, 100349.3, 100620.7, 99122.48, 
    100219.4,
  100729.8, 100622.4, 100612.5, 100694.4, 100663.8, 97136.84, 100475.3, 
    100533.9, 100406.2, 100349.5, 100399.5, 100596.7, 100920, 101220.6, 
    101620.7,
  100933, 100864.2, 100828.8, 100820.8, 100882.9, 100657.2, 96918.36, 
    100489.6, 100613.5, 100660.1, 100711.7, 100864, 101167.1, 101551.7, 
    101913.1,
  101101.2, 101059.3, 101028.5, 101011.7, 101010.2, 101022.5, 100886.7, 
    94677.49, 94048.63, 100785.7, 101021.3, 101142, 101401.2, 101685, 102113.5,
  101268.6, 101230.3, 101188, 101166.6, 101144.2, 101126.6, 101165.3, 
    101126.3, 100961, 101222.7, 101295.4, 101394.4, 101627.9, 101917.3, 
    102265.1,
  101405.5, 101396.1, 101351.8, 101337.1, 101319.7, 101322.4, 101293.5, 
    101360.6, 101428, 101442.8, 101532.7, 101653, 101827.2, 102080.8, 102387,
  101556.9, 101546.7, 101510.2, 101481.9, 101435, 101430.6, 101441.1, 
    101442.1, 101480.2, 101614.6, 101760.2, 101887.9, 102053.3, 102277.8, 
    102548.1,
  101701, 101701.6, 101682.9, 101667, 101647.6, 101616.2, 101594.5, 101642, 
    101707.9, 101796.9, 101929, 102079.3, 102219.7, 102421.1, 102660.7,
  101854.8, 101852.3, 101835.5, 101827.6, 101801.2, 101816.8, 101834.2, 
    101847.5, 101895.2, 101966.2, 102094.7, 102246.5, 102373.6, 102559, 
    102759.1,
  100628.5, 100465, 100375.5, 100278.3, 100217.6, 100145.7, 99986.81, 
    99856.74, 99804.44, 99611.55, 99902.02, 100501.8, 100628, 100499.4, 100576,
  100602.7, 100477, 100332.9, 100206.7, 100089.1, 99797.42, 99879.91, 
    99692.3, 99602.45, 99854.79, 100132.6, 100506.1, 100765.2, 99172.52, 
    100109.8,
  100638.4, 100494.2, 100337.7, 100175.5, 99856.27, 96335.68, 99626.51, 
    99742.22, 99678.09, 99891.75, 100145.1, 100491.9, 100850.9, 101127.5, 
    101418.9,
  100655.5, 100517.4, 100378.3, 100181.2, 100001.6, 99580.81, 95923.34, 
    99457.01, 99644.83, 99909.08, 100206, 100513.3, 100885.5, 101284.1, 
    101606.8,
  100701.6, 100571.9, 100444.7, 100267.9, 100070.8, 99847.27, 99600.41, 
    93606.07, 93093.51, 99810.66, 100284, 100578.6, 100963, 101303, 101737.3,
  100760.6, 100650.2, 100517.5, 100370.6, 100166.3, 99931.4, 99810.04, 
    99767.23, 99613.07, 100089.5, 100346.4, 100684.2, 101063.7, 101464.8, 
    101845.8,
  100850.6, 100759.6, 100636.1, 100502.6, 100327.4, 100126.4, 99918.5, 
    99955.42, 100072.9, 100192.6, 100460, 100815.6, 101180.1, 101571.6, 
    101944.3,
  100968.6, 100889.3, 100774.1, 100651.3, 100471.4, 100305.8, 100171.6, 
    100087.8, 100127.5, 100339.5, 100649.4, 100972.9, 101346.9, 101725.2, 
    102156.4,
  101100.2, 101045.3, 100954.6, 100845.1, 100703.5, 100544.4, 100418.8, 
    100410, 100485.5, 100633.2, 100904.5, 101207, 101551.2, 101948.5, 102379.7,
  101264.4, 101203.2, 101131.4, 101042.2, 100914.1, 100794.7, 100707.1, 
    100664.7, 100724.4, 100887, 101179, 101486.3, 101821.5, 102229.4, 102579.2,
  101102.3, 100968.4, 100913, 100815, 100785.3, 100814.2, 100967.7, 101229.6, 
    101476.6, 101386.6, 101627.2, 102207.3, 102351.5, 102147.4, 102113.1,
  100910.8, 100802.4, 100756, 100703.5, 100704.4, 100579.9, 100866.7, 
    101068.5, 101291.5, 101625.7, 101893.1, 102274.1, 102538.9, 100813, 
    101658.5,
  100787, 100727.6, 100704.3, 100663.3, 100516.3, 97133.28, 100668.9, 
    101050.4, 101332, 101640, 101936.6, 102306.9, 102654.6, 102850.2, 102981.4,
  100669.7, 100652.6, 100626.8, 100580.1, 100550.3, 100390.8, 96920.89, 
    100806, 101277.3, 101659.6, 102034.8, 102355.8, 102694.4, 102960.3, 
    103119.3,
  100611.1, 100611.5, 100572.9, 100528.8, 100481.3, 100522.8, 100618.9, 
    94897.48, 94547.84, 101582.3, 102155, 102440.7, 102756.5, 102922.1, 
    103177.4,
  100574.1, 100568.5, 100503.4, 100446.4, 100408.8, 100417.5, 100779.9, 
    100991.9, 101146.6, 101849.8, 102203.5, 102523.9, 102807.2, 103018.6, 
    103236.3,
  100559.4, 100549.6, 100468.4, 100399.6, 100385.6, 100443.9, 100724.8, 
    101199.9, 101630.1, 101906.1, 102281.5, 102612, 102851.5, 103098.6, 
    103326.2,
  100573, 100538.9, 100438.2, 100348.1, 100344.9, 100471, 100829.9, 101155.5, 
    101523.5, 101965.5, 102376.8, 102682.8, 102968.5, 103244.1, 103512.3,
  100610.4, 100580, 100463, 100377.5, 100407.2, 100586.5, 100939, 101352.6, 
    101741, 102088.1, 102482.9, 102799.9, 103103, 103405.7, 103705.2,
  100674.2, 100626.7, 100494.2, 100429, 100493.2, 100744, 101088.1, 101407.8, 
    101771.6, 102188.7, 102612, 102947.4, 103286.2, 103622.9, 103899,
  102304.9, 102268.4, 102314, 102330.4, 102373.2, 102475.9, 102726.4, 
    103068.2, 103348.8, 103229.7, 103472.1, 103973.6, 103948.8, 103549.4, 
    103339.3,
  102071.6, 102032.6, 102041.2, 102077.5, 102267.2, 102358.4, 102831.1, 
    103084, 103286.2, 103577.3, 103800.7, 104047.4, 104143.2, 102191.2, 
    102902.4,
  101852.6, 101842.2, 101877.4, 101965.3, 102144.1, 98947.41, 102729.1, 
    103200.1, 103457.2, 103647.6, 103859.8, 104087.3, 104260.3, 104255.6, 
    104245.6,
  101656.5, 101671.6, 101738.4, 101854.5, 102196.9, 102246, 98853.62, 
    102898.7, 103361.6, 103647.4, 103947.5, 104125, 104297.1, 104371.8, 104388,
  101446.6, 101531.7, 101640, 101809.3, 102107, 102420.9, 102558.8, 96755.73, 
    96354.45, 103500.6, 104022.2, 104191.4, 104365.7, 104364.6, 104441.1,
  101278.2, 101410.6, 101554.7, 101739.3, 102016.6, 102282.7, 102718, 
    102918.7, 103036.4, 103748.3, 104028.8, 104251.8, 104404.5, 104464.8, 
    104495.8,
  101142.8, 101343.4, 101515.1, 101717.1, 101968.1, 102214.1, 102591.7, 
    103063.1, 103476, 103744.5, 104052.8, 104322.7, 104441.9, 104514.4, 
    104544.5,
  101048.9, 101292.6, 101482.4, 101685.1, 101890.3, 102139.5, 102586.6, 
    102921.6, 103309.6, 103719.4, 104118.3, 104363.6, 104500.6, 104582.9, 
    104645.3,
  101007.4, 101292.8, 101501.1, 101697.9, 101894.6, 102149.6, 102597.4, 
    103041.7, 103446.3, 103786.7, 104166.5, 104406.5, 104540.3, 104638, 104718,
  101006.8, 101298.2, 101498.9, 101691.1, 101902.4, 102218.5, 102679.4, 
    103024.9, 103414.4, 103817.7, 104213.5, 104444.3, 104598.3, 104727.2, 
    104799.7,
  103276.3, 103369, 103545, 103679.1, 103891.3, 104065.9, 104233.9, 104514, 
    104740.8, 104510.3, 104592.5, 104828.6, 104518.1, 103920.3, 103673.9,
  103084.7, 103187.5, 103361.6, 103523.7, 103777.9, 103837.1, 104251.1, 
    104476.5, 104638.3, 104845.5, 104913.3, 104904.4, 104722.9, 102611.2, 
    103268.3,
  102903.5, 103038.8, 103210.2, 103381.4, 103576, 100309.8, 104124.5, 
    104618.2, 104807.5, 104890, 104940.7, 104941.1, 104829, 104687.6, 104601.5,
  102748.3, 102875, 103054, 103209.6, 103547.1, 103620.9, 100162.9, 104226.6, 
    104636.8, 104853.9, 104982.8, 104956, 104871.7, 104763.5, 104736.5,
  102588, 102726.5, 102902.9, 103066.8, 103368.5, 103763.7, 103860.1, 
    97953.4, 97457.62, 104576.4, 105008.7, 104977.8, 104927.6, 104786.5, 
    104773.9,
  102411.9, 102553.8, 102730, 102900.6, 103183.8, 103542.9, 103941.9, 
    104139.7, 104156, 104807.3, 104950.3, 104996.6, 104942.6, 104884.5, 
    104835.4,
  102217.9, 102396.6, 102576.3, 102754.7, 103051.9, 103412, 103748.1, 
    104208.9, 104544.9, 104726.5, 104905.6, 105020.1, 104970.4, 104944.3, 
    104884.8,
  102010.2, 102216.4, 102400.3, 102611, 102914.3, 103261.6, 103636.4, 
    103940.5, 104270.2, 104634.7, 104900.7, 105006.6, 105007.5, 104996.6, 
    104955.5,
  101835.4, 102077.4, 102283.1, 102509.2, 102849.9, 103172.8, 103551.9, 
    103965.8, 104346.6, 104572, 104872.8, 105006.9, 105046.8, 105038.1, 
    104994.9,
  101681.7, 101926.9, 102170.8, 102422.2, 102771.7, 103099.2, 103489.6, 
    103815.1, 104164.2, 104483.3, 104843.2, 105000.2, 105068.7, 105069.6, 
    105015,
  103759.6, 103860.2, 104067.4, 104235.8, 104476.9, 104644.1, 104719.7, 
    104802.3, 104780.9, 104312.4, 104219.7, 104357, 104166, 103709, 103522.2,
  103626.9, 103729.1, 103935.5, 104150.2, 104422.8, 104437.4, 104734.8, 
    104795, 104748.2, 104717, 104576.7, 104473.6, 104377.3, 102413.7, 103143.1,
  103475.2, 103622.1, 103828.9, 104069.9, 104278.4, 100837.1, 104597, 
    104919.1, 104938.3, 104814.3, 104691, 104563.6, 104500.7, 104500.9, 
    104487.7,
  103316.2, 103484.1, 103699.5, 103941.2, 104302.1, 104248.4, 100639.9, 
    104555.7, 104812, 104856.4, 104798.6, 104646.9, 104577.7, 104580.8, 
    104627.2,
  103127.3, 103333, 103560.1, 103842.5, 104157.1, 104466.8, 104448.3, 
    98348.58, 97636.8, 104644.7, 104878, 104740, 104670.5, 104590.9, 104628.3,
  102924.6, 103142.6, 103382.4, 103693.2, 104018.8, 104280.7, 104583.6, 
    104603.8, 104506, 104879.4, 104896.6, 104833.9, 104746, 104697, 104661.1,
  102697.6, 102954.3, 103228.7, 103549.3, 103914.9, 104202.2, 104405.9, 
    104652.8, 104795.9, 104845.3, 104928.8, 104918.8, 104833.5, 104780.8, 
    104743.7,
  102462, 102735.1, 103037.6, 103389.8, 103741.7, 104064.9, 104303.5, 
    104447.5, 104612.9, 104831.8, 104971.2, 104974.2, 104922.4, 104852.9, 
    104817.4,
  102248.6, 102568.7, 102894.8, 103257.4, 103643.3, 103960.2, 104182.5, 
    104390.8, 104638.2, 104770.3, 104979.8, 105030.4, 105004.7, 104932, 
    104872.7,
  102060.8, 102375.1, 102726.6, 103108.9, 103483.5, 103827.2, 104065.3, 
    104207.8, 104451.2, 104672.2, 104951.6, 105041.3, 105063.1, 105006, 
    104938.3,
  103193.1, 103300.4, 103550.5, 103705.6, 103901.7, 103975.6, 103946.9, 
    103961, 103999.4, 103724.5, 103878.3, 104252.3, 104148.4, 103721.8, 
    103567.5,
  102986.9, 103108.9, 103390, 103605.1, 103862.6, 103802.8, 103997.9, 
    103973.4, 103960.8, 104064.6, 104151.6, 104289.9, 104329, 102403.7, 103171,
  102762.4, 102945.7, 103254.2, 103522.3, 103713.8, 100226.2, 103879.4, 
    104063.2, 104079.1, 104082.1, 104167.3, 104273.7, 104411, 104473.8, 
    104514.3,
  102569.1, 102779.1, 103114.1, 103396.1, 103748.6, 103644, 99957.77, 
    103786.7, 104005.3, 104102.4, 104179.2, 104267.7, 104397.2, 104532.8, 
    104627,
  102432.6, 102674.9, 103014, 103320.3, 103628.8, 103859.5, 103795, 97625.81, 
    96979.18, 103907.8, 104203.5, 104269.5, 104411.3, 104486, 104621.3,
  102351.6, 102595.2, 102916.1, 103236.6, 103529.9, 103696.1, 103946.2, 
    103926.8, 103814.8, 104112.1, 104203.5, 104270.9, 104392.8, 104482, 
    104574.9,
  102330.5, 102564.9, 102870.3, 103155.8, 103458.8, 103668.4, 103818.7, 
    103962.5, 104046.7, 104106.1, 104211, 104302, 104394.7, 104477, 104548.2,
  102292.8, 102505.9, 102769.5, 103060.3, 103336, 103563.9, 103783.5, 
    103872.4, 103965.9, 104119.4, 104249.2, 104325.7, 104413, 104513.6, 
    104603.1,
  102212.2, 102430.5, 102692.5, 102957.4, 103253.3, 103492.3, 103712.8, 
    103894.4, 104010, 104162.9, 104295.7, 104381.1, 104459.2, 104556.4, 
    104637.2,
  102069.9, 102268.6, 102526.6, 102821.1, 103118.2, 103379.9, 103635, 
    103816.2, 103954, 104139.8, 104314.3, 104429.4, 104511.1, 104609.2, 
    104670.3,
  102369.4, 102545.6, 102884.8, 103142.5, 103401.9, 103586.6, 103762.8, 
    103955.5, 104095.9, 103807.4, 103881.5, 104151.8, 103938.6, 103417.9, 
    103175.7,
  102214.1, 102386.4, 102736.4, 103040.6, 103353.3, 103395.6, 103762.7, 
    103932.7, 104045.2, 104196.7, 104238.6, 104278.1, 104202.2, 102184.5, 
    102809.8,
  102102.3, 102269.1, 102626.6, 102961.2, 103193.6, 99820.82, 103592.5, 
    103999.3, 104161.2, 104234.6, 104293.2, 104332.1, 104330.9, 104284.5, 
    104179,
  102023.8, 102165.7, 102539.1, 102853.9, 103260.8, 103182.2, 99665.33, 
    103614.1, 104032.3, 104203.5, 104329.6, 104349.8, 104384.5, 104375.5, 
    104326.7,
  101953, 102110.8, 102473.4, 102803.1, 103145.5, 103446.8, 103410.1, 
    97432.34, 96833.93, 103866.9, 104314, 104338, 104413.4, 104369.2, 104384,
  101917.8, 102090.1, 102434.4, 102770, 103051.2, 103246.8, 103549.2, 
    103601.5, 103552.9, 104033.5, 104202.4, 104311.6, 104392.8, 104410.3, 
    104413.9,
  101958.4, 102130.6, 102447.1, 102741.9, 103025.1, 103211.5, 103370.1, 
    103615.9, 103784, 103911.6, 104102.2, 104266.4, 104356.5, 104402.4, 104404,
  102010.8, 102193.3, 102463, 102740.4, 102954.5, 103129.2, 103300.3, 
    103394.5, 103542.2, 103785.7, 104040.7, 104198.9, 104326.5, 104399, 
    104446.3,
  102075.1, 102254.1, 102486.2, 102719.8, 102935.7, 103098.9, 103242, 
    103390.9, 103521.4, 103702.6, 103966.4, 104140.9, 104283.7, 104380.6, 
    104458.7,
  102083.9, 102236.4, 102454.2, 102685.2, 102875.5, 103017.9, 103179.8, 
    103279, 103395.3, 103607.3, 103895.3, 104081.8, 104239.6, 104372.3, 
    104477.4,
  102968.5, 103160.6, 103404.4, 103522.8, 103672.1, 103746.2, 103750.1, 
    103744.6, 103680.4, 103243.1, 103167.5, 103272.7, 102959, 102360.7, 
    102081.7,
  102918.8, 103093.1, 103336.6, 103534.5, 103732.3, 103634.2, 103845.9, 
    103819, 103735, 103703.2, 103567.8, 103445.4, 103228.2, 101138.1, 101674.3,
  102861.6, 103060.4, 103298.2, 103537.7, 103595.9, 100129.6, 103785.4, 
    104002.6, 103963.8, 103835.9, 103713.9, 103579.1, 103414, 103242.2, 
    103041.6,
  102810.4, 103009.6, 103263.6, 103455.2, 103745.3, 103569.3, 99880.36, 
    103685.7, 103866.9, 103929.6, 103851.3, 103704.6, 103564.6, 103410, 
    103247.5,
  102758.1, 102965.2, 103220, 103398.8, 103623.6, 103828.7, 103742.4, 
    97520.19, 96799.41, 103723.3, 103960.4, 103815.8, 103717.8, 103531, 
    103449.2,
  102727, 102915.4, 103145.9, 103343.8, 103530.6, 103656.3, 103843.4, 
    103833.9, 103711.7, 103940.8, 103993.7, 103926.6, 103851.4, 103723.7, 
    103621.2,
  102676.3, 102855.9, 103073.7, 103244.1, 103436, 103568.8, 103703.3, 
    103806.9, 103911.1, 103949.6, 104015.1, 104026.2, 103971.6, 103892.9, 
    103815,
  102625.5, 102775.8, 102971.7, 103142.8, 103314.9, 103432.8, 103564.1, 
    103658.4, 103734, 103891.3, 104039.5, 104084.7, 104096.3, 104061.6, 
    104024.5,
  102525.8, 102674.2, 102868.3, 103022.9, 103185.8, 103323.9, 103437.2, 
    103557.9, 103697.6, 103825, 104023.6, 104125, 104180.3, 104196.7, 104192.7,
  102407.9, 102520.1, 102700.9, 102879.7, 103063.4, 103176.8, 103316.1, 
    103416.5, 103516.2, 103699.6, 103955.9, 104122.5, 104228.5, 104300, 
    104328.6,
  103828.1, 103860.8, 103953.7, 103879.3, 103895.7, 103802, 103650.5, 
    103528.5, 103380.5, 102831.4, 102722, 102826.5, 102567.1, 102021, 101766.4,
  103768.9, 103787.6, 103859.4, 103875.6, 103923.1, 103620.6, 103765.5, 
    103550.1, 103387.1, 103261.8, 103079.7, 102966.2, 102806.1, 100781.3, 
    101350.2,
  103702.4, 103767.3, 103813.8, 103884.4, 103751.7, 100191.9, 103601.4, 
    103809, 103620.3, 103413.1, 103211.4, 103081.8, 102956.2, 102850, 102682.1,
  103637, 103701.2, 103772.9, 103814.8, 103882.4, 103590.8, 99810.02, 
    103428.6, 103562.9, 103540.9, 103376.5, 103218.3, 103103.6, 103001.5, 
    102880.3,
  103567.6, 103641.5, 103730.7, 103762.4, 103827.4, 103810.9, 103649.9, 
    97399.87, 96731.63, 103456, 103563, 103380.9, 103302.7, 103155.5, 103091.6,
  103443.2, 103531.8, 103611, 103683.5, 103728.3, 103744.7, 103745.4, 
    103726.3, 103572.8, 103762.9, 103695.1, 103569.1, 103490.5, 103387.5, 
    103292.3,
  103253.6, 103354.8, 103455.4, 103545.9, 103619.9, 103677, 103711.3, 
    103769.6, 103882.3, 103863.6, 103817.1, 103748.4, 103672.3, 103599.5, 
    103507.5,
  102999.5, 103087.1, 103195.1, 103315.9, 103426.2, 103527.1, 103603.8, 
    103644, 103738.1, 103884.7, 103933.9, 103893, 103854.8, 103795.6, 103726.2,
  102689, 102759.2, 102871.8, 103049.4, 103219.6, 103369, 103475.8, 103589.5, 
    103740.6, 103920, 104005, 104021.5, 104004.6, 103974.6, 103913.6,
  102347.1, 102375.8, 102452.7, 102662.4, 102945.5, 103171.8, 103350.6, 
    103459.7, 103604.3, 103825.5, 104001.3, 104099.8, 104126.3, 104127.8, 
    104073.6,
  104309.2, 104264.7, 104244.9, 104149.1, 104154.9, 104097.1, 103942.7, 
    103812.8, 103673.4, 103185.6, 103093.6, 103161.3, 102826.4, 102199.7, 
    101861.8,
  104193.5, 104169.9, 104088.2, 104039.3, 104083.5, 103869.4, 104019, 
    103859.4, 103708.6, 103605.2, 103438.7, 103288.1, 103045.2, 100925.3, 
    101379.8,
  104050.8, 104074.8, 104027.6, 104012.3, 103841.2, 100363.6, 103857.5, 
    104009, 103871.4, 103734.3, 103564.3, 103406.2, 103198.4, 102976.5, 
    102667.5,
  103889.9, 103933.5, 103951.1, 103918.7, 103877, 103678.8, 99996.54, 
    103733.4, 103876.9, 103830, 103705.6, 103529.4, 103339.7, 103112.9, 
    102820.3,
  103731.7, 103770.4, 103803.2, 103799.1, 103821.7, 103816, 103822, 97610.8, 
    96937.23, 103701.9, 103837.6, 103659.1, 103494.2, 103236.1, 103004.4,
  103508.1, 103558.1, 103617, 103665.7, 103690, 103731.1, 103854.9, 103940.9, 
    103800.3, 103976.9, 103918.4, 103796.1, 103631.7, 103409.3, 103167.3,
  103219.2, 103326.2, 103377.4, 103463.9, 103537.6, 103637.7, 103750.1, 
    103951.6, 104040, 104025.6, 103990.4, 103910.2, 103770.1, 103572.9, 
    103337.7,
  102802.4, 102947.8, 103103.5, 103260, 103347.9, 103479.3, 103617.5, 
    103777.2, 103895.7, 104003, 104040.1, 103991.4, 103897.6, 103736.1, 103534,
  102616.9, 102652.6, 102726, 102875.8, 103084.9, 103292.9, 103453.3, 
    103610.7, 103765.1, 103941.4, 104028.3, 104043.7, 103990.5, 103868.3, 
    103690,
  102722.2, 102683.4, 102643.2, 102670.7, 102796.5, 103027.3, 103257.9, 
    103413.8, 103554.4, 103741.6, 103941, 104026, 104036.5, 103973.9, 103836.7,
  104226.1, 104281.9, 104324.6, 104238.4, 104264.7, 104307.1, 104293, 
    104218.9, 104073.2, 103545, 103362.1, 103321.6, 102853.2, 102112.4, 
    101715.2,
  104166.2, 104200.7, 104151.2, 104073.2, 104149.8, 104075, 104262.1, 104194, 
    104056.7, 103928.7, 103690.1, 103437.2, 103065.2, 100861.9, 101239,
  104056.8, 104142.5, 104150.6, 104083.2, 103934.2, 100506.6, 104035, 
    104262.8, 104162.6, 104003.8, 103780.6, 103526.7, 103208.3, 102910.4, 
    102535,
  103922.4, 104036.3, 104082.2, 104061.7, 103972.1, 103834, 100106.4, 
    103868.3, 104037.9, 104030.8, 103869.7, 103615.8, 103338, 103031.4, 
    102698.3,
  103773, 103891.7, 103962, 103988.1, 103933.4, 103895.5, 103893.3, 97734.18, 
    97016.82, 103816.3, 103928.8, 103694.8, 103471.2, 103155.1, 102885.9,
  103602.4, 103729.6, 103803.3, 103856.3, 103839.6, 103795.9, 103881.1, 
    103929.6, 103823.5, 103994.2, 103923.5, 103755.8, 103563.4, 103303.4, 
    103031.4,
  103377.1, 103529.6, 103619.8, 103705.7, 103738.3, 103737.5, 103749, 
    103844.7, 103946.9, 103953.6, 103882.3, 103772.3, 103625, 103421.5, 
    103170.7,
  103127, 103315.5, 103421.9, 103526.9, 103560.7, 103589.8, 103604.9, 103659, 
    103697.8, 103766.5, 103771.1, 103718.2, 103629, 103493.5, 103307,
  102884.5, 103044.8, 103166.5, 103275.5, 103356.3, 103412, 103422.9, 
    103462.5, 103510.2, 103538.7, 103565.4, 103575.4, 103557.6, 103496.5, 
    103372.3,
  102777.8, 102872.5, 102942.7, 103024.4, 103080, 103130.7, 103174.1, 
    103200.1, 103225.2, 103245.3, 103318.7, 103368.4, 103397, 103410.4, 
    103362.6,
  102873.3, 103161.6, 103462.9, 103712.8, 103920.3, 104055.1, 104104, 
    104141.4, 104083.2, 103639.4, 103553.8, 103583.8, 103190.3, 102506.4, 
    102166.3,
  102965.5, 103195, 103452.3, 103677.1, 103860.5, 103836.2, 104051.3, 
    104047.5, 103988.1, 103951.9, 103824.3, 103656.9, 103379.4, 101230.4, 
    101667.1,
  103014.3, 103210.1, 103417.7, 103648.1, 103711.5, 100257.2, 103828.8, 
    104081.6, 104049.1, 103942.6, 103824.7, 103674.5, 103447, 103211, 102918.7,
  103058.7, 103236.1, 103422.4, 103580.6, 103752.5, 103601.2, 99929.71, 
    103663.4, 103805.8, 103851.2, 103799.5, 103662.3, 103461.7, 103244.8, 
    102986.9,
  103094.5, 103266, 103440.9, 103575.2, 103677.9, 103755.1, 103665.2, 
    97565.35, 96834.14, 103536.7, 103742.6, 103603.9, 103434.1, 103215, 103052,
  103093.8, 103269.4, 103417, 103546.5, 103615.6, 103652.7, 103682.9, 
    103635.6, 103490.9, 103651.3, 103634, 103520.8, 103371.8, 103186.2, 
    103049.7,
  103063.1, 103229.7, 103364.5, 103480.1, 103554.3, 103600.3, 103584.8, 
    103559.1, 103526.9, 103509.2, 103466.3, 103382.1, 103250.1, 103120.3, 
    103007.6,
  102993.4, 103151.7, 103261.4, 103362.1, 103400, 103430.3, 103430.2, 
    103401.4, 103347.2, 103311, 103262.5, 103190, 103104.6, 103027.4, 102958.9,
  102879.9, 103015.7, 103110.9, 103191, 103231.1, 103245.1, 103221.1, 
    103198.7, 103153.3, 103103.4, 103052.2, 102998.2, 102940.4, 102898.1, 
    102852.7,
  102709.5, 102825.6, 102896.1, 102946.2, 102956.6, 102960.6, 102950.4, 
    102917.3, 102868.4, 102808.6, 102803.1, 102776.1, 102746.9, 102730.6, 
    102713.4,
  102067.3, 102302.3, 102630.2, 102941.8, 103285.7, 103564.2, 103730.3, 
    103857, 103904.6, 103519.8, 103458, 103523.7, 103105.5, 102396, 102107.5,
  102063, 102278.6, 102602.6, 102958.5, 103269, 103385.8, 103723, 103828.8, 
    103784.7, 103778, 103642.6, 103498.3, 103206.1, 101079.7, 101632.3,
  102008, 102257.2, 102584.5, 102973.3, 103152.1, 99864.4, 103550.5, 
    103843.1, 103835.2, 103714.1, 103581, 103427.2, 103187.1, 103000.8, 
    102899.9,
  101969.5, 102226.3, 102568.8, 102904.1, 103258.2, 103189.8, 99653.16, 
    103441.5, 103635.3, 103600, 103535.9, 103368.9, 103165.6, 103004.6, 
    102983.3,
  101964.1, 102223.7, 102566.2, 102886.6, 103195, 103477.4, 103385.4, 
    97375.17, 96658.69, 103363.1, 103486.7, 103334.6, 103161.9, 102974.7, 
    103011.6,
  101982.8, 102247.6, 102556.5, 102861.5, 103103.7, 103312.5, 103543.8, 
    103508, 103437.3, 103524.9, 103430.1, 103299.3, 103144.4, 102991.1, 
    102956.1,
  102027.2, 102289.9, 102580.4, 102842.5, 103087.6, 103261.2, 103403.1, 
    103505.7, 103516.7, 103440.8, 103352.2, 103240.2, 103105.2, 102975.9, 
    102915,
  102088.2, 102335.1, 102583, 102812.2, 102996.2, 103168.4, 103292.5, 
    103350.4, 103339.3, 103317.4, 103246.1, 103156.4, 103047.8, 102937.5, 
    102859.8,
  102171.6, 102391.2, 102606.6, 102802.6, 102962.3, 103085.5, 103163, 
    103218.3, 103201.6, 103158.2, 103096, 103017.6, 102929.1, 102843.5, 
    102777.7,
  102242, 102416, 102580, 102729.8, 102846.6, 102940.7, 103000.1, 103005.5, 
    102978.4, 102919.8, 102890.2, 102829.7, 102758.7, 102700.1, 102646.5,
  102315.4, 102574.7, 102857, 103100.8, 103356.3, 103547.2, 103648.7, 
    103700.9, 103618, 103137.4, 103049.8, 103245.3, 103069.7, 102555.1, 
    102288.9,
  102295.6, 102546.5, 102837.4, 103121.7, 103348.4, 103381.8, 103665.6, 
    103708.1, 103605.4, 103506, 103333, 103250.5, 103182.2, 101182.6, 101741.8,
  102251.9, 102529.7, 102792.4, 103101, 103217.6, 99840.76, 103527.6, 
    103773.6, 103709.2, 103548.5, 103407.7, 103263.6, 103167.7, 103084.6, 
    102926.9,
  102217.8, 102479.6, 102729.9, 102990.6, 103275.2, 103185.2, 99605.99, 
    103400.6, 103610.5, 103555.1, 103475, 103323.8, 103169.9, 103060.4, 
    102948.5,
  102178.4, 102414.7, 102645.6, 102898.9, 103140.8, 103405.8, 103341.9, 
    97318.23, 96647.69, 103394.6, 103521.3, 103385.4, 103231.6, 103050.2, 
    102950.1,
  102126.9, 102337.2, 102535.9, 102777.9, 102984.8, 103194.2, 103427.9, 
    103444.6, 103395.5, 103614.2, 103539.1, 103426.8, 103278.3, 103089.5, 
    102943.6,
  102042.3, 102231.7, 102420.6, 102640.7, 102865.9, 103066.2, 103247.9, 
    103440.7, 103571.7, 103585.4, 103536.9, 103441, 103302.7, 103119, 102935.3,
  101951.8, 102113.1, 102290.5, 102497.9, 102698.3, 102908.5, 103098.9, 
    103236.6, 103369.9, 103475.1, 103487.7, 103414.6, 103287.9, 103127.8, 
    102948.2,
  101869.6, 102012.4, 102185.3, 102376.3, 102573.9, 102763.1, 102949.3, 
    103131.1, 103263.8, 103348.8, 103370, 103324.9, 103230.3, 103083.2, 
    102927.9,
  101829, 101957.3, 102115.3, 102280.3, 102453.1, 102627.4, 102795.2, 
    102936.1, 103047.9, 103127.9, 103205.1, 103194.9, 103122.5, 103014.6, 
    102890.9,
  102862, 103056.2, 103268.4, 103405.2, 103557.1, 103624.7, 103620.3, 
    103541.5, 103413.7, 102880.9, 102733.1, 102702.1, 102237.2, 101546.9, 
    101323.7,
  102841.3, 103021.8, 103227.9, 103414.2, 103544, 103467.8, 103643.5, 
    103541.8, 103411.5, 103266.3, 103057.1, 102824.1, 102476.6, 100351.5, 
    100932.7,
  102768.8, 102972.5, 103147.8, 103358.7, 103374.2, 99878.82, 103432.9, 
    103639.4, 103507.6, 103309.2, 103135.3, 102920.9, 102623.6, 102399, 
    102271.1,
  102681, 102881.5, 103053.5, 103213.4, 103387.6, 103243.2, 99524.21, 
    103163.1, 103350.8, 103315.1, 103191.9, 103003.6, 102747.9, 102549.1, 
    102447.4,
  102589.9, 102773.8, 102938.5, 103080.7, 103205.2, 103309.8, 103216.4, 
    97134.6, 96372.83, 103064.3, 103234.7, 103069.9, 102867.9, 102622.1, 
    102601.7,
  102474.2, 102652, 102802.7, 102939.7, 103028.4, 103096.9, 103169.6, 
    103143.2, 103035, 103232.8, 103211.4, 103114.8, 102964.3, 102754.2, 
    102707.8,
  102367, 102529.3, 102659.1, 102774.3, 102854.3, 102914.5, 102949.1, 103020, 
    103067.9, 103103.3, 103154, 103126.9, 103020.3, 102829.1, 102767.6,
  102255.2, 102388.2, 102496.4, 102599.6, 102659, 102714.7, 102758.9, 
    102778.5, 102820.9, 102934.8, 103039, 103079.6, 103053.8, 102917.5, 102834,
  102141.2, 102258.5, 102339.9, 102411.9, 102474.5, 102523, 102562.5, 
    102643.4, 102692.9, 102772.5, 102892.7, 102995.2, 103020.5, 102945.1, 
    102837.8,
  102037.4, 102101.3, 102160.3, 102213.7, 102250.3, 102298.9, 102350.4, 
    102387.4, 102458.8, 102530.2, 102712.8, 102857.6, 102938, 102943.6, 
    102860.9,
  103046.7, 103179.9, 103321.9, 103388.1, 103456.4, 103402.6, 103288.8, 
    103196.4, 103085.9, 102658, 102671.1, 102940.2, 102828.3, 102369.1, 
    102157.2,
  103108.6, 103232.1, 103361.5, 103451.5, 103456.3, 103203.4, 103314.3, 
    103125.1, 103010, 103020.8, 102995, 103044.2, 103056.8, 101102.2, 101801.8,
  103110.3, 103251.4, 103337.5, 103443.1, 103290.3, 99743.12, 103102.5, 
    103277.1, 103121.8, 103060.9, 103034.3, 103117.6, 103195.3, 103265.5, 
    103211.4,
  103094.5, 103226.1, 103290.8, 103327.4, 103315.6, 103069.5, 99267.49, 
    102788.4, 102911.4, 103053.5, 103069.1, 103137.8, 103246.8, 103379.6, 
    103383.6,
  103058.7, 103150.9, 103207.8, 103212.8, 103189.4, 103116.9, 102897.9, 
    96830.1, 96084.48, 102706.5, 103094.5, 103123.9, 103291.6, 103375.9, 
    103478.4,
  102942.5, 103042.1, 103072.3, 103083.6, 103022.5, 102968.5, 102890.8, 
    102779.6, 102596.4, 102808, 103043.5, 103095.8, 103270.5, 103401.4, 
    103493.4,
  102837.7, 102888.9, 102911.9, 102904.9, 102861.2, 102795.4, 102730.1, 
    102722.9, 102716.5, 102746.9, 102954.1, 103065.2, 103212.8, 103374.5, 
    103485.8,
  102708, 102735.5, 102725.9, 102718.5, 102661.5, 102621.2, 102593.4, 102572, 
    102590.4, 102669.7, 102861.5, 103004.9, 103137.7, 103320.6, 103460.4,
  102540.5, 102578.3, 102579.5, 102552.2, 102519.6, 102500.7, 102491, 
    102516.6, 102556, 102601.5, 102730.7, 102946.5, 103072.7, 103219.9, 
    103387.9,
  102347.6, 102379.6, 102386.2, 102382.6, 102372.8, 102366.3, 102367.5, 
    102338, 102354, 102417.7, 102585.9, 102801.4, 102974.1, 103126.8, 103230.6,
  103667.3, 103709.7, 103729.4, 103650.1, 103553.1, 103410.3, 103218.3, 
    103225.4, 103328.2, 103037.4, 103117.1, 103357.1, 103090.8, 102396.2, 
    101992.4,
  103682.3, 103712, 103710, 103642.3, 103506.5, 103139.9, 103181.1, 102991.7, 
    103079.5, 103255.6, 103321, 103340.8, 103219.6, 101068.7, 101524.1,
  103644.2, 103691.7, 103655.3, 103633.1, 103319.6, 99728.31, 102899.8, 
    103035, 103040.6, 103144.7, 103195.4, 103273.6, 103218.6, 103090.1, 
    102804.6,
  103573.9, 103640.2, 103619.2, 103547.4, 103370.8, 102987.4, 99118.8, 
    102555.6, 102809.9, 103029.5, 103122.8, 103173.8, 103185.8, 103106.2, 
    102877.3,
  103513.3, 103552.7, 103543.9, 103437.6, 103293.9, 103086.4, 102750.3, 
    96701.6, 95944.53, 102588.6, 103034.4, 103072.9, 103161.3, 103041.9, 
    102940.3,
  103387.8, 103430.3, 103411.6, 103314.6, 103159.2, 102981.5, 102832, 
    102667.7, 102486.6, 102718.6, 102936.7, 103003.1, 103087.7, 103043.7, 
    102954,
  103264.2, 103272.7, 103251.7, 103184, 103075.9, 102910, 102776, 102719.6, 
    102696.5, 102694.8, 102843.9, 102935.3, 103014.7, 103008.5, 102938.1,
  103159.8, 103164.5, 103129.8, 103075.7, 102949, 102824, 102734.8, 102642.3, 
    102599.9, 102634.2, 102747.8, 102828.7, 102919.9, 102970.9, 102948.1,
  102982.8, 103004.7, 102983.2, 102933.7, 102844.1, 102756.7, 102684.7, 
    102636.5, 102596, 102556.3, 102611.3, 102710.9, 102812, 102902.2, 102917.1,
  102779.7, 102806.9, 102811.4, 102774.9, 102710.6, 102667.4, 102616.8, 
    102538.2, 102465.5, 102393, 102421.4, 102518.9, 102655.2, 102803.4, 
    102888.8,
  103850.7, 103922.2, 103945, 103866.1, 103721.8, 103484.5, 103159, 102961, 
    102820, 102364.8, 102300.2, 102417, 102131.7, 101470.8, 101123.1,
  103761.4, 103818.7, 103821.1, 103762.3, 103602.6, 103182.4, 103154.2, 
    102846.6, 102669, 102581.1, 102460, 102354.2, 102202, 100118.3, 100586.6,
  103611, 103697.4, 103676.1, 103636.2, 103357, 99744.48, 102868.9, 102980.2, 
    102767.2, 102547.7, 102381.8, 102282.2, 102166.2, 102032.8, 101793.8,
  103471.1, 103551.7, 103540.2, 103494.5, 103359.4, 102966.5, 99122.48, 
    102479, 102518.3, 102465.8, 102325.5, 102212.4, 102126.5, 102024.5, 
    101824.5,
  103304.1, 103370.8, 103381.1, 103323.9, 103223.2, 103059.5, 102734.2, 
    96655.23, 95815.66, 102152.5, 102275.1, 102138, 102082.5, 101972.8, 101863,
  103186.8, 103196.8, 103186.5, 103145.9, 103029.4, 102910.6, 102781.3, 
    102548.8, 102258.8, 102306.6, 102201, 102092.4, 102028.9, 101979.7, 
    101877.3,
  103065.5, 103058.1, 103020.6, 102963.5, 102885.4, 102774.5, 102633, 
    102529.4, 102394.2, 102225.6, 102109.2, 102024, 101949.4, 101964.6, 
    101887.7,
  102899.4, 102887, 102843.8, 102789.6, 102692.6, 102591.6, 102471.1, 
    102322.6, 102190.7, 102117.8, 102034.2, 101947.4, 101896.1, 101960.3, 
    101919.1,
  102665, 102667.7, 102618.9, 102557.4, 102480.6, 102387.2, 102275, 102199.5, 
    102098, 102005.3, 101940.5, 101873.5, 101824.6, 101929.2, 101933.4,
  102439, 102414.5, 102363.7, 102319, 102221.5, 102131.5, 102047.4, 101937.6, 
    101851.2, 101802.7, 101825.8, 101796.8, 101748.6, 101871, 101948.7,
  103578, 103660.5, 103739.6, 103742.9, 103727.9, 103637.3, 103451.9, 
    103270.8, 103044.5, 102409.8, 102196.2, 102185.8, 101810.9, 101260, 
    101212.9,
  103410, 103469.4, 103497.3, 103520.2, 103476.2, 103196.3, 103248.1, 
    102957.9, 102701.2, 102527.6, 102277.2, 102070.6, 101847.4, 99876.09, 
    100667.2,
  103163.8, 103233.8, 103247, 103246.9, 103068.1, 99528.12, 102717.8, 
    102875.6, 102595.6, 102338.1, 102100.8, 101920.8, 101728.9, 101687.9, 
    101859.7,
  102995.6, 103009.6, 102994.9, 102967.5, 102880.3, 102580.7, 98790.79, 
    102115.5, 102199.1, 102121.6, 101916.1, 101736.7, 101597.4, 101629.8, 
    101865.2,
  102837.5, 102814.6, 102787.6, 102712, 102628.6, 102496.6, 102190.7, 
    96162.55, 95272.59, 101579.6, 101718.1, 101532.7, 101441.9, 101479.7, 
    101788.3,
  102700.6, 102631.6, 102534.3, 102447.4, 102292.1, 102167.8, 102015.9, 
    101786.2, 101504.5, 101572.2, 101431.8, 101315.4, 101263, 101370.3, 101702,
  102509.5, 102433.1, 102305.2, 102170.5, 102009.4, 101829.9, 101648, 
    101520.8, 101361.9, 101206.7, 101110.6, 101059.4, 101047.6, 101237.5, 
    101609.1,
  102236.6, 102120.9, 101948.7, 101806, 101605.6, 101441.3, 101257.8, 
    101090.3, 100956.8, 100895.3, 100810.7, 100780.4, 100829, 101118.3, 
    101554.8,
  101912.5, 101812.4, 101654.8, 101491.7, 101303.5, 101112.5, 100923.6, 
    100845.5, 100717.8, 100609.7, 100534, 100535.8, 100618.9, 100995.6, 
    101476.5,
  101637.6, 101507.8, 101337.9, 101179.7, 100958.2, 100781.1, 100683.8, 
    100545.3, 100411, 100319.2, 100292.6, 100331.5, 100462.9, 100908.6, 
    101415.1,
  102847.8, 102916.6, 103006.2, 103051.1, 103109, 103112.5, 103058, 103004.1, 
    102892.3, 102350, 102176.8, 102175.1, 101782.4, 101161.2, 101008.5,
  102585.7, 102635.2, 102695.9, 102764.6, 102801.4, 102633.8, 102764.6, 
    102583.7, 102388.9, 102237, 102024.1, 101783.1, 101554.3, 99559.16, 
    100260.8,
  102210.7, 102262, 102341.5, 102399, 102328.9, 98893.01, 102172.4, 102387.1, 
    102179.1, 101869.7, 101601.5, 101381.8, 101199.6, 101124.2, 101294.5,
  101823.5, 101876.3, 101955.7, 102013.6, 102064.1, 101860.8, 98167.88, 
    101526.4, 101557.7, 101445.4, 101200.8, 101001.3, 100939.9, 100893.4, 
    101240,
  101378.9, 101467, 101562.3, 101638.6, 101700.9, 101714.6, 101522.7, 
    95573.28, 94636.77, 100800.7, 100919.8, 100760.4, 100723.2, 100690.5, 
    101176.1,
  100899.3, 101005.1, 101120, 101229.7, 101281, 101314, 101290.1, 101093, 
    100812.2, 100830, 100703.8, 100611.6, 100542, 100568.9, 101138.2,
  100388.6, 100498.4, 100633.3, 100785.9, 100875.6, 100924.7, 100903.7, 
    100876.5, 100738.9, 100633.4, 100562, 100500.1, 100389.1, 100522.6, 
    101184.6,
  99937.68, 100002.3, 100107.4, 100288.8, 100416.1, 100530.6, 100562.6, 
    100536.2, 100510.7, 100524.3, 100451.6, 100395.6, 100302.9, 100555.5, 
    101280.5,
  99521, 99553.77, 99653.82, 99838.8, 100026, 100183.8, 100257.7, 100345, 
    100360.7, 100367.9, 100322.6, 100304.7, 100293.4, 100705, 101445.3,
  99159.09, 99145.91, 99225.46, 99405.06, 99610.88, 99815.99, 99961.91, 
    100072.9, 100139.4, 100192, 100211.7, 100238.7, 100385.2, 100887.5, 
    101531.2,
  101439, 101570.2, 101780.2, 101971.7, 102200.2, 102383.5, 102505.1, 
    102630.7, 102716.7, 102375.4, 102368.1, 102500.4, 102166.4, 101453.8, 
    101031.1,
  101009.8, 101121.1, 101338.1, 101556.3, 101790.4, 101819.7, 102145.5, 
    102239.5, 102279.7, 102376.3, 102340.3, 102268.2, 102086.3, 99959.77, 
    100411.9,
  100415.8, 100615, 100850.4, 101088.2, 101263.8, 98015.41, 101456.6, 101996, 
    102014.7, 102019.1, 102011.9, 101957.7, 101838.8, 101683.9, 101660.2,
  99899.41, 100091.8, 100348.1, 100562.3, 100857.6, 100838.2, 97445.66, 
    101082.9, 101554.3, 101674.7, 101719.2, 101654.8, 101637.5, 101596.4, 
    101768.8,
  99486.94, 99661.64, 99855.02, 100083.7, 100304, 100617.5, 100653.6, 
    95021.98, 94279.92, 100894.5, 101392.5, 101369.6, 101442.8, 101479.4, 
    101792.8,
  99209.64, 99340.76, 99456.8, 99612.22, 99773.03, 99978.74, 100307, 
    100392.1, 100480.7, 100973.4, 101087.4, 101164.3, 101290.8, 101478.1, 
    101820.4,
  99081.93, 99151.56, 99174.73, 99222.6, 99319.52, 99464.31, 99687.24, 
    100045.1, 100355.3, 100609.2, 100821.1, 100990.4, 101179.6, 101497.7, 
    101859.1,
  99044.73, 99041.7, 98965.03, 98921.07, 98897.24, 98987.54, 99165.36, 
    99420.09, 99776.75, 100228.3, 100567.5, 100812.9, 101110.1, 101524.9, 
    101933.4,
  99084.45, 99020.41, 98872.49, 98733.05, 98611.27, 98592.38, 98715.34, 
    99009.27, 99376.88, 99829.11, 100269, 100626.4, 101034.1, 101545.8, 
    102013.5,
  99155.59, 99023.45, 98821.36, 98615.36, 98383.07, 98233.92, 98291.94, 
    98545.89, 98946.53, 99429.63, 99992.58, 100451.9, 100974.4, 101566.5, 
    102042.4,
  100051.4, 100376.4, 100805, 101163.6, 101573, 101945.2, 102247.2, 102563.7, 
    102853.9, 102717.1, 102919.5, 103278.9, 103161.9, 102677.9, 102448.5,
  99718.92, 100030.5, 100450.2, 100887, 101298.4, 101520.8, 102021.4, 
    102304.3, 102547.7, 102824.5, 102995.9, 103141.2, 103197.1, 101246.6, 
    101879.8,
  99350.23, 99677.2, 100113.2, 100588.2, 100937.4, 97823.4, 101538.4, 
    102187.2, 102397.7, 102574.9, 102734.5, 102913.4, 103023, 103086, 103103.5,
  99003.02, 99361.84, 99783.64, 100203.3, 100759.2, 100806.7, 97564.94, 
    101471.6, 102040.7, 102296.2, 102512.6, 102642.6, 102847.8, 102956, 
    103104.6,
  98789.85, 99102.15, 99536.95, 99964.09, 100465.7, 100933.4, 100974, 
    95346.34, 94789.91, 101529.1, 102205.8, 102323.5, 102605.7, 102757.2, 
    103014.7,
  98935.91, 99001, 99365.5, 99755.54, 100178.6, 100542.8, 100934.9, 100989.6, 
    101080, 101624.1, 101836.5, 102025.1, 102331.9, 102591, 102887.4,
  99204.07, 99187.12, 99379.93, 99671.82, 100045.5, 100346.7, 100607, 
    100929.3, 101174.8, 101329.5, 101525.5, 101774.5, 102079.3, 102413.7, 
    102782.8,
  99509.89, 99439.94, 99465.11, 99625.92, 99851.39, 100082, 100305.4, 
    100501.3, 100712.3, 101030.2, 101312.6, 101571.1, 101901.1, 102273.6, 
    102715.6,
  99940.8, 99824.79, 99769.68, 99804.75, 99891.66, 99964.66, 100034.5, 
    100203.7, 100419.6, 100697.1, 101027.4, 101365.5, 101728, 102160.7, 
    102662.6,
  100269.6, 100209.4, 100156.8, 100110.3, 100051.9, 100015.1, 99939.05, 
    99921.28, 100035.3, 100290.9, 100721.6, 101144.9, 101577.2, 102072.1, 
    102617.6,
  100310, 100662.6, 101071.4, 101431.7, 101889.8, 102316.1, 102692.9, 103118, 
    103484, 103368.4, 103602.9, 103983.3, 103875.1, 103437.7, 103286.7,
  100216.8, 100543.1, 100960.1, 101376.5, 101801.1, 102091.8, 102644.6, 
    103045, 103354.2, 103676.9, 103868.8, 104023.3, 104071, 102105.2, 102885.7,
  100085.9, 100434.7, 100850.6, 101315.3, 101623.5, 98542.49, 102438, 
    103069.9, 103401.9, 103618.8, 103829.4, 103995.6, 104119.2, 104179, 
    104221.6,
  99955.05, 100305.7, 100724.8, 101157.8, 101673, 101697, 98547.7, 102614.4, 
    103231.8, 103551.2, 103789.9, 103923.3, 104099.4, 104200.8, 104338.6,
  99864.38, 100209.1, 100609.8, 101047.1, 101505.2, 101979.6, 102036.9, 
    96488.73, 96077.12, 103088.2, 103694.7, 103823.6, 104039.4, 104123.6, 
    104310.9,
  99818.57, 100149.1, 100507.1, 100926.9, 101348.3, 101723.1, 102188.7, 
    102315.8, 102483.6, 103191.6, 103484.7, 103695.4, 103910.6, 104069.9, 
    104230.9,
  99830.46, 100097.9, 100445.6, 100812, 101237.3, 101592.5, 101934.3, 
    102386.3, 102746.8, 102993.5, 103258.9, 103519.1, 103740.3, 103950.7, 
    104126.9,
  99929.55, 100148.7, 100411, 100738.5, 101094, 101438.7, 101773.8, 102030.6, 
    102317.2, 102716.9, 103048, 103305.9, 103562.9, 103810.6, 104041.6,
  100119.1, 100236.7, 100424.7, 100693.3, 101002.2, 101297.8, 101591.4, 
    101927.6, 102220.1, 102533.3, 102826.9, 103114.4, 103382.5, 103658.8, 
    103932.5,
  100479.5, 100498.7, 100561.3, 100717.5, 100937.2, 101169.8, 101421.1, 
    101667.2, 101928.8, 102240.8, 102621.5, 102933.8, 103210.4, 103520.3, 
    103828.2,
  101502.2, 101848.5, 102254.5, 102630, 103035.1, 103359.7, 103617, 103895.8, 
    104085.6, 103859.8, 104010.9, 104353.4, 104191.8, 103703.8, 103488.8,
  101566.2, 101913.7, 102323.6, 102744.7, 103108.2, 103290.6, 103770.8, 
    103991.5, 104114.3, 104319, 104402.6, 104518.9, 104464.7, 102487.6, 
    103145.1,
  101585, 101988.2, 102397.5, 102853, 103035.5, 99891.08, 103729.8, 104198.6, 
    104376, 104464.8, 104541.4, 104653.8, 104694.2, 104682.1, 104587.1,
  101578.2, 101991, 102413.4, 102826.7, 103266.7, 103224.9, 99947.38, 
    103938.1, 104348.8, 104548.2, 104686.1, 104748.1, 104826.2, 104854.1, 
    104803.3,
  101572, 101986.9, 102408.9, 102824.5, 103226.6, 103669, 103646.7, 97775.12, 
    97329.95, 104400.5, 104802.9, 104834.8, 104932, 104908.2, 104942.6,
  101542.3, 101956.3, 102354.2, 102784.4, 103158.5, 103534.2, 103930, 
    104020.7, 104080.9, 104655.6, 104798.4, 104898.4, 104986.6, 105006.5, 
    105012.2,
  101525.7, 101934.8, 102337.2, 102747.5, 103138.6, 103507, 103802.2, 
    104182.6, 104476.1, 104659.1, 104798.9, 104945.1, 105007.1, 105042.5, 
    105026.4,
  101487.9, 101882.1, 102273.1, 102676.6, 103053.7, 103427.8, 103755.4, 
    103998.7, 104258.7, 104585.4, 104788.9, 104929.9, 105018.7, 105074.9, 
    105076.2,
  101479.9, 101873, 102269.2, 102662.5, 103022.5, 103367.7, 103681.5, 
    104001.6, 104271.5, 104537.6, 104735, 104896.7, 104991.9, 105060.9, 
    105071.1,
  101458.7, 101828.3, 102209.9, 102596.4, 102966.2, 103308.4, 103600.5, 
    103847.5, 104094.2, 104375.4, 104627.1, 104812.4, 104932.2, 105024.4, 
    105064.6,
  102520, 102833.7, 103196.6, 103515.4, 103847.8, 104070.7, 104196.1, 
    104308.4, 104335.9, 103953.8, 103960, 104164.4, 103934.9, 103392.1, 
    103177.5,
  102579.6, 102911.9, 103293.3, 103683.1, 103958.1, 104018.9, 104382.2, 
    104432, 104417.4, 104467.6, 104407.2, 104390, 104232.7, 102197.6, 102829.1,
  102644.1, 103049.7, 103429.3, 103849.1, 103908.6, 100626.4, 104347.6, 
    104707.2, 104745.1, 104684.1, 104624.7, 104580, 104502.1, 104401.5, 104253,
  102726.3, 103143.5, 103540, 103885.2, 104227.3, 104057.8, 100618.7, 
    104482.9, 104760.2, 104854.3, 104840.9, 104739.7, 104680.3, 104580.6, 
    104473.7,
  102843.4, 103247.5, 103627.5, 103949.3, 104254.4, 104609.2, 104429.5, 
    98353.45, 97830.88, 104796.9, 105038.2, 104908.4, 104866.6, 104704.5, 
    104658,
  102971.6, 103347.6, 103692.2, 104018.1, 104268.7, 104523.5, 104832.8, 
    104808.3, 104783.9, 105152.8, 105155.3, 105088.6, 105008.7, 104888, 
    104777.6,
  103098.8, 103455.5, 103787.4, 104090.8, 104378.5, 104607.6, 104786.9, 
    105077.7, 105258.1, 105279.6, 105298.4, 105255.4, 105154.9, 105037.6, 
    104904.1,
  103208, 103547.4, 103876, 104159.4, 104413.6, 104660.9, 104887.4, 105060.2, 
    105220.4, 105392.9, 105436.5, 105390.3, 105302.6, 105178.4, 105039.2,
  103336.1, 103676.4, 103994.7, 104271.1, 104526.4, 104753.7, 104968.6, 
    105205.6, 105405.8, 105512, 105527, 105499, 105413.3, 105300, 105149.6,
  103428.5, 103754.7, 104066.8, 104344.8, 104599.7, 104829.8, 105040, 
    105219.1, 105397.1, 105496.1, 105567.5, 105552, 105487.3, 105399.2, 
    105272.7,
  103579.6, 103805.6, 103984.6, 104082.4, 104167.7, 104186.6, 104148.4, 
    104173, 104173.3, 103840.1, 103902.2, 104202.2, 104038, 103550.3, 103357.8,
  103589.4, 103834.7, 104034.6, 104228.9, 104294.6, 104122.5, 104324.5, 
    104250.2, 104179.7, 104219.6, 104215.9, 104249.4, 104193.2, 102169.8, 
    102828.2,
  103581.3, 103897.8, 104108.7, 104352.1, 104213.6, 100742.2, 104286.6, 
    104504.3, 104473.8, 104365, 104304.9, 104290.3, 104264.1, 104200.8, 
    104097.5,
  103567.4, 103898.6, 104152.3, 104349.2, 104521.3, 104236, 100583.1, 
    104293.4, 104407.7, 104473.2, 104415.1, 104330.7, 104287.9, 104219.8, 
    104164.4,
  103579.2, 103920.6, 104201.8, 104386.9, 104526.6, 104688.9, 104421.6, 
    98171.65, 97631.75, 104391, 104577.1, 104423.9, 104393.8, 104266.1, 104273,
  103578.1, 103942.9, 104224.9, 104466.9, 104600.1, 104713.8, 104865.5, 
    104792.4, 104592.3, 104769.8, 104701.1, 104582.4, 104506.2, 104417.3, 
    104376,
  103598.5, 103992.2, 104298, 104543.6, 104733.8, 104860.1, 104916.5, 105033, 
    105075.9, 104992.8, 104889.4, 104792.7, 104691.6, 104610.7, 104546,
  103619.7, 104012, 104342.9, 104621.4, 104821.8, 105010.9, 105141.1, 
    105187.7, 105198, 105191, 105105.6, 105001.8, 104904.2, 104820.5, 104761.8,
  103678.2, 104077.8, 104436.3, 104723.4, 104963.1, 105139.6, 105283.8, 
    105400.5, 105447.3, 105400.5, 105319.8, 105232.6, 105129, 105033.3, 
    104951.6,
  103719.6, 104117, 104479, 104790.8, 105054.5, 105278.2, 105453.6, 105541.5, 
    105552.9, 105496.2, 105484.5, 105445, 105354, 105266.1, 105177.4,
  103949.9, 103989.2, 104068, 104105.7, 104204.5, 104284.5, 104352, 104455.6, 
    104533.5, 104224.3, 104300.5, 104589.8, 104377.2, 103878.5, 103658.4,
  103965, 104031.6, 104107.9, 104210.8, 104279.3, 104162, 104412.7, 104456.3, 
    104469.5, 104594.8, 104642.2, 104713.6, 104647.5, 102654.5, 103339,
  103949, 104078.2, 104128.7, 104286.7, 104145.7, 100627.5, 104256.4, 
    104536.9, 104609.1, 104624, 104672.7, 104742.6, 104786.4, 104763.5, 
    104716.9,
  103943, 104051.6, 104116.1, 104212.2, 104319.2, 104084.4, 100378.4, 
    104205.9, 104458.3, 104589.2, 104700.1, 104743.1, 104820.8, 104861.1, 
    104897.9,
  103973.8, 104051.9, 104099.8, 104143, 104198.3, 104341.2, 104177.1, 
    98011.18, 97421, 104347.3, 104711.7, 104731.3, 104837.4, 104835.8, 104958,
  103995.7, 104088.3, 104123.5, 104184.2, 104215.6, 104271.4, 104390.3, 
    104386.8, 104217.2, 104589.1, 104680.1, 104746.9, 104851.3, 104922.5, 
    105009.4,
  104038.2, 104163.4, 104235.6, 104310.3, 104354.6, 104399.3, 104424.9, 
    104542.1, 104646, 104674.9, 104742.5, 104834.1, 104912, 105001.6, 105071.7,
  104092.9, 104262.7, 104374.6, 104475.4, 104525.1, 104581.7, 104633.2, 
    104663.9, 104715.8, 104801.1, 104871.9, 104945.1, 105030.1, 105111.1, 
    105176.6,
  104179, 104385.7, 104551.6, 104684.5, 104767.2, 104818.3, 104861.7, 
    104941.5, 105003.6, 105027, 105064.3, 105120.5, 105188, 105259.5, 105314.8,
  104256.7, 104508.1, 104719, 104882.8, 104988.9, 105073.3, 105123.5, 
    105144.6, 105173.8, 105188, 105279.2, 105341.9, 105391.5, 105453.1, 
    105494.2,
  104110.3, 104189.1, 104300.8, 104350.7, 104441.5, 104455.3, 104384.8, 
    104382.8, 104380.2, 104036.8, 104108.5, 104420.7, 104298.4, 103887.6, 
    103742,
  104097.1, 104197.3, 104316.3, 104440.4, 104514.7, 104327.9, 104516.9, 
    104452.4, 104405.4, 104484.7, 104496.2, 104587.3, 104547.5, 102665, 
    103408.4,
  104038.4, 104190.8, 104317, 104518, 104392.9, 100874.7, 104473.4, 104719.2, 
    104737.1, 104686.7, 104691.8, 104739.3, 104797.1, 104832.3, 104831.1,
  103977.8, 104135.8, 104292.4, 104440.2, 104639.6, 104338.4, 100717.7, 
    104497.2, 104734.6, 104840.5, 104900.2, 104893, 104966.5, 105036.7, 
    105094.2,
  103934.8, 104067.4, 104236.9, 104398.4, 104523.5, 104750.1, 104521.6, 
    98358.59, 97833.09, 104775.3, 105094.7, 105060.5, 105150.4, 105154.8, 
    105301.3,
  103884.3, 104023.7, 104146.5, 104328.1, 104441.2, 104602.5, 104844.9, 
    104782, 104654.7, 105103.7, 105180.2, 105223.4, 105299.1, 105358.6, 
    105455.6,
  103844.2, 103946.1, 104088.8, 104256.9, 104421.3, 104596.7, 104712.3, 
    104948.4, 105137.3, 105206.3, 105292.5, 105385.9, 105463.9, 105547.2, 
    105629.6,
  103802.3, 103929, 104062.8, 104223, 104360.1, 104561.8, 104754.4, 104878.2, 
    105061.9, 105271.6, 105411, 105514.6, 105621.7, 105733.9, 105843.9,
  103833.6, 103961.3, 104087.8, 104245.6, 104406.6, 104582.7, 104759, 
    105014.4, 105259.9, 105388.8, 105503.6, 105629.2, 105763.1, 105893.2, 
    106001.6,
  103926.5, 104062.5, 104190, 104318.6, 104451.2, 104636.7, 104839.8, 
    105028.7, 105238.4, 105381.5, 105573.9, 105738, 105890, 106034.8, 106152.1,
  104294.9, 104329.4, 104400.2, 104405, 104450.1, 104438.5, 104414.9, 
    104505.4, 104593.5, 104254.6, 104315.1, 104633.3, 104513.4, 104073.2, 
    103940.7,
  104232.1, 104270.6, 104318.2, 104375.2, 104373.5, 104212.9, 104428.9, 
    104479.4, 104512.1, 104622.4, 104690, 104801.8, 104817.8, 102923.1, 
    103732.6,
  104090.5, 104173, 104221.8, 104306.3, 104202.5, 100637.8, 104299.9, 
    104612.5, 104735.1, 104733.3, 104805.2, 104930.3, 105083, 105191.6, 
    105277.6,
  103969.5, 104031.9, 104099.8, 104133.9, 104293.5, 104066.3, 100469.8, 
    104305.8, 104643.2, 104799.1, 104969.8, 105073.9, 105293.2, 105496.8, 
    105607.8,
  103863.7, 103929.7, 103987.4, 104033.4, 104111.2, 104386.5, 104210.7, 
    98200.62, 97637.49, 104683.2, 105112.7, 105229.8, 105464.2, 105613, 
    105868.1,
  103793.5, 103885.4, 103918.1, 103967.9, 104042, 104212.3, 104492.2, 
    104453.7, 104387.4, 104950.2, 105162.8, 105365, 105594.8, 105788.4, 
    106003.1,
  103739.6, 103843.2, 103913.1, 103960.3, 104079.8, 104216.8, 104364.1, 
    104639.8, 104860.3, 104986.4, 105217.1, 105465.2, 105685.6, 105892.1, 
    106089.3,
  103691.9, 103822, 103928.8, 103989, 104080.4, 104235.7, 104405.3, 104497.3, 
    104717.8, 104997.5, 105276.5, 105517.6, 105763.8, 105981.1, 106187,
  103653.6, 103808.7, 103961.1, 104068.3, 104188, 104286.2, 104438, 104663.4, 
    104913.7, 105095.9, 105321.2, 105562.8, 105808.6, 106034.9, 106230.3,
  103595.8, 103761.8, 103948.5, 104085.9, 104209.4, 104345.8, 104500.2, 
    104654.2, 104874.6, 105059.3, 105334.1, 105581, 105827.7, 106061.4, 
    106247.9,
  104194.1, 104193, 104216.1, 104159.8, 104143.8, 104062.5, 103984.3, 
    104010.6, 104104, 103866.9, 104049.9, 104475.4, 104441.9, 104125.3, 
    104046.6,
  104126.5, 104135.1, 104141.6, 104145.3, 104136.7, 103902.1, 104078.3, 
    104011.8, 104048.1, 104220.5, 104360.2, 104559.2, 104672.5, 102833.2, 
    103675.4,
  103951.9, 104016.1, 104039.3, 104080.9, 103981.5, 100365.4, 103975.3, 
    104186.5, 104226.7, 104289.2, 104417.2, 104608, 104807.6, 104946.2, 
    105090.8,
  103772.9, 103840.2, 103884.4, 103904.3, 104001.3, 103840.4, 100079.2, 
    103940.4, 104194.1, 104348, 104534.4, 104696.8, 104928, 105171.7, 105349.2,
  103601.6, 103661.6, 103717.9, 103748.5, 103789.4, 103960.3, 103930.2, 
    97681.84, 97153.17, 104242.9, 104677.8, 104803.9, 105059.2, 105225.4, 
    105521.2,
  103434.7, 103483.6, 103535, 103592, 103639, 103764.7, 103994.6, 104066.6, 
    103964.5, 104498.3, 104721.9, 104913.6, 105160.1, 105370.5, 105600.3,
  103262.3, 103320.9, 103354.1, 103430.7, 103504.2, 103645.6, 103814, 
    104073.9, 104326.3, 104533.5, 104739.5, 104995.4, 105212.7, 105436.8, 
    105637.4,
  103092.7, 103157.1, 103195.9, 103272.7, 103349.1, 103502, 103724, 103928.4, 
    104181.5, 104480.6, 104753.7, 105017.8, 105253.7, 105487.5, 105693,
  102968.2, 103036.9, 103066.4, 103147.7, 103243.7, 103394.6, 103589.3, 
    103852.7, 104182.8, 104479.1, 104731.4, 105000.4, 105241.6, 105479.9, 
    105676.2,
  102858.8, 102942.8, 103014.6, 103087.8, 103171.1, 103314.9, 103504.9, 
    103731, 104061.2, 104344, 104650, 104925.1, 105175.3, 105423.9, 105623.6,
  103912.8, 103979, 104032.9, 104000.4, 104040.5, 104050.6, 104110.6, 
    104266.7, 104438.5, 104214.1, 104407.3, 104797, 104724.3, 104351.5, 
    104248.5,
  103768.6, 103862.5, 103937.1, 103956.1, 104035.6, 103887.5, 104148.2, 
    104219.9, 104364.4, 104535.9, 104686.6, 104835.7, 104914.7, 102987.6, 
    103780.7,
  103517.5, 103684, 103786.7, 103876.4, 103802.2, 100286.7, 103965.6, 
    104279.6, 104417, 104526.6, 104665.8, 104802.8, 104945.3, 105017, 105105.6,
  103221.5, 103449.2, 103573, 103680.9, 103749, 103670.4, 99929.32, 103912.7, 
    104279.3, 104448, 104626.1, 104749.1, 104919.8, 105078, 105221.3,
  102944.3, 103199.5, 103359.2, 103486.4, 103511.1, 103557.7, 103685.8, 
    97488.48, 96953.84, 104052.9, 104568.1, 104672.1, 104892.4, 104988.9, 
    105207.1,
  102663.5, 102939.1, 103118.9, 103285.9, 103356.1, 103362.5, 103535.2, 
    103762.6, 103649.2, 104132, 104384.8, 104570.7, 104797.6, 104965.2, 
    105149.7,
  102396.7, 102690.6, 102899.8, 103089.2, 103182.5, 103242.5, 103276.5, 
    103511.9, 103771.3, 103966.3, 104189.8, 104460.3, 104672.6, 104868.8, 
    105048.4,
  102140, 102443, 102668.2, 102875.3, 102997.8, 103090, 103148.1, 103289.5, 
    103516.8, 103810.1, 104064.6, 104313.7, 104539.6, 104758.3, 104965,
  101937.5, 102252.5, 102490.7, 102685, 102811.5, 102917.4, 102981.8, 
    103120.4, 103358.8, 103653.4, 103912.5, 104162.1, 104395.4, 104614.8, 
    104823.3,
  101768.5, 102070.3, 102301.5, 102490.6, 102626.1, 102749.1, 102843, 
    102967.1, 103186.5, 103440.3, 103728.9, 103988.5, 104221.3, 104465.2, 
    104679.1,
  102734.3, 103001.9, 103336.5, 103571.8, 103788.9, 104000.9, 104198.1, 
    104363.7, 104542.6, 104289.1, 104414.6, 104748.9, 104622.9, 104214.9, 
    104082.2,
  102500.4, 102738.5, 103102.5, 103392.6, 103657.3, 103746.3, 104137.9, 
    104281.4, 104412.5, 104587.8, 104692.4, 104773.8, 104812.3, 102819.6, 
    103603.9,
  102180.8, 102478.7, 102873.9, 103224.5, 103400.3, 100047.3, 103896.9, 
    104345.1, 104484.3, 104540, 104644.2, 104739.2, 104814.1, 104874.2, 
    104921.9,
  101794.9, 102159.3, 102565.4, 102951.1, 103362.8, 103347.1, 99836.62, 
    103863.4, 104289, 104462.4, 104605.9, 104678.3, 104789.6, 104895.2, 
    105016.5,
  101417.4, 101816.2, 102260.1, 102696.1, 103093.6, 103493.2, 103519.3, 
    97517.63, 96924.37, 103965.9, 104522.1, 104585.4, 104751.5, 104809.6, 
    104996.6,
  101096.1, 101481.8, 101922.2, 102411, 102815, 103161.6, 103514.7, 103609.3, 
    103587.8, 104047.6, 104295.8, 104453.8, 104647.2, 104773.6, 104913.3,
  100800.1, 101186.8, 101652.1, 102153.1, 102590.5, 102960.6, 103215.4, 
    103530.6, 103753.6, 103851.8, 104052.7, 104292.2, 104487.6, 104650.2, 
    104793.9,
  100559.8, 100916.1, 101363.3, 101886, 102326.2, 102724.9, 103015.7, 
    103214.3, 103413.3, 103667.2, 103901.1, 104123.5, 104322.1, 104501.9, 
    104662.8,
  100371, 100727.1, 101185.7, 101692.6, 102144.2, 102536.4, 102838.9, 103078, 
    103281.4, 103468.9, 103689, 103928.4, 104125.5, 104305.7, 104473.7,
  100232.7, 100547, 100980.8, 101491.9, 101941.3, 102338.1, 102656.9, 
    102888.1, 103065.1, 103234.8, 103462.5, 103691.6, 103900.9, 104101.8, 
    104274.6,
  101503.2, 101603.3, 101849.8, 102216.1, 102590.6, 102933.8, 103184.5, 
    103414.2, 103600, 103368.5, 103510.3, 103918, 103841.4, 103493.1, 103397.1,
  101253.6, 101377, 101634.6, 102044.5, 102420, 102641.5, 103096.7, 103311.8, 
    103446.7, 103676.7, 103784.4, 103944.4, 104023.6, 102092.4, 102897.7,
  100952.2, 101110.3, 101445.9, 101893.4, 102159.4, 98942.05, 102848.1, 
    103382.3, 103561.3, 103648, 103766.6, 103907.1, 104054, 104144.5, 104219.9,
  100683.5, 100811.7, 101205.6, 101645, 102135.4, 102150.4, 98834.71, 
    102884.3, 103372.3, 103589.7, 103758.5, 103858.8, 104025.8, 104173.9, 
    104322.5,
  100441.9, 100553.7, 100934.4, 101414.1, 101895, 102380.7, 102402, 96631.14, 
    96084.91, 103193.6, 103729.2, 103808, 104010.6, 104092.8, 104312.7,
  100256.3, 100338.7, 100662.1, 101157, 101607.8, 102062.7, 102523.1, 
    102620.3, 102694.1, 103329.9, 103579.9, 103746.9, 103944.3, 104089.5, 
    104266.8,
  100080.4, 100149.3, 100435.1, 100932.9, 101415.5, 101865, 102244.6, 
    102736.5, 103058.2, 103206.3, 103414.6, 103658, 103857.4, 104032.1, 
    104189.1,
  99960.6, 100014.7, 100239.1, 100725.3, 101176.4, 101653.4, 102051.6, 
    102394.2, 102706, 103040.9, 103323.9, 103558.3, 103766.2, 103958.1, 104128,
  99898.88, 99932.29, 100118.2, 100598.5, 101043.9, 101496.9, 101890.6, 
    102304.1, 102674.3, 102954.5, 103207.3, 103447.1, 103655, 103848.7, 
    104015.9,
  99910.28, 99907.87, 100049.7, 100465, 100906.4, 101347.9, 101734.3, 
    102096.4, 102481.1, 102783, 103072.4, 103309, 103520.9, 103721, 103891.2,
  100708.2, 100602.6, 100582.7, 100736.4, 101048.5, 101380.9, 101650.2, 
    101935.6, 102214.6, 102091.9, 102315.5, 102773.4, 102722.2, 102404.4, 
    102329.7,
  100498.5, 100377.8, 100387.3, 100614.6, 100994.8, 101166.4, 101643.9, 
    101885.2, 102118.4, 102380.3, 102563.1, 102764.3, 102882.5, 100993.4, 
    101816,
  100281.4, 100156.8, 100214.8, 100511.7, 100788.2, 97609.75, 101480, 
    101991.9, 102212.7, 102375, 102534.6, 102722.8, 102894.8, 103018.6, 
    103121.8,
  100054.8, 99954.93, 100016.3, 100344, 100781.4, 100817.4, 97509.61, 
    101590.4, 102075, 102323.6, 102523.6, 102678, 102883, 103074.6, 103236.2,
  99815.18, 99772.21, 99807.21, 100165.5, 100593.6, 101025, 101074.1, 
    95346.08, 94840.7, 101988.2, 102517.6, 102646.8, 102869.9, 102997.5, 
    103232,
  99610.56, 99603.66, 99616.02, 99961.7, 100391, 100799.5, 101230.6, 
    101386.2, 101484.9, 102145.9, 102414.4, 102618.2, 102842.6, 103015.9, 
    103204.4,
  99450.7, 99469.38, 99463.06, 99773.45, 100237.2, 100659.1, 101046.7, 
    101517.8, 101851.6, 102062.7, 102313.4, 102583.3, 102795.2, 102990.5, 
    103157.6,
  99395.54, 99411.27, 99371.24, 99637.97, 100099.2, 100525.9, 100922.3, 
    101294.8, 101606.8, 101974, 102279.2, 102547.4, 102771.7, 102974.5, 
    103144.8,
  99383.8, 99354.18, 99301.6, 99553.62, 100050.7, 100468.2, 100862.2, 101251, 
    101636.3, 101960.8, 102234.8, 102504, 102730, 102939.6, 103112.2,
  99393.2, 99303.12, 99248.07, 99551.05, 100044.3, 100416, 100789.4, 
    101172.6, 101562.2, 101872.7, 102190.2, 102462.1, 102685.1, 102904.5, 
    103085.8,
  99867.93, 99921.52, 100033, 100122.8, 100261.8, 100422.4, 100628.5, 
    100889.8, 101213, 101159.7, 101453.8, 101920.1, 101856.3, 101447.4, 
    101278.4,
  99530.75, 99604.08, 99758.73, 99896.12, 100078, 100189.9, 100629.3, 
    100838.5, 101104.2, 101444.4, 101679.4, 101910.7, 102023.9, 100094, 100830,
  99143.97, 99237.88, 99428.46, 99648.85, 99813.97, 96761.77, 100511.6, 
    101024.5, 101205.4, 101430.8, 101642.2, 101858.4, 102029.5, 102119.2, 
    102177.4,
  98808.94, 98907.12, 99084.11, 99342.16, 99732.41, 99824.95, 96621.56, 
    100617, 101123.7, 101386, 101612.1, 101802.9, 102020, 102199.5, 102310.8,
  98501.77, 98601.58, 98788.12, 99059.38, 99505.54, 99928.38, 99988.44, 
    94388.58, 93923.08, 101027.8, 101609.1, 101759.1, 102011.3, 102136.5, 
    102347.6,
  98271.64, 98344.7, 98528.79, 98821.31, 99270.46, 99745.88, 100104.7, 
    100245.7, 100371.3, 101140.2, 101480, 101719.4, 101989.8, 102168, 102359.3,
  98211.87, 98233.64, 98382.45, 98667.94, 99141.48, 99641.69, 99994.1, 
    100390.1, 100727.4, 101052.8, 101377.8, 101704.4, 101957.2, 102170.5, 
    102344.5,
  98238.72, 98270.78, 98379.96, 98662.52, 99121.3, 99581.28, 99965.95, 
    100281.1, 100627.2, 101061.7, 101396.5, 101709.5, 101962.7, 102191.5, 
    102368.1,
  98380.3, 98395.19, 98510.27, 98774.51, 99234.82, 99639.07, 100007.4, 
    100375.3, 100776.6, 101127.9, 101441.3, 101735.5, 101979.1, 102198.2, 
    102370.5,
  98529.79, 98565.74, 98696, 98975.49, 99396.82, 99741.23, 100118, 100482.3, 
    100884.9, 101173.6, 101496.9, 101772.8, 102002.9, 102216.9, 102388.3,
  99539.72, 99563.6, 99652.27, 99744.77, 99887.99, 100033.7, 100170.7, 
    100341.9, 100547.1, 100451.5, 100772.8, 101311.9, 101371.3, 101084, 
    100975.1,
  99192.59, 99231.55, 99344.41, 99476.48, 99615.67, 99649.31, 100004.4, 
    100147.8, 100354.2, 100672.8, 100947.8, 101255.6, 101475.2, 99612.24, 
    100346.3,
  98861.69, 98892.7, 99031.38, 99222.29, 99323.53, 96170.95, 99750.77, 
    100216.5, 100388.6, 100636.2, 100901.3, 101190.1, 101426.4, 101546, 
    101576.1,
  98632.57, 98647.28, 98751.74, 98979.59, 99284.66, 99303.27, 96047.91, 
    99871.64, 100347.7, 100632.4, 100882.5, 101143, 101403.6, 101574, 101585.7,
  98408.2, 98428.48, 98530.59, 98764, 99122.38, 99499.16, 99526.56, 93929.32, 
    93415.54, 100356.4, 100930.8, 101124.9, 101400.2, 101514.9, 101614.7,
  98243.81, 98240.07, 98337.62, 98622.98, 98997.47, 99369.77, 99711.02, 
    99796.13, 99860.33, 100527.7, 100845.3, 101117.7, 101397.8, 101542.3, 
    101625,
  98146.73, 98159.77, 98234.74, 98556.36, 98979.19, 99332.91, 99617.23, 
    99971.26, 100196.8, 100448, 100784.9, 101131.4, 101392.2, 101568.7, 101631,
  98135.73, 98160.47, 98258.97, 98648.59, 98993.9, 99351.94, 99622.72, 
    99847.86, 100099.2, 100489.8, 100830.3, 101171.8, 101423, 101617.9, 
    101685.6,
  98323.52, 98333.3, 98496.75, 98832.57, 99141.12, 99439.01, 99683.31, 
    99995.4, 100306.9, 100623.5, 100931.4, 101238.8, 101480.9, 101669.1, 
    101738.9,
  98837.12, 98790.72, 98896.74, 99129.02, 99335.96, 99590.23, 99867.42, 
    100188.4, 100480.3, 100741.7, 101036.6, 101334.9, 101550.5, 101735, 
    101802.9,
  100072.7, 100102.1, 100175.4, 100265, 100398.1, 100527.5, 100608.6, 
    100721.1, 100829.5, 100586.4, 100719.8, 101091.1, 101062, 100828.4, 
    100914.2,
  99716.95, 99748.09, 99827.89, 99948.54, 100047.7, 100038.4, 100345.2, 
    100441.4, 100525.6, 100686.2, 100782.5, 100959.3, 101114, 99403.55, 
    100300.6,
  99375.43, 99355.21, 99422.86, 99560.19, 99642.89, 96440.2, 99859.12, 
    100319.8, 100367.7, 100490.6, 100626.9, 100824.8, 101044.9, 101256.2, 
    101516.8,
  99163.98, 99083.56, 99081.81, 99159, 99401.87, 99413.68, 96072.98, 
    99757.03, 100218.6, 100366.2, 100536.3, 100726.1, 101024.2, 101313.6, 
    101601.3,
  99056.21, 98934.2, 98893.7, 98927.77, 99113.62, 99446.52, 99508.88, 
    93928.21, 93333.06, 100065.5, 100547.9, 100710.6, 101032.6, 101263.5, 
    101621.3,
  99074.99, 98894.2, 98787.45, 98804.73, 98950.43, 99298.72, 99643.61, 
    99713.31, 99764.02, 100299.2, 100497.7, 100750.5, 101077.7, 101332.1, 
    101646.5,
  99216.65, 99038.7, 98851.38, 98843.82, 99084.22, 99418.68, 99668.35, 
    99959.24, 100129.6, 100280.1, 100518, 100828.7, 101126, 101385.5, 101634.2,
  99431.89, 99355.08, 99294.89, 99303.16, 99439.83, 99608.22, 99789.32, 
    99928.11, 100141.5, 100396.1, 100634, 100932.5, 101203.3, 101459.1, 
    101659.9,
  99622.84, 99586.24, 99546.42, 99580.9, 99665.94, 99805.74, 99955.8, 
    100176.2, 100398, 100555.5, 100793.8, 101052.5, 101290.9, 101507.2, 
    101641.3,
  99842.53, 99783.9, 99789.88, 99823.65, 99888.9, 99995.59, 100152.4, 100348, 
    100529.3, 100681.1, 100918.6, 101162.5, 101371.3, 101542.8, 101617.4,
  100618, 100592.6, 100570.2, 100592.7, 100668.8, 100802, 100886.5, 101025.4, 
    101191.9, 101001.2, 101189.9, 101598.1, 101561.9, 101264.4, 101216.5,
  100424.9, 100341.9, 100267.1, 100274.3, 100319.1, 100325.6, 100638.8, 
    100767.3, 100889.2, 101100.8, 101244.5, 101413.2, 101521, 99742.28, 
    100507.3,
  100353.8, 100203.3, 100059.1, 99984.11, 99943.11, 96716.49, 100159.1, 
    100636.9, 100734.5, 100883.2, 101035.1, 101210.2, 101366.6, 101501, 
    101653.6,
  100344.2, 100150.6, 99951.65, 99779.59, 99776.74, 99749.21, 96335.45, 
    100038.8, 100509.7, 100692.5, 100870, 101018.8, 101226.4, 101434, 101641.3,
  100371.1, 100191.7, 99984.91, 99756.82, 99671.18, 99806.17, 99833.83, 
    94157.84, 93539.2, 100185.8, 100735.5, 100872.2, 101126.4, 101308.1, 
    101622.3,
  100415.8, 100271.8, 100055.6, 99877.48, 99692.65, 99742.94, 99968.38, 
    99954.07, 99906.52, 100287.4, 100529.7, 100769.2, 101057.5, 101312.8, 
    101630.9,
  100490.6, 100418.8, 100283.5, 100148.7, 100046.7, 99981.73, 100032.6, 
    100137.1, 100189.5, 100199.5, 100451.5, 100743.4, 101054.1, 101352.5, 
    101686.6,
  100532, 100514, 100436.1, 100356.5, 100262.9, 100230.7, 100229.5, 100212.5, 
    100234.2, 100327.6, 100536.6, 100814.6, 101129.7, 101459.9, 101803.6,
  100588.3, 100622.5, 100594.8, 100548.6, 100504.4, 100468, 100455.6, 
    100523.5, 100538, 100551.6, 100722.7, 100964.1, 101276.1, 101612.1, 
    101944.2,
  100657.7, 100701.4, 100720.4, 100701.3, 100664.2, 100647.8, 100667.3, 
    100707.8, 100733.6, 100772.3, 100937.6, 101171.4, 101453.1, 101774.2, 
    102069.3,
  101630.1, 101557.7, 101447.6, 101315.9, 101172.7, 101074.2, 101021.3, 
    101056.8, 101147, 100914.8, 101043.6, 101389.6, 101311.2, 101039.7, 
    101030.5,
  101605.5, 101530.5, 101412.4, 101269.6, 101082.7, 100780.6, 100929.3, 
    100906.1, 100954.1, 101113, 101203.4, 101319.6, 101400.7, 99610.41, 
    100412.6,
  101599.2, 101537.1, 101420.2, 101285.1, 100975.6, 97442.48, 100722.3, 
    100928.9, 100913.1, 100957, 101054.5, 101190.5, 101325.5, 101464.8, 
    101607.8,
  101591.6, 101549.3, 101444.2, 101287.9, 101140.2, 100797.6, 97075.26, 
    100604.5, 100845.2, 100888.1, 100953.9, 101060.9, 101231, 101436.8, 
    101620.8,
  101573.2, 101574.2, 101497.5, 101355, 101204.9, 101062.2, 100843.5, 
    94789.48, 94034.33, 100521.5, 100840, 100930.6, 101142.4, 101307.2, 
    101574.9,
  101550.9, 101565.1, 101493, 101380.1, 101220.8, 101100.8, 101027.1, 
    100891.1, 100661.9, 100713.9, 100718.3, 100835.2, 101066.9, 101276.4, 
    101534.1,
  101518.8, 101552.9, 101491.2, 101374.3, 101230.5, 101102.9, 101020.6, 
    101005.8, 100876.7, 100672.9, 100669.5, 100829.1, 101032.6, 101265.8, 
    101521.6,
  101500.6, 101511, 101414.9, 101300, 101161.7, 101054.7, 100990.6, 100963.4, 
    100880.9, 100766.9, 100731.5, 100868.3, 101067.1, 101315.7, 101585.7,
  101470.1, 101454.7, 101348.7, 101217.4, 101112, 101013.5, 100955.9, 
    101014.8, 100969.5, 100843.1, 100813.4, 100947.8, 101140.7, 101410.6, 
    101703.7,
  101421.3, 101317.2, 101183.9, 101101.1, 100997.2, 100925.5, 100918.4, 
    100967, 100959.1, 100876.3, 100897, 101045.2, 101254.9, 101545.3, 101805.4,
  102874.6, 102880.3, 102879, 102793, 102666.3, 102482.2, 102237, 102052.9, 
    101886, 101411, 101426.3, 101648.9, 101484.3, 101036.2, 100896.1,
  102843, 102844.2, 102794.3, 102675.2, 102489.9, 102075.2, 102090.3, 
    101777.3, 101586.7, 101539.5, 101499.9, 101516.8, 101497.7, 99578.39, 
    100236.1,
  102771.6, 102774.8, 102662.2, 102540.1, 102162.3, 98563.86, 101558.6, 
    101739, 101487.6, 101373.5, 101339.9, 101372.1, 101370.4, 101389.7, 
    101389.2,
  102675.9, 102633.7, 102503.1, 102295, 102032.6, 101557.7, 97721.52, 
    100934.1, 101152.3, 101217, 101245, 101242.5, 101284.2, 101326.9, 101401.7,
  102569.2, 102505.9, 102340.9, 102087.9, 101785.7, 101467.9, 101071.7, 
    95105.04, 94305.59, 100816.9, 101183.4, 101140.1, 101196.5, 101243.3, 
    101400.3,
  102489.5, 102369.4, 102123.5, 101849.9, 101504.8, 101228.7, 101026.8, 
    100861.5, 100745.6, 101050.8, 101106.1, 101100.1, 101111.9, 101209.2, 
    101381.6,
  102394.5, 102217.1, 101944.4, 101675.9, 101351.5, 101112.7, 100989.3, 
    100961.6, 100973.3, 101048.4, 101090.2, 101092.3, 101075.1, 101202.4, 
    101379.5,
  102276.9, 102065.4, 101772.8, 101511.8, 101195.4, 101071.2, 101013.7, 
    100861.5, 100885.7, 101067.5, 101118, 101101, 101109.1, 101244, 101420,
  102184.9, 101953.2, 101683.2, 101446.4, 101197.4, 101132.3, 101071.5, 
    100966.7, 101017.9, 101110.8, 101126.5, 101146.6, 101187.9, 101335.9, 
    101512.1,
  102105, 101843.5, 101584.7, 101381.3, 101162.8, 101133.6, 101129.8, 
    100957.6, 101014.1, 101084, 101152, 101217.3, 101286.1, 101445, 101591.6,
  102796.4, 102876, 102889.3, 102776, 102651.6, 102474.8, 102238.1, 102035.6, 
    101826.7, 101210.1, 100995.3, 101047.7, 100820.9, 100490.2, 100491.2,
  102851, 102840.9, 102763.6, 102613.6, 102438.6, 102016.6, 102111, 101771.3, 
    101516.4, 101300, 101000.4, 100833.1, 100778.1, 99047.38, 99890.6,
  102831.1, 102787.4, 102631.3, 102490.6, 102132.7, 98615.88, 101721.8, 
    101888.9, 101599, 101293, 100971.2, 100886.8, 100926.7, 101079.1, 101220.3,
  102790.1, 102707.4, 102547.9, 102382.9, 102224.5, 101844.4, 98128.26, 
    101422.7, 101463, 101413.4, 101234.2, 101190.2, 101257.7, 101374.4, 
    101451.7,
  102793.4, 102701.9, 102567.3, 102416.6, 102254.7, 102154.5, 101866.8, 
    95699.83, 94907.25, 101409.2, 101549.2, 101431.5, 101444.1, 101444.7, 
    101574.3,
  102794, 102699.1, 102572.7, 102461.7, 102262.6, 102162.9, 102092.7, 
    101929.2, 101650.9, 101783.5, 101708.6, 101616.9, 101573.8, 101567.9, 
    101659.2,
  102811.6, 102744.4, 102621.6, 102497.5, 102335.4, 102208.8, 102074.4, 
    102064.9, 102021.9, 101913.4, 101803.5, 101731.5, 101638.8, 101652.8, 
    101765,
  102858, 102771.7, 102634.2, 102503, 102308.7, 102188.2, 102089.8, 101975.1, 
    101930.7, 101941.2, 101893.1, 101813.8, 101758.6, 101817.2, 101892,
  102915.6, 102828.2, 102690.5, 102534.9, 102371.4, 102205.8, 102063, 
    101988.9, 101963.7, 101941.1, 101915.4, 101885.3, 101856.2, 101912, 
    101987.3,
  102948.9, 102820.4, 102668.3, 102488.9, 102283.6, 102128.1, 102007, 101857, 
    101761.8, 101787.2, 101866.4, 101921.4, 101940.9, 102003.5, 102055.3,
  102911.3, 103039.9, 103157.6, 103134.1, 103101.3, 102945.2, 102704.1, 
    102515.6, 102401.1, 101941.6, 101796, 101783.1, 101311.1, 100624.1, 
    100452.3,
  103014.7, 103128.2, 103196.8, 103169.1, 103081.1, 102666, 102734.7, 
    102359.1, 102164, 102221.8, 102109.4, 101921.5, 101608.6, 99468.09, 
    100028.6,
  103085.6, 103219.1, 103204.5, 103187, 102876.5, 99370.75, 102430.8, 
    102618.5, 102398.4, 102272.5, 102154, 102034.7, 101854.2, 101688.5, 
    101512.8,
  103143.8, 103207.5, 103186.1, 103121.8, 103047.8, 102617.2, 98829.99, 
    102017.9, 101995.3, 102186.2, 102184.1, 102092.2, 101995.5, 101926.4, 
    101844.7,
  103206.1, 103241.7, 103217.6, 103128.1, 103024.5, 102864.1, 102500.1, 
    96325.79, 95485.45, 101757.5, 102201.1, 102107.9, 102107.6, 102021.5, 
    102055.2,
  103206.1, 103236.5, 103205.9, 103158.7, 103017.9, 102846.3, 102658.6, 
    102358.4, 101929.5, 101952.5, 102067.4, 102087.9, 102119.7, 102134.3, 
    102153.5,
  103233.6, 103288.1, 103245.8, 103174.2, 103056.3, 102885.6, 102655.2, 
    102428.4, 102170.6, 101921, 101904.8, 102013.5, 102076.5, 102166.9, 
    102225.4,
  103252.7, 103287, 103255.8, 103179.1, 103029.5, 102863.4, 102662.9, 
    102378.8, 102047.5, 101815.2, 101736.6, 101858.1, 101974.6, 102131.6, 
    102231.8,
  103276.6, 103319.1, 103288.3, 103178, 103043.5, 102854.8, 102641.2, 102398, 
    102087.5, 101771.4, 101608.4, 101669.9, 101813.6, 102013.2, 102172,
  103278.3, 103276.6, 103227.4, 103123.7, 102948.8, 102769.3, 102575.9, 
    102290.6, 101953.8, 101616.1, 101455.8, 101476.5, 101607.3, 101833.2, 
    102045.1,
  103320.2, 103526, 103662.4, 103640.8, 103617.7, 103522.3, 103368, 103284.7, 
    103302.6, 102902.6, 102848.7, 102980.8, 102724.4, 102178.8, 101974.2,
  103442.1, 103598.3, 103692, 103692.2, 103667.2, 103390.8, 103480.5, 
    103229.6, 103115.3, 103238.7, 103185.1, 103138.7, 103001.7, 100989.7, 
    101656.3,
  103536.3, 103691.5, 103726.9, 103780.1, 103593.1, 100142.2, 103374.5, 
    103507.6, 103296.1, 103213.2, 103193.4, 103196.9, 103144.2, 103113.2, 
    103032,
  103597.2, 103700.5, 103758.1, 103794.3, 103818.9, 103498.2, 99757.32, 
    103147.3, 103135.3, 103149.7, 103129.6, 103175.9, 103169.2, 103193.6, 
    103161.5,
  103652.3, 103742.4, 103803.8, 103815, 103814.2, 103773.8, 103508.3, 
    97386.36, 96602.5, 102924.4, 103078.5, 103040.8, 103136.5, 103114.9, 
    103157,
  103672.6, 103755.3, 103786.3, 103820, 103778.4, 103715.6, 103650.4, 
    103458.8, 103145.8, 103153.7, 102997.7, 102895.2, 102948.7, 103005.7, 
    103060.8,
  103664.8, 103745.7, 103783.6, 103777.9, 103745.7, 103673.7, 103554.5, 
    103481.2, 103338, 103124.6, 102925.7, 102798.8, 102756.5, 102811, 102889,
  103631.8, 103678.8, 103693.5, 103702.6, 103624.8, 103540.5, 103438.4, 
    103299.1, 103146.2, 103003.2, 102831.3, 102681.8, 102577.2, 102596.6, 
    102664,
  103561.4, 103587.9, 103572.6, 103552.1, 103482.9, 103399.8, 103271.3, 
    103169.1, 103037.6, 102860.3, 102677.7, 102531.7, 102413.3, 102363.6, 
    102415,
  103442.2, 103423.3, 103382.8, 103352.2, 103250.9, 103153.3, 103037, 
    102894.8, 102740.6, 102574.6, 102460.2, 102330.7, 102224.1, 102141.5, 
    102146.6,
  103828.5, 104071.9, 104310, 104431, 104549.6, 104569.9, 104562, 104590.3, 
    104573.3, 104181.3, 104157.2, 104363.8, 104128, 103584.5, 103321.3,
  103944.8, 104149, 104345.8, 104449.5, 104524.7, 104370.5, 104549, 104383.9, 
    104270.5, 104285.3, 104239.8, 104212.1, 104148.6, 102105.2, 102671.5,
  104055.7, 104257.4, 104398.3, 104508, 104393.8, 100918.4, 104269.7, 
    104510.3, 104334.1, 104116.9, 104002.6, 103963.3, 103904.7, 103846.1, 
    103740.3,
  104116.7, 104278, 104375.3, 104430.1, 104469.5, 104207.6, 100432.8, 
    103819.9, 103944.5, 103942.8, 103787, 103662.7, 103602.2, 103549, 103485.9,
  104151.8, 104268.2, 104335, 104345, 104317.6, 104249.9, 103990.2, 97889.24, 
    96999.2, 103326.8, 103533.9, 103332.2, 103253.6, 103162.3, 103124.9,
  104119.3, 104194.9, 104183.7, 104171.2, 104069.2, 103979.1, 103852, 
    103615.7, 103286.2, 103320.1, 103157.5, 102982.2, 102864.8, 102735.6, 
    102673.6,
  104039.2, 104071.3, 104014.2, 103942.2, 103821.5, 103673, 103488.1, 
    103335.5, 103145.2, 102893.9, 102701.4, 102548.3, 102397.5, 102272.8, 
    102169.7,
  103889.6, 103845.8, 103733.4, 103621.1, 103442.4, 103260.9, 103056, 
    102826.6, 102594.3, 102420.2, 102236.2, 102048.9, 101894.4, 101771.7, 
    101679.5,
  103696.2, 103602.3, 103452.2, 103274.3, 103069.8, 102842.1, 102583.7, 
    102358.4, 102137.1, 101898.9, 101690, 101515.2, 101371.2, 101265.9, 
    101193.3,
  103387.4, 103217.6, 103012.5, 102799.9, 102536.9, 102282, 102036.9, 
    101777.4, 101532.9, 101293.3, 101142.5, 100994.6, 100877.3, 100809.2, 
    100780,
  104518.3, 104716.7, 104920.6, 105073.6, 105202, 105248.4, 105194.4, 
    105153.7, 104997.7, 104413.2, 104178.4, 104116.4, 103637.1, 102838.8, 
    102349.1,
  104465.5, 104624.2, 104802.9, 104952.3, 105029.7, 104881.1, 105017.2, 
    104811.3, 104562.6, 104382.5, 104090.7, 103791.4, 103456.7, 101243.5, 
    101491,
  104368.1, 104548.5, 104699.8, 104861.1, 104790.8, 101281.5, 104515.1, 
    104774.7, 104539.6, 104125.1, 103766.9, 103441.2, 103082.7, 102741.3, 
    102336,
  104240.4, 104412.9, 104547.7, 104658.2, 104731.7, 104483.7, 100682.8, 
    103848.2, 103797.8, 103689.7, 103421.2, 103057.7, 102733.5, 102381.6, 
    101983,
  104118, 104283.1, 104402.5, 104473.1, 104504.9, 104468, 104165, 98033.19, 
    96979.96, 103012.9, 103080, 102665.9, 102357.1, 101955.7, 101603,
  103975.7, 104126.5, 104209, 104271.6, 104216.5, 104144.3, 103993.8, 
    103667.2, 103222, 103053.8, 102709.2, 102340.2, 101990.5, 101563, 101169.5,
  103829.4, 103960.7, 104019, 104034.9, 103974.7, 103835.2, 103613.4, 
    103375.5, 103046, 102655.7, 102357.3, 102013.9, 101607.4, 101178.5, 
    100739.3,
  103681.5, 103757.3, 103774.5, 103753.2, 103630.5, 103454.1, 103201.3, 
    102893.4, 102581.3, 102352.1, 102046.5, 101673.6, 101257.2, 100812, 
    100344.6,
  103525, 103566.2, 103541.2, 103459.1, 103313.1, 103089.8, 102821.3, 
    102557.5, 102324.4, 102050.7, 101698.1, 101322.1, 100898.1, 100427.6, 
    99936.55,
  103347.4, 103312.8, 103232.4, 103116.7, 102903, 102665.1, 102414.9, 
    102199.7, 101972.9, 101686.6, 101369.8, 100986.5, 100535.7, 100054, 
    99571.75,
  104041.6, 104119.7, 104253.2, 104374.4, 104544.2, 104667.7, 104731.2, 
    104805.5, 104797.7, 104374.5, 104297.7, 104402.6, 104056.8, 103409.9, 
    103061.4,
  103917.3, 103958.1, 104079.8, 104216.1, 104316.7, 104283.7, 104540.1, 
    104516, 104448.9, 104443, 104309.7, 104184.6, 104004.8, 101941.5, 102382.4,
  103727.1, 103793.9, 103892, 104040.5, 104047.3, 100616.5, 104021.7, 
    104413.4, 104292.1, 104156, 104023.4, 103898.9, 103762, 103626.8, 103426.5,
  103534.8, 103582, 103654.5, 103741.9, 103914.2, 103783.5, 100141.5, 
    103592.1, 103876.2, 103871.4, 103744.9, 103583.6, 103501.1, 103404.1, 
    103227.2,
  103305.7, 103359.6, 103419.4, 103496.6, 103582.1, 103742, 103611.7, 
    97680.62, 96705.26, 103208.5, 103475.2, 103299.7, 103243.4, 103110.5, 
    103009.7,
  103093.4, 103138.1, 103171.6, 103249.2, 103289.9, 103348.2, 103438.8, 
    103308.1, 103177.4, 103317.5, 103163.6, 103036, 102949.2, 102821.4, 
    102720.3,
  102873, 102907.7, 102931.3, 102988.9, 103045, 103078.3, 103081.2, 103113.5, 
    103027.4, 102863.1, 102771, 102674.8, 102572.7, 102458.2, 102347.2,
  102663, 102682.5, 102696.6, 102747.5, 102766.9, 102787.4, 102767.9, 
    102689.6, 102605.6, 102530.9, 102422.5, 102311.1, 102207.8, 102102.8, 
    102004.6,
  102475.7, 102494.2, 102493, 102512.6, 102532.6, 102531.5, 102487.7, 
    102434.2, 102319.4, 102169.8, 102044.9, 101939.2, 101841.2, 101742.2, 
    101634.5,
  102276.7, 102302.6, 102318.2, 102334, 102311.7, 102280.8, 102208, 102091.5, 
    101952.8, 101809.9, 101721.5, 101621.6, 101516.6, 101420.9, 101323,
  104208, 104081.4, 103992, 103864.2, 103761.3, 103648.1, 103532.9, 103477.5, 
    103459.1, 103099.4, 103132.4, 103379.6, 103189.4, 102694.2, 102430,
  104034.5, 103873.1, 103775.4, 103637.2, 103508.9, 103223.1, 103368.7, 
    103254, 103193.2, 103222.5, 103188.7, 103189.2, 103132.9, 101132.8, 
    101649.5,
  103808.1, 103662.9, 103539.2, 103413.7, 103186.4, 99686.29, 102951.9, 
    103232.5, 103128.6, 103039, 102962.8, 102939.6, 102873, 102793.5, 102657.6,
  103605, 103455.4, 103314.7, 103171.8, 103073.5, 102829.5, 99134.01, 
    102619.3, 102838.9, 102829.6, 102748.9, 102686.6, 102632.3, 102578.5, 
    102455.6,
  103398.1, 103265.5, 103125.2, 102982.5, 102885, 102816.1, 102647.4, 
    96715.71, 95903.22, 102382.5, 102591, 102502.3, 102484.5, 102417, 102369.4,
  103205.6, 103057.4, 102900.4, 102783.9, 102666.8, 102612, 102592.9, 
    102497.9, 102355.1, 102500.1, 102415, 102365, 102372.8, 102309.6, 102215.7,
  102984.2, 102848, 102697.7, 102599, 102519.5, 102471.5, 102421.6, 102413.5, 
    102362.8, 102279.2, 102263.7, 102296, 102267.9, 102186.8, 102034.4,
  102773.6, 102640.4, 102508.4, 102437.3, 102356.3, 102333.8, 102289.4, 
    102227.4, 102189, 102214.2, 102238.8, 102233.8, 102183.6, 102065.9, 
    101885.9,
  102556.8, 102460.5, 102365.6, 102313.4, 102272.5, 102245.1, 102190.7, 
    102169.6, 102145.9, 102150.7, 102162.4, 102160.8, 102079.8, 101940.6, 
    101714,
  102392, 102294.9, 102231.8, 102201.9, 102158.6, 102129.4, 102091.9, 
    102063.8, 102059.7, 102070.1, 102073.9, 102042.1, 101957.7, 101803, 
    101567.1,
  104790.1, 104682.9, 104582.4, 104407, 104220.9, 103977.5, 103679.3, 
    103460.7, 103260.9, 102705.9, 102632, 102767.9, 102547.2, 102056.3, 101872,
  104644.3, 104519.5, 104404.1, 104224.4, 104002.9, 103534.9, 103556.8, 
    103200.5, 102971.5, 102888.8, 102761.4, 102665.4, 102574.4, 100601.8, 
    101175,
  104486.2, 104379.2, 104235, 104075.9, 103697.2, 100118.2, 103092.1, 
    103259.2, 102993.1, 102767.7, 102603.5, 102526.5, 102415.2, 102333.4, 
    102214.8,
  104335.3, 104219.2, 104069.7, 103864.4, 103655.1, 103206.5, 99383.4, 
    102552.7, 102631.6, 102616.7, 102464.9, 102352.7, 102249.5, 102160.3, 
    102037,
  104166.8, 104064, 103906.3, 103697.3, 103494.4, 103257.9, 102888.7, 
    96832.9, 95940.96, 102172.1, 102320, 102161.3, 102075.9, 101951.9, 101871,
  104000.6, 103879.6, 103698.2, 103519.4, 103282.1, 103078.7, 102867.4, 
    102585.2, 102248.9, 102265.9, 102119.3, 101969.3, 101873.1, 101750.3, 
    101701.3,
  103807.5, 103702.9, 103532.4, 103350.2, 103144.5, 102905.9, 102674, 102479, 
    102276.2, 102044.6, 101897.5, 101764.3, 101648.6, 101578.9, 101540.7,
  103623.8, 103499, 103326.4, 103152.4, 102916.1, 102693.2, 102451.7, 
    102197.7, 101978.1, 101828.9, 101677.4, 101548.7, 101486.4, 101486.8, 
    101429.2,
  103417.1, 103312, 103145.4, 102950.1, 102722.1, 102473.3, 102199, 101985.4, 
    101779.3, 101586.1, 101437.7, 101414.8, 101438.3, 101414.3, 101345.9,
  103213.3, 103062.1, 102877.1, 102689.4, 102428.4, 102172.8, 101907.5, 
    101658.7, 101438.9, 101287.6, 101319.3, 101408.3, 101408.5, 101383.2, 
    101279.1,
  105038.2, 104918, 104844.2, 104735.6, 104643.8, 104481.5, 104268.9, 
    104099.4, 103872.2, 103258, 103033.8, 102996.7, 102566.2, 101821.2, 
    101381.6,
  104823.5, 104693.2, 104612.7, 104526.6, 104401.3, 104056, 104100.4, 
    103810.4, 103546.3, 103359.9, 103082, 102817.6, 102511.1, 100360.1, 
    100648.2,
  104555.3, 104442.3, 104350.8, 104294.1, 104065.1, 100551.4, 103593.9, 
    103812, 103512.3, 103176.9, 102865.5, 102586.9, 102264.4, 101951, 101571.7,
  104269, 104161.4, 104071, 103985.7, 103918, 103596.7, 99844.81, 102971.3, 
    103004.5, 102904.1, 102645.1, 102305.8, 101987.9, 101674.8, 101339,
  103913.7, 103846.4, 103772.1, 103707.3, 103640.3, 103550.6, 103257.1, 
    97256.7, 96249.91, 102313.6, 102382.4, 102002.5, 101692.6, 101352.2, 
    101145.5,
  103569.1, 103521.6, 103445.9, 103409.2, 103316.3, 103231.5, 103117, 102833, 
    102479.7, 102407.3, 102083.2, 101721.6, 101383.9, 101084.2, 100946.5,
  103215.6, 103191.9, 103137.3, 103099.1, 103033.1, 102921.6, 102773.3, 
    102632.6, 102386.9, 102063.3, 101748.3, 101408.5, 101073.2, 100868.2, 
    100794.6,
  102938.5, 102892, 102828.9, 102785.8, 102690.4, 102590.2, 102432, 102214.4, 
    101978.2, 101742.4, 101430.8, 101098.5, 100839, 100771.6, 100809.6,
  102639.2, 102589.1, 102525.3, 102457.5, 102366.5, 102243.4, 102075.3, 
    101909.6, 101694.7, 101408.5, 101108.3, 100830.5, 100706.8, 100813.4, 
    100894.9,
  102289.7, 102221.9, 102150.6, 102086.3, 101982.5, 101857.2, 101698.3, 
    101505, 101278.1, 101024.9, 100815.5, 100642.9, 100751.4, 100916.5, 
    100948.2,
  104547.3, 104416.7, 104313.3, 104158.8, 104057.5, 103912.2, 103728.7, 
    103567.2, 103391.4, 102844, 102688.1, 102716.9, 102323.4, 101613.2, 
    101178.5,
  104205.3, 104050, 103945.4, 103823, 103697.4, 103348.3, 103413.4, 103192.5, 
    102990.6, 102861.8, 102649.2, 102464.8, 102215.4, 100121, 100458.4,
  103787.6, 103638.3, 103521.2, 103434.5, 103209.6, 99692.86, 102745.9, 
    103056.5, 102794.4, 102589.3, 102364.7, 102177.4, 101949, 101714, 101410.4,
  103371, 103240.9, 103131.5, 103017.1, 102946.2, 102647.1, 98952.56, 
    102149.4, 102358.3, 102284.4, 102116.9, 101895.6, 101707.8, 101493.8, 
    101214.4,
  102909.1, 102818.7, 102727, 102637, 102573.3, 102496.6, 102238.8, 96350.95, 
    95403.64, 101682.9, 101858.4, 101618.9, 101452.2, 101217.8, 101026.6,
  102469.3, 102406.1, 102310.8, 102268.8, 102178.6, 102128.1, 102069.3, 
    101870.5, 101662.3, 101740.2, 101556.8, 101371.9, 101195, 100984.7, 
    100818.3,
  102034.3, 101999.4, 101922, 101884.2, 101833.1, 101773.7, 101695.3, 
    101666.8, 101542.8, 101374.2, 101248.6, 101092.6, 100906.7, 100727, 
    100625.4,
  101708.6, 101656.4, 101573.8, 101552.8, 101492.2, 101450.6, 101371.5, 
    101265.6, 101165.3, 101085.7, 100955.8, 100800.2, 100643.8, 100501.7, 
    100496,
  101322.3, 101273.3, 101210.9, 101167.7, 101109.9, 101056, 100989.9, 
    100948.4, 100861.6, 100741.4, 100622.1, 100498.4, 100364.7, 100295.2, 
    100334.7,
  100868.6, 100808.5, 100749.2, 100718.3, 100672.1, 100621.5, 100562.8, 
    100486.4, 100413.5, 100324.6, 100272, 100190.3, 100105.5, 100113.6, 
    100193.5,
  103042.5, 103053.4, 103082, 103050.8, 103048.7, 102997.7, 102904.7, 
    102854.4, 102760.3, 102283.3, 102199.4, 102314.3, 102023, 101433, 101108.6,
  102636.5, 102604.9, 102628.9, 102610.9, 102585, 102377.3, 102519.8, 
    102380.2, 102273.5, 102228.5, 102085.7, 102001.1, 101876.9, 99876.31, 
    100309.9,
  102141.9, 102097.3, 102091.2, 102116.4, 102022.4, 98623.49, 101715.9, 
    102137.7, 101938.1, 101827.1, 101707.2, 101635.7, 101527.8, 101413.6, 
    101238.2,
  101656.5, 101620.9, 101596.3, 101586.5, 101601, 101424.1, 97877.58, 
    101147.3, 101502.3, 101471.5, 101400.1, 101279.6, 101230.6, 101145.9, 
    101002.1,
  101154.7, 101129.7, 101108.1, 101107.7, 101123.5, 101157.8, 100998.3, 
    95304.26, 94399.48, 100781.7, 101079, 100950.2, 100940.5, 100849.8, 
    100785.2,
  100704.5, 100683.3, 100653.7, 100676.9, 100669.7, 100704.9, 100750.1, 
    100639.4, 100571.2, 100806.9, 100751.9, 100717, 100690.6, 100621.9, 
    100535.5,
  100299.4, 100277.5, 100236.3, 100241.9, 100260.3, 100286.2, 100314.7, 
    100417.9, 100432.7, 100405.8, 100435.2, 100432.9, 100390.8, 100330.7, 
    100242.2,
  100086.3, 100038.6, 99956.92, 99928.62, 99895.37, 99926.18, 99957.36, 
    99969.45, 100018, 100102.5, 100130.3, 100127, 100108.9, 100061.6, 99988.34,
  99938.02, 99880.28, 99779.02, 99687.3, 99609.95, 99593.2, 99613.74, 
    99696.15, 99747.19, 99772.75, 99800.59, 99816.73, 99801.08, 99768.27, 
    99703.13,
  99890.44, 99791.55, 99655.91, 99533.21, 99427.16, 99362.02, 99324.38, 
    99307, 99344.91, 99399.7, 99472.25, 99500.66, 99499.35, 99478.03, 99416.65,
  101673.6, 101727.5, 101822.6, 101897.7, 102023.1, 102111.8, 102174.5, 
    102250.6, 102306.5, 101979.1, 102005.3, 102217.4, 101994.9, 101463.6, 
    101178.6,
  101333.6, 101376.4, 101471.4, 101557.3, 101625.9, 101556.6, 101801.4, 
    101815.8, 101823.6, 101915.9, 101871.1, 101864.6, 101814.5, 99866.88, 
    100332,
  100918.8, 100965, 101067.7, 101181.1, 101193.2, 97880.38, 101121.4, 
    101582.1, 101487.9, 101467.3, 101467.5, 101446.7, 101407.9, 101331.7, 
    101250.4,
  100559.6, 100568.3, 100640.8, 100698.7, 100828.1, 100713.7, 97252.46, 
    100610.2, 101037.3, 101075.6, 101081.3, 101023.4, 101031.6, 101002, 100948,
  100287.9, 100259.9, 100273.7, 100330.9, 100395.5, 100547.7, 100459.6, 
    94837.89, 93887.41, 100333.9, 100678.4, 100594.3, 100625.8, 100584.8, 
    100598.7,
  100231.1, 100160.3, 100093.2, 100085.5, 100052.4, 100075.2, 100175.3, 
    100117.5, 100085.6, 100368.8, 100321.2, 100312.4, 100329.4, 100312, 
    100308.8,
  100239, 100189.9, 100139.2, 100112.9, 100097.2, 100047.4, 99992.48, 100032, 
    100001, 99951.93, 99997.41, 100008.4, 100002.9, 100000.8, 99999.3,
  100267.8, 100192.1, 100093.8, 100042.9, 99952.7, 99892.91, 99818.95, 
    99729.18, 99703.06, 99751.97, 99749.25, 99737.62, 99731.93, 99713.09, 
    99703.57,
  100352.9, 100268.9, 100153.3, 100067, 99975.84, 99872.03, 99769.07, 
    99722.77, 99637.95, 99547.96, 99498.28, 99481.88, 99474.38, 99464.84, 
    99452.64,
  100493, 100379.7, 100243.2, 100103.8, 99982.3, 99908.3, 99862.54, 99700.8, 
    99485.43, 99332.98, 99283.05, 99254.3, 99231.52, 99210.2, 99194.79,
  101316.2, 101332.2, 101402.6, 101461.9, 101575.5, 101668.6, 101741.6, 
    101846.1, 101942.9, 101671.2, 101777, 102095.9, 101970.8, 101575, 101389.4,
  100964.5, 100986.7, 101047.1, 101121.5, 101184.8, 101115.5, 101369.9, 
    101412.5, 101461.2, 101593.5, 101628.3, 101728.7, 101762.8, 99915.49, 
    100483.5,
  100584.7, 100582, 100642.2, 100744.1, 100763.2, 97410.82, 100730.4, 
    101135.9, 101106.5, 101157.4, 101208.4, 101290.8, 101346, 101372.2, 
    101373.9,
  100358.2, 100266.8, 100241.3, 100236.4, 100353.8, 100319.3, 96828.44, 
    100295, 100689.7, 100749.8, 100807, 100839.3, 100916.3, 100988.9, 101030.7,
  100332.5, 100271.3, 100197, 100122.9, 100067.8, 100159.9, 100135.6, 
    94429.14, 93602.18, 100081.4, 100429.3, 100407, 100498.5, 100521.5, 100623,
  100376.6, 100290.4, 100213.8, 100140.1, 100033.6, 99961.58, 100024.2, 
    99994.57, 99957.16, 100220.8, 100180.1, 100168.7, 100191, 100200.7, 
    100242.2,
  100432.8, 100344.7, 100268.5, 100213.4, 100158.6, 100076.5, 99983.57, 
    100004.5, 99962.62, 99937.65, 99971.01, 99986.65, 99979.44, 99965.39, 
    99959.83,
  100512.8, 100410.4, 100315, 100245.5, 100152.6, 100095.1, 100058.3, 
    99972.8, 99943.43, 99985.33, 99944.27, 99909.38, 99887.38, 99861.62, 
    99838.34,
  100561.5, 100492.6, 100411.7, 100337.9, 100279.2, 100190.4, 100107.8, 
    100072.1, 100005, 99919.47, 99808.41, 99753.93, 99700.98, 99644.05, 
    99587.47,
  100625.5, 100538.5, 100464.9, 100368.8, 100295.5, 100224.7, 100173.5, 
    100061.1, 99943.75, 99839.08, 99758.77, 99671.92, 99567.98, 99479.2, 
    99357.45,
  100915.6, 100923.8, 100975, 101030.8, 101132.8, 101209.3, 101268.2, 
    101368.1, 101477.9, 101267.4, 101434.6, 101826.8, 101774.8, 101466.7, 
    101396.3,
  100616.6, 100628.7, 100678.9, 100735.1, 100792.8, 100713.1, 100949.3, 
    101010.6, 101090.5, 101258, 101364.5, 101529.7, 101640.8, 99858.49, 
    100550.5,
  100289.4, 100242.6, 100300.8, 100385.1, 100441.1, 97098.8, 100451.8, 
    100798, 100799.4, 100894.8, 101004.5, 101144.2, 101278.4, 101382.3, 
    101472.8,
  100082.5, 99995.67, 99977.59, 99966.04, 100059.3, 100044.5, 96515.27, 
    100035.8, 100414.7, 100497.4, 100621.7, 100728.2, 100886.2, 101047.7, 
    101178.8,
  99942.47, 99887.98, 99876.62, 99901.03, 99892.57, 99956.05, 99921.38, 
    94155.7, 93399.55, 99887.39, 100236.5, 100290.4, 100443.9, 100558.5, 
    100746.9,
  99903.91, 99818.62, 99782.41, 99784.86, 99811.5, 99811.29, 99824.29, 
    99767.8, 99695.66, 99940.34, 99958.3, 100017.6, 100117.2, 100218.3, 
    100340.3,
  99937.19, 99855.11, 99811.44, 99839.55, 99840.59, 99824.21, 99800.5, 
    99802.73, 99760.1, 99733.15, 99771.97, 99818.07, 99873.89, 99943.55, 
    100036.8,
  100037.4, 99968.65, 99936.21, 99966.4, 99960.49, 99931.8, 99907.55, 
    99860.67, 99848.46, 99876.51, 99827.34, 99817.19, 99831, 99865.16, 
    99920.47,
  100224.2, 100172.3, 100148, 100182.5, 100198.8, 100155.4, 100084.1, 
    100024.8, 99944.21, 99852.65, 99732.6, 99728.7, 99730.59, 99773.15, 
    99818.82,
  100435.7, 100359.6, 100332, 100348.8, 100339.1, 100285.3, 100233.6, 
    100105.3, 99984.18, 99877.99, 99821.77, 99798.84, 99750.88, 99755.93, 
    99765.8,
  100117.6, 100122.7, 100181.6, 100260, 100385, 100494.3, 100569.8, 100692.3, 
    100828.3, 100631.2, 100806.5, 101211.1, 101185.3, 100928.1, 100921.3,
  99824.75, 99816.73, 99865.04, 99948.07, 100046.4, 99997.8, 100285.7, 
    100398.4, 100509, 100710.5, 100848.8, 101013.1, 101140.9, 99387.05, 
    100134.6,
  99559.73, 99496.7, 99516.67, 99592.94, 99693.49, 96378.05, 99766.23, 
    100200.5, 100295, 100433.8, 100585.4, 100750, 100913.1, 101036.3, 101176.2,
  99440.47, 99340.39, 99256.76, 99194.43, 99292.37, 99308.42, 95864.62, 
    99451.1, 99922.48, 100110.4, 100304, 100451.4, 100646.3, 100837.6, 
    101002.6,
  99421.53, 99398.3, 99318.59, 99212.66, 99112.43, 99211.14, 99216.92, 
    93577.45, 92899.3, 99449.48, 99951.57, 100083.2, 100334.3, 100482.9, 
    100735.5,
  99405.72, 99445.21, 99424.95, 99375.47, 99242.83, 99153.66, 99209.08, 
    99168.94, 99144.98, 99475.85, 99605.36, 99774.87, 99982.93, 100193.3, 
    100400.4,
  99405.03, 99534.53, 99556.3, 99543.16, 99514.91, 99455.35, 99366.67, 
    99362.95, 99385.29, 99341.51, 99404, 99551.84, 99716.24, 99896.93, 
    100070.9,
  99421.76, 99565.48, 99608.66, 99647.85, 99627.12, 99640.09, 99639.86, 
    99601.91, 99576.12, 99562.22, 99464.41, 99487.42, 99578.19, 99712.8, 
    99855.62,
  99406.21, 99587.59, 99653.95, 99708.78, 99733.76, 99752.28, 99719.34, 
    99719.31, 99689.91, 99647.73, 99570.91, 99611.95, 99606.96, 99662.94, 
    99733.22,
  99414, 99614.88, 99715.84, 99764.52, 99772.42, 99822.92, 99818.05, 
    99763.34, 99703.39, 99676.3, 99685.51, 99731.07, 99730.84, 99740.66, 
    99735.35,
  99140.16, 99258.92, 99400.43, 99517.55, 99653.15, 99799.41, 99902.68, 
    100033, 100157, 99948.17, 100105.7, 100478.1, 100420.6, 100140.4, 100091.2,
  98839, 98971.55, 99144.13, 99270.8, 99387.91, 99362.08, 99638.42, 99737.5, 
    99856.75, 100037.7, 100145.5, 100293.9, 100384.8, 98634.61, 99368.34,
  98502.59, 98706.02, 98896.62, 99029.02, 99052.38, 95797.71, 99162.05, 
    99525.59, 99598.21, 99754.11, 99890.62, 100040.4, 100181.9, 100294.5, 
    100408,
  98280.23, 98513.98, 98748.35, 98856.17, 98938.39, 98847.36, 95367.04, 
    98912.1, 99330.38, 99485.73, 99663.94, 99791.15, 99969.47, 100147.3, 
    100313.8,
  98223.2, 98542.23, 98790.73, 98895.9, 98859.04, 98876.87, 98814.09, 
    93100.03, 92438.28, 98966.41, 99395.77, 99519.78, 99734.75, 99871, 
    100119.1,
  98286.48, 98591.77, 98812.75, 98918.11, 98903.52, 98839.98, 98935.91, 
    98943.73, 98961.98, 99207.24, 99200.34, 99299.66, 99490.33, 99683.46, 
    99913.25,
  98290.13, 98602.19, 98862.9, 98987.26, 99059.05, 99074.25, 99118.51, 
    99301.51, 99355.87, 99299.2, 99224.52, 99199.38, 99283.31, 99462.86, 
    99691.62,
  98418.55, 98703, 98889.66, 98941.03, 98938.83, 99024.76, 99152.48, 
    99248.49, 99338.98, 99356.62, 99289.16, 99168.33, 99148.1, 99293.99, 
    99527.42,
  98689.48, 98943.94, 99031.58, 99049.51, 99025.66, 99089.99, 99205, 
    99343.33, 99430.13, 99410.02, 99322.21, 99210.65, 99048.25, 99132.09, 
    99353.91,
  99211.08, 99266.25, 99308.41, 99326.1, 99367.47, 99423.73, 99441.12, 
    99426.95, 99415.49, 99422.8, 99388.54, 99290.39, 99047.05, 99033.08, 
    99241.77,
  98101.26, 98221.14, 98433.01, 98684.23, 99000, 99314.68, 99562.99, 
    99813.76, 100027.8, 99884.82, 100094.9, 100499.5, 100464.6, 100144.9, 
    100054.7,
  97946.26, 98050.83, 98258.2, 98512.23, 98779.84, 98956.1, 99370.89, 
    99595.97, 99797.52, 100040.9, 100202, 100388.4, 100524.1, 98750.98, 
    99496.78,
  97710.31, 97879.75, 98124.34, 98404.59, 98566.02, 95485.41, 99022.2, 
    99501.42, 99668.62, 99851.35, 100020.4, 100194.6, 100381.8, 100516.6, 
    100632.5,
  97570.8, 97733.26, 98029.45, 98312.84, 98637.93, 98607.38, 95265.9, 
    98945.52, 99434.28, 99653.52, 99846.42, 99993.5, 100200.7, 100384.9, 
    100559.4,
  97455.85, 97746.02, 98055.7, 98329.27, 98598.7, 98843.59, 98788.8, 
    93125.64, 92539.81, 99125.52, 99629.25, 99762.27, 99998.58, 100145.1, 
    100372.4,
  97648.48, 97934.74, 98206.02, 98430.12, 98583.28, 98678.62, 98848.72, 
    98858.69, 98857.52, 99257.12, 99408.02, 99563.93, 99766.31, 99944.17, 
    100139.6,
  97846.49, 98112.55, 98374.34, 98561.78, 98698.02, 98732.14, 98708.56, 
    98843.19, 99047.41, 99175.23, 99349.31, 99506.91, 99627.08, 99756.44, 
    99909.73,
  98094.65, 98399.59, 98672.92, 98825.04, 98855.18, 98787.68, 98660.35, 
    98612.72, 98836.16, 99132.36, 99359.03, 99519.65, 99653.44, 99732.12, 
    99794.69,
  98650.11, 98875.78, 99033.85, 99111.61, 99097.31, 98938.29, 98565.44, 
    98517.48, 98763.77, 99057.08, 99320.45, 99513.88, 99647.7, 99723.06, 
    99754.53,
  99137.2, 99246.46, 99334.84, 99387.7, 99325.48, 99218.13, 99009.54, 
    98792.59, 98891.2, 99096.59, 99365.91, 99533.75, 99626.97, 99677.12, 
    99682.4,
  98336.3, 98348.3, 98407.49, 98499.08, 98671.57, 98878.44, 99112.63, 
    99399.73, 99690.29, 99635.85, 99938.94, 100405.1, 100387.4, 100033.2, 
    99852,
  98238.12, 98255.85, 98290.65, 98393.51, 98509.89, 98584.52, 98962.91, 
    99215.45, 99497.91, 99835.14, 100081.6, 100312.9, 100464.9, 98632.11, 
    99282.18,
  98132, 98171.28, 98228.23, 98339.93, 98359.24, 95221.07, 98708.41, 
    99193.94, 99430.01, 99715.59, 99964.35, 100203.5, 100394.2, 100480.4, 
    100489.4,
  98034.77, 98033.23, 98131.67, 98258.98, 98463.8, 98370.57, 95068.89, 
    98792.57, 99350.23, 99638.42, 99889.07, 100078, 100305.1, 100452.4, 
    100502.9,
  98083.34, 98164.65, 98236.3, 98360.32, 98498.73, 98711.7, 98632.26, 
    93080.68, 92571.27, 99272.44, 99813.26, 99970.3, 100205.5, 100336.6, 
    100488.9,
  98356.77, 98408.09, 98465.42, 98550.02, 98611.76, 98721.47, 98898.91, 
    98935.96, 98934.55, 99429.55, 99645.64, 99860.66, 100089.5, 100266.5, 
    100424.9,
  98652.3, 98723.36, 98770.08, 98837.92, 98902.18, 98949.9, 98962.2, 
    99085.91, 99189.16, 99282.05, 99500.6, 99732.16, 99954.39, 100163.1, 
    100343.2,
  99045.41, 99135.89, 99158.77, 99233.16, 99235.87, 99268.09, 99263.94, 
    99173.3, 99096.84, 99157.92, 99348.12, 99582.14, 99828.54, 100059.1, 
    100272.8,
  99354.65, 99421.73, 99455.29, 99511.05, 99537.49, 99516.33, 99426.48, 
    99384.54, 99282.83, 99169.56, 99197.63, 99426.07, 99686.48, 99952.26, 
    100189.1,
  99624.33, 99661.8, 99699.62, 99743.95, 99704, 99662.34, 99554.55, 99353.48, 
    99131.76, 98983.07, 99077.73, 99293.38, 99578.19, 99881.95, 100146.4,
  98904.36, 98960.69, 99047.53, 99150.88, 99295.38, 99429.59, 99607.53, 
    99834.73, 100074.2, 99975.79, 100274.3, 100805.2, 100906.2, 100745.2, 
    100799,
  98806.1, 98844.84, 98894.3, 99014.02, 99108.63, 99143.87, 99448.37, 99614, 
    99828.24, 100117.5, 100347.1, 100652, 100898.8, 99289.39, 100127.4,
  98614.44, 98686.41, 98797.05, 98905.05, 98890.7, 95673.4, 99137.68, 
    99560.98, 99720.05, 99951.78, 100176.8, 100463.2, 100760.8, 100995.2, 
    101223.9,
  98587.76, 98538.23, 98549.3, 98657.61, 98902.31, 98759.52, 95393.23, 
    98987.69, 99491.33, 99759.08, 100038.9, 100288.4, 100627.5, 100943.6, 
    101201.2,
  98768.05, 98690.55, 98589.06, 98576.03, 98665.54, 98926.63, 98821.27, 
    93245.96, 92720, 99327.5, 99909.23, 100147.6, 100510.9, 100787.1, 101121.5,
  99054.7, 98986.53, 98863.17, 98725.81, 98659.41, 98740.66, 98919.13, 
    98911.55, 98902.78, 99454.18, 99733.54, 100046.6, 100412.8, 100737, 
    101063.6,
  99264.55, 99260.21, 99242.4, 99193.18, 99091.46, 99008.61, 98939.04, 
    99085.42, 99234.92, 99346.1, 99620.41, 99970.66, 100333, 100679.2, 
    101007.1,
  99481.54, 99477.45, 99496.17, 99493.7, 99448.23, 99430.25, 99356.98, 
    99133.65, 99121.39, 99314.95, 99597.29, 99928.36, 100303, 100659.7, 
    101000.7,
  99593.98, 99649.45, 99713.05, 99773.45, 99783.3, 99720.93, 99651.23, 
    99620.27, 99484.56, 99451.45, 99616.48, 99932.47, 100295.2, 100659.4, 
    100998.1,
  99722.96, 99846.13, 99906.32, 99997.02, 99983.27, 99965.95, 99873.24, 
    99714.52, 99600.67, 99562.23, 99703.3, 99982.03, 100317.9, 100679.3, 
    101003,
  99058.35, 99042.12, 99069.75, 99019.22, 98965.16, 98915.14, 98888.56, 
    98935.34, 99067.8, 98938.67, 99266.91, 99841.95, 99992.37, 99931.21, 
    100126.9,
  99019.67, 99004.35, 99062.71, 99057.92, 99003.48, 98798.3, 98985.91, 
    98969.73, 99084.22, 99343.62, 99614.63, 99958.72, 100231.3, 98729.44, 
    99722.58,
  99009.18, 98905.74, 99056.52, 99076.8, 98961.95, 95574.34, 98948.84, 
    99188.85, 99320.08, 99485.03, 99734.05, 100054.6, 100393.7, 100679.4, 
    101022.2,
  99132.27, 98879.82, 98912.5, 99033.59, 99166.53, 98900.03, 95427.08, 
    99005.26, 99358.66, 99597.23, 99875.85, 100161.6, 100528, 100909.7, 
    101226.3,
  99409.54, 99141.91, 98919.11, 98942.54, 99114.56, 99266.9, 99106.57, 
    93332.97, 92899.09, 99532.78, 100028.8, 100280.1, 100643.2, 100950.6, 
    101340.1,
  99547.69, 99446.13, 99188.61, 99012.16, 99065.25, 99198.09, 99405.39, 
    99391.25, 99328.23, 99854.6, 100098.6, 100399.6, 100743.9, 101087.5, 
    101427.3,
  99673.48, 99650.55, 99582.26, 99356.11, 99214.17, 99296.23, 99366.2, 
    99610.17, 99828.82, 99948, 100180.5, 100496.5, 100807.7, 101143.7, 
    101465.2,
  99797.26, 99839.59, 99826.68, 99778.8, 99574.7, 99511.01, 99536.95, 
    99556.77, 99705.38, 99976.16, 100255.6, 100556.6, 100872.2, 101203.8, 
    101534.4,
  100007.3, 100036.8, 100069.6, 100080, 100021, 99904.1, 99834.07, 99857.79, 
    99900.12, 100063.3, 100296.8, 100593.4, 100899.8, 101227.1, 101563.8,
  100310.5, 100309.2, 100316.4, 100336.9, 100261.8, 100189.7, 100068.9, 
    99937.23, 99882.05, 100006, 100293.7, 100600.1, 100915.4, 101263, 101611.7,
  99252.1, 99067.85, 98953.34, 98817.25, 98704.61, 98670, 98652.6, 98749.96, 
    98959.76, 98877.42, 99183.61, 99712.84, 99823.09, 99670.59, 99735.35,
  99267.94, 99001.43, 98835.7, 98679.13, 98546.3, 98311.01, 98530.55, 
    98569.75, 98759.93, 99060.76, 99356.88, 99661.55, 99922.77, 98304.35, 
    99178.19,
  99305.24, 98994.62, 98797.4, 98657.63, 98447.84, 95041.2, 98380.09, 
    98637.55, 98885.59, 99085.61, 99349.49, 99631.1, 99933.84, 100154.3, 
    100366.8,
  99445.8, 99054.94, 98799.61, 98662.23, 98675.85, 98391.03, 94888.93, 
    98546.69, 98879.8, 99134.11, 99425.05, 99659.73, 99962.91, 100227.9, 
    100459.6,
  99565.75, 99244.1, 98947.47, 98761.41, 98744.39, 98827.23, 98644.2, 
    92785.29, 92435.61, 99068.97, 99559.91, 99739.28, 100044, 100230.8, 
    100548.3,
  99745.12, 99428.23, 99123.15, 98904.57, 98832.35, 98848.27, 99027.29, 
    99000.85, 98922.84, 99402.95, 99628.63, 99870.16, 100143.9, 100387.8, 
    100661.7,
  99939.64, 99720.56, 99415.71, 99167.12, 99013.97, 99024.25, 99036.23, 
    99251.37, 99430.84, 99548.9, 99764.96, 100034.2, 100280.5, 100557, 
    100842.8,
  100161.7, 99997.92, 99752.89, 99515.23, 99288.37, 99224.95, 99285.3, 
    99336.79, 99481.78, 99709.19, 99971.11, 100225.4, 100518.1, 100840.9, 
    101159.1,
  100441.4, 100320.3, 100128.5, 99953.58, 99737.26, 99592.5, 99561.66, 
    99690.23, 99839.49, 100006.6, 100224.8, 100500.3, 100819.6, 101126.3, 
    101409.2,
  100745.5, 100654.9, 100493.3, 100308.9, 100101.5, 99965.16, 99907.55, 
    99933.3, 100061.2, 100224.5, 100509.5, 100803.2, 101097, 101397.1, 
    101646.4,
  98851.69, 98643.27, 98503.3, 98453.24, 98443.98, 98479.84, 98798.52, 
    99252.91, 99623.51, 99569.07, 99844.84, 100312.4, 100366.3, 100179.4, 
    100235.8,
  98771.82, 98607.28, 98535.14, 98506.91, 98433.57, 98214.27, 98697.99, 
    99172.9, 99529.38, 99879.66, 100138.8, 100398.7, 100612.3, 98944.84, 
    99801.14,
  98776.97, 98580.34, 98552.09, 98518.98, 98338.75, 94967.66, 98622.41, 
    99238.37, 99650.37, 99934.87, 100198.1, 100454.2, 100706.9, 100903.1, 
    101070.8,
  98881.63, 98661.59, 98604.88, 98577.9, 98634.93, 98402.59, 95174.41, 
    99107.48, 99671.02, 99995.02, 100285, 100514.8, 100773.8, 100990.4, 
    101180.3,
  99051.32, 98869.22, 98779.23, 98798.43, 98846.95, 99045.26, 98970.66, 
    93397.38, 93085.69, 99913.84, 100399.6, 100590.4, 100829.4, 100979.9, 
    101207.6,
  99305.15, 99120.66, 99023.05, 99045.63, 99095.98, 99254.56, 99531.44, 
    99623.39, 99686.81, 100242.3, 100468.2, 100688.2, 100881.3, 101048.9, 
    101214.4,
  99585.27, 99433.81, 99323.39, 99332.55, 99415.38, 99547.89, 99713.62, 
    100005.1, 100232.7, 100374.5, 100574.2, 100774.7, 100924.5, 101072.8, 
    101192.2,
  99925.88, 99774.27, 99647.7, 99618.8, 99648.36, 99793.48, 99950.13, 
    100115.3, 100293.8, 100509, 100703.6, 100848.4, 100983.4, 101107.1, 
    101257.4,
  100306.8, 100160.9, 100052.4, 100031.5, 100030.2, 100101.2, 100229.1, 
    100430.3, 100589.5, 100706.9, 100820.2, 100937.5, 101068, 101220.7, 
    101360.2,
  100684.9, 100547.2, 100433.3, 100381.3, 100351.1, 100407.1, 100486.7, 
    100576.9, 100694.7, 100793.2, 100947.3, 101090, 101237, 101394.8, 101515.8,
  99336.01, 99292.65, 99296.56, 99389.95, 99619.47, 99811.76, 99934.55, 
    100042.2, 100181.8, 99947.05, 100023.1, 100290.6, 100169.8, 99835.93, 
    99743.12,
  99458.22, 99420.68, 99428.64, 99504.98, 99626.46, 99600.8, 99932.94, 
    100104.3, 100184.8, 100249.3, 100229.3, 100238.8, 100295.2, 98582.34, 
    99342.48,
  99631.01, 99583.61, 99607.52, 99670.19, 99635.55, 96419.27, 100020.6, 
    100315.7, 100389, 100354.6, 100290.6, 100233.4, 100309.6, 100475.9, 
    100629.9,
  99919.18, 99852.1, 99876.59, 99938.98, 100097.1, 99939.31, 96506.38, 
    100253.3, 100489.9, 100494.8, 100430.2, 100310.1, 100362.6, 100583.8, 
    100796.5,
  100213.8, 100179.8, 100187.5, 100247.1, 100382.2, 100504.1, 100384.5, 
    94369.85, 93829.8, 100469, 100612.5, 100466.2, 100491.5, 100631.1, 
    100945.2,
  100450.8, 100410.6, 100423.7, 100463.7, 100533.7, 100637, 100766.3, 100739, 
    100625.4, 100835.9, 100796.8, 100708.6, 100709, 100862.5, 101114.2,
  100616.1, 100610.1, 100609.5, 100652, 100700.1, 100780.5, 100848, 100969.3, 
    101027, 101026.5, 101012.8, 100986.1, 100982.6, 101106.3, 101298.1,
  100765.4, 100770.1, 100751.4, 100781.9, 100804.4, 100894.7, 100982, 101075, 
    101137.2, 101204.5, 101238.2, 101256, 101292.1, 101397.6, 101546,
  100924.9, 100958, 100985, 101034.4, 101066, 101088.6, 101148, 101245.6, 
    101307.8, 101349.3, 101391.9, 101441.6, 101498.1, 101588.8, 101701.5,
  101127.3, 101143.1, 101179.6, 101236.2, 101235, 101262.6, 101289.9, 
    101316.5, 101351.6, 101373.2, 101466.9, 101546.8, 101622.8, 101726.1, 
    101818.8,
  100789.3, 100827.7, 100912.1, 100974.2, 101044.3, 101048.8, 100982.9, 
    100888.4, 100726.4, 100191.8, 100011.4, 100009.5, 99700.41, 99289.42, 
    99264.91,
  100951.6, 100965.4, 101030.7, 101089.4, 101128.5, 100956.7, 101104.8, 
    101015.2, 100856.6, 100704.9, 100494.7, 100314.3, 100114.4, 98233.87, 
    98975.14,
  101067.9, 101088.5, 101154, 101199.8, 101089, 97630.54, 101134.8, 101249.4, 
    101122.6, 100922.9, 100718.2, 100558.6, 100440.9, 100384.2, 100345.5,
  101138.7, 101156.4, 101222.3, 101279, 101354.2, 101116.4, 97403.62, 
    101060.3, 101120.9, 101078.9, 100911.8, 100745.4, 100652.6, 100638.9, 
    100634,
  101275.1, 101317.5, 101348.6, 101409.2, 101463.5, 101479.1, 101286.5, 
    95073.16, 94393.1, 100972, 101062.9, 100866.8, 100830.9, 100780, 100845.4,
  101336, 101369.5, 101396.1, 101441.6, 101475.7, 101529.9, 101576.5, 
    101488.6, 101255.2, 101305.2, 101137.9, 100960.6, 100909.9, 100950.2, 
    101003.5,
  101336.7, 101390.8, 101420.4, 101473, 101511.4, 101581.8, 101616.2, 
    101684.4, 101636.5, 101475.4, 101254, 101064.3, 100968, 101060.8, 101143.8,
  101332, 101388.8, 101401.1, 101452.3, 101489.5, 101604.8, 101683.6, 
    101735.5, 101704.2, 101618.1, 101438.9, 101228.6, 101126, 101205.6, 101312,
  101381.3, 101467.9, 101520.1, 101589.2, 101643.8, 101683.8, 101750, 
    101835.1, 101839.5, 101756.6, 101624, 101460.9, 101343.2, 101368.9, 
    101447.3,
  101476.1, 101547.3, 101600.6, 101674.8, 101688, 101709.6, 101763.6, 
    101795.4, 101815.4, 101781.4, 101747.8, 101650.5, 101545.1, 101540.6, 
    101574,
  101692.4, 101622.3, 101560.3, 101415.2, 101292.6, 101126.6, 100878.2, 
    100655.3, 100380.2, 99715.3, 99530.26, 99836.68, 99988.98, 99973.04, 
    100130,
  101668.4, 101629.4, 101564.8, 101448.5, 101304.9, 100902.2, 100948, 100586, 
    100222.3, 99902.46, 99599.38, 99665.44, 99997.99, 98547.39, 99573.86,
  101586.2, 101603.4, 101576.2, 101500.8, 101193.9, 97576.3, 100754.6, 
    100826, 100453.1, 99988.45, 99605.89, 99633.83, 99995.41, 100392.2, 
    100765.5,
  101484.7, 101476.4, 101501.4, 101471.4, 101438.5, 100979.1, 97142.5, 
    100392.3, 100262.4, 100136.4, 99827.66, 99809.62, 100128.7, 100546.5, 
    100914.1,
  101397.5, 101441.1, 101480.1, 101446.1, 101459.3, 101350.8, 101021.4, 
    94670.55, 93879.62, 100172, 100171.6, 100088.2, 100344.9, 100597.7, 
    101014.7,
  101216.6, 101280, 101339.9, 101389.4, 101388.1, 101390.4, 101365.1, 
    101112.9, 100723.3, 100654.1, 100480.7, 100419.5, 100583.2, 100799.4, 
    101108.4,
  100989.6, 101075.2, 101142.5, 101239.8, 101334.5, 101405, 101396.9, 101393, 
    101240.8, 100985, 100776.8, 100750.9, 100817, 100977.7, 101187.6,
  100816.3, 100901.7, 100958.2, 101093, 101189.3, 101377, 101491.5, 101465.9, 
    101354.4, 101242.5, 101118.2, 101043.7, 101088.9, 101202.7, 101357.9,
  100678.4, 100804.6, 100898.8, 101068, 101216.7, 101398.7, 101532, 101638.6, 
    101614.4, 101508.5, 101394.4, 101324.3, 101321.7, 101377.4, 101463.1,
  100524.5, 100674.9, 100819.8, 101023.4, 101190.4, 101359.7, 101526.8, 
    101632.8, 101660.1, 101631.5, 101617, 101557.2, 101521, 101552.6, 101583.5,
  101030.3, 101046.8, 101039.3, 100944.1, 100860, 100734.8, 100549.2, 
    100454.4, 100452.1, 100175.8, 100365.8, 100766.6, 100692.1, 100379.1, 
    100347.2,
  100791.8, 100836.3, 100834, 100747, 100637.8, 100262.1, 100368.2, 100196.4, 
    100136.1, 100277.9, 100459.7, 100712.1, 100858.7, 99123.54, 99916.79,
  100486.9, 100593.2, 100604.1, 100559.4, 100268.6, 96729.73, 99872.95, 
    100124.8, 100059.6, 100152.9, 100335.5, 100622.5, 100884.3, 101051, 
    101200.7,
  100273.5, 100364.6, 100353.5, 100246.5, 100130.4, 99770.25, 96153.69, 
    99669.45, 99936.67, 99999.3, 100250, 100565.2, 100910.8, 101177.6, 
    101357.2,
  100154.7, 100246.8, 100227.1, 100095.9, 100042.6, 100059.1, 99887.91, 
    93793.68, 93144.84, 99813.32, 100279.3, 100606.1, 100977.5, 101203.5, 
    101471.6,
  100087.6, 100177.5, 100147.7, 100088.5, 100037, 100120.3, 100093.8, 
    99983.32, 99796.66, 100117.8, 100391.6, 100758.9, 101097.4, 101360.6, 
    101590.9,
  100090, 100218.1, 100198.7, 100169.1, 100168.2, 100205.4, 100150.7, 
    100195.2, 100238, 100355.9, 100621.8, 100967.8, 101254.2, 101509.7, 
    101728.6,
  100182.3, 100306.7, 100317.6, 100358.1, 100385, 100416.3, 100396.6, 100393, 
    100459.3, 100655.4, 100921, 101205.2, 101463.7, 101705.2, 101921.4,
  100325.3, 100458.4, 100553.6, 100670.6, 100740, 100758.7, 100750.1, 
    100795.3, 100873.1, 101019.9, 101222.8, 101456.9, 101671.1, 101884.4, 
    102067.9,
  100536.2, 100689.4, 100853.4, 100982.6, 101035.5, 101076.3, 101083.2, 
    101101.4, 101175.9, 101291.1, 101497.2, 101690.1, 101870.9, 102054, 
    102185.7,
  99915.42, 100124.5, 100392, 100658.6, 100923.1, 101114.9, 101225.3, 
    101290.3, 101342, 101009.5, 101070.9, 101320.6, 101120.2, 100664.9, 
    100510.6,
  99721.41, 99866.35, 100094.5, 100371.6, 100629.1, 100664.2, 100958.8, 
    101010.6, 101023.2, 101055.9, 101095, 101156.2, 101111.1, 99194.38, 
    99867.02,
  99650.04, 99797.12, 99956.51, 100206.2, 100336, 97073.24, 100572.6, 
    100846.6, 100848.7, 100883.1, 100955, 101050.7, 101044.6, 101052.5, 
    101039.3,
  99676.22, 99772.95, 99877.41, 100039.3, 100270.8, 100163.5, 96638.78, 
    100361.9, 100711.3, 100846.4, 100996.9, 101037.7, 101048.1, 101064, 
    101081.9,
  99616.69, 99667.34, 99755.04, 99900.45, 100230.6, 100430.6, 100307.4, 
    94473.02, 93943.81, 100779, 101093, 101078.1, 101096.6, 101068.7, 101119.3,
  99738.12, 99765.87, 99832.98, 99962.8, 100186.4, 100369.1, 100531.3, 
    100596.3, 100674.5, 101079.7, 101158.3, 101183.3, 101182.1, 101178.9, 
    101183.7,
  99959.25, 99975.96, 100014.8, 100149.1, 100312.4, 100494.9, 100686.1, 
    100972.1, 101156.1, 101241.7, 101313.5, 101358.6, 101356.5, 101365.5, 
    101352.6,
  100273.6, 100294.3, 100319.9, 100410.8, 100525.4, 100733.4, 100942.6, 
    101137.2, 101302.5, 101453.5, 101524.8, 101549.8, 101546.8, 101532.9, 
    101514.7,
  100684.5, 100727.8, 100777, 100884.4, 101006.8, 101155.7, 101324.7, 
    101511.3, 101634.8, 101701.9, 101739.6, 101748.3, 101730.7, 101696.7, 
    101655.5,
  101193.2, 101235.3, 101311.1, 101378.9, 101435.6, 101545.8, 101650.7, 
    101736.6, 101822.2, 101866.2, 101935.2, 101944.2, 101912.1, 101870.2, 
    101804.8,
  99852, 99972.51, 100176.5, 100467.2, 100835.3, 101183.7, 101456.2, 
    101701.5, 101899.5, 101689.6, 101820.8, 102116.7, 101969.9, 101524.5, 
    101343.6,
  99781.43, 99837.91, 100003.8, 100306.9, 100656.9, 100873.9, 101348.2, 
    101587, 101734.1, 101903.1, 101950.9, 101989.5, 101947.5, 99980.57, 
    100584.8,
  99643.7, 99783.04, 99916.09, 100226.2, 100440.3, 97362.97, 101064.8, 
    101573.6, 101700.5, 101786.8, 101806.7, 101807.5, 101750.7, 101675.9, 
    101579.8,
  99644.51, 99671.79, 99863.13, 100155, 100566.5, 100559.5, 97279.59, 
    101139.5, 101568.2, 101656.1, 101671.8, 101623.5, 101575.9, 101505.5, 
    101418,
  99712.09, 99780.61, 99941.07, 100247.2, 100622.5, 100951.5, 100917.1, 
    95154.13, 94513.38, 101279.1, 101578.7, 101510.7, 101476.1, 101394.7, 
    101357,
  99936.27, 100021.7, 100166.3, 100432.8, 100688.2, 100934.3, 101190.6, 
    101198.1, 101197.3, 101499.1, 101499.9, 101476.2, 101421.4, 101341, 
    101282.7,
  100169.8, 100285.8, 100418, 100611.8, 100808.3, 101009.8, 101208.1, 
    101435.7, 101525.8, 101506.3, 101514.1, 101465.5, 101397.2, 101338.7, 
    101278.3,
  100417.3, 100532.5, 100624.9, 100788, 100938.3, 101161.1, 101344.4, 
    101481.1, 101561.6, 101625.1, 101570, 101494.9, 101420.1, 101357.6, 
    101306.4,
  100712.8, 100827.1, 100929.4, 101089, 101242, 101409.9, 101552.5, 101684.7, 
    101720.1, 101690.5, 101640.3, 101568.6, 101487, 101420.3, 101362,
  101136.7, 101231.2, 101344.3, 101448.7, 101518.5, 101626.2, 101692.1, 
    101726, 101751.8, 101730.2, 101727.9, 101665.3, 101580.2, 101509.9, 
    101444.7,
  99924.36, 99973.17, 100032.8, 100125.6, 100301.2, 100544.8, 100800.8, 
    101084, 101405.7, 101291.2, 101506.7, 101818.1, 101652.2, 101118.5, 
    100853.9,
  99818.73, 99883.5, 99964.41, 100100.8, 100306.1, 100401.8, 100834.3, 
    101122.7, 101369.1, 101605.9, 101723.5, 101776.9, 101724.9, 99698.72, 
    100243.7,
  99688.64, 99877.88, 99977.02, 100174.3, 100234.7, 97087.33, 100825.4, 
    101294.6, 101474, 101582.8, 101647, 101673.6, 101625.4, 101526.7, 101373.4,
  99659.52, 99856.63, 100004.9, 100214, 100501.1, 100424.7, 97133.67, 
    101011.4, 101428.7, 101543.5, 101598.3, 101560.3, 101520.2, 101412.4, 
    101287.2,
  99758.68, 99923.77, 100080.4, 100322, 100612.1, 100899.5, 100816.5, 
    95031.75, 94398.46, 101170.6, 101486.4, 101444.3, 101409.6, 101327.2, 
    101289.5,
  99917.11, 100050.2, 100201, 100449.7, 100675, 100885.2, 101127.7, 101127, 
    101096.1, 101391.2, 101416.3, 101420.8, 101386.5, 101325.6, 101267.9,
  100123.4, 100255.2, 100393, 100588.9, 100780.5, 100952, 101112.9, 101318.6, 
    101434.5, 101431.7, 101457.7, 101431.9, 101375.4, 101334.6, 101285.6,
  100362.2, 100457.9, 100546.1, 100684.8, 100808.9, 100983.9, 101161.8, 
    101305.1, 101410.9, 101503.4, 101494.2, 101461, 101416.4, 101375.4, 
    101337.6,
  100584.2, 100664.6, 100727.6, 100841.5, 100954.4, 101102.1, 101260, 
    101433.3, 101528.8, 101550.1, 101551.5, 101523.4, 101475.3, 101437.5, 
    101402,
  100918.4, 100954.3, 101010.1, 101078.4, 101136.2, 101236.4, 101341.6, 
    101426.6, 101500.6, 101531.1, 101593.9, 101590.7, 101556.2, 101525.6, 
    101492.7,
  100423.6, 100451.9, 100480.5, 100501, 100532.4, 100542.7, 100492.2, 
    100481.8, 100549.7, 100342.8, 100593.7, 101063, 101094.9, 100826.4, 
    100744.3,
  100395.3, 100405.2, 100407.4, 100456.3, 100520.1, 100414.6, 100560.2, 
    100567.2, 100644, 100842.4, 101040.2, 101259.8, 101371, 99505.62, 100192.8,
  100327.6, 100418, 100476.7, 100551.8, 100482.2, 97115.67, 100625.7, 
    100872.4, 100996.7, 101103.2, 101255, 101387.8, 101471.8, 101474.5, 
    101377.6,
  100336.1, 100399.7, 100500.9, 100594.5, 100760.9, 100546.5, 97062.64, 
    100835.4, 101157.8, 101308.4, 101418.8, 101456.2, 101488, 101450.7, 
    101354.9,
  100448.4, 100514.6, 100596.3, 100726.4, 100868.5, 101035.5, 100871.7, 
    94927.38, 94398.14, 101222.2, 101530.2, 101492.5, 101516.3, 101468.2, 
    101435,
  100562.1, 100630.9, 100711.9, 100858.8, 100975.2, 101102.6, 101266.6, 
    101229.1, 101152.8, 101507.9, 101565.2, 101593.3, 101589.1, 101546.4, 
    101499.7,
  100643.7, 100747.8, 100843.8, 100973.5, 101094, 101211.7, 101332.1, 101506, 
    101615.9, 101619.1, 101670, 101686.8, 101682.9, 101663.6, 101618.1,
  100698.8, 100823.5, 100918.4, 101033.2, 101131.8, 101304.8, 101470.7, 
    101580.7, 101655.6, 101753.2, 101789.2, 101798, 101796.6, 101780.4, 
    101758.8,
  100684.7, 100822.7, 100939.6, 101092.8, 101252.9, 101443.3, 101621.7, 
    101793.6, 101878.6, 101907.6, 101916.8, 101922.7, 101921.6, 101914.7, 
    101901.1,
  100762.1, 100896, 101043.1, 101221.7, 101399.5, 101611.7, 101767.8, 
    101879.6, 101945.6, 101982.2, 102050.9, 102064.6, 102069.3, 102071.8, 
    102058,
  101586.9, 101627.8, 101671.8, 101657.1, 101629.4, 101525.7, 101356.9, 
    101238.5, 101153.3, 100785.7, 100800.1, 101011.8, 100839.6, 100405.4, 
    100247.5,
  101662.1, 101686.8, 101734.4, 101756.6, 101724.3, 101445.5, 101563.7, 
    101399.5, 101283.2, 101262, 101225.7, 101214.8, 101154.2, 99205.45, 
    99876.51,
  101677.8, 101772.9, 101831, 101866.6, 101663.8, 98156.95, 101586.5, 
    101731.6, 101637.2, 101509.6, 101420.7, 101380.1, 101323.2, 101271.5, 
    101184,
  101643.5, 101739.8, 101848.2, 101905, 101950.7, 101618.7, 97919.55, 
    101575.1, 101683.1, 101713.4, 101619.7, 101521.4, 101471.1, 101403.4, 
    101327.2,
  101627, 101749.6, 101887.3, 101961.9, 102025.8, 102025, 101752.9, 95540.44, 
    94959.12, 101681.3, 101864.6, 101716, 101682.6, 101574.8, 101573,
  101636.3, 101791.7, 101915.5, 102033.8, 102070, 102086, 102127.3, 102023.6, 
    101850.1, 102042.2, 102014.9, 101921.6, 101877.5, 101805.6, 101776,
  101643, 101823.9, 101977.2, 102080.5, 102134.9, 102221.2, 102256, 102308.6, 
    102316.5, 102247.5, 102188.2, 102143.9, 102080.6, 102029.4, 101983.7,
  101677.4, 101879.8, 102014.7, 102116.8, 102208.9, 102314.6, 102399.3, 
    102425.1, 102402.2, 102405.9, 102372.7, 102325.1, 102281, 102235.7, 
    102202.3,
  101724.1, 101947.2, 102107.6, 102292.4, 102433.6, 102543.8, 102605.2, 
    102643.8, 102643.6, 102606.3, 102557.7, 102513.7, 102464.1, 102418.7, 
    102380,
  101774.9, 102061.4, 102331.2, 102548, 102649, 102735.4, 102760.2, 102759.6, 
    102743.6, 102712.4, 102723.4, 102694, 102644, 102598.3, 102541.1,
  101910.9, 102035.5, 102190.2, 102301.7, 102414.1, 102478.7, 102494.3, 
    102512.4, 102472.1, 102071.4, 102052, 102209.4, 101914.1, 101343.8, 
    101071.4,
  102161.4, 102257.5, 102369.2, 102475.9, 102541.5, 102409.8, 102625.9, 
    102548.7, 102467.9, 102442.3, 102357.9, 102272.6, 102099, 100008.1, 
    100573.1,
  102319.8, 102438.8, 102511, 102591, 102448.5, 98931.6, 102526, 102750.5, 
    102674.3, 102557.2, 102414.5, 102325.4, 102165.9, 102039.5, 101887.3,
  102369.8, 102456.1, 102525.8, 102580.8, 102609.4, 102378.8, 98626.05, 
    102447.4, 102572.3, 102623, 102511.3, 102366.7, 102234.8, 102112, 102027.7,
  102383.2, 102470.6, 102539.1, 102611.5, 102660.8, 102659.5, 102474.3, 
    96225.42, 95565.39, 102435.8, 102607.2, 102446.5, 102348.3, 102195.3, 
    102193.8,
  102386.1, 102493, 102573.1, 102662.7, 102717.1, 102746.2, 102757.9, 
    102685.8, 102529.9, 102699.1, 102675.6, 102564.8, 102484.3, 102379.2, 
    102343.9,
  102390.6, 102524.4, 102616.6, 102679.5, 102753.5, 102816.9, 102858, 
    102897.2, 102886.7, 102809.9, 102746.9, 102699.2, 102627.2, 102573, 
    102536.9,
  102430.5, 102525.4, 102622.6, 102701.7, 102770.5, 102847.3, 102901.9, 
    102915.8, 102888.9, 102889.6, 102861.1, 102816.4, 102782.3, 102745.7, 
    102725.6,
  102462.9, 102581.9, 102734.5, 102874.8, 102974.6, 103012.5, 103022.8, 
    103031, 103023, 102984.1, 102943.4, 102910.5, 102879, 102857.8, 102840.5,
  102543.7, 102756.5, 102955.9, 103078.8, 103116.7, 103122.9, 103090.3, 
    103032.1, 103008.7, 102984.5, 103012.6, 102994.3, 102964, 102934.1, 
    102893.8,
  101501.5, 101490.3, 101523.8, 101584.9, 101707.6, 101872.3, 102039.6, 
    102229.9, 102407.3, 102213, 102402, 102750.4, 102618.9, 102183.6, 102023.5,
  101860.5, 101855.6, 101898, 101987, 102061.4, 102036.2, 102337.3, 102461.6, 
    102545.6, 102704, 102765.6, 102836.6, 102800.7, 100799.6, 101430.6,
  102125.6, 102167.2, 102201.6, 102304.1, 102191.8, 98776.62, 102476.1, 
    102737.1, 102801.1, 102821.2, 102831.5, 102824.8, 102766, 102718.7, 
    102652.1,
  102193.6, 102254.5, 102338, 102438.4, 102527, 102311.4, 98620.15, 102563, 
    102821.3, 102890.8, 102871, 102786.9, 102727, 102669.3, 102652.6,
  102220.8, 102289.7, 102374.8, 102479.1, 102574.6, 102674.1, 102537.4, 
    96320.02, 95646.94, 102686.8, 102909.7, 102777.9, 102704.9, 102627.8, 
    102705.6,
  102270.7, 102347.5, 102434.7, 102541.2, 102607.4, 102647.4, 102739.1, 
    102737.5, 102679.3, 102930.9, 102931.2, 102854.9, 102799.1, 102752.3, 
    102763.9,
  102268.4, 102354.9, 102446.1, 102526.5, 102611.4, 102725.6, 102812.2, 
    102929.5, 103014.1, 103017.4, 103003, 102960.5, 102900, 102856.5, 102829.5,
  102217.1, 102262.8, 102341.2, 102430, 102496, 102662.8, 102846.5, 102957.6, 
    103022.3, 103076.6, 103067, 103028.2, 102977, 102914.5, 102851.8,
  102191, 102244.6, 102343.7, 102491.7, 102604.7, 102750.3, 102907.8, 
    103046.1, 103113, 103118.4, 103086.4, 103028.6, 102943.8, 102842.3, 
    102730.4,
  102248.1, 102368.8, 102473.3, 102586.3, 102675.4, 102806.7, 102957, 
    103035.3, 103092.7, 103071.6, 103061.8, 102971, 102835.9, 102677.6, 
    102506.3,
  101290.9, 101057, 100857.2, 100701.7, 100646.2, 100650.4, 100686.3, 
    100792.5, 100937, 100789, 101066.8, 101524.2, 101555.7, 101366, 101408.4,
  101611.3, 101437.6, 101255.8, 101196.9, 101124.8, 100995.4, 101194.4, 
    101262.1, 101360.4, 101562.4, 101707.8, 101913.3, 102014.4, 100263.6, 
    101108.6,
  101836.8, 101764.9, 101660.1, 101657, 101399.4, 98055.21, 101607.5, 
    101847.8, 101899.7, 101978.1, 102086.5, 102220.9, 102335, 102436.2, 102534,
  101938.2, 101923.3, 101937.7, 101934.1, 102003.5, 101653.3, 98106.53, 
    101893.9, 102192.4, 102301, 102369.9, 102408.5, 102517, 102618.6, 102694,
  102020.1, 102055.1, 102106.9, 102155.8, 102210.8, 102297.4, 102033.6, 
    95871.72, 95297.28, 102261.2, 102544.7, 102517.5, 102579.4, 102606.8, 
    102727.6,
  102103.1, 102137, 102198.5, 102265.7, 102305.1, 102325.2, 102432.4, 
    102341.9, 102251.3, 102556.1, 102602, 102599.8, 102633.2, 102662.9, 
    102721.5,
  102090.2, 102151.9, 102267.6, 102314.6, 102388.7, 102448.6, 102482.9, 
    102579, 102636.9, 102603.5, 102604.4, 102614.2, 102620, 102648.9, 102679,
  101880.6, 102083.6, 102167.1, 102250.1, 102271.6, 102410.4, 102508.6, 
    102520.8, 102497, 102510.2, 102492.3, 102484.5, 102504.1, 102561.6, 
    102629.3,
  101648.3, 101887.3, 102001.4, 102165.8, 102330.8, 102469, 102478.2, 102488, 
    102417.4, 102315.5, 102223.2, 102185.6, 102193.2, 102269.5, 102385.1,
  101641.5, 101843.1, 102039, 102286.3, 102404.9, 102498.3, 102452.9, 
    102306.8, 102113.2, 101929.8, 101832.8, 101762.3, 101761.7, 101880, 
    102066.5,
  101814.8, 101525.5, 101206.4, 100903.4, 100677.5, 100474.9, 100252.6, 
    100175.2, 100187.8, 99930.71, 100085.4, 100501.5, 100547.4, 100392.7, 
    100468,
  101976.9, 101741.8, 101449.9, 101208.6, 100973.7, 100621.9, 100663.6, 
    100456.5, 100402.9, 100456.3, 100535.6, 100708.8, 100859.6, 99242.69, 
    100112.1,
  102054.5, 101905.8, 101719.3, 101537.7, 101122.8, 97681.36, 100973.5, 
    101026.8, 100882.1, 100831.1, 100849.9, 100967.2, 101130.3, 101298.7, 
    101481.4,
  102102.9, 101970.8, 101898.7, 101751.6, 101669.8, 101195.4, 97545.28, 
    101094, 101253.8, 101298.9, 101275.5, 101318.8, 101461.3, 101650.7, 101788,
  102133.9, 102054.9, 101973.8, 101907.7, 101851.1, 101818.2, 101443.4, 
    95286.99, 94763.75, 101466, 101688.7, 101648.3, 101753.3, 101836.6, 
    102024.9,
  102050.9, 102002.4, 101994.3, 101942.4, 101914, 101875.5, 101909.3, 
    101788.3, 101621.5, 101892.5, 101926.7, 101904.2, 101991.4, 102071.5, 
    102222.1,
  101876.8, 101842, 101928.7, 101887.6, 101893.4, 101889.1, 101862, 101922.7, 
    101997.3, 101969.3, 101997.4, 102062.3, 102127.8, 102209.2, 102324.4,
  101702.4, 101686, 101818.9, 101863.2, 101834, 101802.6, 101782.9, 101726.7, 
    101719, 101802.2, 101905.2, 101995.9, 102131.3, 102277.6, 102411.1,
  101730.6, 101763.7, 101876.6, 101943.5, 101944.2, 101866.2, 101738.5, 
    101655.1, 101596.3, 101570.8, 101638.3, 101812.6, 102001.9, 102180.2, 
    102377.7,
  101938, 102007.2, 102051.3, 102036.4, 101933.7, 101826.5, 101686.2, 
    101543.3, 101424.9, 101336.8, 101346.6, 101479.4, 101721.4, 101998, 
    102265.2,
  102477.1, 102308.9, 102107.3, 101925.8, 101739.5, 101575.2, 101308.4, 
    101147, 101141.3, 100819.5, 100890.4, 101185.8, 101109, 100812.1, 100751.1,
  102448.4, 102308.3, 102136.4, 102021.3, 101833.6, 101499.2, 101544.7, 
    101267.9, 101113.6, 101092.1, 101081.6, 101144.6, 101228, 99483.91, 
    100231.8,
  102355, 102264.3, 102124, 102102, 101814.8, 98270.16, 101596.4, 101674.1, 
    101471, 101304.7, 101182.1, 101168.3, 101217.2, 101291, 101377,
  102233.6, 102164.7, 102054.9, 102060.2, 102072, 101703, 97954.63, 101495.1, 
    101606.4, 101605.7, 101470.3, 101353.1, 101329.4, 101356.7, 101421.3,
  102107.2, 102060.4, 101981.8, 101977, 102063.9, 102036.2, 101792.6, 
    95608.48, 94986.61, 101614.5, 101757.2, 101576.7, 101530.2, 101441.9, 
    101501.7,
  101947.4, 101904.8, 101881.8, 101932.6, 101980.8, 101972.7, 102033.1, 
    101938.7, 101792.6, 101985.8, 101912.5, 101794.5, 101710, 101633.4, 
    101617.4,
  101792.7, 101796.5, 101838.3, 101937.2, 101963.6, 101980.7, 102002, 
    102043.4, 102094.9, 102069.9, 102018.4, 101970.4, 101892.9, 101829.7, 
    101793.2,
  101700.7, 101729.6, 101835, 101978.9, 101978, 102001.2, 102044.2, 102021.4, 
    101995.9, 102007.7, 102033.4, 102062.2, 102050.1, 102038.3, 102028.9,
  101689.2, 101737.8, 101882.9, 102002.7, 102060.7, 102068.4, 102066.9, 
    102070.8, 102090.8, 102062.2, 102025.5, 102072.5, 102124.2, 102160.3, 
    102184,
  101706.3, 101785.8, 101957.6, 102042.9, 102067.6, 102083.9, 102077, 
    102031.4, 102037.8, 102042.4, 102038.4, 102056.2, 102142.9, 102237.6, 
    102297.6,
  102434.1, 102542.3, 102614.5, 102647.2, 102679.6, 102654.2, 102521.6, 
    102369.4, 102221.7, 101793.6, 101812.1, 102024.1, 101804.2, 101313.8, 
    101113.1,
  102288.8, 102410.5, 102514.4, 102556.8, 102600.9, 102451.4, 102605.5, 
    102446.1, 102296.8, 102181.3, 102072.1, 102015.7, 101981.6, 100070.7, 
    100688.6,
  102073.6, 102256.6, 102397.8, 102469.8, 102418, 98953.48, 102442.5, 
    102650.7, 102509.3, 102380, 102219.5, 102115.2, 102020.9, 101974.7, 
    101903.4,
  101824.5, 102043.1, 102218.1, 102331.4, 102417.5, 102292.1, 98564.12, 
    102293.6, 102488.2, 102500.5, 102400.8, 102271.8, 102172.8, 102072.7, 
    101970.5,
  101591.4, 101826.7, 102030.8, 102193.1, 102309.4, 102402.2, 102298.2, 
    96247.2, 95513.33, 102360.2, 102540.8, 102414.1, 102323.5, 102185.1, 
    102092.2,
  101388.1, 101622.1, 101851.1, 102042.2, 102173.1, 102294.9, 102391.5, 
    102378.4, 102295.8, 102602.5, 102599.8, 102541.2, 102459.4, 102332.2, 
    102205.7,
  101211.4, 101451.9, 101693.8, 101926.2, 102084.7, 102217.9, 102373.2, 
    102495, 102597.3, 102630, 102649.7, 102630.6, 102558.6, 102453.4, 102307.4,
  101078.8, 101322.6, 101568.3, 101825.9, 101981.2, 102132, 102346.3, 102447, 
    102548.9, 102633, 102688, 102698, 102648.1, 102551.9, 102405.2,
  100988.2, 101235.5, 101488.8, 101778.3, 101974.2, 102141.2, 102341.3, 
    102507.9, 102636.8, 102695, 102724.8, 102747.2, 102720.5, 102643.9, 
    102503.2,
  100940.3, 101187.8, 101464.8, 101764.2, 101970.6, 102156.5, 102343.7, 
    102478.8, 102609.7, 102674.8, 102739.2, 102799.3, 102798, 102755.4, 
    102644.7,
  101862.5, 101925.9, 102004, 102157.6, 102356.4, 102532.6, 102602.4, 
    102632.8, 102576.3, 102178.1, 102185, 102398.9, 102229, 101746.3, 101532.1,
  101777.5, 101861.4, 101968.8, 102131, 102317.1, 102358, 102606.9, 102612.3, 
    102573, 102578.5, 102492.5, 102462.1, 102409.8, 100458.3, 101068.1,
  101626, 101788.4, 101916.6, 102089, 102176.3, 98855.5, 102444.3, 102757.2, 
    102718.9, 102669.8, 102630, 102603.5, 102561.2, 102507.1, 102368.3,
  101431, 101608.5, 101807.7, 101988.4, 102229.2, 102139.7, 98586.31, 
    102355.9, 102644.4, 102716.4, 102715.2, 102696.1, 102697.4, 102651.3, 
    102538.9,
  101249.4, 101417.7, 101627.8, 101863.3, 102108.1, 102339.5, 102254.9, 
    96335.49, 95596.53, 102447.3, 102803.1, 102755, 102777.5, 102697.2, 
    102656.5,
  101060.2, 101234.1, 101441.7, 101701.8, 101958.7, 102179.3, 102356, 
    102363.1, 102264.3, 102609.2, 102776.8, 102819.6, 102854.8, 102782.2, 
    102696.5,
  100869.9, 101060.5, 101263, 101536.2, 101823.6, 102082.9, 102248.5, 
    102415.6, 102522.7, 102614.3, 102786.3, 102875.1, 102892.8, 102834, 102697,
  100717.6, 100917.4, 101104.1, 101391.6, 101666.6, 101932.1, 102157.8, 
    102347.2, 102527, 102687.4, 102832.3, 102936.9, 102962.4, 102894, 102736.7,
  100648.1, 100823.1, 101005.4, 101291.3, 101579.4, 101857.2, 102112.4, 
    102388.8, 102605.7, 102743.5, 102883.5, 102991.1, 103021.5, 102963.1, 
    102798.3,
  100666.8, 100818.7, 101000.9, 101270.2, 101544.2, 101820.2, 102095.6, 
    102380.8, 102607.9, 102741.1, 102920.5, 103052, 103109.2, 103069.2, 
    102923.4,
  101588.4, 101585.4, 101620.9, 101640.2, 101660.4, 101673, 101652.1, 
    101685.2, 101760.2, 101512.7, 101676.3, 102037.1, 101952.5, 101598.2, 
    101458.2,
  101493.1, 101500.6, 101597, 101664.9, 101730.6, 101597.7, 101773, 101721.5, 
    101757.6, 101874.2, 101971.4, 102085.1, 102172.1, 100286.8, 101008.4,
  101386.3, 101445.8, 101587.7, 101690.2, 101657.9, 98202.57, 101766.5, 
    101937.9, 101954, 101983.2, 102061.2, 102162.2, 102282.6, 102315.3, 
    102299.3,
  101259.8, 101357.1, 101553, 101672.5, 101811.1, 101611.9, 97985.54, 
    101722.5, 101990.9, 102091.5, 102199, 102301.4, 102413.6, 102469.7, 
    102457.6,
  101150.3, 101270.7, 101473, 101648.5, 101785.2, 101902.8, 101760.7, 
    95767.13, 95170.82, 102020.3, 102362.8, 102413.7, 102518.4, 102515, 
    102547.9,
  101071.6, 101201.6, 101429, 101608, 101780.9, 101864.9, 102009.5, 101944.6, 
    101824.7, 102282, 102422.7, 102534.9, 102613.5, 102605.4, 102564.4,
  100994.4, 101128.7, 101379.4, 101559.8, 101766.3, 101887.2, 101971.5, 
    102090.7, 102226.7, 102341.6, 102505.7, 102633.9, 102679.1, 102648.9, 
    102560.2,
  100958.2, 101111.4, 101352, 101535.6, 101714.7, 101863.7, 102019.7, 
    102082.6, 102216.5, 102427.2, 102613.9, 102728, 102765.5, 102705.3, 
    102603.2,
  100925.4, 101076.8, 101307.3, 101529.3, 101697.3, 101883.1, 102060.5, 
    102232.1, 102417.4, 102559.9, 102718.7, 102814.6, 102838.2, 102769, 
    102659.3,
  100929.9, 101046.1, 101263.4, 101499, 101689.4, 101894.8, 102107.4, 
    102274.6, 102454.8, 102587.2, 102798.8, 102903.7, 102928.4, 102863.2, 
    102749.1,
  101522.8, 101524.9, 101603.1, 101708.8, 101855.7, 101934.3, 101855.2, 
    101739.7, 101657.5, 101267.5, 101326.2, 101629.9, 101540.4, 101226.3, 
    101179.5,
  101322.7, 101330.3, 101470.1, 101610.8, 101798.6, 101685.1, 101875.1, 
    101697.9, 101624.8, 101615.8, 101625.7, 101699.5, 101761, 99960.4, 
    100723.2,
  101099.7, 101184.1, 101354.7, 101578.8, 101641.8, 98221.16, 101671.2, 
    101816.8, 101718.7, 101700.4, 101701.9, 101760.1, 101867.1, 101932.6, 
    102027.2,
  100915.4, 101055.5, 101290.3, 101556.8, 101709.3, 101571.2, 97865.04, 
    101573.8, 101778.9, 101806.3, 101842, 101887.6, 101987, 102112.5, 102191.4,
  100796, 100992.7, 101281.8, 101568.8, 101738.3, 101775.3, 101672.2, 
    95593.84, 94996.94, 101776.6, 102039.3, 102062.1, 102152.5, 102205.5, 
    102324,
  100748.5, 101016.8, 101322, 101582.7, 101691.8, 101763.3, 101808.9, 
    101789.7, 101716.3, 102081.6, 102165, 102240, 102311.6, 102368.8, 102434.6,
  100781, 101089.9, 101395.2, 101614.1, 101714.8, 101780.1, 101836.9, 
    101980.2, 102124.8, 102192.1, 102302.1, 102390.4, 102440.9, 102477.5, 
    102509.4,
  100892.9, 101179.5, 101464.7, 101608.6, 101677.8, 101812, 101965.6, 
    102041.8, 102175.4, 102325.3, 102452.2, 102521.7, 102574.6, 102589.7, 
    102609.3,
  101026.3, 101309.2, 101542.1, 101661.1, 101811.3, 101966.1, 102106.9, 
    102251.9, 102402.2, 102499.4, 102587.4, 102646.7, 102675.3, 102682.1, 
    102689.4,
  101176, 101421.3, 101632.8, 101802, 101954, 102096.9, 102238.1, 102352.8, 
    102471.8, 102554.9, 102685.7, 102749.5, 102777.9, 102788, 102782.3,
  101513.7, 101430.7, 101355, 101275.9, 101219, 101205.9, 101267.4, 101365.9, 
    101487.3, 101269.4, 101423.7, 101789.9, 101741.9, 101446.4, 101405.3,
  101409.8, 101291.8, 101222, 101122.3, 101071.2, 101017.4, 101317.8, 
    101384.4, 101472.9, 101579.8, 101637.3, 101754.7, 101836.6, 100051.9, 
    100832.5,
  101339.4, 101231, 101159.6, 101102.6, 101010, 97744.6, 101291.7, 101565.1, 
    101573.4, 101616.6, 101637.4, 101683, 101788.4, 101883.7, 102013,
  101336.7, 101252.1, 101214.4, 101190.6, 101247.6, 101099.1, 97555.92, 
    101326.2, 101642.1, 101669.1, 101661.9, 101642.7, 101746.4, 101904.2, 
    102075.9,
  101452.1, 101410, 101391.5, 101432.3, 101465.7, 101484.2, 101321.6, 
    95377.35, 94701.55, 101519.2, 101706.7, 101651.7, 101754.6, 101879.4, 
    102124.8,
  101631.4, 101627.4, 101606.3, 101609.2, 101601.4, 101596.4, 101619.2, 
    101579.8, 101508, 101760.5, 101746, 101751.2, 101847.8, 102007, 102209.5,
  101832.6, 101827.8, 101799.1, 101794.9, 101783.6, 101795.6, 101794.3, 
    101853, 101882.4, 101852.5, 101872.2, 101908.6, 102002.4, 102161.6, 
    102345.7,
  102038.1, 102015.7, 101967.7, 101937.4, 101908.5, 101948.9, 101987.6, 
    101968.3, 101990.8, 102032.5, 102058.1, 102116.8, 102233.6, 102389.7, 
    102571.6,
  102218.5, 102221.6, 102196.9, 102201.7, 102197.4, 102214.1, 102218.2, 
    102244.8, 102250, 102250.3, 102283.3, 102362.3, 102472.1, 102612.4, 
    102766.1,
  102390.7, 102398.6, 102394.1, 102406.8, 102391.3, 102387.9, 102398.8, 
    102388.2, 102400.7, 102409.4, 102494.7, 102584.4, 102694.6, 102825.8, 
    102941.4,
  102995, 102890.4, 102770.2, 102607.6, 102415, 102257.3, 102100.7, 101944.3, 
    101785.3, 101283.7, 101203.3, 101347.4, 101111.6, 100747, 100720.5,
  103041.1, 102901.4, 102779.8, 102618.4, 102424.8, 102047.2, 102156.2, 
    101927.1, 101744.8, 101635.9, 101486, 101395.5, 101306.3, 99437.46, 
    100224.2,
  103041.8, 102921, 102792.8, 102687.1, 102341.9, 98667.38, 101952.4, 
    102094.6, 101888.5, 101719.5, 101550, 101476.3, 101426.2, 101447.3, 
    101515.1,
  103062, 102939.7, 102804, 102693, 102541.6, 102126.1, 98206.48, 101729.2, 
    101818, 101768.2, 101619.6, 101534.3, 101531.7, 101588.6, 101685,
  103115.7, 103015.9, 102875.7, 102750.7, 102632.2, 102465.6, 102093.6, 
    95761.34, 94963.41, 101562.4, 101685, 101578.5, 101610.6, 101653.1, 101836,
  103167.6, 103071.5, 102944.6, 102809.2, 102649.1, 102541.6, 102382.3, 
    102133.7, 101805.8, 101805.9, 101700.2, 101648.2, 101699.3, 101794.2, 
    101942.9,
  103218.5, 103154, 103043.4, 102934.8, 102770.8, 102667.1, 102499.9, 
    102340.8, 102129.6, 101901.5, 101782.6, 101766.2, 101810, 101930.3, 
    102062.9,
  103265.7, 103209.9, 103119.5, 103051.8, 102891.7, 102772.9, 102633.2, 
    102435.8, 102250.3, 102093.5, 101966.9, 101949.1, 102004.9, 102124.9, 
    102263.8,
  103312, 103276.6, 103219.1, 103190.4, 103111.1, 102982.2, 102804.5, 
    102658.4, 102498.9, 102356.9, 102247.3, 102228.3, 102273.1, 102374.9, 
    102493.1,
  103357.8, 103300, 103252.8, 103252.1, 103182, 103073.9, 102934.5, 102775.7, 
    102649.5, 102538.1, 102516.2, 102509.7, 102541.3, 102618.9, 102688.5,
  102993.3, 102893.6, 102819.4, 102699.9, 102574.2, 102449, 102239.4, 
    102065.3, 101910.5, 101356.9, 101272.2, 101376.9, 101106.2, 100631, 
    100474.5,
  102950.8, 102826.1, 102763.5, 102666.4, 102545.8, 102151, 102290.9, 
    101969.1, 101750, 101610.1, 101450.4, 101305, 101178.5, 99223.28, 99933.62,
  102890.1, 102765.7, 102724.7, 102672.1, 102393.3, 98795.66, 102013.3, 
    102201.7, 101924.4, 101660.6, 101429.6, 101296.5, 101179.5, 101175.5, 
    101177.9,
  102811, 102669.1, 102649.4, 102599.6, 102587.8, 102159.3, 98339.7, 
    101745.9, 101778.6, 101707, 101511.7, 101363.5, 101294.2, 101309.2, 
    101390.2,
  102725, 102603.6, 102592.5, 102574.1, 102585.4, 102527.9, 102174.1, 
    95848.83, 95120.89, 101603.3, 101699.4, 101516.9, 101496.6, 101478.6, 
    101644.3,
  102615, 102468.6, 102459.3, 102523.6, 102518.6, 102529.3, 102473.5, 
    102246.8, 101912.5, 101969.7, 101864.9, 101760.8, 101733, 101750.1, 101856,
  102495.1, 102377.7, 102327.2, 102467.4, 102517.6, 102570.3, 102510, 
    102485.8, 102367.5, 102175.7, 102067.2, 102020.7, 101994.9, 102037.7, 
    102112.1,
  102383.9, 102219.6, 102146.1, 102318.8, 102443.7, 102556.1, 102584.9, 
    102494.5, 102406.3, 102357.8, 102296.4, 102267.8, 102271.8, 102313.7, 
    102388.2,
  102270.2, 102099, 102014.2, 102137, 102376.2, 102552, 102639.6, 102667.7, 
    102642.8, 102574.2, 102521.3, 102512.1, 102522.8, 102565.3, 102618.1,
  102145.1, 101924.2, 101787.4, 101873.1, 102190.2, 102460.7, 102623.1, 
    102646.3, 102668.4, 102659.5, 102705.6, 102712.7, 102727.3, 102754.7, 
    102781.6,
  100784.8, 100619.3, 100791.2, 101068.8, 101226.3, 101339.8, 101268.6, 
    101227.3, 101121, 100661.1, 100658.5, 100930.5, 100860.7, 100522.3, 
    100430.6,
  100717.3, 100580.4, 100808.4, 101097.3, 101280.9, 101145.7, 101358.7, 
    101168.3, 100991.4, 100900.3, 100837.5, 100860.6, 100933.5, 99134.29, 
    99893.66,
  100671.7, 100582.6, 100844.6, 101171, 101154.8, 97799.48, 101188.7, 
    101386.2, 101219.8, 101022.7, 100897.6, 100917.7, 100987.6, 101101.3, 
    101119.3,
  100652.4, 100592.2, 100863.1, 101166.6, 101373.2, 101167.4, 97555.37, 
    101132.9, 101191.9, 101200.5, 101110, 101077.2, 101127.3, 101192.5, 
    101224.9,
  100662.5, 100646.4, 100894.3, 101229.5, 101439.1, 101565.4, 101354.7, 
    95193.13, 94676.02, 101191.2, 101361, 101248.5, 101283.8, 101249, 101334.6,
  100681.4, 100703.2, 100899.7, 101295, 101502, 101666.2, 101762.2, 101685.6, 
    101457.8, 101633.5, 101580.7, 101509, 101498.7, 101482.2, 101498.3,
  100715.5, 100789.2, 100966, 101386.2, 101640.7, 101855.2, 101901.9, 102007, 
    102014, 101912.7, 101836.6, 101802.5, 101755.7, 101744.7, 101722.5,
  100791.7, 100894.8, 101055.6, 101459.7, 101711.3, 101979.7, 102121.5, 
    102146, 102137.2, 102158.3, 102127, 102088.3, 102047.1, 102011.4, 101971.4,
  100888.3, 101016.2, 101205.4, 101589, 101898.5, 102180.4, 102332.5, 
    102437.8, 102473.1, 102444.3, 102406.3, 102365.4, 102320.3, 102261.1, 
    102190.5,
  101003.8, 101127.3, 101334.4, 101701.1, 102040.4, 102332.4, 102519.9, 
    102590, 102626.4, 102620.8, 102661.4, 102630.1, 102586, 102522.6, 102444.4,
  101131.3, 101248.4, 101319.2, 101301.3, 101275, 101197, 101041.9, 100955.8, 
    100951.9, 100590.8, 100693.3, 101038.4, 100978.4, 100690.9, 100663.4,
  101356.8, 101438, 101454.4, 101438.6, 101373.6, 101053, 101200.3, 100948.1, 
    100830.6, 100897.6, 100954.8, 101057.7, 101160.5, 99337.79, 100131.5,
  101564.2, 101643.1, 101629.7, 101613.4, 101305, 97832.73, 101082.3, 
    101276.5, 101121.6, 100975.8, 100953.6, 101039.6, 101146.6, 101257.2, 
    101329.5,
  101708.1, 101756.1, 101797, 101720.3, 101678, 101225.5, 97514.8, 100939.3, 
    100997.6, 101047.5, 100965.5, 100988.9, 101088.4, 101221.9, 101341.2,
  101888.2, 101925.9, 101970, 101933.4, 101857, 101762.1, 101369.6, 95125.34, 
    94435.27, 100866.4, 101022.3, 100905.8, 100988.5, 101052.5, 101249.3,
  102081.6, 102132.6, 102148.5, 102141, 102055.1, 101941.2, 101841.3, 
    101575.8, 101200.8, 101202.6, 101041.6, 100938.2, 100943.5, 100994.6, 
    101131.2,
  102275.1, 102340.4, 102351.4, 102348, 102295.8, 102222.8, 102045.9, 
    101926.4, 101730.5, 101422.2, 101144.7, 100996.8, 100929.4, 100958.4, 
    101039.3,
  102479.1, 102546.2, 102566.8, 102563.4, 102502.7, 102446.9, 102311.4, 
    102102.9, 101875, 101668.1, 101395.1, 101146.3, 101005.6, 100977, 101021.8,
  102714.3, 102805.8, 102856.4, 102881, 102846.9, 102749.7, 102586.1, 
    102431.4, 102222.6, 101968.7, 101702.7, 101413.9, 101181.9, 101070.6, 
    101057.6,
  102974.3, 103080.4, 103143.5, 103145.7, 103074.2, 102981.5, 102832.1, 
    102631.6, 102435.1, 102214.2, 102023, 101766.6, 101483.8, 101289.6, 
    101194.6,
  101960.2, 101882.1, 101798.4, 101624, 101521.4, 101410.7, 101241.8, 
    101153.7, 101141.1, 100756.9, 100792.4, 100993, 100739.6, 100295.6, 
    100144.7,
  102047, 101950.4, 101840.3, 101679.9, 101517.6, 101144.2, 101305.5, 101034, 
    100906.8, 101019.6, 101047.2, 101065.1, 100980.6, 99034, 99704.4,
  102088, 102026.5, 101925.6, 101812.9, 101421.1, 97868.3, 101026.8, 
    101279.4, 101074.1, 100996.1, 101032, 101094.3, 101081.4, 101070.5, 
    101021.2,
  102128.6, 102052.5, 101983.1, 101876.9, 101731.5, 101241.9, 97437.67, 
    100817.7, 100934.1, 100981.5, 100991.2, 101089, 101143.1, 101188.3, 
    101205.3,
  102242.6, 102174.2, 102095.1, 101986.7, 101862.9, 101703.6, 101264, 
    94993.97, 94232.23, 100747.7, 100990.8, 101040.1, 101181.4, 101218.9, 
    101339.3,
  102367.4, 102300.1, 102199.6, 102103.2, 101935.1, 101798.7, 101636.1, 
    101335, 100976.9, 100981.5, 100943, 101019.2, 101162.3, 101271.1, 101389.3,
  102507.4, 102473, 102364.6, 102258.2, 102117.9, 101971, 101739.4, 101590.8, 
    101387.6, 101103, 100951.3, 101019.9, 101116.8, 101260.5, 101395.8,
  102678.4, 102646, 102566.4, 102448.9, 102285.6, 102120.2, 101913.9, 
    101660.1, 101427.8, 101248.1, 101048.1, 100997.3, 101092.1, 101226.2, 
    101380.4,
  102854.6, 102858.2, 102803.8, 102731, 102583.1, 102366.6, 102097.2, 
    101889.4, 101672, 101431.9, 101219.9, 101040.4, 101055, 101175.8, 101312.4,
  103068.3, 103057.5, 103020.4, 102937.7, 102761.5, 102560, 102322.1, 
    102021.4, 101798.8, 101561.9, 101390.3, 101187.8, 101053.2, 101115.5, 
    101238.3,
  101794.4, 101803, 101802.1, 101736, 101716.1, 101686.7, 101574.7, 101518.4, 
    101466.3, 101059.9, 101125.1, 101401, 101229.1, 100770.2, 100576.8,
  101852.8, 101850.9, 101837, 101768.2, 101693.8, 101429.5, 101605.4, 
    101397.4, 101271.3, 101285.1, 101290, 101342.8, 101311.9, 99352.42, 
    99965.08,
  101852.9, 101910.2, 101896.3, 101870.1, 101578.6, 98006.1, 101298.7, 
    101542.3, 101318.6, 101215.5, 101183.4, 101251.3, 101238.7, 101215.4, 
    101100.8,
  101863.6, 101893.7, 101906.2, 101893.1, 101792.4, 101449.4, 97544.16, 
    101050.5, 101203.3, 101165.2, 101116.6, 101149.5, 101166.3, 101150.1, 
    101035.4,
  101958.7, 101979.9, 101973.5, 101942.7, 101869.6, 101734.7, 101401.9, 
    95071.4, 94260.88, 100906.9, 101084.6, 101073, 101109.4, 101055.7, 100990,
  102090.7, 102097.2, 102061.1, 102004.9, 101885, 101797.8, 101617.3, 
    101386.1, 101075.7, 101097.9, 101005.6, 101026.4, 101075.9, 101038.3, 
    100935.1,
  102225.1, 102245.4, 102203.6, 102134, 102016.2, 101877, 101670.8, 101525.2, 
    101333.4, 101085.6, 100966.7, 101031.3, 101067.1, 101042.7, 100936.9,
  102394.7, 102399.6, 102374, 102301, 102169.6, 102015.2, 101783.5, 101544.7, 
    101340.9, 101160.4, 101026.6, 101027.6, 101079.1, 101074.2, 100999.6,
  102543.7, 102591, 102583, 102536, 102425, 102214.2, 101953.2, 101728.1, 
    101518.1, 101281.5, 101103.4, 101024.1, 101090.8, 101098.5, 101052.8,
  102723.1, 102767.2, 102765.3, 102712.7, 102563.5, 102391.3, 102161.1, 
    101879.1, 101651, 101419.6, 101232.6, 101087.1, 101080.3, 101138, 101120.3,
  101878.3, 101892.4, 101894.5, 101875.5, 101876.3, 101850, 101789.6, 
    101793.2, 101795.4, 101425.1, 101493.8, 101791.2, 101668.8, 101261.3, 
    101130.5,
  102054.4, 102042.8, 102006.8, 101960.6, 101902.1, 101686.5, 101863.7, 
    101734, 101660, 101683.2, 101672.3, 101722.4, 101731.3, 99830.93, 100503.6,
  102150.1, 102143.5, 102119.3, 102072.4, 101816.6, 98227.12, 101631.6, 
    101859.3, 101701.1, 101616.1, 101546.7, 101580.1, 101615, 101657.3, 
    101673.7,
  102100.2, 102113.4, 102133.9, 102117.8, 102015.4, 101702.5, 97798.24, 
    101396.4, 101562.3, 101529.3, 101451.6, 101429.8, 101463.6, 101541.6, 
    101580.8,
  102139.5, 102168.7, 102150, 102149.8, 102079.8, 101966.8, 101667.3, 
    95348.98, 94539.79, 101253.1, 101417.4, 101341.1, 101361.2, 101367, 
    101453.4,
  102201.7, 102210, 102177.8, 102152.8, 102063, 101999.6, 101862.5, 101664.7, 
    101396.8, 101456.6, 101347.4, 101273.2, 101269, 101279.4, 101317.6,
  102233.7, 102252.2, 102221.3, 102187.3, 102112.2, 102041.7, 101887.8, 
    101770.5, 101618.9, 101438.2, 101312.6, 101236.4, 101201, 101190.7, 
    101182.6,
  102273.2, 102272.2, 102241.5, 102201.7, 102124.3, 102046.5, 101902.1, 
    101714.9, 101570.2, 101446.8, 101322.3, 101204.8, 101133.9, 101092.8, 
    101042.2,
  102268.1, 102304.6, 102284.5, 102249.5, 102188, 102051.6, 101892.4, 
    101736.2, 101589.9, 101433.5, 101299.8, 101160.4, 101048, 100963, 100873.2,
  102261, 102272, 102247.2, 102204, 102077.9, 101951.9, 101814.3, 101621.8, 
    101487.2, 101350.5, 101267.5, 101123.5, 100975.8, 100869, 100749.2,
  102316.9, 102321.1, 102323.6, 102298.4, 102292.6, 102241.7, 102164.5, 
    102126.4, 102048.2, 101588.9, 101556.4, 101751.9, 101495.5, 100996.5, 
    100793.6,
  102420.4, 102381.9, 102340.8, 102285.9, 102209, 101962.8, 102120.1, 
    101950.9, 101861, 101858.1, 101797.3, 101755.8, 101696.3, 99694.81, 
    100316.1,
  102395.2, 102357, 102300.9, 102238, 102000.5, 98420.38, 101727.5, 101992.4, 
    101853, 101709.5, 101630.8, 101619.7, 101606.5, 101594.3, 101572,
  102219, 102140.9, 102047.8, 101968.3, 101888.6, 101593.1, 97800.76, 
    101203.5, 101449.8, 101477, 101430.7, 101374.6, 101409.4, 101451.3, 101503,
  102097.5, 101972.5, 101810.9, 101696.5, 101588.3, 101496.6, 101257.8, 
    95175.62, 94284.15, 100820.8, 101147.9, 101064, 101140.3, 101166.5, 
    101310.7,
  101961.9, 101767, 101574.8, 101437.3, 101284, 101200, 101110.6, 100921.8, 
    100686.7, 100841.9, 100795.6, 100769.9, 100835.5, 100913.8, 101053.3,
  101762.6, 101570.4, 101390.2, 101272.4, 101125, 100993.6, 100869.2, 100774, 
    100655.6, 100517.8, 100489.8, 100497.8, 100532, 100625.9, 100783.2,
  101581.3, 101410.5, 101279.7, 101119.5, 100960.8, 100822.3, 100669.8, 
    100473.7, 100313.8, 100236.4, 100191.4, 100198.5, 100269.6, 100379.7, 
    100564.8,
  101463, 101355.2, 101220.2, 101070.6, 100945.4, 100750.2, 100545.8, 
    100318.2, 100102.8, 99926.14, 99862.53, 99886.95, 99989.45, 100136, 
    100336.9,
  101419.5, 101288.5, 101149.6, 100997.5, 100818.2, 100626.7, 100426.2, 
    100105.7, 99818.39, 99604.1, 99558.98, 99591.7, 99719.71, 99930.47, 
    100170.8,
  102573.1, 102452.2, 102311.4, 102168, 102085, 102024.8, 102014.6, 102068.4, 
    102099.8, 101739.7, 101816.2, 102115, 101989.4, 101562.3, 101415.1,
  102527.9, 102377.4, 102200.7, 102034.9, 101888.1, 101639.2, 101840, 
    101780.7, 101794.9, 101905.7, 101919.2, 101972.7, 101996, 100102.6, 
    100733.4,
  102417.9, 102253, 102033.9, 101842.2, 101550.4, 98087.77, 101347.6, 
    101708.2, 101604.1, 101573.4, 101601.3, 101654.3, 101689.4, 101715.6, 
    101731.5,
  102276.5, 102056.6, 101780, 101559.1, 101413.7, 101156.8, 97565.23, 101014, 
    101363.8, 101436.6, 101387.5, 101347.8, 101378.1, 101417.3, 101452.6,
  102112.1, 101828, 101559.6, 101357.2, 101349.3, 101317.8, 101133.4, 
    95172.78, 94312.09, 100910.3, 101218.4, 101076.8, 101095.6, 101040.8, 
    101120.3,
  101852.1, 101558.9, 101322.9, 101286, 101233.7, 101230.1, 101197, 101035.7, 
    100895.2, 101088.7, 100984.4, 100891.5, 100846.2, 100771.8, 100775,
  101605, 101375.9, 101280.4, 101238.3, 101182.5, 101120.8, 101094, 101122.6, 
    101018.5, 100820, 100709, 100604.3, 100513.6, 100451.2, 100434.7,
  101457.2, 101331.4, 101231.2, 101191.1, 101129, 101175.6, 101139.6, 
    100956.3, 100777.5, 100605, 100397.3, 100216.4, 100108.4, 100058.2, 
    100065.8,
  101428.5, 101326.6, 101280.7, 101269.5, 101308.1, 101256.1, 101113.4, 
    100916.8, 100628.9, 100294.6, 100042.7, 99860.57, 99745.89, 99702.35, 
    99712.34,
  101441.6, 101366.6, 101331, 101356.2, 101328.9, 101254.8, 101071.7, 
    100743.9, 100404.2, 100076.1, 99817.3, 99595.04, 99477.29, 99454.16, 
    99471.2,
  103096.3, 103029.8, 102918.4, 102719, 102504.8, 102271.1, 102073.9, 
    102014.1, 101974.1, 101542.2, 101513.7, 101702.9, 101479.3, 100963.8, 
    100753.7,
  102980.9, 102873.2, 102713.1, 102501.5, 102253.4, 101855.5, 101954.9, 
    101837.4, 101744.5, 101787.5, 101710, 101669.8, 101596.2, 99641.89, 
    100233.9,
  102760.3, 102654.1, 102447.8, 102254.9, 101907.3, 98397.59, 101647, 
    101986.3, 101800.4, 101698, 101607.3, 101565.6, 101503.8, 101460, 101386.3,
  102558.5, 102394, 102168.5, 101985.8, 101883.3, 101709.6, 98025.77, 
    101373.7, 101650, 101694.6, 101581.1, 101470.8, 101430.1, 101387.9, 
    101350.8,
  102327.3, 102141.8, 101954.3, 101901.4, 102073.4, 102040.2, 101760.5, 
    95576.6, 94687.64, 101295.2, 101520.4, 101322.7, 101291, 101188.3, 
    101204.7,
  102079.9, 101894.4, 101819.5, 102037.6, 102020.9, 102065.8, 102007.4, 
    101741.9, 101514.4, 101605, 101419, 101259.7, 101176.1, 101068.6, 101035,
  101856.8, 101806.1, 101976.3, 102035.7, 102024.2, 102021.6, 101950.8, 
    101891.6, 101697.8, 101431.3, 101283.5, 101152.3, 101031.2, 100919.8, 
    100858.5,
  101793.5, 101952.6, 101953.1, 101993.4, 101990.5, 101988.3, 101858.1, 
    101621.2, 101420.9, 101286, 101124.8, 100975.8, 100839.5, 100702, 100606.1,
  101894.6, 101993.4, 102073.9, 102108.3, 102081.8, 101944.7, 101755, 
    101566.1, 101331, 101104.1, 100947, 100804.8, 100621.4, 100431, 100286.4,
  101988.1, 102099, 102136.6, 102105.2, 101986.8, 101843.8, 101627.8, 
    101355.8, 101126.2, 100988.2, 100851.8, 100665.1, 100419.8, 100189.1, 
    100023.5,
  102899.8, 103061.4, 103223, 103306.5, 103361, 103331, 103221.9, 103161.7, 
    103128.2, 102727, 102746.2, 102958.6, 102707.6, 102088.7, 101775.2,
  102803.3, 102932.6, 103061.1, 103138.9, 103132.2, 102912.2, 103052.4, 
    102927.5, 102874.7, 102976.7, 102941.8, 102904, 102773.3, 100666.5, 
    101124.3,
  102640.7, 102783.4, 102870.1, 102942.4, 102803.8, 99338.18, 102617.6, 
    103041.4, 102934.2, 102868.4, 102783.7, 102748.6, 102605.3, 102462.7, 
    102260.5,
  102478.4, 102576.1, 102634.5, 102667, 102662.1, 102463.1, 98830.02, 
    102367.7, 102708.8, 102768.3, 102675.1, 102537.4, 102441.5, 102305.4, 
    102112.7,
  102303.5, 102372.4, 102413, 102413.9, 102528.7, 102558.3, 102451.1, 
    96426.16, 95552.62, 102243.5, 102533.2, 102332.4, 102249, 102048.4, 
    101941.6,
  102149.7, 102177.8, 102180.6, 102264, 102329.5, 102450.9, 102508.2, 
    102389.1, 102305.7, 102490.4, 102345.9, 102175.7, 102043.1, 101850, 
    101717.4,
  101942.6, 101967.3, 102018.2, 102129.9, 102218.6, 102284.4, 102403.1, 
    102522.1, 102449.8, 102253.2, 102127.4, 101979.1, 101807.1, 101636.5, 
    101469.1,
  101750.4, 101779.5, 101873.1, 102008.1, 102130.5, 102330.6, 102388.8, 
    102302.1, 102197.3, 102106.5, 101953.7, 101792.9, 101636.3, 101451.4, 
    101255.2,
  101478.2, 101625.3, 101804.9, 102002.7, 102198.7, 102295.3, 102311.2, 
    102265.5, 102113.9, 101917.1, 101788.6, 101660.6, 101465.4, 101245.6, 
    101017.7,
  101399.7, 101560.1, 101783.5, 102036.9, 102198.8, 102262.1, 102235.1, 
    102067.3, 101917.3, 101809.5, 101708, 101533.4, 101308.3, 101056.1, 
    100796.4,
  101241.6, 101374.2, 101564.4, 101786.9, 102040.8, 102277.1, 102508.2, 
    102768.7, 102980.8, 102774.1, 102943.7, 103278.9, 103167.7, 102773.3, 
    102617.8,
  101209.9, 101314.7, 101483, 101716.6, 101929.1, 102030.6, 102428.5, 
    102593.8, 102759.5, 102957.6, 103047.8, 103148.8, 103195.5, 101276.4, 
    101886.6,
  101123.2, 101250.6, 101413.2, 101654.7, 101731.5, 98556.63, 102098.1, 
    102591.7, 102651.1, 102748, 102834.6, 102937.3, 102975.8, 102975.3, 
    102952.8,
  101004.6, 101110.7, 101286.4, 101494.1, 101754.7, 101653.9, 98304.05, 
    101959.5, 102441.5, 102563.2, 102651.5, 102685.1, 102757.6, 102783.2, 
    102757.5,
  100874.2, 100970.8, 101124.7, 101338.7, 101584.7, 101826.6, 101748.2, 
    96050.26, 95366.6, 101980.1, 102412.3, 102407.4, 102486.9, 102490.7, 
    102512.5,
  100760.7, 100830.8, 100954.8, 101152.9, 101382.6, 101573.5, 101802.6, 
    101763.2, 101764.6, 102123.1, 102191, 102228.9, 102293.4, 102282.3, 
    102300.2,
  100645, 100721.5, 100839.1, 100994.4, 101217.2, 101397.4, 101558.6, 
    101763.4, 101904.1, 101944.7, 102038.9, 102098.1, 102118.5, 102111.9, 
    102077.6,
  100546.4, 100630.4, 100722, 100866.9, 101015.5, 101208.9, 101380, 101515.4, 
    101687.4, 101867.8, 101969.9, 102008.4, 102016.4, 101964.2, 101878.5,
  100468.5, 100576.6, 100667.7, 100786, 100917.7, 101083.5, 101303.3, 
    101538.8, 101718.6, 101818.5, 101902.9, 101924.2, 101878.8, 101760, 
    101605.3,
  100458.9, 100511.2, 100600.4, 100712.4, 100873.3, 101131.4, 101397.5, 
    101592.5, 101748.3, 101824.2, 101885.5, 101841.3, 101720.6, 101538.7, 
    101325,
  100144.7, 100066.2, 100019, 100011, 100073.8, 100144.7, 100249.9, 100405.8, 
    100593.5, 100463.5, 100740.6, 101254.5, 101350.4, 101201.7, 101263,
  99958.05, 99868.05, 99813.88, 99808.32, 99834.05, 99798.5, 100085.8, 
    100224.2, 100393.3, 100639.6, 100848.9, 101136.2, 101372.6, 99744.09, 
    100561.1,
  99759.93, 99682.14, 99641.36, 99636.18, 99588.66, 96335.98, 99813.62, 
    100190.9, 100343.7, 100535.7, 100744.1, 100985, 101240.1, 101403, 101588.3,
  99646.67, 99571.98, 99523.55, 99502.38, 99624.27, 99477.45, 96115.05, 
    99798.2, 100240.4, 100451.1, 100654.4, 100834.6, 101083.7, 101316.1, 
    101496.3,
  99613.5, 99539.33, 99474.55, 99506.48, 99607.18, 99772.2, 99667.76, 
    94028.91, 93503.78, 100123.1, 100599.7, 100716.2, 100931, 101073.3, 
    101280.6,
  99614.07, 99557.77, 99505.66, 99553.45, 99641.71, 99749.34, 99938.5, 
    99914.55, 99903.06, 100332.1, 100476.9, 100619.6, 100790.6, 100930.5, 
    101073,
  99662.62, 99601.98, 99587.6, 99636.2, 99763.59, 99871.59, 99983.58, 
    100190.6, 100313.6, 100347.2, 100461.8, 100591.3, 100693.6, 100794.3, 
    100887.2,
  99787.33, 99749.42, 99721.03, 99776.76, 99874.38, 100022.8, 100122.3, 
    100185.5, 100274.1, 100406.7, 100510, 100613.4, 100753.8, 100865.2, 
    100952.5,
  100004.3, 99972.62, 99983.42, 100034.5, 100127.6, 100231, 100336.5, 
    100476.6, 100590.1, 100689.4, 100789.4, 100897.6, 100980.6, 101023.8, 
    101028.5,
  100413.9, 100338.7, 100341.8, 100389.9, 100449.5, 100555.5, 100649.5, 
    100727.9, 100806.3, 100890, 100995.2, 101041.5, 101041.4, 101016.7, 
    100956.1,
  99718.15, 99544.93, 99386.27, 99254.33, 99151.25, 99079.59, 99033.12, 
    99051.94, 99101.71, 98839.81, 98937.69, 99223.94, 99083.79, 98698.29, 
    98564.96,
  99586.02, 99387.12, 99217.08, 99061.09, 98916.18, 98655.88, 98808.72, 
    98777.59, 98800.88, 98892.52, 98962.64, 99054.09, 99100.66, 97304.24, 
    97951.45,
  99519.84, 99330.91, 99139.87, 98987.45, 98700.44, 95250.13, 98437.59, 
    98636.88, 98621.94, 98684.96, 98768.86, 98870.46, 98962.3, 99005.02, 
    99026.72,
  99543.36, 99326.98, 99135.8, 98981.81, 98804.53, 98447.43, 94795.49, 
    98244.2, 98507.28, 98574.52, 98651.85, 98733.23, 98839.67, 98935.88, 
    99004.72,
  99612.8, 99440.51, 99271.69, 99110.98, 98943.03, 98761.86, 98469, 92553.81, 
    91902.12, 98333.32, 98622.27, 98655.82, 98761.45, 98809.05, 98944.25,
  99728.93, 99557.35, 99409.68, 99276.14, 99106.25, 98951.95, 98806.37, 
    98659.31, 98460.52, 98628.48, 98642.97, 98686.32, 98782.9, 98857.85, 
    98966.5,
  99875.9, 99735.62, 99605.55, 99502.14, 99384.52, 99256.45, 99100.58, 
    99015.1, 98930.94, 98860.95, 98861.91, 98893.84, 98931.48, 98986.92, 
    99054.59,
  100021.2, 99898.45, 99788.1, 99713.84, 99612.76, 99531.77, 99416.05, 
    99320.52, 99267.22, 99260.44, 99256.53, 99269.73, 99298.32, 99324.2, 
    99345.41,
  100121.3, 100048.7, 99989.24, 99964.14, 99915.6, 99830.69, 99750.09, 
    99716.78, 99679.15, 99653.88, 99642.59, 99638.16, 99625.88, 99616.07, 
    99593.48,
  100176.7, 100080, 100043, 100060.3, 100026.1, 99986.16, 99933.95, 99886.84, 
    99885.52, 99858.3, 99878.63, 99863.48, 99818.54, 99768.43, 99691.63,
  100345.3, 100349.6, 100344.3, 100302.4, 100252.2, 100121.8, 99954.83, 
    99804.43, 99627.25, 99094.61, 98975.74, 99086.52, 98835.13, 98373.87, 
    98213.29,
  100247.3, 100220.9, 100193.8, 100155.3, 100084, 99763.16, 99871.62, 
    99627.35, 99390.28, 99251.01, 99043.01, 98914.98, 98789.01, 96888.3, 
    97458.66,
  100084.6, 100071.2, 100034.5, 100044.3, 99856.62, 96372.05, 99512.57, 
    99680.38, 99399.4, 99206.36, 98968.92, 98837.63, 98692.59, 98601.48, 
    98486.73,
  99884.62, 99857.59, 99831.89, 99851.55, 99861.2, 99606.99, 95855.62, 
    99210.91, 99328.14, 99240.58, 99029.88, 98846.99, 98698.16, 98578.19, 
    98445.62,
  99645.6, 99655.91, 99664.03, 99706.85, 99780.41, 99776.52, 99545.99, 
    93408.88, 92605.99, 99068.01, 99134.05, 98920.9, 98776.85, 98589.57, 
    98470.22,
  99367.05, 99395.67, 99432.59, 99532.59, 99660.22, 99776.72, 99761.06, 
    99602.73, 99376.04, 99406.02, 99247.44, 99054.52, 98880.36, 98682.77, 
    98510.15,
  99062.37, 99142.97, 99211.62, 99409.9, 99691.26, 99821.96, 99820.59, 
    99811.56, 99715.32, 99545.5, 99379.89, 99213.3, 99024.25, 98830.42, 
    98622.69,
  98809.99, 98885.04, 99020.38, 99397.95, 99743.43, 99890.12, 99894.65, 
    99818.32, 99715.71, 99623.27, 99478.31, 99313.38, 99147.07, 98966.62, 
    98772.2,
  98696.07, 98852.63, 99091.67, 99575.16, 99855.05, 99999.58, 99969.59, 
    99940.53, 99828.59, 99698.62, 99548.95, 99414.37, 99253.37, 99083.89, 
    98893.84,
  98833.62, 98995.58, 99263.87, 99721.43, 99954.37, 100076.8, 100045.2, 
    99949.04, 99835.95, 99715.32, 99615.77, 99495.17, 99352.02, 99208.23, 
    99043.34,
  99604.79, 99669.52, 99771.48, 99907.05, 100073.8, 100218, 100361.2, 
    100541.2, 100694.1, 100484.1, 100640, 100963.4, 100825.7, 100378.5, 
    100171.9,
  99679.02, 99723.1, 99799.55, 99933.74, 100055, 100066.2, 100354.1, 
    100446.8, 100561.8, 100721, 100771.6, 100829.5, 100832.9, 98913.57, 
    99474.18,
  99664.61, 99763.02, 99846.4, 99983.12, 99963.34, 96723.54, 100112.9, 
    100459.7, 100464.7, 100524.3, 100588.4, 100651.5, 100646.3, 100613.7, 
    100546,
  99590.88, 99703.26, 99821.65, 99937.45, 100050.2, 99906.94, 96405.45, 
    99950.85, 100370.4, 100487.4, 100518.6, 100501.8, 100527.2, 100490.7, 
    100425.2,
  99487.64, 99625.45, 99737.3, 99855.75, 99954.07, 100015.8, 99897.9, 
    94136.86, 93465.88, 100170.7, 100526.3, 100437.1, 100455, 100355.4, 
    100331.7,
  99450.9, 99600.1, 99737.16, 99905.05, 100016.8, 100104.8, 100278.9, 
    100247.1, 100280.4, 100567.5, 100500.2, 100425.4, 100371.5, 100271.9, 
    100211.1,
  99709.87, 99888.94, 100072, 100259.3, 100409.8, 100511.3, 100587.8, 
    100693.8, 100630.8, 100491.8, 100436.4, 100361.3, 100277, 100202.3, 100098,
  100068.1, 100209.5, 100324.9, 100486.9, 100582.7, 100678.9, 100670.3, 
    100608.9, 100555.1, 100520, 100406.4, 100296.4, 100211.5, 100118.1, 
    100004.5,
  100474, 100594.6, 100691.8, 100814.5, 100885.7, 100866.4, 100811.3, 
    100749.6, 100608.9, 100436.3, 100295.4, 100183.4, 100068.4, 99983.34, 
    99885.11,
  100805.4, 100861.8, 100927.5, 100964.4, 100922.8, 100878.7, 100778.8, 
    100599.3, 100432.4, 100255.5, 100117.1, 99975.63, 99860.24, 99800.84, 
    99733.23,
  99173.34, 98975.45, 98718.85, 98462.74, 98324.17, 98393.62, 98588.52, 
    98821.27, 99100.14, 99065.85, 99433.98, 99972.32, 100103.9, 100018.8, 
    100145.7,
  99425.1, 99250.73, 99045.34, 98905.49, 98762.72, 98658.5, 98901.53, 
    99065.88, 99279.55, 99557.53, 99811.03, 100103.5, 100356.6, 98778.18, 
    99650.55,
  99647.46, 99544.47, 99420.17, 99354.98, 99096.95, 95879.43, 99275.27, 
    99506.33, 99621.23, 99791.9, 100011.3, 100249, 100479.2, 100662.3, 
    100869.2,
  99825.1, 99763.27, 99747.46, 99695.2, 99740.02, 99402.09, 96017.16, 
    99635.36, 100004, 100142.6, 100323.4, 100471.3, 100701.2, 100878.5, 
    101027.4,
  99960.44, 99966.95, 99984.84, 99986.49, 99979.23, 100033.8, 99785.63, 
    94044.05, 93586.66, 100269.6, 100637.4, 100726, 100900.4, 101007.6, 
    101171.6,
  100208.3, 100212.6, 100251.8, 100297.2, 100269.2, 100233.6, 100285.6, 
    100189.9, 100235.9, 100672.7, 100782.7, 100882.7, 101004.5, 101093.1, 
    101206.7,
  100383, 100432.7, 100479.3, 100533.6, 100562.5, 100586.6, 100570.7, 
    100703.1, 100780.4, 100757.6, 100823.8, 100895.5, 100944.9, 101004.3, 
    101072.3,
  100388.9, 100438.9, 100473.4, 100530.8, 100564, 100613.2, 100626.3, 
    100591.1, 100600.7, 100674.7, 100700.5, 100706.3, 100727.4, 100748.8, 
    100810.2,
  100309.9, 100356.7, 100396.6, 100439.8, 100515.3, 100549.9, 100550, 100575, 
    100548.4, 100469.3, 100405.9, 100365, 100338.5, 100343, 100408.4,
  100138.4, 100144.5, 100164.9, 100235.2, 100267.5, 100279.7, 100262.5, 
    100199.2, 100116.4, 100040.5, 100002.3, 99941.75, 99901.84, 99912.72, 
    99980.91,
  99628.99, 99280.81, 98792.82, 98169.91, 97688.3, 97585.23, 97618.05, 
    97756.98, 97953.55, 97916.98, 98292.29, 98869.37, 99022.64, 98907.68, 
    99003.14,
  99658.59, 99338.11, 98903.89, 98404.97, 97862.47, 97449.17, 97606.41, 
    97731.09, 97926.77, 98267.2, 98586.37, 98954.81, 99219.62, 97706.02, 
    98583.61,
  99685.2, 99442.78, 99095.33, 98692.53, 98036.1, 94509.45, 97642.54, 
    97868.02, 98114.55, 98361.47, 98666.88, 98987.8, 99302.75, 99522.92, 
    99773.42,
  99699.66, 99524.8, 99282.97, 98947.37, 98594.66, 97904.73, 94396.41, 
    97827.02, 98187.62, 98438.17, 98743.39, 99014, 99332.12, 99625.31, 99901.6,
  99702.46, 99634.4, 99470.4, 99239.68, 98890.6, 98617.48, 98051.92, 
    92445.16, 92058.91, 98419.14, 98870.19, 99076.34, 99384.73, 99628.44, 
    99978.96,
  99603.48, 99597.41, 99526.23, 99458.88, 99254.47, 98992.16, 98843.98, 
    98566.48, 98422.28, 98830.09, 98995.38, 99215.75, 99487.02, 99767.95, 
    100102,
  99486.68, 99542.46, 99545.45, 99533.73, 99483.69, 99367.37, 99207.56, 
    99204.32, 99163.43, 99125.53, 99229.19, 99422.38, 99644.23, 99922.01, 
    100238.8,
  99254.53, 99294.92, 99316.93, 99395.7, 99481.91, 99548.98, 99504.42, 
    99384.08, 99317.62, 99398.98, 99496.34, 99649.52, 99865.72, 100137.5, 
    100457.9,
  99041.54, 99083.34, 99122.25, 99197.07, 99321.8, 99485.05, 99603.37, 
    99709.05, 99740.48, 99715.3, 99763.23, 99896.24, 100092.7, 100352.4, 
    100643,
  98761.51, 98749.85, 98762.46, 98849.41, 98982.41, 99245.55, 99490.27, 
    99627.16, 99711.61, 99790.62, 99933.72, 100085.5, 100284.8, 100541.1, 
    100786.9,
  99749.81, 99709.17, 99638.67, 99439.08, 99177.74, 98826.91, 98666.93, 
    98701.38, 98791.39, 98528.92, 98686.41, 99068.88, 99068.83, 98811.47, 
    98764.91,
  99609.87, 99564.35, 99506.28, 99309.78, 99052.8, 98492.97, 98664.09, 
    98698.77, 98740.72, 98823.66, 98962.48, 99139.53, 99254.06, 97565.2, 
    98316.09,
  99412.02, 99407.96, 99388.47, 99258.62, 98907.69, 95276.77, 98456.09, 
    98730.18, 98789.87, 98893.52, 99033.19, 99192.8, 99336.95, 99440.46, 
    99518.62,
  99269.59, 99264.38, 99278.27, 99185.44, 99037.35, 98545.91, 94879.89, 
    98504.04, 98766.79, 98938.59, 99119.02, 99246.2, 99391.34, 99552.8, 
    99656.8,
  99164.68, 99146.68, 99202.38, 99169.2, 99077.38, 98839.12, 98461.37, 
    92859.91, 92421.44, 98842.75, 99206.55, 99314.23, 99481.83, 99596.32, 
    99770.85,
  99142.52, 99090.25, 99109.05, 99116.62, 99079.93, 98932.78, 98719.12, 
    98725.28, 98663.41, 99119.7, 99246.48, 99418.25, 99568.5, 99728.12, 
    99889.33,
  99151.55, 99080.72, 99053.5, 99093.8, 99091.79, 99059.81, 98870.91, 
    98896.65, 99071.26, 99206.84, 99334.5, 99521.81, 99669.98, 99856.2, 100058,
  99219.38, 99098.79, 98994.23, 98977.18, 99000.95, 99105.88, 99029.88, 
    98964.46, 99044.45, 99234.55, 99421.59, 99607.04, 99798.22, 100021.3, 
    100270.9,
  99354.97, 99194.66, 99025.1, 98935.98, 98947.66, 99087.47, 99120.97, 
    99152.64, 99230.41, 99331.6, 99483.36, 99682.39, 99907.9, 100166.3, 
    100439.7,
  99598.9, 99409.62, 99162.64, 98938.77, 98861.4, 99033.36, 99175.59, 
    99205.68, 99247.16, 99322.61, 99514.39, 99729.41, 99983.98, 100284.2, 
    100570.7,
  100239.9, 100064.4, 99898.19, 99760.26, 99619.79, 99532.1, 99438.38, 
    99425.12, 99457.43, 99149.86, 99225.01, 99503.94, 99417.86, 99140.75, 
    99147.92,
  100267.4, 100040.1, 99858.73, 99714.73, 99575.52, 99327.98, 99464.23, 
    99446.73, 99479.52, 99473.55, 99491.45, 99547.02, 99613.12, 97902.93, 
    98697.06,
  100306.2, 100039, 99830.62, 99709.47, 99457.76, 96011, 99288.86, 99527.98, 
    99494.55, 99488.72, 99521.34, 99580.91, 99693.44, 99805.52, 99931.07,
  100363.3, 100086, 99817.1, 99681.35, 99544.43, 99271.75, 95625.64, 
    99222.24, 99464.4, 99477.21, 99566.45, 99640.61, 99765.32, 99932.27, 
    100069.9,
  100389.6, 100166.5, 99873.86, 99677.97, 99529.3, 99437.57, 99225.75, 
    93439.75, 92801.37, 99300.2, 99616.86, 99713.68, 99855.05, 99987.67, 
    100181.8,
  100440.5, 100210.5, 99902.73, 99675.09, 99470.51, 99381.84, 99264.04, 
    99279.24, 99187, 99497.64, 99637.68, 99793.41, 99942.2, 100098.8, 100273.2,
  100472.1, 100261, 99954.3, 99700.19, 99466.27, 99347.32, 99258.48, 
    99331.34, 99420.27, 99533.88, 99689.66, 99869.39, 100021.5, 100203.9, 
    100508.7,
  100541.6, 100324.7, 99991.12, 99703.99, 99363.73, 99285.79, 99269.56, 
    99337.61, 99420.31, 99574.92, 99761.78, 99955.52, 100157.9, 100490, 
    100824.9,
  100618.1, 100414.2, 100113.6, 99834.21, 99428.6, 99310.9, 99301.18, 
    99410.68, 99520.72, 99676.33, 99862.97, 100088.9, 100397.4, 100756.8, 
    101060.3,
  100724.4, 100529.7, 100233.5, 99903.95, 99448.98, 99347.18, 99373.87, 
    99469.47, 99579.84, 99732.62, 99972.5, 100275.3, 100622.2, 100966.5, 
    101249.4,
  100733.2, 100595.3, 100434.8, 100289.3, 100081.2, 99834.8, 99755.99, 
    99699.46, 99569.23, 99094.99, 98994.99, 99070.63, 98776.02, 98227.48, 
    97982.35,
  100762.2, 100573.6, 100414.6, 100289.9, 100086.8, 99663.1, 99812.2, 
    99712.12, 99554.48, 99471.88, 99339.23, 99267.66, 99146.18, 97254.51, 
    97868.75,
  100808.6, 100573.2, 100411.1, 100330.5, 100003.7, 96432.97, 99636.4, 
    99838.62, 99692.72, 99556.56, 99468.72, 99430.99, 99416.2, 99410.31, 
    99390.1,
  100883.8, 100619.4, 100418, 100317.8, 100195.8, 99777.41, 96048.68, 
    99549.76, 99689.37, 99662.89, 99630.12, 99614.56, 99657.75, 99734.63, 
    99784.63,
  100977.3, 100738, 100504.9, 100370.2, 100218.8, 100087.8, 99768.13, 
    93815.21, 93188.87, 99624.8, 99834.2, 99827.45, 99927.88, 99991.83, 
    100164.2,
  101095.5, 100852.6, 100600, 100423, 100254.7, 100144.4, 100043.2, 99950.71, 
    99794.55, 100005.1, 100055.7, 100108.3, 100231.8, 100345.2, 100508.8,
  101213.2, 101026.5, 100763.9, 100538.5, 100364.1, 100291.3, 100201.5, 
    100220.6, 100254.6, 100265.6, 100317.9, 100422.9, 100554.1, 100709.1, 
    100864.2,
  101355.7, 101192.4, 100965.2, 100713.3, 100474.9, 100422.8, 100387.9, 
    100395.6, 100426.8, 100513.5, 100620.2, 100764.2, 100936.2, 101095.4, 
    101227.4,
  101495, 101384.2, 101190.1, 100991.8, 100708.1, 100592.7, 100573.2, 
    100635.5, 100710, 100806.2, 100929.1, 101089.7, 101248.5, 101381.9, 
    101489.7,
  101640.7, 101537.2, 101368.6, 101196.9, 100917.6, 100724.1, 100708.8, 
    100768.7, 100857.5, 100980.9, 101185.1, 101367.3, 101524.3, 101657.6, 
    101734.5,
  101889.1, 101750.5, 101578.8, 101345.3, 101168.2, 101036.1, 100844.5, 
    100672.8, 100479.7, 99918.52, 99758.91, 99748.3, 99376.19, 98806.06, 
    98591.52,
  101941.8, 101791.9, 101644.1, 101455, 101255.2, 100893.3, 101032.3, 
    100778.7, 100577.3, 100421.2, 100191.8, 99963.15, 99641.3, 97624.3, 
    98173.98,
  101972.8, 101835.3, 101720.1, 101607.6, 101226, 97703.26, 100950.9, 
    101113.9, 100901.6, 100689.9, 100457.2, 100250.6, 100007.9, 99798.18, 
    99606.74,
  101998.7, 101869.1, 101773.8, 101680, 101558.4, 101105.5, 97365.34, 
    100863.5, 100941.2, 100922.6, 100766.4, 100561.1, 100391.7, 100214.4, 
    100049.1,
  101998.4, 101921.5, 101839.4, 101777.2, 101665.9, 101547.1, 101189.7, 
    95035.88, 94411.24, 100940.2, 101078.6, 100885.8, 100775.2, 100600.3, 
    100537.5,
  101980.9, 101923.3, 101831.9, 101801.6, 101731.7, 101643.4, 101573.2, 
    101407.6, 101173.3, 101336.7, 101282.6, 101165.6, 101076.2, 100956.2, 
    100872.1,
  101937.5, 101947.4, 101845.4, 101796, 101775.1, 101759, 101661.6, 101657.5, 
    101624.4, 101538.2, 101461.4, 101395.9, 101303.2, 101221.5, 101129.2,
  101883.7, 101896.4, 101849.9, 101773.6, 101696.9, 101751.6, 101746.5, 
    101701.1, 101653.9, 101648.4, 101608.7, 101544.8, 101476.2, 101397.1, 
    101310.1,
  101807.1, 101856.8, 101833.3, 101802.3, 101708.1, 101678.7, 101713.7, 
    101752.5, 101775.1, 101747.4, 101703, 101651.1, 101586.4, 101510.8, 
    101411.6,
  101734.4, 101751.2, 101734.5, 101717.4, 101627.2, 101567.4, 101623.2, 
    101642.5, 101672.4, 101674.7, 101716.5, 101708, 101659.9, 101597.8, 
    101489.3,
  102163.1, 102092.1, 102009.6, 101894.9, 101801, 101709.4, 101543.6, 
    101457.4, 101331.4, 100806.9, 100702.3, 100765, 100428.7, 99858.77, 
    99620.54,
  102018.9, 101920.5, 101818.8, 101714.5, 101592.9, 101254.8, 101428, 101185, 
    101046.2, 101026.1, 100904.6, 100815.7, 100624.6, 98611.18, 99161.39,
  101883, 101770, 101656.9, 101581.7, 101329.2, 97838.8, 100905.3, 101286.4, 
    101036.2, 100883.4, 100803.8, 100780.5, 100692.4, 100591.3, 100471,
  101766.8, 101626.1, 101494, 101386, 101297.5, 100947.8, 97207.39, 100423, 
    100718.6, 100762.8, 100709, 100683.6, 100713.7, 100669.7, 100602.2,
  101662.7, 101525.5, 101384.2, 101254.2, 101173, 101023.4, 100738.6, 
    94658.74, 93736.16, 100209.3, 100565.7, 100526, 100667.5, 100669.3, 
    100723.6,
  101582.6, 101422.6, 101252, 101114.2, 100945.9, 100827.9, 100674.6, 
    100380.9, 100107.9, 100289.8, 100300.5, 100356.5, 100538.5, 100651.5, 
    100734.2,
  101527.7, 101366, 101201.6, 101025.1, 100869.7, 100651.6, 100423.4, 100243, 
    100072, 99948.88, 100001.1, 100146.8, 100368.2, 100566.4, 100691,
  101520.7, 101328.1, 101149.3, 100957.9, 100728.9, 100478.4, 100175.8, 
    99820.48, 99631.16, 99628.61, 99734.02, 99922.55, 100212.8, 100460.8, 
    100631.2,
  101540, 101373.6, 101207.7, 100987.1, 100766.1, 100416.4, 100022.2, 
    99638.88, 99414.4, 99348.87, 99480.64, 99759.73, 100086.6, 100361.3, 
    100541.8,
  101591.4, 101391.4, 101220.1, 100999.7, 100728.1, 100353.5, 99926.03, 
    99416.66, 99148.18, 99119.88, 99344.82, 99685.03, 100015.9, 100288.3, 
    100457,
  101657, 101472.5, 101274.5, 101022, 100782.8, 100494.4, 100163.6, 99906.59, 
    99683.83, 99105.18, 99037.57, 99274.81, 99146.79, 98818.51, 98821.62,
  101724.7, 101520.8, 101325.5, 101090.1, 100792.3, 100192.5, 100235.1, 
    99741.81, 99397.54, 99257.63, 99129.38, 99128.84, 99142.38, 97362.22, 
    98155.25,
  101786.9, 101587.3, 101395.7, 101218, 100712.6, 97031.34, 99821.85, 
    99987.37, 99552.23, 99232.87, 99047.67, 99017.08, 99005.9, 99097.33, 
    99263.02,
  101850.6, 101651, 101492, 101265.7, 100996.4, 100324.3, 96374.01, 99285.25, 
    99239.05, 99164.4, 99037.41, 98934.17, 98912.55, 99065.58, 99294.47,
  101917.6, 101756.8, 101618.9, 101390.5, 101109.1, 100734.4, 100084.3, 
    93727.1, 92784.12, 98941.44, 99112.43, 98939.63, 98942.84, 99094.54, 
    99406.36,
  101959.9, 101824.6, 101681.3, 101491.7, 101171.1, 100808.1, 100425.9, 
    99885.48, 99356.2, 99307.59, 99219.16, 99109.55, 99142.59, 99322.4, 
    99541.03,
  101991.7, 101911.7, 101785.8, 101603, 101358.3, 100982.9, 100530.2, 
    100164.3, 99817.88, 99513.64, 99412.6, 99358.41, 99401.88, 99575.44, 
    99727.7,
  101994, 101926.6, 101833.4, 101687.9, 101422.4, 101114.2, 100744.8, 
    100320.7, 99981.18, 99775.76, 99669.03, 99634.48, 99706.01, 99846.89, 
    99966.73,
  101979.9, 101956.1, 101901.1, 101801.9, 101601.5, 101285.5, 100939, 
    100634.2, 100356.4, 100104.3, 99957.28, 99926.01, 99973.6, 100063.7, 
    100130.6,
  101942, 101894.5, 101836.1, 101737.7, 101565.2, 101362, 101121.3, 100805.5, 
    100559.7, 100365.7, 100282.3, 100223.6, 100219.2, 100245, 100253.9,
  102326.8, 102224.4, 102110.1, 101919.7, 101756.7, 101567.4, 101324, 101141, 
    100941.5, 100331.8, 100201.1, 100309.1, 100058.6, 99508.04, 99277.77,
  102219.1, 102105.2, 101989.6, 101843.8, 101665.7, 101215, 101356.6, 
    101021.1, 100811.2, 100701.8, 100512.5, 100358.8, 100184.6, 98168.05, 
    98725.2,
  102063.1, 101950.1, 101820.8, 101740.9, 101414.3, 97921.68, 100944.6, 
    101262.3, 101030.4, 100768.8, 100560.5, 100406.6, 100227.2, 100091.2, 
    99929.68,
  101900.9, 101772, 101640.1, 101523.1, 101422.7, 101052.5, 97336.37, 
    100560.7, 100694.1, 100773.2, 100631.4, 100454.9, 100309, 100159.8, 
    100033.8,
  101706.8, 101584.9, 101452.2, 101331.6, 101225.9, 101134.9, 100867.2, 
    94849.33, 94044.93, 100404.6, 100668.8, 100496, 100418.2, 100240.3, 
    100162.7,
  101499.8, 101362.2, 101198.3, 101097.8, 100966.4, 100876.5, 100824.5, 
    100645.5, 100408.3, 100604.9, 100572.4, 100504.3, 100457.8, 100352.6, 
    100263.1,
  101275.1, 101131.6, 100964.1, 100847.1, 100743.5, 100648.1, 100542.9, 
    100539, 100512.9, 100431.1, 100423.6, 100457.2, 100438.9, 100400.6, 100331,
  101052.9, 100872.7, 100687.9, 100571.2, 100428.4, 100334.5, 100253.4, 
    100150.3, 100101.6, 100158.4, 100254.2, 100335.7, 100382.5, 100380.4, 
    100340.1,
  100831.6, 100644.8, 100465, 100315.6, 100183.2, 100062.4, 99959.11, 
    99922.22, 99912.92, 99921.45, 100029.3, 100199.1, 100297.7, 100327.2, 
    100298.3,
  100620.2, 100390, 100196.4, 100043.2, 99881.65, 99752.86, 99657.94, 
    99566.17, 99531.73, 99598.3, 99833.2, 100067.9, 100201.3, 100256.2, 
    100225.6,
  101018.9, 100754.7, 100509.8, 100285.5, 100156.8, 100066, 99984.39, 
    99975.69, 100017.5, 99763.44, 99913.73, 100267.6, 100217, 99882.55, 
    99782.63,
  100937.5, 100633.7, 100377.3, 100130.4, 99963.35, 99665.53, 99807.94, 
    99670.88, 99650.79, 99741.48, 99852.88, 100003.2, 100134.2, 98377.96, 
    99063.98,
  100864.2, 100564.9, 100297.5, 100069.7, 99748.23, 96372.34, 99425.54, 
    99613.94, 99500.84, 99479.61, 99533.98, 99682.08, 99845.37, 99977.53, 
    100078.8,
  100814.2, 100517.8, 100249.7, 100004.8, 99819.09, 99465.83, 95854.77, 
    99064.92, 99246.73, 99264.59, 99279.29, 99363.82, 99552.49, 99765.24, 
    99942.08,
  100786.2, 100509.7, 100245.6, 100008.8, 99820.76, 99653.97, 99341.14, 
    93524.52, 92732.95, 98838.71, 99047.31, 99053.6, 99233.66, 99465.58, 
    99756.18,
  100770.5, 100502.8, 100244.5, 100031.2, 99805.71, 99647.74, 99465.11, 
    99233.49, 98942.67, 98963.41, 98830.91, 98805.58, 98965.77, 99238.12, 
    99596.93,
  100769.6, 100533.3, 100293.1, 100095.2, 99899.88, 99695.84, 99481.64, 
    99305.39, 99081.16, 98827.99, 98654.52, 98601.86, 98755.21, 99108.8, 
    99528.49,
  100793.9, 100561.2, 100341.9, 100168, 99952.86, 99762.96, 99531.97, 
    99294.91, 99058.62, 98842.13, 98607.13, 98530.6, 98771.86, 99223.94, 
    99602.98,
  100819.9, 100615.8, 100430.6, 100285.9, 100099.6, 99881.69, 99648.54, 
    99438.41, 99200.8, 98960.71, 98773.31, 98798.84, 99143.93, 99466.59, 
    99735.27,
  100829.4, 100613, 100444.1, 100326.9, 100154.1, 99974.91, 99773.97, 
    99545.69, 99341.46, 99165.05, 99113.8, 99245.86, 99472.19, 99696.32, 
    99878.84,
  101164.9, 100942.8, 100734.9, 100534.1, 100402.7, 100268, 100140.7, 
    99998.65, 99868.95, 99401.41, 99368.71, 99584.41, 99520.69, 99286.52, 
    99309.2,
  101122.8, 100877.5, 100677.1, 100492.9, 100362.9, 100025, 100190.9, 
    99933.62, 99772.8, 99705.38, 99589.89, 99523.13, 99533.22, 97825.34, 
    98559.54,
  101053.6, 100809.9, 100615.6, 100472.7, 100217.2, 96818.66, 99922.05, 
    100144.5, 99956.29, 99772.02, 99577.2, 99455.42, 99386.95, 99447.02, 
    99541.53,
  100950.4, 100714, 100529.9, 100382.5, 100311.4, 100022.6, 96369.07, 
    99679.14, 99783.12, 99797.88, 99582.39, 99370.24, 99251.58, 99264.66, 
    99378.16,
  100830.6, 100609.4, 100432.9, 100298.9, 100239.7, 100212.4, 100004.8, 
    94022.12, 93281.91, 99553.68, 99578.48, 99273.5, 99125.1, 99053.95, 
    99187.7,
  100687.9, 100461.6, 100274.1, 100165.5, 100079.9, 100074.3, 100101.8, 
    99972.66, 99755.8, 99821.41, 99563.45, 99248.85, 99016.19, 98927.27, 
    98998.06,
  100540.7, 100331.4, 100132.9, 100011.3, 99938.31, 99930.53, 99932.26, 
    100019, 100011.8, 99860.13, 99639.23, 99377.23, 99109.96, 98984.16, 
    99093.49,
  100402.4, 100167.8, 99941.62, 99810.96, 99709.89, 99724.83, 99760.26, 
    99798.61, 99827.91, 99856.28, 99780.97, 99646.14, 99528.43, 99472.82, 
    99515.12,
  100276, 100036.1, 99809.2, 99639.23, 99539.52, 99532.98, 99571.2, 99681.39, 
    99779.21, 99817.45, 99812.7, 99784.9, 99735.4, 99730.71, 99765.25,
  100146.4, 99864.02, 99618.2, 99430.02, 99306.25, 99301.17, 99361.16, 
    99415.28, 99503.05, 99603.47, 99734.13, 99808.19, 99841.64, 99880.14, 
    99896.62,
  100475.5, 100156.2, 99877.51, 99649.2, 99565.97, 99583.12, 99622.38, 
    99733.62, 99845.58, 99539.59, 99585.15, 99787.21, 99531.85, 99057.68, 
    98940.45,
  100489.2, 100125.8, 99849.9, 99611.38, 99486.87, 99309.33, 99562.84, 
    99582.66, 99673.59, 99780.01, 99786.2, 99771.79, 99682.86, 97777.17, 
    98400.09,
  100494.2, 100114.9, 99835.29, 99612.73, 99335.22, 96027.43, 99253.66, 
    99587.02, 99636.62, 99661.62, 99687.04, 99689.14, 99643.91, 99568.97, 
    99518.39,
  100484.1, 100107.8, 99817.4, 99583.98, 99427.27, 99144.46, 95618.81, 
    99091.96, 99440.06, 99537.48, 99578.82, 99561.15, 99543.93, 99484.67, 
    99475.74,
  100480.1, 100117.3, 99833.98, 99599.9, 99427.42, 99301.91, 99113.7, 
    93426.14, 92742.66, 99039.34, 99404.74, 99396.18, 99422.93, 99356.65, 
    99374.68,
  100476.1, 100107.3, 99819.47, 99607.77, 99405.75, 99271.2, 99172.45, 
    99080.19, 98964.21, 99189.22, 99238.46, 99272.77, 99314.59, 99276, 
    99248.76,
  100464.8, 100123, 99835.59, 99645.06, 99460.43, 99288.59, 99138.96, 
    99075.97, 99036.9, 99025.8, 99087.32, 99157.66, 99204.11, 99190.95, 99139,
  100439.5, 100100.2, 99815.25, 99667.88, 99484.36, 99319.91, 99148.48, 
    99010.55, 98936.35, 98949.51, 98989.04, 99041.59, 99097.38, 99155.92, 
    99146.55,
  100406.8, 100092.8, 99852.13, 99736.26, 99593.95, 99415.11, 99238.45, 
    99108.7, 98985.98, 98906.85, 98893.38, 98913.41, 98956.75, 99041.71, 
    99117.84,
  100353.6, 100031.6, 99820.07, 99743.3, 99648.55, 99504.57, 99348.91, 
    99171.45, 99029.67, 98902.6, 98847.23, 98812.14, 98818.74, 98911.5, 
    99031.14,
  100815, 100516.5, 100256.7, 100045.2, 99865.19, 99687.63, 99523.85, 
    99419.33, 99402.66, 99124.03, 99275.55, 99591.68, 99460, 99043.52, 
    98850.77,
  100833.6, 100507.9, 100271, 100089.5, 99905.95, 99486.11, 99580.57, 
    99323.32, 99275.43, 99323.7, 99398.06, 99503.23, 99571.48, 97736.17, 
    98340.09,
  100838.1, 100522, 100298.2, 100170.5, 99862.41, 96346.3, 99393.7, 99491.86, 
    99343.54, 99294.42, 99285.2, 99352.54, 99429.91, 99519.83, 99494.84,
  100823.7, 100544, 100331.4, 100215, 100107.7, 99701.76, 95924.55, 99176.17, 
    99356.84, 99357.62, 99260.58, 99211.17, 99253.12, 99373.69, 99456.99,
  100820.3, 100589, 100394, 100308.5, 100216.7, 100066.5, 99701.66, 93634.68, 
    92864.22, 99164.31, 99282.02, 99117.09, 99073.95, 99101.7, 99283.37,
  100817.6, 100615.8, 100444.2, 100392.5, 100289, 100189.6, 100002.2, 
    99796.11, 99526.34, 99541.98, 99362.16, 99185.2, 99061.81, 98981.91, 
    99071.02,
  100823.1, 100680.9, 100542.8, 100518.1, 100461.9, 100321.7, 100156.5, 
    100029, 99856.5, 99653.55, 99477.78, 99296.24, 99102.77, 98982.73, 98915.4,
  100846.6, 100742, 100640.8, 100652.1, 100552.1, 100453.2, 100273.1, 
    100097.6, 99934.31, 99799.69, 99628.89, 99423.47, 99210.34, 99007.72, 
    98885.8,
  100914.5, 100847.1, 100820.3, 100846.1, 100760, 100602.4, 100416.5, 
    100256.7, 100074.7, 99881.96, 99712.84, 99529.15, 99312.18, 99079.13, 
    98888.15,
  101010.2, 100937.2, 100927.1, 100935.8, 100824.9, 100705.7, 100522.7, 
    100301, 100104.8, 99918.98, 99778.77, 99604.08, 99384.16, 99165.95, 
    98927.91,
  101161.4, 101084.7, 100946.8, 100747.1, 100582.1, 100436.4, 100250.5, 
    100078, 99880.43, 99271.27, 99110.43, 99179.99, 98938.35, 98574.35, 
    98456.34,
  101225.4, 101110.9, 101011.5, 100850.6, 100675.7, 100308.1, 100446.4, 
    100153.5, 99971.92, 99824.39, 99561.51, 99346.99, 99173.44, 97298.11, 
    97923.45,
  101248.1, 101124.7, 101024.7, 100962.9, 100619.8, 97048.16, 100267.4, 
    100481.4, 100226.6, 100010, 99761.61, 99540.4, 99291.65, 99184.25, 
    99073.59,
  101273.7, 101145.2, 101035.5, 100966.3, 100850.9, 100469.9, 96615.33, 
    100003.1, 100111.7, 100100, 99908.81, 99675.12, 99445.84, 99246.95, 
    99132.95,
  101280.1, 101160.9, 101044.1, 100960.9, 100841.7, 100742.8, 100431, 
    94177.78, 93333.22, 99868.52, 100003, 99763.05, 99581.7, 99294.16, 
    99156.06,
  101282.5, 101144.2, 101004.7, 100922.8, 100776.3, 100692.1, 100550.5, 
    100312.4, 100036.8, 100104.6, 99976.52, 99802.56, 99625.59, 99418.19, 
    99179.38,
  101282.7, 101150.5, 100995.2, 100896.9, 100787.2, 100637.8, 100452.8, 
    100318.9, 100159.6, 99989.59, 99890.07, 99785.06, 99643.44, 99433.56, 
    99219.05,
  101302.5, 101140.2, 100961.8, 100868.7, 100702.4, 100541.4, 100335, 
    100117.1, 99942.94, 99855.04, 99785.55, 99720.45, 99629.32, 99459.9, 
    99262.19,
  101339.3, 101173.9, 101002.1, 100872.7, 100706.1, 100481.5, 100249.9, 
    100052.8, 99868.98, 99729.11, 99670.39, 99655.47, 99589.22, 99476.41, 
    99246.89,
  101392.3, 101174.9, 100978.4, 100807.2, 100595.3, 100385.3, 100152.4, 
    99887.36, 99689.92, 99576.47, 99571.98, 99579.91, 99549.19, 99478.59, 
    99294.3,
  100532.8, 100311.6, 100093.8, 99935.43, 99837.3, 99888.18, 100043.1, 
    100234, 100327.2, 99976.94, 99955.71, 100071.3, 99647.29, 99031.26, 
    98759.79,
  100387.9, 100114.4, 99891.88, 99733.23, 99649.9, 99568.93, 99972.3, 
    100090.9, 100182.5, 100293.2, 100255.5, 100204.8, 99986.2, 97919.91, 
    98416.81,
  100249.9, 99972.52, 99736.58, 99620.54, 99448.57, 96153.6, 99643.81, 
    100101.9, 100143, 100210.9, 100233.8, 100251.5, 100142.5, 99985.29, 
    99736.2,
  100142.9, 99890.7, 99644.52, 99546.5, 99495.04, 99345.32, 95848.87, 
    99550.61, 99986.4, 100093.9, 100184.6, 100221.5, 100224, 100106.1, 
    99942.02,
  100081.4, 99849.71, 99604.8, 99528.09, 99498.69, 99481.22, 99405.5, 
    93619.49, 92951.55, 99659.98, 100058.1, 100148.5, 100251.1, 100156.8, 
    100075.4,
  100073.5, 99839.84, 99610.98, 99523.63, 99440.41, 99470.55, 99492.55, 
    99493.78, 99476.76, 99798.38, 99913.01, 100075.5, 100220.8, 100222.4, 
    100139.5,
  100103.7, 99911.76, 99686.52, 99587.12, 99537.11, 99529.98, 99480.26, 
    99582.09, 99641.65, 99684.81, 99813.35, 100009.1, 100181.1, 100229.6, 
    100178.2,
  100184.1, 99997.3, 99781.19, 99675.5, 99510.77, 99465.66, 99462.02, 
    99466.08, 99524.43, 99637.27, 99755.18, 99949.62, 100156.3, 100238.4, 
    100203.8,
  100302.8, 100136.4, 99931.76, 99753.48, 99579.78, 99440.45, 99384.82, 
    99432.8, 99508.58, 99580.7, 99707.84, 99923.09, 100142.9, 100233.8, 
    100209.8,
  100435.8, 100257.2, 100030.1, 99806.41, 99547.79, 99381.07, 99325.55, 
    99312.88, 99411.2, 99521.43, 99721.03, 99951.33, 100158.1, 100245.8, 
    100222.6,
  100042.1, 99843.7, 99663.52, 99520.59, 99383.73, 99224.8, 99157.98, 
    99287.7, 99553.8, 99469.96, 99727.72, 100077, 99858.16, 99318.34, 99081.52,
  99983.04, 99736.91, 99534.47, 99370.73, 99172.22, 98875.58, 99052.34, 
    99217.07, 99505.92, 99831.58, 100022.5, 100131.7, 100016.4, 98015.77, 
    98593.77,
  99949.59, 99682.92, 99455.39, 99294.77, 98991.68, 95555.12, 99021.44, 
    99419.65, 99723.52, 99941.88, 100104.6, 100173.3, 100110.9, 99929.38, 
    99793.61,
  99960.95, 99709.32, 99477.59, 99334.65, 99259.23, 99022.02, 95487.15, 
    99342.36, 99815.83, 100055.8, 100193.4, 100209.5, 100147, 100009.9, 
    99913.45,
  100018.4, 99766.12, 99535.86, 99452.44, 99361.97, 99410.95, 99185.84, 
    93550.28, 93032.58, 99888.13, 100264, 100275.6, 100234.2, 100053.6, 
    100022.6,
  100134.4, 99871.83, 99627.85, 99501.23, 99417.57, 99443.57, 99499.82, 
    99542.98, 99605.16, 100146.7, 100274.1, 100348.4, 100298.4, 100173.6, 
    100094.9,
  100279.5, 100044.1, 99774.38, 99599.92, 99509.57, 99493.48, 99466.77, 
    99822.27, 100072.9, 100220.2, 100353.2, 100432.9, 100372.4, 100275.9, 
    100202.6,
  100475.8, 100284.6, 100025.8, 99807.95, 99609.9, 99612.45, 99693.69, 
    99881.83, 100090.4, 100337.4, 100467.8, 100524.1, 100482.1, 100410.8, 
    100365.6,
  100678.4, 100539.5, 100361.9, 100178.5, 100006.5, 99956.37, 100028.9, 
    100229.9, 100393.7, 100512.5, 100605.6, 100655.6, 100624.6, 100557.9, 
    100504.8,
  100888.5, 100770.5, 100607.7, 100455, 100313.9, 100285.3, 100334, 100406.1, 
    100518.2, 100623.9, 100751.6, 100805.1, 100790.4, 100729.1, 100659.1,
  100660.2, 100484.8, 100301.6, 100095.1, 99744.18, 99433.34, 99281.87, 
    99369.56, 99458.31, 99035.3, 99235.7, 99734.87, 99866.98, 99739.97, 
    99784.02,
  100636.7, 100460.3, 100299.4, 100076.8, 99683.41, 99122.26, 99201.33, 
    99271.98, 99362.91, 99404.37, 99617.53, 99899.87, 100153.4, 98512.91, 
    99321.3,
  100643, 100481.4, 100349, 100186.1, 99673.49, 95976.7, 99141.09, 99333.26, 
    99473.39, 99562.11, 99797.3, 100050.4, 100293.5, 100444.2, 100537,
  100669.1, 100543.4, 100446.5, 100293.9, 100062.9, 99558.91, 95814.96, 
    99423.2, 99618.73, 99795.65, 100011, 100180.2, 100358.2, 100489.8, 
    100598.7,
  100718.6, 100630, 100569.7, 100481.3, 100277.6, 100158, 99722.92, 93730.13, 
    93281.52, 99887.66, 100234.2, 100262.4, 100376.5, 100399.7, 100577.6,
  100808.1, 100713.7, 100666.4, 100635.1, 100492.2, 100370.2, 100332.9, 
    100159.2, 99991.84, 100302.4, 100317.3, 100321.4, 100333.3, 100376.7, 
    100512.2,
  100926.6, 100844.8, 100800.7, 100787.2, 100713.7, 100624.6, 100491.4, 
    100519.7, 100507.4, 100391, 100321.1, 100277.2, 100252.1, 100318.7, 
    100446.9,
  101093.2, 101038, 100970.7, 100945, 100866, 100790.6, 100688.2, 100543, 
    100421.1, 100378.7, 100272.8, 100204.5, 100209, 100323.6, 100457.5,
  101240.2, 101229.1, 101200.9, 101136.1, 101057.5, 100963.3, 100814.9, 
    100712.9, 100578.5, 100405.4, 100256.2, 100213.4, 100262.4, 100387.4, 
    100488.9,
  101392.4, 101389.9, 101330.2, 101285.5, 101187.9, 101096.3, 100962.6, 
    100759.2, 100580.1, 100431.7, 100381.3, 100366.2, 100408.3, 100494.7, 
    100542.2,
  101300.9, 101361.6, 101303.3, 101079.8, 100700.1, 100265.2, 99773.6, 
    99282.45, 98999.77, 98566.04, 98636.91, 98867.38, 98745.48, 98509.42, 
    98575.08,
  101313.5, 101387.3, 101308, 101111.5, 100735.8, 100102.7, 99971.18, 
    99465.13, 99135.13, 99021.12, 98947.04, 98962.75, 99007.96, 97389.71, 
    98227.61,
  101341.9, 101401.1, 101352.6, 101228.6, 100731.6, 97014.12, 100051.2, 
    99960.57, 99700.93, 99519.59, 99432.61, 99407.41, 99452.09, 99542.84, 
    99618.9,
  101417.1, 101433.6, 101422, 101280.9, 101102.6, 100512.6, 96679.07, 
    100028.6, 100021.7, 100016.7, 99942.16, 99892.66, 99909.09, 99935.16, 
    99951.54,
  101508.2, 101508.7, 101503.7, 101395.9, 101223.4, 101063.4, 100585.5, 
    94438.13, 93867.71, 100286.4, 100440, 100339.5, 100338.5, 100283.9, 
    100316.7,
  101618.7, 101591.6, 101544.9, 101474, 101312.7, 101146.7, 101074, 100863.6, 
    100597.1, 100742.4, 100706.3, 100646.4, 100631, 100604.4, 100596.5,
  101756.9, 101729.6, 101669.9, 101560.1, 101428.7, 101267.6, 101072.9, 
    101048.4, 101030.9, 100922.6, 100859.8, 100845.7, 100812.3, 100789.1, 
    100763.7,
  101897.3, 101866, 101797.9, 101677.4, 101464, 101291, 101109, 100951.6, 
    100868.1, 100893.5, 100901.7, 100895.4, 100889.3, 100885.9, 100858.7,
  102016.1, 102007, 101954.1, 101818.3, 101615.3, 101369, 101090.5, 100930.3, 
    100867.8, 100836.1, 100822.9, 100843.1, 100872.1, 100870, 100850.1,
  102124, 102113.7, 102035.5, 101913.7, 101712.6, 101488.1, 101205.8, 
    100914.4, 100736.1, 100665.7, 100698, 100738.2, 100787.3, 100827.2, 
    100839.3,
  102668.8, 102515.7, 102351.1, 102124.8, 101882.7, 101628.9, 101329.8, 
    100987.2, 100619.8, 99905.87, 99662.17, 99816.96, 99654.98, 99203.61, 
    99044.73,
  102649.4, 102491.4, 102345.9, 102166.3, 101910.3, 101432, 101442.4, 101059, 
    100712.2, 100422.3, 100057.3, 99857.95, 99896.32, 98011.88, 98688.66,
  102610.8, 102467.6, 102337.5, 102226.4, 101841.4, 98171.23, 101236.1, 
    101305.9, 100953.4, 100621.7, 100288.4, 99967.12, 99897.92, 100001.2, 
    99982.63,
  102574.5, 102448.7, 102332.1, 102209.8, 102034.9, 101569, 97634.19, 
    100843.7, 100838.9, 100735.3, 100496.5, 100169.3, 99869.98, 99982.94, 
    100076.2,
  102526.8, 102438.7, 102325.3, 102207, 102036.8, 101850.5, 101432.1, 
    95149.9, 94250.5, 100615.2, 100653, 100376.5, 100119.6, 99963.55, 100100.7,
  102465.6, 102393.1, 102277.7, 102164.2, 101987.9, 101808.2, 101587.5, 
    101267.4, 100880.5, 100889, 100750.9, 100526.1, 100271.1, 100094, 100096.4,
  102388.1, 102342.4, 102228, 102131.3, 101995.3, 101792.3, 101540.3, 
    101305.6, 101049.4, 100872.6, 100766.7, 100637.4, 100433.1, 100242.1, 
    100161.5,
  102290.4, 102210.1, 102117.4, 102053.1, 101919, 101754.4, 101516.5, 
    101200.7, 100939.5, 100817.8, 100768, 100670.1, 100543.4, 100382.5, 
    100287.1,
  102113.7, 102062.9, 102018.6, 101978.9, 101909, 101747.5, 101519.9, 
    101228.4, 100971.7, 100782.4, 100732.3, 100689.6, 100599.7, 100478.8, 
    100374.4,
  101910.9, 101876.5, 101868.2, 101880, 101807.3, 101713.1, 101521.8, 101203, 
    100916, 100703.4, 100683.3, 100665.4, 100606.8, 100533.9, 100452.9,
  102480.1, 102345.6, 102218.4, 102056.2, 101929.1, 101759.6, 101527.2, 
    101354.8, 101197.4, 100596.6, 100421, 100407.8, 100094.4, 99348.5, 
    98901.69,
  102255.9, 102103, 101985.3, 101836, 101708, 101313.3, 101431.6, 101207.7, 
    101043.3, 100889.5, 100659.1, 100466.6, 100291.8, 98195.65, 98571.84,
  102036.6, 101901.5, 101778, 101675.6, 101400.3, 97917.67, 100990.3, 
    101294.5, 101112.1, 100913.1, 100677, 100492.3, 100362.2, 100252, 99967.73,
  101846.4, 101728.7, 101609.8, 101471.5, 101334.5, 100981.2, 97340.35, 
    100794.1, 100982.4, 100891.2, 100720.5, 100502.7, 100396.9, 100347.5, 
    100220,
  101690.9, 101580, 101466.5, 101322.6, 101220.7, 101110, 100994.8, 94996.91, 
    94227.94, 100676.3, 100731.9, 100520.6, 100376.7, 100319, 100318.7,
  101573.5, 101453.1, 101335, 101218.8, 101118.5, 101131.3, 101200.1, 
    101077.2, 100850.5, 100892.5, 100719.4, 100529.8, 100331.2, 100243.7, 
    100235.6,
  101482.9, 101375.5, 101279.4, 101193.9, 101169.7, 101235, 101214.4, 101159, 
    101066.2, 100838, 100707, 100549, 100324.6, 100169.4, 100082.7,
  101423.5, 101317.8, 101251.6, 101214.5, 101243, 101278.7, 101222, 101052.3, 
    100915.3, 100797.3, 100698.1, 100552.7, 100339, 100164.7, 100012,
  101374.1, 101328, 101299.9, 101331.3, 101372.9, 101347.3, 101238.4, 
    101073.9, 100908.7, 100774.7, 100688.3, 100563.2, 100359.5, 100175.4, 
    100022.8,
  101361.6, 101340.3, 101338.8, 101366.5, 101379.6, 101375.3, 101253.5, 
    101020.6, 100824.4, 100709.7, 100680.9, 100565.7, 100378.3, 100202.6, 
    100074.9,
  101715.8, 101619.2, 101509.1, 101361, 101229.3, 101097.3, 100981.3, 
    100921.2, 100963, 100677.7, 100749.2, 100915.4, 100616.6, 99981.49, 
    99588.8,
  101673.1, 101559, 101467.2, 101343.3, 101223.4, 100884.1, 101042.7, 
    100899.3, 100913.4, 100998.3, 100955.5, 100883.4, 100694.1, 98639.79, 
    99058.79,
  101651.6, 101572.4, 101489.9, 101429.9, 101161.2, 97668.13, 100882, 
    101154.8, 101067.3, 101014, 100908.6, 100813.4, 100620, 100427, 100175.5,
  101650, 101599, 101537.7, 101506.8, 101422.4, 101084.8, 97317.83, 100780.2, 
    100976.4, 100995.2, 100867.7, 100724.8, 100532.1, 100334, 100111.7,
  101646.3, 101646.5, 101612.6, 101592.9, 101537.1, 101451.5, 101117.4, 
    94991.81, 94181.02, 100684.3, 100817.5, 100631.4, 100434, 100199.5, 
    100013.9,
  101624.7, 101644.6, 101611.2, 101609.4, 101521.1, 101460.7, 101338.2, 
    101089.9, 100808.8, 100882.5, 100719.4, 100540, 100324.9, 100086.8, 
    99905.42,
  101580, 101603, 101564.3, 101585.2, 101556.8, 101471.2, 101325.6, 101175.2, 
    100973.1, 100766.7, 100613.3, 100440, 100208.9, 99978.69, 99823.97,
  101535.3, 101511.2, 101455.3, 101481.1, 101471.2, 101459.3, 101314.6, 
    101071.4, 100846.9, 100709, 100543.1, 100351.7, 100122.5, 99927.75, 
    99820.34,
  101490.2, 101450.4, 101395.6, 101393.3, 101443.8, 101468, 101333.5, 
    101124.6, 100873.4, 100671.4, 100483, 100293.3, 100083.3, 99945.7, 
    99863.92,
  101459.9, 101379.2, 101310.8, 101283.2, 101365.8, 101460.2, 101342.9, 
    101075.7, 100824.8, 100621.2, 100467.1, 100301.1, 100135.1, 100045.2, 
    99980.63,
  101954.4, 101947.6, 101882.8, 101761.1, 101650.9, 101560.1, 101430.3, 
    101331.4, 101196.3, 100694.1, 100640.5, 100817.7, 100597.3, 100131.8, 
    99926.66,
  101936.7, 101882.1, 101805.4, 101683.6, 101557.3, 101254.4, 101450.6, 
    101212.8, 101039.5, 100968.1, 100843.5, 100774, 100675, 98721.66, 99259.05,
  101851.7, 101783.7, 101684.6, 101598.8, 101324.5, 97896.49, 101133.4, 
    101389.3, 101151.9, 100929, 100731.4, 100636.1, 100496.1, 100401.5, 
    100243.7,
  101737.4, 101668, 101565.6, 101448.1, 101369.6, 101151.6, 97483.35, 
    100824.8, 100895.8, 100840.9, 100629.3, 100466.5, 100300.4, 100153.3, 
    99967.55,
  101648.2, 101582.9, 101487.9, 101341, 101301.2, 101352.4, 101174.8, 
    95058.34, 94222.48, 100505, 100547.4, 100312.6, 100124.4, 99914.4, 
    99756.49,
  101583.6, 101520.5, 101412.6, 101273.1, 101266.1, 101337.3, 101332.5, 
    101098.5, 100733.8, 100689.3, 100455.5, 100209.4, 99968.98, 99723.79, 
    99524.2,
  101546.2, 101513, 101422.4, 101288.5, 101342.9, 101384.7, 101294.1, 
    101153.8, 100919.7, 100657.2, 100411.5, 100132.8, 99816.02, 99523.97, 
    99251.69,
  101527.8, 101515.2, 101454.9, 101347.7, 101389.1, 101419.2, 101297.3, 
    101069.4, 100870, 100697, 100443, 100129.7, 99767.49, 99411.98, 99061.11,
  101513.2, 101544.2, 101545.8, 101480.7, 101544.5, 101486, 101331.7, 
    101150.6, 100992.4, 100794.7, 100557.7, 100244.6, 99859.65, 99467.01, 
    99093.58,
  101506, 101536.4, 101565, 101558.2, 101610.7, 101520.8, 101368.1, 101162.7, 
    101033.6, 100887.6, 100724.6, 100446.6, 100084.4, 99714.72, 99339.08,
  101929.5, 101920.3, 101879.2, 101793.6, 101719, 101658.5, 101607.9, 
    101581.5, 101492.2, 100980.5, 100868.1, 100961.1, 100687.2, 100179.3, 
    99986.33,
  101919.8, 101912.5, 101889.5, 101816.4, 101731.4, 101476.8, 101696.4, 
    101485.1, 101307.1, 101189.1, 101014.2, 100858.7, 100694, 98729.49, 
    99323.62,
  101927.9, 101952, 101936.5, 101918.2, 101673, 98258.18, 101509.5, 101681.8, 
    101460.2, 101201.3, 100926.6, 100742.4, 100535.1, 100418.1, 100319,
  101934.8, 101984.2, 101995.4, 101975, 101945.4, 101631.9, 97886.84, 
    101238.7, 101188.8, 101144.8, 100874.2, 100612.3, 100380.9, 100215.2, 
    100128.7,
  101952, 102014.2, 102047.6, 102054, 102055.5, 101972.1, 101673.3, 95500.23, 
    94702.64, 100886.2, 100843.9, 100473.3, 100199.6, 99942.75, 99886.34,
  101932.8, 102033.3, 102067.6, 102108.9, 102073.1, 101997.4, 101902.7, 
    101660.2, 101281.6, 101152.7, 100806.7, 100405.8, 100051.7, 99743.14, 
    99577.85,
  101894.7, 102046.9, 102094.8, 102144.2, 102141.4, 102049.2, 101912.3, 
    101792.5, 101552, 101185.3, 100805, 100408.4, 100000.7, 99649.16, 99395.49,
  101874.2, 102041.1, 102095.9, 102161.5, 102127.5, 102065.9, 101956.7, 
    101767.9, 101509.5, 101224.7, 100875.8, 100474.5, 100052.2, 99661.1, 
    99351.98,
  101823.4, 101998.2, 102107.5, 102166.4, 102170, 102085.6, 101983.8, 
    101858.5, 101636.2, 101317.7, 100970.5, 100575.2, 100134.4, 99716.09, 
    99355.65,
  101774.1, 101910.6, 102046.3, 102101.5, 102109.1, 102061.2, 101982.9, 
    101835.4, 101629.7, 101350.3, 101063.7, 100694.9, 100246.9, 99806.58, 
    99410.66,
  102885.8, 102894, 102884.5, 102897.7, 102890.1, 102825.7, 102727.7, 
    102652.4, 102515.6, 101989.8, 101863.2, 101928.4, 101565.2, 100915, 
    100622.5,
  102888.4, 102890.2, 102891, 102880.4, 102849.1, 102604.7, 102739.8, 
    102530.4, 102370.2, 102277.9, 102104, 101937.2, 101700.5, 99602.21, 
    100059.2,
  102790.5, 102820.9, 102857.8, 102878, 102687, 99184.15, 102466.2, 102686.4, 
    102498.8, 102267.6, 102058.2, 101893.5, 101664.2, 101450.4, 101180.9,
  102613.5, 102668.4, 102725.9, 102764.3, 102762.9, 102495.8, 98740.24, 
    102113.2, 102193.5, 102200.3, 102011.5, 101803.6, 101594.5, 101372.6, 
    101108.4,
  102432.5, 102514.6, 102569.5, 102621.1, 102628.6, 102623.5, 102407.1, 
    96303.18, 95462.02, 101805.5, 101938.8, 101685.8, 101487.5, 101220.3, 
    101001.7,
  102294.8, 102349, 102378.6, 102435.3, 102432.8, 102432, 102404.9, 102219.2, 
    101930.8, 101977.8, 101782.2, 101563.2, 101342.6, 101086.5, 100827.1,
  102190.4, 102223.6, 102234.6, 102258.1, 102261.3, 102242.8, 102164.8, 
    102116.4, 101980.2, 101757.2, 101570, 101398.7, 101172, 100930.9, 100627.6,
  102095, 102098.6, 102065, 102086, 102046.3, 102009.2, 101922.9, 101786.8, 
    101632.3, 101518.5, 101374.3, 101213.9, 101020.6, 100779.7, 100469.1,
  102029.9, 102013.8, 101971.6, 101927.9, 101862.1, 101780.7, 101670.4, 
    101583.1, 101465.4, 101311.4, 101175.1, 101050, 100876.8, 100629.1, 
    100315.6,
  101991.6, 101905.2, 101801, 101716.1, 101603.7, 101497.4, 101410.8, 
    101286.8, 101178, 101066.7, 101011.8, 100916.6, 100752.3, 100504.9, 
    100202.7,
  102917.3, 102837.7, 102775.4, 102710.2, 102713.8, 102725.9, 102707.6, 
    102710, 102665.6, 102200.4, 102156.6, 102322.5, 102107.6, 101577.5, 
    101342.3,
  102672.1, 102573.4, 102528.6, 102492.8, 102505.8, 102329.9, 102566.8, 
    102444.8, 102352.5, 102320.5, 102232.3, 102191.3, 102151.7, 100204.6, 
    100783.2,
  102444.7, 102358.6, 102330, 102322.8, 102262.8, 98909.93, 102114.6, 
    102424.1, 102276.3, 102125.9, 102013.3, 101966.9, 101931.6, 101917.4, 
    101857,
  102272.4, 102204.5, 102182.2, 102187.2, 102194.3, 102018.3, 98398.41, 
    101700.1, 101859, 101836.5, 101755.8, 101666.9, 101641.9, 101642.4, 
    101656.3,
  102161.2, 102140.1, 102126.8, 102096.6, 102091.9, 102039, 101831.1, 
    95936.28, 95084.24, 101279.8, 101482.8, 101344.3, 101315.5, 101264.6, 
    101312.6,
  102117.2, 102084, 102036.3, 102011.9, 101900.9, 101823.6, 101713.8, 
    101517.7, 101254.4, 101324.7, 101187.9, 101070.3, 100999, 100939.9, 100948,
  102040.6, 102012.8, 101954.7, 101891.2, 101795.1, 101651, 101491.8, 
    101373.9, 101237, 101069.2, 100927.9, 100805.6, 100684.7, 100611.7, 
    100583.7,
  101940.1, 101897.3, 101824.5, 101743.5, 101588.1, 101458.6, 101309.5, 
    101185.6, 101043.5, 100905.9, 100742.5, 100598.9, 100480.7, 100402.9, 
    100364.7,
  101841.6, 101813.5, 101733, 101624.3, 101505, 101382.9, 101278.1, 101161.4, 
    100969, 100781.9, 100642.4, 100499.9, 100337.7, 100232.8, 100162.8,
  101780.9, 101725.4, 101607.6, 101525.1, 101403.7, 101381.5, 101258.5, 
    101058.8, 100881.1, 100715.1, 100555.1, 100342.5, 100137.4, 100026.3, 
    99951.62,
  101899.8, 101851.3, 101781.4, 101687.6, 101632.9, 101571.2, 101514.2, 
    101534.5, 101579.2, 101224.6, 101264.6, 101465.5, 101265, 100780.9, 
    100569.9,
  101860.8, 101776.1, 101703.1, 101625.9, 101577.7, 101328.8, 101521.3, 
    101403.7, 101369.3, 101422.6, 101362.3, 101329.9, 101279.8, 99399.9, 
    99977.28,
  101832.4, 101760.3, 101690.8, 101648.2, 101462.3, 98097.89, 101241.1, 
    101532.8, 101412.6, 101303.2, 101205.4, 101148.1, 101074.7, 101042.2, 
    101003.9,
  101855, 101790.9, 101738.3, 101680.1, 101619.6, 101351.1, 97736.43, 
    101052.5, 101275.4, 101283.3, 101166.2, 101046.4, 100981, 100933, 100885.3,
  101921.9, 101879.8, 101839.3, 101779.9, 101739.5, 101654.6, 101396.6, 
    95443.89, 94641.66, 101042.4, 101239.8, 101104.1, 101093, 101017.6, 
    100986.1,
  101997.3, 101968.6, 101920.4, 101892.6, 101801.5, 101765.1, 101670.3, 
    101465.9, 101244.6, 101387.7, 101282.1, 101178.9, 101109.5, 101010.9, 
    100967.4,
  102064.1, 102075.8, 102053.9, 102039.5, 102000.2, 101900.1, 101799, 101734, 
    101589.5, 101387.4, 101256.6, 101136.9, 101014.6, 100905.8, 100818.3,
  102142.1, 102163.3, 102169.1, 102181.6, 102118.1, 102049.1, 101901.5, 
    101686.1, 101493.2, 101352.9, 101198.4, 101039.8, 100887.2, 100750.1, 
    100632.8,
  102225.1, 102287.9, 102331.6, 102341.5, 102279.4, 102151.6, 101973.1, 
    101779.5, 101540.3, 101299.6, 101099.7, 100926.6, 100739.2, 100580.6, 
    100426.4,
  102324.2, 102360.7, 102391.1, 102379.5, 102279.3, 102178.6, 101991.2, 
    101716.3, 101450.7, 101213.3, 101020.2, 100815.2, 100603.9, 100430.8, 
    100268.2,
  102620.5, 102538.4, 102425.5, 102286.1, 102183.8, 102117.2, 101965.1, 
    101839.3, 101676.3, 101110.6, 100955.6, 101002.2, 100663.6, 100109.2, 
    99862.08,
  102762.8, 102676.7, 102586.6, 102457.1, 102321.3, 101986.7, 102167.4, 
    101881.8, 101685.2, 101559.8, 101334.7, 101143.2, 100902.4, 98872.55, 
    99385.46,
  102845.5, 102787.2, 102714.2, 102657.3, 102323.2, 98808.26, 102001.6, 
    102224.1, 101965.9, 101714.4, 101459.7, 101283, 101047.6, 100863.1, 
    100607.1,
  102892.9, 102837.9, 102784.5, 102736.1, 102638.7, 102229.3, 98402.62, 
    101762.9, 101808.8, 101771.9, 101549.4, 101360.7, 101176.5, 101008.4, 
    100783.7,
  102900.1, 102866.4, 102816.7, 102781.7, 102704.4, 102602.3, 102237.8, 
    95988.6, 95170.7, 101570.1, 101625.1, 101391, 101240.4, 101058.5, 100969.6,
  102862.9, 102820.5, 102765.9, 102757.2, 102672.2, 102581, 102459.1, 
    102172.9, 101822.5, 101818.2, 101625.3, 101420, 101252.3, 101095.7, 
    100999.2,
  102810.8, 102773, 102719.9, 102720.5, 102680.1, 102576.8, 102426.8, 
    102297.2, 102100.4, 101826.6, 101619.4, 101433.3, 101239.2, 101085.6, 
    100971.5,
  102744.3, 102672.1, 102613.8, 102627.6, 102560.4, 102505.9, 102393.5, 
    102194.3, 101981.9, 101805.2, 101622.3, 101427.6, 101242.3, 101073.3, 
    100938.8,
  102678.2, 102599.7, 102561.4, 102544.8, 102500.6, 102436.7, 102340.7, 
    102217.7, 102031.4, 101796.3, 101612.9, 101431.6, 101236.4, 101059, 
    100912.2,
  102588.9, 102480.4, 102395, 102359.1, 102302, 102294.4, 102267.8, 102121.1, 
    101935.8, 101734.6, 101593, 101419.5, 101226.4, 101056, 100896.2,
  102935.2, 102935.3, 102907.9, 102796.9, 102699.8, 102559.8, 102375.4, 
    102315.8, 102263.7, 101760.6, 101682.1, 101770.6, 101406.4, 100742.3, 
    100393,
  102764.9, 102742.6, 102716.4, 102634.6, 102506.6, 102128, 102298.9, 
    102048.7, 101977.8, 102019.4, 101918.3, 101815.1, 101620.3, 99539.59, 
    99992.23,
  102557.8, 102543.4, 102494.8, 102451.2, 102180.9, 98715.37, 101792.3, 
    102159.5, 102009.2, 101919.4, 101856, 101799.6, 101649.7, 101513.4, 
    101270.3,
  102343.2, 102336.4, 102279.1, 102190, 102091.7, 101775, 98082.53, 101397.2, 
    101701.9, 101821.9, 101799.8, 101732.4, 101651.6, 101523.7, 101360.9,
  102163.3, 102159.8, 102090.1, 101987.8, 101880.4, 101773.3, 101538.4, 
    95615.09, 94805.85, 101356.6, 101719.9, 101647.2, 101624.2, 101484.1, 
    101402.6,
  102004.1, 101990.1, 101891.7, 101799.9, 101640.6, 101528.6, 101448.4, 
    101296.5, 101196, 101533.1, 101582.6, 101584.4, 101554.5, 101454.7, 101360,
  101865.2, 101857.2, 101757.4, 101653.9, 101489.9, 101342, 101235.5, 
    101261.7, 101409.3, 101443.5, 101486.5, 101504.4, 101461.2, 101398.5, 
    101302.3,
  101754.2, 101740.3, 101633.5, 101507, 101297.7, 101184.8, 101074.8, 
    101071.4, 101241.8, 101388.7, 101425.2, 101404.2, 101371.5, 101328.1, 
    101247.1,
  101665.9, 101656.2, 101559.9, 101390.4, 101218.8, 101097.3, 100998.6, 
    101118.5, 101304.8, 101320.5, 101330.4, 101315.9, 101278.6, 101234.7, 
    101171.7,
  101616.5, 101550.5, 101428.9, 101280.2, 101148.5, 101057.3, 101007.2, 
    101094.7, 101203.8, 101238.9, 101302.2, 101257.7, 101186.3, 101144.8, 
    101087.4,
  100951.2, 100869.8, 100791.2, 100698.4, 100648.7, 100602.4, 100526.3, 
    100482.6, 100455.7, 100106.8, 100206.1, 100573, 100576.6, 100301.2, 
    100163.8,
  100865.3, 100741.9, 100635.9, 100524.2, 100447.4, 100220.6, 100426.6, 
    100268.7, 100187.8, 100199.6, 100225.5, 100388.7, 100616.2, 98934.71, 
    99644.1,
  100804.6, 100684.6, 100572.1, 100481.2, 100288, 96994.54, 100154.3, 
    100412.3, 100255.8, 100116.8, 100080.8, 100252.5, 100548, 100783.5, 100858,
  100793.1, 100685.9, 100592.2, 100512.6, 100472.9, 100207.6, 96636.22, 
    99951.47, 100143.4, 100128.3, 100074.7, 100261.5, 100616.8, 100854.7, 
    100937.2,
  100810.8, 100745.4, 100686.3, 100627, 100633, 100534.9, 100305.1, 94403.77, 
    93685.2, 99994.33, 100276.8, 100444.7, 100717.9, 100862.6, 101008.8,
  100857.1, 100822.4, 100774.7, 100787.8, 100723, 100723, 100658.6, 100497.3, 
    100330.4, 100429, 100485.3, 100632.8, 100825.5, 100951, 101059,
  100902.7, 100924.4, 100923.8, 100940, 100939.7, 100888.4, 100852.9, 
    100843.5, 100780.5, 100668.3, 100686.9, 100793.1, 100886.1, 100983.5, 
    101065.2,
  100984.2, 101031.6, 101050.6, 101090.4, 101067.8, 101074.2, 101009, 
    100940.2, 100886.8, 100877.3, 100862.1, 100876.3, 100913.2, 100974.2, 
    101045.2,
  101095.4, 101161.4, 101245.7, 101283.5, 101296.8, 101246, 101191.8, 
    101154.6, 101068.8, 100979.1, 100930.1, 100907, 100896.6, 100912.9, 
    100953.4,
  101261.5, 101313.3, 101389.6, 101444.5, 101443.3, 101419.9, 101344.5, 
    101219.9, 101124.1, 101029.3, 100989.5, 100935.2, 100891.3, 100880.5, 
    100878.6,
  101215.4, 101110, 100972.7, 100796.9, 100688.7, 100598.3, 100400.7, 
    100207.5, 99987.09, 99384.48, 99196.94, 99278.75, 99127.03, 98864.66, 
    98924.62,
  101357.1, 101244.5, 101143.1, 100962, 100804, 100491.4, 100624.2, 100301.2, 
    100053.9, 99787.52, 99453.96, 99173.59, 99167.27, 97508.64, 98363.6,
  101460, 101369.7, 101298.8, 101182, 100831.4, 97305.16, 100510.5, 100626.3, 
    100328.7, 99955.02, 99504.94, 99157.65, 99085.88, 99272.99, 99520.46,
  101547.8, 101482.1, 101442.9, 101328.4, 101199.3, 100759.9, 96963.42, 
    100287.7, 100252.5, 100102.1, 99737.82, 99332.47, 99251.45, 99475.1, 
    99687.7,
  101635.4, 101606.1, 101582.3, 101480.9, 101367.8, 101193.3, 100816.2, 
    94604.46, 93843.66, 100133.5, 100103.4, 99773.01, 99660.98, 99698.85, 
    99872.48,
  101708.8, 101716.6, 101682.6, 101608.3, 101459.9, 101308, 101144.8, 
    100877.2, 100539, 100553.2, 100367.4, 100158.2, 100073.3, 100074.9, 
    100153.9,
  101779, 101834.8, 101799.1, 101743.4, 101617.2, 101441.6, 101228.9, 
    101087.5, 100926.7, 100741.7, 100580.4, 100473.3, 100389.8, 100366.2, 
    100378.5,
  101894, 101946.6, 101902.1, 101841.3, 101678.1, 101531.5, 101333.8, 
    101114.9, 100935.6, 100833.2, 100726.3, 100634.3, 100590.3, 100580.8, 
    100575,
  102020.5, 102066.3, 102037.4, 101941.7, 101806.9, 101635.5, 101419.6, 
    101236.8, 101069, 100925.7, 100818.6, 100751.9, 100701.5, 100677.8, 
    100665.5,
  102168.7, 102145.7, 102077.8, 101961.4, 101815.9, 101673.3, 101488.7, 
    101247.1, 101068.5, 100925.2, 100846.8, 100785.4, 100775.6, 100768.8, 
    100741.6,
  102182, 102020, 101799.1, 101556.7, 101379.1, 101225.4, 101045.7, 100875.5, 
    100693.5, 100111.1, 99906.78, 99880.07, 99539.02, 99098.16, 98969.47,
  102172.2, 101951.5, 101740.9, 101517.7, 101331.4, 100940.4, 101066.7, 
    100767.4, 100540.8, 100349.6, 100027.3, 99697.73, 99458.93, 97602.05, 
    98277.55,
  102154, 101920.5, 101695.9, 101532.2, 101192.5, 97650.47, 100770.2, 
    100924.8, 100651.5, 100362.8, 99948.88, 99571.12, 99208.12, 99189.25, 
    99272.78,
  102138.5, 101909.2, 101689.1, 101501.7, 101344.2, 100949.7, 97133.11, 
    100448.5, 100461.7, 100357.2, 100010.3, 99575.23, 99148.69, 99072.09, 
    99211.75,
  102125.7, 101923.5, 101709.7, 101525.9, 101377.3, 101227.6, 100879, 
    94687.91, 93895.2, 100210, 100151.2, 99754.3, 99367.28, 99138.85, 99279.85,
  102123.9, 101923.4, 101716.6, 101544.5, 101362.4, 101221.9, 101083.6, 
    100837.2, 100534.9, 100537.2, 100296.5, 100005.6, 99768.7, 99556.6, 
    99522.19,
  102122.7, 101952.4, 101757.3, 101609.3, 101437.8, 101282.6, 101101.2, 
    100988.4, 100872.5, 100670.3, 100451, 100231.3, 100012.5, 99881.89, 
    99806.45,
  102129.1, 101963.4, 101788.8, 101637, 101448, 101319.9, 101165.8, 100991.2, 
    100868.2, 100772.8, 100620.9, 100449.4, 100262.9, 100104.2, 99969.59,
  102148.3, 102014.3, 101873.7, 101735.6, 101585.4, 101423.1, 101250.9, 
    101122.5, 101016.8, 100900, 100765.6, 100620, 100447, 100268, 100070.5,
  102163, 102022.9, 101886.5, 101770.5, 101619.1, 101491.3, 101354, 101181.4, 
    101061.5, 100956.6, 100892.3, 100786.1, 100623.7, 100430.3, 100171.6,
  101819.2, 101827.6, 101814.2, 101693.9, 101540.7, 101419.3, 101261.1, 
    101118.6, 100966.8, 100428.1, 100273, 100298, 99892.34, 99235.83, 98921.89,
  101798.2, 101824.8, 101830, 101737.8, 101575.6, 101220.7, 101348, 101060, 
    100849.8, 100735.6, 100546, 100357.2, 100136.4, 98116.73, 98645.57,
  101770.7, 101830.8, 101841.8, 101834.9, 101524.9, 97963.41, 101151, 
    101310.5, 101089.2, 100801.5, 100547.4, 100356.3, 100145.9, 100005.2, 
    99902.7,
  101753.8, 101835.8, 101862.3, 101846.2, 101774.2, 101356, 97551.16, 100869, 
    100841.2, 100802.3, 100558.4, 100328.1, 100139.6, 99971.65, 99967.8,
  101758.5, 101880.1, 101916.5, 101918.7, 101845.7, 101732.7, 101356.7, 
    95134.77, 94345.61, 100585.3, 100587.9, 100267.6, 100099, 99909.55, 
    99905.87,
  101773.1, 101911, 101946.3, 101966.6, 101874.2, 101753.1, 101629.6, 
    101342.9, 100942.7, 100866.4, 100572.8, 100245, 100023.2, 99914.88, 
    99856.56,
  101802.2, 101958.5, 102035.4, 102063.4, 101991.2, 101854.9, 101655.5, 
    101502.6, 101264.4, 100927.4, 100577, 100203.2, 99879.43, 99760.88, 
    99781.53,
  101841.8, 102007, 102088.9, 102109.8, 102021.1, 101911.1, 101737.8, 101508, 
    101246.2, 100980.3, 100632.5, 100209.7, 99805.05, 99612.09, 99611.45,
  101875.7, 102065.4, 102174.9, 102200.5, 102150.3, 102022.2, 101821.4, 
    101644.9, 101404.8, 101097.9, 100733.3, 100298, 99824.54, 99479.03, 
    99417.27,
  101925.9, 102088.2, 102198.6, 102221.1, 102162.8, 102080.7, 101920.4, 
    101700.1, 101466.9, 101183.3, 100885.6, 100469.3, 99999.53, 99571.11, 
    99310.03,
  101037.1, 101361.9, 101656.1, 101734.9, 101750.5, 101648.9, 101457.3, 
    101259.7, 101060.4, 100495.5, 100338.3, 100381, 99984.49, 99223.11, 
    98800.73,
  101196.9, 101541, 101714.9, 101790.4, 101733.4, 101402.4, 101457.8, 
    101095.2, 100809.8, 100684, 100515.7, 100384.7, 100168.1, 98096.54, 
    98426.68,
  101438.2, 101686.8, 101809.5, 101892.2, 101641.3, 98090.86, 101171.4, 
    101304.7, 101011.2, 100686.3, 100414.9, 100307, 100172.1, 100042.1, 
    99692.51,
  101639.4, 101774.5, 101901.3, 101909.8, 101882.3, 101428.7, 97601.46, 
    100736.4, 100667.5, 100590.4, 100333.2, 100176.4, 100124.3, 100079.5, 
    99863.88,
  101782.2, 101909.8, 101989.9, 102004.7, 101936.9, 101763, 101346.5, 
    95107.65, 94270.71, 100349.4, 100289.1, 100024.4, 100056.8, 100040.8, 
    100014,
  101900.2, 102004.2, 102059.1, 102072, 101964.4, 101801.8, 101607.4, 
    101245.7, 100786.1, 100622.8, 100257.4, 99969.67, 99975.34, 100050.7, 
    100057,
  101980.7, 102095.1, 102164.3, 102174.5, 102078.7, 101894.7, 101654.4, 
    101435.2, 101140, 100725.5, 100321.3, 100021.7, 99921.98, 100032.4, 
    100084.4,
  102033.5, 102164.8, 102234.9, 102228.4, 102115.9, 101978.9, 101759.8, 
    101466.7, 101156.4, 100840.7, 100482.6, 100151.8, 99991.32, 100066, 100115,
  102080.4, 102241.3, 102318.3, 102319.4, 102231.4, 102089.3, 101877.4, 
    101645.9, 101376.1, 101031.8, 100673.2, 100338.8, 100097, 100083.4, 100152,
  102126.9, 102273.6, 102337, 102316.3, 102236, 102155.5, 101992.1, 101739.5, 
    101478.1, 101175.8, 100874.2, 100549.5, 100249.7, 100109.1, 100163.7,
  101449.8, 101577.4, 101634, 101612.6, 101538.2, 101435.3, 101295.3, 
    101170.4, 101017.4, 100494.3, 100370.8, 100488.5, 100234.9, 99695.25, 
    99376.9,
  101707.7, 101759.3, 101738.2, 101682, 101540.2, 101206, 101307.1, 101051.7, 
    100827, 100669.9, 100489.2, 100367.7, 100257.1, 98301.84, 98740.15,
  101862.6, 101870.8, 101847.6, 101804.9, 101473.5, 97932.66, 101080.8, 
    101227.4, 100975.7, 100677.6, 100425.8, 100305.8, 100201, 100117.3, 
    99822.2,
  101975.3, 101965.6, 101930.3, 101864.5, 101765.5, 101332.5, 97519.21, 
    100795.1, 100766.9, 100676.9, 100438.2, 100292, 100195.8, 100079.2, 
    99741.62,
  102050.2, 102066.2, 102029.9, 101964.2, 101855.1, 101713.2, 101318.8, 
    95132.78, 94352.87, 100503.5, 100505.1, 100297.1, 100223.3, 100033.6, 
    99784.95,
  102100.1, 102127.3, 102101.7, 102052.6, 101919.6, 101780.9, 101607.4, 
    101302.3, 100907, 100794, 100553.9, 100355.7, 100257.8, 100087.8, 99837.57,
  102104.1, 102159, 102170.5, 102140.1, 102027.2, 101878.2, 101670.9, 101489, 
    101257.1, 100928.5, 100646.1, 100430.2, 100302.1, 100161.6, 99944.63,
  102068, 102147.7, 102192.2, 102182, 102064.7, 101962.5, 101777, 101527, 
    101282, 101043.8, 100789.2, 100534.9, 100371.7, 100249.7, 100073.3,
  102000.1, 102109.1, 102206, 102216.5, 102119.9, 102043.6, 101873.9, 
    101682.8, 101472.7, 101213.7, 100952.2, 100676.9, 100472.2, 100349.5, 
    100207.2,
  101914.4, 102018.4, 102138.9, 102169.1, 102105.1, 102086.6, 101966.5, 
    101755.3, 101546.8, 101321.7, 101113.2, 100860.4, 100607.1, 100457.3, 
    100367.1,
  102058.3, 102060.5, 101978.2, 101853.1, 101727, 101631, 101510, 101412.1, 
    101271.8, 100785.1, 100660.3, 100774, 100524.3, 100070.5, 99891.38,
  102089.4, 102065.2, 102018.6, 101912.3, 101765.1, 101450.3, 101562.6, 
    101338.4, 101162.4, 101052.8, 100857.5, 100725.1, 100611.7, 98678.81, 
    99259.67,
  102074.6, 102078.2, 102042.7, 102020.6, 101705.8, 98164.38, 101372.7, 
    101512.2, 101294.2, 101072.8, 100824.9, 100661, 100506.6, 100427.2, 
    100301.6,
  102060.4, 102087.1, 102063, 102041.4, 101958.2, 101582, 97740.53, 101125.6, 
    101144, 101070.9, 100814.9, 100599.5, 100429.6, 100303, 100139.9,
  102025.8, 102104.8, 102100.8, 102089.5, 102006.7, 101895.2, 101541.7, 
    95377.13, 94593.67, 100865.2, 100841.8, 100551.1, 100369.8, 100178.9, 
    100033.5,
  101976.1, 102083.8, 102104.6, 102119.2, 102026.5, 101921.1, 101762.1, 
    101508.6, 101174.6, 101116.2, 100852.7, 100552.9, 100337.1, 100112.2, 
    99922.29,
  101915.2, 102062.4, 102116.4, 102157.9, 102085.5, 101978.1, 101786.4, 
    101642.3, 101443.6, 101178.2, 100889.9, 100588.5, 100321.8, 100089.3, 
    99884.12,
  101878.9, 102036.1, 102082.6, 102163.8, 102095.5, 102024.7, 101842.9, 
    101644.4, 101440.1, 101248.2, 100976.5, 100654.7, 100357.5, 100107.2, 
    99894.34,
  101838.8, 101960, 102081.6, 102187.7, 102153.5, 102090.5, 101933.9, 
    101760.8, 101565.6, 101342.8, 101079.8, 100754.4, 100423.4, 100161.6, 
    99947.23,
  101819, 101923.9, 102029.7, 102139.4, 102151, 102132, 102011.7, 101816.9, 
    101634.2, 101421.5, 101213.5, 100891.1, 100530.4, 100262.9, 100060.7,
  102310.7, 102367.8, 102339.7, 102253, 102170.1, 102064.2, 101937.8, 
    101834.8, 101704.5, 101207.4, 101091.6, 101125.1, 100758.5, 100173.1, 
    99917.84,
  102345.1, 102345.2, 102351.2, 102278.7, 102171.8, 101849.2, 101971.4, 
    101740, 101585.9, 101502.1, 101327.7, 101132.4, 100890.7, 98859.03, 
    99370.86,
  102329, 102360.8, 102352.4, 102342.5, 102075.4, 98514.95, 101750.4, 
    101912.6, 101725.2, 101543.7, 101325.5, 101119.5, 100873.8, 100685.7, 
    100492.1,
  102296.4, 102351.1, 102371.5, 102348.9, 102277.5, 101913.1, 98084.62, 
    101497.4, 101556, 101541.5, 101324.8, 101087.9, 100828.1, 100627.6, 
    100457.6,
  102308.2, 102393.3, 102404, 102393.1, 102315.5, 102199.9, 101869.3, 
    95722.78, 94927.41, 101303.4, 101332.6, 101039.8, 100769, 100534.6, 
    100390.8,
  102341.1, 102413.5, 102410.6, 102424, 102321.3, 102210.7, 102081.8, 101852, 
    101540.1, 101538.1, 101300.2, 100997.3, 100685.9, 100456.9, 100292.6,
  102380.9, 102440.2, 102442.8, 102464.1, 102382.5, 102250.2, 102086, 
    101967.6, 101786.7, 101540.6, 101274.1, 100951.2, 100611.6, 100397.2, 
    100225.5,
  102429.4, 102441.9, 102433.4, 102461.7, 102366.5, 102267.1, 102105.3, 
    101919, 101732.1, 101532.9, 101269.6, 100915, 100578.3, 100377.6, 100227.9,
  102457.7, 102457.9, 102434.1, 102452.2, 102377.8, 102267.8, 102128.1, 
    101985.6, 101805.1, 101560.8, 101283.6, 100908.1, 100573.9, 100395.3, 
    100262.1,
  102500.8, 102431.1, 102375, 102333.1, 102254, 102189.9, 102116.3, 101958.1, 
    101799.5, 101569.9, 101322.5, 100933.3, 100608.6, 100440.2, 100325.5,
  102430.6, 102406.4, 102362.3, 102267.4, 102192.2, 102095.2, 101987.1, 
    101928.2, 101856.3, 101412.1, 101382.5, 101535.2, 101239.6, 100634.2, 
    100328.2,
  102443.3, 102367, 102310.2, 102220.3, 102111, 101813.5, 101966, 101775.9, 
    101678.8, 101675.4, 101576, 101509, 101344.5, 99300.91, 99793.88,
  102393.6, 102315.5, 102213.2, 102158.8, 101901.1, 98394.14, 101612.1, 
    101874.6, 101712.4, 101610.1, 101498.8, 101429.5, 101272.4, 101117.4, 
    100926.8,
  102327.1, 102240.9, 102114, 102016.3, 101913.3, 101608.5, 97862.5, 
    101262.7, 101461, 101508.1, 101419.8, 101314.6, 101178.1, 101029.9, 100871,
  102284.9, 102145.1, 101995.2, 101871, 101758.5, 101657.2, 101411, 95426.94, 
    94625.76, 101102.8, 101318.6, 101178, 101057, 100891.4, 100790.9,
  102187.3, 102001.9, 101834, 101700.1, 101556, 101458, 101369.8, 101221.7, 
    101052.1, 101231.6, 101150.3, 101044.4, 100906.4, 100756.8, 100669.3,
  102086.4, 101904.3, 101735.3, 101596.5, 101460.3, 101309.8, 101168.1, 
    101125.2, 101094.4, 101040.2, 100980.9, 100892.4, 100736.9, 100612.8, 
    100532.3,
  102022.5, 101841.6, 101665.2, 101501.2, 101318.4, 101155.3, 101003.9, 
    100876.5, 100855.7, 100889, 100848.1, 100735.1, 100588.8, 100476.7, 
    100397.2,
  102000.5, 101836, 101663.4, 101477.2, 101288.3, 101085.3, 100914.6, 100866, 
    100867.5, 100820.3, 100724.1, 100582.1, 100427.1, 100330.4, 100265.3,
  102021.1, 101826.2, 101635.8, 101467, 101265.3, 101072.1, 100938.9, 
    100843.7, 100818.2, 100727.6, 100617, 100429.8, 100260.5, 100177.8, 100120,
  101732.1, 101736.1, 101740, 101720.7, 101721.3, 101682.3, 101639.4, 
    101655.5, 101685.4, 101360.2, 101447.2, 101738, 101591.9, 101132.3, 
    100892.1,
  101659.6, 101605, 101562, 101516, 101463.7, 101249.9, 101417.2, 101360, 
    101380.2, 101488.5, 101530.9, 101639.9, 101694.9, 99806.32, 100416.8,
  101589.7, 101489.9, 101401.7, 101344.8, 101128.8, 97689.5, 100888.3, 
    101163.1, 101087.3, 101168.8, 101297.7, 101454.4, 101600.8, 101675.3, 
    101648.6,
  101507.4, 101398.1, 101300.4, 101205, 101110.3, 100793.1, 97144.42, 100499, 
    100835.6, 100905, 101063.1, 101241, 101469.4, 101613.2, 101677,
  101486.5, 101376.6, 101287.1, 101182.2, 101073.6, 100956.5, 100675.2, 
    94773.78, 93972.67, 100402.7, 100813.7, 101013.9, 101317.7, 101498.8, 
    101657.1,
  101511.8, 101400.1, 101294.8, 101183.8, 100987.1, 100848.9, 100742.4, 
    100559.6, 100409, 100653, 100651.5, 100859.4, 101172.2, 101417.8, 101589.6,
  101558.4, 101455.9, 101327.6, 101174.4, 100945.3, 100714.2, 100538.3, 
    100495.4, 100421.8, 100407.4, 100533.5, 100748, 101058.3, 101337.6, 
    101519.1,
  101601.3, 101471.1, 101314.5, 101121.1, 100829.9, 100587.4, 100378, 
    100247.2, 100225, 100306.7, 100443.6, 100664.6, 100987.8, 101271.5, 
    101465.4,
  101648.5, 101523.2, 101361.7, 101144.9, 100855.1, 100530.9, 100283, 
    100215.5, 100248, 100242.9, 100368.6, 100622.1, 100936.3, 101218.1, 
    101413.3,
  101725.1, 101553.5, 101369.5, 101136.9, 100823.8, 100494.2, 100225.2, 
    100030.7, 100097.4, 100192.9, 100349.5, 100604.1, 100904.4, 101186.1, 
    101383.1,
  101504.5, 101462.9, 101418.2, 101372.8, 101345.6, 101311.7, 101300.7, 
    101349.3, 101438, 101190.8, 101350.7, 101705.7, 101655.8, 101311, 101152.6,
  101489.7, 101399.7, 101341.2, 101279.6, 101236.7, 101039.1, 101244.4, 
    101182.9, 101234.1, 101388.9, 101501.7, 101640.7, 101768.4, 99974.41, 
    100653.1,
  101368.3, 101264.2, 101178.8, 101125, 100989, 97599.8, 100926.5, 101221.5, 
    101152.2, 101213.1, 101364.6, 101529.8, 101704.3, 101834.8, 101882.9,
  101245.8, 101119.6, 101000.7, 100924.6, 100901.4, 100724.4, 97158.04, 
    100734.4, 101081.5, 101099.5, 101212.4, 101394.3, 101619, 101824.7, 
    101939.1,
  101131.3, 100991.9, 100880.4, 100803.8, 100825, 100794.4, 100656.9, 
    94878.2, 94216.48, 100814.6, 101105.3, 101267.9, 101534.9, 101765, 
    101975.8,
  101050.4, 100905.3, 100789.8, 100784.8, 100714.5, 100666.3, 100651.5, 
    100624.3, 100600.1, 100984.9, 101017, 101185, 101472.7, 101773.6, 101973.7,
  101001.6, 100865.1, 100775.8, 100734.7, 100635.9, 100529.1, 100442.2, 
    100510.9, 100671, 100867, 101001, 101140.3, 101455.8, 101792.1, 101986.8,
  100983.2, 100844.2, 100742.5, 100648.1, 100487.1, 100371.1, 100292.8, 
    100301.8, 100482.7, 100822.1, 100984.4, 101138, 101496.9, 101841.7, 
    102037.7,
  101004.2, 100861.3, 100733.9, 100580.8, 100388.9, 100245.8, 100200.7, 
    100276.2, 100501, 100811.5, 100980.1, 101195.4, 101581.8, 101907.3, 
    102098.4,
  101050.6, 100874.7, 100706.5, 100530.2, 100326.5, 100204.2, 100187.2, 
    100257, 100547.3, 100800.4, 101006.7, 101319.9, 101703.6, 102002.7, 
    102165.6,
  100781.7, 100775.6, 100802, 100830.6, 100931.7, 100993, 101036.4, 101091.8, 
    101108.1, 100830.2, 100994.1, 101364.3, 101307.7, 100982.2, 100846.2,
  100690.5, 100652.6, 100652.6, 100655.9, 100704, 100637.6, 100929.4, 
    100982.7, 101034.9, 101136.5, 101234.5, 101406, 101522.2, 99737.03, 
    100425.1,
  100644.4, 100571.5, 100541.6, 100513.1, 100420.1, 97134.23, 100505.8, 
    100934.2, 101028.7, 101114.6, 101237.7, 101413.3, 101580.9, 101671.5, 
    101704.7,
  100572.8, 100484.8, 100441.6, 100403.1, 100417.3, 100246.4, 96762.59, 
    100424.8, 100927.7, 101077.6, 101242.6, 101396.6, 101597.6, 101745.2, 
    101825,
  100508.3, 100431.9, 100400.3, 100402.4, 100453.8, 100502.7, 100265.8, 
    94674.02, 94186.16, 100795.9, 101245.1, 101397.1, 101618, 101737.9, 
    101909.9,
  100477.2, 100382.2, 100329.6, 100384.9, 100416.1, 100471.8, 100507.7, 
    100438.5, 100494.9, 100991.4, 101190.8, 101411.5, 101626.2, 101793, 
    101935.2,
  100453.2, 100373, 100344.2, 100335.2, 100383.8, 100450.2, 100454.2, 
    100589.9, 100822.5, 100977.7, 101202.6, 101441.8, 101646.7, 101822.4, 
    101914.6,
  100486.9, 100409.7, 100352.4, 100298.5, 100282.3, 100412.5, 100463.2, 
    100543.7, 100757.8, 101025.1, 101263.9, 101487.5, 101700, 101865.5, 
    101921.9,
  100546.5, 100461.6, 100384.4, 100306, 100302.9, 100404.6, 100512.2, 
    100708.1, 100922.6, 101124.6, 101337.9, 101562.2, 101761.6, 101891.3, 
    101948.5,
  100650.6, 100546.3, 100454.8, 100374.9, 100367.3, 100467.2, 100599.6, 
    100763.4, 100976.8, 101183, 101433.4, 101657.5, 101837.3, 101949.6, 
    101960.3,
  100763.4, 100793.4, 100788.5, 100754.8, 100705.2, 100689, 100732.8, 
    100848.2, 100924.5, 100630.2, 100751.7, 100932.6, 100621.4, 100039.2, 
    99699.1,
  100767.9, 100723.2, 100703.1, 100646.4, 100593, 100427.6, 100686.4, 
    100778.2, 100855.2, 100927.6, 101010.4, 101009.2, 100877.3, 98894.06, 
    99397.94,
  100692.2, 100627.4, 100584.4, 100549.4, 100407, 97056.89, 100441.7, 
    100793.9, 100880.1, 100940.6, 101042.5, 101083.5, 101025.5, 100927.9, 
    100745.4,
  100618, 100546.1, 100485.3, 100461.5, 100434.9, 100225.8, 96722.55, 
    100411.1, 100792.2, 100931.8, 101079.1, 101138.2, 101140.2, 101096.5, 
    101020,
  100539.2, 100465.2, 100399.7, 100379.7, 100432.3, 100443.7, 100261.2, 
    94648.28, 94134.31, 100718.6, 101124.1, 101211.7, 101265.9, 101224.8, 
    101249.5,
  100506.7, 100396.2, 100361.6, 100335.7, 100400.1, 100487.8, 100522.6, 
    100455.4, 100472.1, 100939.4, 101141.7, 101294.1, 101372.7, 101399.9, 
    101416.2,
  100447.8, 100364.5, 100366.7, 100364.1, 100413.5, 100526.8, 100566.2, 
    100606.7, 100788, 100978.7, 101202, 101392, 101495.6, 101559.6, 101592.2,
  100459, 100383.1, 100372.4, 100352.5, 100384.4, 100528.4, 100563.1, 
    100578.6, 100766.1, 101055.6, 101289, 101492.5, 101624.7, 101704.7, 
    101762.5,
  100511.1, 100446.7, 100401.1, 100390.6, 100461.6, 100547.9, 100577.9, 
    100718.5, 100935.5, 101186.5, 101401.1, 101610.8, 101737.9, 101827.7, 
    101887.2,
  100637.6, 100571.5, 100533.7, 100508.5, 100529.2, 100587.1, 100659.4, 
    100811.3, 101050.8, 101272.3, 101514.5, 101708.8, 101841.4, 101942.5, 
    102002.6,
  101198.6, 101249.6, 101248.2, 101253.6, 101262.4, 101256.8, 101231.1, 
    101221.1, 101223.4, 100880.9, 100961.1, 101204.4, 100978, 100407.3, 
    100010.6,
  101194.5, 101174.9, 101186.9, 101155.7, 101140, 100950.7, 101128.9, 
    101075.6, 101076.1, 101106.3, 101137.6, 101157, 101058.4, 99036, 99438.2,
  101145.1, 101111.3, 101077.3, 101047.8, 100911.1, 97537.73, 100812.8, 
    101025.9, 101042.9, 101071.4, 101119.2, 101098.5, 100975.2, 100791.4, 
    100571.8,
  101077.6, 101021.5, 100953.1, 100920.8, 100892.9, 100713.4, 97105.95, 
    100685.7, 101022.3, 101050.8, 101093.9, 100996.1, 100881.3, 100718, 
    100655.1,
  101001.5, 100922.6, 100865.1, 100820.4, 100833.6, 100866.1, 100712.3, 
    94916.98, 94282.88, 100787.2, 101045.7, 100913.8, 100818.6, 100703.7, 
    100808.5,
  100941.5, 100857, 100819.2, 100829.1, 100827.1, 100828.6, 100823.6, 
    100806.8, 100720.3, 101008.6, 100970.6, 100879.5, 100827.9, 100844.2, 
    100952.9,
  100896.2, 100844.1, 100846.8, 100867.3, 100862.6, 100882.1, 100811.8, 
    100917.3, 101020.4, 101035.5, 100980.9, 100946.2, 100963.9, 101043.1, 
    101162.4,
  100901.7, 100871.3, 100881.8, 100869.4, 100878.1, 100895.9, 100885.7, 
    100969.3, 101081.2, 101127.6, 101124.6, 101144.2, 101218.7, 101325.4, 
    101438.6,
  100933.8, 100914.1, 100933.8, 100953.4, 100965.6, 100983.8, 101026.5, 
    101171.4, 101282.6, 101314.9, 101340.2, 101399.2, 101479.3, 101573, 
    101653.3,
  101020.6, 100990.1, 101005.4, 101021.2, 101045.7, 101099.8, 101200, 
    101320.5, 101428.6, 101472, 101568, 101649.5, 101722.8, 101807.3, 101868,
  101202.2, 101280.7, 101390.4, 101451.9, 101508.7, 101537, 101550.7, 
    101596.7, 101656.5, 101345.6, 101420.6, 101690.1, 101562.1, 101197.7, 
    101061.3,
  101319, 101382.7, 101432.8, 101426.4, 101433, 101251.3, 101463.9, 101426.8, 
    101447, 101516.7, 101529, 101589.1, 101632.2, 99823.18, 100465.1,
  101401.7, 101404.3, 101406, 101399.4, 101265.9, 97878.16, 101110.5, 
    101357.1, 101283.8, 101333, 101372, 101458.5, 101532.2, 101586.7, 101569.4,
  101413.4, 101410.8, 101355.8, 101313.4, 101270.9, 101064.6, 97451.43, 
    100900.8, 101206.1, 101243.8, 101300.1, 101349.2, 101437.7, 101501.2, 
    101498,
  101380.5, 101336.2, 101280.8, 101254, 101281.4, 101253.2, 101035.6, 
    95153.67, 94422.91, 100908, 101206.7, 101244.2, 101325.9, 101341.3, 
    101396.9,
  101328.8, 101289.6, 101253.9, 101279.2, 101195.6, 101145.3, 101108, 
    101014.9, 100875.3, 101066.6, 101074.8, 101138.8, 101191.3, 101239.9, 
    101299.2,
  101302.5, 101270.8, 101283.3, 101230.5, 101142.2, 101052.4, 100956.4, 
    100986.8, 100981, 100971.7, 100992.6, 101033.5, 101073.8, 101164, 101269.5,
  101309.5, 101307.7, 101272.4, 101168.7, 101033.4, 100961.3, 100931.4, 
    100880.2, 100849.7, 100837.2, 100888.5, 100962.4, 101078.5, 101228.8, 
    101381.8,
  101354, 101359.8, 101289.2, 101167.3, 101062.4, 100989.2, 100898.4, 
    100834.3, 100743.6, 100793.4, 100902.3, 101053.3, 101214.5, 101380.8, 
    101499.6,
  101439, 101408, 101339.7, 101222.7, 101086.2, 100979.9, 100886.5, 100816, 
    100825.3, 100901.1, 101083.4, 101257.1, 101414.6, 101555.2, 101652.9,
  101184.3, 101406.8, 101600.7, 101760, 101899.8, 101940.7, 101902.8, 
    101911.1, 101903.3, 101504.7, 101523.5, 101738.1, 101548, 101162.1, 
    101011.5,
  101096.3, 101302.6, 101534.2, 101713.6, 101815.9, 101659.5, 101880.5, 
    101756.1, 101719.2, 101739.5, 101673.1, 101694.6, 101698.8, 99859.62, 
    100527.5,
  101013.5, 101262, 101478.8, 101639.3, 101617.3, 98277.12, 101511.2, 
    101811.1, 101661.4, 101626.8, 101577.8, 101596.4, 101635.2, 101704, 101697,
  100951, 101253.6, 101426.5, 101573.8, 101596.3, 101462.3, 97866.43, 
    101304.6, 101570.1, 101551.8, 101514.3, 101503.8, 101558, 101661.4, 
    101719.9,
  101025.5, 101259.4, 101398.9, 101488.6, 101606.2, 101597.3, 101429, 
    95546.48, 94774.73, 101248.1, 101467.2, 101449.2, 101503.7, 101587.4, 
    101721,
  101100, 101290.7, 101368.6, 101479.7, 101454.3, 101474.9, 101446, 101359, 
    101248.9, 101451.7, 101402.5, 101432.9, 101470.4, 101570.7, 101685.7,
  101198.4, 101326, 101375.4, 101414.6, 101377.4, 101319.5, 101277.6, 
    101340.2, 101355.4, 101374.6, 101414.3, 101439.4, 101480.7, 101565.8, 
    101655.8,
  101297.3, 101343.9, 101352.1, 101309.1, 101177.4, 101138.6, 101148.5, 
    101176.6, 101241.1, 101354.1, 101412.1, 101448, 101495.1, 101557.4, 
    101625.4,
  101351.4, 101341.1, 101290.8, 101169.9, 101045.7, 101010.1, 101070.7, 
    101181, 101253.2, 101309.7, 101369.7, 101424.5, 101453.4, 101510.5, 
    101561.3,
  101363.7, 101292.5, 101211.1, 101048.6, 100906.8, 100926.9, 101007.1, 
    101089.8, 101168.8, 101221.2, 101300.1, 101375.3, 101420.1, 101489.3, 
    101540.3,
  100125.6, 100123.8, 100167.3, 100205.2, 100291.1, 100381.9, 100514, 
    100695.5, 100904.6, 100767.9, 101038, 101474.3, 101476.7, 101221.6, 
    101166.9,
  99892.7, 99850.91, 99880.05, 99929.31, 100015.1, 100034.3, 100385, 
    100539.4, 100737.8, 100995.6, 101217.1, 101458, 101625.2, 99907.09, 
    100647.9,
  99632.46, 99581.59, 99620.45, 99720.76, 99764.83, 96758.48, 100182.6, 
    100634.1, 100786.9, 101035.3, 101271.2, 101505.3, 101644.8, 101754.8, 
    101820.8,
  99414.69, 99351.25, 99431.15, 99604.07, 99840.08, 99873.26, 96796.83, 
    100479.3, 101001.7, 101199.5, 101400.4, 101540.4, 101690.1, 101792.2, 
    101855.1,
  99318.1, 99319.45, 99497.76, 99770.98, 100098.9, 100380.6, 100388.9, 
    94906.98, 94435.12, 101086.1, 101496.4, 101585.1, 101706.8, 101761.3, 
    101897.6,
  99682.98, 99730.4, 99909.59, 100158.5, 100368, 100640.8, 100861.4, 
    100902.2, 101022.4, 101430, 101529.4, 101615.9, 101703.4, 101788.8, 
    101893.7,
  100167.5, 100234.4, 100364.9, 100528.1, 100729, 100882.6, 101068.5, 
    101298.2, 101434.8, 101494, 101589.1, 101619.5, 101678.7, 101794.1, 101905,
  100527.5, 100606.8, 100718, 100833.1, 100958.2, 101109.2, 101238, 101332.6, 
    101471.9, 101603.7, 101643.3, 101661.7, 101741.5, 101847.7, 101951.4,
  100805.1, 100885.1, 100965.8, 101051.6, 101161.2, 101277.1, 101416.2, 
    101559.3, 101636.8, 101671.4, 101714.6, 101766.8, 101827.2, 101913.4, 
    101991.6,
  100977.1, 101034, 101112, 101191.5, 101300.7, 101419.6, 101516.2, 101580.3, 
    101640.1, 101673.6, 101758.3, 101829.8, 101888.5, 101958.8, 101989.5,
  101608.9, 101409, 101157.7, 100861.7, 100621.3, 100452.1, 100351.5, 100292, 
    100263.8, 99925.76, 99951.53, 100185.7, 100039.3, 99710.74, 99673.91,
  101507, 101187, 100860.7, 100516.6, 100249.4, 99918.66, 100054.6, 99979.9, 
    99924.66, 99917.49, 99888.18, 99908.11, 99949.71, 98287.91, 99069.94,
  101333.6, 100978.3, 100604.6, 100251.3, 99909.52, 96566.76, 99792.02, 
    100011.2, 99903.75, 99852.97, 99783.58, 99774.59, 99841.29, 99978.74, 
    100208.9,
  101242.6, 100880.6, 100490, 100196.8, 100018.2, 99781.43, 96434.88, 
    99904.04, 100087.3, 100042.5, 99937.59, 99883.79, 99933, 100135.4, 
    100387.3,
  101244.2, 100956.8, 100650.3, 100462.6, 100337.6, 100321.8, 100135.1, 
    94366.67, 93812.78, 100117.9, 100257.6, 100168.1, 100236.5, 100372.2, 
    100651.6,
  101362.6, 101185.4, 100984.1, 100833.7, 100729.3, 100728.2, 100728.2, 
    100613.8, 100490.6, 100642.7, 100609.1, 100585.5, 100644.8, 100758.5, 
    100944.6,
  101472.9, 101401.2, 101295.7, 101210.5, 101133.8, 101080.5, 101050.8, 
    101069.1, 101029.6, 100941.3, 100920.3, 100937.8, 100982.5, 101076.2, 
    101201.9,
  101608, 101597.2, 101545.1, 101485.1, 101411.2, 101374.2, 101315.1, 
    101243.8, 101206.4, 101203.7, 101194.1, 101214.6, 101262.5, 101337.2, 
    101416.7,
  101685.2, 101740.2, 101736.5, 101712.2, 101674.1, 101620.9, 101557.9, 
    101522.4, 101459.4, 101405.4, 101392.3, 101420.1, 101457.7, 101497.2, 
    101518.7,
  101771.8, 101834.1, 101852.1, 101832.5, 101796, 101765.4, 101717.6, 
    101634.5, 101583.1, 101544.7, 101586.7, 101612.1, 101631.9, 101644.2, 
    101620.7,
  101479.8, 101626.3, 101796.5, 101895.2, 101918.6, 101887.6, 101867.8, 
    101805.6, 101686.5, 101155.3, 101008.6, 101043, 100692.2, 100127.9, 
    99897.57,
  101331.3, 101479.9, 101686, 101816.4, 101865.8, 101700.4, 101910, 101727, 
    101593.1, 101456.2, 101206.8, 100947.5, 100691.4, 98694.35, 99200.38,
  101180.9, 101387.2, 101622.6, 101808.1, 101745.4, 98393.71, 101699.5, 
    101899.5, 101705.7, 101470.8, 101183.8, 100867.4, 100540.5, 100313.8, 
    100190.7,
  101038.5, 101342.3, 101613.2, 101820.4, 101915, 101701.8, 98063.83, 
    101483.9, 101596.6, 101500.4, 101195.4, 100802.8, 100424.9, 100119.5, 
    100059,
  101247.7, 101524, 101745.2, 101908.6, 101998.3, 102000.4, 101786.1, 
    95792.65, 94994.87, 101269.3, 101258.1, 100804.8, 100384.2, 99974.18, 
    100001.3,
  101576.2, 101735, 101875, 102001.8, 102014.5, 102022.4, 101981.9, 101805.9, 
    101566.6, 101567.9, 101290.7, 100885.3, 100458.5, 100072.1, 100057.8,
  101742.6, 101895.9, 102001.9, 102076.1, 102084.6, 102044.2, 101961.6, 
    101919.1, 101778.1, 101580, 101328.6, 100978.9, 100610.6, 100352.4, 
    100319.1,
  101876.5, 101972.3, 102053.3, 102095.9, 102064.4, 102029.6, 101941.4, 
    101817.1, 101721.7, 101603, 101385.1, 101074.3, 100817.4, 100681.3, 
    100639.2,
  101897.4, 102017.3, 102100.7, 102088.5, 102047.9, 101977.2, 101891.9, 
    101839.7, 101744.8, 101606.6, 101419.7, 101171.1, 100981.9, 100893, 
    100878.8,
  101957, 102052, 102052.6, 102015.8, 101940.2, 101877.8, 101810.6, 101735.3, 
    101664.8, 101559.6, 101440.4, 101259.6, 101131.6, 101089.2, 101095.6,
  101595.9, 101229.4, 100836, 100468.8, 100234.6, 100148, 100273.8, 100514, 
    100819.5, 100766.8, 101095.4, 101550.9, 101506.4, 101100.2, 100880.7,
  101496.4, 101055, 100627.7, 100278.2, 100031.6, 99876.52, 100190.9, 
    100437.2, 100752.3, 101099.9, 101361, 101580.8, 101632.7, 99757, 100253.7,
  101430.7, 100976, 100565, 100250.2, 99947.68, 96693.96, 100142, 100611.4, 
    100926.9, 101217.9, 101438.2, 101584.4, 101581.5, 101473.7, 101259.3,
  101489.7, 101082.6, 100747.5, 100468, 100371.3, 100110.9, 96941.76, 
    100684.2, 101174.5, 101386.1, 101542.2, 101549.3, 101477.5, 101276.4, 
    100993.1,
  101668.5, 101411.3, 101163.9, 100977.2, 100871.4, 100928.9, 100726.2, 
    95102.84, 94663.11, 101255.5, 101589.2, 101475.6, 101333.2, 101005, 
    100704.9,
  101797.5, 101672.2, 101514.7, 101389.9, 101251, 101232.3, 101344.3, 
    101257.5, 101239.3, 101573.9, 101550.2, 101408.2, 101174.9, 100816.6, 
    100630.5,
  101853.6, 101815.4, 101730.2, 101647.6, 101580.2, 101530.3, 101493.1, 
    101606.7, 101660.1, 101582.9, 101503.7, 101312.1, 101057.5, 100809.6, 
    100705,
  101860.6, 101860.1, 101827.3, 101766.5, 101682.6, 101672, 101655.5, 
    101594.4, 101585.7, 101572.5, 101449, 101217.7, 101063.6, 100940, 100855.6,
  101829.1, 101835.2, 101828.5, 101776, 101720.9, 101684.4, 101657.6, 
    101683.3, 101655.1, 101558.4, 101369.4, 101199.8, 101109, 101038.7, 
    101011.8,
  101808.8, 101762.9, 101727.9, 101698.3, 101659, 101667.5, 101646.3, 101597, 
    101556.4, 101481.7, 101347.3, 101259, 101218.9, 101195.9, 101186.2,
  102627.4, 102579.5, 102527.9, 102443.2, 102200.8, 101823, 101424.7, 
    100956.9, 100504.6, 99839.8, 99736.05, 99954.95, 99916.12, 99683.07, 
    99675.6,
  102501.1, 102464.6, 102486.2, 102422.8, 102188.7, 101618.4, 101576.9, 
    101077.2, 100654.8, 100380.2, 100257.4, 100321.7, 100368.7, 98694.68, 
    99442.49,
  102386.1, 102402.9, 102453.1, 102444.8, 102099.3, 98456.71, 101469.3, 
    101480.4, 101113.4, 100834.8, 100700.4, 100718.5, 100759.9, 100799.4, 
    100808.2,
  102269, 102324.1, 102434.3, 102418.8, 102302.6, 101834.6, 98030.23, 
    101314.6, 101292.8, 101206.6, 101075.4, 101023, 101016.4, 101038, 101004,
  102173.8, 102292.6, 102397.1, 102421.6, 102345.9, 102173.6, 101817.5, 
    95681.36, 94983.41, 101233.6, 101313.1, 101177.1, 101122, 101029.2, 
    100985.5,
  102148.5, 102247.5, 102324.5, 102389.4, 102317, 102228.8, 102125, 101924.2, 
    101576.8, 101587.3, 101417.8, 101286, 101175.2, 101085.8, 101048.2,
  102132, 102163.2, 102193.4, 102266.2, 102272.8, 102237.2, 102125.3, 
    102061.2, 101933.5, 101694.4, 101498.9, 101364.8, 101252, 101178.4, 
    101144.4,
  102074.1, 102044.3, 102024.1, 102090.4, 102120, 102163.4, 102151.8, 102056, 
    101900.1, 101744.5, 101577.9, 101441.9, 101348.1, 101290.5, 101269.4,
  102019.1, 101970.7, 101930.8, 101932.2, 101987.4, 102074.6, 102095.9, 
    102078.2, 101997.1, 101804.2, 101644.7, 101543.3, 101459.5, 101417.5, 
    101382.5,
  102000.9, 101918.1, 101851.3, 101808.1, 101847.3, 101964.8, 102071.7, 
    102026.6, 101923.8, 101768.2, 101709.5, 101652, 101577.4, 101540, 101506.5,
  102259.2, 102336.5, 102383.7, 102464.1, 102673.7, 102753.6, 102679.4, 
    102553.1, 102356.1, 101711, 101475.5, 101457.1, 101041.6, 100365.4, 
    100006.1,
  102263.3, 102297.5, 102368.7, 102517.5, 102697.7, 102529.6, 102742.1, 
    102494.5, 102292.2, 102057.5, 101768.9, 101560.9, 101289.7, 99244.57, 
    99657.34,
  102287.6, 102378.9, 102463.1, 102616.2, 102578.2, 99186.85, 102481.2, 
    102651.2, 102392.5, 102137.2, 101834.8, 101627.7, 101400.4, 101205.2, 
    100921.8,
  102374.1, 102405.3, 102513.2, 102676.6, 102734.7, 102544.6, 98837.55, 
    102255.2, 102319.2, 102173.1, 101911.3, 101677.6, 101475.2, 101297.8, 
    101085.7,
  102422.8, 102479.6, 102563.4, 102664.5, 102766.4, 102765.1, 102582.2, 
    96494.87, 95716.64, 102013, 101985, 101736.5, 101560.8, 101370.7, 101235,
  102477.6, 102521, 102521.8, 102627.3, 102646.2, 102721.8, 102721.7, 
    102586.9, 102305.2, 102262.1, 102017.9, 101794.9, 101615.7, 101452.8, 
    101301.1,
  102524.4, 102561.3, 102541.3, 102528.1, 102511.8, 102569.1, 102598.9, 
    102644.5, 102528, 102294.8, 102066, 101851.9, 101672, 101513.8, 101355.5,
  102550, 102589.8, 102565.1, 102523.6, 102421.1, 102451.9, 102535.4, 
    102579.2, 102465.4, 102317.9, 102110.7, 101914.2, 101742.6, 101577.2, 
    101408.3,
  102649, 102673.8, 102629.8, 102540.4, 102457.7, 102467.9, 102577.2, 
    102627.6, 102524.9, 102352.9, 102162.7, 101984.1, 101819.2, 101649.9, 
    101476,
  102725.1, 102720.4, 102634.7, 102537.4, 102482.2, 102532.9, 102646.4, 
    102610.6, 102483, 102330.4, 102202.8, 102055.4, 101903, 101748.7, 101582.8,
  101833, 101970.3, 102120.3, 102248.6, 102396.9, 102488.8, 102456.4, 
    102410.6, 102312, 101793.9, 101636.4, 101635.6, 101261, 100630.1, 100303.9,
  102035.4, 102151, 102319.2, 102421.3, 102537.6, 102352, 102577.3, 102386.5, 
    102265.5, 102115.4, 101889.5, 101663.5, 101410.1, 99384.85, 99838.89,
  102200.7, 102386.9, 102478.5, 102596.9, 102473.3, 99110.44, 102404.7, 
    102552.1, 102402.8, 102184.4, 101893.9, 101665, 101415.3, 101248.5, 
    101003.1,
  102372.7, 102546.1, 102624.4, 102710.7, 102723.1, 102482.6, 98773.98, 
    102214.2, 102237.7, 102191.3, 101916.9, 101665.2, 101431.1, 101257.4, 
    101060.1,
  102571, 102703.2, 102775.7, 102790.5, 102821.2, 102787.9, 102539.8, 
    96445.09, 95705.38, 101978.4, 101961.9, 101674.4, 101471.6, 101263.5, 
    101127.3,
  102688.5, 102808.8, 102842.5, 102855.9, 102797.1, 102784.7, 102746.2, 
    102578.5, 102243.2, 102211.4, 101969.4, 101720.6, 101517.6, 101316.3, 
    101161.6,
  102835.9, 102960.5, 102993.2, 102975.9, 102923.1, 102852.9, 102738.8, 
    102633.2, 102462.7, 102233.8, 101994.5, 101774.5, 101567.7, 101380, 
    101197.5,
  102971.9, 103072.8, 103106.6, 103090.4, 103018.4, 102944.3, 102820.2, 
    102626.1, 102409.2, 102245.3, 102038.4, 101829.2, 101634.8, 101454.8, 
    101257.6,
  103081.4, 103182.9, 103222.6, 103211.2, 103157.9, 103040, 102854.8, 
    102671.9, 102481.3, 102284.7, 102090.6, 101892.3, 101700.5, 101526.3, 
    101315.8,
  103191.6, 103289.8, 103310.9, 103295.9, 103221, 103100.4, 102910.2, 
    102690.3, 102488.4, 102286.9, 102148.4, 101961.3, 101773.1, 101598.6, 
    101382.2,
  102378.7, 102533.3, 102641, 102658.9, 102650.9, 102591.4, 102508.7, 
    102420.9, 102270.1, 101728.3, 101566.9, 101588.8, 101232.2, 100634.9, 
    100333.6,
  102562.6, 102680.5, 102745.9, 102750.6, 102684.9, 102428.9, 102552.3, 
    102318.9, 102133.9, 101999.6, 101792.9, 101587.4, 101366.7, 99356.46, 
    99814.4,
  102686.9, 102820.5, 102854.4, 102870.3, 102622.5, 99134.75, 102324.9, 
    102486.7, 102270.8, 102018.4, 101764.2, 101567.6, 101345.4, 101171.3, 
    100933.5,
  102769.8, 102892.9, 102940.6, 102919.4, 102848.3, 102482.1, 98689.25, 
    101991.1, 102018.7, 101998.7, 101748.2, 101524.4, 101309.1, 101122.2, 
    100896.9,
  102843.5, 102982.3, 103014.8, 102981.5, 102880.9, 102740.8, 102397, 
    96307.66, 95506.45, 101721.6, 101744.3, 101469.1, 101259.1, 101024.1, 
    100840.8,
  102908.5, 103038, 103070.6, 103036.9, 102882, 102725, 102552.3, 102296.7, 
    101956.1, 101935.2, 101697.1, 101439.4, 101204.5, 100963.9, 100754.2,
  102980.9, 103134.6, 103152.1, 103077.8, 102924.3, 102737.1, 102530, 
    102387.3, 102182.1, 101925.1, 101682.3, 101427.3, 101166.1, 100934.9, 
    100709.9,
  103061.1, 103183.7, 103184.1, 103096.1, 102925.5, 102746.6, 102544.6, 
    102324.8, 102107.6, 101922.2, 101698.9, 101432.8, 101183.5, 100951.3, 
    100731.9,
  103160.2, 103250.3, 103235.8, 103136.9, 102987.4, 102784.6, 102583.4, 
    102399.4, 102189.5, 101959.9, 101731.2, 101482.1, 101233.7, 101008.6, 
    100792.7,
  103243.3, 103282, 103240.3, 103141.8, 102996.5, 102808.3, 102614.3, 
    102387.3, 102166.4, 101950.6, 101779.5, 101555.3, 101323.5, 101111.8, 
    100906.5,
  102545.3, 102625.7, 102651.2, 102601.7, 102535.5, 102438.8, 102322.2, 
    102220.7, 102098.2, 101613.5, 101523.3, 101610.2, 101284.3, 100687.3, 
    100407.2,
  102689.2, 102724.3, 102715, 102639.9, 102524.4, 102193.9, 102327.1, 
    102080.5, 101923.9, 101850.4, 101693.2, 101539.8, 101326.9, 99316.32, 
    99790.8,
  102762.4, 102809.8, 102767.3, 102707.3, 102425.2, 98894.34, 102043, 
    102208.3, 102007.3, 101831.7, 101627.5, 101437.6, 101207.8, 101034.5, 
    100842.6,
  102808.4, 102854.1, 102797.8, 102705.6, 102576.9, 102202.9, 98410.48, 
    101716.9, 101810.7, 101773.1, 101565.7, 101331.2, 101118.9, 100949.9, 
    100773.9,
  102860.1, 102889.5, 102833.2, 102739.1, 102590.9, 102429.6, 102090.1, 
    96032.2, 95217.23, 101489.6, 101517.2, 101243, 101051.5, 100875.7, 
    100754.5,
  102886.3, 102911, 102841.1, 102738.6, 102548.3, 102392, 102222, 101976.9, 
    101648.9, 101655.6, 101422.6, 101188, 101014.5, 100854.9, 100709.7,
  102908, 102930.6, 102850.8, 102737.7, 102565.8, 102363.7, 102152.3, 
    101993.4, 101793.4, 101560.4, 101343.8, 101148.6, 100978.2, 100828.2, 
    100669.4,
  102933, 102915.8, 102824.4, 102694.2, 102508, 102317.1, 102089.7, 101844.1, 
    101631.3, 101468, 101280.9, 101110.9, 100960.6, 100807.2, 100645.2,
  102965.8, 102918, 102807.1, 102679.3, 102520.8, 102286.6, 102034.1, 101808, 
    101600, 101389.7, 101214.2, 101069.5, 100925.9, 100784.2, 100623.2,
  102981.1, 102881.7, 102743.5, 102621.3, 102441.4, 102220.8, 101962.7, 
    101681.3, 101446, 101249.8, 101135.1, 101022.7, 100894, 100769.2, 100616.7,
  102739.4, 102803.9, 102785.6, 102696, 102591.6, 102456.5, 102310.8, 
    102202.3, 102095.1, 101622.5, 101590.9, 101749.5, 101507.2, 100990.6, 
    100755,
  102827.7, 102825.4, 102777.6, 102676.7, 102529.8, 102164.8, 102290.9, 
    102022.3, 101866.8, 101826.2, 101742.1, 101690.3, 101597.1, 99667.88, 
    100217.5,
  102843.3, 102848.2, 102758.8, 102667.2, 102360.8, 98842.12, 101899.6, 
    102105.2, 101873.7, 101709.4, 101610, 101584, 101512, 101463.5, 101343.9,
  102835.9, 102819.2, 102711.7, 102570, 102425.3, 102019, 98253.02, 101427, 
    101549, 101560, 101473.2, 101419.8, 101389.6, 101372.6, 101314.6,
  102835.5, 102786.9, 102657.9, 102504, 102336.7, 102138.1, 101758.1, 
    95761.35, 94883.77, 101118.8, 101322.9, 101240.8, 101239, 101215.6, 
    101234.5,
  102790.9, 102722.8, 102563.9, 102415.5, 102194.3, 101996.9, 101769.3, 
    101463.5, 101135.2, 101195.9, 101093, 101046.2, 101052.6, 101060.6, 
    101094.8,
  102746.4, 102668.3, 102506.2, 102351, 102149.3, 101890.1, 101623.1, 
    101413.5, 101191.5, 100987.6, 100887.7, 100857, 100851.5, 100881.6, 
    100923.3,
  102713.9, 102601.3, 102436.7, 102277.5, 102055.6, 101813, 101536.1, 
    101245.3, 101015.6, 100876.9, 100764.1, 100695.4, 100688.3, 100719.3, 
    100770.2,
  102706.8, 102580.5, 102433.3, 102273.7, 102070.2, 101792.6, 101505.6, 
    101255.8, 101018.9, 100816.3, 100675.2, 100599.9, 100562.8, 100569.9, 
    100614,
  102716.8, 102552.4, 102399.1, 102247.1, 102044, 101792.2, 101524.6, 
    101236.8, 100989.2, 100778.3, 100658.2, 100558.8, 100494.2, 100480.8, 
    100498.5,
  102197.2, 102317.1, 102352, 102277.3, 102161, 102027.9, 101877.3, 101781.4, 
    101703.3, 101268.9, 101286.1, 101546.2, 101420.9, 101053, 100899,
  102314.2, 102356.9, 102312.4, 102194, 102044.4, 101695.4, 101810.5, 
    101580.7, 101453.5, 101427.5, 101385.9, 101438.2, 101504.9, 99724.75, 
    100390.6,
  102352.7, 102356.5, 102244.2, 102148.5, 101847.9, 98380.82, 101438.4, 
    101608.8, 101399.5, 101287.2, 101245.7, 101294.9, 101406.8, 101505.2, 
    101543.6,
  102350, 102304.4, 102188.9, 102057.5, 101913.6, 101535.9, 97814.47, 
    101063.8, 101206.1, 101196.2, 101152, 101171, 101286.1, 101445, 101551.5,
  102353.8, 102277.1, 102173, 102039, 101874.5, 101669.4, 101336.9, 95409.26, 
    94594.52, 100873, 101068.6, 101054.4, 101178.8, 101323.4, 101527.5,
  102315.6, 102255.9, 102151.6, 102008.5, 101764.5, 101563.8, 101359.6, 
    101136.2, 100901.3, 101016.7, 100955.3, 100965.5, 101069.4, 101251.3, 
    101459.5,
  102313.5, 102277, 102180.8, 102002.5, 101761.7, 101482.8, 101236.9, 
    101094.4, 100990.3, 100905.5, 100861.4, 100889.1, 100983.8, 101179.3, 
    101395.6,
  102337.3, 102280.8, 102178.1, 101969, 101688.4, 101413.9, 101142.2, 
    100913.9, 100819.4, 100828.3, 100795.9, 100828.4, 100929.8, 101135.6, 
    101365.8,
  102375.3, 102325.8, 102222.4, 102020.1, 101747.8, 101419.5, 101105.4, 
    100886.1, 100774.8, 100752.6, 100732.6, 100790.6, 100910, 101119.4, 
    101350.7,
  102417, 102338.6, 102222, 102020.3, 101729.8, 101436.1, 101123.3, 100835.9, 
    100671.6, 100638.4, 100695.7, 100765.4, 100930.2, 101144, 101366.1,
  101463.9, 101510.6, 101502.7, 101430.9, 101366.5, 101287.7, 101197.1, 
    101183.2, 101216.3, 100906.8, 101026.6, 101369.9, 101317, 100971.5, 
    100816.5,
  101600.9, 101564.3, 101508.9, 101415.9, 101309.3, 100984.9, 101164, 
    101066.6, 101077.2, 101144.1, 101206.3, 101353.4, 101482.9, 99731.84, 
    100406,
  101639.7, 101584.6, 101498.5, 101408.9, 101116, 97678.57, 100791, 101041.7, 
    101013.2, 101096.9, 101171.3, 101331.5, 101514.8, 101609.4, 101624.1,
  101650.6, 101586.2, 101487.5, 101339.7, 101148.2, 100798.6, 97138.27, 
    100625.9, 100940.7, 101034.7, 101168.8, 101321.4, 101526.7, 101687.4, 
    101748.6,
  101667.2, 101603.9, 101486, 101292.4, 101092.6, 100885.2, 100649.7, 
    94860.59, 94341.12, 100818.5, 101201.4, 101346.1, 101570.7, 101706.1, 
    101839.8,
  101680.6, 101618.9, 101473.6, 101282.8, 101023.9, 100849.4, 100724.9, 
    100722.9, 100676, 101064.3, 101213.8, 101409.4, 101617.4, 101796.2, 
    101913.1,
  101713, 101660.9, 101512.4, 101320.6, 101104.5, 100914.8, 100784.1, 
    100845.7, 101003.2, 101141.3, 101292.9, 101489.4, 101682, 101869.4, 
    101995.1,
  101759.7, 101704.4, 101569.6, 101398.1, 101198.4, 101048.8, 100959.1, 
    100970.3, 101085.1, 101251.1, 101392.6, 101576.6, 101779, 101969.4, 
    102114.4,
  101836, 101794.9, 101681.4, 101532, 101382.1, 101247.4, 101168.7, 101206.3, 
    101293.7, 101386.8, 101510.3, 101690.7, 101888.7, 102073.1, 102211.9,
  101924, 101876.4, 101786.7, 101657.2, 101514.8, 101419.8, 101368.2, 
    101363.1, 101404.2, 101465.1, 101631.3, 101820.6, 102017.9, 102196.3, 
    102326.1,
  101312.4, 101355.5, 101349.5, 101294.5, 101245.3, 101189.4, 101130.8, 
    101160.5, 101208.1, 100926.8, 101063.5, 101387.3, 101252.7, 100801.9, 
    100519.9,
  101341.6, 101325.7, 101315.5, 101242.1, 101171.1, 100891.9, 101073.8, 
    101053.6, 101116.6, 101210.6, 101306.1, 101434.8, 101436.2, 99557.81, 
    100081.8,
  101308.2, 101301.8, 101267.7, 101211.6, 100986.6, 97581.09, 100830.6, 
    101059.8, 101143.9, 101230.4, 101322.4, 101451.5, 101482.6, 101445.3, 
    101250.9,
  101267.4, 101295.6, 101246.7, 101170.8, 101044.4, 100817, 97192.12, 
    100859.1, 101113.1, 101237.5, 101381.5, 101479, 101522.8, 101485, 101334.2,
  101282.9, 101313.2, 101263.1, 101152.5, 101061.9, 100999.1, 100872.9, 
    95116.43, 94628.09, 101109.4, 101454.1, 101517.8, 101551.5, 101475.9, 
    101421.2,
  101317, 101356.7, 101302.7, 101214.6, 101094.8, 101041.5, 101053.8, 
    101089.3, 101017.4, 101395.7, 101506.1, 101592.8, 101597.6, 101566.4, 
    101512,
  101368.6, 101436.5, 101386.3, 101323.9, 101245, 101213.8, 101197.9, 
    101314.3, 101442.2, 101523.4, 101611.9, 101673.7, 101688.6, 101695.1, 
    101675,
  101464.8, 101522.1, 101495.1, 101449.3, 101383.6, 101371, 101390.2, 
    101436.2, 101521.5, 101658, 101756.2, 101818.9, 101863.6, 101880, 101873.9,
  101579.3, 101626.4, 101617.6, 101592, 101573.4, 101569.7, 101592.8, 
    101686.6, 101782.8, 101872, 101946, 102017.2, 102049.1, 102069, 102050.6,
  101703.1, 101737.1, 101739.7, 101733.9, 101724.2, 101748.4, 101799.7, 
    101851.7, 101923.8, 102004.1, 102138.2, 102222.4, 102260, 102292.5, 102268,
  100584.6, 100766.2, 100936.7, 101082.4, 101240.6, 101345.9, 101396.4, 
    101475.2, 101512.3, 101176.1, 101229.3, 101535.7, 101366.2, 100875.7, 
    100573.7,
  100686.9, 100855.5, 101021.3, 101148.5, 101237.5, 101127.9, 101364, 
    101386.9, 101436.3, 101502.7, 101500.5, 101585, 101546.3, 99638.54, 
    100117.3,
  100770.9, 100962.6, 101091.4, 101202.4, 101131, 97799.85, 101121, 101396.9, 
    101417, 101497, 101517.8, 101576.1, 101560.7, 101480.2, 101259,
  100860.4, 101052.9, 101128.6, 101206.6, 101217.9, 101063.3, 97465.11, 
    101076.2, 101392.7, 101454, 101516.7, 101539.9, 101533.2, 101444.6, 
    101248.2,
  100980.1, 101133.1, 101182.8, 101203.7, 101225.2, 101240.2, 101089.1, 
    95349.53, 94737.65, 101215.1, 101494.9, 101499.4, 101470.9, 101333.4, 
    101217.7,
  101109.8, 101217.2, 101223.9, 101231.2, 101155.3, 101181, 101220.6, 101207, 
    101110.2, 101408.1, 101438.7, 101449.1, 101392.7, 101270.5, 101193.3,
  101242.4, 101305.2, 101308.7, 101289.9, 101264.2, 101244.1, 101249.3, 
    101343.4, 101381, 101391.7, 101417.8, 101402.8, 101315.3, 101257.7, 
    101241.5,
  101357.2, 101394.1, 101378.1, 101346.1, 101300.8, 101313.1, 101322.8, 
    101319.9, 101320.8, 101354.9, 101357.4, 101341.4, 101319.3, 101333.2, 
    101360.2,
  101484.9, 101507.5, 101486, 101451, 101423.6, 101391.7, 101371.4, 101395.2, 
    101392.4, 101361.8, 101348.7, 101364.2, 101386.5, 101435.5, 101482.9,
  101637.7, 101642.9, 101618.7, 101564.9, 101499.6, 101475.9, 101466.3, 
    101441.8, 101401.5, 101371.4, 101426.5, 101470.4, 101517.1, 101585.6, 
    101640.8,
  99784.87, 99978.18, 100173.3, 100477.2, 100802.9, 101098.9, 101370.5, 
    101584.5, 101747.9, 101488.9, 101593, 101841.3, 101625.4, 101152.5, 
    100864.9,
  99882.52, 100080.4, 100322.7, 100653.7, 100948, 101118, 101488.6, 101670.8, 
    101775.4, 101877.7, 101878.3, 101923.8, 101849.3, 99891.12, 100352.3,
  100059, 100279.6, 100524.7, 100825.1, 100931.1, 97921.99, 101442.1, 101820, 
    101865.6, 101934, 101953.7, 101918.4, 101843.6, 101722.2, 101460.7,
  100301.1, 100517.3, 100726.6, 100961, 101175.8, 101105.3, 97816.82, 
    101478.3, 101846.7, 101920.3, 101926, 101876.1, 101802.3, 101648, 101372.2,
  100586.9, 100760.7, 100930.3, 101114, 101302.7, 101480.7, 101351.4, 
    95775.01, 95137.41, 101638.5, 101886.8, 101832.2, 101742.9, 101514.3, 
    101331.1,
  100852.1, 100976, 101078, 101226, 101306.9, 101459.4, 101604.5, 101574.5, 
    101552.2, 101812.1, 101834.7, 101798.5, 101651.7, 101442.7, 101298.6,
  101069.4, 101152.7, 101221.7, 101296.2, 101390.5, 101466.5, 101562.9, 
    101725.9, 101794.8, 101808.9, 101836.2, 101749.9, 101559.3, 101418.9, 
    101367.8,
  101190.8, 101232.3, 101281.8, 101332.2, 101362.5, 101468.5, 101571.8, 
    101654.7, 101773.4, 101849.7, 101801.1, 101668.3, 101530.1, 101489.8, 
    101495.9,
  101247.4, 101283.1, 101308.9, 101345.5, 101405.8, 101476, 101579.8, 
    101718.9, 101820.4, 101799.2, 101733.2, 101622.6, 101581, 101596.4, 
    101632.2,
  101296.2, 101269.5, 101271.4, 101304.1, 101349.6, 101451.9, 101572.1, 
    101658, 101715.2, 101695.5, 101665.6, 101653.9, 101673, 101741.7, 101816.2,
  99731.52, 99891.48, 100076.9, 100314.5, 100573.1, 100858, 101200.4, 
    101488.7, 101759, 101628, 101865.1, 102204.2, 102092, 101677.7, 101480,
  99728.07, 99909.41, 100128.7, 100440.5, 100732.3, 100940.1, 101400.3, 
    101673.8, 101865.8, 102096.3, 102238.6, 102342.6, 102337.3, 100418.9, 
    100995.6,
  99741.09, 99963.86, 100242.2, 100593.1, 100741.7, 97939.48, 101533.4, 
    101933.4, 102134.2, 102257.6, 102348.2, 102378.6, 102349.4, 102285.4, 
    102130.8,
  99794.8, 100051, 100377.7, 100705, 101046.6, 101052, 98035.19, 101790.4, 
    102220.4, 102323, 102367.9, 102352.3, 102291, 102167.4, 102039.9,
  99919.41, 100200.9, 100542.1, 100893.7, 101234.4, 101623.4, 101542.2, 
    96093.52, 95571.13, 102115.8, 102369.6, 102289.4, 102174, 101992.8, 
    101925.8,
  100109, 100388.8, 100710.4, 101078, 101382.2, 101714.7, 101967.6, 101954.2, 
    102022, 102336.8, 102358.3, 102219.6, 102042.4, 101886.7, 101824.6,
  100374.4, 100635.9, 100940.9, 101266.3, 101582.1, 101844.6, 102040.1, 
    102288.9, 102406.5, 102408.3, 102330.5, 102150.9, 101988.3, 101880.1, 
    101850,
  100669.8, 100897.6, 101170.3, 101450.6, 101723.6, 101967.2, 102164.2, 
    102292.7, 102388, 102415, 102290.2, 102118.2, 102019.1, 101962.5, 101959.2,
  100958.9, 101184.7, 101426.9, 101671.1, 101898.5, 102115, 102305.6, 
    102452.3, 102519.1, 102412.3, 102274.3, 102140.8, 102072.5, 102050.2, 
    102050.4,
  101183, 101369.2, 101590.4, 101815.8, 102025.4, 102224.5, 102395.4, 
    102460.3, 102458, 102362.6, 102257.7, 102173.1, 102151.4, 102157.2, 
    102177.6,
  99498.84, 99540.32, 99690.33, 99911.15, 100177.7, 100435.4, 100699, 
    100991.4, 101303.4, 101290.6, 101641.5, 102119.7, 102142.9, 101853.2, 
    101701.5,
  99416.8, 99465.38, 99643.88, 99911.36, 100188.5, 100360.5, 100779.7, 
    101088.6, 101363.7, 101696, 101964.5, 102232.4, 102354.5, 100597.8, 
    101250.7,
  99454.24, 99553.34, 99754.52, 100047.6, 100191.4, 97389.22, 100920, 
    101355.1, 101620.6, 101864.8, 102092.5, 102302.5, 102422.4, 102482.5, 
    102451.5,
  99645.58, 99756.89, 99977.18, 100223.8, 100539.1, 100538.1, 97604.85, 
    101321.4, 101812.3, 102033.6, 102205.7, 102337.1, 102431.8, 102459.1, 
    102432.8,
  99883.91, 100042.9, 100260.7, 100530.7, 100813.6, 101176.7, 101068.6, 
    95778.59, 95353.21, 101886.8, 102297.6, 102324.5, 102358.8, 102287, 
    102287.7,
  100135.6, 100322, 100526.2, 100816.1, 101051.3, 101327.5, 101537, 101499.9, 
    101617.8, 102157.8, 102239.8, 102262.3, 102203.4, 102116, 102085.6,
  100353.2, 100582, 100822.2, 101079.5, 101345, 101575.6, 101739.3, 102010.7, 
    102179.4, 102189.7, 102204.1, 102168.5, 102087.1, 102044.2, 102046.5,
  100572.8, 100830.6, 101073.6, 101342.1, 101553.6, 101783.4, 101936.7, 
    102024.7, 102112.5, 102198.8, 102180.1, 102151, 102108.2, 102098.1, 
    102117.8,
  100812.1, 101106.8, 101402.6, 101663.3, 101875.3, 102040.2, 102171.6, 
    102284.6, 102307.5, 102257, 102230.6, 102193.7, 102155.6, 102147.7, 
    102151.7,
  101088.8, 101377.4, 101647.8, 101883.8, 102078.4, 102231.7, 102317.2, 
    102322.2, 102314.8, 102284.2, 102299.1, 102264, 102226.5, 102237.5, 
    102266.5,
  100085.2, 100252.1, 100392.1, 100534.5, 100526.9, 100552.3, 100575.1, 
    100613.8, 100703.3, 100607.2, 100936.1, 101490.8, 101660.2, 101486.9, 
    101462.5,
  99837.4, 100043, 100260.1, 100453.3, 100512.7, 100464.5, 100670.9, 
    100671.7, 100727, 100931.8, 101195, 101529.7, 101838.8, 100269.2, 101044.4,
  99583.05, 99854.16, 100141.8, 100395.8, 100423.2, 97317.74, 100583.8, 
    100787.1, 100827.7, 100954.1, 101233.6, 101551.9, 101886.3, 102072.9, 
    102259.3,
  99487.93, 99753.48, 100068.7, 100302.8, 100531.6, 100391.9, 97119.81, 
    100541.5, 100870.5, 101021.9, 101289.6, 101593.7, 101942.3, 102189.7, 
    102356.9,
  99647.86, 99857.3, 100104.9, 100340.2, 100528.6, 100713.7, 100575.7, 95100, 
    94601.23, 100930, 101397.3, 101661.9, 101983, 102180.7, 102375.9,
  99931.93, 100077.6, 100235.4, 100435.4, 100562.9, 100696.4, 100823.5, 
    100769.9, 100779.4, 101265.3, 101491.6, 101775.2, 102049.9, 102225.2, 
    102344.9,
  100271.8, 100364.1, 100470.7, 100610, 100731.7, 100850.9, 100954.2, 
    101178.8, 101359.8, 101471.8, 101685.7, 101918, 102074.2, 102184.8, 
    102252.5,
  100623.2, 100683.9, 100759.1, 100867.2, 100971.2, 101105.6, 101230.5, 
    101343, 101498.5, 101693, 101860.5, 101986.9, 102092.8, 102172.7, 102220.8,
  100977.3, 101051.1, 101128.2, 101221.3, 101321.4, 101427.5, 101543.1, 
    101686.3, 101801.1, 101879.5, 101965.2, 102047.5, 102111.5, 102168.4, 
    102177.1,
  101295.9, 101361.4, 101436.2, 101517.8, 101603.6, 101703.7, 101793.7, 
    101855.1, 101911.7, 101965.3, 102063.6, 102133, 102199.5, 102246.3, 
    102221.6,
  100281.9, 100398.7, 100434.2, 100493.5, 100458, 100391.4, 100417.3, 
    100509.5, 100686.2, 100502.1, 100695.2, 101081.3, 101144, 100953.5, 
    100959.6,
  100365.1, 100445.3, 100467.3, 100481.6, 100338, 100108.2, 100286.9, 
    100388.9, 100527.5, 100714.9, 100914.1, 101151.5, 101354.7, 99800.48, 
    100588.6,
  100470.2, 100503.7, 100485.9, 100452.4, 100140.1, 96855.13, 100087.9, 
    100366.5, 100541.4, 100696, 100916.5, 101172.6, 101445.5, 101613.4, 
    101824.3,
  100550.3, 100538.9, 100507, 100375.7, 100283.6, 99891.65, 96655.41, 
    100097.8, 100483.6, 100670.7, 100944.6, 101207.8, 101529.4, 101803, 
    102008.4,
  100633, 100600.1, 100526.8, 100423.3, 100273.9, 100308.7, 100029, 94661.88, 
    94225.52, 100501.9, 101006.6, 101266.5, 101596.8, 101841.1, 102117.6,
  100726.4, 100689.4, 100596.2, 100511.7, 100377.8, 100339.4, 100459.8, 
    100372.7, 100298.5, 100785.5, 101037.9, 101357.5, 101676.5, 101956.7, 
    102202.9,
  100850.4, 100810.6, 100737.9, 100640.7, 100561.5, 100507.2, 100505.3, 
    100673.4, 100805.7, 100905, 101148.8, 101472.9, 101780.8, 102056.1, 
    102266.6,
  101017.7, 100994.1, 100933.1, 100869.7, 100793.3, 100774.8, 100788.4, 
    100796.9, 100894.9, 101114.5, 101373.1, 101653.8, 101927.1, 102174.4, 
    102372.1,
  101274.7, 101275.8, 101252.4, 101217.2, 101186.8, 101158.7, 101173.8, 
    101261.9, 101358.4, 101462.9, 101638, 101859.3, 102077.9, 102277.9, 
    102435.6,
  101555.4, 101557.8, 101554.5, 101535.3, 101515.5, 101516, 101526.2, 
    101532.8, 101589.6, 101691.6, 101881.9, 102054.1, 102216.3, 102371.9, 
    102494.8,
  100870.9, 100800.7, 100735.2, 100731.2, 100781, 100861, 100939.9, 101079.4, 
    101236.3, 101086.4, 101146.4, 101393.4, 101308.4, 101085.1, 101062.1,
  100825.7, 100698.7, 100615.4, 100617.6, 100619.6, 100600.5, 100879.5, 
    100982.3, 101121.9, 101365.4, 101399.2, 101449.4, 101487.2, 99893.2, 
    100640.5,
  100701.2, 100515.7, 100412.6, 100407.3, 100384.5, 97252.24, 100637, 
    101027.7, 101184.6, 101357.4, 101410.7, 101469.2, 101551.8, 101654.2, 
    101794.3,
  100590.2, 100349.1, 100183.4, 100102.9, 100270.5, 100195.5, 97044.02, 
    100624.8, 101087.5, 101337.1, 101434.1, 101476.7, 101574.9, 101742.4, 
    101922.5,
  100507.8, 100204.1, 99935.44, 99800.12, 99932.91, 100318.4, 100295.7, 
    95090.31, 94688.66, 101053.1, 101438.4, 101493.9, 101597.8, 101736.7, 
    101997.5,
  100488.7, 100119.1, 99761.2, 99542.89, 99644.96, 100059.7, 100479.5, 
    100577.1, 100662.1, 101247, 101364.4, 101496.1, 101628.5, 101803.2, 
    102060.5,
  100553.1, 100158.3, 99775.06, 99536.68, 99627.58, 100017.7, 100377.3, 
    100810.7, 101077.8, 101205.7, 101332.4, 101502.1, 101654, 101848.6, 
    102094.3,
  100711.3, 100336.1, 99953.31, 99715.39, 99765.62, 100113.8, 100429.7, 
    100659.2, 100880, 101161, 101341.1, 101520.1, 101712.8, 101925.2, 102185.7,
  100948.6, 100632.8, 100309.5, 100106.3, 100127.4, 100327, 100564.5, 
    100856.5, 101072.3, 101235.9, 101385.4, 101579.3, 101782.5, 102016.1, 
    102266.3,
  101215.8, 100967.9, 100696.3, 100511.7, 100481.4, 100603.8, 100762.8, 
    100913.7, 101070.9, 101254.8, 101469.8, 101677.4, 101893.7, 102144.7, 
    102358.9,
  101538.9, 101510.4, 101470.2, 101415.4, 101379.1, 101327.8, 101271.7, 
    101237.8, 101190.2, 100857.3, 100882.5, 101112.5, 100943.4, 100581.6, 
    100484.9,
  101450, 101364.8, 101301.8, 101234.8, 101173.5, 100992.3, 101171.4, 
    101104.1, 101046, 101090.6, 101079.9, 101090.7, 101079.1, 99362.9, 
    100059.2,
  101276.9, 101159, 101067.1, 101003.5, 100870.1, 97574.2, 100821.9, 
    101092.1, 101040.6, 101038.9, 101051, 101038, 101085.4, 101139.3, 101248.2,
  101089.3, 100924.4, 100791.3, 100709.5, 100730.1, 100586.5, 97187.71, 
    100636.3, 100916.5, 100992.6, 101037, 100998, 101086.9, 101228.3, 101415.9,
  100869.7, 100667, 100492, 100422.9, 100449.6, 100599.1, 100538.4, 95047.64, 
    94478.2, 100732.5, 101033, 100987, 101117.2, 101278.7, 101568.7,
  100660, 100404.2, 100182, 100108.3, 100156.9, 100339.2, 100604.6, 100651.3, 
    100582.8, 100958.8, 100973, 101015.6, 101183.4, 101406.8, 101677,
  100486.8, 100182.1, 99915.42, 99842.87, 99958.57, 100184, 100458.7, 
    100773.6, 100901.2, 100955.3, 100971.4, 101085.4, 101267.5, 101494.1, 
    101758.2,
  100405.2, 100066.2, 99777.13, 99684.27, 99828.88, 100134.6, 100437.8, 
    100650.3, 100780.3, 100965.2, 101033.4, 101172.4, 101374, 101607, 101888.4,
  100442.7, 100131.4, 99868.57, 99805.91, 99963.35, 100229.9, 100503.5, 
    100745.6, 100923.1, 101037.6, 101126.6, 101281.6, 101482, 101730.8, 
    102001.2,
  100589.2, 100340.1, 100145.2, 100088.7, 100197.9, 100405.4, 100623.4, 
    100791.4, 100956.8, 101069.3, 101226.7, 101394.4, 101596.1, 101859.9, 
    102101.9,
  101536.8, 101595, 101651.8, 101697.7, 101768.9, 101794.5, 101813, 101836.1, 
    101848.9, 101491, 101487.6, 101632.9, 101364, 100796.5, 100469.2,
  101464.8, 101495.7, 101533.9, 101565.4, 101584, 101446.9, 101665.7, 
    101624.4, 101588.2, 101618.8, 101564.2, 101522.6, 101417.1, 99498.52, 
    99951.44,
  101432.1, 101435.6, 101426.2, 101428.5, 101313.9, 98050.13, 101229, 
    101538.2, 101444.6, 101424.9, 101383.8, 101367.3, 101297.5, 101218.9, 
    101056.5,
  101371.2, 101299, 101221.9, 101164.7, 101157.4, 100985.6, 97541.16, 
    100923.6, 101236.8, 101242.8, 101228.6, 101194.4, 101178.5, 101137.4, 
    101068.6,
  101184.8, 101056.6, 100928.9, 100847.6, 100840.3, 100908.9, 100820, 
    95263.77, 94535.41, 100845.7, 101098.6, 101075.5, 101076, 101043, 101102.4,
  100966.5, 100783.3, 100608.5, 100514.5, 100483.9, 100567.4, 100737.2, 
    100763.7, 100762.6, 101033.4, 101018.8, 101011.8, 100997.1, 101044.2, 
    101141.2,
  100760.6, 100554.2, 100375.7, 100254.7, 100247, 100332.2, 100489, 100731.1, 
    100871.1, 100881.1, 100908, 100900.1, 100946.8, 101064.6, 101236.2,
  100641.7, 100442.2, 100237, 100097.1, 100065.1, 100193.9, 100369, 100535.4, 
    100673.7, 100781.1, 100786.3, 100837.7, 100975.3, 101168.5, 101419.7,
  100620.5, 100436.4, 100257.8, 100145.6, 100146.1, 100227.6, 100382.7, 
    100560.1, 100653.9, 100678, 100723.8, 100885.9, 101089.3, 101346.7, 
    101596.5,
  100674.2, 100506.5, 100350.3, 100254.9, 100243.4, 100326.9, 100438.3, 
    100514.1, 100556.3, 100595.3, 100787.4, 101024.4, 101271.3, 101540.4, 
    101763.1,
  100524.3, 100731.4, 100935, 101139.3, 101342, 101502.1, 101676.1, 101855.2, 
    101988.6, 101746.2, 101896.1, 102168.3, 101989.8, 101411.2, 101014.7,
  100529.4, 100727.6, 100921.6, 101129.1, 101306.6, 101362.6, 101690.6, 
    101810.6, 101934.9, 102086.4, 102140.6, 102167.1, 102065.3, 100097.2, 
    100424.4,
  100647.7, 100841.9, 101006.7, 101187.3, 101206.2, 98168.18, 101502.4, 
    101902.6, 101943.3, 102025.2, 102078, 102084.4, 102019.6, 101836.3, 
    101503.6,
  100938.5, 101013.9, 101118.8, 101230.8, 101356.5, 101233.5, 97965.94, 
    101429.9, 101872.4, 101964.3, 102030.3, 101989.3, 101972.2, 101824.4, 
    101534.8,
  101132.1, 101147.2, 101181.2, 101244, 101319.2, 101442.3, 101329.5, 
    95872.95, 95229.05, 101599.6, 101941.3, 101919.2, 101957.2, 101809.3, 
    101658.9,
  101139.8, 101121.6, 101113.1, 101146.2, 101170.1, 101246, 101379, 101372.5, 
    101408.3, 101780.6, 101839, 101948.8, 101988.8, 101867.4, 101739.6,
  101066.8, 101024.3, 100993.6, 100994.6, 101025.1, 101072.1, 101156, 
    101377.2, 101557.6, 101666.6, 101802.5, 101956.6, 101986.1, 101922.1, 
    101886.8,
  100953.7, 100887.2, 100820.7, 100805, 100794.1, 100855.4, 100955.7, 
    101090.2, 101317.1, 101574.9, 101764.9, 101938.9, 102005.6, 102005.9, 
    102053.3,
  100845.4, 100750.8, 100667, 100622.1, 100632.5, 100678.6, 100799.5, 101020, 
    101265.1, 101504.4, 101727, 101935.4, 102011.6, 102093.5, 102193.5,
  100731.8, 100566.5, 100448.9, 100424.8, 100473, 100550.5, 100691.4, 
    100887.2, 101155, 101419.5, 101703.8, 101924.4, 102032.4, 102197.9, 
    102327.3,
  100310.5, 100026.7, 99920.98, 99953.88, 100034.6, 100207.8, 100533.8, 
    100878.9, 101208.2, 101180.4, 101525.9, 101957.6, 101896.6, 101469, 
    101215.4,
  100283.8, 100006.5, 99962.85, 100069.2, 100181.4, 100266.9, 100716, 
    101020.2, 101295.5, 101630.1, 101895.9, 102092.6, 102132.7, 100249.5, 
    100764,
  100350.6, 100084, 100060.3, 100220.9, 100256.4, 97364.22, 100841.5, 
    101242.4, 101541.5, 101811.1, 102029.6, 102175.5, 102213, 102127.6, 
    101945.2,
  100533.5, 100213, 100186.9, 100325.9, 100584, 100522.7, 97535.45, 101190.1, 
    101720.8, 101955.4, 102148.1, 102210.9, 102265.7, 102173.5, 102050.9,
  100791, 100432.6, 100336.7, 100500, 100709.5, 101024.3, 101005.7, 95774.62, 
    95384.93, 101835.8, 102230.3, 102263.4, 102310.2, 102221.7, 102202.8,
  101024, 100747, 100559.2, 100694, 100858.5, 101093.6, 101387, 101440.4, 
    101555.2, 102090.6, 102235.8, 102347.4, 102353.9, 102330.7, 102312.7,
  101140.4, 101003.5, 100837, 100897.8, 101048, 101265.1, 101469.6, 101768.4, 
    102006.4, 102141.7, 102296.6, 102417.1, 102432.9, 102467.9, 102480.2,
  101188.5, 101176.8, 101052.6, 101084.1, 101176.1, 101364, 101557.9, 
    101724.4, 101930.5, 102194.9, 102364.3, 102479, 102541.8, 102605.8, 
    102640.5,
  101182.6, 101216.3, 101193, 101202.4, 101287.5, 101439.5, 101627.5, 
    101866.6, 102087.5, 102277.5, 102409.6, 102551.3, 102626.9, 102713.1, 
    102750.3,
  101124.8, 101146.7, 101184.5, 101229, 101314.6, 101459.2, 101647.1, 
    101843.3, 102049.7, 102244.6, 102445.2, 102614.7, 102712.3, 102819.3, 
    102864.9,
  101630.9, 101345.1, 100934.2, 100604, 100380.8, 100376.3, 100438.9, 
    100574.3, 100771.2, 100651.7, 100928.5, 101357.5, 101371.3, 101096.4, 
    101004,
  101642.1, 101369, 101026.7, 100798.7, 100618.6, 100467.5, 100729.5, 
    100859.2, 101020.9, 101229.3, 101417.1, 101617, 101705.9, 99981.74, 
    100673.6,
  101607.6, 101413.9, 101144.7, 101033.1, 100779, 97644.89, 100981, 101256.5, 
    101419.4, 101544.1, 101686.2, 101830.1, 101925.4, 101966.7, 101956.5,
  101565.6, 101446.4, 101236.6, 101175.1, 101233, 100973.5, 97761.55, 
    101328.4, 101644.5, 101797.4, 101919.3, 101991.9, 102079.9, 102130.1, 
    102126.1,
  101514.7, 101464.6, 101291.2, 101304.3, 101381.3, 101554.3, 101335.5, 
    95817.59, 95386.42, 101816.6, 102137.4, 102166.5, 102262.4, 102276.7, 
    102326.5,
  101459.8, 101440.4, 101277.5, 101354.3, 101423, 101557.1, 101694.3, 
    101669.2, 101683.7, 102135.6, 102237.2, 102343.4, 102412, 102457.6, 
    102476.5,
  101415.4, 101418.4, 101272.9, 101334.3, 101483.1, 101648.3, 101740.8, 
    102001.3, 102197.7, 102281.7, 102387.2, 102498.4, 102565.3, 102612.4, 
    102611.5,
  101390.9, 101382.3, 101229.4, 101281, 101445.2, 101665.1, 101856.7, 
    102030.5, 102189.4, 102393.1, 102530.7, 102636.1, 102704.3, 102730.2, 
    102713.2,
  101354.2, 101375.9, 101240.3, 101257.5, 101447.9, 101682.6, 101924.9, 
    102192.2, 102401.7, 102553.1, 102653.9, 102757.9, 102799.5, 102814.1, 
    102771.4,
  101331.4, 101336.8, 101232.5, 101204.6, 101406.6, 101683.9, 101989.2, 
    102233.1, 102430.2, 102562.7, 102742.8, 102844.9, 102897, 102908.2, 
    102854.3,
  101343.5, 101402.8, 101476.3, 101523.1, 101580.6, 101570.3, 101561.9, 
    101583.4, 101615.9, 101339.3, 101465.4, 101748, 101645.1, 101289.6, 
    101157.4,
  101278.5, 101313.8, 101397, 101466.1, 101543.6, 101463.5, 101692.3, 
    101693.8, 101728.6, 101824.8, 101875.3, 101975.7, 101984.9, 100207.9, 
    100863.7,
  101169.4, 101200.2, 101277.5, 101398.2, 101395.7, 98308.05, 101671.3, 
    101939.8, 101968.5, 102004.6, 102066.8, 102144.8, 102201.1, 102220.5, 
    102180.8,
  100985.9, 101023, 101112.8, 101243, 101451.4, 101352.5, 98147.23, 101721.2, 
    102043.6, 102140.7, 102224.4, 102291.7, 102358.1, 102389.8, 102344.7,
  100784.5, 100823.8, 100921.7, 101104.2, 101350.6, 101618.3, 101562.3, 
    96090.59, 95535.07, 102019.1, 102357.1, 102430.7, 102504.4, 102503.7, 
    102515.8,
  100633.5, 100646.7, 100709.6, 100928.6, 101194.7, 101493.2, 101759.1, 
    101758.8, 101761.7, 102267.6, 102406.4, 102541.6, 102601.2, 102619, 
    102581.5,
  100666.8, 100608.4, 100593.3, 100797.8, 101124.2, 101448.3, 101685.3, 
    101984.6, 102192.4, 102335.7, 102489.7, 102625.4, 102668.4, 102671.5, 
    102619.8,
  100830.1, 100697.1, 100601.4, 100730.1, 101052.8, 101420.7, 101698.4, 
    101916.4, 102137.9, 102393.3, 102575.9, 102677.4, 102715.5, 102678.5, 
    102608.7,
  100974.8, 100858.5, 100759.5, 100849.5, 101135.4, 101460.6, 101742.4, 
    102039, 102291.3, 102504, 102641.4, 102733.5, 102738.9, 102688.3, 102604.1,
  101077.8, 100991.2, 100901, 100982.7, 101203.2, 101506.5, 101799.9, 
    102075.6, 102317.5, 102508.9, 102686.8, 102778, 102777.7, 102722.3, 
    102640.3,
  101478, 101580.9, 101633.9, 101641.1, 101612.7, 101610.3, 101631.1, 
    101692.7, 101743.6, 101428.7, 101565.5, 101884.5, 101777.3, 101411.5, 
    101247.8,
  101624, 101688.5, 101720.6, 101704.3, 101611.8, 101434.6, 101651.7, 
    101584.3, 101619.4, 101730.8, 101780.9, 101926.7, 102005, 100225, 100857.4,
  101724.1, 101762.4, 101757.6, 101745.5, 101555.7, 98216.69, 101392.5, 
    101688.4, 101604.2, 101649, 101746.4, 101909.9, 102030, 102098.9, 102095.3,
  101756.8, 101768.8, 101731.3, 101681.6, 101629.4, 101374.4, 97854.8, 
    101170.8, 101519.1, 101627.6, 101721.4, 101869.2, 102042.1, 102156.9, 
    102176,
  101758, 101723.4, 101648.6, 101577.6, 101505.3, 101479.9, 101273.3, 
    95669.16, 94961.65, 101308.2, 101718.5, 101842.1, 102044, 102146.6, 
    102248.6,
  101665.1, 101584.1, 101440.7, 101339.1, 101219.5, 101189.1, 101237.1, 
    101160, 101121.1, 101524.3, 101650.1, 101825.1, 102039.4, 102175.4, 
    102277.2,
  101505.9, 101374, 101190.9, 101031.4, 100902.3, 100861, 100911.6, 101119.2, 
    101272.1, 101379, 101583.2, 101821.3, 102031, 102187.4, 102277.5,
  101316.3, 101127.1, 100867.4, 100618.4, 100412, 100431.1, 100572.9, 
    100753.8, 100987.8, 101284.6, 101553.5, 101813.5, 102045, 102194.8, 
    102280.5,
  101141.8, 100890.5, 100573.1, 100224.5, 99962.23, 100025, 100282.2, 
    100634.2, 100953.9, 101253.6, 101559.3, 101853.6, 102065.2, 102200.3, 
    102277.7,
  100994, 100682.4, 100336.9, 99827.92, 99550.27, 99717, 100089, 100505.1, 
    100901.5, 101259.3, 101623.7, 101919.4, 102098, 102240.8, 102298.5,
  99950.98, 100070.1, 100199.4, 100342.3, 100519.3, 100681.1, 100812.8, 
    100922.8, 100985.9, 100717.7, 100840.4, 101150.5, 101091.2, 100824, 
    100747.9,
  100050.3, 100191, 100356.1, 100545.6, 100706.3, 100759.9, 101028.3, 
    101040.2, 101086.9, 101165.7, 101147, 101169.3, 101204.6, 99537.02, 
    100222.6,
  100389.4, 100507.3, 100636.9, 100778.5, 100728.8, 97604.99, 100966.4, 
    101233.4, 101127, 101134.3, 101145.4, 101161.7, 101190.6, 101263.5, 
    101335.1,
  100733.7, 100822.9, 100907.8, 100996.9, 101049.6, 100867.5, 97425.6, 
    100876.8, 101201.2, 101251.3, 101190.3, 101127.5, 101146.5, 101224.5, 
    101334.3,
  100959.1, 101019.1, 101054.5, 101095.5, 101119.5, 101171, 100992.7, 
    95317.49, 94544.19, 100912.9, 101202.6, 101096.9, 101096.1, 101128.2, 
    101298,
  101073.3, 101087.3, 101061.5, 101058.4, 101011, 101007.6, 101021.4, 
    100930.2, 100874.8, 101154.5, 101145.5, 101107.9, 101078.5, 101108.9, 
    101269.9,
  101074.2, 101059.1, 101000.3, 100943.2, 100863, 100784.4, 100722.1, 100776, 
    100819.8, 100865.2, 100990.5, 101053, 101056.3, 101128.9, 101277.1,
  101040.2, 100992.7, 100888.5, 100774.8, 100624.1, 100491.5, 100381.5, 
    100341.5, 100450.6, 100672.6, 100853.7, 100951.3, 101033.4, 101157.2, 
    101353,
  100998.4, 100911.8, 100770.1, 100629, 100421.5, 100200.6, 100043.5, 
    100051.8, 100189.5, 100409.7, 100669.4, 100859.6, 101006.3, 101209.5, 
    101407.6,
  100938.1, 100789.5, 100645.6, 100508.8, 100247.2, 100024.1, 99886.62, 
    99901.07, 100059.8, 100320.4, 100622.9, 100843, 101057.2, 101297.7, 
    101455.4,
  100641.7, 100469.6, 100307.9, 100128, 100001.4, 99899.73, 99819.97, 
    99800.4, 99833.71, 99581.11, 99682.06, 99976.55, 99872.99, 99568.47, 
    99537.22,
  100505, 100220.2, 99997.21, 99810.05, 99649.8, 99416.02, 99544, 99518.91, 
    99550.71, 99689.34, 99784.98, 99908.25, 99937.49, 98272.73, 98933.01,
  100524.6, 100197.6, 99908.45, 99675.14, 99384.16, 96182.72, 99241.2, 
    99485.16, 99449.77, 99581.41, 99724.73, 99873.55, 99954.83, 99971, 
    100054.4,
  100690.9, 100429.5, 100154.6, 99890.01, 99698.74, 99310.04, 95961.77, 
    99281.3, 99572.81, 99659.34, 99807.8, 99913.59, 100035.6, 100095.5, 
    100157.2,
  100778.1, 100601.8, 100406.8, 100201.5, 100028, 99890.27, 99502.3, 93935.4, 
    93402.2, 99663.23, 100007.6, 100060.9, 100175.2, 100172, 100290.6,
  100853.7, 100714.4, 100542.5, 100372.3, 100172.4, 100060.7, 99984.05, 
    99810.1, 99717.4, 100087, 100164.6, 100251, 100310.7, 100316.9, 100368.9,
  100879.5, 100780.2, 100657, 100505, 100365.1, 100213.4, 100100.9, 100151.1, 
    100171.9, 100180.9, 100269.6, 100375.9, 100398.3, 100399.6, 100434,
  100909.5, 100827.7, 100716.8, 100578.7, 100411, 100293.2, 100188.5, 
    100095.3, 100108.9, 100240.7, 100356.8, 100440.5, 100486.2, 100503.8, 
    100587.8,
  100915.9, 100865.9, 100788, 100677.2, 100538.2, 100384.4, 100261.3, 
    100230.3, 100225.3, 100260.7, 100385.8, 100515.9, 100580.4, 100658.6, 
    100780.1,
  100936.9, 100891.5, 100851.6, 100752.8, 100619.2, 100504.1, 100385.4, 
    100283, 100274.5, 100337.1, 100498.1, 100628.4, 100707.1, 100833.1, 
    100927.8,
  101039.3, 101161.2, 101298.1, 101403.7, 101462.8, 101450.4, 101393.5, 
    101316.3, 101167.3, 100650.2, 100489.2, 100534.1, 100189.1, 99579.97, 
    99258.83,
  101315.4, 101373.5, 101436.4, 101477.2, 101434, 101206, 101346.9, 101112.7, 
    100879, 100733.4, 100473.7, 100266.4, 100029.8, 98103.91, 98482.46,
  101474.4, 101507.7, 101516.4, 101529.5, 101332.6, 97951.36, 100976.9, 
    101158.3, 100849.6, 100589.5, 100273.2, 99994.98, 99706.49, 99521.41, 
    99397.93,
  101530.7, 101529.6, 101529.6, 101502.2, 101433.6, 101111.3, 97461.34, 
    100547.2, 100641.6, 100480.1, 100136.8, 99772.2, 99507.11, 99372.67, 
    99326.43,
  101534.2, 101520.8, 101513.9, 101460.5, 101402.8, 101268.4, 100948.3, 
    95079.91, 94224.22, 100255.7, 100137.1, 99727.17, 99455.81, 99303.81, 
    99353.57,
  101484, 101476.4, 101450.1, 101419.8, 101277, 101182.6, 101074.9, 100858.6, 
    100603.3, 100549.3, 100206, 99916.59, 99685.77, 99546.11, 99565.13,
  101427.5, 101428.3, 101426.3, 101358.5, 101256.1, 101120.2, 101015.5, 
    100989.8, 100818.7, 100553.7, 100329.8, 100169.1, 100012.7, 99940.36, 
    99944.05,
  101372.6, 101410.5, 101392.3, 101311.7, 101180.4, 101095.6, 101010.8, 
    100887.4, 100767.5, 100643.4, 100468.5, 100377.2, 100314.4, 100280.4, 
    100291.7,
  101380.1, 101434.6, 101384.3, 101305.8, 101211.8, 101112.7, 101026.8, 
    100984.6, 100876.8, 100724.7, 100621.9, 100570.4, 100544.6, 100539.4, 
    100550,
  101430.9, 101447, 101389.1, 101312.7, 101210.2, 101133.3, 101053.3, 
    100950.4, 100870.1, 100785.5, 100757.2, 100743.3, 100743.5, 100760.4, 
    100776.2,
  99768.73, 99802.19, 99884.43, 100012.5, 100192.3, 100400.1, 100683.6, 
    100971.3, 101239.6, 101132.4, 101368.4, 101706.9, 101548.1, 101027.5, 
    100710.9,
  99969.32, 99851.24, 99945.44, 100119.5, 100271.1, 100403.3, 100781.5, 
    101008.9, 101231.2, 101496, 101631.1, 101740.6, 101681.1, 99764.4, 
    100166.2,
  100420.5, 100211.5, 100193.1, 100341.8, 100312, 97413.94, 100824.4, 
    101245.1, 101377.5, 101555.8, 101663.5, 101720.4, 101655.8, 101516.3, 
    101260,
  100781.7, 100657.5, 100585.9, 100599.8, 100728.6, 100548, 97466.95, 
    101035.4, 101506, 101626.9, 101692.3, 101676.1, 101645.5, 101474.3, 
    101250.9,
  101062.2, 100989.3, 100945, 100930.3, 100996.2, 101137.2, 100950.6, 
    95520.34, 94966.63, 101391.3, 101691.2, 101658, 101624.3, 101431.5, 
    101299.6,
  101257.5, 101228.7, 101195.1, 101201.1, 101184.1, 101252, 101380, 101275.2, 
    101285.2, 101664.5, 101639.8, 101673.1, 101612, 101483.2, 101371.4,
  101397.9, 101406.2, 101400.3, 101391.5, 101415.7, 101425.8, 101461, 
    101624.4, 101672.1, 101613.7, 101644.5, 101663, 101603.3, 101521.8, 
    101449.9,
  101490.1, 101533.5, 101523, 101520.4, 101503.8, 101551.9, 101574.5, 
    101562.3, 101603.4, 101666.1, 101676.4, 101677.9, 101631.8, 101574.9, 
    101553,
  101583.3, 101619.1, 101609.2, 101612.2, 101612.7, 101629.9, 101660.5, 
    101724.5, 101730.2, 101700.5, 101694.9, 101710.8, 101658.6, 101619.4, 
    101602.7,
  101663.2, 101659.2, 101644.7, 101640.6, 101640.9, 101655.8, 101675.6, 
    101663.9, 101664.7, 101696.8, 101733.3, 101742.1, 101707.1, 101699.8, 
    101689.9,
  100729.6, 100635.7, 100559.2, 100518.2, 100510.6, 100465.3, 100536.8, 
    100724, 100899.6, 100745.8, 100990.8, 101438.4, 101522.8, 101350.6, 
    101298.1,
  100826.1, 100640.8, 100507.7, 100495.7, 100418.9, 100277.2, 100509.2, 
    100593.2, 100742.2, 100952, 101135, 101412.8, 101653.8, 100089, 100792.9,
  100926.7, 100701.4, 100489.5, 100438.1, 100289.1, 97168.02, 100321.4, 
    100665.3, 100739.7, 100888.3, 101089.7, 101378.8, 101655.6, 101831.6, 
    101955.9,
  101027.8, 100799.3, 100559.9, 100342.8, 100362.4, 100069.6, 96939.6, 
    100246.3, 100669.9, 100873.1, 101093.3, 101345.5, 101661.7, 101890.7, 
    101996,
  101148.8, 100934.5, 100691.7, 100450.5, 100293.9, 100353.5, 100130, 
    94962.39, 94430.73, 100593.4, 101136.8, 101350.2, 101670.7, 101866.5, 
    102052.9,
  101258.8, 101084.8, 100834.4, 100597, 100353.6, 100255.2, 100355.4, 
    100232.8, 100238.6, 100847, 101121.7, 101406, 101709.3, 101929.4, 102094.6,
  101363.1, 101222.4, 101023.9, 100786.9, 100563, 100398.3, 100339.8, 
    100547.8, 100756.4, 100904.5, 101175, 101492.4, 101763.2, 101982.8, 
    102127.9,
  101455.4, 101352.5, 101171.2, 100975.4, 100735.8, 100586.3, 100478.8, 
    100503.3, 100715.2, 101028.6, 101327.8, 101606.1, 101850.7, 102048.2, 
    102203.8,
  101523.9, 101468.8, 101348, 101198, 101008.4, 100856.5, 100784.4, 100884.8, 
    101054.8, 101258.6, 101504.8, 101744.2, 101941.4, 102114.4, 102245.4,
  101571.2, 101526.5, 101470.3, 101362.2, 101250.2, 101152.8, 101094.2, 
    101122.2, 101250.8, 101442, 101691.7, 101885.4, 102035.6, 102184.6, 
    102300.4,
  101191.1, 101077.6, 100924.2, 100802.1, 100704.6, 100625.3, 100678.9, 
    100829.9, 100966.6, 100757.4, 100920.7, 101257.3, 101216, 100982.1, 
    100976.9,
  101409.5, 101272.1, 101116.7, 100988.9, 100777, 100613.8, 100754.8, 
    100748.4, 100853.5, 100992.1, 101065.3, 101204.4, 101301.5, 99733.41, 
    100456.8,
  101563.3, 101464.9, 101308.9, 101203.2, 100881.5, 97565.78, 100716.9, 
    100885.7, 100870.7, 100936, 101002.6, 101121, 101252.6, 101359.7, 101505.4,
  101694.8, 101576.6, 101470.2, 101309, 101231.3, 100842.1, 97346.47, 
    100565.6, 100848.4, 100936.9, 100993.6, 101052.1, 101185.8, 101344, 
    101515.3,
  101764.1, 101689.9, 101570.6, 101445.8, 101294, 101251.9, 100921.9, 
    95262.53, 94615.13, 100676.2, 100972.9, 100990.9, 101106.5, 101241.7, 
    101477.2,
  101767.1, 101715.4, 101606.7, 101485.3, 101315.3, 101199.1, 101137.9, 
    100957.1, 100745.1, 101018.9, 100966.7, 100972.6, 101051.8, 101194.7, 
    101437.2,
  101722.7, 101698.7, 101632.8, 101493.7, 101336.3, 101178.5, 101034.4, 
    101026.2, 101016.8, 100920.4, 100913.2, 100943.9, 101002.8, 101151.8, 
    101396.1,
  101636.1, 101636, 101581.3, 101453.6, 101263.9, 101107.1, 100932.5, 
    100747.8, 100671.9, 100721.7, 100785.3, 100852.6, 100962.6, 101140.5, 
    101409.3,
  101530.3, 101578.1, 101561.5, 101436.8, 101261.5, 101060.3, 100834.3, 
    100682.3, 100599.7, 100561.8, 100613.1, 100734.8, 100910.8, 101150.8, 
    101443.2,
  101441.6, 101502.5, 101500.1, 101393.3, 101230.2, 101043.5, 100808, 
    100540.8, 100389.3, 100357.9, 100476.9, 100647.8, 100881.5, 101171.1, 
    101473.3,
  100062.1, 99795.45, 99658.91, 99739.14, 99866.6, 100061.9, 100279.7, 
    100523.7, 100737.3, 100635.9, 100880.6, 101278.4, 101264.4, 101024.6, 
    100979.6,
  100536.3, 100249.6, 100004.9, 99950.02, 99977.09, 100036.9, 100360.9, 
    100539.5, 100720.6, 100926.5, 101089.5, 101284.3, 101400.1, 99822.05, 
    100489.4,
  100974.2, 100699.2, 100468.7, 100299.4, 100075.6, 97139.49, 100399.6, 
    100736.8, 100867.6, 100995.1, 101130.7, 101281, 101417.7, 101485.9, 
    101538.1,
  101338.2, 101114.9, 100905.5, 100708.9, 100597.9, 100277.2, 97188.24, 
    100617.5, 101001.8, 101161.6, 101251.9, 101321.8, 101415.3, 101510.8, 
    101554.9,
  101585.1, 101454.6, 101296.3, 101111.9, 100968, 100932.6, 100604.9, 
    95318.4, 94891.87, 101111.6, 101393.8, 101389.2, 101443.3, 101458.6, 
    101547.2,
  101717.9, 101666, 101563.7, 101468, 101302.8, 101230.7, 101223.3, 101058.4, 
    101038, 101452.7, 101486.1, 101496, 101491, 101483.1, 101508.5,
  101771.3, 101750.4, 101736.4, 101691.5, 101622.4, 101545.9, 101496.6, 
    101604.2, 101640.7, 101564.6, 101567.5, 101591.9, 101565.9, 101541.9, 
    101489,
  101752, 101747.5, 101747.1, 101802.4, 101758.8, 101743, 101699.3, 101605.8, 
    101584.2, 101650.3, 101658.6, 101639.4, 101614.2, 101587.7, 101547.7,
  101662.9, 101690.9, 101726.1, 101803.9, 101840.9, 101830.5, 101820.2, 
    101851.4, 101821.9, 101741.9, 101684.9, 101660.2, 101629.8, 101593.1, 
    101539,
  101556.7, 101568.4, 101618.6, 101711.1, 101791.7, 101836, 101813.4, 
    101745.4, 101687, 101649.6, 101653.8, 101618, 101563.1, 101525.9, 101489.9,
  99569.21, 99431.12, 99570.66, 99815.08, 99968.28, 100002.9, 100107.6, 
    100288.7, 100516.3, 100463.4, 100785.3, 101251.7, 101326.2, 101151.8, 
    101143.4,
  99768.34, 99454.27, 99545.59, 99771.43, 99862.57, 99822.52, 100075.4, 
    100253, 100463.2, 100733.4, 100991.9, 101273, 101479.6, 99976.55, 100695.2,
  100073.6, 99699.89, 99633.35, 99786.44, 99731.19, 96725.53, 99982.36, 
    100355.4, 100566.2, 100742.9, 100992.3, 101251.1, 101493, 101638.8, 
    101751.4,
  100415.7, 100001.9, 99794.61, 99783.47, 99871.14, 99632.79, 96637.77, 
    100042.3, 100527.3, 100754.5, 100997.2, 101214.6, 101472.4, 101658.4, 
    101781.6,
  100739, 100375.3, 100076.2, 99933.37, 99878.87, 100005.7, 99831.9, 
    94830.52, 94461.4, 100537.2, 101011.8, 101188.1, 101436.7, 101604.6, 
    101778.4,
  100995.7, 100734, 100415.3, 100185.6, 99980.74, 99963.45, 100152.2, 
    100102.1, 100173.6, 100729.6, 100941.1, 101169.6, 101401.8, 101596, 
    101762.6,
  101204.5, 101023.8, 100776.1, 100526.9, 100297.6, 100142.3, 100184.7, 
    100434.5, 100637.4, 100740.2, 100935.3, 101170.4, 101390.8, 101590.1, 
    101749.4,
  101370.8, 101237.4, 101061.4, 100864.7, 100637.6, 100427.7, 100350.7, 
    100368.9, 100515.3, 100757.2, 100982.2, 101201.5, 101413.4, 101614.3, 
    101780.6,
  101490.4, 101399.8, 101281.6, 101167.8, 101002.8, 100822.9, 100679.8, 
    100716.5, 100809.7, 100928.1, 101094.3, 101301.1, 101493.5, 101680.6, 
    101835.2,
  101564.4, 101468.4, 101408.3, 101325.1, 101251, 101149.3, 101019.9, 
    100916.2, 100936.6, 101043.1, 101239.5, 101413.6, 101581.9, 101758.1, 
    101895.6,
  100882.2, 100569.7, 100520, 100668, 100861.4, 100937.5, 101021, 101001.1, 
    100838.6, 100517.3, 100795.1, 101235.8, 101291.8, 101052.3, 101008.3,
  100833.6, 100464.9, 100377.3, 100546.2, 100711.6, 100719.1, 100959.4, 
    100926.3, 100786.6, 100844.2, 101070.1, 101350, 101538.4, 99989.77, 
    100720.9,
  100875.8, 100472.3, 100327.9, 100490.1, 100538.8, 97448.47, 100762.8, 
    100979.7, 100924.8, 100904.2, 101143.8, 101403.6, 101663.7, 101801.4, 
    101906.1,
  100965.8, 100580, 100387.3, 100417.1, 100648.6, 100436.1, 97247.5, 
    100543.8, 100781.6, 100932.3, 101192.8, 101436.6, 101721.5, 101912.7, 
    102035.3,
  101092, 100755.5, 100516, 100454.6, 100540.7, 100752.7, 100516.8, 95188.45, 
    94675.66, 100751.8, 101226.1, 101455.3, 101743.9, 101922.5, 102098.7,
  101213, 100940.6, 100639.9, 100493.4, 100449.6, 100519.8, 100740, 100620.1, 
    100528.5, 100978.8, 101180.5, 101449.8, 101717.2, 101929, 102100,
  101328.1, 101106.2, 100831.2, 100599.7, 100446.7, 100455.8, 100535.9, 
    100807.4, 100967.9, 100987.1, 101139.6, 101397.9, 101652.9, 101871, 
    102041.6,
  101425.9, 101240.1, 100990, 100740.6, 100486.3, 100351.8, 100433.1, 
    100525.9, 100679.3, 100910.9, 101096.2, 101312, 101556.5, 101780.3, 
    101971.7,
  101488.2, 101364.3, 101161.8, 100934.9, 100674.2, 100409.1, 100318.6, 
    100510.6, 100711.3, 100869, 101033.1, 101232.8, 101449.8, 101664.8, 101855,
  101507.3, 101430.5, 101273.6, 101081.4, 100847.3, 100589.6, 100321.6, 
    100323.4, 100485.9, 100691.4, 100934.2, 101132.4, 101332.2, 101540.4, 
    101729.5,
  101951.6, 101806.6, 101631.8, 101548.9, 101550.3, 101558.9, 101534.5, 
    101546.6, 101440.5, 100939.4, 100821, 101087.8, 100967.6, 100613.5, 
    100442.3,
  101855.8, 101643.6, 101431.3, 101354.6, 101310.6, 101220.4, 101417.6, 
    101400.1, 101271.8, 101218.9, 101134.5, 101227.4, 101236.3, 99568.5, 
    100197.7,
  101746.5, 101497.2, 101267.5, 101185.4, 101081.3, 97862.98, 101134.6, 
    101380.7, 101309.5, 101214.9, 101210.2, 101314.7, 101416.2, 101459.7, 
    101432.6,
  101659.9, 101404.8, 101186.5, 101046.8, 101118.6, 100872, 97546.36, 
    100852.4, 101068.5, 101130.5, 101271.4, 101399, 101535.3, 101606.1, 101627,
  101596.9, 101385.9, 101128.9, 101029.9, 101021.2, 101159.2, 100897.9, 
    95333.2, 94736.14, 100896.3, 101336.6, 101473.7, 101634.4, 101675.6, 
    101783.5,
  101568.1, 101399.4, 101117, 100995.6, 100974.7, 101004.2, 101138.5, 
    100920.6, 100710, 101129.8, 101329.1, 101535.2, 101699.8, 101794.9, 
    101893.6,
  101566.3, 101447.4, 101176.7, 100994.4, 101002, 101020.5, 101030.4, 101082, 
    101071.4, 101116.9, 101342, 101570.9, 101751.4, 101877.8, 101992,
  101603.6, 101502.1, 101254.7, 101032.6, 100941.4, 100978.1, 101031, 
    100915.1, 100895.6, 101097.6, 101358.6, 101580.6, 101788.8, 101940.1, 
    102085.4,
  101644.5, 101587.5, 101402.7, 101180.4, 101014.3, 100964.6, 100984.5, 
    101013.4, 101030.6, 101156, 101367.4, 101592.5, 101799.4, 101961.7, 
    102105.1,
  101684.9, 101649.3, 101528.3, 101351.4, 101121.4, 100996.2, 100961.9, 
    100915.4, 100954.7, 101110.5, 101367.7, 101586.3, 101783.6, 101954.3, 
    102098.1,
  102276.5, 102341.9, 102326.4, 102289.6, 102240.3, 102118, 102027.3, 
    101942.6, 101814, 101286, 101149.3, 101156.9, 100907.2, 100569, 100484.4,
  102230, 102270.5, 102270.2, 102241, 102142.1, 101893.7, 102023.5, 101841.6, 
    101686.2, 101606.6, 101419.9, 101258.2, 101160.2, 99492.55, 100184.6,
  102174.7, 102192.4, 102179.3, 102160.7, 102011.8, 98591.86, 101760.1, 
    101944.3, 101768.3, 101598, 101431, 101303.1, 101292.7, 101365.4, 101411.1,
  102123, 102094.3, 102079.9, 102035.4, 102014.8, 101759.8, 98166.34, 
    101430.8, 101621, 101583.1, 101449.7, 101354.6, 101384.3, 101507.4, 
    101615.1,
  102032.2, 102001, 101965.7, 101937.6, 101888.8, 101891.5, 101646.5, 
    95933.95, 95124.55, 101376.7, 101497, 101413.1, 101458.9, 101576.1, 
    101765.7,
  101934.6, 101900, 101833.6, 101768.9, 101675.8, 101643.8, 101696.5, 
    101575.8, 101457.2, 101664.4, 101536.8, 101483, 101503.5, 101671.5, 
    101843.1,
  101850.1, 101788.8, 101682.1, 101573.7, 101482.7, 101454.2, 101452.5, 
    101601.9, 101666.8, 101574.3, 101556.1, 101498.7, 101526.8, 101713.1, 
    101896.5,
  101761.2, 101638.2, 101494.6, 101362.4, 101216.7, 101204.8, 101248.5, 
    101299.6, 101387.6, 101489.4, 101516.7, 101480.4, 101546.5, 101745.4, 
    101956.7,
  101652.4, 101509.2, 101366.5, 101227.7, 101058.7, 100998.9, 101050.5, 
    101200.4, 101337.7, 101390.2, 101436.9, 101463.7, 101544.5, 101757.2, 
    101971.1,
  101575.8, 101387, 101270.4, 101117.2, 100867, 100746.2, 100822.2, 100936.4, 
    101091.2, 101205.9, 101354.8, 101424.2, 101534.2, 101765.3, 101974.5,
  102345.6, 102452.4, 102473.4, 102481.4, 102450.4, 102387.9, 102300.5, 
    102163.2, 101958.1, 101424.7, 101280.8, 101348.3, 101092.4, 100646.4, 
    100436.6,
  102371.5, 102480.1, 102535.6, 102547.8, 102487.5, 102310.9, 102429.8, 
    102243.2, 102080, 101921.5, 101667.2, 101556.1, 101433.2, 99667.96, 
    100244.8,
  102333.3, 102455.9, 102536.4, 102578.7, 102453.3, 99071.81, 102358.7, 
    102513.8, 102306.1, 102117.2, 101877.2, 101713, 101654.1, 101601.8, 
    101514.1,
  102285.6, 102389.6, 102475.4, 102529.9, 102542.1, 102384.6, 98741.38, 
    102168.3, 102321, 102306.6, 102089.9, 101918.7, 101797.8, 101790.2, 
    101736.5,
  102335.6, 102352.5, 102394.4, 102450.1, 102489.6, 102551, 102402.2, 
    96570.4, 95820.41, 102180.1, 102296.8, 102092.6, 101945.6, 101892.9, 
    101913.2,
  102317.1, 102311.2, 102293.2, 102313.4, 102330.8, 102383.1, 102457.4, 
    102403.5, 102287.5, 102469.9, 102384.9, 102246.6, 102060.5, 102025, 
    102031.7,
  102202.7, 102177.9, 102152.4, 102151.5, 102169.7, 102208.7, 102256.3, 
    102397.4, 102445.8, 102429.1, 102415.4, 102337.9, 102162.6, 102100.7, 
    102125.9,
  102090.7, 102035.8, 101966.6, 101936.2, 101917.9, 101960.9, 102029.6, 
    102087.2, 102181.8, 102314, 102359.4, 102330.2, 102247.2, 102165.7, 
    102213.4,
  102015.3, 101918.2, 101810.7, 101715.3, 101678.4, 101694, 101773.6, 
    101914.8, 102054.9, 102146.3, 102239.1, 102285.7, 102262, 102206.7, 
    102248.2,
  101952.7, 101777.5, 101598.8, 101466, 101411.2, 101422.5, 101500.3, 
    101594.5, 101741, 101885.7, 102079.5, 102180.3, 102221.4, 102226.6, 102266 ;

 rlut =
  186.7222, 194.2757, 192.7097, 204.8557, 198.6682, 190.0629, 195.1854, 
    191.2768, 191.5528, 171.4344, 170.7977, 171.6754, 164.1939, 168.8092, 
    158.8546,
  188.569, 199.0868, 195.0602, 191.7088, 181.9433, 179.9996, 189.8094, 
    194.9452, 195.5129, 190.2661, 178.1034, 177.6634, 174.888, 163.1884, 
    156.7982,
  193.3486, 200.4762, 196.3385, 189.6511, 183.9561, 169.8442, 185.0716, 
    196.8983, 203.4032, 199.4102, 192.038, 180.4719, 175.3746, 171.045, 
    163.5138,
  190.5482, 197.5287, 194.6769, 197.7034, 193.525, 190.0928, 167.2314, 
    191.3926, 197.0063, 197.2567, 192.7287, 184.7601, 180.4041, 172.0914, 
    169.2234,
  192.428, 201.084, 203.5893, 202.3525, 199.8602, 197.9088, 196.4487, 
    164.582, 171.6045, 186.5409, 189.5247, 182.4898, 178.1878, 175.7353, 
    172.4164,
  198.1227, 199.3893, 200.0807, 206.8369, 208.3036, 210.6583, 201.5773, 
    197.7393, 198.9808, 189.6227, 179.2669, 175.1239, 174.4442, 166.9892, 
    170.521,
  205.4943, 208.1395, 198.7731, 194.4453, 196.5861, 208.0246, 196.0914, 
    193.8118, 195.6661, 187.9236, 179.3095, 173.8251, 169.6132, 169.3038, 
    172.2475,
  215.1657, 204.3699, 198.1151, 200.5763, 199.3142, 206.8559, 199.336, 
    195.6741, 191.0237, 177.6417, 178.0886, 169.8724, 167.5806, 163.5483, 
    169.0258,
  201.2531, 199.6181, 199.9539, 204.4133, 203.1487, 205.023, 201.4388, 
    196.647, 187.41, 188.539, 178.0096, 170.9474, 166.5488, 166.2778, 171.542,
  201.4429, 205.7095, 200.5584, 205.5298, 196.558, 200.9058, 194.6199, 
    198.8224, 189.6818, 182.9379, 179.0433, 176.0473, 166.2269, 167.8445, 
    167.78,
  184.7233, 195.8312, 191.2898, 205.2937, 203.5549, 190.8419, 176.6682, 
    166.258, 163.1609, 163.4114, 162.5, 155.1787, 151.9681, 154.7532, 158.0946,
  200.022, 193.3197, 195.9277, 202.2185, 196.451, 189.8699, 181.7442, 
    172.3282, 167.4415, 167.909, 159.9196, 163.2513, 155.8603, 157.4274, 
    158.1145,
  201.2159, 198.2912, 203.312, 197.6499, 201.1906, 170.627, 185.5983, 
    174.022, 172.6525, 171.4199, 167.3178, 159.9857, 163.6272, 163.937, 
    163.6401,
  210.726, 202.0393, 209.5648, 205.1411, 203.255, 204.7584, 169.032, 178.09, 
    178.5542, 173.3483, 167.4994, 164.3115, 165.7402, 162.9797, 164.9045,
  216.2454, 212.5307, 199.1647, 203.931, 206.988, 209.2002, 204.23, 171.1328, 
    164.2349, 172.6315, 170.6471, 170.0926, 167.533, 168.3033, 169.2719,
  211.3516, 209.5372, 202.0083, 203.5089, 190.5234, 198.7406, 199.4697, 
    201.1189, 187.692, 178.8015, 173.9836, 172.0318, 169.8255, 170.5081, 
    171.135,
  210.6067, 205.5921, 208.4576, 206.919, 199.6504, 192.5153, 196.7047, 
    194.6034, 196.2474, 190.4058, 185.8932, 175.952, 176.5656, 173.8887, 
    174.6303,
  215.4309, 210.3895, 201.1946, 202.4957, 200.5618, 202.9854, 198.5481, 
    196.2984, 189.4414, 189.1752, 184.6711, 179.7362, 179.278, 176.5906, 
    179.7525,
  213.7549, 212.1475, 206.0556, 204.1759, 199.4206, 199.6671, 200.9135, 
    194.9045, 189.8655, 197.6914, 188.2903, 178.6505, 178.0285, 178.926, 
    178.8849,
  217.2834, 210.082, 208.3664, 204.8511, 199.734, 195.168, 194.8864, 
    196.0617, 198.2664, 186.7502, 186.24, 180.73, 180.5617, 183.3732, 184.4637,
  189.6529, 196.1631, 195.0582, 202.9131, 196.1674, 183.4075, 183.5612, 
    189.7891, 190.1398, 176.9493, 178.3311, 183.3206, 180.3806, 178.702, 
    168.7405,
  192.0303, 204.6477, 202.7372, 196.7122, 183.9797, 177.4079, 173.6509, 
    186.49, 189.1751, 182.0827, 180.9524, 186.2009, 186.3264, 173.3558, 
    172.2489,
  193.5036, 198.8956, 205.4256, 199.5666, 182.3115, 167.3545, 177.3315, 
    179.7782, 181.0047, 179.0688, 186.0652, 184.5729, 182.8174, 182.6535, 
    182.8483,
  192.5618, 203.5035, 206.7883, 198.4347, 186.7669, 178.7205, 167.3269, 
    176.7122, 175.3115, 177.5633, 182.7944, 184.0048, 181.6175, 180.6633, 
    185.6208,
  191.9871, 202.7338, 205.5755, 203.6465, 197.3231, 190.5532, 175.9481, 
    170.1742, 176.0128, 177.5989, 180.6221, 181.9673, 178.3699, 181.3714, 
    184.5762,
  188.7365, 194.889, 202.9477, 205.0181, 200.4332, 189.939, 174.4878, 
    168.9975, 181.8043, 187.5904, 181.6445, 179.0583, 176.2176, 176.8677, 
    183.0909,
  191.852, 191.8294, 198.1012, 205.9717, 201.8825, 189.0352, 181.4689, 
    170.9267, 173.006, 182.1028, 183.6269, 173.4653, 174.6311, 178.6035, 
    187.5443,
  196.8191, 200.2873, 198.2163, 200.2031, 196.425, 190.5728, 177.0167, 
    177.9075, 171.4627, 172.7506, 178.0359, 173.8857, 173.3276, 178.2831, 
    184.1537,
  195.8696, 199.3202, 201.0211, 196.7089, 192.886, 182.4494, 183.0689, 
    180.098, 173.5388, 172.5543, 172.9055, 166.4972, 168.6031, 171.1896, 
    175.5643,
  193.8489, 198.014, 201.3718, 199.5975, 191.0545, 187.8248, 180.3439, 
    182.5317, 180.0779, 176.3932, 171.9, 164.298, 160.4768, 166.2088, 171.9181,
  178.21, 189.6674, 193.4578, 190.1511, 186.7158, 178.1618, 184.3498, 
    191.1536, 191.4254, 177.2012, 178.1212, 179.4348, 173.3155, 174.8007, 
    162.3042,
  185.5631, 196.5712, 201.0572, 200.3667, 181.3515, 179.0037, 189.1129, 
    192.302, 193.1843, 189.1101, 182.0591, 185.0364, 187.4249, 169.6404, 
    164.0162,
  193.2972, 204.9, 212.5006, 201.6777, 187.9576, 172.5871, 191.0068, 
    191.9142, 192.4579, 188.8043, 188.8459, 186.595, 185.9883, 189.9301, 
    180.7668,
  206.7185, 212.9506, 214.8423, 210.1007, 199.5133, 192.1976, 180.6362, 
    195.2039, 194.4796, 187.8724, 187.6271, 186.9634, 186.7268, 187.7769, 
    186.713,
  208.4145, 216.6991, 208.2877, 211.8591, 211.0705, 204.2927, 199.106, 
    182.32, 181.3149, 186.5441, 188.1573, 187.9528, 188.7668, 190.919, 
    190.6857,
  212.7972, 214.187, 209.9382, 204.509, 210.2691, 208.455, 205.8527, 
    204.3872, 204.2013, 203.823, 191.3185, 189.576, 191.0996, 192.2801, 
    192.5249,
  213.585, 209.2566, 210.0099, 211.2687, 210.9932, 203.2493, 203.4936, 
    192.1752, 189.966, 187.8583, 199.4037, 193.064, 193.5826, 194.106, 
    195.1924,
  214.3189, 208.6735, 208.989, 206.1106, 210.7313, 205.0695, 202.3956, 
    182.2422, 181.2571, 187.5807, 199.9992, 195.6059, 195.5839, 196.2396, 
    196.5947,
  212.9668, 213.5696, 207.2896, 199.1766, 198.5658, 201.7014, 201.9837, 
    185.3644, 190.3381, 184.8422, 203.6237, 197.211, 197.2937, 195.6932, 
    196.8702,
  214.7295, 211.0367, 199.7714, 189.9033, 194.6543, 200.6186, 199.0499, 
    192.5262, 192.3605, 204.7978, 201.9819, 198.5388, 197.8454, 195.8987, 
    197.4881,
  183.8251, 184.5343, 185.6517, 182.2028, 185.2313, 185.8823, 192.1637, 
    189.0338, 186.1033, 176.9804, 173.1203, 176.1617, 168.8056, 168.8001, 
    159.3069,
  183.2041, 187.2525, 183.7998, 178.0948, 183.782, 193.5636, 193.6224, 
    191.0232, 188.1986, 184.6943, 177.2116, 182.8356, 184.6137, 165.2372, 
    157.7709,
  179.8858, 191.1798, 188.2583, 189.8261, 196.5146, 188.3292, 191.7613, 
    188.5183, 187.4629, 186.8656, 186.8172, 184.3006, 182.9824, 184.021, 
    173.2089,
  185.2762, 190.5429, 194.0299, 195.6798, 205.7625, 204.2292, 183.4012, 
    188.7171, 187.6075, 186.5285, 185.3798, 182.3423, 182.3359, 183.1618, 
    180.7804,
  192.4728, 189.3161, 192.6808, 195.5852, 205.5567, 207.6953, 208.2173, 
    179.2886, 176.6615, 182.9436, 184.477, 182.7782, 184.4384, 185.9309, 
    188.8512,
  190.6599, 193.4204, 201.6325, 207.1298, 206.4667, 206.5201, 209.3751, 
    213.3174, 201.2946, 198.39, 185.79, 184.5507, 185.1239, 188.2639, 190.2789,
  197.3387, 200.5914, 208.646, 210.0501, 206.5598, 201.4171, 208.5033, 
    208.4221, 194.0596, 182.8011, 192.4233, 185.4347, 187.6548, 190.7095, 
    191.9543,
  200.726, 203.6435, 212.7498, 208.8255, 210.5148, 202.947, 208.6291, 
    196.7516, 181.062, 180.3868, 190.2836, 187.4228, 190.1459, 192.426, 
    193.6748,
  196.3068, 210.7412, 215.6006, 210.2402, 207.7432, 201.9706, 206.0927, 
    194.6734, 180.1466, 179.0952, 193.2456, 190.0428, 192.7361, 193.9766, 
    194.1563,
  202.5395, 218.167, 212.6049, 210.0103, 204.8958, 208.571, 209.6059, 
    200.3778, 187.3386, 200.6711, 193.5994, 191.4284, 194.4434, 193.7843, 
    194.4785,
  174.8817, 179.179, 184.5674, 201.6878, 191.7131, 191.0393, 190.244, 
    185.993, 186.3615, 174.7225, 169.1858, 175.9149, 169.1531, 169.7152, 
    160.6719,
  186.1062, 182.6237, 190.2538, 198.4079, 191.7784, 192.8273, 189.9063, 
    189.7682, 188.7966, 185.2857, 174.2711, 184.7956, 186.6108, 166.05, 
    160.6142,
  189.5703, 185.3344, 199.7036, 203.1022, 190.5415, 187.7236, 192.1384, 
    190.1754, 189.0283, 188.0257, 189.0256, 188.5426, 186.096, 183.9939, 
    171.4182,
  193.7685, 196.7892, 201.871, 198.9587, 195.3203, 203.2772, 183.6691, 
    188.7187, 188.3186, 188.2539, 188.1181, 188.5257, 189.469, 187.2016, 
    180.6187,
  194.1763, 200.2747, 202.2044, 199.0602, 190.0157, 199.1076, 210.1085, 
    177.4644, 171.3307, 180.1859, 186.8474, 190.0231, 191.1842, 190.6071, 
    192.1458,
  190.4062, 205.7716, 202.8627, 194.291, 195.3471, 204.1333, 205.1304, 
    215.9129, 201.5482, 195.912, 187.2534, 191.6686, 192.7213, 192.9477, 
    190.2757,
  206.3174, 197.7324, 198.4649, 193.6992, 201.7589, 207.0463, 207.3078, 
    195.9633, 197.5324, 201.4737, 198.8005, 193.6389, 193.7423, 194.7128, 
    193.3201,
  209.7284, 198.1629, 196.9394, 194.0919, 200.5297, 211.1079, 209.5643, 
    212.9722, 191.923, 199.0704, 196.3184, 194.4492, 195.3504, 195.1813, 
    196.5733,
  206.5737, 199.5023, 194.3421, 196.5642, 201.8413, 209.2943, 213.4621, 
    211.9773, 185.4158, 193.9403, 195.4361, 194.786, 195.5128, 195.6523, 
    195.4365,
  201.3146, 197.7581, 194.9565, 197.9901, 199.4324, 209.8519, 208.6528, 
    208.4963, 197.4283, 196.1465, 194.9733, 194.8639, 195.4819, 196.2189, 
    195.1501,
  201.7088, 202.6943, 202.6483, 215.489, 195.8579, 189.8722, 192.7155, 
    189.0985, 181.0121, 165.3829, 162.0921, 158.5541, 158.9541, 160.5423, 
    156.686,
  197.6376, 202.911, 211.3022, 208.5738, 194.6554, 190.103, 193.2992, 
    189.5504, 181.3312, 173.0132, 163.4924, 165.4354, 167.8232, 159.7534, 
    158.4227,
  191.8219, 197.687, 197.4951, 191.5084, 202.3217, 186.0701, 193.2486, 
    190.1486, 182.838, 174.7247, 166.8676, 164.1086, 166.2188, 167.7323, 
    163.6642,
  182.0518, 198.2945, 197.1869, 191.0258, 195.9575, 202.5276, 184.3849, 
    185.6718, 183.7984, 173.6453, 166.6696, 166.9883, 167.4416, 176.4176, 
    172.5551,
  173.4191, 191.4585, 202.5588, 213.7998, 204.6155, 195.2953, 203.0484, 
    177.9341, 166.6492, 169.2371, 165.8742, 170.9322, 176.7742, 182.6738, 
    189.6656,
  169.7825, 178.2912, 192.2476, 213.0121, 210.2611, 197.866, 197.747, 
    201.2321, 189.1348, 179.0758, 173.6582, 176.9107, 181.7083, 185.5632, 
    192.8004,
  187.0834, 175.131, 182.3041, 209.444, 212.1446, 216.1978, 197.5943, 
    197.4542, 193.0072, 198.2351, 185.4937, 183.5379, 184.1958, 188.7384, 
    192.6646,
  193.9768, 184.5837, 183.5229, 202.2667, 213.6675, 215.1996, 208.9732, 
    202.4516, 195.9422, 188.9591, 187.6601, 184.8729, 186.9081, 189.4638, 
    194.0591,
  192.7118, 189.9535, 189.1092, 195.5499, 210.8157, 214.0344, 212.6297, 
    196.36, 201.9595, 194.3313, 191.6078, 190.0383, 188.0192, 187.7234, 
    191.2823,
  199.4868, 191.9271, 188.1425, 192.9143, 209.2627, 211.5701, 213.4476, 
    211.7982, 205.6748, 198.4872, 194.69, 191.7188, 192.1942, 190.0605, 
    191.2882,
  166.076, 184.9417, 188.6756, 206.9754, 193.3423, 182.0441, 180.8298, 
    177.7563, 178.0731, 170.7606, 169.3409, 172.1099, 167.9636, 170.9668, 
    166.2264,
  157.3606, 170.229, 190.9027, 194.6674, 190.2905, 181.2477, 184.5648, 
    174.7771, 176.5346, 176.937, 171.9126, 176.5008, 178.1026, 165.2915, 
    161.0782,
  161.5049, 166.1855, 180.222, 192.276, 199.2684, 180.388, 184.6894, 
    174.3119, 175.9337, 176.2188, 180.1569, 180.4059, 180.2237, 178.2646, 
    170.4398,
  161.9946, 159.9536, 177.5155, 188.1383, 195.1164, 199.9819, 171.9908, 
    174.0584, 174.1649, 172.5758, 176.6618, 179.9837, 179.0603, 181.2479, 
    177.5644,
  157.6088, 158.2175, 172.2316, 205.6689, 197.1091, 191.7651, 193.7255, 
    170.5627, 168.0935, 169.9499, 175.5994, 183.4982, 184.2977, 184.7478, 
    184.4049,
  164.2867, 159.3405, 173.7874, 211.0625, 193.44, 193.9403, 186.731, 
    175.4471, 171.7916, 174.3836, 178.7774, 186.2961, 188.4492, 186.1325, 
    188.307,
  196.1517, 167.1112, 177.6304, 209.1248, 214.1675, 192.6037, 187.5827, 
    175.9857, 174.5636, 176.0134, 181.7739, 183.5895, 186.7948, 185.6145, 
    182.9503,
  214.2456, 196.2383, 185.8192, 208.3351, 211.5965, 213.7927, 186.642, 
    177.4766, 169.4874, 171.4282, 180.9191, 183.4135, 186.4716, 183.5255, 
    183.9451,
  198.9928, 208.7713, 203.7015, 212.4762, 212.0638, 214.5126, 209.9119, 
    179.7587, 168.8001, 174.8251, 178.7294, 179.1827, 182.1116, 182.7077, 
    177.1404,
  182.6478, 194.3455, 208.2619, 208.5341, 207.5265, 212.2813, 207.3, 
    184.5354, 170.9606, 172.0572, 177.7166, 178.1848, 176.4654, 175.5421, 
    176.2809,
  173.2276, 161.3723, 163.0906, 186.7729, 183.1713, 179.2021, 183.9904, 
    181.3428, 182.7025, 168.8303, 168.565, 174.4652, 169.1282, 172.1268, 
    163.6497,
  182.9226, 165.5657, 167.0094, 182.0475, 180.4076, 176.1895, 183.5619, 
    186.3634, 184.8493, 184.1581, 173.3033, 185.637, 187.863, 164.2473, 
    160.6998,
  188.0504, 167.3659, 167.2691, 179.2697, 192.1143, 170.6736, 183.8467, 
    185.1459, 187.4739, 188.4836, 189.0277, 189.6186, 189.2434, 185.0499, 
    173.403,
  187.9035, 185.7293, 168.2432, 174.7856, 195.6918, 190.5326, 173.6239, 
    182.5948, 187.02, 187.3914, 187.8515, 188.5096, 186.4774, 184.2864, 
    176.346,
  190.1111, 183.7605, 176.854, 183.707, 187.0469, 189.8557, 193.5996, 
    175.6428, 173.6584, 180.2408, 186.7348, 186.6415, 181.9238, 182.8264, 
    183.3579,
  188.1999, 188.1763, 186.0405, 190.7193, 190.3402, 195.6658, 188.3818, 
    197.1132, 191.8534, 190.3849, 186.5618, 186.987, 183.0535, 186.3058, 
    185.0368,
  192.4191, 187.8146, 188.3535, 196.3148, 204.3493, 183.4546, 192.8885, 
    188.9318, 196.0884, 200.6286, 192.3218, 188.0825, 186.3844, 186.454, 
    183.5217,
  196.5435, 187.4131, 191.7962, 201.4636, 208.1957, 193.8644, 184.3074, 
    189.3703, 193.5583, 196.6341, 190.9362, 189.6597, 188.7623, 188.3534, 
    183.0527,
  205.3039, 196.6926, 200.926, 209.3853, 209.3591, 197.0709, 190.7253, 
    190.9836, 194.0313, 190.3247, 189.8556, 188.5905, 189.8682, 187.0935, 
    181.0382,
  204.9118, 204.2001, 207.2708, 210.8457, 210.3475, 207.9162, 195.489, 
    188.1134, 192.5571, 190.9594, 191.0692, 187.8173, 189.2667, 185.3636, 
    178.4503,
  188.934, 200.821, 187.4682, 188.3904, 180.5279, 177.7551, 183.7192, 
    183.4645, 185.1236, 175.8962, 175.3545, 175.9209, 172.4807, 171.9983, 
    165.5004,
  185.6548, 188.0735, 188.186, 186.9599, 178.8437, 175.9348, 185.044, 
    186.1467, 186.9168, 185.7652, 177.1852, 183.4397, 184.6355, 170.3863, 
    170.2388,
  189.6214, 182.3493, 186.935, 179.7603, 193.1126, 173.6465, 180.8497, 
    187.037, 185.3866, 186.3601, 185.8911, 183.614, 183.4504, 182.4693, 
    174.1892,
  204.325, 188.732, 180.4052, 182.8837, 188.1198, 198.7395, 175.5086, 
    180.3053, 186.7526, 184.7734, 184.1062, 183.3428, 183.4613, 184.7524, 
    179.8795,
  207.0408, 199.9482, 194.4389, 188.7801, 190.7837, 190.9457, 197.147, 
    173.9213, 170.3479, 176.6638, 182.4624, 184.2108, 182.2973, 181.6445, 
    180.6794,
  216.063, 208.2541, 208.0411, 205.847, 186.679, 193.1036, 191.6099, 
    199.6998, 195.131, 188.4659, 179.993, 186.4297, 184.4947, 182.995, 
    183.3602,
  209.2601, 211.9514, 213.3434, 214.3397, 211.5965, 200.2002, 193.0322, 
    192.9276, 195.49, 197.8728, 188.7867, 187.9631, 184.3412, 184.2043, 
    183.6076,
  219.4777, 217.632, 217.629, 211.1228, 210.0728, 205.7138, 206.6063, 
    191.665, 194.28, 195.976, 192.7955, 188.0094, 185.2325, 184.7254, 184.886,
  221.87, 217.9739, 214.9557, 208.5705, 211.2607, 201.9245, 206.2405, 
    209.702, 195.4254, 194.3584, 193.1107, 188.1396, 186.2349, 184.2061, 
    184.8286,
  193.0493, 217.2848, 213.7271, 211.1086, 205.2314, 198.696, 196.8908, 
    203.8765, 209.0978, 200.2059, 197.3472, 189.5519, 186.5868, 185.7033, 
    181.9763,
  191.539, 208.6926, 191.2934, 199.0369, 189.3, 182.183, 184.4153, 180.8613, 
    178.3468, 174.7244, 174.1073, 174.4007, 170.3137, 172.5731, 168.9137,
  191.4263, 200.5252, 204.6564, 207.5146, 182.6718, 179.0712, 188.1112, 
    183.3826, 180.7789, 177.5035, 172.105, 171.9558, 174.4845, 169.558, 
    167.9124,
  193.5044, 192.5537, 195.9114, 197.5862, 197.2098, 177.3335, 185.3286, 
    182.1664, 175.4053, 174.2233, 173.2455, 172.927, 172.3201, 171.3065, 
    166.4761,
  192.0758, 187.5826, 186.6785, 192.3, 198.9267, 200.576, 177.7638, 178.8467, 
    176.5012, 172.1426, 173.5802, 175.1517, 170.4685, 169.0404, 164.9067,
  194.0689, 193.2643, 186.9946, 187.5069, 191.2813, 198.9488, 198.717, 
    176.8536, 176.7901, 176.5642, 173.4284, 177.785, 175.0312, 176.6739, 
    168.1625,
  211.1549, 197.4732, 191.3837, 187.108, 187.3987, 191.5348, 198.3495, 
    197.0457, 184.6314, 176.1112, 174.074, 180.471, 182.4063, 182.3427, 
    176.337,
  217.2793, 215.8339, 203.0276, 210.2057, 211.3779, 196.0707, 199.542, 
    199.4352, 188.9895, 184.4576, 183.0769, 176.8983, 177.9009, 181.0144, 
    176.3956,
  200.0313, 198.7886, 201.3724, 203.3671, 208.6075, 212.3199, 211.5008, 
    201.5463, 189.8024, 187.4907, 183.9646, 179.164, 178.1839, 181.7654, 
    179.4436,
  173.2891, 174.6065, 181.6508, 193.154, 200.5069, 211.9413, 211.7699, 
    209.5006, 199.6327, 182.8431, 186.8041, 184.3533, 182.9286, 180.0809, 
    182.4582,
  173.8513, 172.1703, 180.5692, 185.2931, 190.5521, 205.7306, 211.4211, 
    211.3106, 202.129, 187.1164, 189.0537, 184.7108, 185.2221, 182.9504, 
    184.4198,
  190.2779, 206.9267, 191.9235, 198.3234, 189.8681, 179.9279, 184.1884, 
    184.4073, 183.0509, 176.7965, 171.0303, 168.1196, 164.9808, 164.3602, 
    162.6673,
  203.1012, 191.0945, 197.7007, 198.6754, 185.8931, 177.5896, 181.0383, 
    185.2747, 188.1756, 183.0195, 173.3847, 166.9397, 166.1354, 163.3392, 
    158.3423,
  193.5648, 189.0574, 194.1327, 196.0754, 193.8328, 180.3467, 180.3545, 
    183.4409, 184.9285, 184.7803, 180.0012, 173.9763, 167.3802, 166.1703, 
    162.1734,
  196.099, 189.8256, 188.8339, 193.5038, 201.4222, 196.3123, 172.3728, 
    179.2793, 184.1731, 184.6138, 181.6742, 175.1756, 171.5051, 166.0675, 
    157.3137,
  197.7281, 196.0939, 192.6023, 195.0307, 195.5399, 204.0678, 195.2647, 
    174.4324, 178.3878, 182.2867, 184.9639, 180.8918, 173.4573, 170.7905, 
    164.5887,
  179.1168, 177.528, 194.418, 199.8675, 202.9964, 203.3924, 196.2744, 
    202.1637, 190.0349, 187.472, 183.6829, 186.4576, 181.1109, 177.8504, 
    169.9155,
  177.3992, 178.0928, 173.5652, 186.4276, 203.5207, 213.2989, 208.1127, 
    194.1243, 205.2435, 193.1502, 192.5308, 189.2345, 186.8977, 181.6392, 
    175.2123,
  173.2111, 177.4987, 182.2862, 186.6988, 198.5153, 209.9547, 214.8831, 
    204.888, 192.6885, 194.421, 192.9108, 190.9265, 187.7727, 182.1708, 
    179.3132,
  195.7237, 203.7303, 197.272, 195.8132, 195.0307, 197.0305, 214.6418, 
    206.6343, 201.8808, 191.7219, 193.4454, 191.7779, 188.814, 186.5283, 
    184.8577,
  197.7352, 209.2023, 203.3156, 207.5623, 200.9688, 186.7694, 207.5675, 
    212.5427, 206.7309, 197.7148, 195.0233, 193.4537, 190.8465, 190.7657, 
    187.9041,
  189.1118, 202.6919, 191.2866, 196.9572, 192.7179, 185.1651, 191.1037, 
    191.1155, 186.4114, 176.1277, 168.8121, 165.7881, 161.5901, 167.7887, 
    167.8637,
  207.9876, 208.238, 200.9083, 201.2402, 188.4911, 183.5559, 189.7091, 
    191.1924, 188.0278, 183.9507, 171.5903, 171.1809, 164.9429, 163.6056, 
    169.2648,
  195.2335, 200.6788, 206.5734, 208.3878, 194.6127, 183.441, 188.8175, 
    190.1809, 188.7024, 187.4935, 180.8628, 173.1349, 165.51, 166.6562, 
    167.1033,
  202.9236, 198.7798, 198.6815, 214.0885, 207.8145, 193.9601, 185.9942, 
    184.9595, 189.5082, 188.6744, 186.0479, 179.3066, 170.8574, 166.3533, 
    163.9173,
  198.3771, 196.8521, 214.4223, 205.1841, 210.991, 215.3413, 201.7614, 
    179.8303, 178.5747, 187.5612, 189.6694, 184.1885, 175.774, 166.4607, 
    167.7899,
  203.1481, 195.9865, 216.1398, 215.1722, 213.4606, 213.3652, 205.2635, 
    210.0112, 194.218, 188.8678, 190.1746, 188.9659, 179.8946, 173.1909, 
    167.7636,
  214.9069, 216.7763, 202.1035, 200.5341, 211.5348, 215.7548, 207.3631, 
    205.3095, 202.3671, 198.5458, 193.8876, 190.8078, 187.234, 181.9306, 
    170.2581,
  206.0312, 215.9694, 203.3045, 207.0577, 216.7719, 216.5951, 211.1518, 
    204.3382, 205.6378, 194.9829, 192.2779, 191.1115, 189.7112, 184.6546, 
    180.631,
  212.9707, 210.7908, 221.9066, 219.5805, 218.6066, 217.9916, 214.9345, 
    212.5769, 204.237, 194.5401, 192.9726, 192.7673, 191.4551, 188.9988, 
    188.8947,
  190.3286, 199.8, 203.3082, 211.4465, 212.346, 217.4321, 214.3662, 214.9485, 
    211.8521, 196.6359, 195.3888, 194.658, 192.8974, 191.8474, 190.0191,
  165.2533, 178.4529, 177.2005, 181.4824, 181.7382, 182.6407, 186.3513, 
    189.8624, 190.8417, 187.8826, 186.1933, 184.4137, 179.7713, 173.6317, 
    166.946,
  175.509, 176.0062, 181.4209, 181.4068, 181.4524, 181.4847, 187.7519, 
    193.1375, 192.3437, 189.6066, 186.5142, 185.7233, 181.1935, 174.7439, 
    164.9356,
  187.9284, 190.0651, 188.3955, 189.7057, 185.6272, 179.5002, 191.8866, 
    192.9891, 192.0276, 191.0057, 190.7862, 186.4778, 180.1253, 174.0546, 
    164.8372,
  192.0261, 200.6218, 195.1545, 196.8809, 203.0953, 193.537, 189.1175, 
    193.379, 195.1037, 190.6804, 192.5102, 188.4762, 182.5804, 173.1547, 
    164.2885,
  206.6716, 204.9406, 204.091, 210.9838, 210.9729, 202.9218, 202.0164, 
    192.525, 189.4348, 189.1668, 190.9154, 187.522, 182.063, 176.5793, 
    168.8369,
  213.782, 207.8969, 212.7731, 214.654, 213.713, 216.1317, 213.8341, 
    210.5972, 203.0097, 189.767, 188.4258, 187.3327, 183.4897, 177.148, 
    167.7473,
  216.0424, 214.6789, 212.421, 215.6198, 216.2265, 214.869, 215.0583, 
    213.1655, 211.4482, 188.7411, 188.312, 187.4764, 182.8526, 176.1702, 
    173.6766,
  219.6542, 215.0727, 213.6823, 212.2219, 217.0063, 217.6018, 215.9996, 
    216.858, 216.4377, 198.8608, 188.7064, 188.224, 183.8566, 177.6899, 
    174.8143,
  216.0741, 219.6943, 219.4004, 218.9009, 214.6531, 218.4779, 218.6609, 
    217.8375, 217.5972, 209.9975, 198.9702, 196.4576, 188.4718, 176.656, 
    179.6082,
  219.1145, 218.3588, 219.5549, 221.2919, 218.4946, 218.156, 219.0985, 
    218.3952, 215.0217, 204.7028, 198.7357, 196.4281, 190.3377, 175.849, 
    172.676,
  169.2758, 165.2463, 162.6013, 163.7714, 165.0899, 169.1855, 173.6555, 
    183.9417, 189.3531, 187.2271, 186.282, 184.5567, 177.6854, 177.3265, 
    170.1574,
  174.0717, 167.1447, 165.6304, 164.1332, 164.2652, 165.5533, 172.9399, 
    183.6012, 190.4371, 193.1544, 189.9911, 187.0189, 180.6231, 176.817, 
    174.9484,
  180.8024, 169.2946, 164.2207, 164.7915, 166.3336, 163.7399, 171.4155, 
    181.7446, 190.1767, 192.5861, 188.0089, 184.1148, 179.9477, 176.2458, 
    177.2515,
  180.7212, 171.6034, 162.4245, 158.3489, 169.0285, 170.977, 167.5759, 
    175.1742, 184.8063, 187.1844, 184.9518, 181.3437, 172.6017, 172.3905, 
    178.8779,
  176.3234, 166.6619, 163.6437, 163.7082, 162.2913, 175.6711, 179.9435, 
    177.3138, 182.9214, 184.5158, 184.5133, 182.0537, 172.879, 169.7491, 
    180.0712,
  171.5766, 167.5782, 163.2173, 168.4171, 168.6897, 174.0273, 179.982, 
    194.973, 192.7306, 185.3004, 185.8874, 183.1784, 173.0467, 163.035, 
    172.3277,
  175.5389, 170.4462, 172.7724, 174.7863, 174.2304, 184.7669, 182.8113, 
    192.9625, 200.8519, 187.1605, 187.0488, 185.5979, 176.1782, 164.6527, 
    169.9735,
  184.2969, 180.6272, 181.4081, 185.0746, 184.0093, 188.5266, 197.3014, 
    202.1012, 208.9711, 208.9369, 200.5926, 193.5981, 182.9159, 164.9072, 
    166.6589,
  196.3732, 191.4736, 192.3886, 193.2507, 197.9694, 200.6913, 206.6003, 
    208.4176, 213.4786, 211.4764, 201.1225, 193.8455, 188.5177, 172.2649, 
    168.471,
  206.0662, 206.4526, 206.6734, 206.3634, 206.8135, 211.7848, 214.6548, 
    214.1902, 214.0784, 201.4858, 200.1131, 191.9208, 191.8499, 183.8163, 
    175.184,
  186.2418, 186.2841, 183.6533, 182.6848, 177.4935, 178.5286, 186.3084, 
    189.4813, 188.7428, 187.8136, 185.9529, 189.6053, 179.688, 172.3625, 
    157.814,
  196.2221, 196.816, 195.3049, 181.4514, 171.1182, 172.009, 181.5841, 
    187.355, 190.3468, 187.5449, 184.6568, 187.8333, 188.6687, 174.3643, 
    161.7683,
  202.1295, 195.6837, 179.8632, 172.5015, 174.6628, 165.9041, 173.3671, 
    176.2865, 186.3928, 185.028, 183.8764, 183.8559, 187.4793, 183.0415, 
    163.4868,
  194.6346, 187.0524, 173.8048, 170.1725, 171.652, 174.7365, 165.1047, 
    169.6508, 183.3181, 181.9808, 183.7155, 183.9138, 183.5579, 186.8924, 
    167.364,
  196.2689, 191.8822, 181.0731, 170.6799, 166.5229, 172.5234, 180.8582, 
    166.11, 179.7921, 176.493, 182.9961, 183.8551, 183.8965, 192.7905, 
    177.7161,
  201.0526, 192.847, 185.8321, 175.8838, 172.4556, 170.0161, 172.4615, 
    179.8232, 172.7159, 168.438, 179.1637, 183.6331, 184.3034, 192.5748, 
    182.206,
  211.3275, 200.0469, 184.5618, 171.5271, 168.4639, 168.4126, 169.4649, 
    177.5485, 174.387, 169.0289, 176.8016, 183.1974, 189.6668, 190.3488, 
    187.6776,
  203.4536, 195.3213, 182.404, 175.1599, 168.6779, 161.2367, 162.1138, 
    164.7289, 166.0221, 177.8747, 182.0099, 184.7293, 189.1575, 187.8921, 
    186.9809,
  194.2136, 191.8772, 185.8458, 171.7708, 167.0375, 161.8872, 163.3751, 
    164.9324, 168.2198, 179.0144, 188.7, 198.9432, 191.8923, 192.7713, 
    185.7705,
  193.3021, 184.7134, 179.7683, 170.3887, 167.1714, 159.6148, 165.2173, 
    166.7761, 173.555, 178.8953, 193.8543, 201.718, 199.077, 188.4205, 182.887,
  194.8262, 200.4311, 195.0319, 195.8924, 190.0945, 185.5752, 186.8303, 
    187.9595, 186.145, 181.1482, 181.1306, 180.4779, 181.0514, 170.5244, 
    166.1931,
  211.9855, 212.4895, 206.3439, 199.3666, 181.5332, 177.8288, 184.8847, 
    184.2905, 185.6841, 182.3524, 182.1743, 182.4543, 177.306, 177.3772, 
    167.542,
  212.8447, 213.2739, 200.5416, 199.4122, 190.2845, 168.1677, 177.3422, 
    178.2285, 180.4905, 181.6264, 183.1907, 183.668, 178.3122, 176.7221, 
    168.6892,
  212.2586, 203.4768, 188.5104, 183.0762, 189.4041, 188.3934, 170.5299, 
    166.6823, 175.9231, 179.1574, 181.3671, 182.6392, 179.6454, 176.489, 
    176.9953,
  204.0921, 192.088, 184.3533, 184.4099, 179.7171, 174.1815, 182.4747, 
    170.8789, 171.4262, 172.4639, 178.7619, 188.6771, 182.2159, 175.8059, 
    176.1615,
  192.868, 185.6618, 180.6396, 182.4153, 177.4951, 176.0919, 174.7869, 
    175.5098, 170.4958, 168.4687, 176.8392, 186.8061, 185.9138, 176.6085, 
    173.9448,
  187.9469, 182.9293, 189.7625, 182.4494, 179.0619, 178.9165, 177.9902, 
    172.704, 170.5662, 176.6267, 175.0379, 183.5256, 188.4028, 175.1901, 
    174.3503,
  186.7109, 184.7137, 176.9147, 178.0262, 179.0817, 173.8292, 175.9043, 
    173.5556, 173.6007, 168.0305, 170.0645, 177.0175, 191.1975, 184.6884, 
    171.8362,
  185.7611, 182.8329, 178.6387, 179.9008, 180.6966, 179.199, 176.5831, 
    175.6449, 171.9264, 168.3266, 169.0205, 171.7658, 187.2198, 197.5059, 
    174.3906,
  206.1961, 201.9148, 196.7274, 193.1594, 187.7871, 186.4101, 178.1886, 
    170.3633, 170.6319, 163.3091, 171.2311, 168.624, 178.6277, 197.2972, 
    173.9022,
  198.4365, 202.33, 197.3578, 196.6746, 190.6805, 184.2547, 190.6456, 
    187.7199, 186.4632, 182.2782, 184.6362, 184.0091, 173.506, 169.2287, 
    159.429,
  208.5546, 201.2317, 202.8913, 199.7446, 180.8575, 178.9517, 182.6068, 
    185.2363, 181.6768, 186.3224, 185.7745, 187.9847, 183.61, 164.275, 
    157.1149,
  204.0539, 197.5654, 196.9797, 198.3163, 196.074, 180.299, 178.021, 
    171.7178, 172.6866, 179.7681, 188.0078, 188.421, 185.7224, 181.0636, 
    169.165,
  196.9866, 198.0177, 196.3371, 194.5579, 194.9428, 189.3194, 180.8293, 
    169.1816, 173.1808, 176.8346, 185.056, 189.9918, 185.6719, 182.272, 
    175.9344,
  198.0096, 200.6001, 193.9093, 193.9494, 187.8861, 183.6682, 178.1486, 
    172.6183, 182.5368, 173.905, 180.1117, 190.7641, 184.595, 184.2305, 
    181.5503,
  197.1755, 193.4578, 193.0074, 185.2733, 185.91, 182.7886, 172.7478, 
    175.0358, 177.5299, 173.6591, 175.8212, 187.5528, 184.7809, 184.169, 
    183.0905,
  214.7843, 196.9034, 196.5821, 187.4521, 178.35, 177.3399, 175.3113, 
    179.7416, 179.805, 182.0367, 176.4297, 183.7932, 185.6361, 183.8808, 
    183.1911,
  191.6417, 184.0259, 182.0909, 176.5012, 172.7036, 176.6303, 181.3334, 
    186.3817, 193.1479, 186.8362, 178.1542, 182.8472, 185.5318, 182.0379, 
    180.9657,
  178.7415, 172.9741, 171.5943, 171.2801, 184.2493, 193.7505, 197.2864, 
    196.4104, 193.8369, 192.1252, 183.849, 179.2492, 186.3297, 182.757, 
    179.8451,
  175.7146, 178.2124, 189.5334, 199.4802, 206.5596, 206.6257, 204.4745, 
    200.8259, 190.8041, 189.206, 192.2515, 181.153, 184.6692, 188.1195, 
    179.6614,
  198.3133, 202.3608, 192.853, 197.0658, 193.6001, 188.8903, 187.6415, 
    188.9239, 186.8085, 170.7703, 166.9621, 168.8718, 162.7319, 162.7355, 
    155.4132,
  199.9964, 201.9128, 211.3546, 202.4641, 189.1576, 186.6713, 185.414, 
    187.2579, 189.8794, 183.3739, 173.1267, 178.877, 176.9809, 159.8787, 
    156.1708,
  194.9319, 197.8029, 202.7699, 208.2709, 197.2042, 187.6537, 183.5554, 
    176.7893, 185.6271, 188.4052, 185.6494, 182.4368, 179.3593, 175.2784, 
    162.7216,
  195.051, 194.8905, 199.6693, 195.8272, 205.8271, 192.2855, 179.9698, 
    182.3951, 188.7271, 189.9846, 186.8913, 184.0161, 180.9351, 175.839, 
    167.5706,
  193.4557, 196.4745, 195.5321, 189.2719, 194.4339, 190.4945, 191.0637, 
    184.0028, 188.941, 190.9426, 188.6937, 185.9256, 182.0762, 178.2221, 
    168.841,
  192.2419, 195.1391, 188.7382, 196.3601, 194.5855, 194.0226, 191.3609, 
    200.6403, 196.4115, 195.0711, 189.119, 188.2584, 184.0555, 179.6807, 
    171.2893,
  213.6053, 216.6031, 201.7092, 189.5748, 189.4432, 194.5253, 204.1782, 
    206.5475, 204.8182, 201.0106, 193.6968, 190.0038, 186.6519, 181.4342, 
    176.4589,
  220.7885, 211.7127, 190.6715, 184.2857, 187.3717, 196.774, 207.9901, 
    211.061, 206.8722, 200.0683, 193.6272, 191.7737, 189.7828, 185.3368, 
    177.5756,
  213.5569, 201.3064, 184.4688, 181.5368, 187.1048, 201.7882, 207.8099, 
    205.0501, 195.293, 193.3549, 193.2062, 192.5366, 192.5255, 189.3771, 
    179.4742,
  202.9296, 185.6923, 180.0671, 180.4313, 191.4523, 196.5375, 205.3776, 
    192.9335, 189.7696, 186.5182, 197.0189, 192.6759, 192.2541, 190.5428, 
    186.8102,
  189.4944, 197.8191, 192.874, 197.9619, 197.2111, 193.9381, 193.8143, 
    196.4439, 193.6008, 191.4528, 183.5755, 177.5059, 166.4829, 164.3737, 
    160.0684,
  202.0676, 202.2384, 205.4062, 203.5286, 194.3508, 193.8628, 194.9048, 
    198.1333, 195.7691, 197.541, 185.1947, 179.9506, 171.5597, 162.2416, 
    160.6941,
  194.0029, 195.8513, 192.6258, 194.4584, 200.1541, 192.2019, 193.9623, 
    192.1482, 189.1429, 189.6903, 187.7087, 182.6432, 174.6563, 163.1245, 
    159.8253,
  189.4022, 199.6018, 194.6466, 188.2378, 196.894, 193.9406, 188.7021, 
    189.1441, 189.9941, 184.7584, 183.68, 181.3032, 177.9266, 165.6406, 
    159.9864,
  196.4259, 199.7608, 196.2785, 187.0576, 193.0667, 184.8748, 187.8812, 
    188.3107, 192.6352, 184.4912, 181.8309, 181.0989, 178.6995, 163.827, 
    157.4989,
  212.087, 207.5476, 203.3911, 198.8126, 190.4983, 185.7838, 182.2111, 
    189.6783, 187.7343, 182.1647, 179.8853, 183.5388, 182.1395, 167.7111, 
    159.2271,
  216.8755, 214.4136, 210.9103, 200.9534, 189.8396, 184.5159, 186.511, 
    183.7677, 184.9241, 181.7896, 183.2433, 185.2811, 187.864, 175.5894, 
    162.3388,
  220.9754, 219.2921, 215.0511, 205.4892, 198.0127, 188.4801, 190.0009, 
    191.7361, 186.2218, 178.8327, 183.1956, 188.1859, 189.4162, 176.0858, 
    163.216,
  219.5797, 220.0316, 219.4546, 209.0383, 200.9991, 197.4437, 188.0664, 
    180.178, 175.6636, 176.4205, 184.0927, 189.9131, 192.2658, 184.9361, 
    163.044,
  222.7669, 216.103, 211.3195, 208.8976, 193.2335, 189.5139, 182.3237, 
    178.9765, 174.3038, 169.4682, 185.4081, 192.1393, 193.6432, 185.2891, 
    169.0737,
  153.3472, 162.5296, 164.9339, 170.3727, 173.1503, 170.8525, 170.516, 
    176.2973, 171.9738, 173.389, 173.8581, 176.4021, 168.9418, 165.4267, 
    160.2303,
  178.1378, 180.2607, 177.6008, 174.9805, 169.8706, 170.9018, 176.8314, 
    176.363, 177.059, 179.2044, 174.8219, 177.962, 168.7903, 165.2242, 
    159.1773,
  197.7071, 182.8584, 182.8479, 184.0473, 181.3797, 175.7322, 180.3107, 
    173.8244, 177.3938, 181.6133, 181.3444, 178.5832, 172.8096, 168.2126, 
    156.4176,
  191.4079, 183.7307, 186.3373, 196.3289, 196.8625, 195.2593, 179.9218, 
    184.3219, 180.3711, 176.1037, 184.1617, 180.4128, 171.4518, 166.3307, 
    155.315,
  193.9382, 200.3034, 207.1947, 203.6073, 203.5979, 196.033, 189.696, 
    182.198, 185.3183, 183.909, 181.3298, 178.1342, 172.097, 166.4096, 
    155.6296,
  206.5, 210.3633, 213.9089, 210.4296, 202.6017, 197.1974, 186.4321, 
    183.8294, 184.7466, 180.5215, 180.4179, 175.1759, 169.5288, 161.9444, 
    156.2621,
  207.5664, 212.5146, 210.1103, 199.6134, 189.1614, 191.4791, 185.9259, 
    185.1052, 183.4617, 183.0018, 175.7289, 170.1607, 165.5104, 160.9487, 
    157.0114,
  203.5136, 201.3331, 201.9566, 196.0707, 189.4582, 184.9046, 185.5128, 
    188.1687, 184.8209, 180.8178, 178.4627, 164.7238, 160.6022, 161.3341, 
    159.1743,
  201.5272, 193.7462, 190.299, 189.7858, 187.5457, 181.7655, 187.0465, 
    190.2728, 192.9836, 185.9024, 172.0347, 165.2719, 160.1821, 164.1456, 
    161.1334,
  185.2352, 184.3079, 179.3137, 186.6869, 184.5291, 188.7864, 191.4946, 
    189.9297, 191.7534, 179.4854, 174.2086, 165.3855, 164.9781, 167.0766, 
    161.816,
  193.9835, 195.4347, 193.9062, 193.0161, 191.3153, 191.4431, 191.1877, 
    190.057, 186.2222, 178.5727, 171.8582, 166.5643, 164.4466, 162.5044, 
    157.7741,
  211.1569, 211.9404, 213.9922, 203.1856, 191.1732, 192.7339, 196.1349, 
    190.9007, 184.4232, 173.1083, 163.8551, 163.8621, 163.6621, 161.2274, 
    155.0986,
  209.1981, 208.8561, 204.6883, 201.4523, 205.3879, 194.4271, 199.7494, 
    178.7084, 164.9818, 160.9671, 157.3644, 158.0455, 163.071, 163.533, 
    158.9816,
  204.6537, 200.3432, 200.6742, 197.8432, 203.5007, 206.9757, 188.8759, 
    173.3499, 155.1075, 150.8471, 151.2596, 154.9707, 163.5273, 165.1442, 
    163.5807,
  204.004, 205.6955, 199.6323, 204.5704, 198.5276, 192.5081, 184.6078, 
    172.3479, 162.1083, 150.6903, 148.1582, 159.2293, 169.892, 170.054, 
    163.2526,
  200.8267, 201.5223, 198.4015, 197.4085, 190.0678, 175.315, 166.8175, 
    153.8752, 153.3762, 155.2252, 157.5341, 175.231, 176.0594, 170.5038, 
    163.328,
  198.4407, 194.0272, 184.7698, 185.1655, 178.8489, 164.5555, 161.5624, 
    158.0942, 155.3404, 158.2511, 174.4962, 186.7164, 180.2653, 168.0059, 
    168.2823,
  190.8552, 176.5267, 176.1805, 167.9453, 168.393, 161.6864, 161.6671, 
    160.513, 167.3493, 176.8013, 186.577, 192.3339, 178.7278, 171.7121, 
    170.0065,
  181.7217, 172.0506, 170.6438, 157.8166, 163.8315, 160.6148, 159.0227, 
    164.9082, 175.2626, 183.2996, 188.8611, 190.3459, 186.4523, 177.4098, 
    169.6212,
  181.1813, 173.4784, 162.2457, 161.1062, 160.7365, 161.6879, 163.0975, 
    165.1094, 176.998, 179.414, 190.2444, 194.8649, 190.6905, 180.7194, 
    172.2895,
  189.1165, 199.1396, 198.1536, 196.8206, 191.2343, 191.877, 194.2181, 
    190.7916, 188.9005, 183.9791, 174.0448, 160.3396, 152.2369, 147.4534, 
    160.6581,
  188.8595, 200.1219, 207.6391, 204.7547, 190.9577, 197.1172, 199.2335, 
    193.7983, 191.6195, 184.0676, 171.5411, 162.0963, 151.741, 150.2903, 
    173.3407,
  176.9414, 184.774, 191.2454, 194.2811, 198.2547, 190.4045, 204.0444, 
    196.2632, 190.3715, 184.3643, 172.4596, 160.479, 152.6097, 164.5542, 
    183.6097,
  175.6193, 177.9324, 180.5417, 183.2904, 187.1977, 196.0927, 189.2478, 
    195.5163, 193.932, 185.6738, 171.5308, 163.637, 157.0104, 167.2382, 
    186.9925,
  170.2421, 169.8405, 170.1984, 174.1335, 179.0401, 178.3079, 184.7817, 
    180.0565, 187.3179, 178.4003, 168.5792, 163.3335, 165.2236, 177.4098, 
    185.827,
  173.4674, 170.3157, 171.0112, 168.1058, 168.6876, 165.5007, 171.7928, 
    174.1299, 173.177, 170.8677, 168.1661, 166.5713, 164.4486, 183.0667, 
    184.2491,
  174.3835, 172.8481, 170.7845, 173.4449, 173.9176, 171.645, 166.3259, 
    161.0625, 165.3654, 164.931, 167.783, 160.8358, 170.0369, 177.9919, 
    188.9279,
  179.8237, 180.9603, 184.6557, 186.8017, 184.3945, 184.7178, 173.8145, 
    168.8472, 164.1461, 165.686, 161.6862, 163.49, 171.5238, 177.5186, 
    184.1923,
  196.8211, 207.9463, 215.2351, 207.9642, 200.3037, 189.1441, 184.5355, 
    177.6167, 170.9522, 168.6292, 164.3853, 161.5715, 170.6037, 181.3272, 
    179.1474,
  213.9892, 219.8231, 213.9325, 203.8914, 191.2803, 185.9542, 181.4257, 
    176.5075, 174.2416, 169.7009, 165.6408, 161.8992, 171.9443, 182.2398, 
    180.3065,
  173.0043, 171.7373, 180.0117, 193.9452, 191.0222, 191.271, 194.7402, 
    189.5405, 186.5872, 177.1851, 176.1414, 166.2379, 158.1705, 151.8894, 
    163.7258,
  171.9753, 171.8735, 174.9962, 186.883, 189.8127, 197.3239, 198.9882, 
    192.3161, 189.8513, 184.768, 179.719, 171.5167, 161.4599, 151.8815, 
    166.6584,
  175.3174, 172.3201, 168.1729, 179.2893, 190.8561, 187.8643, 204.2561, 
    196.269, 192.2754, 188.1845, 185.5211, 175.1786, 166.985, 160.9124, 
    177.5961,
  176.8101, 172.4795, 166.7232, 168.0827, 179.6427, 197.4194, 186.2313, 
    198.3932, 196.4805, 191.6503, 184.8075, 180.1965, 170.1374, 165.5132, 
    182.9863,
  176.8221, 167.4477, 164.5184, 162.0576, 162.8466, 177.9813, 196.6335, 
    183.1945, 188.1461, 193.9529, 191.4148, 186.3446, 179.5371, 170.4291, 
    186.6782,
  191.5152, 171.8565, 165.1173, 162.8769, 164.3685, 167.2734, 169.5338, 
    189.297, 187.6538, 185.0505, 184.2298, 187.5463, 183.7334, 178.4741, 
    187.7953,
  209.1904, 189.2918, 168.4385, 160.198, 159.0061, 159.9008, 163.4924, 
    167.9121, 173.2945, 182.1081, 181.3336, 184.9075, 180.0045, 179.5552, 
    188.1044,
  223.4055, 210.0673, 187.9349, 172.2579, 165.1919, 162.4435, 163.843, 
    161.8414, 166.3418, 170.1346, 171.0543, 176.5931, 179.0768, 182.072, 
    187.9223,
  218.3782, 217.4454, 208.5655, 194.7637, 187.9887, 185.0271, 176.655, 
    175.8318, 168.238, 168.4006, 167.1225, 165.9649, 176.4486, 178.8705, 
    184.8378,
  213.0721, 214.5636, 204.4108, 202.9416, 196.6358, 193.7866, 190.3804, 
    189.3169, 182.5971, 174.866, 167.6769, 160.908, 172.3004, 174.9701, 
    184.6366,
  174.226, 173.7092, 175.3793, 187.8489, 186.7557, 190.4792, 193.5173, 
    186.2728, 183.4426, 174.4716, 170.4035, 171.2718, 165.827, 165.6843, 
    161.3136,
  174.3027, 180.8568, 185.5477, 191.7577, 186.5282, 195.6215, 195.2847, 
    188.1021, 185.7478, 181.5081, 174.1823, 179.3985, 176.1113, 162.2484, 
    159.8541,
  182.9073, 182.2676, 198.9533, 203.5592, 198.0123, 188.122, 197.3589, 
    190.1315, 186.9606, 184.0933, 183.463, 178.6331, 177.4741, 174.5299, 
    168.5569,
  173.2727, 180.2356, 191.7766, 195.0783, 217.364, 209.0488, 187.7279, 
    192.4384, 189.7396, 184.7529, 182.5898, 181.0487, 180.4701, 178.5933, 
    176.0029,
  174.3616, 174.981, 183.975, 190.6678, 198.2263, 218.0876, 216.7689, 
    185.3404, 182.7288, 188.6602, 187.767, 186.193, 180.4914, 180.7072, 
    184.1138,
  171.1583, 170.7266, 177.8987, 187.1908, 190.536, 201.0586, 215.8463, 
    218.0311, 200.3532, 193.1721, 191.5662, 191.5871, 184.3368, 183.1961, 
    183.7815,
  177.0586, 165.4442, 170.0357, 176.9415, 186.8708, 193.5122, 204.6136, 
    210.7657, 213.4549, 202.8059, 196.2174, 191.0216, 186.0342, 186.0749, 
    185.2253,
  186.9747, 172.6884, 167.8805, 168.2531, 178.7767, 184.8073, 190.7353, 
    198.327, 199.1413, 201.6906, 196.0451, 191.5428, 190.038, 186.7048, 
    184.6086,
  193.7421, 181.5769, 174.5547, 170.4774, 172.0788, 176.0258, 180.7731, 
    183.8956, 189.6388, 200.2272, 192.223, 191.6749, 191.4616, 187.3901, 
    183.7181,
  198.8093, 199.1425, 189.3396, 177.7165, 173.972, 173.1108, 176.6228, 
    180.585, 183.5295, 188.7572, 193.2247, 191.2735, 192.2253, 190.0414, 
    186.3558,
  191.4523, 194.877, 188.9674, 188.8836, 186.9893, 187.7108, 191.8572, 
    182.987, 183.3859, 172.4389, 168.858, 171.173, 166.7355, 168.9818, 
    165.3349,
  200.4228, 197.008, 196.7599, 192.8029, 186.7012, 190.5902, 189.0764, 
    184.3944, 182.3049, 180.5838, 174.6865, 179.7727, 180.1466, 164.9603, 
    162.2336,
  211.6138, 204.1566, 205.0653, 199.2075, 196.9643, 181.0085, 187.3661, 
    183.8012, 182.8223, 182.4568, 184.4734, 180.247, 178.4912, 178.1351, 
    169.1747,
  205.2451, 201.1271, 206.0682, 212.6165, 214.3631, 203.6098, 178.3907, 
    183.0455, 183.1804, 182.6989, 182.0114, 180.3459, 179.0313, 178.6443, 
    176.5701,
  190.6794, 195.5198, 203.6477, 208.2529, 215.0573, 214.3768, 212.0152, 
    178.653, 173.2293, 179.5543, 184.2051, 183.6625, 181.1855, 182.1426, 
    182.9749,
  188.7524, 188.026, 199.8544, 201.8757, 214.9886, 211.9271, 215.0909, 
    211.9131, 197.8357, 189.7394, 186.2969, 188.4028, 183.8386, 182.696, 
    181.3596,
  179.5586, 183.3569, 197.1217, 204.3035, 211.6056, 208.6309, 209.0157, 
    214.9004, 211.7189, 200.6723, 194.2259, 189.7124, 186.3906, 184.5111, 
    182.1139,
  179.7699, 182.4229, 197.9197, 211.2712, 212.9184, 212.8874, 205.2758, 
    201.1329, 200.8494, 200.8281, 193.0845, 189.5054, 188.4359, 184.8657, 
    182.0146,
  172.2781, 180.0896, 196.5966, 210.1201, 206.4706, 204.8093, 211.0178, 
    208.5628, 203.2354, 199.9059, 193.5956, 191.1036, 190.0223, 185.9972, 
    182.0577,
  172.7432, 180.9424, 195.1625, 205.847, 196.9971, 205.0667, 200.0922, 
    197.488, 205.2673, 197.5632, 199.2826, 193.4229, 191.5241, 188.4516, 
    185.6316,
  183.6155, 186.883, 178.7236, 179.7959, 184.1502, 184.3273, 187.4774, 
    181.9222, 184.4205, 175.6584, 174.1519, 178.798, 175.7397, 174.7343, 
    171.6342,
  189.4834, 186.0762, 183.2206, 183.6286, 184.4469, 183.0422, 183.8428, 
    181.3985, 180.887, 184.5557, 178.9971, 184.1733, 186.1787, 172.496, 
    169.2006,
  200.5318, 193.1449, 191.9442, 195.5059, 196.7336, 174.9945, 181.4867, 
    177.9786, 178.0687, 183.3763, 185.753, 183.9774, 184.7134, 183.3227, 
    173.896,
  201.7761, 194.4471, 192.7186, 210.5842, 214.1496, 199.495, 171.3894, 
    176.0189, 176.7251, 181.4928, 182.951, 183.0216, 183.3402, 183.1775, 
    178.4046,
  193.3799, 188.6629, 199.8605, 212.2552, 218.7214, 206.5946, 194.2186, 
    173.2717, 167.5683, 177.2692, 184.0219, 185.1105, 182.4613, 185.0729, 
    183.6841,
  194.3347, 196.7087, 193.5658, 213.9323, 219.6339, 208.7191, 194.9735, 
    194.4725, 192.3898, 189.5458, 184.2537, 187.9522, 185.3064, 184.7746, 
    182.8128,
  203.8227, 212.8628, 213.3336, 210.2157, 209.5909, 205.7026, 205.4434, 
    205.8891, 207.2284, 200.0319, 192.9757, 189.3607, 186.847, 185.8918, 
    185.3273,
  215.6507, 215.4161, 218.2705, 217.9305, 207.7403, 195.4014, 202.7187, 
    207.7191, 209.8561, 197.497, 191.8386, 189.9294, 189.0816, 185.6151, 
    184.0702,
  215.5389, 219.2113, 217.6764, 214.8607, 210.4617, 201.0638, 202.6569, 
    212.0387, 208.5573, 195.2643, 192.2273, 192.2111, 191.6046, 187.7214, 
    185.9819,
  214.351, 216.5083, 215.0208, 212.5471, 209.419, 204.7521, 200.6383, 
    201.3004, 200.2381, 191.7247, 196.9601, 194.6843, 192.9724, 190.856, 
    187.9057,
  181.7213, 195.8928, 193.1602, 194.5111, 188.1861, 185.1388, 188.748, 
    185.7639, 186.8969, 177.8025, 174.481, 174.8196, 171.4453, 173.725, 
    174.3334,
  184.2675, 201.5151, 203.5131, 194.6415, 184.9451, 182.3143, 185.9649, 
    183.7809, 183.1386, 181.4378, 174.905, 174.0084, 175.9677, 173.0198, 
    174.09,
  189.0346, 204.7656, 210.7811, 200.2444, 197.8706, 174.0996, 185.3045, 
    182.3377, 178.4605, 176.3711, 175.3629, 172.7123, 174.3217, 177.5799, 
    178.3447,
  188.9248, 202.2532, 215.7323, 211.9905, 212.0578, 201.0593, 173.1058, 
    182.1985, 179.6736, 174.2623, 171.2354, 169.8906, 172.5474, 176.1421, 
    179.618,
  183.7342, 194.2949, 211.3244, 211.1665, 214.4812, 208.505, 205.6532, 
    176.1261, 178.106, 177.3061, 173.1408, 171.8656, 173.9899, 177.7859, 
    180.4816,
  177.5148, 193.8829, 206.3459, 207.157, 213.1353, 209.5508, 205.7912, 
    200.7652, 184.891, 184.7812, 175.576, 175.7761, 173.4363, 175.4045, 
    178.705,
  176.6763, 185.5393, 189.023, 204.1786, 206.5079, 204.7169, 206.7396, 
    201.0054, 198.9392, 192.5531, 182.2859, 178.2471, 175.2876, 175.6396, 
    177.6632,
  172.7525, 190.1222, 198.2178, 199.5094, 199.5536, 196.4691, 199.084, 
    208.2099, 205.7448, 194.0135, 188.2792, 183.6326, 181.7716, 178.3152, 
    177.0345,
  172.4729, 185.8739, 205.8303, 208.3937, 198.1143, 190.0565, 197.4044, 
    204.8541, 208.8704, 198.084, 195.3475, 190.8644, 185.6201, 181.4451, 
    180.4616,
  178.6779, 188.0746, 206.7685, 211.9832, 206.5609, 188.8045, 196.005, 
    202.2576, 200.4702, 196.1644, 199.2428, 195.3363, 190.7352, 186.2399, 
    184.2978,
  193.6615, 198.046, 191.3411, 193.7809, 188.0198, 184.74, 187.4393, 
    186.8427, 187.475, 177.315, 174.6763, 177.4551, 176.6796, 177.3021, 
    172.4327,
  204.8925, 202.5065, 201.1731, 193.8773, 185.2501, 181.8757, 185.4863, 
    186.558, 184.9431, 184.8285, 178.7294, 183.0846, 183.7694, 173.3228, 
    168.6955,
  205.0101, 202.185, 203.0231, 196.5565, 192.4316, 173.7433, 182.5883, 
    181.1636, 182.1831, 182.8658, 183.7023, 184.2014, 183.47, 180.6591, 
    175.3649,
  200.6576, 200.3941, 198.207, 192.1689, 185.2926, 175.9664, 173.0143, 
    176.6536, 180.5058, 181.7962, 183.4835, 184.5518, 183.7963, 184.1476, 
    181.5623,
  197.0143, 194.1781, 190.5018, 184.6711, 178.6877, 169.2953, 171.1375, 
    172.9538, 177.8391, 181.9554, 184.4601, 188.9794, 187.095, 188.3465, 
    185.7906,
  196.3148, 192.0714, 187.8259, 182.62, 179.017, 180.5146, 177.7933, 
    179.3923, 184.4324, 186.9946, 187.3797, 192.1851, 191.6176, 188.1638, 
    185.5548,
  202.933, 196.7691, 192.3923, 184.5956, 179.6826, 179.3493, 180.4668, 
    180.5308, 185.0113, 185.9227, 189.9478, 192.9423, 192.6573, 187.5946, 
    184.2321,
  208.7392, 197.175, 192.9355, 189.9849, 187.7627, 184.3719, 184.3187, 
    184.1891, 186.8693, 185.7943, 187.1693, 190.1848, 190.8249, 188.1092, 
    190.444,
  213.3862, 209.6021, 215.9852, 192.5348, 191.3121, 190.4923, 190.2818, 
    189.8109, 186.6438, 185.2873, 185.0495, 184.6613, 179.2652, 185.2687, 
    184.0035,
  206.2672, 209.3208, 211.471, 197.9399, 195.0805, 193.9385, 192.9729, 
    195.4935, 187.392, 190.7573, 187.3557, 183.9469, 180.8974, 179.1785, 
    178.3268,
  189.7838, 192.4921, 184.0575, 189.058, 184.1556, 181.7685, 184.4979, 
    187.2234, 188.6491, 192.1171, 191.5202, 190.4724, 180.867, 178.4074, 
    174.4711,
  199.7157, 197.9028, 194.1885, 187.7502, 178.2681, 178.5197, 181.3391, 
    184.5654, 187.1655, 190.0006, 184.2255, 180.3544, 177.4215, 173.8859, 
    172.7713,
  199.1261, 203.4028, 202.4711, 193.5291, 188.8161, 171.2806, 177.5103, 
    177.2629, 181.325, 177.6391, 172.5046, 174.3574, 175.4242, 174.5335, 
    175.7656,
  195.0494, 200.2965, 194.1044, 196.0038, 193.4257, 186.0077, 170.7738, 
    176.29, 175.9639, 171.0777, 170.7299, 172.2955, 170.7483, 176.6958, 
    176.2381,
  192.1901, 189.9599, 186.5612, 188.5769, 194.5298, 189.2774, 190.5614, 
    175.122, 166.6527, 166.4098, 166.8294, 167.9368, 168.8698, 176.7465, 
    181.8684,
  191.4094, 184.9544, 182.7028, 183.4969, 186.6073, 189.7722, 188.2233, 
    183.0965, 176.2375, 171.6458, 166.0624, 167.9887, 170.3061, 175.4221, 
    185.8347,
  177.6781, 183.1834, 185.2181, 185.0586, 188.0355, 190.5729, 192.111, 
    182.171, 177.2255, 172.0433, 168.6484, 168.9583, 172.802, 179.7758, 
    188.2496,
  178.5495, 177.8623, 180.0632, 189.6208, 192.7448, 198.0733, 189.8246, 
    183.3239, 179.9694, 176.6782, 168.088, 168.2183, 174.3936, 184.8563, 
    189.0553,
  180.4996, 177.3455, 182.4762, 189.3645, 194.5961, 196.5651, 192.6966, 
    186.4068, 181.4233, 172.6552, 169.5232, 170.128, 173.9651, 185.3082, 
    190.5813,
  190.3352, 191.0338, 194.2709, 192.6325, 195.1435, 196.3162, 193.3251, 
    184.4517, 179.9957, 173.8134, 173.0538, 172.4844, 178.2707, 186.4831, 
    192.058,
  184.0011, 190.1458, 185.5066, 192.0797, 185.5515, 187.5529, 189.1314, 
    188.4082, 190.2542, 184.8807, 186.7612, 190.2979, 187.5332, 184.2947, 
    179.891,
  194.5829, 195.151, 194.4393, 192.16, 184.3461, 187.5128, 189.7784, 
    189.1936, 188.2545, 188.0604, 184.5069, 188.639, 189.7836, 180.0554, 
    178.34,
  194.8192, 194.3008, 198.621, 196.1927, 191.698, 187.7841, 190.0387, 
    187.1541, 185.3528, 184.7411, 188.746, 189.419, 190.3109, 191.3601, 
    184.6953,
  186.8414, 187.134, 189.1374, 191.4109, 189.866, 191.3793, 187.6022, 
    185.5372, 179.111, 180.588, 182.1594, 185.416, 187.9262, 189.2903, 
    189.3836,
  180.1524, 186.292, 181.8226, 183.4068, 186.8555, 187.8641, 192.5138, 
    178.5129, 172.8776, 176.2587, 180.3398, 184.4538, 187.9694, 190.5872, 
    190.7588,
  186.945, 185.9155, 186.4963, 180.184, 184.2965, 188.1466, 182.1671, 
    175.9793, 175.0591, 178.1543, 178.5147, 184.4614, 189.6466, 190.3737, 
    190.7692,
  197.1106, 184.2548, 181.775, 176.8723, 182.6404, 185.286, 179.543, 
    167.5047, 170.8187, 175.5381, 180.9978, 186.4739, 190.2431, 189.767, 
    190.1047,
  193.3516, 190.8282, 180.6833, 182.2506, 182.0594, 178.241, 171.458, 
    165.6688, 168.5853, 176.9563, 179.6596, 186.0811, 189.9815, 189.8238, 
    190.1864,
  186.4531, 195.1767, 182.679, 185.3985, 182.8993, 178.2176, 169.7039, 
    164.8071, 164.5462, 169.3711, 171.4186, 184.396, 189.2061, 189.5989, 
    190.6674,
  190.7117, 191.5193, 187.8814, 185.4689, 183.1621, 182.3788, 170.2858, 
    163.6579, 161.4396, 162.7649, 172.3977, 179.3494, 187.8633, 190.2466, 
    191.9059,
  183.81, 192.2092, 179.4305, 176.2797, 170.0126, 170.5082, 177.2402, 
    183.5609, 189.8173, 189.5783, 187.6196, 186.4028, 182.6086, 178.6495, 
    173.3182,
  199.5395, 198.8638, 195.3278, 180.8607, 169.2387, 170.3681, 176.4356, 
    185.1772, 190.7498, 191.7815, 189.5671, 190.4663, 190.5412, 176.3493, 
    173.5064,
  216.1432, 202.662, 202.8724, 187.8491, 178.7561, 169.4633, 177.2818, 
    185.9002, 190.8141, 190.9365, 191.8882, 189.213, 188.8994, 189.5668, 
    181.4555,
  205.5648, 198.5452, 196.2006, 192.9586, 180.4125, 176.6387, 174.3305, 
    182.3283, 189.9989, 190.4409, 188.1295, 185.4015, 185.4718, 185.5125, 
    186.5947,
  201.5891, 214.4656, 211.1084, 195.0356, 184.4937, 179.0104, 185.202, 
    176.1729, 178.397, 184.8009, 185.9049, 184.4273, 184.5133, 186.1711, 
    187.4643,
  195.9348, 210.4459, 208.1397, 203.946, 192.2815, 179.7162, 181.0757, 
    196.4434, 197.3809, 194.6633, 185.9625, 184.5714, 184.3345, 185.1022, 
    185.9084,
  199.3089, 209.1952, 212.8332, 213.8449, 209.1742, 186.851, 179.1143, 
    190.1855, 195.2004, 193.1187, 189.2471, 185.4999, 184.7785, 184.2248, 
    185.0802,
  206.3103, 198.8073, 210.074, 209.437, 206.5927, 183.4142, 175.1222, 
    185.1892, 194.6791, 190.4868, 186.8972, 185.0007, 184.1116, 182.8951, 
    184.0399,
  201.4758, 192.5716, 201.3339, 208.5398, 204.9791, 188.8174, 176.989, 
    177.972, 189.7123, 187.4151, 185.9045, 184.8194, 182.9433, 182.9662, 
    184.1239,
  199.001, 184.7259, 188.4149, 202.0248, 205.1451, 188.186, 175.6545, 
    178.7069, 185.5152, 187.7138, 189.7325, 186.1385, 184.0986, 183.804, 
    183.3752,
  185.2715, 192.6319, 186.0857, 185.2472, 177.3334, 175.7768, 182.5788, 
    183.3665, 183.0627, 172.0358, 170.942, 179.5115, 180.8765, 172.6329, 
    165.6677,
  191.8002, 197.9002, 196.536, 188.527, 174.7984, 173.004, 181.765, 184.8028, 
    182.7025, 182.4227, 175.521, 182.9742, 186.2656, 170.4446, 165.881,
  199.4068, 205.3376, 207.2247, 196.7202, 181.6298, 169.6892, 178.2972, 
    183.6144, 183.6794, 183.9042, 183.516, 183.8793, 185.6754, 185.6741, 
    177.0113,
  187.4877, 196.952, 201.6185, 197.2723, 193.7216, 184.3435, 171.1503, 
    181.5565, 185.4904, 184.5421, 182.2552, 181.5976, 183.1473, 184.5173, 
    182.5516,
  177.299, 187.2764, 209.6947, 210.3493, 198.4312, 188.9372, 188.2046, 
    174.9776, 173.1912, 182.6593, 182.1205, 181.2908, 182.3511, 183.9216, 
    184.5588,
  166.8648, 189.2411, 202.6355, 213.2393, 215.2116, 195.8716, 188.3834, 
    196.1351, 193.6355, 193.7698, 186.3372, 183.078, 182.2228, 181.9905, 
    183.0242,
  165.2561, 189.2827, 202.1444, 206.4252, 215.1063, 203.8137, 194.1149, 
    188.2348, 189.9771, 192.5319, 189.039, 184.0099, 182.9106, 181.8342, 
    182.8427,
  179.3326, 186.5064, 195.9398, 200.7243, 205.1757, 207.9202, 194.1519, 
    186.5748, 188.0854, 187.9611, 187.1273, 184.3461, 182.9546, 181.6173, 
    181.7536,
  182.7208, 187.2477, 191.9195, 196.2721, 200.2917, 204.6595, 199.8637, 
    189.8464, 185.8597, 183.8984, 185.1208, 184.3305, 182.8548, 181.4494, 
    182.2802,
  182.4231, 184.7164, 184.0787, 191.0428, 199.0865, 200.7153, 195.7757, 
    187.9166, 183.8364, 182.4843, 187.3459, 184.7582, 183.4005, 183.4628, 
    182.9584,
  160.7696, 168.2033, 174.7543, 184.5515, 187.6063, 183.6973, 180.9739, 
    179.9174, 178.0426, 165.0125, 164.6252, 169.9594, 169.318, 165.9119, 
    159.9372,
  161.1606, 162.7562, 173.5098, 180.1268, 183.3852, 180.773, 181.0321, 
    179.4662, 176.8211, 174.9496, 168.4965, 176.3308, 179.9657, 162.9606, 
    159.9603,
  160.6807, 158.2667, 168.7054, 177.0484, 186.5096, 174.1678, 179.9176, 
    179.05, 176.2417, 176.2727, 176.9124, 178.198, 179.2894, 178.0894, 
    168.7063,
  159.6525, 157.2713, 163.305, 172.9014, 191.7647, 194.4458, 172.2727, 
    177.6585, 177.4691, 175.2641, 176.2605, 177.5812, 178.9767, 177.7379, 
    172.6407,
  161.082, 157.4058, 159.5945, 169.708, 188.3278, 198.2341, 202.0635, 
    171.8451, 167.9776, 175.3985, 175.5549, 177.9821, 181.3066, 180.8059, 
    175.2428,
  163.8017, 160.2509, 160.4445, 163.7538, 178.4066, 195.9815, 195.8282, 
    201.5042, 192.3412, 190.3525, 182.9935, 180.1291, 179.6023, 179.0416, 
    175.7888,
  180.8083, 174.5976, 167.3491, 160.1775, 176.4186, 193.7973, 202.1306, 
    196.8275, 193.1261, 192.5486, 187.4941, 180.7532, 179.4657, 179.8012, 
    177.3868,
  174.3613, 171.3915, 164.9117, 164.3994, 169.3242, 191.0569, 201.0918, 
    201.8215, 198.0089, 190.5064, 186.7572, 182.9666, 179.7763, 178.814, 
    177.3264,
  178.2391, 172.6751, 169.4738, 163.0239, 166.5253, 176.1024, 192.0115, 
    201.4451, 198.6069, 195.2388, 190.4303, 187.0963, 182.2645, 177.9681, 
    177.2734,
  180.1445, 171.8622, 168.9377, 165.4529, 164.4344, 168.858, 175.8394, 
    186.6412, 188.6385, 194.1017, 192.5347, 189.5122, 186.0781, 183.5708, 
    178.9665,
  172.7105, 171.013, 168.1794, 167.8967, 163.4906, 169.0422, 176.4349, 
    178.5678, 176.3661, 163.7409, 162.6645, 168.3547, 165.8123, 165.247, 
    157.4241,
  172.9319, 171.0119, 170.8714, 168.799, 162.9783, 167.9005, 177.1131, 
    177.7816, 173.8795, 167.7878, 166.1994, 174.5796, 175.8729, 161.7503, 
    157.8817,
  173.1839, 170.7466, 179.8717, 171.0692, 166.1791, 163.8876, 176.2432, 
    176.9522, 171.7772, 168.8341, 170.9987, 174.3366, 176.0363, 176.0501, 
    169.5111,
  175.3279, 176.2291, 174.8303, 183.4836, 174.0567, 178.1009, 168.7421, 
    174.355, 171.6029, 163.4464, 167.1507, 169.1012, 172.9753, 174.2393, 
    171.6865,
  177.4659, 177.274, 175.0711, 171.4964, 176.5712, 187.0158, 191.7296, 
    170.3708, 165.7416, 165.9286, 164.4967, 168.2312, 171.0267, 174.0667, 
    173.3419,
  182.1756, 178.0024, 187.2613, 186.7654, 174.8166, 179.9364, 203.5338, 
    199.9397, 189.1569, 178.9454, 170.5795, 170.0508, 171.9428, 170.9724, 
    170.0706,
  182.6353, 179.546, 183.438, 183.7675, 180.8604, 176.552, 203.6301, 
    201.7583, 195.3739, 185.1497, 175.1388, 169.1233, 170.8676, 170.2886, 
    171.7896,
  189.6633, 176.854, 177.9618, 188.6273, 190.4259, 178.8497, 185.3236, 
    202.5344, 199.422, 185.4647, 175.5232, 169.9192, 169.7804, 170.9393, 
    169.7312,
  190.1446, 177.1702, 174.2009, 182.2984, 185.8141, 187.6646, 180.5325, 
    188.544, 195.4005, 186.9103, 181.4668, 174.0757, 171.9969, 169.8589, 
    169.4613,
  196.5093, 180.4438, 176.5299, 180.9852, 183.9937, 192.9175, 188.472, 
    200.8427, 192.5629, 189.521, 189.4718, 181.3754, 177.0409, 174.57, 
    172.8329,
  191.1314, 186.0858, 178.2341, 171.78, 169.3315, 168.35, 172.7629, 172.4496, 
    172.8654, 162.974, 162.344, 163.9885, 160.448, 160.6003, 155.4696,
  191.3018, 188.4957, 180.8428, 173.2546, 168.7653, 169.4185, 172.077, 
    173.9566, 172.6877, 169.519, 165.0847, 171.2766, 171.2203, 157.3017, 
    154.1853,
  193.4494, 189.4702, 181.43, 171.9501, 173.1947, 169.3873, 174.5515, 175.47, 
    172.4792, 169.3426, 172.4804, 172.8482, 172.5421, 170.7704, 164.1956,
  194.7932, 193.1214, 182.4025, 178.6543, 172.2573, 177.1042, 168.1005, 
    173.2547, 170.9781, 168.4058, 170.5358, 172.2842, 171.7785, 170.3385, 
    167.9155,
  197.3885, 195.6236, 187.7349, 180.6966, 185.9074, 175.4245, 192.182, 
    167.6088, 162.4939, 166.0145, 170.4191, 172.8645, 171.7757, 170.0492, 
    169.183,
  204.2597, 196.6863, 188.6802, 178.229, 183.6552, 182.311, 195.4764, 
    197.0228, 185.8171, 178.866, 175.0182, 175.3308, 172.9148, 168.8975, 
    165.3789,
  208.326, 205.1787, 192.4909, 174.5362, 190.7074, 183.7381, 196.2157, 
    199.4155, 187.3912, 182.0283, 179.0285, 175.8509, 173.6871, 167.434, 
    164.1853,
  222.7256, 212.4416, 188.4799, 179.4864, 185.0863, 190.9214, 182.3547, 
    209.5815, 195.7054, 179.4009, 175.6127, 175.1866, 172.5941, 168.2175, 
    163.0484,
  224.1189, 210.8874, 188.6246, 172.3206, 180.0033, 194.3289, 188.9953, 
    202.7226, 189.148, 179.9143, 174.1509, 172.6102, 171.1512, 166.1735, 
    163.3572,
  220.4164, 209.6077, 178.6585, 176.6035, 184.4393, 190.468, 201.4509, 
    199.7828, 186.8988, 180.292, 179.2207, 173.0174, 171.7145, 166.1812, 
    163.7532,
  166.478, 168.3862, 169.8067, 175.9836, 176.5101, 174.7259, 177.251, 
    175.5779, 171.1313, 164.6014, 163.6918, 164.2197, 158.4053, 158.2165, 
    152.872,
  166.3453, 167.4509, 170.938, 175.3896, 176.7599, 175.5866, 177.1751, 
    177.6281, 170.6422, 167.9009, 166.8473, 171.292, 169.5581, 154.6752, 
    151.4978,
  167.1715, 170.1705, 172.8959, 173.2699, 175.7718, 178.1778, 174.6215, 
    176.3746, 172.8412, 169.3549, 170.9169, 171.6648, 171.1552, 168.618, 
    162.0596,
  166.9486, 167.0254, 172.278, 176.586, 176.3252, 181.4615, 173.6335, 
    172.795, 172.9247, 170.9401, 169.8536, 170.4418, 169.6595, 168.8453, 
    166.7471,
  164.2107, 166.6663, 170.2965, 173.6707, 179.1263, 178.1682, 180.2076, 
    169.8504, 164.7814, 168.3439, 170.6266, 170.6496, 169.9096, 169.636, 
    168.8548,
  172.5625, 169.7837, 176.4495, 176.6185, 179.5857, 178.1681, 175.0277, 
    188.685, 187.5836, 185.2083, 176.127, 172.5782, 170.742, 168.873, 168.3482,
  207.748, 186.4121, 182.7258, 181.3929, 178.6824, 186.4522, 186.3622, 
    186.029, 182.2762, 184.7952, 180.039, 173.2177, 171.2159, 168.6822, 
    168.0824,
  224.4503, 212.0718, 196.5245, 179.3752, 178.8491, 191.0355, 195.6415, 
    191.4267, 190.9167, 178.1439, 176.0505, 172.8553, 170.7317, 168.2554, 
    167.9697,
  215.6465, 214.8938, 195.6672, 182.2483, 180.881, 194.1808, 196.2609, 
    192.6431, 186.2635, 177.5661, 174.3692, 172.4847, 170.634, 167.2253, 
    166.7652,
  216.1772, 204.2723, 186.8994, 179.3907, 187.6693, 193.1129, 192.6436, 
    195.8208, 179.6184, 177.1568, 179.8493, 173.58, 171.067, 168.4861, 167.578,
  181.4006, 177.7977, 170.0664, 167.6595, 166.7792, 164.2089, 162.3689, 
    163.2138, 165.8722, 166.4436, 164.9159, 167.6619, 162.2676, 160.0512, 
    155.9764,
  170.7948, 170.4935, 167.2454, 164.5576, 163.0405, 165.4556, 164.4396, 
    166.7002, 166.6079, 167.8258, 165.9678, 172.1952, 172.9225, 157.0754, 
    152.9166,
  174.7279, 175.446, 173.7182, 170.4279, 167.8543, 165.6625, 163.322, 
    163.6646, 165.3363, 170.076, 169.3496, 172.6266, 174.3069, 172.233, 
    161.9637,
  192.6327, 191.8683, 183.5416, 173.6685, 169.6862, 170.2331, 165.3626, 
    163.1304, 165.8917, 169.2088, 171.884, 172.4113, 172.683, 171.1699, 
    167.9096,
  205.8485, 200.4671, 188.4624, 176.7874, 171.393, 169.3466, 175.4502, 
    168.0029, 169.8813, 169.0382, 171.7255, 172.701, 172.1432, 171.7009, 
    171.9468,
  210.0247, 206.9654, 197.1485, 186.0815, 177.5789, 177.9721, 176.2605, 
    186.9721, 182.1529, 182.0581, 178.8422, 175.013, 172.6799, 170.366, 
    169.9454,
  221.623, 213.7257, 199.0602, 186.5241, 176.5657, 180.1266, 195.7169, 
    186.3241, 183.0362, 187.5292, 182.7426, 175.054, 172.7569, 169.4143, 
    168.8446,
  220.8308, 212.7672, 190.6584, 182.2237, 170.1011, 174.2356, 194.1763, 
    191.7615, 187.6423, 180.7034, 177.8784, 174.5887, 172.0444, 168.6006, 
    167.7076,
  212.2419, 201.0372, 188.2444, 171.725, 165.0232, 174.9545, 183.4708, 
    183.6317, 182.6427, 177.2662, 174.9308, 173.2552, 170.817, 168.2425, 
    166.745,
  216.0289, 208.2375, 193.3187, 178.4707, 174.0358, 183.5513, 183.8379, 
    187.9964, 177.0219, 175.6666, 178.2328, 173.3955, 171.4536, 169.5648, 
    168.562,
  185.9361, 184.4274, 184.1617, 183.1974, 181.4623, 179.8279, 178.2845, 
    172.8754, 171.5522, 170.6972, 168.1136, 168.8416, 165.3358, 161.4097, 
    159.9989,
  178.5915, 177.119, 170.7689, 175.3925, 180.229, 181.2983, 176.4449, 
    177.0169, 171.9814, 169.0875, 167.8306, 167.1469, 168.3191, 162.4476, 
    160.4049,
  190.8187, 184.378, 175.3083, 167.825, 167.8108, 174.5708, 172.5, 171.5925, 
    174.3074, 170.0639, 171.661, 168.9249, 165.5687, 165.9458, 164.2476,
  214.3379, 203.3923, 194.4197, 182.1098, 173.034, 175.7978, 170.189, 
    171.045, 171.0753, 172.3801, 171.6471, 169.6376, 168.7343, 165.7007, 
    165.1032,
  219.1346, 214.8444, 204.4563, 198.2721, 181.3595, 175.2894, 179.45, 
    175.1653, 179.8508, 169.7688, 169.8957, 169.153, 168.1687, 167.8366, 
    168.1967,
  223.2824, 216.0713, 204.5733, 195.9732, 180.5418, 174.6087, 179.8774, 
    181.3522, 178.1612, 175.8398, 172.8416, 171.8243, 169.5244, 168.642, 
    168.7205,
  224.9825, 215.9173, 207.1808, 194.4066, 179.79, 183.7701, 189.974, 
    178.6213, 182.139, 183.0663, 175.862, 171.0129, 169.1711, 167.1716, 
    168.9124,
  222.8335, 216.1134, 212.9346, 202.4344, 183.7906, 192.569, 183.3448, 
    183.0964, 181.9746, 178.2222, 175.2475, 172.023, 170.3252, 168.074, 
    168.5882,
  220.1729, 217.8751, 212.8803, 198.5538, 190.181, 189.497, 183.0446, 
    184.8053, 182.4112, 177.9495, 174.1245, 173.2157, 171.0472, 168.8431, 
    168.3259,
  222.1404, 215.1173, 210.426, 199.0352, 186.9793, 184.6302, 180.9359, 
    188.6669, 179.8921, 176.6857, 178.0779, 173.7811, 172.5935, 170.4701, 
    169.2114,
  201.137, 200.598, 197.7709, 195.1946, 191.07, 189.1099, 188.3615, 188.4368, 
    186.9038, 177.2177, 176.1898, 175.7781, 175.2661, 173.0575, 170.8612,
  204.6354, 203.6681, 201.2054, 196.7982, 189.3214, 186.8484, 186.854, 
    187.7634, 185.8832, 184.6823, 180.1917, 180.1934, 180.8129, 173.4452, 
    171.8294,
  218.9124, 215.113, 208.6862, 200.3769, 194.062, 183.5244, 178.0446, 
    177.9584, 180.8443, 182.474, 182.6483, 182.6546, 179.4995, 177.375, 
    174.9554,
  220.3008, 221.6018, 219.3554, 208.8725, 199.479, 190.2938, 177.1996, 
    171.5239, 172.6688, 177.7074, 178.5134, 178.5735, 179.6869, 177.7137, 
    175.9337,
  222.6054, 221.6855, 213.3962, 218.2912, 203.3975, 186.7951, 183.3094, 
    175.2561, 170.4503, 164.0727, 169.0855, 174.4894, 175.4616, 176.326, 
    175.9172,
  223.0204, 220.0336, 214.4631, 215.946, 204.9157, 185.8612, 177.6879, 
    171.9068, 163.6384, 161.201, 166.2855, 173.0065, 172.8644, 171.9967, 
    171.5938,
  221.4343, 221.9093, 216.0124, 207.9754, 202.5792, 200.5546, 189.9064, 
    178.9131, 170.5401, 169.2531, 169.168, 169.4072, 170.0011, 168.9229, 
    171.1932,
  223.5081, 223.2796, 218.5562, 212.4082, 211.1415, 205.6401, 191.8141, 
    190.2662, 189.0375, 177.2652, 168.8704, 168.4955, 167.5969, 167.3934, 
    171.2308,
  222.9599, 217.2496, 216.5479, 217.7561, 212.9341, 199.1613, 192.4662, 
    186.1935, 184.1102, 176.6313, 168.2029, 166.5806, 164.4353, 166.7077, 
    168.2617,
  218.0827, 219.0242, 216.8354, 210.4279, 211.8744, 190.5135, 184.6609, 
    185.3878, 180.9941, 175.7982, 172.5324, 165.5814, 163.4525, 165.2198, 
    167.3323,
  198.939, 200.4755, 201.2559, 195.9594, 194.5145, 191.8964, 191.0119, 
    183.6259, 181.5524, 176.84, 169.8398, 164.7493, 164.1519, 166.0679, 
    167.644,
  204.4088, 204.2846, 204.301, 200.1799, 195.0274, 195.1188, 188.2293, 
    188.5228, 186.6232, 184.6713, 181.0763, 178.8566, 171.4597, 166.9815, 
    167.7378,
  205.2804, 217.3899, 212.8153, 202.8078, 199.3296, 190.6413, 188.9784, 
    185.2427, 186.6859, 184.898, 182.7755, 184.8805, 178.4239, 172.678, 
    171.6138,
  214.7155, 220.7104, 215.3476, 213.5023, 204.3632, 200.0417, 190.6676, 
    191.5457, 189.2368, 188.8189, 186.197, 186.0777, 183.5424, 180.1349, 
    175.5511,
  216.7589, 221.4525, 216.5313, 217.0653, 209.6936, 210.4752, 201.8719, 
    187.39, 186.8803, 180.205, 178.9237, 179.7358, 181.5675, 180.2549, 
    177.7995,
  208.8435, 222.1394, 213.649, 208.644, 206.8466, 204.8896, 194.3791, 
    196.5057, 193.6647, 188.3182, 178.4833, 173.4153, 174.6557, 175.7855, 
    173.4257,
  213.9571, 225.0484, 212.1274, 201.9658, 200.428, 188.2744, 191.5245, 
    193.9815, 196.364, 192.4842, 179.888, 170.6204, 172.0434, 168.6493, 
    171.9727,
  222.0314, 224.4347, 209.8405, 194.7057, 193.8001, 198.0221, 190.1376, 
    192.0837, 193.2535, 189.7954, 180.3781, 168.6829, 168.1433, 167.8034, 
    166.4569,
  225.8037, 212.5829, 189.6076, 185.7094, 187.9337, 182.7154, 188.747, 
    189.5729, 189.61, 185.6216, 177.9126, 168.9242, 165.1539, 163.5357, 
    166.6832,
  210.1907, 196.6497, 175.9524, 174.5143, 183.2454, 182.1584, 188.9381, 
    186.3952, 183.6035, 178.3698, 177.8573, 166.5419, 161.9963, 161.2855, 
    172.1433,
  201.3077, 206.9236, 199.1504, 200.8688, 197.2352, 194.3553, 187.0318, 
    181.707, 179.6975, 180.8202, 182.3737, 183.5744, 181.1294, 176.8055, 
    174.016,
  208.7455, 204.8034, 200.7045, 200.3814, 195.2201, 189.8144, 182.3432, 
    176.4996, 179.0598, 180.827, 183.721, 186.6646, 185.8595, 177.636, 
    172.6492,
  210.9603, 211.2, 210.6733, 199.338, 188.4558, 175.935, 179.6363, 169.0557, 
    173.8833, 181.5927, 186.0819, 188.7775, 187.0974, 180.554, 172.6246,
  210.323, 215.5924, 199.9531, 193.6235, 169.2417, 164.6452, 162.9282, 
    173.6653, 176.143, 179.3794, 186.2676, 188.9195, 187.9163, 183.1179, 
    175.159,
  221.3375, 214.7017, 196.2718, 169.9489, 154.6029, 157.1804, 165.5013, 
    169.4212, 177.8594, 181.4758, 188.1699, 189.3836, 187.4433, 183.9132, 
    180.7028,
  206.2656, 203.5202, 177.3271, 154.6332, 153.0301, 165.1969, 169.5224, 
    178.4566, 187.6683, 190.3321, 189.6664, 188.4615, 186.3886, 184.8781, 
    181.8454,
  202.1028, 188.7193, 156.3155, 153.0055, 155.6083, 173.3039, 181.2402, 
    185.8304, 186.4222, 189.0144, 189.7861, 185.5667, 183.3308, 180.1756, 
    179.682,
  196.9222, 164.4534, 149.7614, 148.3932, 159.7646, 181.1273, 190.8602, 
    193.8705, 188.3065, 184.2405, 184.2908, 182.5663, 181.8146, 176.757, 
    177.1372,
  186.9677, 156.4128, 143.8653, 151.5721, 162.6754, 185.3759, 196.259, 
    195.6034, 184.2768, 183.8835, 182.7102, 181.8069, 179.593, 173.3635, 
    173.6883,
  170.5959, 155.8853, 148.7005, 157.2275, 177.7543, 191.084, 193.8798, 
    194.0478, 184.4082, 180.5956, 179.7107, 182.0059, 176.9849, 172.695, 
    170.8642,
  202.229, 207.7352, 199.7722, 200.0305, 178.258, 167.9727, 171.8902, 
    174.5194, 174.3485, 173.67, 176.3847, 176.4626, 177.6967, 180.3743, 
    180.0861,
  209.692, 205.4255, 202.285, 183.504, 165.4036, 168.7363, 171.9462, 
    175.9943, 181.0437, 184.0869, 181.6712, 178.2309, 179.7339, 178.4809, 
    180.3243,
  212.6818, 206.4642, 199.6864, 170.7939, 161.1975, 167.659, 183.7512, 
    184.3246, 184.2103, 187.7095, 182.1074, 175.687, 176.2946, 179.8106, 
    183.955,
  205.1552, 204.4346, 177.9214, 166.353, 164.4437, 179.5303, 186.5881, 
    196.0936, 193.6555, 185.3309, 178.5414, 179.5888, 184.3356, 186.7566, 
    187.5929,
  207.7267, 199.3423, 172.8016, 168.349, 171.3702, 188.1026, 199.9558, 
    191.7853, 185.5161, 187.1343, 184.366, 186.8019, 188.8631, 188.718, 
    185.7857,
  205.7931, 193.2303, 176.9594, 169.4131, 169.4384, 185.6118, 196.4596, 
    189.5744, 193.5157, 192.2303, 186.6828, 187.6247, 187.5094, 185.9406, 
    186.8201,
  202.2805, 192.4953, 182.9661, 174.6081, 170.0408, 174.9957, 185.5143, 
    187.1301, 188.3983, 190.6951, 186.8669, 186.0805, 187.4975, 185.5372, 
    181.8047,
  203.4386, 194.6193, 185.8916, 180.3146, 168.8974, 165.273, 174.3004, 
    181.9896, 181.029, 183.6129, 182.7975, 184.0866, 182.307, 180.696, 
    179.4954,
  204.3684, 197.5087, 189.776, 178.8448, 165.6551, 166.0237, 165.437, 
    172.1369, 174.8944, 176.4722, 177.8181, 179.2517, 179.6257, 178.1369, 
    177.9933,
  202.291, 196.5675, 190.6381, 188.9395, 172.8465, 166.3956, 164.3654, 
    165.6178, 167.8132, 170.2978, 172.5614, 177.3634, 178.7883, 177.8752, 
    177.5699,
  204.3727, 205.5432, 199.3987, 198.9084, 193.8961, 192.6417, 192.5794, 
    183.1397, 177.3069, 181.0682, 187.8699, 188.6855, 184.3013, 183.8764, 
    180.2226,
  207.5947, 204.7762, 200.3936, 197.3153, 190.2737, 193.1381, 194.1724, 
    181.4731, 173.5026, 181.1958, 185.42, 192.2168, 189.6246, 180.7171, 
    178.1054,
  215.2231, 216.1561, 208.3902, 197.3712, 190.7881, 186.937, 187.9907, 
    169.6847, 167.3338, 171.829, 183.2462, 191.8826, 192.0362, 188.0683, 
    181.5404,
  211.6674, 201.018, 200.0387, 199.7684, 194.7812, 192.5815, 185.5556, 
    175.3914, 172.2125, 168.5348, 175.9574, 188.866, 192.1782, 188.6927, 
    185.2937,
  204.2196, 201.9737, 198.8891, 196.0486, 194.2234, 194.4142, 194.1829, 
    188.4, 172.6079, 166.0823, 167.6786, 183.4937, 187.7873, 189.3134, 188.219,
  214.3451, 218.6251, 203.0727, 197.956, 199.788, 197.7984, 185.9522, 
    177.9344, 168.7334, 165.0383, 165.6364, 176.9911, 183.9811, 185.7419, 
    185.0041,
  219.4479, 205.6696, 208.705, 215.0612, 201.0552, 197.6209, 187.2055, 
    175.0476, 170.7408, 170.0706, 169.5007, 172.2345, 180.5729, 181.9111, 
    180.3616,
  210.5738, 217.401, 212.567, 216.581, 200.4428, 197.1111, 186.4124, 180.507, 
    181.767, 177.2554, 170.9701, 172.705, 177.4881, 181.7496, 177.5605,
  209.698, 209.2333, 202.8481, 214.1317, 196.703, 194.0285, 190.3497, 
    186.2864, 182.9395, 181.927, 178.0585, 176.2387, 177.434, 175.8529, 
    176.841,
  202.8332, 202.9368, 205.486, 208.5965, 204.7287, 201.9749, 193.7406, 
    193.1904, 192.0376, 189.1043, 185.0792, 178.5037, 176.8747, 179.0568, 
    177.8408,
  175.2228, 187.9012, 199.4427, 202.8709, 201.0859, 201.243, 201.117, 
    198.5177, 193.4387, 180.7805, 184.1809, 188.3084, 184.9035, 178.4158, 
    176.7191,
  180.8177, 195.5332, 201.7409, 202.7208, 200.9991, 201.2199, 201.0866, 
    203.3819, 197.7207, 190.9062, 181.575, 188.6385, 187.1126, 176.2471, 
    174.2617,
  199.4154, 199.6942, 201.122, 201.374, 203.6178, 200.2581, 203.4118, 
    197.6539, 193.4328, 192.4292, 189.5847, 187.593, 188.1203, 187.4241, 
    185.0393,
  202.9856, 201.5832, 202.8405, 203.3266, 203.4547, 203.193, 199.2478, 
    206.0317, 199.7365, 193.7758, 190.7253, 187.7478, 183.7887, 185.9355, 
    186.8797,
  202.9508, 202.4919, 202.9273, 203.0552, 203.1005, 201.3, 199.0299, 
    194.7399, 192.5831, 193.4093, 191.316, 190.5727, 186.5332, 184.0633, 
    188.6682,
  203.0346, 204.4895, 203.5004, 202.9516, 201.9325, 199.3391, 191.577, 
    190.2457, 192.2038, 192.986, 193.0688, 193.6853, 189.0792, 185.6307, 
    183.9385,
  200.5421, 209.4431, 202.6678, 204.719, 199.9878, 194.8788, 189.0722, 
    186.5546, 189.4042, 190.1202, 194.4409, 195.579, 193.1849, 187.5262, 
    184.7669,
  209.5017, 214.1681, 210.0848, 202.4665, 193.6355, 190.9653, 187.7468, 
    187.3191, 190.6036, 192.3267, 193.9281, 196.555, 195.3041, 192.0236, 
    186.1132,
  212.9641, 212.6061, 210.7861, 200.2177, 196.9084, 190.7924, 190.5083, 
    186.0294, 193.236, 194.9742, 195.0412, 199.3432, 196.3987, 193.3738, 
    189.6475,
  211.8967, 209.1337, 207.1206, 190.0883, 186.3555, 188.077, 187.0372, 
    193.7527, 192.7626, 195.1213, 196.451, 195.7617, 195.502, 194.8823, 
    191.3828,
  180.5681, 197.4022, 202.8646, 205.2315, 200.6681, 198.2383, 196.1381, 
    190.4534, 186.1688, 187.789, 181.6593, 185.4892, 175.3155, 178.5193, 
    179.6768,
  193.4261, 200.9077, 204.8512, 206.325, 201.7239, 198.7204, 195.6855, 
    189.1102, 182.2368, 185.87, 183.6016, 184.5618, 185.2551, 183.1731, 
    181.3422,
  199.9434, 204.8558, 207.0419, 204.7372, 202.0381, 198.4895, 199.144, 
    183.1518, 178.6062, 179.9622, 185.0804, 180.9255, 184.7184, 184.611, 
    179.2007,
  205.6835, 208.2839, 206.2828, 205.3035, 203.5209, 201.899, 195.7424, 
    184.8091, 182.9083, 179.9218, 180.7608, 178.5344, 178.1389, 175.5392, 
    177.0741,
  209.7725, 210.6791, 208.097, 207.0191, 204.3085, 200.0119, 192.8599, 
    188.0676, 186.7369, 179.4064, 178.2937, 175.7941, 174.5933, 173.1417, 
    174.3118,
  212.9328, 213.0701, 213.1094, 209.8327, 208.7395, 197.0592, 184.8454, 
    181.6285, 176.9969, 169.0521, 170.1604, 174.007, 171.2271, 171.1843, 
    171.2754,
  216.3716, 212.2275, 211.2487, 211.6117, 210.0223, 191.7839, 175.2406, 
    168.5055, 167.9942, 167.3295, 167.7045, 170.8378, 168.7739, 167.1587, 
    166.608,
  217.3408, 212.1824, 211.6674, 211.7829, 195.1115, 186.458, 172.9527, 
    166.6086, 162.4677, 159.8269, 163.2548, 162.4606, 164.9411, 161.734, 
    166.3529,
  215.849, 211.6161, 204.9158, 196.1373, 193.8128, 182.7525, 170.9818, 
    161.9824, 160.8105, 155.2305, 159.7045, 156.8757, 158.2725, 161.5821, 
    163.2784,
  204.4634, 193.6946, 187.5359, 185.9227, 185.8037, 182.2688, 173.2864, 
    164.7658, 160.7758, 157.7911, 155.5839, 157.878, 154.6056, 155.4387, 
    160.9957,
  195.1595, 208.9485, 206.2002, 201.516, 194.9736, 194.6325, 197.1393, 
    189.4294, 184.9838, 178.838, 177.5581, 173.2391, 172.0721, 177.2769, 
    169.7825,
  199.7376, 206.7042, 208.0409, 202.2363, 195.9175, 196.1006, 195.9254, 
    195.8199, 193.74, 183.4486, 176.0206, 171.5843, 173.3012, 175.5407, 
    176.5692,
  206.2942, 209.5781, 211.9361, 206.3188, 200.4786, 191.2077, 202.2846, 
    192.4264, 185.4487, 190.4058, 187.384, 176.2435, 174.6687, 175.4193, 
    177.5896,
  215.2034, 216.5201, 219.4892, 216.9355, 210.6898, 203.2328, 199.0992, 
    189.8642, 175.9258, 170.9038, 182.4126, 180.3271, 176.3693, 174.1982, 
    177.2271,
  214.9829, 218.7109, 220.7153, 220.0223, 214.8723, 209.5607, 195.8073, 
    190.9946, 183.7964, 174.774, 173.7272, 178.9706, 181.161, 185.8334, 
    178.9015,
  214.9785, 216.341, 218.3452, 220.1233, 218.6875, 209.5947, 199.0288, 
    193.7593, 183.7805, 180.7762, 186.8007, 190.6015, 186.4295, 189.9576, 
    188.6447,
  214.162, 213.5255, 216.9039, 217.4697, 217.4894, 204.8481, 199.3594, 
    188.9763, 187.5625, 195.3712, 196.5189, 196.7485, 199.5254, 194.7963, 
    192.7882,
  215.8695, 215.2139, 218.06, 219.3787, 210.5606, 203.5757, 199.2202, 
    193.6647, 202.8627, 203.8951, 201.635, 204.1803, 202.0417, 198.9839, 
    194.488,
  218.153, 218.1477, 212.7593, 205.4177, 196.3853, 200.1575, 197.9361, 
    203.5179, 205.2466, 209.4538, 209.926, 208.4253, 200.5834, 196.0922, 
    193.2495,
  215.2352, 209.2097, 202.705, 189.4467, 190.3101, 197.1825, 204.411, 
    206.7478, 210.7153, 208.396, 211.2988, 206.5797, 199.3755, 196.8396, 
    191.1571,
  199.3675, 201.1226, 205.6254, 205.941, 203.6208, 201.4194, 203.0839, 
    196.8361, 193.4968, 189.1066, 189.6252, 191.409, 189.5607, 189.2242, 
    186.7863,
  198.1215, 197.5201, 204.0715, 204.9231, 202.3248, 200.7848, 203.187, 
    198.8969, 197.0233, 193.7061, 193.1524, 194.2577, 194.6769, 196.7068, 
    192.155,
  191.4934, 193.6052, 197.0729, 198.1019, 203.1504, 200.6148, 205.0927, 
    201.3496, 202.6083, 200.5159, 199.7475, 193.6334, 194.6892, 198.05, 
    193.0619,
  191.9844, 189.1718, 190.9985, 191.6094, 193.0647, 196.3823, 197.3743, 
    195.7983, 200.6351, 198.7643, 198.9138, 195.3037, 194.6776, 195.8422, 
    194.123,
  187.0397, 185.6533, 187.6708, 180.1113, 185.5917, 186.6537, 185.9754, 
    192.9188, 196.7262, 192.7933, 195.9791, 192.6514, 191.6884, 191.1816, 
    188.3362,
  193.832, 189.9705, 186.9846, 184.2106, 182.2473, 180.6964, 184.7343, 
    184.9767, 191.1676, 191.1402, 190.5094, 188.8005, 190.4292, 186.9472, 
    184.0062,
  197.6391, 193.0078, 189.6459, 185.701, 182.0988, 187.7043, 185.1615, 
    187.702, 185.4539, 188.537, 184.0391, 184.6243, 188.2104, 186.1781, 
    182.6918,
  200.5696, 193.4866, 195.1906, 192.8872, 193.7604, 195.3397, 201.3712, 
    206.2444, 201.4651, 191.3162, 187.7361, 187.9473, 186.8998, 185.3306, 
    184.7978,
  202.1246, 199.4647, 200.6838, 201.0996, 210.3558, 210.8041, 212.4534, 
    204.6093, 196.4145, 191.2971, 190.7847, 189.1697, 187.8546, 183.2923, 
    178.8963,
  207.0369, 214.2264, 212.1416, 216.2019, 215.1626, 207.341, 197.7375, 
    194.6712, 189.4048, 188.9298, 187.5429, 186.7601, 184.3527, 177.8828, 
    176.936,
  186.362, 199.4793, 204.4702, 201.5064, 200.9714, 198.0721, 197.2128, 
    191.3372, 186.1103, 180.7702, 177.5011, 177.1512, 177.032, 174.6706, 
    177.3747,
  198.9951, 208.3084, 204.928, 201.9433, 198.3788, 195.7711, 193.3657, 
    189.4035, 190.3139, 180.7467, 173.2765, 173.6443, 172.2686, 171.9184, 
    173.7342,
  208.3218, 207.1472, 205.8305, 200.477, 194.9472, 191.8591, 189.5906, 
    182.7503, 182.7979, 174.8036, 169.4035, 167.3845, 170.3148, 175.5756, 
    178.6121,
  211.4587, 208.8453, 201.3408, 196.66, 192.9271, 192.1318, 187.2817, 
    185.3737, 176.5682, 169.3788, 165.625, 167.7254, 171.9588, 176.3671, 
    177.5774,
  212.6144, 206.0544, 201.8606, 200.7211, 196.0599, 189.3698, 186.0064, 
    184.7909, 179.0144, 166.0368, 168.0686, 174.5596, 178.9288, 181.0039, 
    181.012,
  210.4932, 211.0325, 206.5338, 202.2629, 198.7729, 194.9131, 189.5288, 
    181.8054, 181.213, 179.1825, 175.6949, 181.6176, 179.8876, 182.4542, 
    183.66,
  212.5768, 213.3143, 210.4922, 204.1836, 202.3413, 191.6201, 194.6022, 
    185.5224, 185.6086, 179.5456, 180.3904, 181.6888, 182.6557, 183.3702, 
    187.0869,
  210.0654, 210.2057, 208.9992, 207.6762, 204.8127, 198.8187, 199.2979, 
    197.7268, 185.0305, 183.9921, 182.5292, 184.6395, 182.7209, 183.4508, 
    185.7516,
  217.0168, 210.9196, 211.1508, 206.816, 203.9684, 204.7011, 207.6609, 
    188.7431, 188.9583, 185.7445, 188.0872, 181.944, 181.5333, 180.5652, 
    181.7822,
  219.5653, 213.1706, 206.275, 203.5226, 206.5217, 203.1616, 192.1717, 
    190.0592, 186.2073, 184.2043, 182.0421, 181.5229, 178.2556, 177.5312, 
    178.4748,
  188.1551, 199.5356, 210.9589, 212.2143, 205.8541, 197.4967, 196.0619, 
    194.8857, 197.1316, 192.7615, 193.874, 186.9998, 184.1326, 181.1009, 
    177.6371,
  193.5579, 203.9705, 213.9953, 210.2984, 204.2813, 199.4047, 193.8535, 
    195.0812, 200.8097, 199.6451, 196.5206, 190.0514, 184.8982, 181.1631, 
    180.0778,
  209.0441, 216.5441, 217.0527, 207.4774, 203.1293, 199.1783, 204.5163, 
    195.4631, 197.0341, 198.7757, 196.5691, 194.3801, 187.6492, 185.0584, 
    180.9437,
  218.3556, 220.5432, 218.5039, 206.1816, 199.313, 202.1966, 201.5242, 
    207.4261, 201.4429, 195.5987, 195.0572, 193.8889, 190.0438, 185.2631, 
    186.2272,
  222.7526, 218.9823, 216.5507, 208.0488, 205.0717, 201.4885, 198.3603, 
    200.2304, 198.5838, 197.257, 195.4655, 193.645, 190.8728, 188.6018, 
    182.8673,
  222.1099, 220.2137, 216.4978, 210.8326, 210.036, 202.8661, 194.303, 
    196.872, 196.9413, 196.795, 195.4931, 189.0912, 189.0091, 188.0452, 
    183.6048,
  220.0483, 218.3685, 216.6132, 214.2702, 213.0801, 203.7045, 196.4167, 
    193.0627, 191.0088, 190.3575, 189.8581, 187.7747, 190.4066, 186.8241, 
    187.4658,
  225.8829, 220.6426, 216.2462, 214.022, 210.948, 200.2318, 194.0554, 
    193.0922, 187.0437, 183.5318, 181.9597, 185.6269, 184.9256, 186.3759, 
    184.0785,
  226.9079, 221.7666, 218.354, 212.527, 203.7512, 195.1725, 191.9288, 
    187.9048, 184.0441, 180.1928, 181.0595, 184.6977, 185.4875, 180.4512, 
    179.3387,
  226.2915, 222.0146, 211.9372, 199.5522, 189.097, 187.0114, 188.011, 
    178.7499, 176.3721, 177.513, 179.159, 180.4532, 180.5079, 178.5222, 
    179.251,
  185.9149, 188.3181, 199.3785, 210.5087, 210.395, 212.3794, 212.0359, 
    208.886, 199.2099, 198.5671, 198.2734, 196.7849, 194.15, 181.9129, 
    175.3031,
  187.7746, 192.6179, 204.3523, 206.7214, 213.4958, 217.6848, 215.1716, 
    209.6732, 209.3009, 199.589, 194.2669, 191.1259, 185.0802, 180.769, 
    176.0489,
  202.8151, 204.829, 211.2661, 213.43, 216.2475, 215.2336, 214.1919, 
    193.4666, 184.5062, 188.7486, 186.9967, 188.7548, 180.3971, 172.3213, 
    171.8293,
  207.7875, 215.682, 218.4554, 220.1885, 218.5678, 218.0806, 208.1086, 
    197.1832, 185.8992, 178.8485, 188.45, 184.189, 175.3887, 178.9883, 
    176.5416,
  216.1966, 218.3795, 220.6631, 221.7017, 220.093, 217.6751, 213.8169, 
    201.3846, 196.9154, 192.8242, 184.3258, 187.4557, 180.0593, 177.9717, 
    173.393,
  217.8552, 222.2033, 221.0446, 223.0901, 220.0845, 219.04, 213.0298, 
    203.3393, 201.4414, 191.5633, 188.7326, 190.3646, 184.772, 178.2007, 
    175.171,
  220.6161, 220.7248, 221.0257, 219.7534, 220.9865, 215.8641, 211.5527, 
    202.1963, 195.4531, 195.9601, 188.3924, 189.3708, 184.065, 175.176, 
    171.4156,
  220.2152, 220.8093, 220.712, 220.1187, 219.5198, 214.3557, 213.1702, 
    206.5105, 203.2709, 198.9028, 193.9539, 189.1464, 177.3031, 171.926, 
    171.4735,
  221.4151, 220.1815, 221.0228, 221.0107, 217.2341, 214.086, 214.6173, 
    209.7948, 203.3855, 196.9648, 195.5969, 184.2618, 174.4667, 174.3918, 
    164.8985,
  219.0371, 218.5253, 218.734, 216.261, 209.3667, 207.6123, 212.1129, 
    208.5496, 201.3807, 196.8587, 191.5772, 177.5129, 173.7161, 168.7015, 
    168.2911,
  185.263, 189.3972, 184.8334, 188.2115, 189.9402, 193.9083, 199.182, 
    204.6864, 204.3806, 203.1179, 202.3388, 204.4013, 204.1433, 203.9069, 
    198.6311,
  188.7037, 193.7925, 190.3229, 192.3455, 192.8994, 199.8355, 194.5164, 
    203.6855, 209.5079, 205.6751, 201.8598, 205.1437, 203.918, 203.0058, 
    200.1215,
  197.0851, 203.4668, 201.6777, 199.301, 198.8813, 200.8195, 204.9384, 
    196.4906, 203.0505, 207.86, 206.6772, 202.1154, 201.8179, 200.7634, 
    201.6575,
  201.8477, 208.0236, 203.3499, 207.2957, 201.8767, 201.1818, 199.702, 
    202.9147, 203.475, 204.6156, 204.9855, 200.9662, 202.9842, 197.1034, 
    198.6453,
  203.0317, 201.4774, 202.471, 201.8698, 201.1205, 198.2115, 193.5309, 
    200.2123, 202.5489, 207.5608, 201.3658, 199.985, 199.9132, 197.8718, 
    195.7849,
  201.6191, 199.2109, 199.2513, 199.6915, 197.9969, 195.262, 195.3896, 
    194.2996, 197.7719, 197.5937, 198.877, 199.3745, 198.8498, 197.9802, 
    193.4639,
  203.9602, 201.154, 200.3845, 202.477, 200.2919, 196.2676, 197.3933, 
    191.9687, 192.8766, 194.7937, 198.4357, 199.1927, 197.0148, 195.1748, 
    188.6887,
  206.2727, 201.5273, 205.0945, 198.8967, 198.1327, 192.8392, 192.4631, 
    191.7218, 192.3332, 193.7006, 196.0991, 200.4682, 195.2203, 190.6307, 
    184.0941,
  199.5171, 197.4179, 193.1552, 195.7651, 194.9076, 192.8708, 196.2324, 
    193.4482, 192.9446, 192.7763, 194.7507, 198.1013, 192.28, 187.8305, 
    174.7474,
  185.0881, 179.587, 183.4568, 184.689, 188.4131, 185.7643, 190.2995, 
    195.9391, 191.3693, 194.7953, 195.9634, 192.6451, 185.1119, 180.6057, 
    169.7119,
  189.1532, 199.0325, 189.6304, 182.3546, 175.6521, 174.9652, 174.4733, 
    173.4325, 176.7643, 181.2953, 179.9637, 183.8737, 184.9358, 189.0773, 
    186.827,
  173.6711, 182.6187, 178.3466, 171.832, 173.5172, 175.9695, 171.443, 
    172.7857, 179.2971, 181.3095, 179.9008, 180.8605, 182.4645, 190.0738, 
    185.1553,
  166.3784, 176.1279, 177.085, 171.5612, 165.6576, 172.118, 177.8602, 
    166.6158, 173.0886, 180.61, 186.5015, 180.1453, 181.6271, 185.3178, 
    187.3187,
  167.0392, 166.5454, 171.8719, 167.8862, 176.3772, 174.3398, 181.7343, 
    176.1407, 174.8461, 174.6083, 182.3814, 189.4779, 187.0962, 188.6461, 
    188.9084,
  170.1871, 166.1966, 167.8872, 167.9942, 169.7317, 170.228, 174.3819, 
    184.9376, 189.3236, 181.7934, 185.459, 191.9905, 195.149, 192.3968, 
    189.9054,
  166.9809, 168.3841, 171.9784, 176.9073, 181.7313, 183.3409, 181.9389, 
    193.6015, 192.7685, 186.6442, 191.0166, 197.0186, 191.8262, 194.0912, 
    189.1374,
  190.8308, 187.5918, 191.8385, 192.3919, 197.8343, 194.8331, 199.9394, 
    198.0772, 199.3761, 195.2043, 196.6242, 194.7293, 192.2725, 190.9979, 
    189.8168,
  200.7285, 196.9603, 196.7591, 200.2925, 200.6962, 199.346, 202.9022, 
    203.5256, 202.2992, 195.9187, 192.9168, 193.0513, 193.6865, 191.9198, 
    185.6594,
  191.2745, 191.0385, 189.2875, 183.1393, 182.3921, 186.3139, 190.5548, 
    191.2983, 190.2853, 183.6925, 187.2854, 183.0737, 182.78, 179.1937, 
    179.6217,
  198.6954, 198.9019, 193.6618, 188.0897, 180.5537, 177.6429, 174.0471, 
    173.7123, 175.9299, 175.1497, 171.751, 169.5542, 169.9831, 172.7162, 
    172.1098,
  191.3736, 195.0507, 190.6013, 191.5699, 189.7399, 191.0518, 195.992, 
    194.9349, 190.6955, 191.4325, 191.2973, 188.5169, 185.9338, 180.9052, 
    179.009,
  196.9728, 197.9207, 196.3939, 192.9644, 188.0449, 193.9179, 198.1392, 
    192.3967, 191.8536, 188.9495, 192.8283, 189.5754, 184.6782, 178.8152, 
    181.68,
  182.9255, 198.5889, 198.7511, 197.8758, 191.3747, 190.2848, 205.0328, 
    193.5398, 192.8436, 190.0915, 191.6345, 190.1419, 189.0019, 184.0932, 
    186.4572,
  173.399, 174.3815, 182.5743, 189.3062, 196.3173, 192.4206, 188.4939, 
    206.3878, 199.546, 191.3821, 193.0001, 196.9856, 190.8637, 189.7408, 
    193.3532,
  173.2329, 173.0533, 173.6056, 181.0025, 185.6984, 196.5918, 191.2878, 
    194.3407, 199.8802, 199.5283, 196.4122, 194.704, 192.8439, 195.7807, 
    196.1954,
  206.8889, 200.122, 188.4038, 178.3052, 177.2521, 174.9745, 179.2434, 
    198.0718, 202.068, 191.0545, 196.9013, 197.8477, 196.156, 197.1338, 
    196.1947,
  216.6859, 217.5269, 210.1161, 207.4043, 206.6415, 205.144, 198.3163, 
    200.0006, 202.5024, 195.9793, 192.6263, 195.3279, 197.7153, 197.6788, 
    198.3524,
  209.526, 214.8769, 216.0057, 214.6892, 218.6358, 211.9373, 211.9629, 
    209.0345, 204.6608, 195.5496, 190.0709, 191.355, 190.2866, 188.0936, 
    186.0567,
  211.443, 213.815, 211.9946, 208.5591, 216.6936, 217.5327, 213.9811, 
    205.8303, 200.2417, 195.4962, 195.7987, 192.3038, 191.249, 188.5243, 
    182.4504,
  206.595, 213.6675, 211.847, 211.6419, 213.2375, 212.6455, 205.7096, 
    196.1222, 194.8399, 191.7971, 189.1377, 183.5325, 185.7356, 182.438, 
    178.5729,
  180.0439, 180.5445, 180.3074, 184.7195, 180.0104, 184.2719, 189.6471, 
    187.8432, 190.8158, 191.9866, 192.2198, 192.7216, 191.7106, 190.9876, 
    188.7547,
  193.471, 192.1008, 187.5037, 185.5649, 184.567, 191.2122, 189.9866, 
    188.0821, 191.8379, 191.7738, 192.8606, 192.9734, 193.377, 189.303, 
    187.3243,
  204.4913, 200.3465, 194.2158, 190.5903, 188.3594, 187.2592, 192.3814, 
    188.1735, 189.788, 190.2133, 190.3686, 192.1752, 188.1215, 188.2339, 
    186.2939,
  206.8165, 204.6275, 199.0605, 193.2615, 187.0893, 188.9789, 186.418, 
    193.1604, 194.4234, 189.9918, 187.6513, 189.5129, 186.4167, 187.2093, 
    183.9772,
  202.8523, 206.4774, 204.1592, 197.497, 194.8391, 184.1793, 186.8071, 
    189.9691, 194.8651, 184.6659, 184.889, 188.1406, 183.5092, 184.2552, 
    185.4344,
  202.5473, 208.3004, 214.7621, 212.1723, 203.5574, 193.148, 182.4755, 
    187.5728, 190.7053, 183.8016, 184.6027, 184.4091, 182.5167, 184.4076, 
    184.1376,
  205.4354, 211.0607, 210.4166, 213.0109, 214.5069, 212.521, 206.6057, 
    195.5356, 196.715, 197.3407, 194.2361, 189.9701, 189.4438, 187.1324, 
    188.9443,
  205.7802, 199.2917, 204.6766, 211.1331, 208.801, 210.6762, 207.0723, 
    206.191, 205.3701, 196.9095, 197.3457, 196.3582, 197.7568, 199.5831, 
    198.7907,
  204.8037, 206.6963, 203.3938, 192.8141, 200.2944, 193.9765, 200.2788, 
    193.8431, 192.0547, 192.0992, 199.5014, 195.6145, 195.9186, 196.0623, 
    198.797,
  195.4574, 194.3308, 185.8765, 195.4966, 193.4245, 192.6344, 192.9656, 
    188.5645, 189.9329, 184.2695, 191.2838, 188.42, 189.3435, 189.9725, 
    192.8107,
  194.3575, 194.9478, 190.4254, 189.1392, 182.0735, 181.0458, 179.088, 
    170.1591, 168.9705, 166.0673, 164.2255, 167.4073, 167.7351, 174.0048, 
    174.2676,
  202.3378, 197.1005, 193.7604, 188.5478, 182.9544, 185.2925, 180.5147, 
    178.3773, 175.4833, 172.6473, 165.6229, 168.7782, 170.4633, 171.395, 
    170.4494,
  190.0944, 192.9684, 188.4733, 190.3919, 187.8796, 188.4827, 187.0135, 
    172.5683, 176.9828, 176.397, 175.2886, 172.3458, 172.8163, 173.1509, 
    172.4482,
  182.6933, 183.515, 187.7257, 186.1363, 183.6788, 185.5775, 183.3129, 
    180.6714, 181.6911, 180.947, 183.2011, 181.0525, 176.9923, 175.2939, 
    174.7851,
  187.4331, 183.9528, 188.8189, 188.3152, 187.8625, 178.4524, 181.5308, 
    184.962, 190.7359, 188.6494, 185.921, 189.336, 186.7755, 181.8557, 
    177.9449,
  193.3789, 190.3285, 187.2268, 183.6884, 186.6902, 186.4588, 177.888, 
    182.8923, 184.4246, 180.8839, 189.0917, 190.6247, 189.9738, 187.9718, 
    183.4842,
  199.8055, 202.2712, 198.5254, 197.2434, 190.1997, 187.1487, 186.9246, 
    180.897, 182.9483, 181.7626, 181.9302, 181.2603, 186.4107, 184.9473, 
    183.3737,
  200.9528, 206.1272, 204.6245, 202.6836, 201.8865, 201.7699, 196.4392, 
    201.7543, 189.7981, 182.5363, 179.5485, 181.2569, 182.8735, 184.1633, 
    183.6538,
  209.9834, 209.192, 205.5868, 209.6667, 204.9581, 205.8777, 193.7304, 
    203.0969, 195.9376, 191.137, 195.5746, 181.9213, 179.3828, 179.2018, 
    179.5053,
  210.1353, 209.8971, 206.467, 210.0753, 208.1539, 201.2595, 193.6904, 
    189.6973, 190.9131, 185.5063, 187.9221, 181.465, 180.1774, 179.0254, 
    177.3906,
  193.5452, 194.5109, 194.4209, 194.8378, 189.3527, 188.5192, 185.0185, 
    177.2049, 170.2388, 165.0171, 163.4391, 159.7028, 157.4546, 157.9586, 
    156.0098,
  196.5618, 196.2551, 190.4772, 189.7025, 190.193, 191.6678, 191.5045, 
    188.5996, 179.9248, 177.2753, 174.7106, 168.4868, 164.5108, 159.7905, 
    159.7547,
  194.638, 196.2798, 189.2915, 184.0682, 180.6282, 185.6796, 192.4268, 
    190.882, 188.1469, 183.5108, 183.5476, 180.738, 176.2931, 171.5517, 
    167.0896,
  197.8166, 205.0684, 196.7597, 187.741, 179.4731, 178.6634, 181.7225, 
    188.6986, 191.8822, 191.0407, 188.1704, 186.6345, 182.4889, 175.5088, 
    174.0602,
  198.2188, 203.754, 207.8797, 199.0466, 187.4065, 178.0133, 173.5364, 
    185.1189, 193.6276, 189.2953, 186.4847, 188.0704, 185.9702, 184.8845, 
    180.5852,
  190.6474, 200.7119, 203.4954, 200.5741, 197.2249, 187.7793, 179.3575, 
    177.1801, 178.2027, 177.7739, 187.6695, 192.446, 188.3352, 188.1834, 
    186.3195,
  190.991, 191.8747, 197.2957, 198.2598, 202.4013, 203.6498, 194.6668, 
    184.0837, 181.5137, 181.6653, 185.4124, 188.1271, 188.4719, 190.5362, 
    189.3023,
  182.9642, 183.6981, 192.553, 192.0436, 197.5926, 209.5319, 211.4371, 
    204.1457, 192.6557, 181.7688, 178.3195, 179.3293, 184.0813, 187.4676, 
    189.1676,
  181.8637, 181.5878, 186.6069, 189.5163, 191.5157, 192.807, 204.5025, 
    199.0683, 191.7021, 187.6637, 185.1637, 176.9807, 178.3127, 181.2648, 
    184.2678,
  166.4474, 170.7079, 176.6206, 181.0146, 183.141, 184.1381, 184.3907, 
    184.3234, 183.9118, 178.2811, 180.7632, 175.1425, 175.1821, 175.292, 
    181.507,
  170.9951, 176.3864, 181.1867, 185.6512, 187.2139, 191.1738, 194.9611, 
    191.122, 187.505, 184.2131, 178.6134, 174.2045, 169.144, 166.2398, 
    163.0371,
  168.6696, 172.6027, 176.4006, 181.9088, 183.4083, 194.0686, 194.2991, 
    191.7407, 189.8429, 184.7371, 182.1753, 175.9844, 170.6271, 162.8195, 
    159.3493,
  170.0861, 167.8402, 172.4878, 180.5566, 184.1029, 191.7682, 192.6031, 
    189.0331, 189.2886, 185.713, 183.7565, 176.035, 171.1142, 167.7273, 
    161.4996,
  166.7607, 165.999, 176.0896, 190.1608, 187.3549, 186.8306, 183.4437, 
    183.5415, 185.5007, 187.5394, 184.7824, 179.5435, 172.3, 169.5328, 
    161.6663,
  170.5308, 190.5073, 207.0987, 203.9237, 199.9768, 191.0368, 181.3228, 
    183.2352, 185.1689, 176.2612, 178.5762, 182.6796, 174.7822, 170.7245, 
    163.9557,
  202.1693, 211.6776, 214.5526, 212.8448, 206.7327, 199.584, 189.4709, 
    184.4483, 180.5048, 178, 184.8602, 185.6691, 179.4287, 175.0048, 168.091,
  200.9852, 203.646, 209.6626, 204.4483, 208.6484, 202.9958, 201.3426, 
    194.245, 187.7283, 187.9081, 185.6488, 183.6006, 183.1209, 179.7031, 
    172.7433,
  160.1943, 174.6086, 183.6203, 183.6284, 184.6397, 190.2129, 200.7662, 
    211.206, 196.4279, 185.9926, 182.8776, 181.2562, 182.9316, 182.5243, 
    175.2576,
  155.6238, 165.0574, 173.861, 172.7699, 170.0208, 169.6957, 177.3113, 
    189.6948, 192.4549, 189.8443, 188.7967, 179.0156, 178.7287, 178.8162, 
    178.3978,
  163.821, 169.4422, 177.5611, 179.4589, 180.9984, 173.8019, 171.1379, 
    174.9388, 179.8671, 177.6945, 179.6306, 176.3815, 175.7674, 174.1035, 
    175.8919,
  173.9761, 170.9433, 168.9139, 172.957, 175.3272, 179.322, 183.0667, 
    189.217, 185.5069, 185.7988, 185.6699, 184.8867, 179.6684, 176.6664, 
    170.9432,
  174.564, 173.6158, 171.8421, 171.1468, 170.4611, 178.0225, 179.8922, 
    182.3411, 187.8089, 184.6557, 185.4592, 185.1967, 187.171, 181.7, 174.8967,
  183.4676, 179.2804, 176.2269, 168.7809, 171.0841, 172.8593, 172.8969, 
    175.7671, 184.9691, 189.1648, 185.0255, 185.3833, 185.0972, 184.551, 
    182.834,
  186.1531, 177.9675, 173.6805, 171.3141, 167.4457, 170.1649, 170.0259, 
    179.3563, 183.1828, 188.0283, 189.6531, 189.5164, 186.4077, 185.8473, 
    186.4215,
  178.619, 177.5958, 180.317, 187.3125, 188.1865, 183.7229, 183.1345, 
    187.4137, 190.4119, 187.9588, 189.8352, 192.7536, 189.4966, 188.4555, 
    187.3902,
  199.5958, 201.1477, 190.7292, 194.8851, 199.9876, 203.4756, 204.4056, 
    199.7377, 193.213, 186.0859, 189.7494, 191.9109, 190.5634, 190.6514, 
    188.3796,
  210.6659, 206.0981, 203.2759, 195.1476, 207.3604, 210.9804, 210.9209, 
    206.4044, 199.7215, 194.1551, 191.4779, 187.4481, 187.6948, 189.1311, 
    189.8216,
  180.3836, 184.0511, 189.2475, 195.7267, 198.7722, 200.1316, 191.5031, 
    192.2018, 193.7549, 191.7028, 186.2061, 184.3755, 182.5902, 182.9866, 
    185.2204,
  150.3053, 162.5483, 167.1646, 185.9125, 204.6383, 200.6617, 195.9242, 
    180.7821, 174.244, 179.1723, 182.3572, 180.572, 179.3466, 178.5072, 
    180.5997,
  163.1222, 172.2766, 179.1166, 201.5027, 198.384, 191.527, 186.8879, 
    176.4588, 168.822, 166.4916, 170.5522, 173.9369, 174.6774, 176.5042, 
    178.8535,
  187.468, 181.3252, 172.3279, 168.9456, 160.2596, 163.448, 167.8819, 
    173.3927, 177.1664, 183.6606, 185.9617, 185.8512, 176.9566, 171.7944, 
    168.3595,
  193.7198, 183.6902, 175.3087, 166.9447, 163.35, 162.7152, 167.5466, 
    170.8436, 175.2939, 179.5694, 185.5204, 187.096, 181.8233, 171.1909, 
    165.1284,
  196.6339, 186.1681, 181.7159, 173.2963, 168.3845, 167.7318, 165.2634, 
    169.2686, 173.7506, 176.729, 182.3, 187.5475, 179.7592, 176.4331, 166.4301,
  168.202, 168.3641, 172.8048, 177.9468, 173.3377, 169.6723, 165.2095, 
    168.5098, 174.1797, 175.0671, 181.1294, 185.349, 181.2084, 177.8092, 
    170.0101,
  163.0762, 161.8517, 167.2612, 170.3604, 172.2222, 166.6529, 171.7621, 
    172.5753, 178.0899, 172.6945, 177.1248, 183.6295, 183.9717, 180.6315, 
    173.417,
  192.039, 195.2359, 193.7854, 191.7515, 189.8394, 181.5246, 172.2704, 
    171.6801, 170.1765, 171.392, 179.4952, 184.5881, 183.3146, 180.0867, 
    177.9488,
  210.4074, 212.4534, 214.7941, 210.1601, 210.8736, 207.0144, 198.7915, 
    186.2612, 183.5438, 183.6883, 183.4155, 182.0804, 183.2549, 179.251, 
    177.5217,
  210.9323, 213.7947, 210.1346, 217.4707, 212.4225, 208.8701, 206.8582, 
    205.6968, 200.1453, 193.5967, 188.8528, 185.6625, 182.6559, 181.0528, 
    177.6094,
  210.9656, 214.3378, 215.7994, 218.0444, 215.4727, 209.5173, 207.1434, 
    201.1929, 195.6868, 194.1513, 192.9025, 187.7963, 181.4904, 180.4565, 
    177.8231,
  213.0766, 215.8465, 209.6788, 206.5231, 195.3648, 188.2145, 186.845, 
    190.1488, 187.0994, 188.0965, 189.8602, 187.2382, 180.9689, 179.5878, 
    174.4476,
  194.8555, 203.0503, 199.8906, 196.3454, 186.9354, 182.1518, 178.0423, 
    177.3517, 181.8477, 183.6989, 188.7491, 188.8363, 188.9824, 191.0364, 
    192.3882,
  196.3372, 192.9512, 194.0932, 193.8326, 185.267, 189.9087, 183.5253, 
    176.138, 178.3382, 182.9104, 185.6692, 189.8785, 190.1777, 190.4312, 
    191.1823,
  200.6285, 189.6073, 177.3503, 180.1066, 186.5087, 183.7227, 184.0933, 
    174.4476, 173.7854, 177.7881, 179.8506, 181.8683, 182.4713, 188.8798, 
    187.5495,
  194.4012, 187.5913, 178.5701, 177.685, 181.0848, 182.7728, 177.6051, 
    176.1762, 174.5686, 174.3793, 173.5903, 177.6192, 178.5571, 182.0818, 
    187.7985,
  193.539, 202.0384, 188.5733, 176.36, 170.6141, 177.7761, 176.6167, 
    176.8894, 178.9847, 172.6861, 168.541, 173.189, 177.2877, 180.2678, 
    183.2906,
  202.5933, 221.4307, 207.5448, 179.1573, 167.4173, 166.7058, 167.0955, 
    178.5692, 174.8004, 166.8243, 169.903, 172.562, 176.392, 178.9203, 
    181.3796,
  207.1799, 218.3813, 216.9678, 211.9812, 196.0112, 178.804, 169.547, 
    170.1274, 168.2135, 168.9051, 169.6283, 168.2316, 175.3535, 178.5935, 
    180.6621,
  218.7665, 217.3066, 218.3995, 220.1784, 217.9611, 203.0164, 181.0711, 
    177.4723, 175.6505, 169.9225, 166.9185, 166.3647, 172.3534, 175.1233, 
    179.606,
  214.1981, 220.6456, 217.2378, 219.9272, 213.1797, 207.0127, 195.5802, 
    184.1027, 173.0745, 169.0316, 167.5521, 167.5885, 170.2878, 175.9214, 
    180.9459,
  208.1366, 216.3656, 213.8476, 204.0291, 192.4827, 187.0121, 185.0988, 
    183.6396, 176.2014, 169.5215, 168.7293, 171.3245, 172.4548, 177.1901, 
    180.09,
  191.7419, 186.2571, 181.7882, 176.3015, 168.4169, 165.7953, 170.0126, 
    171.9245, 179.1095, 177.2927, 179.5728, 178.141, 180.0869, 174.1352, 
    174.3478,
  199.9294, 190.6165, 190.694, 179.3701, 167.4408, 170.7471, 168.4906, 
    173.9144, 177.0192, 178.1506, 176.4346, 178.4019, 177.0489, 172.8537, 
    175.1835,
  207.4193, 201.4024, 196.8356, 183.4293, 173.2626, 173.646, 173.6802, 
    170.4439, 173.5949, 174.7541, 177.3581, 173.3667, 173.6102, 169.8268, 
    171.6106,
  211.4085, 204.8984, 207.6392, 201.4775, 183.6618, 177.6876, 174.5361, 
    173.6881, 172.1139, 173.2654, 170.3277, 173.0399, 174.2377, 170.5974, 
    177.0813,
  221.1262, 203.4158, 213.1809, 206.0869, 203.1026, 183.9143, 181.4579, 
    183.6914, 180.903, 175.3434, 173.1759, 171.7834, 173.896, 176.8697, 
    185.0939,
  218.1419, 214.9327, 208.5983, 201.82, 199.5215, 195.8379, 182.5486, 
    180.3153, 177.268, 176.64, 178.7555, 174.6647, 176.0173, 176.9626, 
    183.3093,
  202.8385, 217.3463, 221.135, 203.6904, 195.6653, 194.4474, 195.0909, 
    183.9854, 178.5199, 183.659, 177.2494, 172.7683, 175.1467, 177.544, 
    188.3062,
  201.8344, 218.3994, 214.4901, 212.8411, 201.7678, 202.367, 199.2786, 
    198.752, 187.4089, 181.4128, 177.2801, 176.453, 174.5045, 177.3427, 
    185.2074,
  212.6017, 211.3826, 219.2709, 212.0651, 195.6221, 198.3009, 192.9984, 
    188.498, 186.0993, 184.5359, 182.2274, 180.7241, 176.7597, 178.5473, 
    180.3568,
  217.5199, 211.1701, 207.8267, 202.9643, 190.6611, 186.7148, 186.1938, 
    187.3647, 184.8801, 184.8463, 184.7648, 180.296, 177.424, 174.4404, 
    179.1041,
  194.5956, 174.7085, 167.3259, 165.5976, 161.5631, 157.644, 162.3848, 
    168.7565, 172.8748, 176.6428, 182.8895, 190.4568, 190.6579, 188.6509, 
    185.2728,
  206.8752, 182.0612, 166.9656, 162.2061, 159.4678, 161.727, 171.545, 
    181.6573, 181.8004, 184.8339, 185.8098, 195.2655, 195.5197, 184.9023, 
    178.8348,
  212.3283, 193.1465, 170.6207, 165.8626, 167.5186, 173.1093, 185.3353, 
    187.7108, 186.2874, 186.2487, 191.1878, 191.1426, 185.8855, 183.3801, 
    176.7938,
  215.0081, 199.1404, 183.7034, 174.5121, 173.3729, 181.0314, 180.789, 
    190.2742, 188.021, 184.6603, 189.9133, 186.4931, 181.207, 179.462, 176.014,
  213.0343, 202.5644, 189.2363, 178.8223, 178.0475, 181.2428, 188.7393, 
    184.7093, 185.1888, 182.0691, 184.7321, 184.9735, 179.5699, 178.7897, 
    175.5748,
  215.6955, 207.0263, 191.0228, 182.9282, 177.0388, 181.4142, 179.5642, 
    183.5247, 186.9886, 188.6591, 184.7519, 183.6156, 175.3759, 174.2714, 
    175.8428,
  219.7469, 207.0625, 192.2356, 184.7761, 178.5896, 177.292, 180.9476, 
    180.3098, 180.5456, 181.2554, 177.6621, 175.7739, 170.4616, 169.9967, 
    174.5609,
  220.4991, 210.5155, 201.5868, 188.9492, 179.8327, 173.4744, 177.0154, 
    182.2615, 184.2964, 180.5414, 180.5548, 174.874, 172.1887, 176.5495, 
    180.2452,
  221.1065, 216.2256, 205.2593, 192.8899, 186.6308, 181.1485, 181.497, 
    178.9241, 180.467, 179.4752, 177.1958, 176.2488, 177.3219, 179.9451, 
    185.6373,
  226.3563, 206.924, 206.4135, 194.6553, 185.7991, 180.0376, 179.8206, 
    184.094, 177.9917, 176.4969, 173.26, 175.334, 177.3441, 182.9352, 187.0312,
  171.197, 164.3833, 163.2176, 165.369, 168.5007, 166.8522, 166.8158, 
    180.064, 191.4901, 184.6717, 180.5326, 180.6636, 180.5561, 178.9751, 
    179.4201,
  178.4886, 171.4635, 174.3205, 182.8532, 180.7774, 173.5981, 166.8796, 
    175.5613, 185.8259, 183.2051, 184.4003, 188.4834, 187.3916, 182.808, 
    183.0976,
  180.9193, 181.1993, 184.3194, 190.5679, 189.7545, 176.2382, 172.0868, 
    176.3125, 181.4996, 183.036, 191.8704, 191.9502, 191.1071, 191.5621, 
    187.3787,
  186.2118, 187.6296, 195.0054, 197.5463, 188.1183, 185.3801, 175.9723, 
    179.6839, 180.1144, 186.1001, 192.7164, 193.7829, 193.8223, 192.091, 
    192.5299,
  187.309, 189.405, 200.2723, 201.4403, 202.7877, 189.8524, 192.3743, 
    186.8449, 185.9734, 190.5601, 192.4503, 193.3222, 192.952, 194.1419, 
    189.9418,
  190.4317, 192.2786, 195.1188, 205.4875, 211.1324, 210.3913, 202.7469, 
    203.9469, 201.7585, 200.1782, 194.9493, 194.655, 193.4579, 187.0476, 
    183.845,
  192.8028, 194.3836, 198.5182, 201.6464, 209.7506, 212.0816, 215.4922, 
    202.7339, 201.8455, 201.1452, 195.1731, 192.6686, 188.5477, 181.2259, 
    178.2781,
  202.175, 201.0174, 202.8888, 203.9556, 207.1086, 207.6344, 214.5611, 
    205.5533, 199.4555, 195.9303, 192.3593, 185.4325, 181.1214, 178.2279, 
    179.6075,
  204.1972, 201.444, 202.4429, 196.1664, 201.3338, 200.3114, 203.4073, 
    200.6906, 195.5022, 188.8413, 185.8732, 186.1036, 182.1511, 183.664, 
    182.6333,
  199.1332, 203.9206, 206.866, 201.0634, 201.1615, 199.8278, 199.6554, 
    199.6199, 194.6295, 190.5771, 188.2266, 191.1494, 189.7319, 188.2382, 
    189.9348,
  195.3734, 201.1696, 195.969, 194.183, 190.171, 186.3177, 188.173, 186.4463, 
    193.1582, 188.2651, 186.3093, 193.0541, 189.4306, 181.4644, 166.9055,
  202.832, 201.1681, 200.6843, 197.1251, 189.0069, 182.6447, 178.3502, 
    183.4562, 191.497, 192.4301, 185.638, 188.778, 191.1798, 183.2326, 172.673,
  210.5948, 203.6172, 202.6949, 196.5469, 187.104, 177.097, 181.2694, 
    190.2001, 191.0623, 184.1185, 183.8554, 182.2961, 184.8946, 186.9524, 
    178.201,
  216.2551, 214.6951, 212.6876, 200.5653, 187.4412, 195.7196, 188.1638, 
    189.1957, 186.6345, 180.2565, 179.6396, 179.353, 181.3102, 183.1789, 
    179.8736,
  223.2972, 218.3756, 218.0056, 218.8054, 204.6476, 200.2183, 206.1223, 
    181.4877, 185.3423, 183.5919, 180.0975, 178.5196, 182.405, 183.8219, 
    182.3238,
  225.869, 221.38, 222.2462, 222.1653, 218.8843, 202.9469, 197.0741, 
    203.0045, 197.5186, 194.2743, 184.9138, 181.8285, 182.9055, 182.2076, 
    182.9126,
  223.6087, 223.0316, 218.0009, 218.3619, 218.6912, 217.123, 205.1109, 
    199.2788, 197.2109, 197.152, 189.4112, 185.7605, 180.8535, 181.1551, 
    181.679,
  218.5858, 223.932, 223.6051, 214.9822, 215.3789, 212.845, 201.6196, 
    196.6245, 194.4825, 192.8337, 189.2824, 185.9077, 182.6125, 179.9205, 
    177.6567,
  207.0224, 222.0286, 226.0964, 197.0115, 198.9303, 196.7651, 196.628, 
    195.3004, 189.4705, 184.6161, 182.6182, 183.2798, 181.6389, 175.9881, 
    177.6087,
  186.314, 189.6746, 203.278, 200.6603, 199.2188, 196.2441, 194.7383, 
    194.4484, 186.5339, 180.8766, 178.8728, 181.8847, 178.3757, 177.5099, 
    178.6763,
  199.797, 201.7819, 199.4316, 200.8895, 196.1165, 192.9035, 189.4536, 
    182.3407, 177.5789, 171.15, 169.1264, 170.1316, 173.0433, 176.6358, 
    181.186,
  203.6119, 199.2973, 200.2505, 198.812, 195.7861, 195.1181, 194.6783, 
    186.3874, 184.0848, 180.6742, 177.3438, 174.9862, 178.2787, 176.0164, 
    175.9583,
  208.9002, 204.0729, 201.716, 197.0573, 193.5902, 185.952, 194.1217, 
    193.3698, 192.4736, 188.4555, 182.9837, 182.4489, 178.9464, 178.1537, 
    176.156,
  220.4574, 223.2654, 212.3555, 198.158, 198.8283, 202.355, 187.0896, 
    188.4617, 192.9265, 190.7422, 188.6771, 187.2672, 183.3596, 182.703, 
    178.0122,
  222.1016, 224.0761, 221.6834, 217.5455, 202.2222, 200.153, 201.8595, 
    189.1699, 189.8472, 191.1338, 191.1971, 189.9729, 186.6833, 187.3413, 
    183.0607,
  227.6292, 222.6831, 221.8184, 219.6743, 215.6598, 203.1287, 200.2948, 
    198.2095, 198.244, 199.3667, 193.9574, 195.0437, 191.759, 190.2812, 
    186.5719,
  224.3068, 222.0267, 221.3375, 220.1656, 222.4919, 218.7029, 203.6309, 
    199.7187, 199.4093, 197.5083, 194.3807, 196.8517, 197.3376, 194.0477, 
    189.6871,
  225.8552, 224.6564, 218.4799, 219.8759, 219.9884, 200.3281, 202.2436, 
    202.2102, 195.839, 191.5767, 190.5451, 192.4426, 194.8649, 197.3541, 
    192.9692,
  223.334, 224.3169, 208.2013, 199.5337, 200.817, 201.9631, 200.0153, 
    198.0043, 192.3457, 189.7561, 188.2343, 187.5383, 188.9801, 194.3206, 
    192.9981,
  203.1053, 203.6799, 208.9617, 200.9492, 198.719, 191.9781, 191.088, 
    192.2898, 189.2552, 187.9337, 185.1313, 186.7303, 186.0417, 188.3649, 
    188.6961,
  199.8121, 201.2456, 198.2047, 196.513, 182.3428, 173.0681, 171.733, 
    168.0191, 167.1481, 171.0089, 180.3289, 186.8919, 192.7164, 198.1297, 
    201.4737,
  208.2661, 203.9149, 202.3382, 200.6307, 197.3693, 182.6776, 172.637, 
    170.2557, 167.9324, 173.7899, 181.2374, 188.9809, 194.2839, 199.5469, 
    199.9757,
  210.1265, 212.5956, 206.024, 202.0464, 200.2056, 189.7281, 183.0624, 
    168.1035, 168.7167, 174.0857, 180.7965, 191.2182, 199.8374, 206.9182, 
    203.2074,
  229.635, 211.1904, 214.8066, 205.7059, 205.5246, 203.7896, 183.763, 
    175.4445, 172.0393, 174.9279, 181.5213, 193.0796, 199.5138, 203.4444, 
    203.0802,
  223.354, 227.434, 225.9752, 218.9784, 208.3983, 204.0699, 198.2151, 
    180.0085, 174.3687, 177.1745, 181.4429, 192.5242, 198.1215, 201.2132, 
    200.5358,
  208.81, 218.5958, 218.6597, 216.2645, 212.3411, 205.3796, 201.2736, 
    193.6904, 185.756, 183.2722, 182.8274, 189.1457, 194.7152, 195.2356, 
    196.6314,
  205.7084, 212.4816, 217.0057, 217.8616, 214.6037, 217.3271, 209.3491, 
    196.9566, 188.4582, 187.2294, 189.0522, 189.7774, 192.8277, 192.723, 
    193.8214,
  195.3238, 200.0783, 206.6588, 212.3006, 222.1564, 218.6227, 214.9471, 
    202.8846, 194.357, 191.4544, 192.7924, 192.2323, 191.6218, 190.3697, 
    189.6127,
  189.075, 194.7336, 193.115, 201.9235, 207.8447, 213.6391, 209.8791, 
    200.135, 196.0329, 191.9142, 192.7831, 195.1018, 194.3688, 190.0454, 
    189.6421,
  178.8668, 180.7314, 185.6809, 190.0342, 197.8311, 200.6312, 199.4927, 
    197.7561, 193.0638, 192.6045, 187.9501, 191.295, 190.9037, 193.7319, 
    193.6049,
  199.0569, 202.6416, 199.277, 194.7791, 185.3346, 175.0707, 171.3688, 
    171.6584, 174.5322, 177.4572, 189.0253, 193.4778, 190.882, 193.0443, 
    195.0684,
  206.8937, 205.077, 200.8874, 194.6149, 180.2122, 171.4185, 169.9152, 
    172.961, 177.0396, 180.0327, 189.0543, 196.7174, 197.4431, 194.0473, 
    194.4257,
  222.4707, 215.0526, 204.8285, 192.5821, 180.8043, 171.5994, 171.3153, 
    170.1019, 176.6763, 181.5168, 192.3235, 197.9685, 198.0709, 198.8382, 
    195.4235,
  226.6365, 221.5781, 215.7916, 189.6907, 177.6295, 181.5632, 172.7744, 
    174.0496, 176.5763, 184.6717, 193.5114, 199.5451, 198.4098, 198.5097, 
    195.2724,
  223.2429, 225.3949, 208.2448, 189.2372, 186.0022, 190.324, 187.9747, 
    177.2771, 185.3935, 189.4913, 194.5205, 198.5718, 198.9998, 198.6543, 
    196.3606,
  224.5451, 218.6613, 209.1096, 193.8911, 201.239, 200.9499, 191.5636, 
    193.3966, 191.1359, 197.2668, 197.2737, 198.3937, 197.9803, 198.2065, 
    196.5344,
  218.806, 219.4223, 209.5042, 203.4149, 209.3864, 209.2659, 208.8026, 
    196.7433, 195.7259, 198.5919, 199.0606, 198.4754, 199.0782, 197.8848, 
    197.6537,
  218.2696, 210.7349, 207.4343, 206.2764, 211.2095, 206.555, 211.9616, 
    206.1291, 200.2526, 199.0775, 197.8857, 197.522, 199.1892, 198.3925, 
    199.2221,
  220.0624, 206.8602, 209.8062, 214.4534, 213.5585, 209.8206, 206.3567, 
    200.4602, 199.167, 197.6586, 196.7328, 197.0872, 197.8378, 198.2511, 
    198.9724,
  212.5697, 208.12, 213.0477, 208.5536, 203.7413, 200.0699, 198.3721, 
    199.3784, 196.1056, 194.0419, 193.2001, 195.4277, 196.2104, 195.7525, 
    196.5425,
  181.2627, 178.2878, 176.9413, 179.0678, 175.5317, 175.9386, 178.195, 
    178.299, 179.172, 177.5467, 182.3519, 184.697, 183.0424, 187.611, 188.0748,
  196.9567, 194.4328, 189.652, 184.4459, 177.3373, 180.2624, 176.3796, 
    179.1051, 180.349, 177.9239, 180.5097, 185.9571, 187.0477, 186.1714, 
    189.4426,
  205.0443, 204.0752, 198.2661, 187.9885, 184.65, 180.7037, 178.1223, 
    176.4433, 181.2562, 179.7392, 188.0917, 192.3795, 192.1889, 195.7556, 
    195.5702,
  223.9456, 208.4402, 204.2251, 191.3521, 186.5237, 188.8437, 178.0118, 
    181.3486, 182.5305, 181.7208, 194.5328, 195.7482, 192.0765, 196.0988, 
    196.9969,
  211.8919, 209.3282, 202.9176, 202.0149, 193.0613, 190.1222, 187.3682, 
    179.7259, 189.4698, 191.0343, 191.281, 192.7299, 191.6322, 192.1467, 
    194.6327,
  208.5676, 206.6174, 208.3075, 207.2255, 198.3253, 194.0818, 189.652, 
    192.7358, 200.0106, 198.0837, 191.3377, 187.167, 185.2503, 186.9737, 
    187.9733,
  216.2635, 210.5245, 210.1439, 201.5357, 201.8145, 207.9079, 210.3428, 
    198.8392, 198.8951, 194.5245, 188.2225, 185.0184, 182.9709, 184.1383, 
    186.2497,
  222.84, 214.2724, 213.6237, 210.8629, 212.9106, 215.6727, 199.8415, 
    203.4465, 196.869, 192.2762, 188.9932, 186.6977, 186.403, 185.4148, 
    187.4777,
  219.905, 213.3136, 212.7732, 212.2942, 208.707, 210.271, 202.7314, 
    198.9398, 195.734, 193.5004, 192.6689, 190.953, 190.6144, 192.8928, 
    193.6334,
  210.2898, 211.1845, 206.9639, 202.0292, 200.2443, 199.0959, 197.9139, 
    198.8709, 194.9643, 192.4353, 191.7318, 192.8738, 195.6996, 193.0655, 
    196.021,
  190.5823, 179.0372, 175.1193, 170.6223, 170.2758, 173.5225, 180.9314, 
    181.4496, 179.7045, 179.82, 184.5379, 188.2639, 184.5707, 184.0839, 
    180.5591,
  205.0443, 193.041, 182.8089, 175.7015, 169.7554, 170.1872, 172.0442, 
    174.0654, 175.075, 177.4228, 185.1508, 190.6814, 192.1921, 183.2975, 
    179.2971,
  216.601, 200.7852, 193.1923, 178.6272, 175.181, 168.8753, 169.5983, 
    170.8048, 174.0173, 181.4078, 190.8843, 193.8074, 193.5394, 189.575, 
    187.7067,
  219.83, 222.5122, 205.5247, 188.306, 177.7879, 174.0697, 169.7207, 
    174.4902, 181.0359, 188.866, 194.7044, 193.2266, 190.2288, 190.6588, 
    190.4997,
  217.4789, 215.7915, 209.4003, 190.5259, 187.1957, 182.106, 190.4978, 
    182.0506, 184.2387, 187.3728, 187.8996, 186.7023, 185.689, 188.7645, 
    191.8169,
  218.8761, 217.2128, 207.9619, 199.7363, 208.9713, 205.4325, 200.7815, 
    206.5807, 198.0265, 195.7845, 181.3551, 179.0547, 180.2971, 181.6648, 
    185.2359,
  218.4905, 220.1732, 220.014, 216.0909, 215.8223, 216.1573, 212.4034, 
    200.4131, 192.9801, 183.9364, 177.0567, 174.661, 174.8334, 174.5272, 
    178.8994,
  217.5867, 222.0862, 219.9929, 218.8904, 215.1432, 213.892, 200.0455, 
    199.9202, 191.0638, 180.6071, 178.076, 177.2626, 176.0683, 176.9516, 
    176.9903,
  225.112, 218.2671, 221.8647, 207.8023, 202.6807, 199.7385, 198.1108, 
    194.9887, 189.0435, 184.1391, 182.9513, 184.3465, 182.832, 182.7359, 
    183.6455,
  224.7277, 217.4059, 204.74, 202.3323, 200.0887, 197.193, 194.6336, 
    195.6679, 188.8543, 181.8527, 181.0348, 185.6436, 186.0802, 185.8227, 
    187.2318,
  197.8028, 195.5686, 189.9723, 187.6948, 182.1245, 177.9415, 185.4049, 
    186.2199, 184.3384, 179.2358, 179.2672, 183.082, 178.6544, 178.8042, 
    176.1148,
  202.1614, 194.6644, 187.9958, 182.8189, 178.4135, 176.9373, 181.6903, 
    184.4016, 183.9948, 181.8925, 181.5004, 186.3402, 186.1068, 176.4785, 
    176.1016,
  211.9183, 202.3353, 188.3718, 181.1284, 178.2063, 174.9886, 179.9337, 
    184.5225, 180.9304, 185.1603, 187.0117, 187.1946, 180.9445, 180.3874, 
    177.3297,
  213.1831, 206.3433, 191.3357, 186.3673, 173.7928, 179.684, 175.6319, 
    179.218, 178.7881, 183.408, 187.2148, 185.4459, 180.8035, 174.3099, 
    174.8797,
  209.2901, 207.0281, 196.5032, 191.6565, 180.9893, 177.0768, 188.2785, 
    179.8835, 175.6913, 183.5629, 183.5975, 182.0508, 181.4005, 177.5293, 
    173.4691,
  205.2597, 208.6967, 205.8517, 204.2844, 199.1921, 193.8151, 193.2166, 
    202.5582, 195.2455, 191.364, 181.7968, 180.3696, 179.9172, 179.1025, 
    178.3813,
  212.7064, 213.5099, 216.0176, 216.9162, 216.1969, 216.8152, 209.4794, 
    198.4453, 190.7543, 186.0919, 183.5796, 179.0883, 178.6095, 176.9335, 
    175.9675,
  219.3443, 217.9579, 215.1366, 217.6015, 218.9309, 214.914, 210.0468, 
    199.2135, 188.4924, 182.032, 177.3127, 176.8214, 175.2201, 175.783, 
    176.9779,
  223.9405, 221.6421, 216.0594, 217.8581, 201.5609, 200.0446, 199.319, 
    191.8215, 185.1871, 179.1049, 177.4043, 176.2772, 175.8517, 175.0358, 
    176.5871,
  214.4781, 214.0224, 203.6649, 200.6969, 197.0946, 195.6637, 194.2949, 
    190.7038, 184.4178, 176.5382, 174.1634, 178.5075, 178.0492, 179.0451, 
    178.546,
  202.3568, 201.3032, 199.1195, 199.6137, 196.7598, 190.8554, 183.3017, 
    177.2131, 178.025, 177.6407, 174.7542, 176.0531, 174.9778, 179.2719, 
    176.9421,
  203.6206, 201.7196, 200.6154, 197.4436, 191.0792, 183.2524, 175.9746, 
    175.221, 176.2099, 177.7408, 175.8166, 180.8487, 186.4651, 176.7982, 
    176.2988,
  214.2226, 205.4051, 200.3831, 198.4614, 195.6671, 182.9622, 180.097, 
    173.6838, 172.8908, 176.5627, 181.9656, 186.978, 189.0941, 189.6056, 
    179.7652,
  214.3607, 208.2127, 205.2987, 203.8618, 195.7134, 190.8942, 179.423, 
    178.0158, 177.9725, 179.4106, 184.6749, 187.5381, 189.8443, 183.3077, 
    172.9237,
  220.3593, 204.2152, 205.215, 204.9453, 196.9608, 185.1863, 192.1759, 
    176.3766, 169.3092, 177.2884, 183.7947, 186.1604, 185.6435, 177.728, 
    172.5074,
  219.6887, 222.0261, 215.7732, 209.981, 206.1807, 197.5449, 186.2921, 
    197.8071, 191.4539, 188.2041, 182.1609, 182.7903, 180.3931, 176.7356, 
    171.5107,
  213.303, 213.7867, 219.4842, 217.421, 208.0836, 217.5483, 203.8165, 
    192.8837, 188.537, 186.7301, 184.4674, 182.2919, 179.6334, 176.7218, 
    173.5821,
  202.377, 210.3834, 213.5296, 214.613, 215.0053, 215.9208, 208.9186, 
    195.9329, 187.501, 184.1306, 182.5483, 181.298, 178.6775, 177.0682, 
    176.6568,
  187.2005, 193.8458, 207.3526, 207.3667, 211.3207, 203.5164, 196.9201, 
    187.4334, 183.0964, 181.2111, 180.0664, 179.2795, 178.1126, 178.2882, 
    176.6134,
  183.3078, 183.496, 188.4079, 194.6811, 195.7603, 194.6539, 191.4745, 
    186.226, 179.8941, 174.872, 173.5787, 175.6979, 174.5893, 174.4631, 
    174.4561,
  204.2265, 203.9353, 201.111, 198.7422, 192.8348, 190.0801, 191.4442, 
    188.7973, 190.5993, 186.652, 184.7131, 184.3015, 186.156, 182.2953, 
    180.6136,
  204.3822, 203.0076, 199.9568, 195.8763, 188.188, 185.6854, 186.6997, 
    186.6389, 186.5883, 189.7133, 185.9768, 189.3271, 189.514, 174.7497, 
    170.5341,
  207.6176, 205.5175, 200.5558, 196.0251, 193.9175, 179.1741, 184.2713, 
    183.7287, 183.3114, 186.5471, 186.2744, 186.7089, 188.0637, 186.6861, 
    183.1501,
  215.7973, 209.713, 206.266, 201.6098, 196.9098, 200.2535, 174.9546, 
    181.2624, 180.3372, 179.824, 183.2563, 183.7608, 186.0245, 187.0779, 
    183.3072,
  211.8937, 199.1488, 199.8114, 211.7841, 196.2314, 196.942, 199.2883, 
    172.7166, 173.515, 178.7057, 177.9771, 180.2744, 183.221, 185.2679, 
    186.7528,
  219.2129, 201.5728, 197.4408, 203.9528, 205.7403, 199.2395, 195.3326, 
    195.9047, 185.2383, 178.5098, 175.2565, 178.4603, 180.9575, 184.4456, 
    185.3201,
  216.8781, 222.4372, 220.1246, 199.5465, 208.7652, 203.6681, 199.6637, 
    190.8855, 184.9431, 182.2718, 179.3663, 176.5162, 177.6907, 179.113, 
    182.0443,
  215.674, 217.8851, 220.6354, 216.5362, 196.3068, 201.5505, 201.5777, 
    191.3987, 185.1316, 181.1344, 177.5387, 176.5011, 175.058, 175.5397, 
    177.7036,
  220.5876, 215.1028, 218.5635, 212.8132, 201.0471, 202.9637, 195.8556, 
    187.7738, 182.8208, 179.5112, 176.6315, 174.9484, 174.3412, 175.8395, 
    177.9473,
  217.0534, 209.3171, 214.9909, 199.6217, 193.5389, 189.7075, 188.0836, 
    187.2879, 181.653, 175.1739, 173.1258, 175.4195, 175.2219, 176.29, 
    175.7079,
  181.5276, 187.1077, 184.8672, 188.764, 187.318, 184.8295, 190.019, 
    189.6926, 191.3616, 182.8333, 181.0008, 184.31, 183.3081, 179.5677, 
    176.9631,
  196.6148, 198.0101, 195.3923, 192.8048, 185.6138, 181.9079, 185.553, 
    186.0545, 187.1424, 189.9879, 182.2993, 186.6708, 187.7082, 171.7494, 
    168.5622,
  208.8716, 203.6399, 199.3414, 195.1041, 192.1614, 174.9433, 180.7309, 
    182.5345, 182.6243, 185.6282, 186.7291, 186.6688, 187.6447, 186.0008, 
    177.1906,
  215.0587, 206.5278, 205.587, 200.6997, 195.8939, 198.1754, 173.1338, 
    178.755, 182.1991, 180.9707, 183.5453, 185.1673, 186.6604, 185.9279, 
    180.8138,
  224.4995, 201.5605, 200.2026, 202.191, 195.1663, 196.7291, 199.8976, 
    171.2095, 172.8728, 179.36, 180.2621, 182.2935, 184.6636, 185.1378, 
    184.4669,
  222.3416, 201.7448, 203.2927, 199.8149, 199.7574, 195.9923, 195.9765, 
    195.348, 183.953, 180.5874, 178.4831, 180.9002, 182.3045, 183.1053, 
    184.2743,
  219.4342, 219.4457, 202.3115, 200.8956, 197.8514, 197.3494, 194.0029, 
    185.0003, 179.7287, 180.2375, 179.3129, 180.1497, 180.2362, 179.5888, 
    181.9008,
  222.1038, 221.2808, 216.9879, 211.7312, 200.6143, 194.1405, 194.5982, 
    181.9982, 179.2066, 177.8836, 178.6496, 179.2902, 178.5396, 178.9212, 
    181.222,
  220.092, 221.8883, 215.5396, 197.0444, 194.7097, 190.2355, 186.7475, 
    178.5477, 176.328, 176.1364, 177.3678, 178.2763, 178.2287, 178.7737, 
    179.8362,
  219.7522, 218.337, 205.4196, 195.5247, 186.6022, 181.2369, 179.6496, 
    179.1925, 177.9537, 173.7295, 171.9262, 176.0262, 176.6542, 176.6331, 
    178.3445,
  180.7321, 180.2982, 177.2731, 176.7409, 174.4086, 174.2065, 174.4981, 
    176.175, 179.8864, 177.6496, 177.3698, 179.8712, 177.2785, 175.3249, 
    170.7048,
  183.326, 179.5008, 177.3912, 178.6249, 176.1282, 174.8792, 179.7917, 
    180.4505, 182.9612, 186.0388, 179.6237, 184.3382, 185.7749, 171.9733, 
    170.0372,
  199.4625, 191.713, 186.6339, 185.7827, 187.5058, 173.5946, 178.7959, 
    181.2462, 182.55, 184.6491, 185.0254, 185.0801, 186.7584, 186.6923, 
    178.0689,
  212.9232, 206.8423, 203.4625, 200.4789, 195.5, 196.5443, 173.6529, 
    178.4517, 180.9633, 179.3116, 181.7443, 183.9112, 186.4589, 186.7536, 
    182.1709,
  215.7653, 214.059, 204.1934, 197.3044, 194.9107, 197.6663, 199.1387, 
    172.894, 169.7666, 175.2351, 178.6077, 181.7775, 185.1346, 185.5034, 
    185.619,
  217.5457, 214.5767, 202.9972, 201.7875, 198.9015, 196.1884, 197.4584, 
    198.767, 187.5264, 181.8811, 175.6102, 179.6997, 182.5374, 183.7088, 
    184.358,
  220.1148, 218.3965, 215.0846, 212.0027, 211.8445, 203.5704, 194.859, 
    190.6834, 184.9395, 181.6562, 178.7617, 178.1369, 178.305, 179.5213, 
    181.035,
  209.9906, 203.7852, 198.08, 196.3765, 197.485, 203.3499, 198.5914, 
    188.5816, 183.8653, 179.4625, 177.1316, 176.4005, 175.4971, 177.7071, 
    181.2147,
  209.8544, 201.6188, 191.3275, 185.5189, 187.6454, 193.2167, 193.3138, 
    187.1429, 182.5408, 177.6745, 176.2299, 175.2287, 174.8148, 175.5471, 
    177.2943,
  197.9276, 195.7261, 182.787, 181.6879, 184.2368, 186.9417, 188.5193, 
    187.0046, 180.2757, 172.0553, 170.1284, 173.7448, 171.268, 170.6713, 
    171.7303,
  174.1403, 177.652, 169.7721, 166.5591, 158.1076, 161.6245, 163.6142, 
    166.1344, 168.6401, 168.1886, 167.1174, 166.4598, 168.0479, 169.8888, 
    170.1189,
  174.6875, 169.1498, 166.6902, 162.0888, 162.8303, 161.3598, 160.4452, 
    164.0219, 166.8204, 166.7691, 167.7434, 170.1992, 173.5139, 171.2355, 
    170.1209,
  189.7098, 176.4777, 169.0679, 167.0823, 164.4296, 162.8756, 160.8504, 
    165.0672, 166.8017, 169.2475, 174.8855, 177.5492, 180.0211, 182.2953, 
    177.5696,
  207.0546, 192.2872, 190.9906, 180.1647, 172.8395, 172.2541, 163.4881, 
    167.9035, 172.3878, 174.1495, 177.8393, 181.8508, 185.4793, 186.3904, 
    183.8161,
  220.7477, 205.9878, 200.8925, 208.444, 193.4014, 189.1732, 189.8909, 
    170.8614, 168.5211, 173.4047, 177.0094, 182.7612, 185.3516, 186.7373, 
    187.4113,
  223.4205, 211.1638, 208.5799, 208.2674, 202.4673, 196.65, 197.2749, 
    199.0772, 186.8986, 181.353, 176.8004, 181.0265, 182.8509, 184.2948, 
    184.7134,
  205.3863, 221.8398, 223.4176, 213.3462, 208.9752, 204.6768, 198.7218, 
    191.1293, 185.2413, 183.3642, 181.4797, 179.5028, 179.3192, 180.6995, 
    180.7307,
  182.1926, 206.1967, 208.9126, 211.0399, 217.2932, 213.361, 205.0248, 
    190.1253, 185.1965, 182.2708, 179.9452, 178.7614, 176.8527, 177.0379, 
    180.1426,
  191.6264, 191.9969, 199.5299, 201.6374, 212.102, 203.062, 193.7051, 187.31, 
    182.9162, 178.0486, 175.1608, 173.8268, 172.7789, 172.1434, 178.6772,
  205.1578, 202.2347, 197.7755, 198.3329, 191.116, 184.3563, 178.0921, 
    177.284, 172.5321, 169.0066, 169.9273, 170.0058, 171.3513, 170.116, 
    172.4123,
  191.8797, 172.4679, 165.78, 162.128, 161.4488, 168.0554, 169.4108, 173.097, 
    178.2959, 182.2269, 181.7848, 177.8884, 173.0213, 169.1976, 171.8897,
  194.7186, 171.941, 162.9502, 160.5026, 160.5179, 164.1039, 165.4049, 
    168.7602, 173.2535, 178.7719, 180.7983, 176.8419, 175.5257, 170.7876, 
    167.9316,
  208.8365, 177.9945, 163.9677, 160.404, 161.0271, 163.6497, 167.1552, 
    166.1893, 169.1266, 172.8715, 172.0888, 173.6548, 174.9678, 172.8487, 
    173.4129,
  221.286, 207.6732, 174.8444, 169.0141, 163.8445, 161.6085, 167.9532, 
    168.5948, 174.9326, 174.7695, 174.4425, 175.9934, 174.272, 171.6768, 
    168.903,
  215.6852, 222.0273, 190.5289, 181.1621, 170.9537, 174.5095, 177.8293, 
    177.7846, 175.4522, 178.3082, 180.6812, 182.4458, 180.2531, 178.4639, 
    177.3367,
  212.0103, 222.1426, 202.0755, 194.7847, 188.3327, 184.0757, 187.7715, 
    193.0453, 185.0636, 181.2436, 180.1984, 183.5699, 183.7933, 180.7124, 
    178.0194,
  194.1331, 222.1178, 211.9075, 207.2153, 202.4243, 201.5385, 196.8145, 
    191.7554, 187.4535, 186.0908, 183.0766, 182.7047, 183.4109, 184.9086, 
    182.7532,
  199.9136, 214.1159, 211.2629, 205.8051, 207.4335, 205.9065, 204.5709, 
    196.3447, 195.386, 190.2249, 184.9384, 182.2933, 180.491, 179.8389, 
    185.228,
  203.151, 207.7253, 182.7829, 187.4811, 185.6253, 196.5609, 196.4506, 
    194.1934, 192.6182, 190.8574, 187.6796, 182.9501, 178.4992, 176.2565, 
    177.8235,
  194.2058, 183.5125, 174.7105, 173.3927, 178.038, 184.2901, 187.7076, 
    188.7746, 187.6971, 184.7359, 187.0724, 181.7457, 174.6925, 170.1038, 
    169.5671,
  201.6525, 201.8776, 195.3951, 186.5685, 188.6191, 190.4816, 194.8047, 
    194.9406, 192.3328, 190.1147, 192.7289, 200.7106, 204.5211, 208.4085, 
    197.5681,
  201.6096, 201.0307, 197.2174, 186.3891, 184.9546, 184.3486, 183.5989, 
    186.6424, 184.5232, 189.3092, 189.6463, 194.2046, 198.2745, 202.8293, 
    204.3876,
  202.8183, 202.6517, 199.4008, 187.7103, 182.0743, 179.1118, 180.3832, 
    181.2365, 183.2868, 183.7384, 184.5596, 186.5099, 190.2519, 196.1053, 
    196.9893,
  204.7243, 212.0728, 205.2871, 193.9684, 179.3449, 179.0198, 174.2656, 
    178.2351, 180.0626, 180.2428, 180.8884, 178.7112, 180.9897, 185.8235, 
    190.2125,
  201.2288, 208.1985, 206.4192, 197.8872, 180.7469, 176.5979, 180.0667, 
    178.0385, 177.8094, 179.615, 185.4983, 185.9868, 182.2399, 176.5291, 
    177.9191,
  198.4319, 204.9152, 204.819, 198.2235, 179.0267, 172.8015, 180.3136, 
    187.6078, 187.7601, 188.3226, 186.6101, 191.2196, 192.4153, 185.358, 
    174.9696,
  196.3313, 207.4481, 212.594, 192.8587, 180.3057, 177.6377, 186.9452, 
    193.6792, 195.2596, 194.1264, 188.4051, 186.9734, 189.0879, 192.0139, 
    186.8131,
  205.4941, 214.2446, 219.0854, 184.8709, 178.1594, 183.7851, 194.8868, 
    196.7426, 199.3704, 197.897, 196.3916, 186.4456, 183.6415, 184.906, 
    189.3171,
  212.9934, 215.1125, 202.8448, 189.9155, 188.6364, 194.2937, 195.8987, 
    194.8225, 193.9744, 192.3344, 190.8111, 189.9198, 186.9812, 183.1738, 
    182.9016,
  208.3536, 213.4464, 190.9846, 180.6644, 185.1595, 192.678, 194.8181, 
    194.1691, 190.8195, 188.1794, 190.9153, 188.512, 184.376, 181.656, 
    179.4535,
  192.1277, 190.8304, 194.226, 199.1403, 203.5314, 196.5553, 199.3831, 
    204.1155, 208.5618, 207.1992, 204.5284, 205.5101, 202.1098, 192.3255, 
    185.5832,
  194.411, 191.5038, 189.7686, 200.1048, 202.9639, 191.009, 194.8356, 
    198.2501, 203.9086, 207.1817, 203.7286, 203.4154, 204.2614, 204.5851, 
    203.6009,
  197.9759, 191.067, 186.7546, 194.0473, 203.1536, 192.6702, 190.7614, 
    193.4689, 196.0272, 198.8466, 202.075, 205.8061, 204.0972, 206.0494, 
    206.3428,
  198.4609, 192.2543, 194.154, 197.1667, 205.8589, 205.9644, 189.6186, 
    187.0266, 192.2674, 192.0637, 195.4112, 201.3785, 204.8433, 206.3019, 
    206.0459,
  197.223, 194.2936, 188.3133, 200.1915, 198.3463, 198.2781, 202.3094, 
    185.6572, 180.6397, 180.5973, 187.2497, 193.7769, 200.201, 203.6154, 
    205.2465,
  187.8895, 179.9904, 185.0038, 196.8508, 197.2874, 195.8904, 196.7046, 
    193.2522, 184.1376, 183.5846, 184.2147, 189.0005, 193.0483, 197.8174, 
    202.0299,
  181.8339, 177.4182, 181.6439, 191.5338, 198.2796, 198.658, 192.9967, 
    185.5621, 183.4396, 189.3827, 189.8832, 186.6895, 187.4138, 189.7169, 
    195.6015,
  178.8888, 173.9389, 186.2757, 187.43, 193.2697, 196.6568, 187.0721, 
    183.9836, 185.5888, 188.9262, 193.2211, 186.0089, 183.0291, 185.0291, 
    189.8886,
  177.1645, 176.2365, 185.967, 183.1008, 191.8534, 189.7155, 183.493, 
    180.3344, 184.4435, 188.8566, 192.2835, 186.8151, 182.3428, 183.0292, 
    186.1,
  173.2892, 180.519, 181.6652, 186.0594, 185.4473, 182.1912, 181.6501, 
    182.3462, 182.6513, 188.1457, 190.6801, 188.6739, 181.3195, 180.9385, 
    182.8487,
  186.4416, 182.6546, 177.6624, 176.2234, 178.1267, 176.3343, 178.0038, 
    186.4982, 197.7954, 197.6635, 198.4101, 200.4038, 207.2717, 197.8835, 
    189.271,
  187.1, 182.8798, 178.8649, 175.6482, 177.7782, 174.5121, 177.1832, 
    182.3715, 190.1238, 198.4158, 200.4604, 198.9971, 207.0303, 202.2549, 
    199.2244,
  202.2327, 191.4902, 182.3328, 178.8737, 180.6938, 181.0517, 175.3644, 
    177.5543, 182.7474, 188.8247, 195.1125, 201.4209, 204.2873, 204.7121, 
    199.7551,
  216.7649, 199.4703, 184.3308, 178.284, 177.5201, 181.9483, 180.8586, 
    179.0506, 179.1778, 183.743, 189.3917, 194.0828, 196.9195, 198.7012, 
    198.5348,
  216.4598, 212.0903, 197.9039, 182.6912, 177.7621, 180.2496, 186.1127, 
    188.7821, 192.5664, 179.9433, 183.0609, 187.0788, 192.9522, 194.4037, 
    196.3439,
  208.8405, 210.772, 205.0301, 189.7238, 180.4364, 181.5788, 185.3478, 
    188.9689, 185.581, 184.0758, 180.0471, 184.0789, 187.8509, 190.8141, 
    194.2983,
  192.4556, 195.8193, 198.6141, 194.0206, 183.2027, 185.1877, 180.425, 
    180.1148, 186.5477, 186.2835, 182.4242, 181.1414, 184.3757, 186.8034, 
    192.6277,
  193.2009, 186.3424, 185.5117, 189.6018, 192.0114, 185.6877, 181.7076, 
    182.6563, 181.2923, 184.276, 182.2435, 184.8354, 181.7989, 184.9717, 
    191.6187,
  197.8976, 187.1821, 183.2541, 184.2041, 180.8023, 183.4249, 181.4732, 
    179.5973, 177.922, 180.7039, 179.7657, 185.5637, 180.59, 183.9715, 
    189.6538,
  201.2573, 189.7372, 182.6545, 179.3111, 177.1869, 175.3123, 174.6021, 
    181.0791, 178.284, 174.3518, 178.3907, 182.9357, 179.5763, 181.7564, 
    186.1342,
  209.422, 206.7191, 204.5699, 204.4464, 193.1169, 183.9183, 174.8185, 
    169.5212, 169.8159, 169.4341, 175.1407, 181.3226, 191.8552, 195.8062, 
    201.0238,
  209.5802, 206.1155, 205.8176, 201.3164, 188.5312, 179.5703, 172.4389, 
    166.2462, 171.6452, 170.2886, 177.4569, 179.2085, 189.9144, 191.6799, 
    197.7344,
  210.9085, 206.6048, 206.4819, 199.8777, 189.6939, 176.1031, 170.0983, 
    170.9682, 169.0779, 170.1573, 172.6125, 179.4348, 187.1723, 194.3035, 
    188.793,
  219.2169, 212.1106, 207.1633, 199.3451, 187.2048, 174.6897, 169.1881, 
    169.9559, 169.3503, 171.3316, 171.7424, 178.0132, 183.6144, 188.4992, 
    188.3344,
  223.9728, 222.1454, 213.8666, 198.1226, 182.3363, 171.0794, 167.6697, 
    168.5391, 171.6953, 168.1019, 170.8697, 176.4021, 182.1919, 186.85, 
    190.2881,
  219.9579, 221.693, 215.6719, 201.8702, 179.6665, 174.8329, 169.0797, 
    165.9514, 167.1994, 168.1119, 169.7775, 177.1544, 181.4188, 185.0549, 
    188.9249,
  223.1821, 219.5367, 220.6396, 205.0846, 175.8131, 169.084, 170.0201, 
    169.1106, 170.2573, 170.8611, 173.0435, 177.0536, 179.6823, 183.5549, 
    189.052,
  226.9763, 225.1246, 218.594, 203.1095, 176.895, 169.2182, 169.0666, 
    172.0283, 169.6297, 172.5907, 173.3745, 176.1488, 177.414, 182.8257, 
    189.3158,
  227.4112, 220.5415, 214.9541, 200.3667, 180.3908, 169.5089, 168.3082, 
    168.5568, 169.4378, 170.359, 172.3161, 174.9566, 177.7767, 182.7306, 
    187.3366,
  223.986, 214.3238, 200.2357, 201.898, 189.6801, 175.0623, 167.1596, 
    165.7115, 169.1655, 167.7475, 169.6653, 175.0422, 177.9524, 181.1494, 
    185.0252,
  177.7808, 187.2497, 187.1118, 191.1398, 192.1384, 191.0068, 198.3058, 
    195.1664, 186.5433, 177.2551, 170.7641, 166.6559, 165.8177, 170.7195, 
    175.9651,
  179.9859, 182.7905, 181.7752, 188.4994, 192.274, 188.7237, 193.4153, 
    191.9776, 185.0021, 177.4688, 167.6414, 164.9576, 163.1899, 166.2775, 
    169.1413,
  183.1883, 187.4147, 184.9257, 195.498, 196.5056, 186.8245, 189.8645, 
    186.049, 178.2227, 170.3313, 161.6859, 161.2063, 162.8366, 167.6788, 
    170.1672,
  181.8501, 188.5013, 189.8258, 193.6138, 197.4038, 201.24, 188.7817, 
    182.4833, 178.2656, 168.3593, 163.0038, 159.6824, 159.8563, 164.3938, 
    170.3569,
  183.3203, 190.7544, 195.271, 194.3314, 195.6134, 202.3792, 194.5072, 
    180.3673, 175.1871, 164.1241, 160.6236, 158.9994, 165.4525, 170.1677, 
    175.743,
  185.1218, 196.1248, 205.6074, 198.0473, 205.534, 198.6898, 191.2049, 
    176.4573, 168.2779, 165.5106, 161.9649, 161.4668, 163.4334, 169.2535, 
    179.5417,
  197.0657, 198.9782, 211.1451, 204.6885, 212.4112, 198.0465, 184.8051, 
    173.161, 168.7745, 163.9112, 162.234, 165.4418, 166.9627, 175.0854, 183.64,
  199.4532, 214.2532, 224.0986, 217.8399, 210.2823, 197.8576, 175.9353, 
    173.7687, 167.1243, 165.5179, 164.5124, 167.226, 171.6023, 177.6644, 
    185.5881,
  226.2233, 228.9855, 217.1336, 218.9796, 200.749, 184.5674, 173.0771, 
    170.5001, 167.9747, 167.3706, 168.6726, 168.5701, 173.6382, 181.1239, 
    185.5519,
  230.1905, 226.9771, 221.9065, 212.4043, 196.9157, 174.5933, 170.3761, 
    170.2577, 167.0728, 168.6066, 167.5488, 169.6739, 176.6584, 180.6081, 
    183.6328,
  175.4584, 188.2339, 194.165, 191.8641, 189.4005, 185.4291, 185.6629, 
    190.3109, 189.0249, 188.8349, 186.7469, 187.566, 185.6886, 185.4733, 
    187.384,
  192.2849, 201.02, 199.7946, 192.4526, 188.6829, 188.3526, 187.7222, 
    187.3619, 184.7169, 184.0461, 184.2112, 187.9948, 184.7512, 181.4653, 
    184.0092,
  206.571, 202.4653, 198.9588, 195.8322, 191.0052, 188.9903, 183.3024, 
    183.1047, 182.1681, 183.1865, 186.5293, 185.7953, 182.4896, 179.5032, 
    184.6703,
  209.0897, 208.2248, 200.5569, 196.785, 189.3008, 189.8422, 179.2347, 
    179.648, 179.5033, 183.806, 183.2845, 182.448, 177.4642, 175.709, 174.9501,
  214.6229, 209.321, 202.3601, 196.086, 188.4903, 187.882, 187.8197, 
    182.1058, 177.1012, 180.2513, 180.6781, 179.7039, 172.29, 169.7612, 
    167.969,
  217.5185, 209.9171, 203.8099, 198.2489, 187.6535, 189.2487, 190.4721, 
    195.6792, 187.517, 185.1481, 177.8391, 173.5447, 168.9726, 166.0794, 
    163.6357,
  214.5037, 204.2678, 210.89, 198.2039, 195.2577, 200.0091, 197.0963, 
    190.4293, 186.3372, 180.5367, 173.5459, 167.9129, 161.9869, 159.0444, 
    160.6872,
  219.9657, 217.2604, 209.9165, 209.7764, 216.5612, 208.8831, 189.0681, 
    184.5278, 177.6165, 172.2974, 166.1186, 161.5255, 158.6023, 159.0933, 
    161.6066,
  223.997, 217.6409, 221.048, 211.1664, 210.6879, 186.8392, 178.0889, 
    176.2238, 169.934, 165.7708, 163.102, 160.2863, 160.5039, 159.8845, 
    164.4415,
  218.3812, 218.3553, 215.1566, 204.6494, 192.0743, 177.0975, 173.574, 
    173.0873, 168.036, 164.2487, 163.2917, 160.8365, 161.1642, 166.3965, 
    170.1999,
  206.1765, 204.1543, 204.3807, 203.4323, 201.4415, 197.4061, 195.6129, 
    195.7228, 197.8419, 197.8883, 197.89, 196.7553, 195.676, 190.7888, 
    186.5936,
  209.8355, 208.9012, 206.7326, 202.5564, 200.614, 195.4823, 193.996, 
    192.6768, 194.7986, 193.4258, 191.9444, 191.7768, 189.8136, 182.967, 
    183.5834,
  214.6915, 209.7609, 205.426, 202.7356, 200.6813, 191.8138, 192.539, 
    189.2757, 189.6126, 190.822, 188.3038, 186.5623, 183.9077, 179.2395, 
    179.7404,
  218.7212, 220.2169, 214.6793, 201.7687, 198.9868, 199.4737, 187.6509, 
    188.101, 186.5, 185.8032, 183.6206, 181.2951, 177.0575, 173.9221, 176.1809,
  220.9061, 222.4162, 216.6557, 204.5893, 197.2962, 192.8881, 196.8743, 
    180.1994, 181.2935, 180.0954, 180.1652, 179.7982, 175.6273, 174.9317, 
    176.0736,
  223.675, 220.0511, 212.2786, 206.9741, 200.7177, 191.2416, 189.2952, 
    189.7969, 189.7028, 184.6666, 179.9044, 180.1325, 178.013, 176.1462, 
    179.3594,
  219.4816, 223.6316, 210.7162, 208.3869, 207.2451, 193.9574, 190.4064, 
    187.9931, 189.067, 190.0562, 186.1892, 181.8128, 179.4178, 178.62, 178.763,
  214.8067, 216.2103, 209.4253, 200.4069, 207.2391, 200.3663, 188.8402, 
    186.4552, 186.4579, 187.1601, 185.7038, 179.7189, 176.7205, 175.9194, 
    170.1212,
  210.0465, 208.5195, 211.261, 216.0239, 211.0324, 197.7082, 188.1933, 
    184.471, 183.261, 182.3387, 179.4912, 175.9525, 172.0383, 169.9188, 
    162.4115,
  207.614, 204.1844, 203.0097, 202.194, 194.9243, 192.6925, 188.6157, 
    186.1813, 183.3391, 179.0205, 175.343, 171.6695, 168.2728, 164.1575, 
    162.7574,
  201.2073, 202.5183, 201.5204, 198.6586, 195.8504, 188.038, 188.2944, 
    187.0298, 183.7845, 183.9623, 181.3068, 181.9502, 183.7874, 189.6862, 
    192.218,
  199.9692, 202.4924, 202.799, 199.5121, 194.6779, 187.4271, 187.0413, 
    187.8912, 187.7009, 186.1497, 181.9887, 181.7605, 186.0166, 185.1205, 
    191.6568,
  200.4354, 201.6213, 202.6483, 201.7889, 200.0364, 186.2268, 188.2144, 
    182.816, 185.0643, 186.1322, 186.8597, 185.6998, 188.8878, 193.4686, 
    194.2547,
  200.8542, 206.053, 203.5512, 205.0079, 201.7583, 199.9458, 183.8261, 
    186.1957, 186.6254, 186.2153, 185.6448, 188.6731, 190.611, 194.0893, 
    195.4149,
  191.1793, 197.434, 197.9363, 204.4181, 203.8045, 201.7204, 199.5818, 
    179.2429, 185.9633, 188.7621, 185.8773, 188.2806, 188.8226, 193.2107, 
    192.9886,
  182.2586, 190.9751, 190.9045, 205.6993, 205.6288, 201.0269, 198.7921, 
    196.4053, 193.0249, 188.8237, 187.5978, 187.2474, 188.7806, 189.9819, 
    191.0394,
  178.0202, 188.1959, 185.8291, 200.0192, 210.4141, 206.412, 198.5726, 
    193.8051, 192.5863, 193.897, 192.9697, 190.9809, 190.5922, 190.3668, 
    190.3596,
  176.6122, 173.2716, 184.3507, 194.1424, 209.4889, 210.3278, 198.0795, 
    193.6121, 191.4348, 191.4185, 191.5776, 191.1826, 189.8961, 188.5744, 
    187.314,
  172.5305, 173.5165, 175.6244, 188.4975, 203.2316, 207.0844, 198.3879, 
    193.3186, 190.3197, 188.4564, 188.3522, 188.4422, 188.0485, 187.6564, 
    186.5033,
  177.8272, 176.2357, 173.399, 182.5946, 191.591, 197.7204, 197.2228, 
    195.2343, 189.5217, 184.0423, 184.581, 187.2677, 186.6772, 187.0748, 
    187.3168,
  181.3122, 172.8061, 175.4204, 193.2381, 198.2117, 190.4581, 187.8414, 
    187.625, 184.175, 182.7755, 177.264, 177.2463, 180.3289, 185.4226, 
    185.5235,
  186.893, 176.3516, 174.2383, 191.0622, 196.1385, 189.7611, 189.1045, 
    189.0291, 192.0206, 188.6164, 183.1695, 183.4663, 183.1958, 185.5764, 
    182.7498,
  193.2647, 180.7224, 175.801, 194.7932, 202.445, 188.1396, 189.2165, 
    190.6302, 192.5042, 193.0184, 193.6705, 194.1587, 195.3777, 195.4565, 
    192.5081,
  194.7833, 184.4443, 180.6074, 193.4084, 205.2182, 202.3185, 183.8918, 
    189.8564, 193.1226, 194.3613, 195.9238, 195.6189, 195.2376, 189.8194, 
    183.7461,
  201.882, 189.436, 183.7791, 192.3323, 203.3766, 202.8162, 203.0356, 
    182.4108, 187.7006, 192.4307, 190.4942, 187.1128, 184.0701, 178.5345, 
    170.2016,
  208.1871, 196.4398, 186.9081, 190.8345, 202.4723, 202.2345, 200.6079, 
    198.5957, 192.4594, 192.8505, 190.2271, 185.3691, 180.1289, 177.9322, 
    172.6982,
  213.1001, 200.9404, 191.037, 191.8199, 204.6129, 204.3296, 199.3151, 
    194.3181, 191.3724, 191.6362, 187.8837, 184.0284, 180.4398, 178.8521, 
    172.6735,
  218.4086, 208.4498, 193.8074, 192.4225, 201.4922, 204.8501, 199.4067, 
    194.6616, 190.365, 187.8261, 184.4878, 183.1358, 178.9841, 176.2617, 
    175.5963,
  220.8072, 215.9298, 199.4257, 190.3047, 200.6512, 204.1368, 199.1878, 
    194.3309, 189.7982, 186.0827, 183.9416, 180.2155, 179.814, 176.033, 
    175.1174,
  221.0298, 217.2798, 206.2156, 195.5849, 196.2638, 200.3458, 198.8198, 
    195.8584, 191.1759, 185.5907, 182.4509, 182.831, 180.9373, 176.128, 
    171.7421,
  197.0297, 197.0882, 196.4754, 196.4634, 194.2195, 191.8851, 192.4098, 
    187.0173, 188.7753, 182.5882, 181.9909, 184.0269, 180.5782, 182.2473, 
    176.8518,
  203.4268, 200.7888, 200.6891, 197.3743, 194.2031, 190.4745, 190.1341, 
    189.3991, 189.4162, 189.354, 187.6823, 192.2753, 191.8553, 180.007, 
    178.2256,
  207.3172, 203.0769, 202.243, 200.3921, 199.9882, 186.193, 186.2694, 
    181.1395, 180.5933, 187.536, 191.898, 193.7614, 192.6531, 191.1225, 
    186.1605,
  202.6124, 207.0887, 202.7695, 202.3216, 196.6862, 192.0591, 180.0917, 
    177.7865, 175.2661, 172.8724, 174.5628, 186.5307, 190.4008, 192.744, 
    191.2878,
  200.2502, 202.9844, 203.7359, 199.4717, 194.3445, 191.5145, 188.7687, 
    179.7079, 178.6518, 169.7533, 167.1225, 166.7607, 175.2126, 182.8703, 
    187.5894,
  204.8522, 203.2451, 205.1686, 201.06, 196.5261, 190.1428, 183.562, 
    180.9042, 175.1787, 166.0287, 165.0635, 166.9887, 168.3669, 176.6479, 
    183.7668,
  210.8932, 201.219, 198.6422, 199.5891, 205.577, 192.2598, 182.3307, 
    177.0838, 173.1962, 170.7138, 169.083, 168.8454, 167.1189, 172.1119, 
    176.9921,
  213.2895, 204.9826, 199.4793, 202.0855, 205.2218, 201.1027, 185.571, 
    178.8332, 173.4778, 169.353, 167.2961, 167.2771, 170.7706, 171.6818, 
    177.0555,
  217.6589, 200.3952, 200.8691, 203.2906, 201.9847, 199.1976, 191.696, 
    182.6423, 173.7606, 171.5393, 169.3698, 167.7574, 167.1947, 171.496, 
    171.618,
  206.4963, 201.2977, 206.0458, 201.6467, 199.023, 198.4476, 196.8924, 
    192.9734, 185.5861, 175.7395, 173.5044, 170.1239, 167.4517, 166.7139, 
    169.2438,
  201.4759, 200.1817, 195.9441, 196.1738, 193.3175, 187.3806, 187.5127, 
    183.9977, 183.4039, 181.0211, 181.167, 185.8054, 184.1031, 185.4805, 
    184.5573,
  203.8995, 200.5071, 197.4914, 196.5561, 193.5471, 186.4848, 184.6363, 
    184.5228, 183.0477, 184.0768, 182.1015, 187.7302, 186.4448, 180.5885, 
    180.7119,
  204.7708, 202.5616, 200.3803, 197.3582, 196.9138, 186.485, 184.4082, 
    182.3965, 180.1953, 183.0414, 186.9198, 189.202, 187.601, 183.432, 
    183.1387,
  200.6683, 198.922, 201.869, 196.9793, 194.7055, 197.5726, 180.9105, 182.9, 
    185.2673, 183.6947, 184.9027, 190.0698, 189.6139, 186.2251, 184.8252,
  198.938, 202.1162, 198.2733, 198.4146, 194.9988, 194.2046, 195.6296, 
    181.0363, 183.072, 183.9784, 185.2983, 189.7097, 190.6532, 189.1327, 
    187.0978,
  196.7562, 193.628, 195.1482, 195.252, 192.6156, 191.7914, 190.5706, 
    189.7821, 180.5298, 179.3225, 182.6644, 189.6722, 190.7981, 189.9488, 
    188.1071,
  195.1327, 193.5524, 193.3155, 193.7772, 191.8537, 195.0052, 191.3329, 
    187.0974, 180.95, 177.0147, 180.7363, 188.1722, 189.1324, 190.276, 
    188.6513,
  197.2421, 191.7166, 188.7575, 187.6915, 189.8987, 197.9525, 193.4707, 
    191.082, 184.7734, 176.4439, 172.8731, 177.669, 186.4629, 191.8916, 
    189.4043,
  199.0786, 192.2804, 196.6199, 192.3214, 198.7101, 192.5029, 194.1369, 
    192.9801, 186.6806, 176.2668, 172.0304, 169.8515, 174.4681, 184.3171, 
    190.4321,
  200.2659, 198.6425, 195.4038, 189.2566, 185.3941, 190.8121, 192.4108, 
    196.4297, 191.2801, 178.5928, 171.8651, 169.7597, 167.4496, 170.5181, 
    185.4452,
  199.0611, 199.4225, 197.4025, 196.287, 192.6373, 188.2792, 187.701, 
    189.0852, 189.637, 185.9214, 185.967, 186.5867, 183.3076, 182.0262, 
    181.025,
  202.4155, 199.56, 196.5945, 196.183, 193.8083, 185.5081, 185.4889, 
    187.6519, 188.9164, 188.9794, 185.9666, 188.0868, 189.8028, 182.2522, 
    182.3155,
  202.6139, 200.7874, 197.884, 198.2497, 196.3915, 184.9135, 186.6555, 
    186.6784, 185.0167, 186.8266, 187.883, 187.8035, 188.7741, 190.3358, 
    188.5039,
  203.4902, 202.0183, 201.5873, 198.6306, 199.7358, 198.3315, 183.0619, 
    186.133, 185.4182, 183.9733, 187.4046, 187.998, 187.9147, 188.2047, 
    189.0284,
  207.452, 207.8549, 198.8032, 196.9692, 197.5392, 197.4165, 196.9417, 
    174.4267, 177.2317, 177.9904, 184.3974, 187.3146, 186.3503, 185.8713, 
    186.9243,
  212.359, 209.0754, 196.7191, 200.6569, 196.1291, 192.7539, 188.2559, 
    186.5867, 178.7621, 176.7676, 182.0818, 187.0157, 184.5446, 181.9718, 
    182.88,
  212.1478, 203.5444, 193.4381, 200.6783, 204.4351, 193.9405, 184.4509, 
    180.6897, 173.226, 179.1631, 183.3579, 184.2804, 182.4115, 179.3764, 
    179.2827,
  205.8821, 203.9648, 192.343, 187.6089, 198.9204, 196.6113, 182.2183, 
    177.1127, 172.6557, 176.7033, 181.1505, 181.7618, 183.0107, 179.3501, 
    175.9847,
  206.4869, 190.9883, 190.9433, 215.4908, 204.6474, 191.377, 183.2605, 
    175.6276, 170.1499, 173.4521, 179.647, 181.3096, 178.9855, 178.099, 
    177.0284,
  199.8535, 203.0448, 214.0098, 196.6858, 188.7, 187.745, 184.7324, 179.9863, 
    170.5118, 170.0246, 176.555, 178.3419, 179.6209, 177.9077, 176.6414,
  193.2948, 192.7634, 192.4054, 190.7909, 190.8712, 186.8376, 185.4915, 
    183.5173, 183.675, 181.8976, 184.769, 186.2371, 185.0234, 182.8189, 
    183.0036,
  196.8354, 195.2075, 195.8649, 193.7381, 191.2082, 181.7831, 183.3434, 
    185.2311, 186.2246, 188.952, 187.9117, 189.3583, 188.6323, 185.5763, 
    181.9354,
  209.6112, 197.2912, 195.5608, 197.7439, 196.9061, 180.6879, 183.3094, 
    183.3342, 183.961, 186.861, 190.2815, 190.3096, 188.9301, 187.8184, 
    184.1956,
  221.1894, 214.9953, 209.1069, 196.7916, 197.946, 195.4755, 175.8115, 
    183.6236, 184.9138, 186.8899, 189.506, 189.991, 189.2881, 188.2778, 
    186.6003,
  220.586, 213.2316, 210.7904, 198.0043, 196.3436, 196.7437, 191.9709, 
    170.1113, 173.9652, 173.9815, 180.9515, 185.0806, 186.4129, 189.0219, 
    189.2828,
  222.5867, 208.0061, 214.6861, 204.3337, 199.5179, 193.2449, 182.6477, 
    177.7981, 175.5038, 175.0305, 176.8729, 181.6836, 183.8709, 187.3294, 
    188.6869,
  221.401, 219.9608, 216.8485, 206.6669, 208.0113, 194.1023, 181.7194, 
    176.5427, 172.8514, 177.8433, 180.6012, 180.7043, 182.446, 184.7743, 
    186.7316,
  214.3021, 213.4672, 207.311, 200.2789, 202.4896, 194.2708, 184.7812, 
    180.4762, 177.1483, 179.5835, 182.6301, 182.6967, 182.7803, 184.4209, 
    184.9277,
  216.1685, 199.5396, 199.6585, 206.4742, 194.4012, 186.3305, 184.5944, 
    181.8437, 180.7426, 181.3744, 182.0167, 183.2885, 182.8111, 183.6137, 
    181.6826,
  201.3629, 196.8153, 200.6962, 186.4743, 181.2384, 179.3517, 178.5927, 
    189.9055, 185.1394, 178.1663, 177.4303, 181.3289, 181.7429, 180.9881, 
    179.038,
  192.879, 194.0937, 192.9948, 192.9334, 189.6584, 184.6402, 185.813, 
    186.641, 186.0597, 181.1461, 181.7133, 180.2811, 175.776, 174.5251, 
    172.0895,
  199.289, 197.4346, 196.361, 195.3602, 191.7786, 185.9512, 187.6653, 
    188.3156, 189.7696, 188.0287, 186.4957, 184.9578, 180.7032, 173.1723, 
    170.6459,
  212.4552, 199.5335, 197.6473, 199.2762, 198.6094, 186.8921, 187.6262, 
    186.0432, 186.174, 187.6471, 190.0497, 191.2819, 187.568, 184.2184, 
    179.2484,
  222.8221, 218.8947, 209.5273, 199.1495, 202.2784, 198.0194, 187.8325, 
    190.0295, 186.8657, 186.2764, 189.2319, 191.4931, 191.0041, 190.6934, 
    185.5299,
  223.361, 216.3871, 210.2399, 195.9017, 192.7051, 190.106, 185.0868, 
    176.9468, 179.8392, 181.7688, 182.0802, 187.574, 187.219, 188.8313, 
    188.953,
  216.3437, 205.4845, 201.9131, 192.4739, 184.0405, 179.2755, 171.3549, 
    171.6667, 173.1012, 173.9308, 176.3836, 176.1603, 178.063, 180.9705, 
    184.7526,
  207.2042, 193.0873, 193.0872, 183.6573, 178.8036, 166.9513, 166.9028, 
    164.0345, 168.0555, 171.8047, 173.2953, 173.2836, 173.9452, 175.5051, 
    178.7475,
  195.0806, 183.1454, 180.683, 174.577, 163.3183, 163, 165.399, 167.0688, 
    168.8226, 172.6209, 170.7822, 172.1627, 173.5109, 176.0944, 178.5801,
  187.9074, 176.8064, 174.8991, 165.569, 157.6248, 163.1845, 167.5657, 
    166.7779, 173.0708, 173.8404, 171.5603, 171.0433, 169.3999, 173.1908, 
    176.0987,
  187.9552, 175.3199, 166.391, 160.5803, 160.8388, 168.6614, 172.7126, 
    178.2058, 176.2504, 169.7468, 167.2177, 166.836, 168.4869, 170.3521, 
    176.1474,
  203.4455, 197.5849, 192.9584, 193.5665, 189.4288, 185.9384, 187.0372, 
    183.6749, 183.631, 182.8144, 184.7827, 186.9264, 183.549, 185.0564, 
    182.0269,
  206.648, 204.8944, 203.4356, 202.9545, 199.61, 199.9445, 200.0645, 
    198.4658, 196.2363, 195.2196, 194.1623, 194.0348, 193.5177, 189.5557, 
    187.7598,
  217.0681, 207.5434, 203.1175, 199.9576, 205.9986, 203.3546, 202.3241, 
    193.872, 192.9202, 193.0999, 192.4213, 192.0178, 191.3522, 190.071, 
    188.8286,
  223.676, 203.6582, 189.0004, 186.2558, 192.787, 203.757, 196.8429, 
    193.9371, 185.1943, 180.9124, 182.9126, 185.4368, 183.5237, 183.1749, 
    183.6492,
  208.4018, 179.9112, 171.2866, 175.8804, 177.2888, 182.4454, 189.4646, 
    186.6656, 185.8121, 184.3467, 184.5131, 184.1693, 180.5591, 181.001, 
    179.9336,
  183.0184, 169.1715, 173.4755, 173.3092, 179.8583, 180.4233, 178.3434, 
    180.6593, 184.3298, 184.8082, 187.5794, 188.2508, 184.8733, 183.6202, 
    179.8014,
  170.274, 171.7675, 175.7733, 170.6997, 177.0344, 181.2912, 185.6857, 
    187.7958, 187.5947, 185.3861, 184.7367, 185.5756, 186.4284, 184.7189, 
    181.5467,
  173.6319, 176.1769, 177.1855, 175.9179, 182.8811, 186.0348, 189.2124, 
    187.3512, 185.5414, 183.9594, 183.4015, 183.2119, 183.8963, 184.6433, 
    182.2189,
  177.7234, 175.4656, 177.1894, 181.647, 181.8687, 187.4649, 188.056, 
    187.192, 187.1673, 186.7398, 183.1809, 181.1837, 181.2084, 180.6428, 
    179.245,
  178.9196, 178.324, 180.9008, 180.6722, 184.2582, 187.9392, 185.4897, 
    191.869, 189.8582, 182.1712, 181.8752, 179.8845, 177.0288, 177.6187, 
    176.0389,
  203.698, 204.7941, 204.752, 203.2768, 206.3322, 206.9298, 207.7653, 
    204.0455, 201.6803, 195.7861, 195.3962, 193.8073, 188.1258, 186.4405, 
    177.3138,
  203.4373, 205.192, 204.5062, 203.2435, 205.7351, 201.7262, 205.4418, 
    201.8218, 200.7231, 198.5527, 196.4328, 196.3096, 196.5216, 194.3336, 
    193.431,
  218.5046, 210.4923, 205.9746, 204.2568, 206.6875, 202.0924, 204.0591, 
    198.25, 197.4817, 195.1077, 194.2413, 194.9966, 195.0462, 194.0471, 
    192.7638,
  227.6316, 220.5382, 202.3081, 193.9413, 193.3715, 200.5331, 192.475, 
    195.8553, 192.2943, 188.7582, 190.9691, 192.7808, 192.1539, 191.5059, 
    191.9608,
  220.9264, 202.1477, 186.1066, 184.0643, 183.4674, 191.7728, 197.6772, 
    186.1227, 186.8082, 190.0055, 190.7211, 190.3591, 189.3017, 190.0123, 
    189.8422,
  204.0083, 186.8368, 181.3364, 181.3769, 188.9064, 192.007, 193.4688, 
    189.7762, 187.376, 183.7859, 186.2677, 188.3793, 188.3247, 188.5132, 
    187.8925,
  179.8406, 178.8681, 181.5255, 188.7315, 201.4154, 194.9526, 188.5332, 
    185.9574, 184.3379, 182.9764, 182.681, 183.332, 183.9682, 184.1818, 
    184.7243,
  178.0218, 182.391, 189.9794, 200.5109, 207.6874, 194.062, 187.4719, 
    185.5172, 184.6647, 183.5055, 182.519, 182.5199, 182.3783, 182.0706, 
    182.6985,
  180.7932, 177.6302, 193.5374, 209.7236, 198.4612, 190.4696, 187.313, 
    187.254, 187.6267, 187.8567, 182.6129, 180.6252, 182.4954, 183.6318, 
    182.2022,
  174.6005, 189.5168, 197.4576, 195.4514, 190.3929, 188.4501, 186.9479, 
    192.3763, 191.6478, 182.5442, 182.0813, 180.523, 181.57, 183.5173, 
    180.1484,
  165.8037, 166.9411, 172.921, 184.2728, 192.664, 197.0789, 203.9912, 
    202.3659, 198.9507, 194.142, 193.5679, 191.6068, 189.2819, 189.4507, 
    187.5408,
  164.7304, 166.2028, 174.0295, 181.1014, 189.4603, 193.2471, 196.6232, 
    197.481, 193.2639, 190.6624, 188.2358, 189.0836, 189.5046, 187.2245, 
    187.7218,
  167.5193, 169.6432, 176.576, 186.6681, 190.7526, 194.0839, 192.1912, 
    185.8013, 188.6205, 189.7124, 189.2587, 188.6663, 188.381, 187.8029, 
    187.3188,
  178.6872, 184.299, 181.2594, 185.6818, 186.1418, 193.5122, 188.2378, 
    187.9797, 188.1214, 188.0338, 189.615, 188.6808, 187.303, 186.3755, 
    185.4943,
  183.3752, 187.004, 185.2288, 187.5147, 183.1965, 185.1993, 194.6394, 
    186.5739, 182.7247, 189.1091, 191.2632, 188.0388, 185.9443, 185.4091, 
    184.9043,
  197.0555, 191.1945, 184.7901, 187.6426, 187.9609, 193.3773, 194.0258, 
    191.4704, 186.824, 182.5341, 182.657, 185.1642, 185.0478, 184.6479, 
    183.6626,
  199.4241, 191.8275, 186.3942, 188.2659, 195.5728, 195.9071, 191.7956, 
    187.5401, 185.3858, 184.2403, 184.9552, 184.5701, 184.4661, 183.3748, 
    182.6577,
  187.2778, 181.7834, 192.2384, 195.9761, 203.1218, 193.6956, 189.1349, 
    186.5941, 187.1024, 186.1955, 185.3904, 183.8513, 182.2661, 181.1439, 
    182.0542,
  173.9458, 177.8582, 185.6353, 198.838, 195.1174, 190.134, 187.631, 
    188.6525, 190.2169, 189.4721, 183.1472, 180.1629, 180.1477, 180.8486, 
    179.4622,
  172.8392, 170.4421, 183.7975, 186.4865, 184.4824, 185.8975, 186.0195, 
    192.2196, 193.24, 182.9839, 180.2023, 176.2758, 176.527, 176.636, 174.2554,
  175.9724, 170.1823, 169.0076, 172.0991, 172.5313, 177.8594, 172.755, 
    176.9474, 181.1617, 182.3493, 182.3746, 187.3828, 186.8717, 185.4085, 
    186.4053,
  170.935, 175.1809, 171.5361, 174.6407, 169.4853, 171.1913, 172.5718, 
    174.3307, 176.6905, 178.5474, 181.2594, 184.1145, 182.533, 185.2641, 
    183.9534,
  172.2829, 170.6905, 176.0199, 171.0109, 173.5424, 171.7806, 169.7609, 
    166.1398, 173.3748, 179.324, 178.5391, 180.6191, 180.0367, 180.9823, 
    184.8625,
  178.4072, 173.7473, 173.1023, 177.9476, 170.7591, 171.1565, 169.3613, 
    171.5146, 172.7391, 177.1159, 177.903, 180.8407, 179.1794, 177.7621, 
    180.4059,
  188.6908, 179.7524, 170.0943, 166.9552, 167.8453, 167.9778, 167.7243, 
    170.2038, 174.8921, 172.3541, 175.1221, 179.6303, 180.4308, 177.9227, 
    179.1429,
  203.6853, 187.6783, 177.6452, 166.02, 168.9252, 171.3779, 172.0182, 
    171.3037, 176.3115, 176.9317, 177.3873, 179.0479, 177.6431, 179.4252, 
    179.272,
  206.6603, 202.5974, 187.1301, 176.4722, 171.3234, 168.0705, 168.117, 
    166.9624, 171.0743, 173.3039, 173.2609, 174.7323, 178.2703, 182.5717, 
    181.2728,
  194.3049, 193.6693, 190.8722, 176.3098, 169.5545, 170.7807, 172.5495, 
    172.2711, 172.5486, 175.4115, 177.7385, 180.4432, 182.7721, 181.438, 
    179.7469,
  195.3456, 190.9581, 181.1118, 181.37, 175.5643, 176.3934, 172.2247, 
    172.7838, 178.1026, 182.2856, 182.4391, 182.4893, 180.5638, 178.9189, 
    175.2539,
  179.2244, 175.1221, 171.8582, 175.7705, 173.2271, 177.939, 178.6609, 
    183.9888, 187.2278, 182.9587, 178.052, 177.2991, 176.3703, 173.7308, 
    169.6646,
  195.0473, 193.8904, 192.1766, 195.2281, 197.0502, 201.212, 203.3583, 
    204.8846, 201.4613, 191.9978, 184.7503, 182.6694, 178.1173, 174.2206, 
    173.7825,
  197.6055, 194.53, 188.3891, 188.2334, 186.9963, 194.246, 195.8322, 
    196.5314, 197.2489, 190.3758, 186.8757, 181.9993, 180.8324, 177.702, 
    174.7088,
  203.899, 195.601, 188.1731, 177.2586, 180.033, 180.5697, 188.3338, 
    189.6632, 190.5788, 189.5828, 188.7641, 183.0281, 175.9838, 178.8563, 
    175.1958,
  204.931, 202.1861, 172.4725, 169.0663, 170.0751, 170.3818, 171.7466, 
    181.5319, 185.3092, 188.1175, 186.0085, 181.4956, 176.9446, 178.6691, 
    170.5425,
  205.7077, 210.0772, 175.1592, 164.5215, 165.8003, 169.2233, 172.9726, 
    180.127, 184.6207, 180.6509, 182.3663, 179.3003, 177.9847, 180.2404, 
    173.3096,
  202.1619, 198.7329, 177.0881, 165.7779, 167.589, 166.1295, 170.5104, 
    173.75, 174.0217, 174.2319, 177.6499, 176.285, 181.1286, 176.2346, 
    175.4601,
  196.8982, 205.5072, 183.2338, 161.1537, 165.2906, 164.9489, 171.1175, 
    173.1415, 175.664, 178.4346, 177.3499, 179.1379, 180.8688, 178.4733, 
    177.9778,
  185.8076, 192.8932, 185.6583, 173.1818, 164.8153, 167.8316, 173.1913, 
    174.9047, 181.3646, 180.6768, 181.1641, 180.7062, 181.7431, 180.1363, 
    178.8606,
  182.7444, 180.8779, 181.2178, 174.9573, 167.2835, 167.732, 170.8304, 
    174.3061, 179.7703, 181.7611, 184.0684, 183.6026, 183.0338, 181.2152, 
    178.9916,
  195.2567, 189.8289, 187.3477, 179.4894, 178.1899, 180.4626, 185.5876, 
    192.9387, 191.5158, 183.0182, 177.9607, 177.6675, 176.4342, 176.405, 
    176.7906,
  211.1582, 201.2314, 192.21, 190.9015, 190.7246, 195.9061, 197.4973, 
    196.9973, 198.211, 195.2218, 191.8974, 188.8972, 181.4788, 180.6371, 
    173.5666,
  198.0408, 191.1052, 190.4038, 193.3737, 193.0758, 192.2793, 192.0026, 
    193.9542, 198.0124, 198.1255, 192.3994, 187.5974, 182.4949, 176.4474, 
    173.2506,
  191.7298, 188.0948, 187.7289, 187.2083, 186.9821, 187.0859, 189.2558, 
    190.1509, 196.141, 199.2657, 197.7272, 188.8804, 184.8727, 177.7821, 
    174.9608,
  192.8403, 189.1593, 188.0968, 182.1205, 181.8763, 186.9468, 184.3866, 
    187.8653, 194.5699, 198.6384, 200.0407, 194.8546, 186.449, 173.0294, 
    169.8802,
  192.7774, 190.848, 191.0492, 183.7603, 182.1624, 181.5578, 184.0132, 
    183.2904, 187.4171, 192.2341, 197.8826, 200.081, 190.4089, 182.2698, 
    170.0603,
  195.0422, 193.0343, 190.6078, 184.5845, 184.4958, 181.9583, 182.3214, 
    178.4117, 174.267, 176.6995, 187.4745, 190.5031, 189.2083, 184.1991, 
    174.0286,
  205.9436, 199.1663, 196.2679, 189.6174, 192.937, 188.2265, 186.0726, 
    181.3143, 176.6483, 174.5353, 173.8455, 179.2177, 182.9965, 181.4037, 
    175.9942,
  201.4093, 203.7824, 195.9498, 198.0084, 197.8262, 188.6454, 188.149, 
    187.7664, 181.6098, 179.3689, 175.9437, 174.156, 175.9268, 176.9624, 
    177.2788,
  202.0795, 196.5435, 196.9605, 208.9071, 196.7721, 191.6227, 191.5574, 
    190.5792, 187.6101, 184.4386, 181.3407, 182.9269, 182.976, 181.9198, 
    180.9646,
  190.207, 194.8529, 202.2791, 195.3906, 191.4731, 189.7639, 189.9741, 
    194.6783, 188.0473, 180.4166, 178.407, 179.7249, 179.5831, 179.8807, 
    179.3984,
  213.2501, 209.2171, 207.3422, 204.8987, 201.1767, 199.6264, 201.6566, 
    201.6128, 198.4798, 196.039, 196.3783, 194.7146, 192.0163, 191.0388, 
    191.632,
  212.4831, 209.8946, 206.8614, 205.2307, 200.3608, 201.0571, 200.091, 
    201.6436, 200.8164, 197.2898, 196.2481, 193.3149, 189.8572, 188.8, 
    190.9027,
  220.4382, 213.8515, 208.3307, 203.4736, 201.0902, 195.8116, 200.8262, 
    198.6904, 196.861, 194.3918, 192.2133, 187.423, 189.311, 190.1357, 
    191.2712,
  215.7072, 216.0476, 210.8148, 199.8289, 196.4942, 198.5416, 190.1566, 
    194.1673, 187.1902, 186.3387, 189.4488, 190.3893, 188.9978, 191.9963, 
    191.295,
  204.0372, 198.5404, 196.0299, 190.2188, 193.0098, 194.7516, 196.4725, 
    181.9566, 181.3638, 186.5569, 185.9071, 188.9048, 190.6958, 191.6147, 
    192.4659,
  189.6338, 182.453, 184.1494, 185.0027, 187.6817, 192.8857, 191.0249, 
    186.7435, 182.6324, 181.2301, 182.4555, 185.2003, 185.3336, 185.1837, 
    182.3287,
  174.3138, 172.8847, 174.3706, 180.3568, 191.3509, 191.3983, 188.4997, 
    179.2331, 176.9433, 176.9189, 178.8563, 178.4296, 179.5502, 180.5643, 
    177.008,
  167.7712, 168.0853, 167.0448, 180.0647, 197.9975, 190.9579, 187.7836, 
    182.5043, 178.7821, 175.712, 176.0041, 179.3674, 179.3137, 177.8877, 
    176.733,
  171.9935, 167.8152, 169.0724, 189.3402, 197.3664, 190.4265, 186.2913, 
    181.5532, 177.9054, 174.27, 175.7898, 178.6743, 180.1462, 180.1505, 
    178.7406,
  178.0375, 180.1216, 182.7555, 187.6555, 192.6759, 188.1304, 185.5641, 
    185.3185, 179.1481, 173.5217, 173.4362, 176.764, 178.4381, 179.685, 
    180.6543,
  199.0387, 193.6236, 187.2969, 188.8604, 183.2292, 185.7798, 187.3188, 
    186.5186, 186.0714, 187.3301, 189.0245, 189.2046, 190.3439, 191.1498, 
    188.9473,
  203.1738, 204.786, 201.801, 196.7251, 193.7576, 196.8145, 196.7695, 
    196.9174, 193.2587, 187.7165, 191.8048, 192.2285, 189.329, 187.0855, 
    184.8053,
  206.5806, 203.6965, 205.1178, 202.3385, 198.8382, 198.6575, 198.1588, 
    194.3238, 188.3757, 193.2907, 192.3797, 188.1315, 184.0288, 181.297, 
    180.5675,
  189.3358, 190.7166, 199.4414, 199.6082, 193.7332, 195.5061, 191.271, 
    187.7237, 181.4388, 177.9048, 182.224, 183.6301, 182.8295, 180.8739, 
    180.5563,
  181.7194, 186.1921, 183.5311, 186.195, 185.1217, 184.1566, 180.3755, 
    174.9898, 176.4294, 178.8802, 178.8124, 180.978, 180.6255, 181.9902, 
    181.5706,
  188.8921, 186.7325, 184.5991, 188.3756, 184.19, 180.6051, 178.6224, 
    179.8964, 177.0512, 176.3884, 176.4528, 179.3245, 178.4441, 179.8074, 
    180.2309,
  195.1518, 191.1468, 195.3132, 192.5768, 190.4631, 186.0378, 183.324, 
    182.418, 181.4535, 180.8266, 179.5871, 177.0391, 177.9108, 178.2299, 
    179.0569,
  209.7012, 205.5916, 207.4209, 211.0058, 202.3643, 192.0643, 188.1506, 
    184.7942, 182.9542, 179.8536, 177.5604, 176.5299, 174.3839, 175.8665, 
    179.634,
  219.2544, 216.2653, 216.8841, 218.4255, 197.5431, 190.3763, 186.3409, 
    184.1428, 181.094, 178.059, 173.5414, 172.3276, 171.6897, 172.5961, 
    176.4926,
  219.2993, 215.562, 214.0694, 195.5348, 188.4339, 186.0586, 183.8237, 
    183.9874, 179.2988, 169.9298, 165.9466, 165.1299, 167.7944, 171.2398, 
    174.7382,
  178.2182, 166.8297, 160.7027, 153.4674, 155.4322, 163.9291, 160.2536, 
    158.9073, 166.2605, 160.9301, 167.7852, 165.0563, 161.882, 161.5674, 
    162.9144,
  180.5569, 171.5549, 163.803, 154.5045, 155.2379, 156.2884, 159.9213, 
    156.7358, 162.505, 161.7787, 163.2202, 159.3796, 166.1694, 163.5486, 
    164.3645,
  199.4822, 184.5964, 172.292, 164.352, 160.7784, 161.4958, 161.4015, 
    161.4873, 165.908, 171.6105, 170.5737, 172.1636, 175.1994, 176.7654, 
    174.5726,
  212.6278, 208.4844, 191.7402, 181.4222, 174.3748, 173.6277, 170.3663, 
    173.4536, 175.6678, 174.8177, 181.8926, 179.2737, 183.4687, 182.8028, 
    182.9862,
  224.0311, 218.3398, 211.1674, 197.2795, 190.4216, 183.5983, 179.8698, 
    177.3942, 175.7668, 174.2644, 176.401, 177.8056, 178.73, 179.8649, 
    182.8785,
  215.3927, 214.7924, 210.6829, 203.9511, 199.3966, 191.459, 189.2414, 
    186.4735, 183.0037, 176.0839, 174.5914, 179.0778, 178.8637, 181.4592, 
    180.5697,
  218.5253, 217.3448, 220.3326, 211.6675, 206.1669, 196.804, 191.7075, 
    186.4072, 181.2953, 179.4017, 180.9735, 179.2766, 181.4333, 182.9627, 
    180.7952,
  216.6057, 209.3589, 209.6937, 222.6092, 213.247, 194.9563, 189.6891, 
    185.6875, 186.4211, 185.4215, 184.958, 184.1588, 182.851, 178.7808, 
    177.597,
  208.4901, 209.4663, 216.1952, 213.335, 202.6828, 196.3709, 193.6952, 
    192.3205, 191.3439, 189.5575, 185.9758, 183.6506, 181.0845, 178.0495, 
    177.1297,
  199.6364, 202.9423, 206.0319, 201.9546, 198.4615, 196.686, 194.6076, 
    195.6183, 194.6519, 193.1623, 191.2477, 185.9193, 184.4211, 179.6944, 
    177.2936,
  194.1591, 181.1367, 172.0923, 171.2469, 176.552, 181.076, 190.97, 197.5056, 
    199.8702, 202.6452, 209.2944, 210.9494, 213.7527, 213.4485, 210.293,
  202.6046, 185.9823, 173.2072, 164.1327, 172.0783, 178.7055, 189.2227, 
    195.5649, 201.2464, 203.4709, 208.127, 208.8851, 211.5907, 208.1851, 
    199.5859,
  215.7741, 201.5038, 177.4872, 166.6345, 166.3657, 177.482, 188.2132, 
    189.1484, 193.8727, 196.5973, 202.4505, 205.4812, 201.9792, 201.2437, 
    197.7358,
  214.0339, 222.7983, 192.7218, 169.0288, 165.5599, 170.4888, 180.7157, 
    187.5244, 190.2094, 191.2971, 196.5643, 199.4426, 198.7287, 193.9961, 
    191.5769,
  212.9358, 224.3389, 224.3921, 179.2794, 169.2904, 162.7445, 173.8094, 
    182.0568, 183.7382, 188.3349, 188.0842, 190.6845, 191.5944, 190.3799, 
    185.0768,
  222.8227, 228.6058, 228.2855, 197.2769, 171.8252, 165.8776, 164.6752, 
    168.4758, 175.9382, 176.6911, 181.5204, 184.7754, 181.6889, 176.8545, 
    171.6719,
  225.7822, 229.8679, 229.37, 210.2406, 188.5528, 172.3337, 165.6993, 
    163.673, 163.594, 168.105, 169.7374, 171.7867, 169.9828, 168.8968, 
    169.2812,
  231.55, 224.1433, 228.3086, 225.289, 211.9072, 182.879, 170.4435, 165.898, 
    168.2, 164.9935, 164.2826, 166.2699, 164.8733, 164.6624, 166.7689,
  199.6974, 200.5402, 210.5565, 216.504, 208.8414, 199.7448, 184.1326, 
    174.1857, 170.9055, 166.1182, 165.9052, 162.68, 164.232, 166.9447, 
    168.8839,
  174.8295, 180.1929, 186.8212, 196.5608, 201.8821, 203.8685, 197.4621, 
    189.3109, 183.1442, 176.8697, 172.9537, 171.3421, 173.1797, 170.6044, 
    174.7805,
  213.3943, 211.0188, 209.8106, 205.2542, 199.4637, 196.1244, 200.7488, 
    200.5236, 205.5908, 209.164, 206.2279, 208.6277, 208.9902, 208.087, 
    205.3328,
  211.3348, 212.9407, 212.2777, 201.3883, 199.6506, 195.8494, 197.2435, 
    199.3678, 206.3926, 205.3555, 206.4072, 208.8449, 210.2839, 204.9085, 
    200.4804,
  207.816, 214.2308, 214.1386, 196.0677, 193.6502, 196.9324, 196.4996, 
    198.7192, 195.8265, 198.4888, 206.9731, 206.5296, 201.096, 197.5857, 
    202.907,
  201.4476, 209.6789, 210.1581, 198.3493, 189.64, 200.0914, 201.4257, 
    199.0836, 204.6582, 199.3187, 202.41, 199.5095, 199.1516, 203.2815, 
    200.6543,
  197.4025, 210.9788, 219.9155, 201.7307, 188.0165, 188.7502, 197.9314, 
    199.4219, 199.4178, 199.8132, 198.3626, 197.0723, 198.3462, 200.0072, 
    193.5888,
  205.236, 206.3557, 216.4872, 208.7458, 186.1536, 185.3303, 200.2878, 
    209.1946, 212.3397, 205.2155, 197.3193, 193.4359, 194.7285, 195.0403, 
    194.5187,
  207.4823, 203.1948, 212.0434, 212.313, 194.3793, 178.4417, 199.9605, 
    205.3541, 209.1207, 200.5322, 194.6513, 191.1769, 189.3453, 190.7569, 
    198.1822,
  199.7153, 200.5174, 204.9835, 216.6579, 210.4037, 180.7445, 186.6101, 
    205.9223, 207.3468, 198.8806, 191.2061, 189.2209, 190.6059, 188.9207, 
    191.0266,
  208.7983, 204.5156, 198.4743, 203.494, 208.0443, 185.3911, 181.9422, 
    196.1265, 199.9092, 194.1629, 187.8185, 188.605, 189.4031, 184.6687, 
    182.8044,
  219.1218, 212.632, 197.1897, 193.1008, 196.8854, 194.7796, 182.118, 
    189.0598, 194.4812, 194.6082, 185.5191, 185.2569, 183.6892, 180.1673, 
    181.5941,
  208.0718, 204.7877, 204.566, 204.7116, 208.1326, 208.3996, 211.7725, 
    209.8576, 209.6265, 206.0723, 207.0475, 209.7203, 207.9582, 206.7722, 
    204.9932,
  209.619, 205.6825, 201.7329, 202.693, 205.8292, 205.6016, 208.8195, 
    209.0456, 210.2549, 210.0824, 211.1898, 213.0058, 211.6291, 208.5515, 
    208.0545,
  217.0508, 209.9206, 206.1893, 200.9323, 200.8872, 203.2345, 206.0262, 
    206.8214, 202.9014, 204.3939, 202.6637, 202.7618, 206.4901, 212.252, 
    211.4451,
  224.3672, 217.2793, 208.4423, 200.3952, 201.7179, 205.6062, 206.1904, 
    207.2212, 210.8163, 200.0648, 208.2181, 208.0514, 209.3984, 207.3916, 
    207.3069,
  227.8171, 223.2836, 209.2769, 201.2048, 200.6972, 203.1085, 208.5849, 
    203.4252, 201.1201, 205.0045, 204.3685, 204.193, 204.4774, 203.9477, 
    199.6736,
  223.7507, 224.9317, 215.4871, 202.7008, 199.3673, 204.8596, 206.9597, 
    208.5152, 204.7622, 206.267, 207.129, 204.944, 203.2952, 200.8884, 
    197.5327,
  231.1694, 228.6056, 211.6748, 205.5956, 201.4745, 202.3161, 206.261, 
    205.6197, 204.3797, 208.3152, 206.6046, 204.35, 201.4628, 197.5344, 
    199.1696,
  228.0051, 228.6351, 210.4856, 206.2624, 197.1462, 203.1544, 206.3222, 
    209.7564, 203.9024, 205.3805, 204.2566, 197.9907, 196.9738, 197.8127, 
    196.8216,
  226.6243, 225.1416, 207.4115, 201.0277, 198.3049, 200.2801, 203.538, 
    204.6427, 202.0021, 201.5407, 194.0531, 192.0628, 196.921, 196.0727, 
    194.7483,
  216.1275, 211.541, 209.4997, 202.1971, 195.3384, 196.6133, 201.7483, 
    203.2782, 197.5041, 194.5968, 187.0965, 189.8234, 194.9762, 194.237, 
    194.5707,
  212.7554, 209.0363, 206.345, 207.4999, 201.0371, 189.9817, 195.7953, 
    200.3869, 198.304, 196.6361, 193.1138, 190.9524, 188.1336, 188.8806, 
    188.85,
  214.1119, 210.6345, 208.0863, 208.3615, 201.6016, 189.4483, 195.7154, 
    201.4955, 204.9862, 205.9053, 201.8902, 198.7772, 188.3844, 186.1884, 
    186.0048,
  221.3354, 219.1853, 212.0005, 208.3478, 205.2083, 193.5032, 198.4981, 
    203.8123, 204.369, 205.1214, 203.1876, 197.5854, 195.2955, 191.4626, 
    191.3875,
  220.2373, 224.3329, 221.1955, 212.6879, 206.8779, 202.8046, 199.9542, 
    203.3572, 208.5649, 204.6279, 205.3135, 203.4949, 200.0305, 198.4209, 
    194.7919,
  228.5087, 224.9749, 217.0715, 210.2816, 209.6624, 206.8966, 204.6468, 
    200.539, 196.7863, 202.5739, 203.8413, 202.3376, 199.584, 198.0157, 
    196.784,
  226.2711, 225.8771, 220.3606, 207.7498, 206.7045, 208.2719, 207.0613, 
    207.0934, 203.4849, 199.7535, 198.9431, 195.0328, 191.9884, 191.4076, 
    195.1285,
  217.5674, 216.8417, 210.7618, 205.361, 205.6926, 206.7772, 206.3204, 
    206.0931, 203.9896, 201.6948, 194.6477, 189.2499, 190.877, 194.6115, 
    195.5564,
  211.8767, 209.4527, 205.4894, 205.9373, 204.5796, 208.1367, 205.0865, 
    207.7794, 205.9657, 200.2176, 198.1266, 198.1746, 196.1672, 195.9578, 
    194.8609,
  214.0403, 210.9443, 206.8999, 208.0107, 210.6353, 206.8158, 205.063, 
    205.4282, 200.7779, 199.8127, 199.8721, 199.1441, 195.9562, 194.7191, 
    194.3744,
  228.8564, 222.3906, 212.4321, 206.0623, 207.434, 208.177, 206.4892, 
    206.9784, 199.6552, 199.5403, 198.7971, 196.2323, 194.5379, 193.8303, 
    194.848,
  215.5471, 209.1499, 208.8112, 208.716, 209.4644, 203.847, 202.9343, 
    200.0628, 199.9035, 197.5098, 187.1325, 189.9441, 185.3422, 185.5056, 
    190.1249,
  216.3416, 212.653, 210.5705, 210.3302, 210.916, 203.7504, 201.937, 
    201.4099, 203.2399, 199.3893, 194.0335, 194.8913, 189.7563, 187.4277, 
    185.4675,
  216.7312, 218.0803, 211.0146, 208.5181, 210.7986, 202.9909, 201.1182, 
    199.3856, 198.2915, 197.9816, 199.6577, 199.0695, 194.0194, 190.7962, 
    186.0697,
  218.2061, 220.204, 211.6117, 207.5296, 210.941, 209.7895, 198.0226, 
    196.1036, 198.0318, 197.2924, 197.3533, 198.9275, 200.1714, 196.9312, 
    190.1135,
  221.62, 211.0335, 211.4201, 208.8135, 209.6074, 209.6652, 210.1613, 
    196.1643, 193.8476, 194.565, 194.0393, 196.4375, 199.7336, 201.6197, 
    202.4667,
  221.4311, 216.1398, 210.6107, 204.3162, 208.0443, 209.2128, 207.6523, 
    208.7579, 199.1653, 193.0665, 188.9138, 191.6176, 196.2669, 198.7704, 
    201.7332,
  218.0732, 212.062, 208.6717, 202.1997, 203.511, 203.6211, 203.9602, 
    202.2152, 198.4588, 195.3171, 192.1894, 191.6119, 194.2548, 195.3038, 
    197.1856,
  221.1987, 215.5108, 203.4625, 198.0841, 197.4235, 199.6421, 198.4493, 
    197.5248, 195.7643, 193.7066, 191.3095, 191.6795, 194.2629, 194.8562, 
    194.6285,
  225.3464, 213.949, 198.8759, 192.9439, 189.8621, 193.7694, 195.528, 
    193.7759, 192.0289, 189.4976, 189.8908, 191.951, 192.3676, 193.2744, 
    194.0403,
  223.6054, 211.1112, 192.9374, 181.4897, 183.2927, 187.1367, 189.5041, 
    190.2737, 188.5473, 186.015, 187.2753, 188.2077, 189.6561, 190.7012, 
    193.9523,
  212.2133, 205.2256, 192.7721, 187.8679, 186.8231, 180.5524, 184.3181, 
    184.1715, 190.3115, 191.7207, 195.059, 196.9108, 193.5824, 190.1254, 
    185.3641,
  211.533, 200.1018, 190.0509, 186.1538, 182.4719, 178.5062, 176.1806, 
    181.5015, 183.2261, 190.9818, 193.7166, 196.6217, 199.8784, 194.141, 
    185.2676,
  214.5797, 200.7091, 186.47, 182.3882, 176.5902, 173.7014, 178.0034, 
    176.1788, 179.1993, 187.003, 191.3743, 195.7583, 201.0661, 205.3885, 
    196.4309,
  209.1545, 199.7101, 185.8767, 178.1866, 176.2668, 175.4481, 173.8166, 
    183.5345, 185.1948, 185.921, 189.7041, 191.4144, 196.9365, 201.7066, 
    204.629,
  208.2821, 198.4249, 185.515, 173.5555, 173.5856, 170.5376, 179.9713, 
    180.1263, 186.7032, 191.8896, 188.6237, 189.9659, 192.6326, 197.8952, 
    205.1207,
  200.5361, 188.6194, 182.4129, 175.7142, 174.1931, 174.4957, 182.4632, 
    186.4731, 189.5742, 188.8387, 188.3812, 187.0171, 186.431, 192.9768, 
    199.426,
  199.0151, 190.6845, 176.3589, 180.4333, 181.4479, 181.6985, 186.616, 
    187.87, 187.1064, 186.8554, 188.2296, 183.6629, 186.2708, 188.4037, 
    194.0096,
  198.1408, 191.2324, 183.7275, 186.1592, 190.3747, 190.3676, 192.1319, 
    188.353, 187.6899, 186.853, 181.1378, 181.8391, 185.2498, 186.5178, 
    188.7643,
  192.5396, 192.2507, 189.0368, 195.3477, 196.0856, 196.9217, 195.667, 
    191.262, 188.3313, 185.9518, 183.1693, 179.8451, 178.7339, 182.1161, 
    184.972,
  194.848, 190.7295, 198.6147, 197.2165, 200.8614, 202.3081, 200.6524, 
    196.3179, 191.5833, 187.2022, 183.582, 182.166, 178.1148, 176.9188, 
    181.6923,
  197.2846, 194.5761, 191.2558, 190.2468, 193.7702, 189.1576, 186.0648, 
    190.0979, 191.0205, 192.0688, 188.3593, 186.5598, 180.7483, 183.524, 
    175.7054,
  202.4304, 195.2897, 197.4298, 194.9698, 197.2673, 197.9768, 195.2673, 
    194.2302, 199.0659, 201.1964, 195.5134, 191.9749, 188.952, 181.519, 
    177.6234,
  203.7732, 199.7955, 200.1309, 199.1025, 201.9404, 198.0688, 205.3073, 
    195.0487, 199.3402, 203.2325, 200.7648, 198.0732, 190.2898, 186.0965, 
    179.4433,
  203.6285, 202.5577, 208.4182, 204.8752, 204.9686, 203.6425, 199.9263, 
    207.2116, 206.2802, 203.4082, 201.5924, 198.7379, 191.1424, 184.6605, 
    178.8192,
  206.5583, 207.3851, 206.0751, 207.4439, 205.2591, 202.7963, 200.0316, 
    195.0543, 195.886, 202.9286, 202.8312, 200.434, 190.8804, 179.5663, 
    176.4159,
  214.5717, 215.0639, 216.3566, 211.8743, 210.2412, 203.7949, 197.9631, 
    196.3113, 198.2539, 201.2343, 201.1795, 199.0699, 188.6667, 179.0393, 
    176.5224,
  213.5163, 216.7895, 214.3586, 216.7823, 209.0786, 205.0817, 201.3463, 
    198.7269, 200.3741, 203.1837, 202.3811, 200.1532, 192.4277, 179.6873, 
    187.0616,
  212.8973, 221.2099, 216.8221, 210.9735, 207.4065, 202.8363, 201.8147, 
    200.8392, 199.8789, 199.6657, 203.323, 200.8409, 191.2058, 183.4829, 
    188.3327,
  214.1534, 220.0982, 222.1563, 206.7186, 199.6475, 198.843, 198.6032, 
    199.7347, 199.8641, 200.5332, 198.9181, 198.8029, 190.7596, 183.473, 
    184.945,
  213.8044, 211.3777, 210.5211, 200.9383, 198.9007, 194.9827, 196.4594, 
    199.0672, 198.5957, 197.1857, 196.9198, 195.7628, 189.5258, 183.7056, 
    184.1879,
  206.1548, 203.582, 199.237, 199.7803, 200.0005, 197.1013, 196.2447, 
    197.5419, 197.3537, 197.3311, 200.9644, 199.8562, 196.8916, 197.0014, 
    196.8763,
  207.329, 203.9157, 202.7543, 199.3862, 201.2317, 194.4949, 194.4689, 
    195.1013, 194.5415, 196.9037, 198.9519, 199.9515, 202.2198, 197.5529, 
    193.6774,
  209.5594, 203.1128, 203.6109, 199.4383, 196.6102, 193.6378, 194.8535, 
    190.7597, 189.9143, 195.0948, 196.5919, 198.6909, 202.6289, 202.5037, 
    199.1684,
  214.5667, 204.7808, 202.3993, 197.306, 192.4298, 192.6382, 190.6357, 
    193.1039, 191.9202, 191.9717, 193.2602, 195.3747, 199.1501, 199.6533, 
    195.604,
  211.7811, 205.6503, 201.8193, 197.1502, 189.3844, 190.0387, 186.3022, 
    188.032, 189.8829, 189.1175, 188.2929, 190.8253, 195.5651, 197.698, 
    196.788,
  214.4216, 210.0131, 204.4001, 196.6186, 196.1474, 186.0689, 183.1988, 
    184.4669, 182.9789, 181.4974, 182.6479, 185.3961, 188.5101, 194.8584, 
    197.0494,
  213.9065, 208.7681, 205.6155, 195.6528, 193.3751, 189.314, 181.7205, 
    178.0359, 177.1046, 177.5144, 176.1882, 180.2158, 184.5107, 190.2193, 
    194.222,
  220.9957, 208.9547, 204.901, 199.4306, 195.5174, 188.0972, 183.0656, 
    177.5367, 176.2255, 172.434, 170.1585, 176.7494, 180.4561, 186.3611, 
    191.2219,
  218.1633, 208.6102, 207.6151, 198.7008, 193.8356, 187.373, 185.6059, 
    177.224, 174.4514, 170.1162, 169.9896, 172.8855, 177.3304, 183.2366, 
    190.4272,
  223.7778, 215.2543, 210.106, 204.6001, 200.4198, 196.3541, 189.1289, 
    177.7031, 170.9538, 166.4481, 165.3904, 169.0736, 176.3688, 187.3162, 
    189.5292,
  218.457, 213.6357, 204.8449, 197.8309, 187.9187, 184.757, 181.3617, 
    180.0778, 178.0043, 177.048, 184.5824, 181.501, 184.2949, 187.4601, 
    188.5303,
  221.8527, 217.5675, 208.4344, 197.6563, 193.1593, 185.9685, 183.618, 
    186.394, 183.0071, 176.4501, 177.4987, 180.8488, 181.3767, 183.8595, 
    184.1022,
  222.6816, 217.3574, 211.2475, 203.3899, 195.9711, 190.9698, 193.1258, 
    184.6821, 187.5643, 185.573, 181.5459, 175.9687, 175.3812, 176.9337, 
    179.067,
  222.6954, 218.1121, 214.8636, 206.7818, 199.7225, 199.1097, 192.8848, 
    195.7511, 182.9754, 181.2417, 184.7332, 175.0971, 173.7797, 172.9616, 
    175.1645,
  220.0379, 217.1126, 212.4258, 208.8176, 203.5215, 198.6531, 200.9077, 
    195.0869, 188.4066, 183.4005, 183.4851, 179.3611, 174.385, 170.916, 
    169.6342,
  215.8626, 213.8746, 211.3451, 210.4604, 206.8215, 202.785, 199.4277, 
    197.4801, 199.1716, 191.0664, 186.2673, 179.0843, 175.2523, 170.8303, 
    170.1946,
  217.0978, 214.6438, 209.3944, 210.8036, 208.012, 207.9573, 202.9001, 
    199.1569, 197.6122, 196.7782, 187.0616, 175.055, 172.7682, 168.4105, 
    169.0089,
  215.847, 212.1951, 210.1476, 208.3704, 211.417, 212.6128, 206.8757, 
    204.1805, 201.7312, 194.7747, 192.1855, 183.5382, 173.1461, 174.1658, 
    173.1244,
  219.3597, 215.0205, 213.2372, 208.3396, 210.0701, 211.1068, 209.0224, 
    207.8183, 201.0276, 194.139, 191.9995, 188.158, 184.2609, 178.3119, 
    186.7909,
  213.0065, 211.8813, 209.9911, 205.2364, 207.9617, 209.1562, 210.8573, 
    207.7156, 203.461, 197.8076, 195.2593, 191.7159, 189.3639, 194.1521, 
    196.6223,
  196.4029, 195.1645, 196.5609, 198.2817, 196.3573, 198.8232, 202.3237, 
    209.0046, 208.3223, 208.0555, 205.2662, 195.8904, 188.8705, 181.8445, 
    180.0645,
  197.7905, 196.844, 198.9886, 200.1402, 198.619, 202.0556, 203.4714, 
    208.9283, 212.741, 212.0211, 208.5831, 203.1958, 196.05, 188.4479, 
    178.1522,
  200.058, 204.2479, 200.8297, 196.7487, 195.8763, 201.3071, 200.2836, 
    203.2697, 209.072, 209.5098, 211.2498, 208.1571, 199.8144, 188.9184, 
    183.9104,
  199.6066, 203.6787, 200.6364, 200.4637, 194.6313, 199.5814, 201.3082, 
    207.0554, 211.793, 211.8344, 210.1496, 209.3009, 205.6172, 197.8709, 
    189.4307,
  203.2103, 206.9221, 205.8912, 202.2619, 197.3421, 196.1415, 200.9888, 
    202.9394, 206.6921, 211.2986, 211.9455, 210.0143, 206.571, 200.8557, 
    192.1951,
  209.8967, 207.474, 210.5569, 203.1209, 198.826, 194.0652, 194.9598, 
    202.1948, 206.0505, 207.6728, 211.3174, 212.6407, 211.3831, 204.9645, 
    193.6006,
  213.136, 211.2374, 209.0121, 204.0502, 200.6502, 193.1952, 193.0672, 
    196.4949, 201.2057, 203.3779, 207.7755, 211.5303, 212.587, 204.5272, 
    194.8259,
  215.4139, 216.2408, 211.9557, 205.1126, 198.8703, 197.3013, 194.1188, 
    195.7111, 199.1849, 201.2169, 202.2784, 204.0732, 207.4157, 205.3326, 
    200.4943,
  218.2118, 216.9352, 212.1138, 209.0378, 204.1055, 202.266, 202.6251, 
    193.4316, 195.2101, 196.8082, 194.3491, 199.0003, 200.0642, 201.2089, 
    201.573,
  221.7897, 219.8519, 217.0011, 216.5829, 211.4818, 206.892, 206.0479, 
    198.5188, 193.4124, 189.3858, 187.3519, 187.599, 189.4624, 193.5367, 
    195.3238,
  216.7926, 213.8332, 205.2184, 206.7472, 210.8124, 210.318, 208.3993, 
    208.4629, 210.6305, 208.6828, 204.4284, 205.4417, 206.3105, 206.4479, 
    204.9552,
  220.4058, 214.1216, 210.7044, 208.5252, 210.8151, 209.6501, 207.5516, 
    210.1651, 209.8459, 211.1986, 207.233, 205.1331, 206.9386, 209.3401, 
    209.8332,
  220.3985, 213.9716, 211.7566, 210.1564, 213.2037, 209.4326, 210.3644, 
    208.0206, 210.3341, 211.2057, 209.1116, 207.8623, 209.248, 208.2736, 
    207.9359,
  223.7091, 214.9805, 213.003, 211.2856, 212.8218, 212.8381, 210.6554, 
    210.745, 205.1854, 206.5562, 208.221, 208.2988, 211.0334, 209.8315, 
    207.8105,
  226.3378, 217.177, 209.2332, 213.1065, 216.2366, 215.2259, 216.3056, 
    210.6502, 204.3788, 206.647, 206.0729, 205.8401, 204.856, 206.7969, 
    209.866,
  226.4798, 220.0009, 213.989, 211.2061, 216.858, 215.1722, 213.601, 
    214.5273, 207.8196, 203.6124, 198.9297, 201.9949, 200.4452, 204.582, 
    206.2886,
  225.9594, 223.0263, 215.6621, 212.5823, 215.4574, 215.038, 213.4344, 
    209.7626, 204.2532, 202.2407, 195.868, 195.7097, 196.7017, 199.3414, 
    201.2333,
  225.505, 224.0929, 216.7371, 212.9614, 211.8612, 213.5429, 215.2106, 
    211.4165, 205.5958, 201.0989, 197.4512, 194.7704, 190.8714, 190.6754, 
    192.4685,
  225.9865, 223.2644, 219.2199, 214.3232, 213.3814, 213.0958, 210.0631, 
    212.1428, 205.5016, 198.2262, 200.0027, 196.3768, 194.1566, 187.2321, 
    185.2702,
  227.0634, 224.8689, 220.4396, 214.0284, 211.9955, 209.8365, 208.8968, 
    207.4934, 204.0319, 198.9921, 200.5617, 196.0731, 198.2206, 189.906, 
    186.2291,
  220.071, 219.4794, 220.3395, 220.1436, 218.2979, 213.2864, 209.6923, 
    203.8107, 198.9263, 199.6108, 200.2121, 203.8176, 200.0444, 202.7606, 
    205.4812,
  217.7406, 220.7316, 220.9887, 218.8545, 220.8669, 217.0248, 210.2102, 
    207.0806, 199.7111, 196.6764, 194.913, 197.4435, 200.3299, 199.4066, 
    202.0519,
  218.4594, 221.3238, 220.4727, 217.17, 218.8226, 214.1373, 211.3918, 
    207.2835, 198.1527, 198.9811, 190.7534, 191.4247, 190.7962, 199.8952, 
    199.98,
  218.9471, 220.8519, 219.1813, 216.9957, 214.5393, 215.0333, 210.3262, 
    210.4115, 200.6343, 189.3902, 187.154, 185.6843, 186.9435, 187.3808, 
    192.602,
  219.7728, 219.7081, 220.3507, 216.7067, 214.6262, 212.6523, 206.4096, 
    208.2865, 200.4361, 195.8122, 189.5606, 187.9827, 186.2368, 184.8418, 
    185.1542,
  220.9247, 218.7669, 219.3816, 217.315, 216.1405, 212.6808, 206.8356, 
    204.31, 201.7494, 197.0856, 194.6395, 189.8983, 186.3753, 183.669, 
    188.3913,
  221.7177, 217.9392, 218.3888, 218.5031, 215.8748, 210.4025, 208.2803, 
    205.3403, 201.9966, 200.415, 197.6091, 194.2491, 190.7686, 180.5002, 
    183.7312,
  217.3123, 217.1853, 218.8083, 220.6097, 218.0075, 210.0174, 206.8745, 
    204.2085, 201.1959, 200.2345, 197.3829, 197.2351, 194.2593, 189.0504, 
    184.3907,
  215.2104, 216.1831, 220.1309, 217.4695, 211.8417, 208.0337, 206.196, 
    204.4031, 202.0262, 200.5525, 198.0999, 197.4347, 195.2428, 190.2263, 
    191.4353,
  213.2355, 216.3051, 219.0122, 214.4634, 209.1772, 207.0375, 205.3099, 
    204.9041, 203.467, 198.1636, 196.114, 195.9322, 194.4076, 195.8883, 
    190.4465,
  215.2335, 208.3645, 201.3266, 198.6925, 199.0072, 199.6011, 201.4969, 
    204.8097, 204.6427, 197.5349, 195.6283, 186.9837, 186.9985, 186.0259, 
    180.4599,
  217.3603, 213.493, 202.5242, 200.6092, 200.0308, 200.434, 202.825, 
    204.4924, 204.4557, 200.2719, 198.3348, 191.4603, 186.6669, 181.5771, 
    179.8816,
  215.821, 214.8678, 211.306, 200.3921, 200.2895, 199.2348, 202.964, 
    201.7283, 201.8376, 202.443, 201.3091, 196.7617, 192.7219, 182.3438, 
    177.6754,
  218.3663, 208.7902, 211.1221, 206.0158, 199.9848, 200.429, 197.2842, 
    200.3962, 201.229, 201.5334, 200.8326, 201.5893, 195.1049, 188.5195, 
    179.7115,
  219.976, 212.0107, 208.3357, 206.2702, 204.2569, 199.7269, 199.093, 
    191.6789, 194.2277, 202.5747, 200.9102, 199.5272, 200.9065, 195.5229, 
    181.6685,
  217.0789, 209.3474, 209.9499, 210.0464, 211.3492, 200.1397, 195.3924, 
    196.3568, 195.3001, 193.7145, 193.1521, 196.1303, 198.6066, 197.3197, 
    186.5513,
  222.3401, 210.6646, 211.0123, 214.5823, 212.6977, 201.504, 196.4702, 
    194.362, 192.1089, 193.5618, 193.122, 194.2182, 197.285, 198.5886, 
    192.1245,
  223.358, 216.3478, 215.3778, 214.5775, 207.8474, 200.7023, 193.9998, 
    190.9617, 190.4101, 192.0275, 192.8527, 192.891, 194.5462, 196.7044, 
    195.8192,
  220.6798, 214.4574, 214.2575, 209.7445, 204.9503, 196.8745, 192.6568, 
    188.0518, 188.4822, 190.3315, 192.4523, 191.36, 192.1415, 195.1897, 
    198.216,
  224.1641, 217.0551, 211.9125, 206.8682, 205.6498, 198.3155, 193.6344, 
    190.6457, 186.8003, 186.0973, 189.306, 190.2986, 190.166, 193.1424, 
    196.672,
  217.0179, 210.2047, 204.6968, 201.1018, 197.1081, 192.1364, 194.7336, 
    195.5782, 195.3281, 193.6947, 193.4236, 196.7224, 195.4247, 189.9183, 
    180.1431,
  222.2933, 214.7289, 208.3921, 203.5285, 200.5639, 194.3168, 194.9601, 
    197.3974, 196.5188, 196.1645, 192.574, 195.7799, 197.8837, 194.3323, 
    183.8526,
  227.1446, 217.814, 209.9544, 204.6149, 200.0501, 194.5536, 196.13, 
    194.7704, 197.8677, 196.2254, 195.8864, 195.8721, 198.207, 198.3283, 
    189.1069,
  223.7091, 219.0545, 214.2392, 202.5371, 197.7754, 193.8679, 193.9023, 
    194.9404, 197.6578, 198.1724, 197.1432, 195.9009, 197.1202, 197.9625, 
    193.365,
  226.0545, 218.8793, 217.6709, 205.829, 202.0873, 189.7698, 193.7044, 
    191.8797, 195.2371, 199.7893, 198.8742, 195.9623, 195.0056, 197.1653, 
    197.1971,
  219.3335, 217.2442, 214.152, 207.5696, 203.6239, 191.6731, 184.0571, 
    187.1451, 193.6397, 192.3374, 194.7076, 195.3143, 193.6033, 195.3231, 
    198.6337,
  225.6765, 220.5412, 216.2274, 210.4449, 201.4507, 191.4541, 183.9822, 
    183.4693, 188.5721, 195.2594, 196.4034, 195.161, 194.2971, 193.7922, 
    197.8662,
  225.9279, 225.9148, 219.3999, 209.0611, 199.9612, 190.7173, 186.7796, 
    184.014, 185.7819, 190.7825, 195.3424, 194.914, 193.8841, 192.8434, 
    198.1723,
  227.7605, 227.3548, 219.407, 205.6269, 197.1561, 192.8824, 188.3547, 
    185.1122, 185.8449, 191.1102, 194.63, 193.9539, 192.1663, 192.8227, 
    197.7348,
  223.9086, 219.3437, 213.3834, 204.3581, 199.7119, 195.7428, 191.4281, 
    188.9454, 188.273, 188.8949, 193.4888, 193.0312, 190.8104, 191.6044, 
    195.5551,
  214.292, 210.5614, 206.3547, 204.9767, 203.2164, 202.5379, 198.7492, 
    193.8636, 193.7821, 197.1653, 196.256, 195.2692, 190.7118, 194.0483, 
    203.7074,
  218.5629, 217.1502, 205.9849, 202.2066, 199.7419, 196.9294, 187.0257, 
    183.4448, 189.5481, 193.5505, 195.3689, 195.6459, 195.3059, 195.8556, 
    201.212,
  222.4904, 216.0758, 211.0878, 200.5714, 189.2806, 185.3851, 177.8482, 
    174.6591, 185.2332, 192.7563, 197.0313, 196.7845, 194.4326, 191.5277, 
    198.8253,
  221.6661, 223.4129, 213.7645, 202.3492, 187.0446, 187.0911, 172.8561, 
    172.5467, 186.0879, 193.8457, 197.395, 196.3681, 193.2689, 190.5678, 
    197.1632,
  224.7344, 220.9304, 217.5364, 206.4323, 201.9144, 191.5505, 177.8058, 
    173.6808, 190.2628, 195.8011, 198.4633, 194.8384, 189.3319, 191.9705, 
    195.8727,
  228.0436, 221.0902, 217.8596, 209.9271, 211.9952, 199.7446, 179.0413, 
    173.1769, 185.9013, 195.797, 195.1772, 192.3714, 191.0043, 191.783, 
    197.5726,
  228.9958, 220.3911, 219.4967, 209.5213, 209.7151, 199.8394, 183.9307, 
    176.221, 181.7747, 196.5654, 194.8925, 191.3582, 190.6233, 192.2916, 
    197.1513,
  229.2479, 225.0169, 215.1072, 207.709, 200.0168, 193.2786, 189.5224, 
    190.3429, 194.1252, 194.5737, 194.282, 190.7103, 189.692, 194.212, 
    193.2007,
  228.9202, 226.9181, 215.9567, 206.64, 200.4834, 194.7494, 194.6315, 
    197.8137, 194.8112, 193.9961, 192.1856, 191.5606, 192.0083, 195.031, 
    196.0285,
  226.6973, 217.003, 212.6904, 205.3562, 203.6986, 202.7961, 200.8331, 
    200.1687, 196.7096, 192.1779, 191.3356, 190.9895, 193.5187, 194.1897, 
    196.2016,
  214.4465, 210.868, 207.3008, 203.289, 196.4825, 196.7529, 202.7814, 
    203.6153, 190.0631, 178.7191, 183.2891, 192.7206, 195.4894, 200.36, 
    202.6763,
  221.0699, 217.2081, 209.8939, 203.5816, 194.7547, 194.8265, 200.7621, 
    201.1562, 188.5182, 178.7509, 183.1828, 193.2783, 197.1636, 202.8053, 
    202.8679,
  223.8147, 223.4434, 218.5622, 205.239, 192.5612, 186.6533, 196.3008, 
    191.7575, 181.098, 174.6514, 185.8315, 195.1749, 200.5794, 207.0082, 
    206.6506,
  227.5158, 221.8702, 224.3876, 208.8663, 193.2434, 186.8744, 181.9066, 
    182.1765, 175.5237, 175.7475, 194.5734, 200.9908, 202.4412, 207.9859, 
    207.4635,
  225.743, 225.2352, 224.7828, 208.3005, 201.323, 180.6731, 180.5594, 
    182.9059, 182.4098, 190.1138, 198.7113, 201.4998, 205.4601, 207.8024, 
    208.4174,
  229.9282, 225.3691, 219.9906, 209.0173, 208.2468, 191.4774, 182.7218, 
    181.295, 188.974, 195.9832, 196.102, 200.7775, 204.7285, 205.7864, 
    208.9106,
  228.3596, 227.3452, 217.6125, 212.2793, 209.3554, 201.1358, 197.6017, 
    194.0447, 196.3031, 196.1842, 197.2021, 199.5365, 201.7598, 205.4232, 
    210.0318,
  231.0935, 226.5106, 217.6205, 207.4949, 203.9574, 202.255, 199.6285, 
    197.6875, 197.1139, 197.8357, 198.6627, 195.1006, 198.1611, 207.193, 
    207.9164,
  229.8016, 227.2988, 209.5396, 203.4928, 203.0205, 200.1549, 199.809, 
    197.6196, 196.1108, 193.6917, 189.5925, 189.5226, 197.3262, 204.7766, 
    204.533,
  228.563, 218.1, 208.9439, 203.4815, 202.0921, 198.4459, 195.4902, 194.399, 
    186.9175, 183.306, 184.6788, 187.753, 194.9435, 201.2827, 199.2237,
  203.5143, 206.0446, 205.0388, 201.17, 197.4945, 184.3704, 178.625, 
    178.6781, 190.3707, 192.1323, 185.9184, 180.8754, 184.0455, 185.7675, 
    193.6918,
  212.1207, 214.7705, 208.2149, 200.9571, 193.2948, 184.173, 173.6497, 
    169.7446, 178.8963, 180.2898, 180.548, 174.3962, 180.8952, 184.1782, 
    193.7964,
  215.9855, 225.0704, 221.9261, 201.3685, 191.8453, 178.681, 174.1921, 
    167.8884, 168.8806, 170.5006, 179.7452, 180.2897, 181.5222, 180.6459, 
    197.9247,
  222.9097, 228.1147, 222.5803, 207.8345, 192.7634, 181.3592, 173.9854, 
    175.5132, 174.0674, 173.805, 177.741, 185.4231, 189.9476, 195.8418, 
    203.8002,
  225.5943, 221.2764, 223.3723, 208.8014, 202.6061, 186.5293, 182.6719, 
    178.2532, 177.4826, 179.5142, 187.1105, 198.7933, 205.4676, 207.7679, 
    209.2511,
  223.7612, 224.1199, 216.5503, 213.8796, 210.0168, 203.0823, 189.5998, 
    189.448, 191.946, 201.5305, 204.7614, 207.8954, 209.0983, 207.9067, 
    210.1088,
  228.4962, 223.3897, 223.515, 211.0448, 208.7319, 206.2571, 206.7189, 
    205.0444, 205.1569, 205.2114, 206.5767, 208.2175, 210.0591, 209.7116, 
    211.4817,
  224.8844, 224.6911, 206.3974, 209.1878, 207.584, 206.2937, 208.2723, 
    209.2684, 208.6205, 207.9858, 207.8969, 208.0649, 208.8209, 210.2464, 
    211.4027,
  228.4929, 216.8124, 215.4933, 203.6931, 202.7292, 205.279, 207.6046, 
    207.7059, 207.5824, 207.4138, 206.4287, 210.3536, 210.6447, 210.6786, 
    211.3041,
  231.2315, 220.948, 210.5079, 203.1783, 193.5072, 189.8618, 193.7226, 
    199.4582, 205.1021, 195.2464, 203.6221, 209.0799, 211.7205, 212.3867, 
    210.2487,
  216.3712, 208.7606, 199.0186, 192.7905, 192.7878, 191.9724, 192.2158, 
    196.3782, 191.4882, 190.1826, 186.4914, 197.3437, 202.5925, 205.3976, 
    203.0442,
  220.9943, 215.0756, 204.1584, 200.1178, 198.8915, 198.8669, 195.8189, 
    197.142, 195.3243, 189.7857, 182.8786, 186.2141, 202.976, 203.4158, 
    203.2004,
  220.0597, 222.1709, 209.5518, 204.0131, 203.1259, 198.984, 203.9165, 
    199.5844, 197.178, 195.9853, 184.252, 179.2029, 192.3636, 208.1459, 
    206.6915,
  215.1646, 220.6772, 209.5912, 206.5675, 202.7871, 203.9288, 202.8759, 
    207.3942, 206.4289, 200.7083, 192.9867, 182.9892, 183.1239, 196.4857, 
    203.4201,
  211.0051, 212.8074, 211.238, 210.3204, 207.0822, 202.0351, 206.7099, 
    200.9591, 202.1749, 208.0996, 201.9302, 194.5068, 188.6933, 194.909, 
    198.5913,
  210.6426, 199.0356, 204.4802, 208.197, 208.2408, 204.0422, 204.5269, 
    204.1973, 203.9479, 207.9035, 207.0968, 204.2134, 200.3213, 198.8611, 
    199.0072,
  209.5985, 199.3, 198.323, 206.0618, 207.0761, 202.3503, 204.3851, 201.378, 
    202.3553, 210.2022, 209.5144, 207.6566, 205.0944, 205.8004, 202.7188,
  209.1674, 196.3837, 199.9214, 201.9204, 205.7046, 203.6747, 203.0758, 
    202.1399, 197.9777, 211.4191, 211.2928, 210.3399, 208.262, 206.9839, 
    207.7005,
  208.3096, 197.9008, 193.8215, 198.8365, 202.9001, 201.3854, 200.375, 
    202.027, 197.3017, 211.053, 213.1228, 212.1379, 209.7272, 207.6004, 
    204.5805,
  206.2921, 194.7946, 192.1901, 196.9189, 204.5526, 201.9482, 200.3255, 
    204.798, 201.3727, 202.1422, 213.4546, 213.1113, 212.0052, 208.9344, 
    204.2773,
  215.1974, 201.9777, 192.6148, 195.6463, 199.0271, 194.1724, 193.3956, 
    203.857, 204.7444, 198.8199, 194.3218, 200.1299, 203.097, 203.1749, 
    191.2893,
  211.004, 204.7484, 199.6612, 196.2993, 199.4656, 192.1448, 194.2133, 
    208.4339, 203.665, 198.9014, 196.5788, 199.9329, 205.6552, 205.5763, 
    200.1202,
  209.465, 211.3991, 203.1317, 196.3242, 197.5287, 194.198, 201.1141, 
    204.6759, 200.0593, 200.1413, 200.1439, 201.6451, 205.5539, 207.3452, 
    208.1321,
  209.9187, 216.1615, 203.6693, 193.9247, 189.7509, 196.6147, 202.1641, 
    211.7708, 205.6832, 203.818, 200.6839, 202.5205, 201.6587, 200.8994, 
    205.3062,
  216.5579, 217.4366, 206.6708, 190.8752, 194.1979, 203.8737, 210.1583, 
    203.8496, 200.9125, 209.1698, 202.301, 201.4781, 197.5489, 196.3912, 
    195.4422,
  220.8468, 220.6706, 207.3007, 191.2999, 195.524, 207.8983, 207.4733, 
    209.6886, 206.787, 207.2988, 204.8059, 202.6547, 198.706, 196.316, 
    188.6089,
  218.5962, 226.3965, 200.4832, 191.6486, 203.4263, 211.4864, 207.4823, 
    211.3971, 207.8043, 207.65, 206.3488, 202.8849, 199.4843, 194.7917, 
    186.4184,
  221.4837, 218.2825, 197.3994, 194.771, 209.372, 211.3618, 208.7185, 
    211.9778, 210.8335, 208.9263, 204.148, 201.6562, 198.4669, 197.5729, 
    192.0519,
  218.9021, 219.6359, 202.3946, 199.9332, 211.2493, 209.2988, 208.1123, 
    211.9172, 210.0431, 208.4859, 206.2944, 202.2018, 198.3376, 196.9529, 
    196.0341,
  221.5526, 219.6376, 208.7655, 202.492, 212.5191, 207.6433, 207.5515, 
    212.5087, 211.6134, 214.4697, 209.2271, 208.8763, 200.637, 198.9351, 
    194.6666,
  221.4283, 218.7423, 217.2774, 215.8379, 210.4825, 205.6954, 206.5482, 
    206.4134, 207.6723, 209.3322, 208.3925, 203.8851, 199.3304, 201.8508, 
    207.3199,
  220.773, 219.502, 219.5323, 216.2967, 211.2583, 212.3029, 209.7869, 
    211.1734, 209.9158, 211.3909, 207.5015, 204.1617, 200.1847, 201.8656, 
    207.2556,
  222.7271, 222.9871, 220.7523, 215.0454, 214.5021, 213.3181, 212.3441, 
    210.0819, 211.2244, 210.3093, 209.3244, 203.5728, 198.3035, 198.9598, 
    206.1947,
  220.4566, 217.2072, 223.2321, 213.1534, 212.0257, 216.3581, 210.9713, 
    212.5255, 208.8476, 210.0089, 210.5379, 202.154, 196.3617, 198.1373, 
    203.4454,
  217.8723, 215.5782, 220.1119, 215.3938, 213.9859, 212.0663, 212.4025, 
    204.7497, 202.7957, 211.1828, 205.5242, 201.6341, 197.9792, 201.586, 
    202.1794,
  217.088, 215.9673, 211.3587, 219.6226, 212.4005, 211.3394, 207.3227, 
    208.8697, 209.288, 209.7077, 205.5529, 207.8404, 203.7451, 203.2457, 
    202.7007,
  213.8765, 214.6574, 208.8948, 212.6384, 209.4198, 212.008, 208.3386, 
    208.1523, 209.527, 208.1764, 207.1993, 210.005, 203.0856, 206.3874, 
    204.387,
  213.8052, 213.6329, 208.4123, 206.5268, 206.1087, 212.1136, 208.7852, 
    209.3515, 210.592, 207.8976, 208.3396, 210.0488, 207.9467, 205.4444, 
    204.9995,
  218.3973, 214.2665, 209.9097, 206.2223, 205.5788, 211.3121, 209.461, 
    209.0024, 211.8518, 207.8734, 208.4369, 208.5387, 208.8782, 206.4368, 
    206.9441,
  218.5958, 215.6901, 213.453, 208.0023, 205.9565, 211.4395, 209.0589, 
    209.5195, 209.1039, 207.7284, 206.9098, 206.3792, 209.0707, 210.1084, 
    212.4212,
  226.4495, 219.2022, 214.9901, 210.2153, 208.8119, 211.0417, 211.1232, 
    211.0418, 210.5122, 208.759, 209.1054, 208.3499, 206.9655, 205.784, 
    204.7571,
  223.4687, 220.7908, 212.2733, 210.1633, 206.3081, 206.8846, 211.0251, 
    210.5379, 211.3802, 209.9831, 208.2757, 206.2497, 206.2565, 204.245, 
    205.5463,
  219.5023, 216.5967, 211.1857, 209.6049, 205.9632, 206.2887, 210.1828, 
    208.9412, 207.6988, 207.4097, 208.271, 204.9046, 204.74, 204.2362, 
    204.9128,
  219.8314, 214.4139, 206.5877, 207.2273, 204.7843, 208.6506, 208.0974, 
    209.4508, 208.1179, 204.382, 204.7932, 205.086, 204.6656, 204.978, 
    205.1877,
  221.9895, 208.7922, 207.6423, 209.0228, 205.3049, 207.034, 210.8808, 
    206.3621, 204.0633, 204.2222, 205.9109, 206.103, 205.9177, 206.5012, 
    206.5013,
  221.1709, 209.7562, 209.7597, 208.9544, 207.9645, 210.6564, 209.9202, 
    204.9323, 203.5371, 203.8288, 206.8529, 208.6059, 208.2194, 209.3815, 
    210.2743,
  217.1559, 207.9696, 212.3182, 209.4426, 212.1483, 213.348, 210.3474, 
    201.6214, 202.2011, 206.1369, 208.8936, 208.4622, 211.0721, 208.9952, 
    212.7004,
  215.0783, 210.062, 215.8625, 210.1991, 211.5893, 213.6479, 207.6161, 
    203.5205, 206.1047, 205.9129, 208.9799, 208.3484, 207.2304, 208.088, 
    212.3489,
  213.1326, 208.7755, 214.1783, 209.2379, 212.4655, 215.0759, 208.6838, 
    205.457, 206.9546, 208.1858, 204.6175, 203.9207, 205.5847, 206.3062, 
    208.0286,
  207.6298, 211.0819, 213.55, 208.0321, 212.9721, 214.332, 208.846, 208.598, 
    209.4141, 206.7314, 201.8384, 203.1115, 199.7613, 202.2676, 203.9997,
  208.4208, 208.5713, 209.8384, 203.8512, 211.6441, 210.5623, 209.8762, 
    210.1002, 210.7566, 206.2904, 205.4528, 204.3831, 203.2318, 204.8571, 
    204.3227,
  209.4193, 211.0552, 209.2162, 210.1295, 216.2807, 214.4006, 212.8272, 
    211.2071, 211.1767, 207.3837, 207.8058, 202.6086, 200.2924, 199.5676, 
    202.4519,
  210.426, 215.0532, 208.6301, 211.2331, 216.5959, 214.4506, 214.0595, 
    207.9801, 209.9122, 207.2102, 204.9422, 199.4211, 202.118, 204.2839, 
    203.1168,
  208.7014, 216.3897, 209.0013, 209.589, 216.7141, 216.2175, 210.3734, 
    211.6032, 210.6251, 206.7251, 204.1132, 201.6385, 203.072, 204.902, 
    202.9083,
  215.6525, 208.3419, 208.988, 211.9646, 218.9573, 215.696, 214.5499, 
    205.7938, 206.4829, 205.0626, 200.6222, 201.9324, 203.2851, 205.2307, 
    207.6505,
  213.0276, 209.424, 210.6168, 211.2956, 217.8905, 215.7085, 212.1251, 
    208.4742, 203.8643, 200.0789, 200.9479, 194.3124, 199.1577, 206.8313, 
    206.7145,
  211.8381, 209.4611, 210.9905, 212.4401, 216.6739, 216.027, 213.7851, 
    209.1621, 205.1008, 202.5514, 200.2539, 198.1667, 198.9594, 205.0041, 
    211.3379,
  214.8389, 209.902, 226.6417, 214.2281, 216.5925, 217.4871, 215.5411, 
    211.4599, 205.605, 203.4724, 199.6502, 195.0461, 198.6174, 199.6171, 
    208.2754,
  213.5019, 210.4243, 221.7369, 215.2259, 214.8892, 217.4313, 214.8994, 
    212.8468, 208.9116, 204.754, 201.9232, 201.3048, 196.587, 202.445, 
    202.5006,
  212.2641, 211.8798, 216.006, 214.5944, 214.363, 215.9081, 215.0664, 
    219.2161, 212.3759, 207.4195, 204.3024, 196.1763, 192.8184, 196.9203, 
    197.6914,
  221.7586, 218.8247, 217.5538, 214.5744, 210.752, 208.8207, 206.8058, 
    207.2036, 207.4143, 208.892, 207.7984, 207.8372, 207.7112, 205.6353, 
    204.8306,
  223.1312, 221.6472, 218.476, 215.1204, 213.065, 208.7809, 206.4227, 
    206.7616, 206.2264, 207.0051, 204.2823, 205.5485, 207.2723, 207.516, 
    205.3655,
  215.324, 217.017, 219.8907, 217.5352, 213.2409, 208.7311, 207.7394, 
    204.6867, 204.7593, 206.5169, 205.3637, 207.0712, 205.9716, 202.0217, 
    203.3842,
  213.0617, 207.9957, 209.6396, 216.326, 212.713, 209.4567, 206.4468, 
    206.3654, 206.2483, 206.1616, 206.243, 206.7465, 205.1051, 201.9633, 
    199.475,
  211.6616, 205.0328, 210.4075, 214.2746, 213.0138, 206.1067, 206.063, 
    202.6609, 206.2066, 206.0136, 205.9281, 207.6724, 206.5927, 198.7765, 
    198.8179,
  206.4091, 205.1558, 210.5676, 213.0896, 211.4082, 205.7688, 203.1889, 
    204.8793, 202.5792, 200.3276, 200.061, 206.5493, 205.9452, 202.8603, 
    196.8742,
  206.2662, 208.2098, 212.291, 215.1614, 211.8208, 208.9693, 205.067, 
    199.9598, 196.333, 198.3006, 203.56, 206.1389, 205.9676, 200.3827, 196.864,
  206.0578, 211.2836, 219.2206, 211.1092, 208.9361, 206.4354, 204.6296, 
    201.5084, 198.976, 201.3671, 202.2117, 206.75, 206.4825, 200.9277, 
    200.9365,
  209.9196, 215.0152, 213.904, 207.5204, 206.5232, 203.1787, 200.9126, 
    199.1331, 199.1673, 199.7862, 203.7617, 203.4296, 206.5686, 202.7925, 
    197.0316,
  213.8462, 222.4572, 209.9452, 205.5997, 204.1547, 202.6167, 201.601, 
    202.8934, 201.7207, 201.2527, 202.972, 203.6548, 204.052, 201.5012, 
    199.414,
  205.2905, 208.7325, 206.5909, 208.3873, 210.0842, 212.6839, 211.011, 
    210.8793, 211.4076, 210.923, 210.9535, 208.7597, 209.6779, 207.4663, 
    206.1119,
  204.7318, 208.0542, 208.5127, 210.5737, 214.396, 217.941, 214.3382, 
    212.2319, 210.615, 206.7784, 209.0819, 208.5729, 211.194, 207.9205, 
    206.3437,
  206.7175, 212.1747, 216.4656, 215.1968, 218.4201, 217.3128, 212.7713, 
    206.9238, 203.7081, 206.4485, 208.678, 208.1841, 210.7327, 211.5107, 
    209.4193,
  215.182, 219.1766, 220.5238, 217.0623, 218.6312, 215.774, 212.6488, 
    211.0016, 202.8768, 200.556, 205.4508, 206.715, 207.2419, 209.0432, 
    210.0433,
  216.8705, 224.3958, 219.0889, 220.3201, 218.7354, 212.0188, 207.8379, 
    209.0858, 204.3936, 203.2365, 200.0278, 199.7766, 197.4083, 198.2064, 
    199.4951,
  220.9385, 221.9126, 221.2772, 224.9893, 220.361, 207.8941, 203.9642, 
    201.7003, 204.6842, 200.7231, 198.2237, 196.9195, 195.4253, 195.3369, 
    194.0008,
  221.293, 220.5235, 218.3087, 223.0343, 215.442, 206.291, 201.8578, 
    198.3215, 195.7126, 199.1197, 200.3383, 201.0779, 198.0554, 198.8461, 
    194.6202,
  218.1588, 217.8283, 220.8838, 217.8776, 209.2564, 204.0114, 200.6469, 
    200.2542, 203.8262, 205.0877, 204.2076, 203.1349, 201.2232, 198.3282, 
    198.7099,
  217.4681, 219.6633, 224.1386, 212.0292, 207.7375, 205.6066, 206.5114, 
    209.7107, 207.2742, 207.5754, 206.9857, 206.0105, 203.6563, 201.6535, 
    200.8546,
  221.8506, 229.0494, 215.6104, 211.2146, 211.4289, 211.9212, 212.242, 
    212.4491, 209.4376, 208.8131, 209.2789, 208.8392, 206.3357, 203.6508, 
    203.2204,
  208.7178, 200.2657, 197.8855, 196.0196, 198.8531, 212.2521, 221.1295, 
    218.4628, 216.8068, 217.4326, 211.4062, 203.9892, 203.7425, 207.0433, 
    207.0475,
  209.2728, 204.4526, 201.4837, 198.1444, 208.1522, 219.4404, 217.4665, 
    215.5898, 211.4719, 205.2618, 203.3016, 199.9845, 201.1053, 201.3394, 
    204.4057,
  213.6707, 201.9014, 203.1478, 205.5165, 222.4809, 218.8649, 217.9644, 
    212.2103, 210.6914, 202.9394, 200.2245, 195.7047, 194.1911, 198.4397, 
    200.4184,
  211.6335, 207.1632, 207.854, 210.6236, 216.8429, 219.2897, 215.5632, 
    217.2023, 210.5288, 196.8445, 195.8993, 193.674, 190.7869, 193.4489, 
    197.4683,
  211.3414, 206.7121, 214.1833, 218.8034, 215.9249, 213.3207, 212.8326, 
    207.587, 202.9718, 199.1195, 198.503, 200.7573, 199.1279, 203.8644, 
    202.5115,
  211.1175, 211.9548, 222.5787, 221.8089, 217.7428, 213.1049, 210.9174, 
    207.155, 204.0002, 203.3202, 205.1363, 207.0685, 209.2155, 210.0291, 
    209.961,
  214.9498, 220.9496, 224.9108, 219.8656, 216.2037, 214.0844, 212.0972, 
    209.3781, 208.1941, 210.0482, 208.8505, 208.7946, 208.6661, 210.472, 
    211.6743,
  219.5278, 221.5724, 228.6902, 218.2201, 215.1701, 214.9181, 214.2955, 
    212.3184, 208.1051, 206.4038, 205.1864, 205.4891, 204.396, 203.6744, 
    206.5391,
  220.8152, 223.0073, 223.9911, 215.9202, 213.8755, 214.1054, 211.8464, 
    209.3041, 207.5873, 205.8804, 204.2406, 205.9324, 203.4602, 202.8522, 
    202.7489,
  221.0089, 222.4189, 222.3887, 211.65, 213.2933, 212.7563, 210.2966, 
    212.7098, 206.9288, 203.7329, 201.764, 205.2366, 206.6268, 205.0517, 
    205.4792,
  225.6842, 225.1984, 221.9202, 219.1975, 218.5366, 214.1122, 214.1526, 
    212.8243, 213.1184, 208.2603, 205.4632, 201.476, 197.1813, 195.895, 
    187.8942,
  223.4327, 221.6118, 221.9239, 218.5773, 217.1453, 215.4261, 214.424, 
    214.5197, 214.6329, 211.0028, 208.1447, 204.0284, 199.2045, 194.1094, 
    195.0205,
  222.3654, 221.3958, 218.9507, 216.5856, 216.0728, 210.8785, 213.9826, 
    212.2828, 209.9, 212.6102, 212.3651, 209.8047, 206.091, 199.9581, 196.5499,
  220.2886, 220.4129, 220.6428, 212.5916, 212.6932, 212.6005, 208.3446, 
    210.9148, 212.4102, 210.027, 210.8367, 210.7277, 210.4364, 203.375, 
    201.3276,
  220.4326, 217.9833, 219.2173, 213.0257, 211.312, 208.8499, 209.821, 
    204.7531, 203.6665, 207.9755, 209.2261, 207.8924, 208.6635, 209.1296, 
    208.0005,
  218.8983, 216.9592, 216.7886, 214.2413, 211.3727, 210.2749, 206.9124, 
    203.169, 201.2727, 204.481, 208.0195, 206.7687, 206.608, 208.2566, 
    207.1581,
  218.7353, 218.034, 215.5282, 211.707, 209.3167, 208.1299, 205.04, 204.1204, 
    205.3701, 204.3087, 208.6947, 208.1308, 204.8403, 206.2804, 207.5595,
  217.1646, 217.0435, 216.9771, 214.1133, 208.2392, 206.4717, 204.1308, 
    204.2102, 206.5083, 207.3125, 204.2044, 205.6999, 205.7177, 205.6043, 
    204.4301,
  213.6388, 217.5098, 217.3119, 212.8048, 207.5031, 206.1256, 204.1553, 
    202.5688, 204.3644, 205.3341, 204.0077, 202.9769, 208.1369, 210.3567, 
    208.8008,
  211.2041, 215.1341, 215.1602, 210.8642, 203.7152, 201.9358, 202.3982, 
    205.8856, 205.7832, 204.0014, 203.8074, 202.8329, 210.6222, 210.7317, 
    211.5882,
  194.9016, 199.5718, 199.8492, 206.891, 206.8501, 203.9887, 194.4277, 
    197.4158, 200.1229, 205.7645, 209.8279, 207.9146, 211.1421, 205.5823, 
    201.7758,
  194.3294, 195.7458, 196.462, 205.6994, 204.937, 201.366, 193.5338, 190.705, 
    196.9553, 201.0169, 204.8093, 206.7794, 208.4851, 208.7656, 206.7908,
  191.8129, 192.1177, 195.6976, 199.0034, 202.2685, 202.5372, 196.8471, 
    187.1874, 189.5236, 198.5979, 203.4029, 206.7779, 208.55, 211.1342, 
    210.0406,
  191.0989, 188.7255, 193.7277, 197.5811, 196.2113, 197.086, 191.1027, 
    188.5621, 189.2259, 195.3754, 199.4944, 204.2478, 207.8284, 210.679, 
    210.7503,
  186.8399, 190.8367, 190.6777, 197.544, 196.2773, 187.8594, 185.5719, 
    186.0413, 191.5577, 193.422, 199.8663, 201.3698, 205.6294, 210.2421, 
    209.9334,
  193.8723, 188.8303, 190.5712, 197.0023, 201.4165, 189.2908, 180.6966, 
    182.1271, 188.2828, 190.67, 195.6526, 202.4165, 205.9784, 209.2787, 
    207.8446,
  193.3075, 190.9227, 192.8076, 199.0365, 201.8724, 193.7164, 184.9014, 
    186.0846, 189.4639, 197.1359, 195.073, 200.9711, 205.8263, 208.3045, 
    208.6347,
  191.8577, 185.8233, 194.3833, 203.3614, 201.3979, 190.6669, 194.0496, 
    191.9996, 191.9265, 198.2413, 197.8728, 203.3017, 205.2839, 208.4495, 
    209.4296,
  193.6522, 186.0549, 197.8122, 206.4707, 197.3633, 197.0831, 196.2448, 
    194.4493, 196.0529, 196.7994, 199.7858, 203.9715, 204.9, 208.8522, 
    208.9747,
  190.1815, 191.8447, 205.503, 204.6746, 198.915, 203.6635, 200.915, 
    197.9397, 201.887, 200.5729, 202.2691, 204.3232, 205.3697, 207.5764, 
    205.793,
  198.7191, 190.9124, 184.351, 186.5214, 183.2448, 180.4183, 180.4471, 
    183.6386, 183.8327, 186.9158, 188.0655, 193.8343, 205.4789, 212.1704, 
    210.5441,
  198.5887, 197.1272, 195.863, 194.8089, 190.8893, 183.6766, 183.697, 
    188.2243, 190.1003, 193.5676, 194.5255, 193.4834, 201.2501, 209.2324, 
    208.9426,
  207.7044, 205.9643, 204.4274, 199.2424, 193.6254, 190.7629, 197.8586, 
    192.8564, 197.1591, 204.7641, 206.3521, 197.3524, 199.0137, 207.1042, 
    210.0941,
  207.9875, 207.345, 206.1398, 198.4783, 196.8001, 202.6471, 210.3714, 
    209.8868, 207.212, 207.9579, 206.2549, 197.7302, 198.5438, 202.0257, 
    206.7055,
  211.4952, 209.8596, 206.6298, 204.9468, 204.9001, 212.4918, 215.955, 
    213.4783, 208.9282, 211.1626, 202.1527, 195.3865, 193.9271, 198.9678, 
    204.003,
  211.7323, 210.0087, 204.8898, 207.7013, 209.582, 209.4287, 211.0666, 
    214.9365, 214.6613, 210.8009, 204.0862, 195.9405, 190.7563, 193.0249, 
    203.5128,
  215.0042, 206.2391, 208.0084, 214.3159, 215.3561, 214.8432, 215.5105, 
    213.8969, 211.7485, 212.3133, 208.2225, 194.2216, 189.8416, 191.4868, 
    201.3814,
  213.3038, 207.8023, 213.8714, 215.6552, 214.1278, 216.1755, 214.7642, 
    211.7996, 211.6018, 211.446, 206.9653, 201.1332, 192.4281, 195.4709, 
    202.2236,
  207.7593, 202.3087, 210.151, 213.2635, 215.3003, 214.9986, 211.5515, 
    211.4656, 210.3745, 210.3356, 208.3152, 205.4394, 203.9198, 207.1201, 
    208.0226,
  205.2333, 203.6874, 213.76, 214.8438, 215.7258, 214.3247, 213.1901, 
    212.1838, 211.1499, 208.6147, 204.4382, 204.3745, 202.8694, 204.8223, 
    206.4987,
  220.7596, 214.5732, 215.263, 219.7837, 217.706, 216.6887, 216.4428, 
    213.0911, 209.6466, 205.5109, 200.7671, 193.273, 189.1486, 192.0054, 
    198.6525,
  213.6536, 214.862, 217.7604, 216.5249, 220.7441, 215.6041, 213.9485, 
    213.4974, 212.9386, 208.1093, 207.2748, 196.4571, 190.1374, 192.7561, 
    194.7002,
  211.1512, 209.0226, 215.8225, 215.7814, 219.2932, 213.7524, 213.7763, 
    211.8174, 210.8691, 210.67, 214.9053, 210.9226, 191.8097, 189.9304, 
    191.5599,
  210.6299, 207.2696, 212.2875, 214.5802, 216.8806, 215.5794, 208.7538, 
    211.4712, 213.3525, 212.4876, 210.3054, 201.5616, 191.236, 186.0054, 
    190.9271,
  209.5842, 205.0472, 216.2489, 213.4336, 211.7889, 209.7646, 210.8057, 
    205.3203, 202.8699, 209.4677, 203.6555, 198.7172, 191.5714, 188.5697, 
    193.2853,
  216.4931, 205.7927, 210.6579, 212.4288, 210.0544, 208.8206, 206.5964, 
    206.9087, 206.6299, 208.1916, 202.6481, 199.1518, 192.8197, 189.2853, 
    195.7274,
  215.5202, 207.6236, 212.9353, 210.927, 208.3485, 205.2645, 206.1444, 
    205.4946, 205.6832, 208.1703, 202.7826, 192.3991, 193.4556, 193.3426, 
    195.3221,
  213.4, 209.476, 211.8046, 208.0486, 206.1078, 204.1001, 204.0722, 205.7434, 
    205.9095, 209.0577, 207.5007, 199.9039, 189.7436, 192.0814, 197.0455,
  213.5242, 211.3511, 210.6333, 206.3134, 202.5938, 200.996, 201.1556, 
    202.2371, 204.2847, 207.1736, 208.3132, 207.7329, 201.4919, 201.108, 
    204.7219,
  218.8281, 214.151, 208.4927, 203.7653, 200.1267, 198.6495, 198.3658, 
    201.7615, 205.3648, 206.3779, 206.8307, 205.3196, 206.7888, 207.0044, 
    209.459,
  215.8522, 207.3129, 206.2015, 203.0809, 203.2925, 204.8971, 206.7092, 
    206.6793, 207.7493, 208.0136, 208.3296, 209.4715, 213.7303, 213.1624, 
    211.7468,
  210.6851, 211.5652, 206.4701, 201.7822, 206.3891, 205.4568, 205.2224, 
    208.1605, 208.375, 207.944, 209.4372, 209.7869, 210.1781, 213.9753, 
    216.1503,
  211.025, 203.7319, 204.6398, 202.9073, 203.9174, 206.3856, 206.7607, 
    203.8645, 206.6049, 204.7777, 204.9022, 207.0675, 214.7743, 215.0037, 
    211.6801,
  209.1158, 209.716, 205.6328, 202.6223, 202.9918, 203.9452, 205.0354, 
    205.848, 207.7362, 197.4042, 194.6075, 195.0537, 198.5791, 205.6908, 
    202.3943,
  216.3023, 209.9089, 201.1706, 200.0401, 201.5113, 203.6552, 204.7838, 
    204.3591, 204.5481, 196.0882, 188.2726, 190.3833, 192.566, 195.3401, 
    194.2039,
  219.2076, 208.0967, 202.3906, 199.7662, 206.7408, 202.1307, 201.582, 
    207.1471, 205.5693, 194.1148, 185.4245, 185.6745, 186.7332, 189.0249, 
    190.7696,
  219.3987, 208.6119, 203.8756, 200.3358, 205.2919, 203.3964, 204.4867, 
    203.8973, 207.1463, 198.7481, 190.0588, 182.5637, 182.924, 186.2499, 
    189.3397,
  218.0446, 208.7365, 204.5284, 200.0976, 204.9812, 204.3533, 206.3356, 
    206.5802, 209.5686, 202.645, 194.3592, 188.2745, 181.2591, 180.3932, 
    185.2811,
  219.7886, 206.9057, 202.2033, 201.5911, 205.8828, 210.3155, 208.214, 
    208.0145, 209.2691, 207.9871, 199.7842, 191.6134, 190.5717, 188.9513, 
    197.7932,
  217.9955, 210.5536, 210.7611, 206.2036, 208.1569, 210.1306, 210.495, 
    209.135, 209.5898, 209.8201, 207.0321, 201.5923, 198.4763, 202.1124, 
    208.3136,
  209.0685, 208.7702, 215.2573, 213.0664, 212.9187, 208.4389, 206.4749, 
    203.9941, 206.0834, 207.2601, 209.1436, 205.7506, 199.7213, 195.1, 
    198.9284,
  205.7925, 213.3794, 217.1063, 214.1449, 213.1394, 209.5518, 205.5283, 
    203.1317, 206.0806, 207.8746, 210.8396, 207.5723, 208.4881, 204.3869, 
    203.4977,
  206.5654, 214.7948, 215.6559, 216.748, 213.8801, 206.9406, 204.2122, 
    192.9025, 190.5713, 206.3913, 210.7835, 207.8469, 210.0323, 210.6151, 
    208.4829,
  201.9855, 214.1902, 213.5734, 213.103, 212.8657, 210.2094, 199.7311, 
    188.3126, 186.7932, 193.4458, 208.6563, 210.9627, 210.6477, 215.65, 
    212.9475,
  206.088, 216.5516, 213.0279, 212.707, 211.9621, 208.5408, 206.1383, 
    191.0094, 186.1782, 183.207, 192.2671, 211.1273, 212.7745, 209.5003, 
    210.2996,
  203.6873, 218.8093, 215.045, 214.3293, 211.5242, 208.5411, 206.9306, 
    192.0626, 181.1075, 180.3371, 180.7973, 194.5895, 211.3045, 215.2907, 
    212.4467,
  204.5414, 218.7706, 217.3787, 211.1368, 210.6695, 209.4642, 207.4475, 
    199.5916, 183.6523, 177.5881, 172.9659, 182.6044, 196.5864, 213.7842, 
    217.156,
  206.9694, 215.6164, 215.4555, 212.2632, 210.8021, 210.1013, 210.4053, 
    207.568, 194.7158, 181.836, 177.6588, 178.5336, 185.7358, 201.9395, 
    214.2867,
  208.7805, 217.3818, 214.4534, 211.3812, 210.6935, 210.1123, 210.956, 
    209.2254, 205.0367, 189.1124, 180.535, 179.981, 182.271, 187.722, 203.5424,
  204.9276, 218.1244, 221.5201, 210.608, 210.08, 209.7476, 210.1441, 
    210.5074, 210.5765, 203.3786, 188.1952, 186.8497, 189.7676, 188.5345, 
    194.9258,
  197.0694, 198.2854, 205.3055, 214.9963, 212.5647, 210.902, 198.2332, 
    193.6427, 202.3385, 214.0764, 209.8361, 210.0238, 210.4125, 198.689, 
    196.139,
  195.2742, 201.206, 212.9952, 215.7723, 216.0399, 209.2414, 194.5064, 
    195.2895, 201.9547, 211.906, 213.6413, 210.6011, 214.9853, 202.1425, 
    199.9842,
  211.1423, 212.5664, 220.5835, 217.7019, 215.3212, 207.0127, 192.1306, 
    182.4206, 186.6092, 209.0929, 216.4063, 214.9421, 216.1402, 209.8509, 
    203.488,
  213.4397, 218.2731, 216.3437, 213.5824, 211.2128, 208.2319, 187.456, 
    177.4434, 180.9954, 198.2218, 217.9521, 216.5478, 217.1163, 216.4013, 
    209.375,
  215.4642, 214.1613, 213.1483, 212.4865, 209.235, 202.0688, 192.0331, 
    189.1853, 187.3302, 191.1449, 208.5233, 218.2323, 219.3495, 216.782, 
    214.3096,
  214.6111, 214.8374, 212.3195, 213.2235, 208.3005, 202.831, 192.3311, 
    187.0314, 182.9807, 186.547, 202.8702, 216.3342, 218.4983, 219.6666, 
    218.1938,
  216.137, 214.7159, 215.0295, 211.6078, 209.2274, 206.5789, 198.2464, 
    185.461, 183.4485, 188.131, 196.4595, 211.3002, 217.7232, 219.8739, 
    219.765,
  215.05, 214.4536, 214.8123, 210.9172, 209.3953, 208.0072, 205.143, 198.696, 
    193.7811, 189.7205, 192.4577, 205.55, 214.5454, 218.2478, 220.7663,
  216.0124, 217.6954, 218.8454, 211.2732, 209.1041, 212.4701, 212.9417, 
    208.6495, 195.1837, 194.1368, 194.5557, 201.8722, 212.2404, 217.7622, 
    217.7386,
  213.348, 215.9518, 223.1994, 212.8454, 211.6763, 217.0276, 214.1067, 
    213.0676, 208.6017, 201.4146, 197.4155, 202.2979, 207.1913, 208.2644, 
    215.78,
  196.2157, 199.4205, 210.2528, 214.4509, 213.8672, 209.9307, 211.9506, 
    211.5479, 201.0999, 213.8189, 213.9071, 214.2216, 211.2111, 196.3478, 
    188.2366,
  207.565, 209.2685, 218.754, 216.3595, 212.6576, 209.5142, 208.9899, 
    210.3822, 204.4332, 214.4599, 216.1358, 215.1712, 210.3808, 198.6733, 
    191.7217,
  218.5835, 215.4869, 217.4083, 210.886, 208.2714, 208.1452, 196.336, 
    187.2205, 195.6702, 213.9909, 216.2431, 215.3386, 214.2347, 205.6734, 
    190.7057,
  213.5159, 212.6613, 211.2553, 208.9409, 201.2016, 202.2299, 192.0778, 
    186.2434, 198.5907, 208.5878, 215.1411, 215.9507, 214.2709, 210.9501, 
    194.3628,
  212.6126, 211.5296, 210.2832, 208.3455, 202.2261, 199.9406, 200.1153, 
    203.8943, 206.4836, 209.361, 214.5524, 215.8726, 215.1664, 210.8083, 
    200.7159,
  219.7163, 215.0858, 211.4338, 209.4595, 205.7737, 203.1041, 203.3578, 
    203.7728, 201.0675, 205.6675, 213.4613, 214.5643, 216.3401, 210.4604, 
    204.5605,
  215.9014, 217.478, 212.4037, 212.0927, 211.0559, 208.6414, 207.9874, 
    206.6909, 203.6892, 204.458, 211.2326, 212.4583, 218.0647, 213.0264, 
    207.3051,
  215.1698, 220.5681, 223.4768, 216.167, 214.4625, 211.7286, 212.5063, 
    214.4386, 211.8092, 211.5629, 211.1154, 212.7946, 215.6575, 217.4991, 
    215.4267,
  210.9881, 216.758, 223.4097, 217.1986, 217.4516, 213.827, 213.2585, 
    211.9419, 212.0102, 212.3085, 213.7569, 212.6953, 211.8102, 219.0141, 
    219.1197,
  209.3247, 212.1507, 222.1614, 217.2276, 219.6219, 214.5995, 213.3206, 
    213.2823, 212.6062, 213.5008, 216.4608, 214.3952, 211.3873, 212.4298, 
    219.662,
  224.2022, 217.0697, 215.0303, 212.7811, 207.0125, 206.6946, 212.1039, 
    211.4654, 205.6642, 205.9758, 208.1892, 206.796, 208.4263, 209.2131, 
    206.4742,
  226.045, 219.8316, 215.8264, 208.2673, 207.357, 208.6471, 211.9363, 
    212.9409, 211.9349, 207.2056, 205.0787, 206.7276, 208.7455, 207.0184, 
    208.5802,
  214.7582, 212.362, 217.4061, 208.9323, 209.9493, 209.6177, 212.5828, 
    210.2796, 205.4619, 205.1398, 205.9806, 208.5667, 212.7528, 211.7029, 
    208.5358,
  213.9889, 212.7199, 215.6697, 213.2693, 212.1447, 213.8544, 212.6249, 
    212.9329, 210.9354, 204.6485, 205.3298, 209.491, 212.8763, 202.014, 
    200.7272,
  214.1872, 214.5111, 215.1732, 212.7019, 213.0164, 211.3512, 212.4316, 
    209.3743, 205.4886, 205.8624, 205.4847, 208.7379, 214.7069, 202.4986, 
    204.9829,
  212.4975, 213.1349, 215.9144, 213.615, 213.361, 210.7276, 210.0814, 
    211.5853, 210.0984, 206.7216, 205.6568, 207.3988, 209.4267, 203.0713, 
    209.3409,
  212.4052, 214.0043, 222.974, 219.5972, 213.6907, 211.41, 210.2505, 
    210.3854, 209.6939, 206.2025, 206.8994, 206.7585, 209.1839, 204.8557, 
    206.2234,
  211.5714, 213.0585, 230.6784, 218.3671, 213.9584, 211.7385, 209.8097, 
    210.447, 211.049, 211.0251, 205.994, 207.5888, 207.8156, 210.7612, 
    205.6174,
  215.9717, 228.7899, 225.9904, 217.2465, 215.217, 212.4594, 209.8193, 
    210.4095, 210.6, 213.1781, 208.3553, 206.3269, 208.4872, 208.9657, 
    205.3592,
  209.731, 224.2605, 224.3417, 218.0008, 214.3626, 213.1091, 212.751, 
    211.5953, 210.204, 213.5947, 212.5692, 206.9617, 206.6153, 206.7006, 
    208.502,
  223.037, 215.0178, 212.9115, 212.9526, 212.0383, 210.683, 213.1017, 
    213.5104, 214.1809, 207.822, 204.3129, 201.2019, 201.0188, 202.7301, 
    203.3392,
  218.5608, 213.1118, 214.3375, 212.845, 212.6364, 211.9973, 211.5217, 
    216.0548, 215.637, 210.5426, 203.8122, 203.3766, 205.5602, 205.8322, 
    203.3199,
  216.8422, 213.751, 217.0665, 212.169, 212.7775, 208.2226, 215.2076, 
    213.7611, 212.0429, 205.3562, 204.5035, 206.3031, 206.5546, 206.9769, 
    198.8756,
  214.2136, 222.5459, 213.414, 212.969, 211.3132, 212.1591, 209.1992, 
    214.9226, 215.2081, 209.0711, 207.3758, 204.5133, 206.7396, 206.4425, 
    203.4805,
  218.3648, 224.0584, 219.1056, 212.4417, 207.91, 206.5287, 209.0662, 
    208.3097, 207.1057, 211.7787, 207.1835, 207.3237, 206.1763, 214.3905, 
    209.9904,
  215.4926, 224.3323, 222.1235, 212.7329, 207.6615, 205.088, 207.7784, 
    209.8315, 210.7372, 210.7844, 207.9032, 204.338, 204.8314, 212.1427, 
    205.9135,
  211.2994, 220.4236, 224.5214, 212.5994, 204.0244, 203.8468, 207.3807, 
    209.3063, 210.0309, 210.2181, 209.009, 204.6421, 204.3287, 205.6712, 
    215.4712,
  211.2616, 215.0354, 224.2634, 211.5516, 204.5845, 202.6595, 207.6593, 
    209.9332, 211.8508, 210.6221, 210.9691, 206.1843, 204.6785, 217.632, 
    220.8721,
  221.7443, 217.6488, 221.3371, 211.651, 204.3263, 205.1318, 209.9684, 
    209.4133, 211.9019, 213.0734, 211.1704, 209.8037, 206.0469, 219.7171, 
    224.1393,
  218.1155, 221.9149, 210.4233, 209.1394, 205.6104, 205.0342, 207.083, 
    210.2985, 212.1243, 213.7125, 211.8126, 211.6749, 212.2554, 219.6775, 
    221.7265,
  219.7935, 216.4931, 213.7242, 211.06, 209.3122, 207.5599, 206.6559, 
    211.5535, 214.1663, 209.5216, 207.563, 206.9501, 205.573, 205.1104, 
    205.9405,
  220.5802, 214.6479, 213.2159, 209.3116, 208.587, 209.1109, 205.576, 
    210.3263, 211.751, 211.0307, 208.4582, 208.1669, 207.5431, 202.2921, 
    212.3297,
  217.8313, 215.0996, 211.5544, 207.3627, 209.2477, 205.7445, 208.2616, 
    206.6222, 208.1767, 206.7077, 209.098, 206.8116, 204.4963, 203.0217, 
    211.8988,
  222.7907, 215.1099, 208.825, 202.1018, 199.8162, 203.8226, 204.776, 
    206.2338, 203.518, 207.435, 206.4073, 205.6098, 204.6634, 208.2945, 
    212.8286,
  211.5952, 210.9055, 208.3046, 202.1078, 196.962, 198.5471, 201.4013, 
    203.8329, 204.7012, 203.8992, 202.4842, 206.2953, 205.0527, 210.6782, 
    214.0897,
  203.9326, 200.9796, 204.103, 194.4538, 199.1216, 199.3431, 193.9128, 
    198.7809, 201.0845, 196.4387, 200.5128, 204.2256, 205.3964, 217.646, 
    216.1028,
  202.6852, 201.47, 200.595, 202.5873, 201.8895, 200.4232, 197.4003, 
    195.2316, 195.1262, 199.9526, 205.6207, 208.2247, 205.0337, 218.9202, 
    217.0728,
  200.8461, 196.103, 202.2093, 206.0337, 204.0217, 201.6631, 198.5119, 
    198.6699, 198.669, 201.1568, 206.2016, 208.7227, 205.7131, 217.2402, 
    218.0671,
  204.2456, 202.4755, 204.8738, 210.2456, 204.5755, 201.8001, 201.7126, 
    195.7019, 199.3084, 207.8857, 212.133, 211.4362, 215.2668, 218.4953, 
    218.7119,
  206.1239, 207.9067, 211.1269, 209.2946, 206.9813, 205.6031, 200.4088, 
    200.9664, 207.106, 213.7715, 213.9285, 211.813, 218.731, 217.5963, 
    215.7759,
  207.316, 209.7947, 204.4276, 199.3297, 193.6793, 190.7424, 193.6785, 
    195.5197, 191.5431, 196.0655, 202.7892, 206.3157, 207.6167, 208.4638, 
    207.237,
  211.6786, 207.0979, 202.9177, 198.4126, 196.8125, 193.0588, 191.2307, 
    192.0744, 193.9429, 187.0909, 200.1791, 206.6896, 208.6027, 209.5209, 
    210.4777,
  207.8229, 201.156, 200.5137, 197.8471, 194.8683, 195.2773, 192.9464, 
    187.5574, 189.6376, 195.0438, 195.4272, 202.5664, 208.0457, 209.324, 
    211.005,
  209.4027, 204.0332, 201.0862, 197.9585, 199.8032, 200.6465, 197.6366, 
    200.6728, 198.6177, 194.5804, 195.8869, 201.6506, 210.0516, 208.7363, 
    210.8163,
  213.5228, 213.0552, 207.2742, 204.6888, 207.368, 206.1131, 204.9176, 
    204.4799, 208.3794, 208.263, 201.3228, 199.2566, 205.1654, 210.0856, 
    210.7788,
  220.6868, 219.4373, 209.2748, 210.5272, 210.8587, 208.6406, 206.4704, 
    206.3734, 213.5801, 209.387, 212.4053, 206.2499, 207.0409, 210.7639, 
    211.5691,
  221.5443, 219.9509, 215.4996, 211.2072, 212.6826, 211.9238, 214.5089, 
    211.2385, 210.5826, 219.0371, 214.0726, 211.4408, 210.8284, 215.4806, 
    213.1611,
  221.3711, 215.4007, 212.9946, 208.9791, 211.2205, 210.592, 213.6313, 
    214.2648, 214.5532, 218.549, 216.4275, 214.2784, 213.5445, 212.9572, 
    212.0838,
  221.1497, 219.1812, 212.8386, 210.188, 208.3785, 209.4292, 209.1241, 
    213.4736, 215.0046, 219.6732, 213.1584, 217.0598, 215.5152, 211.4998, 
    213.6344,
  224.3634, 213.6673, 214.7446, 213.976, 209.3692, 208.6041, 209.2414, 
    210.5347, 209.1082, 212.2898, 215.3201, 215.8908, 213.3771, 209.9439, 
    214.21,
  228.163, 223.7619, 219.8671, 218.1709, 215.3826, 215.4223, 213.7385, 
    207.213, 204.2332, 201.2055, 194.4662, 189.7794, 196.3265, 202.3045, 
    207.237,
  216.969, 222.2623, 218.0078, 216.1627, 215.7844, 214.5651, 208.8049, 
    210.9438, 207.8828, 198.9349, 194.364, 187.8676, 194.6696, 201.0748, 
    208.1144,
  221.289, 221.868, 218.4788, 213.5304, 214.6245, 207.2484, 207.4129, 
    207.9564, 210.7764, 207.2489, 196.8536, 190.3426, 193.0768, 202.2883, 
    209.5919,
  221.2017, 219.8799, 219.5337, 208.4226, 203.3825, 200.3031, 201.0706, 
    201.0883, 210.5381, 211.8722, 206.4988, 193.4164, 190.7484, 202.4572, 
    210.907,
  220.1007, 222.615, 219.7715, 208.2486, 203.3638, 197.1732, 199.6615, 
    201.7377, 206.5829, 214.1169, 209.0822, 201.1149, 192.7731, 202.1336, 
    211.5928,
  219.2858, 222.776, 211.4922, 202.4949, 202.6719, 200.2001, 197.3168, 
    200.6131, 203.9207, 209.5309, 213.3633, 206.7827, 200.6213, 212.3189, 
    213.6341,
  224.3351, 228.96, 216.7956, 203.3293, 208.3043, 206.4184, 204.9052, 
    200.841, 202.5047, 210.3928, 215.8454, 211.3881, 210.1291, 214.8932, 
    212.6279,
  224.8806, 223.8548, 216.0774, 207.818, 211.3395, 208.5604, 210.9872, 
    210.7014, 206.8775, 207.6837, 215.9495, 215.3462, 215.0561, 217.3015, 
    210.1821,
  229.1772, 222.578, 214.3955, 214.5207, 212.3458, 213.0423, 215.8699, 
    212.8839, 206.6462, 212.1745, 217.5705, 218.3142, 217.0089, 215.8069, 
    208.1368,
  220.6609, 222.7039, 220.387, 217.3416, 215.7116, 216.0781, 217.464, 
    214.6658, 215.1888, 212.5834, 218.0074, 218.1038, 218.015, 215.5262, 
    210.503,
  211.2481, 207.1433, 211.5451, 209.5107, 205.9095, 211.1144, 210.1912, 
    205.0762, 204.2335, 203.7222, 211.2577, 218.3, 212.156, 204.0822, 199.3422,
  218.8948, 216.8476, 211.1788, 207.3802, 204.4419, 210.4356, 206.6609, 
    204.4505, 201.233, 199.7563, 204.3996, 216.8824, 215.1242, 207.9992, 
    201.6625,
  226.4949, 227.7256, 222.2908, 208.4865, 206.2431, 208.7765, 209.3674, 
    200.2409, 201.3909, 199.1088, 203.788, 212.2643, 213.6926, 205.9067, 
    204.8532,
  235.7563, 228.6491, 228.3249, 222.0111, 212.0638, 212.767, 205.7515, 
    206.0341, 204.6784, 202.3847, 207.7566, 214.4346, 213.1252, 208.8429, 
    206.7551,
  233.9359, 232.2256, 221.5985, 221.8222, 215.2261, 213.75, 215.1533, 
    208.3967, 209.2542, 202.2829, 202.7164, 214.716, 214.0012, 207.8091, 
    208.5286,
  235.8354, 232.9117, 231.6117, 209.1195, 214.6173, 216.761, 215.4538, 
    208.5442, 205.3228, 196.8642, 201.2636, 212.8902, 212.11, 209.6544, 
    209.4944,
  234, 233.1147, 228.3883, 214.7649, 214.4272, 217.7071, 216.5067, 207.6446, 
    201.4438, 203.1513, 206.2836, 214.4158, 214.6634, 214.5166, 208.6644,
  229.8629, 230.032, 219.123, 209.0902, 211.1698, 219.008, 214.3171, 
    211.2468, 208.9812, 203.7362, 207.0816, 214.9002, 216.3704, 215.5912, 
    207.5905,
  234.1893, 226.8762, 217.8045, 213.5324, 199.6167, 218.0968, 211.4614, 
    202.5513, 199.8104, 204.581, 214.8756, 216.2709, 214.8952, 209.2616, 
    211.5804,
  232.558, 228.4198, 223.2227, 216.6477, 209.1044, 214.6432, 210.9713, 
    205.1799, 207.8359, 212.1572, 216.5564, 215.3609, 214.1419, 211.4969, 
    208.2373,
  212.5695, 219.7421, 225.518, 229.7187, 223.7138, 219.4532, 212.4679, 
    210.1175, 214.1785, 215.004, 220.9123, 220.2618, 215.5354, 199.4207, 
    190.5981,
  217.7509, 228.1948, 229.2737, 228.6412, 221.2758, 212.2244, 204.0992, 
    209.6618, 211.7582, 213.9164, 215.2931, 220.7169, 211.6562, 200.9314, 
    189.8644,
  238.162, 237.4924, 234.508, 224.1973, 217.1513, 208.9452, 197.3958, 
    206.1822, 212.3657, 209.39, 211.0719, 217.1942, 210.6842, 199.8513, 
    190.7231,
  235.404, 237.3886, 231.4595, 226.279, 215.694, 213.7038, 196.1227, 
    207.2105, 211.5748, 205.7327, 207.8337, 210.1533, 212.4816, 200.7851, 
    197.9568,
  238.2542, 234.6064, 233.1114, 227.7737, 221.2942, 213.5035, 205.4901, 
    197.8547, 208.9217, 205.9143, 206.6445, 211.6341, 208.8594, 205.9336, 
    203.6784,
  234.8663, 233.2114, 230.4946, 217.8773, 214.0678, 214.6123, 210.2767, 
    198.7276, 204.9754, 210.8624, 210.5428, 209.5601, 206.896, 207.8838, 
    207.2945,
  235.574, 235.9308, 230.8619, 215.4472, 214.2468, 211.2916, 218.1086, 
    199.3482, 205.9832, 213.3548, 205.9422, 210.6038, 208.5642, 208.7299, 
    205.3992,
  235.2131, 228.0023, 213.0514, 211.623, 217.1305, 211.5848, 215.1444, 
    204.5953, 211.8817, 216.3346, 208.8786, 208.8521, 212.9266, 210.4088, 
    205.4365,
  229.9277, 225.7198, 223.8508, 210.9392, 214.3094, 210.0029, 205.8545, 
    201.5981, 208.1699, 215.1829, 208.4784, 210.2333, 215.2056, 212.1291, 
    205.1501,
  226.6371, 221.9119, 218.5688, 215.1913, 214.0703, 208.329, 205.6582, 
    206.1157, 213.5944, 215.1478, 209.5141, 210.3571, 214.6356, 210.3859, 
    208.2981,
  225.0866, 216.9262, 218.09, 227.7016, 226.046, 223.9503, 221.9786, 
    213.3997, 208.6301, 204.4868, 216.1064, 224.8701, 223.7198, 217.4907, 
    209.2862,
  225.8957, 231.3658, 229.6155, 230.1043, 223.7142, 221.131, 216.8322, 
    215.7252, 209.2518, 208.7516, 209.9297, 218.4304, 220.7165, 206.5349, 
    201.0858,
  237.8144, 236.4557, 233.9809, 228.0373, 217.5861, 224.4266, 219.4643, 
    211.5553, 211.6299, 220.6462, 218.7814, 221.5289, 211.8167, 197.8187, 
    193.6013,
  238.6414, 236.3002, 229.5206, 223.661, 216.9468, 218.5693, 214.0423, 
    216.1359, 221.6223, 217.5429, 218.0194, 215.8521, 201.7453, 190.3776, 
    192.4788,
  235.0188, 234.038, 224.5334, 225.913, 216.8543, 210.689, 216.8932, 
    211.0024, 216.6587, 211.1721, 213.04, 205.3427, 189.4746, 188.6588, 
    187.1657,
  233.7581, 232.5193, 232.2119, 225.8887, 215.5888, 215.7229, 214.5012, 
    212.8205, 205.3274, 206.2325, 205.2136, 191.8444, 184.0354, 189.7784, 
    190.4256,
  234.9272, 233.345, 228.7811, 218.9635, 215.8298, 215.5962, 210.0077, 
    209.1453, 201.6459, 202.1578, 192.2809, 188.1146, 182.9648, 186.2234, 
    193.2228,
  231.7224, 230.4512, 209.3414, 219.3763, 214.4621, 211.2073, 207.3579, 
    198.9965, 201.2423, 195.1769, 186.7571, 185.3038, 182.9054, 186.2818, 
    192.6018,
  226.5239, 226.2916, 219.5172, 214.118, 214.1541, 213.081, 200.4678, 
    196.2159, 197.7272, 194.7894, 186.628, 182.8728, 188.307, 188.1506, 
    203.1618,
  225.6515, 225.2392, 221.694, 218.4246, 211.7294, 197.5392, 193.5388, 
    193.9182, 197.667, 191.9845, 189.1278, 188.575, 188.1601, 194.3304, 
    205.1772,
  198.5818, 199.4535, 199.4445, 204.6595, 204.9679, 205.7401, 210.1337, 
    213.4252, 213.7738, 217.3971, 220.2371, 217.9346, 217.3262, 218.6717, 
    217.6244,
  203.2925, 205.692, 206.9702, 213.149, 218.8866, 219.2503, 213.2168, 
    215.6978, 217.8894, 215.7687, 218.3138, 211.58, 209.5369, 217.5184, 
    220.2473,
  214.9951, 226.5777, 234.8065, 230.4368, 222.8588, 218.9368, 222.1124, 
    212.4531, 218.753, 220.2439, 217.9069, 212.8602, 219.1443, 221.6384, 
    222.1774,
  241.3406, 236.0667, 236.1747, 231.4216, 224.4767, 223.4677, 216.9579, 
    219.7161, 221.3241, 220.6831, 220.9982, 218.3048, 222.038, 222.5777, 
    219.8766,
  240.2574, 237.8281, 234.0608, 231.0699, 222.6828, 214.1662, 216.4684, 
    214.0467, 215.2635, 222.6529, 223.2338, 223.909, 223.3152, 220.2619, 
    213.487,
  238.752, 234.2122, 230.8713, 227.5982, 218.7595, 215.3232, 212.8648, 
    219.135, 218.9083, 222.2204, 223.0905, 222.3448, 217.0364, 213.6635, 
    204.4164,
  238.7999, 237.6502, 213.3151, 220.3807, 218.5928, 214.8025, 216.1408, 
    221.9441, 220.4107, 220.2265, 218.4393, 212.0207, 208.1512, 205.9273, 
    200.3329,
  238.2474, 234.1961, 214.3372, 219.3093, 216.394, 218.3885, 218.7665, 
    218.511, 216.7672, 209.7567, 207.9309, 203.9929, 201.8003, 204.2004, 
    207.3892,
  232.6276, 228.1061, 222.9386, 211.7939, 204.4367, 204.0617, 205.9434, 
    207.3038, 205.1047, 203.3992, 198.8888, 200.9865, 200.6856, 209.2849, 
    217.4491,
  227.8426, 228.0059, 214.9859, 200.5283, 198.1785, 196.6019, 196.8553, 
    200.7732, 196.6228, 197.2652, 193.1384, 199.4666, 207.209, 215.3352, 
    221.3738,
  211.0041, 215.1125, 214.723, 212.4152, 213.6503, 218.8347, 218.6894, 
    214.232, 211.7363, 214.1539, 210.5261, 209.816, 207.7708, 204.81, 205.1295,
  205.2113, 209.3939, 207.8157, 208.267, 208.8583, 213.579, 213.6861, 
    211.4963, 211.734, 212.1633, 212.3531, 212.9538, 214.6157, 209.7497, 
    211.6445,
  197.8654, 198.8638, 199.4585, 205.1395, 210.808, 213.047, 215.9223, 
    212.8237, 216.1918, 213.3446, 214.5115, 209.6569, 211.2321, 215.167, 
    217.9414,
  190.272, 189.0147, 198.0498, 207.1691, 209.9631, 213.8486, 211.8955, 
    218.4715, 220.7319, 218.0138, 208.8933, 212.0329, 209.3621, 217.9489, 
    215.0079,
  197.188, 205.4528, 213.717, 220.1078, 217.6106, 213.1118, 216.5845, 
    211.5357, 210.8194, 214.9223, 214.4998, 215.4389, 214.0985, 217.7203, 
    219.8879,
  210.9476, 223.7094, 229.3097, 228.3599, 223.7901, 215.6615, 210.6606, 
    214.3161, 215.8788, 213.816, 217.0736, 215.9182, 217.2719, 218.6898, 
    215.8359,
  225.9382, 236.558, 236.4209, 224.0655, 219.1909, 212.1131, 211.7257, 
    209.9121, 213.0345, 221.1064, 215.7789, 212.5575, 213.7672, 219.7795, 
    217.6836,
  238.6289, 239.8914, 232.2345, 223.2561, 214.7477, 214.0352, 219.861, 
    224.1332, 222.7376, 220.8682, 220.0655, 216.6005, 213.4707, 216.6702, 
    215.8206,
  229.3635, 234.0035, 227.7668, 217.8601, 214.4596, 222.8991, 225.8064, 
    225.1497, 222.7309, 220.3339, 220.1337, 218.8023, 214.5488, 213.5363, 
    211.9077,
  222.1114, 230.6321, 220.9616, 215.9385, 221.7896, 227.6839, 227.4009, 
    225.8825, 221.2826, 216.0051, 220.1157, 213.146, 210.2724, 211.1239, 
    210.2942,
  222.0731, 223.0637, 222.1822, 226.7214, 220.7724, 223.4543, 211.3113, 
    199.147, 190.1516, 189.3971, 189.0133, 193.7132, 199.8348, 206.8716, 
    214.0725,
  214.3421, 216.9222, 223.443, 223.1955, 220.7172, 214.5028, 205.3333, 
    198.4571, 191.7567, 194.0879, 193.6264, 197.9292, 207.724, 209.1894, 
    212.4088,
  216.2565, 218.1571, 216.4139, 212.2841, 206.4727, 199.2342, 198.42, 
    191.6404, 193.9168, 196.3484, 198.7849, 206.7669, 209.1385, 215.316, 
    210.5942,
  212.9706, 213.8121, 206.0988, 203.2252, 194.2648, 193.6432, 189.3434, 
    194.3247, 194.2243, 202.072, 208.8757, 213.2673, 211.8521, 214.3781, 
    215.5434,
  225.4324, 209.4492, 205.1291, 193.838, 188.5306, 187.8535, 197.5581, 
    200.0213, 205.0357, 214.8129, 221.4729, 216.0879, 217.7319, 218.966, 
    220.2243,
  205.015, 196.9086, 191.1211, 190.2399, 191.939, 197.8336, 208.5761, 
    221.4567, 224.4263, 223.7997, 223.9862, 223.3705, 218.266, 218.5153, 
    216.9231,
  188.3185, 186.0518, 190.7013, 193.4623, 205.5201, 221.4278, 227.8981, 
    227.6125, 224.7054, 220.3469, 213.7431, 216.6776, 218.3475, 216.436, 
    217.4565,
  186.3064, 194.3729, 198.9139, 211.0256, 226.2996, 223.2341, 227.2909, 
    225.5352, 224.2663, 221.32, 220.4718, 219.3693, 219.762, 219.35, 213.2854,
  189.8851, 196.3016, 215.2556, 222.5934, 222.3289, 226.4389, 224.3979, 
    221.2502, 220.1165, 215.9955, 217.1388, 209.6625, 209.8579, 213.1699, 
    214.4704,
  196.9375, 210.6537, 217.9607, 225.025, 226.5114, 223.4388, 220.9536, 
    219.5308, 218.5926, 218.9305, 218.9712, 211.8275, 212.2799, 216.3695, 
    211.9323,
  239.583, 240.9814, 232.1663, 226.6982, 220.7078, 218.321, 220.7472, 
    221.4798, 218.5379, 219.7009, 217.3344, 215.1808, 214.6494, 212.4756, 
    208.9075,
  238.0891, 231.7826, 218.2886, 211.7831, 210.1019, 204.4226, 203.8256, 
    204.4866, 208.8999, 210.7814, 215.8965, 214.0794, 215.6675, 210.9485, 
    209.5656,
  232.9347, 220.9759, 211.067, 206.4774, 204.5729, 201.2241, 202.3795, 
    203.2028, 204.9898, 207.2632, 209.0526, 208.8824, 211.815, 210.1067, 
    208.4245,
  229.4143, 219.207, 204.8191, 204.7791, 204.0461, 206.4382, 201.4924, 
    203.0791, 199.122, 202.6645, 214.2892, 219.8453, 212.388, 202.0043, 
    201.5336,
  221.6393, 209.2194, 201.7382, 205.2874, 205.2954, 208.5147, 209.6004, 
    205.6748, 212.853, 213.7621, 208.961, 209.1488, 205.0914, 205.582, 
    205.4238,
  212.5311, 195.7263, 202.2771, 205.4727, 208.1357, 206.6543, 211.8932, 
    216.135, 220.7355, 217.2187, 214.8682, 209.3407, 208.4235, 207.8171, 
    207.0221,
  197.2172, 194.4457, 199.9277, 203.9722, 213.9184, 221.7914, 227.024, 
    228.941, 227.7281, 218.3741, 213.9945, 208.6626, 208.01, 207.032, 207.8856,
  189.2079, 196.887, 204.4931, 215.9218, 224.1335, 227.7044, 228.5807, 
    228.5827, 227.8039, 226.2011, 222.7621, 215.8385, 214.2863, 212.9105, 
    212.7821,
  193.8278, 204.0937, 213.0159, 216.4493, 217.8655, 217.7227, 223.1002, 
    223.9275, 223.7586, 222.8101, 221.2495, 219.7973, 217.4764, 218.7453, 
    213.934,
  200.4527, 213.5346, 218.738, 217.37, 216.7138, 215.1113, 216.0496, 
    224.0653, 222.4626, 221.8518, 219.8675, 213.7913, 214.7935, 215.4741, 
    213.2564,
  192.2632, 199.6097, 204.2118, 206.9935, 212.3779, 212.6634, 218.2812, 
    223.449, 222.8922, 219.5968, 217.1295, 216.958, 215.7059, 214.4248, 
    219.3409,
  207.4669, 213.0331, 215.6661, 215.8018, 222.2014, 218.088, 220.8842, 
    221.3464, 219.4068, 216.7935, 215.5365, 211.9586, 209.7153, 208.968, 
    205.4491,
  215.1318, 218.0888, 216.0267, 216.9159, 222.1776, 216.2337, 220.798, 
    224.4591, 222.8175, 223.0934, 220.1383, 216.5042, 210.222, 208.1324, 
    202.8758,
  222.4617, 219.5805, 218.6223, 219.1794, 218.2465, 224.4974, 217.2017, 
    226.789, 226.8401, 223.5374, 224.8038, 220.1367, 213.3015, 209.1939, 
    200.1295,
  212.884, 208.2157, 214.1752, 216.5359, 218.056, 222.2466, 220.9613, 
    219.6197, 217.1853, 224.9368, 224.2143, 223.3469, 212.4997, 211.4682, 
    203.2456,
  205.7159, 202.7924, 208.5292, 221.5565, 222.3524, 223.6889, 219.6283, 
    223.862, 225.2324, 226.7644, 225.2128, 214.4657, 206.1467, 203.106, 
    200.455,
  207.3617, 206.4875, 211.136, 214.6031, 221.6796, 220.9933, 222.2104, 
    222.7068, 224.549, 225.8874, 226.2092, 201.1325, 200.7298, 198.1329, 
    199.7361,
  216.6571, 215.1249, 215.5536, 212.8004, 212.9808, 212.6979, 221.1189, 
    223.2072, 224.9032, 225.3307, 221.8698, 199.6447, 198.0999, 196.6084, 
    199.9774,
  227.4684, 215.0289, 213.3013, 211.3328, 209.39, 210.822, 219.2466, 
    223.1906, 223.9727, 224.0284, 220.2872, 199.9114, 195.6517, 196.1228, 
    198.5151,
  212.0807, 217.0078, 210.9057, 209.4094, 210.6501, 212.7656, 214.45, 
    223.2598, 223.8696, 223.4114, 217.6195, 200.9137, 199.6899, 203.6006, 
    209.3575,
  240.4457, 235.9328, 233.8991, 226.7637, 219.2782, 213.5451, 212.8415, 
    210.7612, 204.2511, 201.4448, 208.9937, 212.2206, 219.4067, 219.0872, 
    223.6749,
  235.4531, 232.9631, 232.1729, 226.5804, 218.7306, 215.6202, 215.1177, 
    207.4467, 200.0753, 196.8956, 205.4597, 212.6769, 219.8919, 221.92, 
    222.8052,
  229.662, 229.2913, 225.9825, 220.359, 217.1777, 210.1755, 207.843, 
    197.8113, 192.1469, 195.1385, 208.134, 217.0483, 224.8977, 223.9298, 
    221.9556,
  224.674, 218.7701, 217.5324, 216.064, 206.9325, 200.5931, 193.8322, 
    193.322, 193.6083, 201.8421, 208.6144, 219.7953, 226.2486, 224.5429, 
    214.2851,
  219.2643, 213.8822, 211.8801, 204.4863, 204.946, 194.5538, 195.4158, 
    196.1398, 195.8335, 209.0358, 216.2815, 223.7648, 226.5791, 215.652, 
    205.1192,
  219.9347, 212.345, 209.4993, 207.8048, 208.6965, 204.8164, 198.17, 201.541, 
    205.7977, 210.1325, 218.7294, 227.8684, 218.0564, 205.1866, 205.4604,
  224.7894, 216.5288, 209.2365, 213.7065, 210.1904, 206.14, 207.3984, 
    207.4622, 209.852, 217.5434, 226.3554, 222.2331, 215.0557, 201.52, 
    204.8674,
  229.8076, 216.3709, 214.5057, 213.2731, 213.0191, 213.7628, 216.4154, 
    221.3781, 221.4958, 226.0279, 227.2896, 218.9399, 207.5572, 198.5019, 
    204.7739,
  236.6472, 223.1279, 214.2779, 210.9723, 211.295, 211.6384, 214.4206, 
    222.2864, 223.841, 226.1396, 215.7845, 209.8311, 198.0552, 196.3316, 
    207.7278,
  230.2661, 219.1377, 211.3073, 214.3971, 214.6891, 220.4655, 221.5174, 
    223.5888, 225.2531, 222.049, 212.5276, 207.8285, 208.9349, 213.9078, 
    216.1398,
  226.455, 223.7621, 224.1277, 224.5548, 226.8165, 220.4225, 210.6919, 
    210.424, 208.9924, 214.383, 216.0986, 204.6591, 192.9572, 189.2671, 
    188.367,
  216.7503, 220.3624, 224.2834, 226.5397, 226.0937, 221.6906, 207.5337, 
    207.3108, 208.4995, 204.3306, 196.409, 189.6473, 190.8267, 188.4646, 
    202.261,
  219.7033, 221.0541, 223.0823, 227.7842, 223.8831, 217.3424, 206.3095, 
    194.4423, 193.4865, 194.3182, 190.2369, 190.8112, 197.8022, 212.0722, 
    229.2041,
  222.1355, 223.5345, 229.5964, 226.3389, 220.5065, 224.066, 197.6353, 
    190.1848, 189.2164, 187.4866, 189.4878, 199.156, 218.5795, 228.459, 
    225.9783,
  230.7126, 226.4826, 235.6084, 222.4415, 219.2988, 214.781, 200.6021, 
    184.8239, 182.0161, 187.1562, 192.1244, 208.223, 224.1435, 225.6683, 
    218.2727,
  241.0979, 224.2644, 222.6034, 218.1281, 216.1895, 215.8382, 207.4493, 
    187.6015, 180.0185, 185.6359, 190.1472, 216.1411, 224.7434, 225.8251, 
    223.7148,
  238.9707, 223.2717, 216.1366, 212.5675, 214.3426, 215.5111, 216.4364, 
    191.5936, 183.7115, 190.814, 202.5434, 220.6899, 224.5458, 222.0512, 
    220.8077,
  240.8967, 221.4279, 214.4814, 210.3796, 210.2324, 212.6087, 216.1009, 
    216.9514, 200.8337, 202.7896, 214.1307, 216.1945, 213.8785, 212.2603, 
    209.5013,
  235.1634, 224.4166, 217.2398, 210.9602, 210.261, 212.0721, 215.1708, 
    224.4232, 217.4882, 212.6871, 218.6636, 213.0975, 213.894, 213.3175, 
    212.6868,
  228.1866, 225.7275, 215.7336, 214.2132, 210.3295, 216.2896, 219.0868, 
    224.9969, 219.8671, 219.1545, 210.8512, 214.4246, 216.2128, 216.4776, 
    219.6658,
  205.3354, 204.8205, 209.4098, 222.996, 228.9578, 229.4076, 225.6271, 
    220.9524, 211.9654, 211.2488, 217.0205, 217.229, 219.5693, 217.5023, 
    204.7886,
  205.4658, 211.5223, 221.1691, 227.8409, 232.4546, 229.3594, 224.6545, 
    221.0524, 213.3839, 209.5108, 215.2376, 216.0513, 220.3429, 219.4498, 
    220.0364,
  211.1997, 221.0112, 229.5426, 232.7094, 230.5896, 228.6913, 224.675, 
    214.9996, 208.0366, 200.6371, 208.5707, 212.0871, 215.4471, 216.8276, 
    217.1167,
  218.1727, 232.3627, 234.3568, 229.8445, 227.4299, 229.9739, 219.9677, 
    216.9938, 206.9393, 199.5299, 207.2362, 209.5184, 212.007, 214.7498, 
    216.5658,
  233.7107, 240.9121, 231.6652, 226.817, 223.6925, 215.5186, 217.57, 
    214.5094, 201.2138, 200.9044, 207.158, 206.6002, 207.3752, 211.5674, 
    214.4332,
  244.3594, 235.7626, 231.6442, 219.3754, 206.5949, 207.6926, 210.348, 
    215.8182, 203.3574, 200.5443, 210.6718, 206.5556, 205.1105, 205.3737, 
    211.5316,
  230.6675, 225.8064, 220.9777, 212.1679, 206.9401, 201.2314, 208.8027, 
    213.6882, 206.6165, 207.2459, 212.4193, 205.6018, 204.056, 203.1955, 
    204.8997,
  244.3157, 239.0143, 230.3249, 224.0439, 215.0963, 213.1403, 212.6331, 
    215.8842, 204.2386, 210.3732, 210.5877, 205.8736, 207.1466, 209.2217, 
    205.2655,
  238.4354, 231.5023, 230.2888, 228.5063, 218.8556, 216.9601, 212.9727, 
    217.7413, 202.3941, 212.8118, 207.2892, 207.844, 206.9593, 207.2349, 
    208.5753,
  234.2861, 228.6725, 228.2104, 227.6684, 227.8868, 219.8043, 215.7671, 
    215.7143, 205.9769, 213.0565, 207.8581, 209.3532, 206.9574, 209.0771, 
    208.6772,
  189.0663, 187.7963, 190.6548, 207.8731, 223.952, 230.1846, 227.865, 
    226.8217, 226.8935, 217.0555, 206.6003, 207.6149, 216.7972, 216.7038, 
    218.3084,
  185.8498, 191.2254, 204.2708, 224.7363, 231.9134, 231.3018, 227.1691, 
    226.1952, 224.5117, 219.4964, 207.065, 209.4756, 218.0284, 217.6447, 
    220.438,
  188.8398, 204.5898, 228.0796, 234.1432, 234.1981, 231.3235, 228.3302, 
    222.4405, 223.0219, 217.7483, 210.1935, 207.5295, 216.0989, 218.971, 
    220.48,
  200.392, 226.514, 238.2897, 238.8881, 232.1096, 232.6681, 220.7524, 
    226.2133, 222.749, 214.3093, 210.0949, 206.1535, 210.8516, 217.0957, 
    217.7695,
  216.5974, 222.1222, 226.6511, 229.0008, 231.7587, 218.0866, 216.3886, 
    216.8223, 214.6785, 217.663, 212.2597, 208.8247, 207.3918, 212.553, 
    213.9301,
  220.6331, 236.6494, 237.1842, 222.7778, 221.4142, 214.7813, 218.7778, 
    219.9398, 219.178, 214.8897, 212.9588, 211.4683, 208.3341, 210.0147, 
    209.0125,
  226.9085, 232.2406, 231.7686, 229.2781, 225.7495, 220.9447, 217.7051, 
    219.7355, 219.8006, 217.8076, 215.1718, 211.7102, 208.1539, 208.4334, 
    209.7989,
  233.0779, 230.4257, 228.1345, 224.9982, 220.6733, 220.9524, 220.3749, 
    222.3723, 216.8952, 215.6545, 210.0126, 208.4455, 208.0343, 208.034, 
    208.9177,
  230.7591, 229.7335, 224.8817, 222.6496, 220.3637, 219.3743, 222.2731, 
    220.6942, 216.6858, 212.2426, 208.6194, 205.8773, 203.7523, 210.3128, 
    206.6286,
  228.0977, 226.3445, 225.2802, 221.568, 220.4291, 220.9762, 218.6628, 
    218.5581, 216.7603, 213.0732, 207.8752, 200.8416, 202.149, 209.0389, 
    210.5874,
  236.2702, 231.6741, 228.8562, 229.3549, 229.6035, 230.8561, 227.9542, 
    225.2523, 222.5036, 219.241, 217.4719, 215.6816, 209.9411, 203.5383, 
    203.474,
  231.0381, 228.3839, 229.5871, 228.881, 231.1015, 228.3773, 225.2018, 
    224.0764, 223.3584, 218.3154, 215.9084, 208.4789, 206.5434, 206.4031, 
    207.0399,
  221.9149, 225.7595, 228.572, 228.558, 230.547, 223.941, 224.8536, 220.9946, 
    217.6937, 216.3658, 210.5712, 202.7602, 202.3805, 207.1345, 206.7608,
  218.1989, 224.7915, 226.5567, 229.4388, 225.0952, 223.9693, 220.0705, 
    224.2037, 218.53, 214.458, 212.2202, 201.3894, 207.8869, 209.289, 205.6318,
  215.375, 221.0231, 224.9027, 230.4999, 225.0543, 221.0771, 220.12, 
    218.1842, 216.9114, 216.2475, 210.7615, 205.6417, 203.1191, 206.5906, 
    205.7374,
  216.1411, 224.7542, 227.1121, 226.0898, 222.3361, 219.7684, 217.6167, 
    217.9378, 218.1969, 213.9035, 210.1515, 205.9918, 205.7131, 211.2835, 
    203.739,
  226.9671, 228.1846, 225.9206, 223.0214, 219.8855, 219.0339, 215.9575, 
    216.1938, 216.9563, 214.7961, 208.9658, 207.1667, 208.9569, 208.8921, 
    206.744,
  228.9657, 227.2202, 225.4281, 222.1926, 218.3553, 216.5654, 215.1459, 
    218.8732, 217.4189, 216.0653, 210.3478, 209.6624, 213.2852, 213.1415, 
    208.7056,
  227.6605, 225.1839, 226.4165, 221.2732, 217.0484, 215.5524, 218.4494, 
    219.3187, 218.7952, 216.3326, 213.6326, 210.9542, 210.0257, 212.3222, 
    213.337,
  225.9254, 228.3143, 225.1857, 220.7538, 217.2746, 216.6169, 216.0199, 
    217.8725, 219.3579, 219.3956, 215.4208, 214.8285, 213.8919, 210.0605, 
    208.0416,
  231.5619, 225.778, 229.9298, 229.8941, 227.81, 225.7989, 223.0863, 
    220.3149, 216.144, 213.9912, 211.4413, 211.0699, 211.0294, 205.5719, 
    204.2776,
  227.9218, 227.351, 229.5474, 227.321, 226.4352, 224.8017, 220.1498, 
    220.3858, 215.6277, 213.5964, 211.9162, 213.0313, 209.3006, 205.9993, 
    206.3805,
  226.8252, 227.9652, 228.3152, 226.5557, 226.9439, 220.381, 220.7993, 
    212.7015, 215.1843, 213.7492, 212.6675, 211.5967, 209.5078, 206.1443, 
    206.4711,
  227.6431, 228.4005, 228.4767, 227.0081, 222.9065, 221.1246, 217.0004, 
    214.2162, 216.9812, 213.5777, 212.0457, 212.3191, 208.3949, 205.3803, 
    204.0422,
  230.9759, 230.0893, 229.0965, 223.8952, 219.7087, 216.1886, 217.0014, 
    216.6974, 216.3035, 215.7579, 208.6967, 209.8423, 209.667, 203.9085, 
    201.6755,
  229.5706, 227.2094, 225.9878, 223.0608, 218.4228, 214.7005, 211.6472, 
    217.0275, 219.272, 216.004, 212.2504, 208.9051, 210.0362, 203.9743, 
    201.7547,
  229.3161, 228.1484, 225.0571, 222.2077, 216.744, 214.5759, 215.061, 
    216.9416, 217.5192, 216.2056, 213.1663, 209.1218, 212.4824, 208.5713, 
    202.0022,
  228.1623, 225.8416, 224.2074, 220.8289, 217.7254, 218.0962, 217.2531, 
    218.2584, 218.4733, 216.5394, 211.0525, 208.5189, 206.1047, 207.1704, 
    210.9856,
  227.5606, 227.3609, 223.5947, 221.0637, 217.3825, 218.5515, 216.9239, 
    214.7637, 214.441, 212.662, 209.3824, 204.4213, 201.2425, 206.281, 
    212.3536,
  230.741, 226.2505, 223.7791, 222.286, 220.4854, 217.4796, 215.1461, 
    213.4611, 210.8371, 208.8579, 208.8563, 205.7603, 203.1136, 208.8192, 
    213.4778,
  240.6207, 231.3828, 231.9231, 228.2804, 226.0684, 222.0991, 218.1428, 
    218.7553, 213.9417, 210.9549, 209.9278, 208.3599, 214.6451, 211.231, 
    205.2709,
  230.89, 235.0695, 230.2151, 227.1026, 223.4028, 220.2887, 213.1876, 
    217.3276, 218.6752, 210.353, 209.3312, 214.478, 215.865, 216.0209, 
    210.5401,
  234.6486, 231.0927, 229.9498, 225.5289, 222.1904, 219.9542, 217.7373, 
    205.9829, 210.0182, 209.8395, 214.5538, 216.8163, 216.0058, 212.3523, 
    208.5404,
  230.8552, 232.0472, 228.4763, 224.6836, 220.9627, 221.6546, 215.999, 
    213.9941, 213.2914, 209.7421, 212.7971, 215.1627, 215.7881, 211.646, 
    208.9312,
  231.6435, 229.8443, 227.3658, 223.8007, 220.9352, 216.7605, 215.1271, 
    213.2371, 213.8739, 212.3447, 212.0123, 213.6851, 211.2207, 209.3148, 
    205.0513,
  237.7118, 229.2269, 226.4643, 223.3558, 221.7098, 216.5831, 210.8529, 
    209.9205, 212.5195, 210.9345, 211.6777, 214.321, 209.7697, 207.9968, 
    206.2176,
  233.6429, 229.4317, 225.621, 225.4959, 223.2296, 215.809, 210.362, 
    211.5758, 207.6388, 209.4863, 213.6897, 211.7564, 207.0936, 206.6877, 
    205.0313,
  232.8828, 229.5423, 226.8939, 225.711, 222.7349, 213.376, 213.1708, 
    211.5718, 210.8878, 207.8383, 210.2057, 209.0491, 208.0143, 209.451, 
    208.8755,
  233.1717, 229.1425, 227.1885, 224.8238, 221.9138, 215.1091, 213.8085, 
    213.4072, 209.7042, 209.5774, 212.0697, 209.5892, 216.331, 216.1381, 
    213.9857,
  233.4263, 231.265, 227.4861, 226.0911, 220.6244, 217.2237, 215.7048, 
    214.8031, 212.5541, 211.1702, 212.2349, 211.0477, 217.364, 213.6738, 
    215.4846,
  241.7833, 236.3028, 232.8217, 227.2216, 225.0049, 221.9755, 217.3262, 
    214.3236, 208.1986, 210.4294, 205.3348, 206.8421, 211.7626, 219.0785, 
    213.7913,
  237.3904, 232.1352, 228.8211, 225.3851, 223.6473, 221.8121, 214.9915, 
    214.3369, 211.9464, 209.6305, 206.6121, 205.2426, 211.6398, 209.0863, 
    217.8465,
  232.869, 231.9451, 227.1778, 223.9242, 222.8797, 218.693, 214.7677, 
    206.6136, 207.0297, 207.7282, 205.7065, 207.8087, 212.3728, 210.0044, 
    211.8726,
  236.009, 230.5449, 226.9095, 223.5545, 221.3558, 214.737, 215.5629, 
    212.1537, 201.8686, 201.5063, 203.4132, 210.3447, 215.0143, 210.1309, 
    211.105,
  232.5709, 229.0312, 225.9835, 223.491, 218.346, 207.3271, 208.7516, 
    211.4218, 203.8304, 203.6785, 204.0104, 206.7275, 214.4888, 211.4755, 
    210.8797,
  234.2854, 228.6971, 225.4477, 222.4491, 216.0997, 205.1227, 200.7823, 
    201.6965, 203.966, 204.2055, 205.315, 206.084, 212.8597, 215.0583, 
    212.3061,
  234.4076, 230.1508, 228.6169, 221.1871, 213.8953, 205.7246, 202.0245, 
    199.5946, 205.5811, 207.6221, 205.3208, 217.4214, 215.6406, 215.8367, 
    215.4494,
  233.4043, 229.6886, 227.2356, 222.6302, 216.4616, 210.6923, 204.0163, 
    201.3356, 204.6434, 208.1654, 208.3552, 218.1385, 212.4942, 217.5944, 
    217.5707,
  233.3437, 229.7491, 227.3567, 222.9921, 217.9675, 211.8129, 206.5038, 
    203.0378, 206.7502, 211.025, 211.6236, 212.0072, 223.4954, 219.9234, 
    219.0208,
  238.3315, 233.5512, 228.52, 227.2717, 220.5416, 215.2054, 208.6886, 
    206.2468, 206.9517, 213.0675, 213.4357, 206.0041, 221.1102, 223.8839, 
    219.812,
  247.1855, 237.1736, 230.9689, 227.1533, 224.8666, 219.8089, 215.7499, 
    212.9151, 208.8975, 205.7041, 215.3627, 222.1007, 217.5473, 220.1398, 
    219.8653,
  235.6483, 231.6397, 229.1231, 228.3934, 223.4273, 215.3681, 209.1436, 
    211.3083, 211.3688, 205.6775, 213.2171, 222.3047, 218.4301, 218.4143, 
    219.1898,
  233.812, 229.1741, 226.475, 221.8522, 218.2374, 213.6617, 206.881, 
    203.3322, 209.6413, 207.4526, 206.0325, 215.7719, 218.3555, 216.1276, 
    216.8572,
  232.4849, 227.6508, 226.742, 222.2089, 215.1147, 211.2968, 202.7569, 
    203.08, 212.5444, 208.4311, 202.3134, 213.8051, 220.9808, 214.5603, 
    218.7986,
  231.6362, 227.5661, 227.5726, 223.7049, 214.5713, 210.5175, 202.4571, 
    199.6688, 204.8576, 209.7724, 203.7443, 208.8172, 213.2381, 215.3402, 
    218.1244,
  231.4345, 227.5716, 229.4234, 224.7126, 219.2972, 210.2629, 202.863, 
    207.341, 208.4641, 204.4191, 200.7039, 206.0158, 210.6038, 214.0351, 
    215.9397,
  230.8819, 230.6953, 228.053, 227.4306, 220.3772, 210.8624, 209.2308, 
    216.6171, 212.9527, 212.0469, 202.6585, 207.6008, 208.8391, 211.0112, 
    217.2872,
  230.3817, 228.9207, 228.2374, 228.009, 223.6791, 211.7218, 211.3244, 
    222.5364, 219.7982, 218.8433, 204.5232, 209.9474, 208.258, 211.4971, 
    215.7463,
  230.1292, 228.4999, 227.9261, 225.9666, 222.622, 212.2015, 209.1969, 
    219.2978, 221.4592, 215.1059, 204.8417, 207.7111, 208.4628, 211.2395, 
    215.1122,
  230.4373, 228.3165, 227.6166, 225.2956, 220.5806, 214.9546, 208.0713, 
    204.9778, 203.126, 203.4341, 205.444, 208.7615, 210.6445, 211.4039, 
    215.369,
  210.9859, 209.0942, 215.7616, 221.839, 225.4461, 221.6109, 213.7504, 
    213.1562, 210.2716, 211.3104, 215.4229, 223.193, 227.9371, 232.5877, 
    218.2008,
  204.3748, 211.7374, 221.0268, 226.7803, 222.7231, 213.6038, 210.9854, 
    211.3954, 211.3795, 209.6823, 212.3467, 222.1862, 226.2722, 220.8046, 
    211.4448,
  201.7142, 214.6877, 226.0302, 227.1544, 218.5021, 210.653, 202.6136, 
    206.9725, 209.252, 202.4084, 213.5247, 219.0382, 224.6202, 215.9122, 
    203.7632,
  207.7872, 222.8659, 227.8482, 227.7992, 215.6775, 207.3998, 211.9518, 
    208.8286, 208.945, 207.904, 212.6114, 218.9083, 220.3216, 210.8955, 
    209.8369,
  220.0807, 226.0784, 228.1912, 228.0181, 208.9211, 206.9981, 205.0788, 
    196.1023, 212.8332, 217.0136, 215.0443, 217.7093, 213.2256, 207.5999, 
    215.3236,
  225.1764, 227.6687, 227.9024, 226.8801, 210.1837, 206.905, 214.8772, 
    220.791, 217.8894, 216.1524, 216.9949, 213.5658, 210.7888, 208.9549, 
    216.0846,
  229.3409, 228.062, 227.4339, 225.4407, 212.2672, 219.778, 228.371, 
    218.1447, 213.2197, 212.4569, 211.7268, 203.5897, 204.1302, 206.3992, 
    211.0612,
  228.611, 228.6537, 226.0733, 210.3668, 205.6517, 209.5777, 216.1083, 
    211.9928, 211.8177, 210.0946, 206.8, 204.4452, 200.0713, 210.4742, 
    209.1929,
  228.6066, 225.1695, 212.284, 206.1761, 205.4841, 206.0928, 207.8786, 
    211.1905, 203.0598, 204.756, 201.8857, 204.4486, 200.4737, 204.0758, 
    208.3694,
  229.8139, 219.2335, 208.8163, 206.493, 205.5705, 209.6048, 207.0402, 
    206.312, 203.1693, 202.7235, 201.1614, 205.4839, 203.565, 204.919, 208.197,
  213.2373, 214.132, 211.1348, 213.0421, 217.0403, 219.8755, 220.4068, 
    219.5668, 222.845, 228.1831, 221.1464, 223.962, 229.0872, 235.4131, 
    214.5815,
  209.6616, 209.7065, 209.4664, 213.674, 218.4324, 218.162, 220.5663, 
    222.0298, 218.8931, 216.4696, 219.311, 226.1541, 232.5364, 231.2745, 
    211.4991,
  202.5523, 200.8199, 208.2617, 214.0445, 222.989, 222.4247, 216.9622, 
    215.0042, 213.0946, 226.7107, 227.969, 223.6619, 232.0784, 227.4648, 
    206.5574,
  193.5884, 200.2625, 211.8401, 220.6575, 228.8938, 223.4897, 227.433, 
    228.5904, 211.4458, 220.7359, 223.7514, 224.4166, 232.48, 221.5208, 
    208.9325,
  198.7116, 215.7977, 224.1859, 226.7412, 225.5772, 208.0179, 213.9202, 
    207.129, 224.5865, 228.5891, 226.0777, 226.6771, 229.7599, 213.6526, 
    210.6634,
  223.2496, 226.8834, 227.1697, 227.4057, 215.1972, 206.7851, 211.2007, 
    222.9944, 218.0025, 227.6266, 231.5293, 231.4414, 220.3948, 210.429, 
    216.294,
  228.0991, 228.0924, 227.0806, 224.3987, 213.5464, 214.7932, 213.3513, 
    219.7507, 220.407, 231.749, 230.814, 223.3108, 213.3141, 212.3636, 
    215.1471,
  230.6999, 230.6018, 226.8853, 219.133, 210.8235, 216.3231, 212.1337, 
    216.1209, 225.3626, 228.4352, 221.1592, 211.4538, 210.6834, 216.0412, 
    222.873,
  236.5971, 221.7711, 207.5591, 206.5909, 208.6271, 213.31, 207.2582, 
    214.9127, 221.2161, 213.2378, 204.4866, 204.2484, 214.4635, 220.8382, 
    224.5087,
  236.6501, 208.3403, 207.0698, 212.2627, 211.558, 208.6376, 214.2631, 
    216.4745, 204.6175, 201.5473, 200.226, 209.9937, 218.6824, 219.4424, 
    225.2406,
  203.7457, 218.2937, 225.2027, 230.4531, 230.2181, 232.4099, 229.1558, 
    224.6168, 223.981, 225.0929, 232.0989, 231.1916, 239.3402, 235.386, 
    228.335,
  192.426, 205.3578, 220.337, 220.2266, 223.4544, 223.1678, 220.4244, 
    223.125, 227.8533, 231.8934, 234.9728, 231.5438, 237.2495, 230.7636, 
    212.8038,
  188.9259, 195.7003, 204.4789, 213.1307, 215.7975, 223.0928, 220.0547, 
    223.3659, 229.2992, 231.909, 233.0383, 231.3192, 236.6853, 221.9878, 
    200.0142,
  189.629, 193.9517, 201.5426, 208.1432, 211.1957, 220.5137, 226.0398, 
    229.4085, 233.5707, 233.3581, 231.2729, 232.1257, 228.1195, 208.9495, 
    202.864,
  196.7724, 199.776, 205.6162, 209.5213, 216.4095, 220.2458, 232.2705, 
    223.5724, 228.3141, 237.0014, 233.2941, 228.5083, 218.7133, 212.2117, 
    213.78,
  207.6611, 213.9254, 220.7713, 221.5681, 226.883, 225.3976, 221.9807, 
    228.8108, 237.0869, 237.1185, 234.0771, 225.6946, 218.118, 219.7881, 
    217.7732,
  224.2646, 224.6653, 225.6839, 228.1309, 225.422, 221.2342, 219.808, 
    224.6714, 236.0761, 236.395, 229.0268, 221.7818, 224.1183, 217.6338, 
    217.8774,
  225.3976, 224.6386, 231.3557, 231.3295, 217.7152, 216.3774, 222.7852, 
    230.9123, 235.5681, 232.2047, 224.6013, 222.739, 220.3784, 215.8074, 
    214.0729,
  240.2464, 226.3723, 224.8843, 214.1663, 222.9687, 221.3297, 230.7922, 
    225.8794, 232.2522, 226.3319, 222.6556, 223.5463, 214.9113, 214.5702, 
    219.2216,
  236.8118, 213.2847, 211.1399, 216.979, 229.2968, 225.4006, 235.6525, 
    233.1236, 228.1358, 223.5305, 214.6175, 214.4284, 212.6275, 220.4531, 
    230.2983,
  243.8565, 239.6293, 232.1072, 218.9565, 209.0144, 220.683, 233.697, 
    240.3847, 233.993, 227.6685, 229.4752, 233.0442, 235.6497, 236.3769, 
    237.3465,
  235.4369, 236.4509, 227.1471, 210.4055, 205.8542, 220.3476, 235.1062, 
    238.6224, 233.5772, 228.9285, 230.1977, 234.057, 234.1379, 234.6812, 
    236.0764,
  234.5907, 229.2842, 222.9052, 208.1306, 206.306, 212.8472, 232.6854, 
    231.5639, 226.2087, 227.6943, 229.3104, 233.9506, 234.542, 234.0641, 
    231.7209,
  225.8043, 227.0661, 213.0736, 198.4529, 198.3759, 210.79, 228.6937, 
    229.7277, 226.5499, 227.8387, 235.0162, 234.8113, 232.7793, 227.6284, 
    231.5097,
  214.0889, 212.9894, 198.9506, 192.1756, 190.366, 195.8284, 211.6333, 
    223.2829, 226.1703, 233.2069, 239.0389, 234.8678, 231.8471, 223.0377, 
    227.7194,
  206.2849, 200.531, 190.801, 182.8051, 188.2599, 195.8225, 202.3677, 
    216.2245, 231.3909, 236.4613, 237.1996, 234.7519, 228.6054, 225.3837, 
    225.0052,
  197.7662, 191.7133, 188.1444, 186.8778, 192.1479, 201.0168, 216.0167, 
    228.4412, 233.9177, 236.7765, 235.2067, 231.354, 227.709, 221.9393, 
    218.3743,
  204.8162, 195.0569, 191.2337, 192.5318, 199.4497, 211.0134, 225.2795, 
    233.4577, 236.1897, 238.9095, 232.4519, 222.0752, 222.3085, 221.4833, 
    220.4265,
  210.6569, 204.6845, 201.0439, 199.9511, 201.645, 214.0589, 226.5197, 
    233.1428, 236.6125, 238.8814, 227.1549, 221.2546, 215.9098, 224.7996, 
    217.9013,
  220.3179, 212.9401, 204.6247, 203.2823, 210.6, 216.9172, 228.2869, 
    240.0453, 240.3805, 236.2143, 221.3556, 220.5387, 220.2273, 225.5343, 
    219.7292,
  181.6585, 198.7924, 216.6106, 222.4678, 218.046, 219.1959, 225.8738, 
    227.6202, 231.5118, 236.4701, 238.6718, 238.3856, 237.4927, 236.6201, 
    237.9839,
  188.2446, 205.4455, 215.3682, 217.9694, 220.1207, 224.435, 227.7275, 
    228.3293, 231.7931, 235.4464, 234.5268, 234.9687, 236.0778, 236.3439, 
    238.7724,
  198.8521, 204.4157, 214.0029, 218.1913, 221.15, 222.9254, 226.7144, 226.93, 
    230.4918, 232.1548, 232.3569, 233.7015, 234.7015, 233.5441, 234.667,
  194.9765, 197.9308, 213.2778, 224.5797, 221.2814, 224.1316, 225.6956, 
    231.7914, 230.6328, 231.42, 233.1374, 233.3122, 233.5928, 227.67, 230.3058,
  189.7827, 199.5837, 215.1391, 228.4765, 224.5775, 216.3709, 220.4955, 
    232.1545, 229.8187, 231.1699, 229.9832, 234.0361, 230.781, 224.8273, 
    223.9925,
  197.5249, 205.7188, 223.0957, 234.3923, 230.7823, 224.9241, 215.018, 
    221.5037, 223.7299, 228.6252, 229.4902, 226.4045, 224.0559, 225.2333, 
    229.668,
  198.5078, 211.0683, 229.3648, 232.2987, 228.1233, 220.9048, 214.1421, 
    219.4823, 223.6599, 226.6963, 231.1955, 224.7373, 225.1243, 222.5994, 
    221.018,
  205.4304, 217.4451, 224.2894, 223.8149, 220.2087, 216.0871, 220.3826, 
    230.738, 236.7273, 235.0435, 226.3578, 222.1478, 225.1112, 224.7474, 
    220.0456,
  203.8147, 215.546, 216.1377, 218.8693, 208.2229, 208.515, 225.8739, 
    236.4676, 237.3652, 227.1704, 219.2214, 216.5932, 216.403, 218.8982, 
    208.6275,
  203.2436, 211.5282, 210.0394, 207.4465, 198.8574, 203.9712, 233.7192, 
    239.9274, 238.7912, 227.2927, 220.9588, 214.678, 214.394, 209.4044, 
    205.0641,
  232.6882, 231.6779, 207.9024, 208.4314, 222.6413, 241.0419, 243.1321, 
    228.8328, 213.2241, 199.4952, 199.3206, 210.6748, 218.8727, 224.8541, 
    235.328,
  216.0068, 223.2119, 213.7029, 217.4036, 232.0557, 244.0977, 244.8031, 
    234.5465, 222.1455, 203.9635, 205.8971, 210.7868, 220.1478, 228.6341, 
    234.7158,
  216.7341, 228.5647, 221.8786, 224.8969, 236.3547, 244.0577, 244.7737, 
    237.0307, 218.8777, 208.3644, 205.8453, 206.9796, 216.4315, 226.7567, 
    231.7699,
  233.8152, 239.5957, 236.6224, 228.976, 239.4872, 243.8667, 239.1826, 
    238.1304, 233.6772, 218.6236, 208.8794, 207.1736, 216.1684, 222.2904, 
    228.3012,
  233.2215, 239.4437, 240.1246, 237.0925, 237.654, 232.756, 230.771, 
    231.3792, 233.6584, 224.7523, 213.2345, 210.6846, 209.9749, 219.2415, 
    215.7571,
  230.1068, 234.294, 237.6518, 237.1971, 236.3952, 230.3783, 222.1225, 
    214.3992, 215.3617, 214.4906, 212.7492, 204.661, 205.1736, 208.5784, 
    215.9089,
  230.1441, 234.8084, 235.6456, 234.4875, 227.4478, 223.257, 220.6962, 
    207.3174, 203.985, 202.3411, 205.1601, 201.5242, 201.8647, 205.9759, 
    215.9808,
  232.3178, 232.5294, 229.4765, 228.4574, 227.7039, 218.1687, 212.1769, 
    210.6068, 211.4833, 215.1991, 212.2529, 210.9911, 220.3148, 226.5552, 
    230.8425,
  234.9531, 231.1423, 228.5243, 223.8066, 225.5167, 224.1611, 232.7816, 
    237.1454, 233.3905, 235.4746, 232.1374, 230.0834, 226.6476, 235.3255, 
    233.7436,
  234.7067, 233.17, 232.0251, 230.8983, 236.3518, 241.7473, 245.9798, 
    245.3116, 237.6274, 225.1715, 222.5594, 220.5778, 229.2917, 232.425, 
    226.1683,
  235.3768, 230.7709, 226.4242, 205.5764, 217.5042, 235.5336, 244.2941, 
    238.4805, 230.3049, 231.4028, 232.5287, 242.6408, 243.1389, 242.303, 
    244.0432,
  230.4418, 216.2142, 199.4302, 193.7354, 205.7857, 233.8514, 239.9915, 
    236.4759, 230.8804, 228.3936, 231.8593, 234.4775, 230.6993, 233.1772, 
    233.9303,
  217.223, 203.5081, 188.1159, 187.9206, 209.1137, 223.5652, 236.6246, 
    228.0824, 221.022, 220.9148, 230.2078, 226.8585, 224.4971, 219.5806, 
    221.6399,
  212.8843, 198.2873, 185.7823, 189.3016, 205.5667, 221.6279, 227.3811, 
    229.6401, 219.3839, 215.5343, 220.1805, 226.2611, 220.312, 216.6954, 
    214.107,
  213.4118, 202.6976, 196.102, 198.1109, 208.107, 225.1616, 232.8544, 
    230.2668, 228.1338, 209.1571, 211.6297, 218.138, 214.6366, 212.708, 
    211.2048,
  231.0715, 231.1264, 223.1455, 218.0734, 222.4079, 231.1216, 238.1221, 
    228.5978, 226.5942, 210.4799, 202.1704, 206.0567, 206.6034, 208.3334, 
    205.6177,
  239.4909, 240.4994, 242.6088, 242.9386, 236.5618, 236.6102, 240.5291, 
    227.38, 225.7691, 215.0191, 203.7264, 198.3769, 200.7869, 197.7175, 
    196.074,
  238.6757, 238.9025, 241.4197, 244.0607, 242.0416, 239.1582, 235.7117, 
    224.8533, 226.0376, 217.9694, 207.2216, 197.4068, 192.9967, 191.8, 
    194.0344,
  226.0499, 226.4744, 225.9908, 226.8324, 228.6597, 230.8997, 228.4283, 
    220.7207, 221.1406, 220.8143, 215.1481, 208.3085, 206.5002, 202.2472, 
    204.6929,
  232.2514, 234.3431, 236.093, 235.898, 234.262, 234.7285, 235.5591, 
    231.4371, 231.0216, 230.5433, 226.02, 220.3843, 219.1606, 215.5879, 
    212.8973,
  221.5739, 223.8502, 223.5961, 224.5466, 216.2454, 216.323, 218.0318, 
    220.0919, 230.8981, 230.5748, 235.7254, 235.2439, 242.2378, 245.1086, 
    248.3774,
  223.0389, 221.011, 217.5643, 220.8911, 222.5843, 230.2139, 225.6295, 
    222.4255, 227.5144, 233.7041, 234.949, 237.8145, 244.5146, 245.8629, 
    248.6919,
  223.9041, 219.8085, 215.0285, 211.8677, 221.0408, 228.2117, 234.5687, 
    223.0089, 227.8452, 235.0489, 235.9532, 239.9815, 245.6449, 246.5942, 
    247.8618,
  228.1338, 221.2574, 206.0034, 209.1508, 208.6004, 230.1185, 230.2399, 
    228.5702, 232.4587, 235.4718, 237.3383, 241.6789, 245.8481, 247.1883, 
    245.8032,
  231.4676, 223.118, 207.0641, 209.6001, 212.9177, 218.7517, 234.0111, 
    230.0776, 233.6869, 240.6306, 238.1806, 244.8391, 246.359, 247.7328, 
    247.8042,
  227.9824, 223.3125, 217.8141, 221.1389, 223.8408, 224.917, 234.5037, 
    238.1592, 237.8811, 237.1283, 240.1087, 244.9962, 247.2524, 247.7467, 
    249.341,
  220.1097, 219.0649, 222.4987, 228.2735, 223.1319, 227.4462, 235.4273, 
    237.3566, 236.4668, 240.371, 243.3092, 245.843, 247.8274, 247.4059, 
    250.6546,
  218.6466, 221.3064, 219.796, 215.99, 220.1438, 222.6598, 236.1132, 
    237.1056, 237.6961, 238.6021, 237.0403, 244.5181, 246.4834, 246.4419, 
    246.4512,
  220.934, 215.3126, 212.957, 213.397, 212.4086, 220.4607, 232.8462, 
    230.1016, 234.3944, 235.5793, 234.7357, 236.3515, 236.6957, 240.5027, 
    239.3039,
  222.404, 218.0735, 215.5591, 212.5752, 216.9552, 221.0264, 226.9513, 
    222.5891, 225.1836, 227.146, 227.0051, 229.8296, 231.6939, 232.8139, 
    229.0707,
  223.2181, 224.2133, 226.9783, 226.7123, 221.8453, 228.3086, 230.5004, 
    225.3742, 227.3695, 224.2677, 226.2319, 222.5804, 212.5746, 216.5136, 
    218.2606,
  225.9468, 229.2014, 228.8574, 228.5586, 225.5347, 224.2658, 224.0867, 
    227.0924, 230.9926, 223.6819, 219.3603, 220.7286, 208.3767, 210.7963, 
    216.4337,
  232.0686, 229.8251, 227.9168, 224.7868, 222.0747, 223.9088, 226.5683, 
    224.6039, 228.3086, 226.5158, 216.5729, 209.1851, 202.9803, 208.3301, 
    215.1453,
  222.7982, 219.4231, 224.6075, 225.8673, 222.646, 224.9226, 223.9399, 
    229.015, 234.6982, 232.8201, 217.5291, 206.6542, 205.7697, 210.319, 
    219.6607,
  215.6062, 220.5843, 225.4134, 223.7922, 224.0085, 219.2366, 221.3192, 
    222.3221, 227.0601, 234.6251, 214.4813, 206.7717, 208.5051, 216.4138, 
    223.8925,
  215.6519, 219.0511, 222.9734, 228.1626, 229.4593, 219.6146, 220.517, 
    222.5368, 235.4279, 231.3696, 211.5207, 211.8406, 217.5041, 223.0186, 
    229.0593,
  215.8557, 217.0025, 215.648, 222.1234, 227.5866, 220.9964, 220.9262, 
    215.5895, 227.9319, 227.3615, 211.9706, 217.301, 223.7324, 227.9672, 
    230.6437,
  216.6077, 209.3486, 207.5897, 227.2168, 224.8757, 217.6021, 219.3861, 
    221.0217, 236.8921, 223.324, 210.5954, 219.2059, 227.3544, 225.7801, 
    229.8036,
  217.0446, 214.73, 205.631, 217.1795, 221.4513, 212.6097, 219.7914, 
    212.8539, 233.4362, 214.4941, 215.5487, 221.7427, 225.6229, 225.277, 
    227.0822,
  216.8705, 214.2807, 208.8815, 209.0054, 211.2098, 213.2782, 212.5953, 
    216.2986, 229.3186, 216.6679, 219.945, 223.2298, 222.3412, 225.5265, 
    229.4496,
  225.1909, 221.3838, 222.9129, 223.0831, 227.1875, 228.0489, 227.2734, 
    226.3473, 229.5252, 231.6224, 233.6955, 232.6559, 233.6245, 238.478, 
    240.302,
  225.0883, 229.3286, 233.5889, 233.5118, 233.5164, 233.9919, 229.3384, 
    228.4121, 232.7984, 229.0032, 227.7078, 235.1154, 234.9569, 236.4529, 
    240.9556,
  236.8054, 237.4704, 232.7117, 229.2994, 228.6291, 225.8955, 228.6353, 
    221.0786, 223.7588, 226.9113, 227.1632, 225.6374, 227.396, 235.8628, 
    238.6774,
  238.4193, 233.4429, 228.1577, 223.1236, 222.4739, 225.8878, 221.7803, 
    225.3293, 224.7804, 224.3093, 225.5303, 222.6926, 230.7321, 234.6483, 
    231.2621,
  229.4424, 221.2874, 213.4487, 214.6297, 216.9206, 217.7792, 222.2825, 
    220.8435, 224.6894, 226.9344, 223.259, 217.8026, 221.6058, 228.951, 
    227.9351,
  215.6023, 209.2676, 208.7603, 209.6087, 210.8537, 216.0055, 220.733, 
    226.219, 227.3817, 230.2271, 223.2472, 216.8539, 221.0178, 228.1045, 
    225.7706,
  209.4623, 208.8334, 203.6755, 203.7921, 209.8112, 222.2481, 222.2976, 
    226.0651, 228.9291, 231.1373, 216.0096, 214.6409, 219.5412, 226.629, 
    227.062,
  206.6279, 206.5443, 212.3997, 211.045, 217.5102, 225.6575, 227.9031, 
    232.598, 231.4825, 219.2182, 210.8541, 212.9316, 222.9839, 230.0175, 
    229.4623,
  205.9138, 210.8678, 213.0966, 214.2885, 222.1289, 221.0086, 229.5746, 
    230.7321, 220.0236, 207.6678, 206.5667, 215.9605, 228.6801, 233.7299, 
    236.2652,
  205.6689, 212.2731, 212.7956, 212.6393, 219.9415, 228.8289, 226.85, 
    221.9415, 206.1372, 203.679, 212.3797, 222.0747, 232.0253, 237.1483, 
    242.9528,
  193.3564, 196.8316, 195.8792, 200.6293, 208.6065, 212.4978, 216.5932, 
    217.701, 221.7605, 224.9422, 242.5103, 240.3171, 238.4062, 239.7228, 
    214.5438,
  189.7324, 194.8593, 204.5413, 206.6967, 216.0488, 220.6978, 224.063, 
    234.4513, 239.0372, 240.1349, 240.5141, 238.7945, 239.0695, 233.9555, 
    205.3163,
  194.8558, 201.3677, 212.8478, 215.4864, 219.7663, 224.127, 228.7536, 
    234.2572, 238.6221, 238.2172, 237.5964, 239.2402, 240.5966, 226.554, 
    194.635,
  210.0652, 215.8045, 222.8542, 230.3336, 229.1755, 234.2607, 233.2152, 
    237.4382, 239.2656, 239.3295, 239.701, 240.0927, 239.2566, 212.8487, 
    189.8219,
  217.5285, 219.9324, 221.4244, 225.4549, 227.0314, 225.5079, 226.9327, 
    226.6002, 234.0328, 235.3242, 235.7077, 237.2438, 232.596, 204.4186, 
    195.0267,
  222.7057, 222.4834, 222.3174, 223.2077, 223.8933, 221.8819, 221.3874, 
    224.4793, 225.4889, 230.9568, 238.7609, 238.6518, 233.8787, 203.149, 
    205.0109,
  230.4989, 226.8032, 227.4189, 226.3541, 221.9274, 216.1709, 214.2803, 
    212.1544, 214.7234, 231.5499, 234.9977, 235.8978, 229.1782, 203.3726, 
    208.2927,
  224.4973, 223.4862, 225.0271, 219.2815, 212.7663, 209.3705, 209.4845, 
    212.7907, 222.6502, 233.857, 234.1572, 235.2937, 227.2332, 206.3295, 
    222.4584,
  224.9667, 222.2244, 217.2674, 214.0194, 209.6598, 205.4804, 207.5286, 
    211.2193, 220.6198, 231.718, 233.9541, 234.3656, 226.3956, 217.7827, 
    229.5496,
  227.8926, 221.1884, 212.1341, 212.2734, 215.6869, 215.159, 214.3885, 
    217.226, 226.3337, 233.0889, 235.3635, 232.6285, 223.4861, 229.3408, 
    230.0187,
  233.8932, 233.5543, 212.5764, 196.9617, 194.0328, 203.2165, 190.5847, 
    189.3407, 183.1716, 199.7603, 209.0072, 227.7322, 242.101, 243.9348, 
    238.3363,
  210.8469, 232.035, 218.9996, 202.1289, 194.4668, 195.1902, 189.7603, 
    190.1082, 192.6819, 205.5416, 215.781, 229.3499, 241.6837, 239.8033, 
    239.4375,
  197.7114, 216.5677, 215.8087, 202.026, 193.6364, 193.8997, 190.0691, 
    187.0832, 198.9636, 205.8053, 217.6404, 235.5489, 240.4572, 240.2, 
    241.9553,
  193.4859, 195.799, 199.4008, 198.7806, 200.122, 198.773, 194.7867, 195.836, 
    199.0319, 210.1746, 221.4202, 236.807, 240.8923, 238.5478, 240.1793,
  191.3618, 186.7668, 188.3304, 192.6219, 198.1673, 193.9007, 204.3202, 
    208.4523, 209.1641, 211.7021, 225.9111, 240.7391, 238.6359, 232.6477, 
    233.809,
  198.1893, 182.8519, 190.7107, 194.0692, 203.8918, 200.378, 200.0233, 
    203.6486, 211.6266, 223.3981, 235.6851, 238.3597, 235.4066, 227.378, 
    224.4807,
  223.4992, 190.825, 190.4183, 199.8686, 203.1287, 205.7682, 210.8393, 
    210.1149, 219.8129, 233.2719, 238.4247, 236.2508, 229.5435, 219.6691, 
    220.1576,
  240.366, 206.6431, 197.3357, 201.8294, 211.9553, 212.6469, 220.4941, 
    234.1641, 238.1142, 237.6395, 236.3813, 234.3936, 225.4068, 211.9786, 
    213.6153,
  233.1075, 227.6909, 206.8587, 204.2009, 211.2674, 216.5997, 223.7946, 
    235.1184, 237.0517, 235.6847, 235.4966, 230.2488, 212.1358, 204.8037, 
    216.4476,
  235.1809, 235.0178, 221.9885, 214.8771, 214.0978, 216.8968, 222.0681, 
    229.7017, 233.6784, 234.4278, 231.6351, 225.3495, 199.6632, 205.8323, 
    225.9479,
  232.9039, 228.8556, 217.0599, 225.2899, 245.4102, 247.7832, 236.7652, 
    212.1138, 197.6374, 197.6371, 192.6161, 190.8188, 194.8118, 200.5932, 
    210.9334,
  223.149, 227.2727, 216.3191, 220.1467, 234.4907, 230.1478, 207.3616, 
    200.0831, 194.2999, 184.8822, 188.4537, 191.5076, 194.8569, 208.6119, 
    230.6464,
  223.0424, 223.1498, 218.3394, 212.3233, 221.8886, 211.9737, 199.9219, 
    192.9056, 194.2996, 186.6134, 185.5662, 191.4894, 205.3145, 226.3326, 
    238.3873,
  220.0286, 222.7027, 224.96, 211.8488, 206.6029, 208.3571, 195.7967, 
    202.0191, 200.598, 194.9612, 189.3714, 197.2842, 223.102, 237.3159, 
    239.3859,
  219.3465, 220.0656, 222.9111, 225.2313, 215.2902, 204.1475, 213.9293, 
    224.812, 206.7223, 191.4599, 195.1757, 212.4457, 234.4577, 236.4772, 
    236.4666,
  223.282, 223.4724, 223.1059, 232.0927, 225.9159, 224.8214, 218.1661, 
    201.7288, 195.9034, 196.6427, 205.0454, 232.6213, 234.5188, 234.0659, 
    234.5161,
  232.0304, 235.6432, 221.3838, 230.8432, 222.7591, 218.3004, 218.7741, 
    203.1881, 199.1821, 210.3647, 233.0433, 234.3983, 233.2983, 233.9695, 
    230.3272,
  229.3644, 231.4822, 216.643, 220.4748, 220.5832, 210.2544, 205.7312, 
    198.8206, 208.3987, 226.6499, 234.3235, 231.9195, 230.3727, 226.7814, 
    226.1358,
  235.267, 236.0991, 214.3447, 210.8741, 207.7775, 200.2338, 197.6147, 
    197.1145, 211.5181, 231.0116, 231.594, 230.5963, 228.2086, 224.3212, 
    228.6074,
  233.6772, 232.319, 212.0986, 200.9548, 199.7484, 197.8598, 190.7153, 
    200.612, 224.5048, 231.2141, 231.2008, 229.2861, 222.7788, 228.445, 
    228.8339,
  227.4355, 211.1537, 204.0038, 214.2346, 225.917, 226.3843, 231.8068, 
    243.3823, 240.6288, 233.0563, 221.1526, 203.2467, 193.7964, 193.4632, 
    204.0321,
  225.5057, 210.7784, 203.8175, 209.8734, 223.4875, 224.5155, 229.1316, 
    238.8689, 240.6045, 239.32, 232.4732, 224.7131, 222.2451, 214.7966, 
    220.8366,
  218.9558, 203.0539, 201.017, 203.5303, 217.5161, 225.0908, 228.6156, 
    227.8936, 238.0003, 237.3331, 224.7188, 218.4689, 215.1792, 224.7515, 
    239.5529,
  227.7529, 218.5411, 207.4715, 207.3308, 209.1351, 216.7082, 225.2754, 
    228.7339, 227.8477, 223.04, 212.5369, 210.2301, 218.6508, 235.3069, 
    239.8385,
  233.8766, 224.6097, 217.5175, 211.513, 214.6207, 213.887, 222.606, 231.147, 
    218.6843, 208.2868, 205.5371, 205.8881, 223.031, 234.584, 237.6301,
  230.1591, 220.5527, 215.9938, 215.6423, 218.6672, 216.5128, 220.8888, 
    215.1958, 213.6073, 214.6389, 210.567, 222.0966, 227.2177, 233.5182, 
    233.1284,
  231.1844, 224.9036, 220.5518, 217.2502, 213.7192, 215.6339, 213.6213, 
    208.732, 209.1436, 209.9981, 215.7522, 221.5368, 232.4788, 233.7131, 
    229.7643,
  220.9905, 214.6154, 212.0433, 214.3004, 208.303, 205.4033, 206.282, 
    204.2368, 207.8163, 208.1599, 219.5637, 230.2452, 230.4217, 229.0341, 
    226.0291,
  205.9721, 197.4445, 198.267, 200.856, 201.9835, 200.6082, 203.2457, 
    204.9884, 206.4667, 212.4509, 226.9346, 230.9226, 229.3438, 222.868, 
    219.3669,
  201.8398, 195.5645, 191.9274, 195.291, 197.5567, 197.7311, 206.5251, 
    210.5964, 210.7793, 225.2542, 230.6246, 230.2162, 226.4344, 218.9104, 
    215.5273,
  212.1373, 211.4645, 209.3459, 214.7063, 217.4784, 216.5102, 216.9803, 
    221.489, 220.2251, 225.4379, 225.2335, 227.3814, 226.0611, 225.0934, 
    224.6414,
  201.6047, 203.7884, 204.1212, 209.1316, 215.6748, 217.6799, 212.4996, 
    219.509, 220.4533, 221.6731, 217.828, 219.6246, 219.8911, 217.3004, 
    218.4618,
  205.1149, 210.1594, 211.3011, 212.7013, 213.9224, 217.6292, 216.8686, 
    216.1225, 215.263, 218.9864, 217.4727, 213.2886, 214.0169, 212.2008, 
    218.0916,
  214.2582, 221.095, 223.552, 229.944, 233.8579, 236.381, 231.1816, 227.1534, 
    219.1246, 208.5629, 210.7301, 207.9856, 210.051, 200.9675, 208.3322,
  228.2875, 231.5012, 236.0602, 239.1767, 240.9201, 240.86, 238.4907, 
    231.2074, 223.8734, 217.7775, 209.8907, 209.8148, 203.0442, 203.7946, 
    208.0577,
  235.7225, 239.1222, 243.4181, 243.437, 245.1461, 246.1259, 241.2783, 
    234.7967, 225.6002, 219.3944, 212.2898, 208.332, 206.5272, 208.9653, 
    216.1288,
  246.4062, 246.4787, 245.0202, 245.3422, 246.1201, 246.0664, 242.6093, 
    234.9075, 222.7189, 219.5014, 217.2791, 211.7906, 208.2614, 212.7231, 
    221.8955,
  249.377, 247.1793, 244.0599, 243.6416, 242.7796, 240.6259, 237.6258, 
    228.871, 226.5476, 221.0791, 212.6879, 215.2787, 214.1404, 217.5267, 
    224.0862,
  245.3155, 242.8262, 236.5745, 232.3473, 232.843, 233.3112, 230.7989, 
    225.3329, 220.7073, 215.342, 215.0272, 216.5005, 215.8082, 222.028, 
    230.0125,
  242.9129, 237.8369, 207.6736, 207.3154, 222.7248, 227.814, 226.2933, 
    219.8578, 217.0526, 213.825, 213.3226, 216.2479, 224.2063, 230.8844, 
    229.5596,
  233.0447, 231.1306, 226.4648, 214.2286, 203.9998, 197.0162, 189.933, 
    184.6035, 191.8851, 196.6282, 198.8411, 198.1552, 201.2751, 202.6329, 
    202.7668,
  213.8008, 212.5733, 207.2597, 201.6803, 201.6925, 194.5819, 192.6786, 
    194.4365, 199.134, 201.5652, 204.327, 203.3835, 206.5298, 209.0508, 
    208.6186,
  203.3674, 198.8929, 198.8288, 197.8212, 204.3573, 197.8343, 196.6916, 
    194.6496, 202.3402, 208.2335, 207.3523, 208.7152, 211.3526, 210.0558, 
    211.0121,
  196.3768, 190.4572, 192.1681, 197.8602, 200.4344, 206.7331, 210.4715, 
    211.8435, 212.7457, 211.1578, 216.3104, 218.5476, 215.6786, 214.3209, 
    215.177,
  199.2659, 199.1958, 200.4466, 212.4091, 214.4592, 220.9709, 225.5859, 
    231.8728, 232.9188, 236.1295, 234.6285, 237.6068, 235.2934, 228.8314, 
    227.9191,
  210.5469, 216.3977, 220.9871, 226.9428, 230.7907, 235.3595, 235.7024, 
    236.8624, 236.1792, 236.087, 236.8812, 238.2792, 236.8324, 232.109, 
    225.3367,
  226.6348, 228.1179, 230.5205, 234.3251, 237.1691, 236.9095, 234.882, 
    233.8998, 234.4252, 232.342, 232.7245, 235.7742, 235.2339, 230.131, 
    222.6708,
  229.9903, 233.9103, 235.5396, 236.4801, 235.6122, 230.4663, 226.0536, 
    221.398, 215.7087, 215.7013, 214.3844, 219.6937, 225.0996, 217.2457, 
    216.9047,
  233.445, 235.6252, 236.3595, 233.6953, 232.3244, 227.8374, 225.0693, 
    220.0182, 216.3441, 213.4326, 215.9727, 221.6668, 220.2735, 214.9733, 
    211.2678,
  239.2115, 237.9176, 230.9167, 235.0964, 237.2668, 233.5022, 235.0778, 
    225.7983, 217.5711, 218.8798, 220.2471, 217.627, 216.0914, 209.4648, 
    207.5628,
  249.9071, 248.5664, 251.6884, 252.6509, 252.7127, 247.6509, 247.998, 
    246.2189, 239.4387, 237.144, 229.4282, 227.8615, 222.9231, 216.3741, 
    206.7218,
  246.9531, 251.9555, 255.6944, 255.9936, 251.4956, 250.9415, 247.0278, 
    240.6621, 232.2897, 225.9182, 219.6294, 218.4546, 215.2915, 214.3331, 
    209.1046,
  239.3121, 247.367, 250.9401, 248.5905, 247.6339, 241.0838, 236.7479, 
    228.838, 226.9431, 218.3115, 219.224, 215.4239, 212.4803, 210.7891, 
    207.5015,
  216.6924, 221.3248, 225.0834, 232.3468, 230.9314, 232.0199, 224.8499, 
    223.1994, 222.3846, 220.06, 216.5169, 213.924, 213.8326, 213.5739, 
    214.2624,
  212.0005, 208.3409, 206.4538, 202.5038, 210.1599, 215.3987, 217.9498, 
    219.7, 220.5663, 220.4049, 217.204, 220.3161, 219.8436, 219.3761, 214.8541,
  211.2268, 199.5826, 192.3951, 192.7706, 191.2525, 194.2412, 200.6974, 
    213.9684, 221.1691, 226.3429, 224.4585, 224.8073, 225.0465, 224.5197, 
    224.7996,
  217.1706, 208.2424, 199.9779, 195.7665, 203.817, 204.2147, 211.3773, 
    212.2904, 216.0026, 215.9601, 220.2485, 224.0361, 225.2097, 232.5794, 
    233.9255,
  220.4095, 222.3795, 224.4276, 221.7343, 228.4421, 231.2455, 233.5798, 
    235.5984, 234.4582, 231.22, 228.4677, 226.853, 228.9155, 234.9863, 
    228.3379,
  225.4346, 228.5003, 230.6781, 229.4978, 232.3746, 234.8038, 235.5926, 
    235.5114, 235.2802, 232.0349, 224.0921, 223.8697, 223.3235, 232.489, 
    224.4708,
  232.1382, 228.3563, 229.984, 230.4785, 231.0706, 234.5507, 237.3251, 
    237.8217, 235.0884, 227.6994, 219.8825, 214.29, 221.0827, 219.9729, 
    221.9068,
  191.5568, 198.1664, 208.1706, 220.466, 229.3293, 235.6639, 240.4408, 
    244.0519, 245.968, 248.9027, 250.7735, 250.9243, 252.3778, 254.0195, 
    254.7836,
  190.2015, 197.9411, 205.0031, 212.7832, 222.1759, 234.9513, 243.0036, 
    244.5457, 246.2313, 248.2635, 251.3577, 250.0071, 250.5658, 249.7991, 
    251.2179,
  198.703, 204.5285, 210.721, 213.9781, 223.0762, 231.6847, 239.7445, 
    242.2293, 244.5381, 245.8599, 248.166, 248.8096, 250.1616, 248.972, 
    247.1322,
  213.9625, 215.4253, 218.5232, 220.869, 224.877, 228.1958, 231.3519, 
    239.991, 241.8349, 244.9668, 246.7101, 248.4741, 249.6021, 248.2326, 
    246.4597,
  226.2503, 226.0314, 226.0698, 226.4966, 227.268, 225.083, 230.0127, 
    233.0823, 232.1731, 239.3133, 241.7297, 245.1665, 247.591, 246.785, 
    242.712,
  233.733, 230.2814, 231.1816, 230.5959, 228.7379, 224.632, 220.6618, 
    226.9778, 224.7347, 229.248, 229.8925, 229.1026, 234.8927, 235.1512, 
    230.4906,
  228.481, 229.3543, 227.4965, 225.3319, 222.9301, 219.5928, 221.0327, 
    223.1704, 225.6817, 223.9911, 218.1671, 213.107, 217.2886, 217.192, 
    209.6563,
  223.8699, 223.6278, 219.8349, 218.908, 219.1218, 220.57, 222.6755, 
    228.6416, 228.5079, 230.0027, 227.4343, 216.287, 209.7374, 206.3083, 
    196.384,
  223.6017, 216.5697, 217.7259, 220.2826, 222.2631, 224.8403, 226.2442, 
    229.4518, 231.7917, 232.5396, 228.1682, 226.3103, 221.8369, 207.5623, 
    196.7935,
  221.1726, 219.7241, 222.3589, 223.7826, 227.2769, 225.9272, 225.7003, 
    224.5132, 230.5492, 221.6938, 228.0397, 229.8901, 226.5563, 218.9919, 
    211.1911,
  236.111, 221.4462, 218.3574, 218.6555, 220.3793, 232.7458, 237.0042, 
    231.4822, 231.4081, 235.8167, 236.1674, 230.2048, 233.3646, 238.6544, 
    242.2753,
  235.6611, 234.8472, 223.4671, 212.4765, 224.0438, 222.1543, 233.8484, 
    231.9486, 236.1199, 232.654, 234.021, 231.1452, 236.5265, 240.2395, 
    241.6925,
  230.4277, 228.9053, 221.8634, 215.9494, 213.6113, 210.8388, 220.6318, 
    221.2444, 225.8657, 229.6191, 230.486, 228.9338, 234.5698, 240.4058, 
    237.404,
  217.855, 217.9902, 213.6703, 210.9823, 207.3353, 204.3744, 204.5234, 
    208.1198, 214.0022, 215.7372, 219.0817, 224.8902, 229.9007, 233.8059, 
    232.4263,
  208.7146, 208.1461, 209.7354, 206.6202, 204.3766, 195.6787, 199.9402, 
    205.8268, 213.1966, 207.6865, 213.6049, 223.0483, 226.4054, 229.1562, 
    228.0958,
  217.3688, 208.5357, 208.8861, 206.4097, 205.7955, 204.1987, 204.8147, 
    204.9479, 211.204, 213.1217, 223.8112, 225.7636, 230.0257, 223.78, 
    224.5456,
  229.901, 222.6174, 215.5976, 212.7705, 212.1714, 213.3423, 213.4075, 
    211.0054, 210.7116, 217.34, 225.3033, 231.8219, 229.6997, 221.6116, 
    211.7631,
  234.629, 232.1327, 222.3859, 220.167, 217.5545, 218.0997, 221.3236, 
    222.6927, 220.2399, 224.8599, 227.7986, 230.9718, 224.098, 213.9267, 
    203.6355,
  229.9635, 226.3661, 225.3363, 224.6664, 222.7647, 224.3887, 228.1673, 
    227.6064, 226.2289, 230.2105, 231.2535, 227.2929, 221.9945, 209.4379, 
    195.3387,
  223.2346, 220.3094, 219.9553, 223.4225, 225.9072, 223.1489, 231.4004, 
    229.3681, 230.0403, 235.416, 234.4647, 223.8793, 215.3262, 199.0314, 
    194.2726,
  234.5627, 233.784, 220.1011, 226.3414, 235.238, 250.7794, 256.2926, 
    259.5032, 261.3705, 267.117, 260.7005, 252.8294, 247.7337, 239.1315, 
    234.6898,
  238.9826, 240.9124, 231.0428, 227.2079, 234.9389, 251.1798, 255.4991, 
    256.2188, 257.7749, 261.2321, 261.7845, 254.1542, 246.3024, 237.5173, 
    233.2184,
  239.3361, 244.0801, 242.8588, 236.8583, 234.0979, 238.8165, 251.7926, 
    251.9655, 256.0924, 256.6736, 256.7635, 250.2411, 241.3942, 232.2763, 
    227.5277,
  236.2406, 243.0542, 247.8731, 242.3559, 240.2651, 236.0866, 233.8911, 
    247.6239, 250.9033, 252.2001, 248.4915, 240.0048, 233.5392, 229.4776, 
    220.2931,
  232.3475, 238.8062, 244.7953, 245.5055, 244.9845, 236.3391, 233.8716, 
    239.4512, 239.0827, 241.1247, 236.1748, 233.8404, 231.6753, 219.5702, 
    206.0323,
  230.8199, 233.2981, 239.7125, 243.5641, 246.5573, 240.6917, 226.6324, 
    227.4739, 226.3906, 221.5511, 222.1232, 217.8808, 208.3131, 200.6836, 
    197.6695,
  231.054, 232.0509, 232.4479, 237.0314, 242.8802, 236.1645, 231.0806, 
    215.1233, 210.0235, 210.5607, 216.6667, 203.6598, 204.6252, 193.285, 
    197.6263,
  234.3469, 232.1318, 231.9555, 228.8881, 234.8873, 240.119, 231.0613, 
    224.5971, 215.6579, 208.6192, 204.4021, 201.7581, 198.7572, 199.2143, 
    205.2776,
  228.0531, 234.0722, 229.9683, 227.7948, 226.0086, 230.1396, 228.8205, 
    220.0034, 218.578, 206.0552, 202.7228, 201.9255, 198.572, 206.432, 
    214.3148,
  218.6391, 222.033, 229.6054, 228.4372, 223.6263, 222.3635, 220.2063, 
    219.9726, 214.424, 206.3552, 203.0524, 200.1641, 208.5983, 215.2362, 
    218.3646,
  199.4574, 196.2631, 205.8965, 224.5815, 231.6651, 237.8209, 241.0139, 
    249.6678, 258.5923, 267.5862, 260.2731, 258.7933, 258.4945, 250.506, 
    242.7901,
  206.2025, 196.2026, 202.1923, 211.999, 227.7428, 233.7495, 236.4157, 
    246.5838, 255.9561, 258.7852, 261.5283, 249.5561, 251.4442, 253.4894, 
    244.0687,
  215.5177, 204.4455, 202.6072, 203.1171, 214.1984, 230.2126, 231.9119, 
    238.8033, 251.7061, 256.9734, 260.0964, 251.3588, 252.7532, 247.7598, 
    245.8393,
  230.4947, 221.1936, 208.4865, 206.698, 206.695, 220.9369, 229.4225, 
    233.3229, 240.7299, 250.9642, 256.3381, 258.2939, 255.2235, 249.6363, 
    245.5338,
  233.5878, 232.5072, 225.9369, 218.762, 208.4444, 214.3677, 228.6588, 
    239.3191, 240.7887, 238.8799, 244.7499, 255.0328, 256.5784, 247.378, 
    234.9985,
  235.191, 235.2614, 233.9913, 233.7472, 226.7883, 218.6109, 224.0387, 
    232.1074, 232.4911, 232.3521, 235.0929, 244.7783, 245.0095, 241.3215, 
    232.5254,
  237.2952, 235.9469, 235.4522, 234.0896, 238.4949, 231.3897, 232.2364, 
    228.1475, 229.4622, 233.5252, 230.7104, 231.5676, 233.2157, 228.211, 
    219.4315,
  236.3364, 238.4751, 236.0143, 236.4175, 240.037, 241.9161, 241.7447, 
    238.6165, 235.192, 233.5356, 226.6246, 229.0442, 227.0808, 217.2172, 
    206.5611,
  218.689, 236.3264, 235.59, 235.2948, 239.971, 241.1875, 245.9939, 245.8584, 
    241.0977, 236.0215, 229.6567, 223.81, 216.1125, 210.8925, 200.01,
  214.5515, 224.4139, 229.4468, 235.4197, 238.2397, 239.723, 243.6559, 
    246.079, 245.4543, 238.2042, 230.0175, 220.2011, 208.1238, 203.2844, 
    195.227,
  180.5534, 206.145, 217.0072, 236.3246, 240.2831, 241.8218, 239.9564, 
    240.456, 248.3438, 264.117, 271.6079, 268.5232, 264.1258, 266.8839, 
    263.7141,
  176.4645, 191.6134, 209.7929, 230.2965, 231.1637, 235.812, 236.4314, 
    239.9538, 250.5803, 264.1349, 269.5805, 267.4523, 267.0102, 266.2644, 
    264.7225,
  177.8796, 180.3837, 200.2013, 217.6124, 231.7065, 232.2059, 231.7889, 
    232.875, 242.0522, 257.3746, 259.4128, 264.0154, 266.0686, 264.2179, 
    260.7179,
  184.5273, 179.2676, 189.5608, 208.3917, 222.5415, 229.6392, 228.1015, 
    230.1653, 233.1365, 249.3527, 247.1602, 257.3311, 262.7585, 265.7847, 
    264.9785,
  198.9484, 186.8194, 184.3707, 194.4436, 212.0589, 222.4718, 227.1492, 
    235.8223, 239.4034, 240.842, 240.189, 248.1551, 254.6402, 259.6753, 
    259.3092,
  213.0233, 200.2903, 193.5917, 194.5337, 198.1615, 210.9357, 220.2358, 
    225.3418, 221.5576, 229.5344, 238.7223, 238.9492, 245.6209, 246.1876, 
    248.195,
  226.2997, 216.5899, 207.0754, 198.6653, 200.4409, 205.248, 212.2786, 
    216.8391, 220.3189, 232.2978, 235.0058, 237.7464, 239.1866, 237.1599, 
    238.9479,
  242.8565, 226.9958, 223.2535, 212.2184, 209.418, 207.8299, 211.9664, 
    216.9185, 222.3967, 230.5937, 229.4084, 233.5357, 233.2316, 234.0868, 
    225.9381,
  247.1685, 237.6983, 233.5363, 225.0871, 218.6576, 213.1272, 215.954, 
    220.2624, 221.093, 223.232, 225.6859, 229.8079, 228.3624, 225.0717, 
    220.0718,
  235.0833, 231.0002, 230.5333, 234.0062, 228.4597, 223.2594, 222.0407, 
    224.703, 226.5773, 228.2859, 231.3071, 232.7978, 226.1349, 221.107, 
    215.2145,
  236.6359, 248.2789, 250.5479, 242.136, 249.3474, 247.4157, 229.5436, 
    222.0291, 238.5788, 270.042, 274.7439, 271.9362, 273.7631, 273.1014, 
    275.0076,
  225.7246, 242.9617, 249.8186, 248.0169, 253.5615, 249.5029, 230.4604, 
    218.1282, 229.1107, 261.9495, 274.9818, 272.3704, 264.2052, 272.052, 
    273.7268,
  218.2738, 231.9518, 246.3734, 246.4992, 252.0228, 244.1496, 229.0929, 
    215.3479, 216.1566, 245.6367, 269.1483, 263.6473, 257.9081, 262.4837, 
    264.7911,
  208.7031, 222.7514, 234.868, 240.2073, 244.6761, 241.9828, 223.3072, 
    217.3318, 215.6174, 235.9465, 252.4947, 262.6743, 262.5494, 261.6198, 
    268.0125,
  196.1335, 206.2195, 223.8137, 233.8872, 237.706, 231.2299, 228.0385, 
    219.2542, 223.8217, 228.8947, 246.8255, 254.7131, 260.5304, 263.2678, 
    262.601,
  190.92, 199.058, 212.7715, 226.1349, 229.9642, 228.1145, 218.9417, 
    213.4656, 214.7299, 225.6483, 237.5632, 239.7039, 246.0636, 254.9085, 
    259.9293,
  201.8233, 196.5874, 205.2793, 218.4914, 222.309, 221.7664, 221.439, 
    213.8795, 213.0959, 220.0217, 226.3548, 228.8249, 232.69, 242.2185, 
    244.6257,
  207.87, 199.3625, 202.9152, 211.03, 218.3318, 216.6996, 223.1269, 216.4991, 
    216.0521, 218.9584, 217.6285, 222.9943, 223.1917, 226.0767, 231.6519,
  228.1712, 212.9107, 204.2232, 206.5377, 212.6403, 216.1958, 216.9594, 
    214.8454, 214.985, 216.1362, 216.9462, 222.6511, 222.3151, 221.1282, 
    228.2869,
  244.8583, 234.3861, 216.1891, 211.1723, 213.8547, 212.0585, 209.6662, 
    210.8457, 212.0568, 212.0336, 220.498, 216.7249, 224.8115, 218.9094, 
    224.8608,
  220.5218, 234.2147, 238.0629, 240.9611, 249.3366, 229.2299, 209.1154, 
    202.0933, 226.3521, 264.2501, 278.97, 274.9008, 276.8175, 275.1948, 
    275.2541,
  213.9538, 237.5028, 242.0008, 235.5128, 249.105, 230.1906, 213.1585, 
    202.7149, 226.6689, 263.1315, 277.7831, 270.7949, 268.3537, 275.0404, 
    275.4844,
  209.0927, 239.1858, 236.7117, 236.0597, 248.0198, 224.0719, 218.3327, 
    202.8442, 229.896, 257.9935, 266.0493, 267.5958, 261.3578, 267.0197, 
    266.7899,
  207.3985, 236.1906, 234.4105, 236.4064, 242.3868, 226.8712, 223.0081, 
    212.7579, 232.9366, 250.4554, 260.1165, 261.3156, 261.8705, 263.3888, 
    264.009,
  205.1525, 231.6814, 233.6273, 235.5393, 242.1454, 221.8463, 226.8334, 
    221.7347, 235.961, 248.2565, 260.9196, 261.5734, 261.2706, 264.0983, 
    264.6234,
  207.6431, 217.5871, 234.5968, 235.1007, 240.499, 225.0429, 223.1901, 
    219.075, 228.7648, 239.8624, 261.5081, 261.2874, 263.2581, 259.1862, 
    259.3053,
  215.031, 209.7635, 228.2228, 236.9808, 234.588, 228.5337, 230.1569, 
    217.3597, 221.6606, 236.4857, 253.7704, 259.5526, 261.2688, 259.3016, 
    253.7011,
  208.1229, 203.419, 216.7387, 224.725, 227.5204, 231.6075, 232.8396, 
    228.3263, 232.2803, 234.4052, 243.0382, 254.4297, 260.6484, 261.1338, 
    253.4228,
  217.596, 222.3463, 212.1731, 221.7749, 225.049, 227.9713, 234.1797, 
    232.3124, 229.856, 233.4745, 237.459, 249.9227, 258.759, 257.1741, 
    250.3958,
  234.5631, 222.1236, 222.445, 223.3408, 221.6558, 223.957, 238.2709, 
    241.2001, 239.476, 231.3938, 236.3692, 236.8792, 243.6516, 246.1664, 
    247.5103,
  231.8349, 234.5791, 237.318, 239.4944, 241.7964, 246.7532, 242.7123, 
    226.749, 222.9822, 250.8469, 272.0692, 273.4205, 268.3123, 246.4048, 
    220.1726,
  228.7959, 233.6604, 237.0271, 238.2746, 242.7077, 246.11, 243.7751, 
    227.7037, 229.7536, 249.9338, 271.118, 268.5411, 259.8788, 227.378, 
    227.593,
  229.7797, 233.5297, 235.6644, 236.9028, 239.8439, 238.8383, 242.6461, 
    226.6886, 228.3225, 249.6333, 261.951, 262.8384, 247.5019, 226.7992, 
    245.1722,
  225.0059, 233.2863, 234.4145, 236.1016, 235.7523, 240.9745, 231.8621, 
    229.8366, 236.3062, 251.9511, 258.4194, 252.214, 238.944, 231.6497, 
    258.1149,
  224.2922, 230.9673, 233.4681, 233.5255, 234.2545, 230.6581, 230.3495, 
    227.8952, 236.8182, 252.2173, 259.8015, 250.4752, 238.1498, 250.778, 
    260.472,
  221.5782, 229.5214, 232.8731, 232.5379, 233.0382, 228.0345, 219.965, 
    222.495, 239.4569, 256.165, 260.3333, 248.584, 242.8983, 255.8011, 255.423,
  221.7128, 225.5606, 231.6822, 234.6011, 232.093, 226.1994, 215.505, 
    215.5064, 238.8571, 260.5901, 257.4875, 250.1138, 249.4276, 251.376, 
    251.1192,
  216.9063, 221.5029, 225.6393, 234.1361, 232.362, 220.0513, 214.1118, 
    220.7338, 242.8821, 260.5422, 256.7117, 249.489, 253.1091, 246.7889, 
    246.824,
  218.0034, 216.1636, 223.9857, 229.7669, 228.6614, 218.6678, 212.7885, 
    217.6864, 242.2143, 260.0143, 259.1034, 254.8306, 251.7899, 251.8527, 
    242.3656,
  224.3624, 220.6311, 217.7755, 224.4346, 223.5302, 213.9463, 214.185, 
    219.0167, 239.4806, 258.6704, 256.6684, 255.0825, 251.3847, 245.5486, 
    246.7536,
  252.9655, 245.5742, 240.2141, 239.973, 239.041, 239.1818, 238.8331, 
    237.2494, 239.8116, 246.0832, 251.8342, 256.5992, 253.1906, 251.9265, 
    267.1861,
  240.86, 241.6926, 239.7943, 241.6694, 240.4916, 240.4405, 239.9438, 
    240.7859, 239.3145, 243.8773, 249.942, 255.1837, 253.7054, 254.2996, 
    264.7396,
  236.008, 235.1404, 237.6151, 240.0407, 242.3601, 239.7492, 242.1114, 
    242.2669, 240.9411, 242.2352, 248.5983, 254.797, 252.4426, 251.0022, 
    260.546,
  233.4656, 231.4221, 236.4257, 237.3183, 239.6095, 242.8121, 239.7907, 
    247.706, 245.7859, 241.9763, 249.0771, 252.8597, 250.6115, 252.0663, 
    257.4886,
  234.4327, 231.6933, 234.1728, 235.553, 237.0779, 240.6003, 243.5789, 
    240.7199, 244.1689, 239.2489, 243.8742, 249.3222, 249.7109, 253.69, 
    254.5539,
  228.241, 230.3715, 231.7026, 232.9852, 236.389, 238.1664, 241.7514, 
    245.3586, 246.1267, 236.246, 238.4616, 242.7088, 251.9364, 254.0342, 
    254.0432,
  223.9172, 224.5577, 223.7686, 226.2202, 231.0787, 236.5314, 241.0754, 
    244.8923, 246.0559, 241.7884, 229.6226, 234.3433, 250.956, 256.4683, 
    253.9469,
  223.8476, 216.9578, 219.9807, 226.7954, 230.8822, 235.9021, 238.6861, 
    246.2643, 248.0165, 242.9058, 227.0118, 236.7857, 254.2268, 257.4297, 
    253.6717,
  217.7197, 215.5569, 217.3441, 217.8736, 225.2115, 234.9481, 239.7014, 
    244.3854, 249.6075, 244.9194, 229.1452, 234.5172, 253.8214, 258.1422, 
    253.8985,
  218.8631, 216.9656, 216.6229, 216.5639, 229.1513, 236.6265, 241.7434, 
    247.6663, 250.7118, 244.0954, 225.8888, 228.758, 252.5748, 254.8409, 
    251.7384,
  234.205, 232.8179, 240.9131, 239.9978, 240.1906, 239.6878, 237.7355, 
    236.4928, 239.2634, 242.7151, 241.9993, 245.3641, 238.2394, 230.4248, 
    238.2418,
  238.8893, 238.8347, 239.4315, 238.2801, 240.3382, 241.5369, 241.0527, 
    238.6052, 239.7303, 238.9651, 245.6306, 243.4711, 234.9494, 231.5994, 
    240.4377,
  233.4594, 240.0672, 241.8719, 238.738, 239.1457, 238.597, 244.5452, 
    239.1143, 241.7387, 240.8024, 245.1597, 245.9566, 231.5506, 225.7306, 
    231.7396,
  228.3762, 229.2777, 238.2759, 241.572, 238.5106, 238.9854, 238.0906, 
    244.2261, 246.6004, 241.0512, 241.3476, 242.1944, 229.9107, 226.8819, 
    234.3665,
  244.1967, 243.028, 237.0155, 238.8395, 238.6758, 237.3685, 238.4566, 
    239.3843, 238.8495, 239.5332, 239.6086, 245.3059, 237.7821, 227.5367, 
    229.9864,
  239.2871, 235.579, 231.3354, 230.2606, 234.6837, 239.8602, 240.842, 
    239.9614, 239.8961, 240.1958, 235.1825, 243.7505, 240.6444, 228.5412, 
    221.5841,
  227.8252, 228.5731, 228.2935, 230.5475, 229.2736, 230.1884, 234.2422, 
    238.0889, 241.9276, 240.8187, 238.543, 240.1321, 248.8992, 236.0924, 
    219.6272,
  229.0299, 229.8016, 229.0027, 230.1527, 229.742, 230.0505, 232.9888, 
    240.861, 241.4668, 241.3854, 239.6404, 238.6757, 247.742, 245.184, 227.952,
  233.36, 231.7883, 230.3364, 229.8862, 226.8472, 225.2549, 230.4318, 
    236.3889, 241.3778, 243.5217, 241.1802, 237.9205, 243.5052, 250.3836, 
    238.6144,
  235.6463, 228.9053, 228.3373, 229.5976, 226.6281, 227.1329, 229.5943, 
    235.0193, 238.9756, 242.1906, 242.0661, 236.5254, 242.9973, 250.2889, 
    244.1418 ;

 scalar_axis = 0 ;

 sfcWind =
  2.676566, 2.237342, 5.129944, 7.198593, 6.214886, 5.142076, 5.013721, 
    5.342939, 6.598415, 5.693856, 5.622478, 6.245234, 5.875058, 4.904199, 
    3.53325,
  4.973601, 3.771099, 2.270533, 4.682699, 4.716466, 3.74073, 3.092965, 
    2.75934, 4.598237, 6.578317, 6.022286, 7.330775, 8.256284, 5.240748, 
    3.802712,
  3.855431, 4.546868, 4.164764, 4.210362, 5.43315, 3.403949, 2.89205, 
    2.496255, 3.092183, 5.056227, 5.617712, 6.300957, 7.660041, 7.941545, 
    6.479714,
  4.966655, 3.692921, 4.051068, 4.372036, 5.392989, 5.326138, 3.071459, 
    3.252526, 3.983122, 3.772166, 3.66767, 4.688342, 6.245932, 7.456203, 
    7.870568,
  6.941166, 5.303833, 4.264295, 4.282642, 4.536706, 5.419481, 5.606862, 
    3.205959, 3.065808, 2.628367, 2.589093, 3.915194, 5.625845, 7.472782, 
    8.621073,
  6.914999, 6.719146, 5.562489, 5.138032, 4.985198, 5.011254, 4.617621, 
    5.058997, 4.676475, 3.63218, 3.231067, 4.280926, 5.34482, 6.706551, 
    7.588317,
  9.013399, 7.674922, 7.054093, 6.491871, 6.205678, 6.325101, 6.473647, 
    6.381407, 5.742992, 5.384028, 5.266144, 5.39699, 5.844362, 6.443192, 
    6.876163,
  9.911755, 8.970157, 7.891126, 7.512885, 7.266252, 7.245043, 7.303005, 
    7.178771, 6.706326, 6.703771, 6.623506, 6.165756, 5.999803, 6.194599, 
    6.206333,
  9.474393, 8.770818, 8.020311, 7.724492, 7.492144, 7.401909, 7.316968, 
    7.447396, 7.518128, 7.371616, 7.084847, 6.765952, 6.731335, 6.728504, 
    6.175414,
  8.760885, 8.395451, 7.938554, 7.524782, 7.155605, 6.99757, 7.205554, 
    7.41612, 6.877507, 5.53698, 5.705801, 6.498296, 6.262331, 5.886835, 
    5.061543,
  2.257151, 5.220962, 2.838068, 5.205431, 7.995394, 8.675356, 12.3755, 
    12.16394, 9.63312, 6.776289, 7.7875, 10.9948, 11.65955, 11.14645, 9.620898,
  6.575763, 3.195955, 3.783875, 4.753549, 5.461802, 6.3886, 11.69327, 
    12.63624, 11.23887, 9.071395, 8.776546, 12.63033, 15.14775, 10.10787, 
    9.168555,
  9.825434, 8.260166, 5.910193, 6.02725, 5.475399, 4.058213, 8.986619, 
    11.64125, 12.21465, 10.91617, 10.77696, 12.52533, 14.3524, 14.37023, 
    11.27739,
  9.613156, 9.986547, 9.359886, 7.890607, 6.406147, 5.643474, 4.02662, 
    8.926245, 12.59436, 11.11136, 10.61069, 11.91677, 13.18163, 13.46354, 
    11.86341,
  8.719664, 9.149869, 8.963287, 8.571285, 7.586767, 7.009469, 6.3846, 
    4.072005, 6.221241, 7.142079, 9.444481, 11.08412, 12.78644, 13.3361, 
    12.57618,
  8.102984, 8.586874, 8.554405, 8.527715, 8.346902, 8.044715, 7.519625, 
    7.674266, 6.548102, 6.508625, 7.037171, 10.19614, 11.75675, 12.38341, 
    11.58002,
  7.718087, 8.182459, 8.219266, 8.237362, 8.095512, 8.13272, 8.097324, 
    7.947407, 7.666409, 8.414713, 9.074242, 9.720152, 10.88356, 11.79967, 
    11.81977,
  7.406002, 7.906741, 8.040468, 8.198955, 7.919717, 7.556585, 7.210545, 
    7.276116, 7.86842, 8.847655, 9.213075, 9.113804, 9.718444, 10.59703, 
    10.84272,
  7.047329, 7.428276, 7.635486, 7.996443, 8.128611, 8.19648, 8.190429, 
    8.373331, 8.649445, 8.615705, 8.546315, 8.317041, 8.571449, 9.340138, 
    9.252439,
  6.512143, 7.03782, 7.28215, 7.445424, 7.638267, 8.044954, 8.534299, 
    8.747893, 7.853069, 6.394479, 6.732209, 7.410385, 7.223111, 7.695226, 
    7.827901,
  5.2674, 6.090342, 4.273342, 4.695629, 5.963855, 6.601816, 9.700163, 
    8.839339, 4.408764, 4.888645, 7.647266, 9.11939, 7.477998, 6.660182, 
    5.65778,
  7.376053, 7.084338, 6.645313, 5.6377, 4.264649, 4.704199, 7.366572, 
    6.447047, 3.591378, 7.363238, 8.841674, 11.42346, 12.37407, 6.711712, 
    5.602903,
  7.002623, 7.223259, 7.447055, 7.105412, 5.579566, 2.889048, 4.97482, 
    4.887989, 5.290305, 9.661407, 11.16408, 12.30538, 12.62315, 12.27331, 
    8.131632,
  6.779916, 7.027283, 7.68712, 8.320389, 8.39426, 5.063607, 2.30301, 4.77946, 
    7.664616, 9.082118, 11.29782, 12.74012, 12.96855, 12.42451, 10.32566,
  7.003661, 7.18357, 7.739654, 8.730014, 9.6057, 8.085889, 5.086749, 
    3.858768, 4.708672, 6.181781, 10.56187, 12.95168, 13.85486, 13.73399, 
    11.98227,
  7.190763, 7.525041, 7.971897, 8.841977, 9.917504, 9.57567, 7.988483, 
    8.191723, 7.275955, 7.621949, 8.440189, 12.91563, 13.96324, 13.85624, 
    12.28858,
  7.590819, 8.147516, 8.477576, 9.163658, 9.901878, 9.979602, 9.673445, 
    9.855131, 10.36388, 11.52177, 12.55323, 13.404, 14.15667, 14.21286, 
    13.99304,
  7.690682, 8.564265, 9.11147, 9.726278, 10.06819, 10.18854, 10.45117, 11.34, 
    12.16793, 13.05649, 13.66135, 13.88352, 14.39873, 15.1386, 15.81145,
  7.743967, 8.592483, 9.317517, 10.08936, 10.42586, 10.41197, 10.68605, 
    11.79595, 12.81554, 13.49295, 14.13357, 14.40852, 15.1885, 16.49484, 
    15.8692,
  7.814574, 8.838723, 9.433667, 10.10335, 10.7061, 10.80058, 10.87085, 
    11.531, 11.3141, 9.841432, 11.23683, 14.59071, 15.215, 15.92125, 14.18395,
  6.447871, 7.524941, 5.377026, 5.605843, 3.546718, 4.462369, 8.367403, 
    9.377589, 8.617589, 5.697855, 5.959538, 8.122555, 6.950385, 5.233516, 
    3.040021,
  7.524348, 5.896281, 4.61349, 3.876809, 2.26205, 2.81425, 5.574991, 
    8.084692, 8.62747, 8.144123, 7.985967, 10.98124, 11.21346, 5.011013, 
    3.149437,
  6.077006, 4.283867, 3.865932, 3.927748, 3.240459, 2.807011, 4.499547, 
    7.008015, 9.320097, 10.77663, 11.45693, 12.13805, 11.06287, 8.004298, 
    4.837331,
  4.338677, 3.42979, 4.02746, 4.361959, 4.085223, 3.814719, 4.605927, 
    6.672979, 9.320237, 10.54159, 11.94661, 12.12127, 10.63051, 7.872997, 
    5.833707,
  3.107805, 3.288079, 4.085297, 4.329671, 3.96828, 4.846987, 9.073192, 
    6.597667, 6.34355, 7.193169, 11.26338, 11.68129, 10.17512, 8.067396, 
    6.273265,
  2.924794, 3.588563, 4.257727, 4.096549, 3.301427, 5.112312, 10.82116, 
    11.65729, 9.809886, 9.038532, 8.636379, 11.24989, 9.57517, 7.713228, 
    7.299282,
  3.108172, 3.866643, 4.332938, 3.621466, 2.941133, 6.060406, 10.66759, 
    11.48594, 12.27331, 12.94169, 12.5756, 11.21897, 9.468002, 8.899949, 
    10.09713,
  3.731552, 4.201309, 4.585914, 3.565553, 4.426233, 8.388972, 12.18073, 
    13.04066, 13.55182, 13.761, 13.02012, 11.20898, 10.19947, 11.06676, 
    12.36287,
  4.420626, 4.695058, 4.820432, 4.634914, 6.892412, 10.66267, 12.92259, 
    13.07367, 13.46644, 13.76475, 13.00175, 11.66208, 11.86162, 13.21751, 
    12.70554,
  4.693767, 5.056462, 5.263218, 6.935612, 9.315482, 11.67645, 13.21455, 
    13.63159, 12.586, 10.19555, 10.17276, 12.55049, 13.14847, 13.50118, 
    12.12362,
  6.325981, 8.535336, 7.156028, 8.130208, 4.946604, 3.856562, 8.939967, 
    10.14307, 8.974958, 6.010798, 5.467537, 6.258366, 4.408255, 2.792312, 
    2.056079,
  8.544291, 8.670268, 7.81982, 6.617763, 4.499989, 6.793281, 9.647645, 
    9.339651, 8.252845, 7.621101, 6.863775, 7.981449, 6.083217, 2.233597, 
    1.348033,
  7.892917, 7.673219, 6.197774, 6.376148, 8.280169, 6.66054, 7.824824, 
    8.572418, 8.987446, 9.30792, 9.303471, 8.356108, 5.227978, 2.933376, 
    2.071805,
  7.849223, 7.122646, 5.945812, 7.706151, 11.17471, 9.253628, 6.610838, 
    7.079964, 7.523088, 8.569442, 9.465666, 8.113613, 5.307953, 3.403818, 
    2.429037,
  8.026664, 7.136493, 6.356838, 7.939669, 10.44839, 11.81648, 11.78, 6.93401, 
    5.026925, 5.933441, 8.810946, 7.68448, 5.09288, 3.252682, 2.30711,
  7.995856, 7.40433, 6.731279, 7.801232, 9.22723, 11.02446, 13.07906, 
    12.26688, 9.225309, 8.261337, 6.971602, 7.685919, 4.953757, 3.11988, 
    3.113241,
  8.33755, 8.01079, 7.149076, 7.741569, 8.425085, 10.21242, 12.07219, 
    11.27063, 11.53649, 11.76125, 10.37759, 7.978199, 4.845638, 3.327373, 
    3.760747,
  9.004086, 8.522618, 7.219384, 7.366332, 8.171852, 10.60426, 12.94846, 
    12.6138, 12.71908, 12.15754, 10.71072, 7.910759, 4.674873, 3.887438, 
    4.306443,
  9.652769, 8.848811, 7.380692, 7.215401, 8.516116, 11.84339, 13.68478, 
    12.59656, 12.19985, 11.86709, 10.66808, 7.587941, 4.962209, 4.835042, 
    4.517015,
  9.903681, 8.538985, 7.028929, 7.673536, 9.786084, 12.6415, 13.79149, 
    12.84947, 11.31579, 8.714995, 7.878811, 7.371952, 5.691524, 5.308788, 
    4.424294,
  5.648944, 7.451566, 6.595611, 7.659402, 6.957153, 5.203731, 6.895168, 
    8.268055, 6.855992, 3.383074, 2.653455, 3.469206, 3.159338, 3.478807, 
    2.94666,
  7.869815, 8.445765, 8.713507, 9.067552, 6.369481, 5.176528, 7.400589, 
    7.656099, 5.889519, 4.048784, 2.698423, 3.797035, 4.388642, 2.820866, 
    1.782141,
  7.768455, 8.741469, 9.274922, 10.21344, 8.982773, 5.953169, 7.003803, 
    7.199245, 6.483496, 4.939179, 3.403181, 3.535324, 4.540225, 3.84253, 
    1.42375,
  8.141805, 9.059665, 9.545518, 10.89802, 12.88613, 10.00992, 6.201511, 
    5.616955, 4.704871, 4.431619, 3.403067, 3.140164, 4.077629, 3.665161, 
    1.837633,
  8.89572, 9.37854, 9.695147, 10.61628, 13.06314, 13.25169, 11.38473, 
    6.015388, 4.074206, 3.812463, 3.627328, 2.721015, 3.454533, 3.453539, 
    2.663993,
  9.692572, 9.641799, 9.672244, 10.3666, 12.69099, 13.40254, 12.7555, 
    11.70638, 7.921458, 6.358003, 4.037633, 2.381596, 2.592621, 3.203698, 
    3.366425,
  10.57005, 10.03754, 9.708907, 10.56092, 12.43096, 12.83623, 11.76435, 
    10.32878, 9.198935, 8.692348, 6.088489, 2.421711, 2.026601, 2.744389, 
    2.936467,
  11.02349, 10.1719, 9.70274, 10.85414, 12.54398, 12.49629, 12.07457, 11.788, 
    11.20112, 9.749838, 6.728385, 2.936096, 1.908122, 2.581881, 2.930777,
  11.27106, 10.30248, 9.952607, 11.28555, 12.69612, 12.39971, 12.10446, 
    11.68048, 10.85529, 9.645205, 7.402756, 3.751693, 2.025494, 2.305043, 
    2.577282,
  11.04034, 10.1821, 9.97564, 11.34453, 12.63061, 12.30932, 12.23036, 
    12.00477, 10.11852, 7.220146, 6.185321, 4.447738, 2.273983, 1.88907, 
    2.342562,
  4.865697, 6.946022, 6.659752, 7.505806, 6.493139, 4.50583, 3.923552, 
    3.803232, 4.072763, 3.807205, 4.5029, 3.919564, 3.122314, 3.640477, 
    3.138391,
  7.859253, 8.060833, 8.839211, 8.832809, 6.302575, 4.117329, 4.175149, 
    3.41256, 3.635052, 4.900749, 4.873224, 5.487565, 4.252197, 2.717789, 
    2.437264,
  8.577957, 8.598182, 9.484961, 10.02961, 7.932535, 4.025171, 4.044272, 
    2.976579, 2.731307, 3.933542, 5.861169, 6.042147, 4.908083, 3.722207, 
    3.336406,
  9.322439, 9.422224, 10.09943, 10.8244, 10.51439, 7.352609, 3.6781, 
    2.532501, 2.294263, 3.093576, 4.923769, 5.627968, 4.973802, 3.761924, 
    3.055209,
  10.53913, 10.4858, 10.89901, 11.47842, 10.78724, 8.982109, 7.367062, 
    3.067693, 2.53794, 2.292643, 3.247794, 5.076087, 4.816714, 4.126807, 
    2.782353,
  11.71333, 11.29907, 11.57267, 11.97376, 11.2571, 9.226321, 7.417449, 
    5.357789, 3.129664, 2.415121, 1.782175, 4.241781, 4.979162, 4.791076, 
    4.009931,
  12.67599, 12.215, 12.35065, 12.7049, 12.00957, 10.05194, 7.794874, 
    5.149667, 3.968252, 3.932776, 2.677155, 3.632612, 4.643477, 4.741834, 
    4.45203,
  12.94792, 12.73088, 12.81961, 13.19706, 12.63462, 10.64016, 8.589883, 
    7.21865, 6.432206, 5.038966, 3.09832, 2.716768, 4.277606, 4.623248, 
    4.440538,
  12.55187, 12.90599, 13.28834, 13.69524, 13.22708, 11.21588, 8.94953, 
    7.688651, 7.050154, 5.662179, 4.046185, 1.935966, 3.464253, 4.373347, 
    4.46021,
  11.93983, 12.59039, 13.1751, 13.59477, 13.2299, 11.31537, 8.767681, 
    8.029303, 7.682194, 5.419854, 4.442766, 2.194334, 2.191396, 3.465152, 
    4.08339,
  5.532729, 7.869373, 6.965435, 7.248662, 5.007086, 1.861451, 3.498797, 
    5.180386, 5.762467, 3.985022, 3.565114, 3.635799, 3.410076, 3.598775, 
    3.04056,
  8.692351, 9.978804, 10.16274, 9.027081, 5.458793, 2.150165, 2.780995, 
    4.400072, 5.292077, 5.036636, 4.095773, 4.66457, 4.93212, 3.237766, 
    2.679876,
  9.006564, 10.8081, 11.28459, 10.2476, 6.843683, 2.55808, 1.830363, 
    2.981696, 4.216638, 5.110519, 5.186659, 5.087273, 4.85446, 4.846385, 
    3.920353,
  8.646903, 10.92272, 11.78848, 10.97309, 8.614044, 5.314394, 2.336986, 
    2.855181, 3.981485, 4.298725, 4.915589, 5.190724, 5.03905, 4.786297, 
    4.252375,
  7.900221, 10.88533, 11.97751, 11.24175, 8.696708, 5.949118, 5.043592, 
    2.421004, 2.060235, 2.489384, 4.108311, 4.955101, 4.880614, 4.698464, 
    4.339772,
  7.364312, 10.7949, 11.93108, 11.19884, 9.150743, 6.488184, 4.372681, 
    2.714844, 2.729831, 3.39158, 3.609378, 4.779891, 4.608314, 4.077835, 
    3.246785,
  8.028172, 10.58799, 11.6433, 11.24037, 9.649682, 7.112318, 4.976859, 
    2.925723, 3.262817, 4.389073, 4.787179, 4.680481, 4.533529, 4.027202, 
    3.190645,
  8.864995, 10.33363, 11.26102, 11.2088, 10.19687, 8.14972, 5.688583, 
    4.055049, 4.133268, 4.792703, 4.890965, 4.729079, 4.714757, 4.41777, 
    3.769854,
  9.207134, 10.243, 11.18481, 11.36409, 10.726, 9.207776, 7.137011, 4.92128, 
    4.538311, 5.034261, 4.75001, 4.655538, 4.961062, 4.881531, 4.16797,
  11.30646, 11.12191, 11.21317, 11.45155, 11.10684, 9.853225, 8.191512, 
    6.33043, 5.333071, 4.657636, 4.402446, 4.652347, 5.018022, 4.986595, 
    4.335745,
  4.706368, 8.607952, 8.798394, 10.00335, 7.598094, 5.279632, 6.941613, 
    6.780446, 5.610685, 3.636719, 3.487492, 3.297128, 3.714339, 4.293313, 
    3.737277,
  5.393965, 9.687178, 11.89757, 11.49464, 6.851958, 4.507771, 6.845479, 
    6.841622, 5.465273, 4.201134, 2.976569, 3.255254, 3.641246, 3.098551, 
    3.00237,
  4.38359, 9.442265, 12.49169, 12.16739, 8.50324, 4.267771, 5.856414, 
    6.503351, 6.164331, 4.744919, 3.579711, 2.960504, 2.957498, 3.192905, 
    2.583782,
  4.580482, 9.290597, 12.56672, 12.31447, 10.71015, 7.545235, 4.362595, 
    4.606547, 4.2617, 4.484294, 3.758394, 2.784984, 2.521631, 2.631073, 
    2.478955,
  5.020181, 9.36693, 12.40666, 11.90942, 10.11958, 9.14231, 8.503239, 
    4.519539, 3.605686, 3.90701, 4.745904, 3.436862, 2.561419, 2.439025, 
    2.74065,
  5.16722, 9.50814, 12.04795, 11.34085, 9.588134, 8.449897, 8.604783, 
    8.472171, 6.05292, 5.275027, 5.041353, 4.552317, 2.930045, 2.525478, 
    2.683289,
  5.806234, 9.719622, 11.59535, 10.67478, 8.810568, 7.547213, 7.140622, 
    6.324478, 5.939044, 7.113808, 7.010445, 5.213098, 3.277083, 2.29127, 
    1.90135,
  5.72582, 9.446876, 10.81135, 9.930005, 8.276264, 7.074458, 6.523122, 
    6.374712, 6.916414, 7.601491, 7.005937, 5.618233, 3.745972, 2.358782, 
    2.072212,
  5.371377, 8.806076, 10.15647, 9.318643, 7.784125, 6.807949, 6.043951, 
    5.317929, 5.843452, 6.940423, 7.041921, 5.992015, 4.473422, 3.438213, 
    3.073272,
  6.160585, 7.876328, 9.300264, 8.953384, 7.664724, 6.621761, 6.029016, 
    5.416363, 5.647261, 5.387189, 5.987144, 6.207534, 5.140503, 4.49659, 
    3.948613,
  5.901932, 8.184597, 6.70495, 6.817003, 5.85981, 4.29058, 5.23857, 5.53484, 
    6.083797, 4.484345, 4.752928, 5.067269, 4.0532, 3.829602, 3.35907,
  9.213236, 9.503554, 9.356365, 8.175788, 5.426669, 3.788155, 4.943905, 
    5.219836, 5.590844, 5.775627, 5.097376, 6.60453, 6.779786, 3.848913, 
    3.394642,
  9.045356, 9.46045, 9.669355, 8.647976, 6.430966, 3.013605, 3.846889, 
    3.847132, 3.905388, 4.917331, 6.233069, 6.93413, 7.218227, 6.908862, 
    4.653176,
  8.799802, 9.466289, 9.605604, 8.509484, 7.296633, 5.226601, 2.38944, 
    3.387752, 3.913159, 3.81198, 4.935904, 6.198584, 6.754334, 6.932894, 
    5.694706,
  9.001707, 9.387442, 9.370314, 8.295838, 6.885045, 5.628635, 4.645867, 
    2.149518, 3.062454, 2.701612, 3.019207, 4.983314, 6.1453, 6.561931, 
    6.907558,
  8.876091, 9.236551, 9.239599, 8.231499, 7.206998, 5.910779, 4.709842, 
    3.716892, 2.430038, 1.905288, 2.328661, 3.699276, 5.232233, 6.177033, 
    7.15176,
  8.075912, 8.943159, 9.204719, 8.438302, 7.404428, 6.294295, 5.105021, 
    3.602925, 2.508403, 2.794819, 2.912813, 3.009692, 4.118124, 5.602052, 
    7.251866,
  7.109616, 8.495394, 9.023877, 8.506646, 7.710736, 6.942384, 6.150697, 
    4.70458, 3.534071, 3.47896, 3.379005, 2.81764, 3.377841, 4.836395, 
    6.278863,
  6.588718, 8.276615, 9.152003, 8.673676, 7.828351, 7.073381, 6.441782, 
    5.631338, 4.440187, 4.445053, 4.876651, 3.60818, 3.121245, 4.086595, 
    4.972872,
  7.456804, 8.054016, 8.939194, 8.805348, 8.053878, 7.227547, 6.637617, 
    6.1798, 5.608046, 4.959473, 5.400912, 4.682501, 3.641682, 3.629661, 
    4.108955,
  4.057718, 4.371275, 2.583485, 2.475929, 3.639771, 4.135655, 5.386626, 
    5.768576, 6.612471, 4.741183, 4.480164, 4.21019, 2.950642, 2.987876, 
    2.428247,
  6.228278, 4.617505, 3.064959, 2.304882, 2.33133, 3.898491, 5.703063, 
    6.055915, 6.789916, 6.554974, 5.012808, 5.560711, 4.942787, 3.210776, 
    3.072376,
  5.919842, 4.378007, 3.093019, 2.084568, 1.782703, 2.19023, 4.689634, 
    4.91202, 5.513291, 6.878586, 6.900951, 6.269884, 6.241178, 5.913092, 
    3.993778,
  5.833354, 4.431814, 3.399728, 1.997557, 1.40587, 1.695324, 1.763151, 
    5.070348, 7.712199, 7.662927, 7.60447, 6.966374, 6.751788, 6.658394, 
    5.361024,
  6.071954, 5.111403, 4.319631, 3.075709, 1.661733, 1.445701, 1.718597, 
    2.187094, 3.515337, 4.843382, 6.473742, 7.001587, 7.270809, 7.111843, 
    7.560399,
  7.513063, 6.697297, 5.876964, 4.677046, 3.117821, 1.399025, 1.643669, 
    2.990526, 1.624298, 2.617321, 4.317072, 6.173604, 6.969302, 7.510973, 
    8.47315,
  9.668384, 9.265064, 8.387494, 7.26918, 5.637989, 3.206583, 1.463917, 
    2.285893, 2.813554, 3.355157, 4.496603, 5.564673, 6.489243, 7.075838, 
    8.42579,
  11.39547, 11.53982, 10.93149, 9.607867, 7.860511, 5.932543, 4.202165, 
    3.15324, 3.586293, 3.70659, 3.610765, 4.652383, 5.772137, 6.71996, 
    7.737216,
  12.74179, 13.27917, 13.23897, 12.03491, 9.779819, 7.459118, 5.297348, 
    4.03539, 4.656116, 4.698279, 3.003331, 3.43322, 4.623632, 6.010536, 
    6.512589,
  10.11545, 11.7453, 12.61547, 12.84353, 11.54505, 9.010182, 6.624331, 
    5.468206, 5.928007, 5.03204, 3.944818, 3.272702, 3.348186, 4.426528, 
    5.709217,
  3.185826, 3.055042, 3.471933, 2.63087, 2.034699, 3.048089, 4.567438, 
    5.192883, 5.315899, 4.059145, 4.250091, 4.739316, 3.802477, 3.624555, 
    3.229285,
  5.394598, 3.540131, 1.932818, 1.44765, 1.414552, 1.892757, 4.212577, 
    4.996297, 5.373487, 5.458049, 5.1103, 6.792465, 6.849403, 4.021681, 
    3.837011,
  5.737999, 4.479711, 2.679182, 2.177775, 2.01553, 1.583456, 2.796303, 
    4.210442, 4.726451, 5.598093, 6.516964, 7.556244, 8.372944, 8.069737, 
    6.138281,
  6.437821, 5.411855, 4.379252, 3.606569, 2.508438, 2.805431, 1.821997, 
    3.815066, 5.464559, 5.756902, 6.345576, 7.372863, 8.594738, 9.102748, 
    8.004222,
  8.106486, 7.105046, 6.180076, 4.860508, 2.989393, 1.734942, 4.675584, 
    2.247838, 2.707774, 3.884666, 5.173265, 6.78941, 8.206013, 9.280378, 
    10.17847,
  10.83737, 9.498386, 8.259811, 6.471676, 4.735497, 2.520827, 3.651876, 
    4.102962, 1.059525, 2.204585, 3.622113, 5.758455, 7.519471, 9.036531, 
    10.81539,
  13.65419, 12.30894, 10.41555, 8.271766, 6.330012, 4.755146, 5.049638, 
    4.533054, 1.990492, 1.799071, 2.824561, 4.5877, 6.635709, 8.319914, 
    10.41706,
  11.21804, 13.10268, 13.07813, 11.36737, 9.074532, 7.144638, 7.012515, 
    7.083934, 4.88706, 2.432069, 1.915253, 3.251232, 5.392658, 7.328416, 
    9.565567,
  4.60875, 5.104574, 8.724586, 11.55767, 11.74736, 9.918619, 8.464067, 
    8.039197, 7.270212, 5.148034, 3.022098, 1.92587, 3.554624, 5.947112, 
    8.429029,
  5.540038, 4.502351, 3.325431, 5.258508, 9.687979, 11.10509, 9.941257, 
    8.68248, 7.785678, 5.764583, 4.813913, 2.726784, 1.816953, 4.148333, 
    7.104447,
  4.132129, 4.190121, 4.445381, 5.242248, 3.410038, 1.618947, 2.467774, 
    4.130494, 5.46928, 4.89977, 5.705835, 7.154598, 5.961607, 5.341382, 
    4.002805,
  7.236729, 4.574401, 2.974372, 2.521932, 3.092771, 1.774487, 2.069048, 
    3.413501, 4.889832, 6.028249, 6.836507, 9.555165, 9.542266, 5.07928, 
    4.593153,
  8.347221, 5.767514, 3.693038, 4.104083, 1.997216, 2.385365, 1.844831, 
    1.975224, 2.582121, 4.97908, 7.798064, 10.23283, 10.93173, 9.661461, 
    6.603491,
  8.720086, 7.366376, 5.184095, 4.739166, 2.774497, 3.692121, 1.55974, 
    2.319139, 4.30456, 5.328059, 6.905702, 9.183935, 10.95638, 11.06059, 
    8.624543,
  9.067961, 8.179012, 6.997211, 5.602832, 4.630503, 2.805287, 5.121317, 
    2.067151, 2.924722, 4.100009, 5.620687, 7.650841, 9.727874, 11.00855, 
    10.79067,
  10.6328, 9.281037, 8.231966, 6.70366, 5.562225, 3.164154, 4.393656, 
    5.007274, 3.440015, 2.901199, 3.905541, 6.046314, 8.158278, 9.975264, 
    11.03907,
  12.26688, 10.59166, 9.171172, 7.771753, 6.599313, 4.765627, 4.72074, 
    4.743708, 4.209733, 3.566037, 4.142251, 4.85421, 6.230748, 8.182841, 
    10.17257,
  12.17749, 11.4874, 10.45289, 9.425303, 8.519662, 7.1299, 6.562028, 
    6.745748, 6.642476, 5.960617, 5.242468, 4.383014, 4.525999, 5.877561, 
    8.096663,
  8.811747, 10.01343, 10.56852, 10.50257, 10.17618, 9.205239, 8.513628, 
    8.463898, 8.297946, 7.074645, 6.335875, 5.377788, 4.010439, 4.185956, 
    5.822001,
  5.614242, 6.755966, 8.06176, 8.928264, 9.627161, 9.617815, 9.465493, 
    9.229988, 8.074474, 5.927775, 6.33911, 7.293045, 5.763407, 4.377142, 
    3.999093,
  8.790821, 10.87337, 8.46753, 8.785545, 6.555889, 3.54414, 2.79087, 
    2.143156, 2.559009, 2.936082, 4.382288, 5.513359, 4.911601, 4.525085, 
    2.934867,
  12.28042, 11.11881, 10.16081, 8.855936, 4.731696, 1.740695, 2.071971, 
    2.324667, 3.472674, 3.847155, 4.50854, 6.382427, 6.880147, 4.29682, 
    3.539824,
  11.5064, 9.930027, 9.541972, 8.758312, 5.654658, 2.094641, 1.045757, 
    1.436186, 2.324188, 3.020412, 4.573555, 6.315518, 7.81246, 7.228889, 
    4.996949,
  10.33953, 8.739219, 8.396926, 7.843716, 6.390952, 4.623681, 1.753466, 
    1.895514, 3.333144, 3.056047, 3.977402, 5.842175, 7.632548, 7.73905, 
    6.041926,
  9.61808, 8.353555, 7.229459, 6.034119, 4.830643, 3.825262, 4.848138, 
    2.309733, 2.964124, 3.397388, 3.753645, 5.898321, 7.228621, 7.136908, 
    6.475379,
  9.157559, 8.37231, 7.231927, 5.838188, 4.61514, 3.576902, 4.036478, 
    4.589216, 3.992766, 3.78842, 4.012321, 6.477111, 7.250192, 6.302297, 
    5.4636,
  9.003205, 8.432755, 7.584352, 6.570775, 5.79601, 5.36318, 5.40706, 
    5.422512, 4.715438, 5.854287, 6.815829, 7.634896, 7.137312, 5.3649, 
    4.19745,
  9.252961, 8.697984, 8.199452, 7.631521, 7.456653, 7.466616, 7.685243, 
    7.623724, 7.432156, 6.981265, 7.907895, 7.823179, 6.482633, 4.563443, 
    3.507407,
  9.589992, 9.230744, 9.193387, 9.134091, 9.252168, 9.344498, 9.422462, 
    9.379038, 9.11223, 7.048235, 7.185032, 7.045774, 6.237112, 4.996377, 
    3.920979,
  9.955256, 9.843093, 9.929488, 10.12981, 10.40565, 10.63203, 10.7732, 
    10.45473, 8.285835, 5.697019, 6.571977, 8.016209, 7.074212, 6.35814, 
    5.282373,
  6.600402, 10.54861, 9.614014, 11.27806, 9.895319, 6.053406, 5.60976, 
    3.416738, 1.239037, 2.302795, 4.047443, 5.57227, 5.828889, 5.388053, 
    3.453009,
  10.25315, 12.41531, 13.29077, 12.61887, 7.921637, 4.503846, 4.859607, 
    2.786997, 2.440202, 4.134914, 4.760657, 6.778001, 7.864617, 4.61875, 
    3.090457,
  10.65678, 12.71357, 13.91716, 13.07893, 8.988732, 4.248497, 3.151658, 
    2.580873, 3.546522, 4.48299, 5.288293, 7.269625, 8.072322, 6.327062, 
    3.597196,
  10.72483, 12.59216, 13.63029, 12.7891, 11.02571, 7.111084, 2.670691, 
    1.308923, 2.363042, 2.057381, 4.402522, 6.980067, 7.753511, 5.378855, 
    3.608131,
  10.91134, 12.3572, 12.93251, 11.96897, 10.17422, 8.414868, 6.38381, 
    2.437881, 1.570135, 2.528992, 4.353723, 6.4067, 7.159794, 4.267031, 
    3.116444,
  10.99601, 11.92786, 12.16169, 11.1583, 9.852296, 8.293519, 7.125976, 
    5.185888, 3.034508, 3.780077, 3.916987, 5.769063, 6.433319, 4.17279, 
    2.136413,
  10.87025, 11.34649, 11.23286, 10.31251, 9.107751, 7.947078, 6.822543, 
    5.811627, 5.084004, 5.273932, 5.195084, 5.604811, 5.717566, 4.48113, 
    1.660885,
  10.28854, 10.4046, 10.00429, 9.152997, 8.284471, 7.46148, 6.952074, 
    6.623979, 6.408046, 5.483312, 5.52109, 5.420407, 5.346097, 4.662166, 
    1.969588,
  9.276164, 9.180963, 8.823153, 8.173213, 7.593825, 7.300504, 7.351593, 
    7.546215, 7.555023, 5.931969, 5.976445, 6.218277, 5.945007, 5.247193, 
    3.174367,
  7.804911, 7.570743, 7.384935, 7.308066, 7.412013, 7.714617, 8.177129, 
    8.451207, 7.099526, 5.002565, 6.039537, 7.670609, 7.142905, 6.473494, 
    5.11342,
  7.779065, 10.28309, 8.312889, 9.222607, 7.619728, 4.541872, 3.736452, 
    2.162892, 3.583177, 3.825232, 2.868859, 3.356904, 3.5267, 3.150054, 
    2.902898,
  12.2899, 12.23329, 11.41615, 10.28042, 6.139679, 3.602959, 3.353292, 
    1.81876, 3.885079, 5.13553, 4.070677, 3.441026, 4.651532, 3.175937, 
    2.862447,
  12.39379, 12.13965, 11.75815, 10.94002, 7.634396, 3.815625, 2.360785, 
    1.224043, 3.278378, 4.558833, 5.292083, 4.615663, 4.196691, 5.097429, 
    4.138512,
  11.78435, 11.49554, 11.32784, 11.05305, 10.22526, 6.982447, 2.836514, 
    1.493469, 2.283121, 3.139354, 4.644488, 5.715745, 4.725369, 5.17896, 
    4.868449,
  10.66312, 10.67112, 10.6809, 10.61881, 10.05158, 9.013443, 7.230655, 
    3.287742, 1.749566, 2.032218, 4.130989, 5.333416, 6.280163, 5.36647, 
    6.058136,
  9.701818, 10.09103, 10.26375, 10.30695, 10.13969, 9.365982, 8.448495, 
    6.895845, 3.541111, 2.189843, 3.199386, 4.779752, 6.064791, 5.506523, 
    6.188756,
  8.898491, 9.635915, 10.12279, 10.08555, 9.985076, 9.447248, 8.493336, 
    7.246181, 5.44777, 3.483685, 3.763382, 4.721004, 5.656883, 6.149603, 
    6.314033,
  7.980174, 8.985055, 9.796532, 9.902767, 9.893684, 9.6695, 9.039845, 8.3488, 
    7.315285, 5.038881, 4.236465, 4.599754, 5.51258, 6.243146, 6.028043,
  6.993393, 8.092615, 9.034041, 9.317954, 9.383353, 9.392653, 9.080052, 
    8.485266, 7.640584, 6.207294, 4.955919, 5.032342, 5.786574, 6.02323, 
    5.479634,
  5.520275, 6.512891, 7.290069, 7.694093, 8.040358, 8.284212, 8.358141, 
    8.083543, 6.943491, 4.755005, 5.18048, 5.648964, 5.739019, 5.9289, 
    5.294306,
  6.208655, 7.860638, 6.183523, 6.169946, 4.426025, 2.446849, 2.639277, 
    4.700215, 5.861772, 4.878762, 5.271228, 7.393245, 6.601018, 5.119331, 
    4.304044,
  9.865131, 9.415935, 8.619508, 7.147533, 3.93151, 1.526987, 1.788892, 
    3.801583, 5.694224, 5.957235, 5.967283, 9.262547, 9.981906, 5.22755, 
    3.367647,
  10.48023, 9.703243, 9.081619, 8.147436, 5.809135, 2.486163, 2.603033, 
    2.995728, 3.90908, 4.892782, 6.314673, 9.486029, 10.89107, 8.631336, 
    4.973754,
  10.69067, 9.884067, 9.260694, 8.520702, 7.9258, 5.899059, 2.390339, 
    2.928794, 4.307277, 4.220223, 4.992903, 8.241857, 10.38847, 9.385479, 
    6.088859,
  10.65756, 10.11478, 9.39032, 8.552647, 8.003577, 7.494781, 6.528172, 
    2.815077, 3.521907, 3.54797, 3.869617, 6.502421, 9.421911, 9.520658, 
    7.258307,
  10.12363, 10.11917, 9.403863, 8.693191, 8.341862, 8.076038, 8.114335, 
    7.539656, 5.486383, 3.608963, 2.646888, 4.944909, 8.195824, 8.918081, 
    7.747339,
  9.269541, 9.579055, 9.235055, 8.709579, 8.429191, 8.170969, 8.04326, 
    7.688241, 6.800319, 4.917179, 3.265575, 3.282548, 6.492876, 8.161367, 
    7.646123,
  8.511911, 8.787011, 8.793075, 8.638118, 8.513451, 8.222715, 7.930278, 
    7.395638, 6.781555, 5.766769, 4.886623, 3.087098, 4.474138, 6.565992, 
    6.924812,
  7.259303, 8.052204, 8.611817, 8.955153, 9.169142, 9.001657, 8.577769, 
    7.935912, 7.023608, 6.189635, 5.957713, 4.475176, 3.067577, 4.531682, 
    5.858045,
  3.855883, 4.996433, 6.162229, 7.064224, 7.714062, 7.922819, 7.865478, 
    7.56415, 6.338286, 4.79563, 5.92213, 6.060116, 3.799678, 3.045186, 
    4.270118,
  5.538321, 6.928534, 5.165935, 4.636313, 3.589536, 3.308949, 3.905955, 
    4.328326, 4.690073, 4.07587, 4.135221, 4.517647, 4.133694, 4.129585, 
    3.565378,
  8.694207, 7.691854, 6.034854, 3.427622, 1.794847, 3.520948, 4.731143, 
    4.703241, 4.700067, 4.500423, 4.262011, 5.11848, 5.078627, 3.102984, 
    2.628716,
  8.221943, 6.661803, 4.823211, 3.169821, 2.556093, 2.565756, 4.52587, 
    4.423487, 3.143924, 4.058448, 4.660714, 5.201233, 5.002546, 4.277793, 
    3.129071,
  7.231881, 5.590473, 4.308237, 3.800709, 4.172708, 4.120535, 3.147422, 
    3.954995, 3.147432, 3.835295, 4.576429, 5.096415, 5.170827, 4.116301, 
    3.174313,
  7.031541, 5.645036, 4.912419, 4.921131, 5.735627, 6.292629, 5.842523, 
    3.105677, 2.750785, 3.052114, 4.561458, 5.04932, 5.53528, 4.384102, 
    2.941453,
  6.977317, 6.516152, 6.371337, 6.623405, 7.291189, 7.601111, 7.012694, 
    5.882077, 3.720795, 3.406317, 3.903628, 4.755113, 5.844177, 5.00506, 
    3.053619,
  7.571508, 7.652897, 7.959709, 8.255311, 8.490312, 7.946927, 6.596362, 
    4.847347, 2.736068, 4.507984, 6.181194, 4.45472, 6.058308, 5.877079, 
    4.02465,
  8.804162, 8.378914, 8.41048, 8.473766, 8.265303, 7.019855, 5.232838, 
    3.736575, 2.683532, 4.288515, 6.726446, 5.042481, 5.728564, 6.514235, 
    4.923511,
  9.407605, 8.783781, 8.372358, 7.782663, 6.843114, 5.508269, 4.797223, 
    4.579159, 4.364179, 4.411908, 6.901412, 6.654984, 5.162101, 6.454079, 
    6.145304,
  7.515796, 6.328261, 5.440392, 4.669532, 4.095718, 3.837441, 3.875902, 
    4.043617, 4.05636, 3.97724, 5.931068, 8.112292, 5.994048, 5.279871, 
    6.199364,
  3.7332, 3.188526, 1.917853, 3.516217, 4.450903, 4.513604, 3.846476, 
    4.666885, 6.436342, 4.048989, 2.998586, 2.869503, 3.359715, 4.248571, 
    4.609026,
  5.846456, 3.298204, 1.77943, 3.03361, 4.148382, 4.995658, 5.6269, 3.923486, 
    6.521902, 5.794692, 3.784827, 3.451952, 3.643369, 3.541471, 4.511229,
  5.578584, 3.172982, 1.773531, 3.623852, 4.570025, 4.592739, 5.952552, 
    3.537456, 6.023265, 6.753618, 5.054025, 3.631426, 3.292591, 4.782893, 
    5.605975,
  5.404241, 3.278581, 2.852871, 4.856116, 7.266408, 6.425317, 4.372542, 
    3.216207, 3.263551, 6.761625, 5.724566, 4.014306, 3.26175, 4.670812, 
    5.573116,
  5.433076, 4.204302, 4.408788, 6.176658, 8.464708, 8.844225, 6.015908, 
    2.616592, 2.91746, 4.745517, 5.321003, 4.380907, 3.284158, 4.183375, 
    6.197893,
  5.965694, 5.686504, 5.80012, 7.05486, 8.530952, 8.57658, 6.243464, 
    3.533121, 2.25743, 3.083743, 3.817334, 4.457064, 3.497009, 3.736851, 
    5.64944,
  6.316249, 6.243423, 6.430296, 7.12244, 8.177827, 7.457987, 5.52041, 
    3.308109, 1.919146, 4.014184, 5.674351, 4.784585, 3.911544, 3.245439, 
    4.442399,
  7.984393, 7.284372, 7.122775, 7.477304, 7.889085, 6.358296, 4.445759, 
    3.064151, 2.826475, 4.507936, 6.134165, 5.389099, 4.249737, 3.016643, 
    3.379075,
  9.764737, 8.97428, 8.358998, 8.012813, 6.947641, 5.042644, 4.187864, 
    3.777682, 4.427526, 4.698042, 6.364714, 6.415745, 5.244319, 3.540995, 
    2.271768,
  10.40785, 9.566898, 8.42308, 7.227278, 5.601775, 4.879311, 4.642848, 
    4.496539, 4.442057, 4.221063, 5.815458, 7.491629, 6.839461, 4.976956, 
    2.447393,
  4.004686, 3.9972, 3.926405, 5.871718, 6.978483, 7.183959, 8.592108, 
    6.662881, 4.486709, 3.762302, 4.300552, 4.685695, 4.269891, 4.203556, 
    3.529917,
  7.432558, 5.794902, 4.989845, 5.8897, 5.396309, 6.106268, 8.134979, 
    6.92132, 5.505276, 4.849803, 4.438756, 5.074315, 4.403376, 3.489138, 
    3.278916,
  8.319006, 6.906734, 6.07531, 6.662998, 5.950323, 5.157122, 6.678599, 
    6.177904, 4.984344, 4.965694, 5.069549, 4.808229, 4.189233, 5.037021, 
    4.017788,
  8.717314, 7.672441, 7.114904, 7.361767, 8.833053, 6.741039, 4.735421, 
    5.367511, 6.31132, 5.603374, 4.514411, 4.035382, 3.934308, 5.106784, 
    3.928055,
  7.965442, 7.936872, 7.85575, 8.141917, 9.27262, 8.875995, 6.427486, 
    3.798233, 5.258554, 5.220373, 4.173136, 3.693727, 3.429929, 4.292402, 
    4.582441,
  7.251875, 7.476181, 7.864942, 8.342365, 8.772647, 8.718006, 7.947182, 
    6.049993, 5.169336, 4.438258, 3.510909, 4.13133, 2.977497, 3.197732, 
    4.098057,
  8.585588, 8.203096, 8.263187, 8.500107, 8.741938, 8.792173, 8.80838, 
    8.293805, 6.388485, 5.018813, 4.937958, 4.449498, 2.283275, 1.593873, 
    3.398224,
  10.02994, 9.565112, 9.44702, 9.375648, 9.520269, 9.516201, 9.122515, 
    8.343999, 6.675958, 5.572744, 4.776005, 4.080215, 2.147667, 1.124103, 
    2.753455,
  10.12261, 10.30658, 10.32753, 10.20971, 10.19173, 10.03105, 9.601027, 
    8.643242, 7.788082, 5.242677, 4.387582, 4.002018, 2.606608, 2.373556, 
    1.807525,
  9.240671, 9.853199, 10.2597, 10.57051, 10.8434, 10.55248, 9.591677, 
    9.296779, 6.62746, 4.02224, 4.584779, 4.041582, 2.873266, 4.081994, 
    2.100235,
  5.21099, 6.832413, 6.028667, 7.288939, 6.944037, 6.644565, 9.463963, 
    10.37342, 9.721254, 7.405952, 7.142209, 6.789349, 5.045526, 2.170166, 
    3.198397,
  9.13701, 9.640193, 9.494046, 9.713114, 5.763348, 5.774864, 9.868049, 
    10.54449, 10.31626, 8.500834, 7.108144, 7.587493, 5.663706, 2.397803, 
    4.46736,
  8.319671, 9.681117, 9.995657, 10.51609, 7.945249, 5.576315, 8.427629, 
    9.736564, 9.64211, 9.270798, 8.546647, 7.989081, 5.571936, 3.79693, 
    7.117565,
  7.023778, 8.357069, 9.371741, 10.29999, 10.90227, 8.621248, 5.733505, 
    6.61775, 8.122284, 8.564598, 8.487993, 7.955941, 5.133623, 4.219114, 
    8.631398,
  6.553926, 7.683639, 9.069385, 10.33825, 11.38407, 11.71075, 9.960735, 
    5.763523, 6.772356, 6.675237, 7.858179, 7.918599, 4.992414, 5.311128, 
    10.42083,
  6.912235, 7.971724, 9.484607, 10.90057, 12.0091, 12.83558, 13.01872, 
    12.2983, 8.912442, 7.263432, 6.78143, 8.05863, 5.00456, 5.793779, 9.951278,
  9.030939, 10.19122, 11.4454, 12.44734, 13.36172, 13.86631, 14.32468, 
    13.99535, 12.91015, 10.66728, 9.561544, 8.33426, 5.262682, 7.68783, 
    10.92901,
  10.98353, 11.92223, 12.73871, 13.09886, 13.82556, 14.12327, 13.55818, 
    12.86476, 11.92045, 10.00703, 9.117327, 7.601912, 6.121493, 10.05697, 
    12.49416,
  11.30817, 11.79304, 12.39173, 12.65334, 13.32368, 12.80299, 11.69232, 
    11.15589, 10.96466, 8.822965, 7.927328, 6.869347, 6.746801, 12.30256, 
    13.67844,
  11.17074, 11.2759, 12.03142, 12.93336, 13.18796, 11.00337, 9.625662, 
    10.24475, 8.881919, 6.30594, 6.512885, 6.333402, 7.595559, 13.65282, 
    13.42782,
  6.625301, 8.89212, 7.762812, 9.343493, 8.273619, 7.272513, 10.20242, 
    10.92672, 11.35407, 8.286463, 8.800984, 10.05715, 9.141253, 6.413385, 
    5.857602,
  11.10184, 12.00258, 11.83468, 11.82875, 6.744306, 6.225551, 10.95487, 
    11.0813, 12.19482, 10.82752, 11.37563, 13.4892, 11.75282, 6.688187, 
    7.140174,
  11.88845, 12.88545, 12.77495, 12.72132, 8.948559, 6.742779, 9.718802, 
    11.55487, 12.49443, 13.21125, 14.10242, 13.10239, 10.99843, 9.067344, 
    9.269227,
  13.14564, 13.50783, 13.33776, 13.10167, 13.04648, 10.38811, 6.174309, 
    7.634704, 11.5601, 12.82986, 12.53022, 10.33705, 9.426074, 8.110437, 
    12.27608,
  14.83334, 14.87486, 14.55936, 14.15139, 14.04841, 13.9235, 11.71986, 
    7.566143, 8.73385, 8.845694, 9.396373, 7.51696, 8.353271, 7.984799, 
    16.57927,
  15.78078, 16.24002, 16.06326, 15.56691, 15.24172, 15.12242, 15.08667, 
    14.58747, 10.03122, 6.683281, 4.61202, 6.281215, 7.817996, 8.154986, 
    17.41802,
  15.89349, 16.76593, 17.30622, 16.98684, 16.26775, 15.31625, 14.71073, 
    13.51446, 10.43163, 6.561673, 4.962882, 5.907629, 5.955707, 10.04854, 
    19.08859,
  15.50494, 16.3693, 17.20816, 17.122, 16.04718, 14.72211, 13.14512, 
    10.50895, 7.604319, 5.194164, 5.005634, 5.334955, 4.294208, 13.39679, 
    19.90398,
  15.78803, 16.1156, 16.29513, 16.08952, 15.34313, 14.1254, 11.85753, 
    9.233651, 6.788835, 5.104608, 4.974497, 4.271122, 5.723792, 17.44167, 
    18.82686,
  15.85969, 15.39067, 14.74842, 14.57602, 14.61853, 13.11474, 10.55615, 
    7.927144, 5.695101, 4.255054, 4.615034, 3.92905, 9.318294, 19.58301, 
    16.78276,
  9.933788, 12.65821, 11.24257, 13.80145, 12.30111, 10.08295, 12.54598, 
    11.56654, 10.57273, 7.667469, 7.511876, 8.302069, 8.129296, 8.534555, 
    6.823736,
  16.15931, 16.56067, 15.89706, 15.84477, 9.499352, 9.026053, 13.88717, 
    13.06617, 12.47969, 10.59854, 8.487925, 11.12936, 11.6029, 7.479361, 
    2.55328,
  15.4835, 17.55622, 17.14722, 16.82355, 12.34301, 8.675146, 12.11704, 
    13.85755, 13.45998, 12.26984, 12.2892, 12.11115, 10.7215, 5.914349, 
    3.309682,
  13.7468, 16.60781, 17.45683, 17.52727, 17.82786, 13.94304, 7.889194, 
    8.076578, 11.69442, 13.14598, 12.52414, 11.35028, 8.017682, 3.895845, 
    6.594779,
  12.15267, 14.20153, 16.06777, 17.17419, 18.1621, 18.51372, 14.7685, 
    8.730231, 7.611857, 8.051073, 10.17735, 9.59194, 5.900697, 4.94134, 
    8.950442,
  9.621774, 11.27717, 13.23008, 15.38003, 17.06361, 18.53966, 19.33559, 
    18.5282, 11.33856, 7.180701, 6.454403, 7.563016, 4.965694, 7.783786, 
    9.817017,
  7.978712, 8.655012, 10.13874, 12.26461, 14.48778, 16.51826, 18.21248, 
    18.66756, 16.13875, 12.36249, 10.16054, 7.253964, 7.470158, 10.66985, 
    11.75867,
  7.375381, 6.939651, 7.243153, 8.736205, 11.58589, 14.15222, 15.54365, 
    16.90335, 16.99602, 14.59442, 11.42233, 8.803438, 10.56639, 12.66793, 
    12.79961,
  7.669841, 8.342712, 8.449548, 8.015173, 9.424589, 12.14788, 14.49074, 
    15.75236, 16.25492, 15.90559, 13.44574, 11.72932, 13.44596, 14.57518, 
    12.67763,
  8.459513, 9.074997, 9.088686, 8.666931, 8.753317, 9.885716, 12.61034, 
    14.35803, 13.47221, 10.88045, 11.18572, 13.90406, 15.6469, 15.80281, 
    13.18674,
  10.53507, 13.81213, 11.94574, 14.3952, 12.73112, 10.17842, 12.92113, 
    11.11664, 9.548328, 6.529075, 5.274692, 5.081461, 3.634202, 2.739154, 
    2.182731,
  15.88103, 16.93533, 16.54018, 15.95482, 9.688957, 8.857731, 13.07265, 
    12.26188, 10.79427, 9.190517, 6.549015, 6.665135, 5.678386, 3.274041, 
    2.123763,
  14.51711, 16.92414, 17.12539, 16.95072, 12.38702, 7.468158, 11.18184, 
    12.92618, 12.55586, 10.66068, 9.277595, 8.236989, 6.963293, 5.707336, 
    4.160754,
  11.50323, 15.65891, 16.74015, 17.42009, 17.0694, 11.99293, 6.821496, 
    8.061968, 11.27119, 13.50099, 11.65208, 9.751763, 7.753398, 6.101208, 
    5.971642,
  4.800111, 12.37525, 15.17382, 16.45342, 16.83398, 15.63193, 12.92802, 
    8.206007, 7.456984, 8.786765, 12.1961, 11.90345, 9.43098, 8.065584, 
    8.629401,
  7.556304, 7.119095, 11.91586, 14.09033, 15.33095, 15.31718, 15.27237, 
    14.98405, 10.06956, 6.930941, 8.036343, 12.0801, 10.76402, 9.751755, 
    9.75551,
  11.18257, 7.292825, 7.969949, 11.25805, 13.42761, 14.13599, 14.1624, 
    13.62214, 11.94475, 10.55749, 10.73747, 10.97221, 11.14944, 11.41392, 
    11.37503,
  13.31545, 10.85856, 7.345004, 7.14051, 9.458675, 11.70789, 13.12237, 
    13.88353, 13.821, 12.61928, 11.03799, 10.44546, 11.52128, 12.06113, 
    12.64196,
  13.23089, 13.32898, 11.66756, 8.843334, 6.047236, 5.511981, 8.925636, 
    11.92062, 13.35341, 13.57493, 13.1056, 12.09149, 12.5753, 13.88732, 
    11.87183,
  10.99145, 11.42238, 11.36731, 10.74871, 9.464702, 7.189464, 4.998818, 
    8.141022, 10.02725, 9.570415, 11.05, 13.82693, 14.06514, 14.96818, 
    13.41595,
  8.795207, 12.3782, 10.89248, 13.71418, 12.61192, 10.3549, 13.1943, 
    11.38179, 9.047009, 5.209124, 3.878651, 3.363887, 2.812159, 2.923683, 
    2.908672,
  13.57544, 14.47375, 14.58335, 14.82623, 9.584759, 8.970145, 12.83235, 
    11.14922, 8.948199, 6.950897, 4.525833, 4.094559, 3.826272, 2.797491, 
    2.421081,
  14.05471, 14.63443, 15.32202, 15.64238, 11.73754, 7.908601, 10.26578, 
    11.25372, 9.197636, 7.852002, 6.289787, 4.660839, 3.808365, 3.942512, 
    3.802051,
  13.94312, 14.36011, 15.37662, 16.20254, 16.25041, 11.95909, 7.943214, 
    7.244525, 7.271747, 7.945628, 7.153072, 5.404304, 4.246294, 4.124661, 
    4.658284,
  12.78901, 13.7561, 14.86176, 15.85335, 15.79478, 15.06526, 13.60314, 
    8.286252, 5.778946, 6.321294, 8.165607, 7.062024, 5.470775, 5.08245, 
    5.468802,
  11.04743, 12.896, 14.12504, 15.1419, 15.4835, 15.11995, 15.32292, 14.94946, 
    9.743924, 7.137143, 7.198562, 8.634337, 7.022544, 5.930345, 5.518452,
  10.00281, 11.135, 12.74005, 13.94611, 14.36927, 14.13364, 13.92173, 
    13.12603, 11.91427, 11.57045, 11.51969, 10.12653, 8.581532, 7.280389, 
    6.559559,
  10.19691, 10.12998, 11.04492, 12.45471, 13.19777, 13.14301, 13.00797, 
    13.01015, 12.85564, 12.44147, 11.85908, 10.4292, 9.298297, 8.161758, 
    7.383453,
  11.15831, 10.26686, 9.981817, 10.82934, 11.82113, 12.27713, 12.41076, 
    12.09671, 11.74651, 11.4739, 11.02807, 10.45074, 9.405952, 8.903625, 
    8.04292,
  11.82749, 10.92708, 10.01278, 9.484623, 9.426197, 9.796538, 10.91043, 
    11.42128, 9.927733, 7.379477, 8.896763, 10.52864, 9.722097, 9.78341, 
    8.922286,
  9.452599, 12.98006, 11.6285, 13.74614, 11.21945, 8.323005, 10.39841, 
    9.045219, 7.354128, 4.862386, 4.209572, 4.464723, 4.251711, 4.472836, 
    3.95018,
  14.68249, 15.29392, 15.18658, 14.50186, 9.284927, 7.911421, 9.568761, 
    8.608979, 6.996227, 5.93079, 4.581549, 4.976616, 5.162025, 3.393904, 
    2.955565,
  15.65843, 15.90995, 15.74732, 15.16291, 10.55319, 7.731636, 7.76302, 
    7.647485, 7.589968, 6.457348, 5.883146, 5.090735, 4.775623, 4.110782, 
    3.120192,
  15.7864, 15.86171, 15.671, 15.11966, 14.49463, 10.68209, 7.240678, 
    6.459886, 5.947434, 4.614757, 5.072705, 4.649437, 4.386581, 4.128977, 
    3.533457,
  15.53266, 15.64848, 15.46731, 14.98409, 13.98057, 13.34422, 11.72714, 
    6.799212, 3.811605, 3.125094, 4.233134, 3.89051, 3.52036, 3.435049, 
    3.333896,
  15.19481, 15.19095, 15.03527, 14.55538, 13.93547, 12.97927, 12.02971, 
    11.04047, 6.953694, 4.986242, 3.9025, 3.738689, 2.898864, 2.619579, 
    2.61129,
  14.81435, 14.86941, 14.7503, 14.32115, 13.58946, 12.62997, 11.27038, 
    9.582026, 8.569566, 7.472483, 5.619496, 3.9083, 2.744471, 2.205692, 
    2.341427,
  14.33465, 14.34855, 14.22182, 13.92814, 13.3228, 12.35214, 11.18641, 
    10.34942, 9.994767, 8.680429, 5.91241, 4.007444, 2.755853, 2.246205, 
    2.374239,
  13.72146, 13.95815, 13.943, 13.61053, 12.97936, 12.15688, 11.19174, 
    10.09951, 9.495514, 8.352731, 6.295392, 4.728595, 3.320777, 2.583535, 
    2.408039,
  12.72478, 13.10186, 13.16407, 12.87173, 12.30914, 11.48973, 10.63854, 
    9.692298, 7.320133, 5.634081, 5.824599, 5.748517, 4.659431, 3.534706, 
    2.900959,
  8.821611, 12.31769, 10.91889, 12.86038, 10.02252, 6.705121, 7.797811, 
    6.838418, 6.829792, 4.689189, 4.53544, 4.800196, 4.31883, 4.469801, 
    3.947755,
  14.1002, 15.03809, 14.99109, 13.73376, 8.286025, 6.528049, 7.763775, 
    7.005268, 6.589719, 6.592489, 5.292912, 6.296979, 6.513326, 3.79323, 
    3.08339,
  15.51298, 15.78437, 15.20941, 13.27638, 9.417426, 5.962482, 6.610176, 
    7.226419, 7.431693, 6.928678, 7.032168, 6.816864, 6.865025, 5.400682, 
    3.295785,
  16.01206, 15.57276, 14.39143, 12.77821, 11.33545, 8.847858, 5.48155, 
    6.614786, 8.295982, 6.737206, 6.354203, 6.196559, 6.254618, 5.917451, 
    4.459803,
  15.89236, 15.08462, 13.54441, 12.17549, 10.63714, 9.866091, 8.73347, 
    5.114034, 3.683734, 3.748237, 5.405107, 5.957911, 6.099414, 6.15745, 
    5.76349,
  15.65649, 14.56016, 13.05368, 11.74521, 10.68734, 9.122016, 7.828803, 
    7.622077, 5.297106, 4.338067, 4.369934, 5.679711, 5.942047, 6.066928, 
    5.988472,
  15.17448, 14.17878, 12.96048, 11.78843, 10.61898, 9.733332, 8.56543, 
    7.376866, 6.768492, 6.00803, 5.178163, 5.336498, 5.786472, 5.984608, 
    5.962976,
  14.46385, 13.51296, 12.48295, 11.53366, 10.68401, 9.919669, 9.342472, 
    8.780301, 7.472868, 5.586813, 4.350157, 4.666945, 5.391687, 5.798042, 
    5.94753,
  13.98966, 13.12837, 12.21381, 11.18881, 10.35981, 9.577111, 8.726908, 
    7.862006, 6.530579, 4.198808, 2.948997, 3.542589, 4.680887, 5.480787, 
    5.507384,
  13.50019, 12.63887, 11.64283, 10.6234, 9.752617, 8.827191, 8.00005, 
    7.216578, 5.085736, 2.495184, 1.612204, 2.128819, 3.494503, 4.711443, 
    4.975122,
  6.728757, 8.147712, 6.170547, 6.799247, 5.704941, 4.880224, 5.902358, 
    5.139315, 5.369965, 3.555717, 2.672221, 2.823961, 2.475358, 2.263283, 
    1.219485,
  11.03688, 10.1212, 8.786245, 7.359347, 4.823533, 5.052986, 6.324285, 
    5.454534, 4.548089, 4.201579, 2.75328, 2.762166, 2.601413, 1.713213, 
    1.72956,
  12.3827, 11.12186, 9.588739, 7.516456, 5.782145, 3.898915, 5.880213, 
    6.28347, 6.118073, 5.070289, 3.999526, 3.133857, 2.641419, 2.422504, 
    2.123543,
  13.29441, 11.89831, 9.998307, 7.939179, 6.252542, 5.361948, 3.260715, 
    6.116264, 9.001148, 6.937958, 5.038215, 3.855915, 3.361399, 3.151822, 
    3.096666,
  13.93069, 12.5054, 10.48552, 8.830971, 7.104262, 6.040783, 5.534213, 
    3.859468, 4.419138, 4.70421, 5.775234, 5.449029, 4.844855, 4.581464, 
    4.610788,
  14.50081, 12.94758, 10.98328, 9.564906, 8.760123, 8.071887, 7.582042, 
    7.867118, 5.221982, 5.173984, 5.091115, 6.64377, 6.575989, 6.054911, 
    6.063668,
  15.11964, 13.5637, 11.73321, 10.30744, 9.303561, 9.088362, 9.097093, 
    8.970995, 8.714294, 8.694756, 8.147498, 7.800386, 7.445484, 6.974812, 
    6.829509,
  15.49419, 13.94308, 12.15519, 10.64832, 9.582995, 9.07359, 8.966394, 
    9.03823, 8.727248, 8.380873, 8.323791, 8.23402, 7.806643, 7.170681, 
    6.938352,
  15.55497, 14.17484, 12.66005, 11.07614, 9.805412, 9.103462, 8.609062, 
    8.14728, 7.362037, 6.406685, 7.636694, 8.296654, 7.964424, 7.547935, 
    6.777685,
  15.28154, 13.9483, 12.46241, 11.06001, 9.786561, 8.774542, 8.040922, 
    6.83439, 4.53103, 3.571654, 5.006527, 6.917425, 7.355923, 7.532188, 
    6.948447,
  2.877916, 3.887151, 4.358409, 5.219018, 5.125987, 3.933498, 4.422589, 
    4.066279, 3.946617, 3.118062, 3.024786, 3.201781, 3.427574, 4.051334, 
    3.923789,
  4.574678, 4.477252, 5.093381, 4.943259, 3.993018, 3.217078, 3.495749, 
    3.420838, 3.000762, 3.160627, 3.072101, 3.616342, 4.245287, 2.848728, 
    2.283664,
  5.453144, 4.988551, 5.161579, 4.788857, 4.436731, 2.8831, 2.556519, 
    2.87751, 3.632665, 3.648766, 3.570765, 3.51329, 3.574361, 3.303128, 
    2.77497,
  6.068575, 5.389724, 4.995412, 4.573144, 4.157423, 3.996412, 2.447966, 
    2.865775, 3.140942, 2.987136, 3.410201, 3.172933, 3.106349, 3.27422, 
    3.366542,
  6.255103, 5.311456, 4.642572, 4.860518, 4.581818, 4.386791, 4.829395, 
    3.106485, 2.432781, 2.629051, 3.312728, 2.789299, 2.640357, 3.063554, 
    3.509854,
  6.742918, 5.675108, 5.306985, 5.710961, 6.147413, 6.150396, 5.453024, 
    5.349364, 4.320163, 4.259852, 3.510707, 3.650672, 3.484182, 3.487159, 
    3.298296,
  7.626903, 6.969211, 7.04009, 7.374471, 7.448542, 7.836269, 7.713606, 
    7.24923, 6.960192, 6.748695, 5.917163, 5.269191, 5.013624, 4.637047, 
    4.016048,
  8.948431, 8.401247, 8.36723, 8.566689, 8.687982, 8.835045, 8.905384, 
    9.047201, 8.748063, 8.120332, 7.305586, 6.819829, 6.133954, 5.496637, 
    5.058713,
  10.34517, 9.777559, 9.673077, 9.543628, 9.553405, 9.775242, 9.861247, 
    9.802382, 9.420077, 8.744149, 8.186292, 7.742255, 6.93927, 6.160931, 
    5.751076,
  11.57132, 10.84821, 10.53247, 10.07726, 9.8829, 9.933119, 9.846784, 
    9.436724, 7.898309, 6.036477, 6.95455, 8.381855, 7.622452, 7.221158, 
    6.963759,
  3.335619, 4.470774, 4.240438, 4.475117, 4.404743, 3.656412, 4.307695, 
    4.945157, 6.081208, 4.609704, 4.137146, 4.379149, 4.53878, 4.615223, 
    3.663192,
  5.104657, 5.293906, 5.612199, 5.084558, 3.922319, 3.767744, 5.58571, 
    5.893099, 6.321672, 6.353576, 5.263125, 6.200865, 6.651719, 3.993236, 
    3.11519,
  6.093085, 5.862292, 6.258246, 5.651607, 4.881969, 3.391047, 5.123896, 
    6.239788, 7.04435, 7.132771, 7.258382, 6.98734, 7.069365, 5.985178, 
    4.283758,
  6.492162, 6.360064, 6.672876, 6.128659, 5.419173, 5.007086, 3.319345, 
    5.481227, 7.113928, 6.227323, 6.47865, 6.409046, 7.118417, 6.70739, 
    5.280425,
  6.309049, 6.368866, 6.675573, 6.663342, 5.698852, 5.427164, 5.721449, 
    3.501919, 2.826425, 3.196538, 5.173428, 5.659424, 6.515531, 7.043604, 
    6.241021,
  6.00472, 6.080722, 6.370679, 6.673189, 6.560117, 6.045398, 4.833586, 
    4.659303, 4.52387, 4.547173, 4.093446, 5.594453, 6.514779, 6.96488, 
    6.897085,
  5.49628, 6.112801, 6.659997, 6.842581, 6.745775, 6.799117, 5.843897, 
    4.935636, 5.962698, 6.091784, 5.652363, 6.026951, 6.635975, 6.838905, 
    7.421294,
  5.266018, 6.45886, 7.065618, 7.290513, 7.159855, 7.001899, 6.609081, 
    7.192396, 7.460733, 6.396111, 5.988758, 6.387019, 6.768728, 6.961679, 
    7.244202,
  6.233857, 6.781129, 7.282741, 7.737492, 7.827112, 7.68272, 7.212209, 
    7.383795, 7.258308, 6.232535, 6.040255, 6.433602, 6.614677, 6.409842, 
    6.276367,
  7.832005, 7.525564, 7.666486, 7.796147, 7.842931, 7.84158, 7.868649, 
    8.127973, 6.695982, 4.71712, 5.111824, 6.397648, 6.084348, 6.121185, 
    6.106122,
  2.727513, 3.057782, 2.41794, 1.614102, 1.070556, 1.344373, 1.845106, 
    3.387569, 3.627873, 2.347124, 2.639998, 3.669566, 4.852737, 5.349071, 
    5.263632,
  4.787024, 4.027852, 3.274884, 2.3795, 1.338347, 1.15243, 2.746649, 
    4.049634, 3.349849, 3.141841, 3.93171, 5.652477, 7.869774, 5.383318, 
    5.544972,
  5.800302, 4.758123, 4.084091, 3.597857, 3.541863, 2.168608, 3.242952, 
    4.555606, 4.826348, 4.607606, 5.934554, 7.274, 8.70306, 9.089025, 6.792384,
  5.839255, 4.787525, 4.250532, 4.435947, 5.194077, 5.141035, 3.571761, 
    4.254959, 4.587669, 4.453236, 6.733381, 8.143724, 9.258108, 8.752545, 
    7.420877,
  5.576928, 4.419581, 3.893764, 4.812487, 6.240184, 7.158648, 7.160936, 
    4.12572, 2.772563, 3.476779, 6.8266, 8.240338, 8.938691, 8.399037, 
    7.210883,
  5.835958, 4.199329, 3.567139, 4.569503, 6.695174, 7.511875, 6.948668, 
    6.925098, 5.686877, 5.928953, 5.977744, 8.414628, 8.409579, 7.936109, 
    6.888884,
  6.596471, 4.598547, 3.828641, 4.777802, 6.320497, 7.555854, 7.326709, 
    6.288394, 7.013359, 8.691356, 9.186293, 8.917722, 8.206024, 7.627962, 
    6.975707,
  7.031204, 5.470532, 4.50556, 4.962167, 5.860204, 6.641663, 7.308558, 
    8.009643, 8.761809, 9.192736, 9.427551, 9.031349, 8.093757, 7.439781, 
    6.734225,
  7.407891, 6.876673, 5.996043, 5.741712, 5.793577, 6.157464, 6.596757, 
    7.247196, 8.008742, 8.454264, 9.010232, 9.04809, 8.247993, 7.366148, 
    6.395943,
  7.071911, 7.25576, 6.71623, 6.238706, 5.799571, 5.756391, 6.326362, 
    7.334568, 6.877538, 5.821237, 6.786254, 8.737785, 8.092598, 7.340611, 
    6.065463,
  2.302125, 1.851819, 1.43337, 1.691342, 2.821304, 2.905954, 2.475193, 
    3.020563, 4.95934, 4.303277, 4.319345, 5.07442, 5.149148, 4.769101, 
    3.759285,
  4.739063, 3.616827, 2.412315, 1.511436, 1.163516, 2.656148, 3.461298, 
    3.600093, 4.990138, 5.762995, 5.622266, 7.177761, 8.256675, 5.00168, 
    4.465124,
  6.193068, 5.320297, 3.821065, 2.925823, 2.113084, 1.456936, 3.406395, 
    4.024582, 5.810246, 7.030046, 7.70363, 8.194421, 8.619103, 8.818347, 
    6.642051,
  6.804006, 6.302518, 5.159836, 4.158542, 4.140164, 3.680923, 2.364603, 
    4.352736, 5.78902, 6.133068, 7.670924, 8.103686, 8.545318, 8.763005, 
    7.892977,
  7.286888, 7.079848, 6.58071, 5.592402, 5.037032, 5.361502, 5.66861, 
    3.163067, 3.014385, 3.962035, 6.896755, 8.268991, 8.837288, 9.00011, 
    8.475509,
  7.603891, 7.391159, 7.330003, 6.611641, 5.831407, 5.834344, 5.295797, 
    5.904655, 6.131726, 6.150195, 5.943997, 8.27549, 8.476727, 8.073443, 
    6.993065,
  7.932022, 7.27595, 7.272453, 6.955346, 6.542816, 6.659534, 6.152423, 
    5.440571, 7.164161, 8.774301, 8.975342, 8.684999, 8.175191, 7.517272, 
    6.867205,
  7.65209, 6.693993, 6.514706, 6.553618, 6.734885, 7.141614, 7.672427, 
    7.74411, 9.04628, 9.599806, 9.044706, 8.639642, 7.784476, 6.970946, 
    6.329457,
  6.939447, 5.886223, 5.239722, 5.541336, 6.292967, 7.104992, 8.107007, 
    8.360312, 9.058558, 9.206329, 9.018354, 8.927591, 7.918163, 7.128999, 
    6.280744,
  6.156184, 5.009859, 3.903802, 3.960182, 4.915304, 6.042461, 7.509832, 
    8.810735, 8.05848, 6.597198, 7.559814, 9.487432, 8.642241, 7.841495, 
    6.766576,
  4.24707, 3.894601, 2.257605, 1.412062, 2.418081, 2.684268, 3.729996, 
    5.40864, 5.728465, 4.12135, 3.710292, 4.140296, 3.732939, 3.581819, 
    2.639356,
  8.12765, 6.287553, 4.109758, 2.954367, 2.078735, 2.182733, 2.738638, 
    4.900996, 5.494711, 5.157476, 4.463889, 5.383476, 5.670745, 3.448851, 
    2.755323,
  10.33105, 8.737659, 6.290479, 5.302821, 4.870192, 2.495605, 1.982876, 
    3.61882, 5.748445, 5.827265, 5.881162, 5.886376, 5.488771, 5.081911, 
    4.41057,
  11.70905, 10.31925, 8.457672, 6.828404, 7.219581, 6.255108, 3.200402, 
    2.874284, 4.292223, 5.46237, 6.106308, 5.568045, 4.932693, 5.041993, 
    5.623415,
  12.81311, 11.34177, 9.970357, 8.445135, 7.387453, 8.007514, 8.260699, 
    4.547458, 3.926958, 4.71793, 6.519042, 6.688731, 6.061857, 6.183039, 
    6.51305,
  13.5727, 12.16886, 10.83936, 9.274436, 7.57396, 6.111149, 9.093417, 
    10.30744, 7.611401, 6.44903, 6.466471, 7.923512, 7.025536, 6.41455, 
    5.949041,
  14.08243, 12.77255, 11.45234, 9.920246, 8.217665, 5.936601, 6.751862, 
    9.201102, 8.607762, 8.500299, 9.558154, 8.859536, 8.173466, 7.32053, 
    6.803397,
  14.10242, 12.61978, 11.36535, 10.1908, 8.88888, 7.12106, 6.104572, 
    7.712955, 9.149765, 8.956078, 8.876501, 8.931355, 8.661837, 7.889489, 
    7.344817,
  13.38115, 12.0087, 11.02439, 10.13095, 9.152685, 7.759895, 6.759411, 
    7.353514, 8.462098, 8.745256, 9.002451, 9.384735, 9.079586, 8.502905, 
    7.934688,
  11.8581, 10.80887, 9.990682, 8.969954, 8.243933, 7.219577, 6.477086, 
    6.94279, 7.350188, 6.579314, 7.762341, 9.787004, 9.474783, 9.361604, 
    8.47613,
  7.861219, 10.5078, 8.471923, 8.400023, 6.682885, 5.462821, 6.454357, 
    6.100238, 5.567243, 3.306887, 2.40759, 2.524601, 2.903514, 3.035965, 
    2.369992,
  12.62517, 13.22704, 12.46056, 10.48392, 6.135742, 4.325557, 6.030329, 
    5.75934, 5.084354, 4.414742, 3.101997, 3.356293, 3.722476, 2.903048, 
    2.515958,
  13.7513, 14.7249, 14.31552, 12.68136, 8.395199, 4.696376, 4.678191, 
    5.187902, 5.561729, 5.330248, 4.680349, 3.756874, 3.046133, 3.941985, 
    4.013772,
  14.32669, 15.53174, 15.44537, 14.62682, 12.93435, 8.589915, 4.747694, 
    3.435293, 2.637201, 5.240236, 5.310302, 4.241799, 3.399225, 3.822554, 
    4.871112,
  14.45116, 16.05655, 16.33157, 15.6313, 13.86455, 12.19911, 10.36315, 
    5.691713, 4.058506, 4.801772, 6.707791, 6.262732, 4.632974, 4.543796, 
    5.110238,
  14.08505, 16.17109, 16.81497, 16.18398, 14.60804, 12.85464, 12.27267, 
    11.49351, 7.336947, 5.568216, 6.701585, 8.143634, 6.276954, 5.205665, 
    4.583521,
  13.49644, 16.1312, 17.20774, 16.71897, 15.21474, 13.13933, 11.26567, 
    10.11699, 8.095286, 7.411946, 9.263832, 8.865833, 7.799305, 6.675035, 
    5.731863,
  12.27765, 15.29707, 17.11963, 16.93466, 15.59037, 13.58174, 11.26251, 
    9.902955, 9.419246, 8.843742, 8.69659, 8.580898, 8.261411, 7.652758, 
    6.772656,
  11.14595, 14.46136, 16.71124, 16.83452, 15.69238, 13.86314, 11.63424, 
    9.066199, 7.607964, 8.788702, 9.423533, 9.392904, 8.729736, 8.148793, 
    7.375465,
  9.550482, 12.98909, 15.63576, 15.93984, 15.07193, 13.63776, 11.61937, 
    8.308141, 5.834369, 5.739212, 7.644213, 10.06318, 9.610602, 9.158321, 
    8.066476,
  5.880562, 7.871939, 8.559533, 12.18568, 10.73283, 7.551363, 7.985775, 
    6.77611, 5.537259, 3.423825, 3.319194, 3.994794, 3.937322, 3.663971, 
    2.818582,
  8.382029, 9.589155, 11.22013, 13.06451, 8.473191, 5.651058, 7.6521, 
    6.743192, 5.300725, 4.45689, 3.800104, 5.020876, 5.765537, 3.504958, 
    2.935683,
  8.732265, 10.3868, 12.72569, 14.28921, 10.89351, 6.518816, 6.19315, 
    6.32078, 6.163787, 5.505935, 4.944619, 5.135676, 5.280081, 5.081861, 
    4.327011,
  8.631247, 10.54086, 13.77115, 15.75401, 15.44275, 10.9664, 6.69433, 
    4.40503, 3.296028, 5.060137, 5.050373, 4.901776, 4.837355, 4.9508, 
    5.269675,
  8.216253, 10.10795, 14.13444, 16.02445, 15.68628, 14.50348, 12.58171, 
    6.979485, 4.281396, 4.338681, 6.006359, 5.717394, 4.86169, 5.377679, 
    5.791367,
  7.993406, 9.435381, 13.91115, 15.94281, 15.80567, 15.08393, 14.66297, 
    13.06109, 7.54801, 5.775455, 6.06388, 7.001246, 5.644043, 5.120922, 
    5.01706,
  7.832979, 8.726234, 13.52898, 15.82017, 15.61249, 14.94724, 13.60779, 
    10.98956, 7.971509, 8.085602, 8.849312, 7.707707, 6.729415, 5.781129, 
    5.259496,
  7.020667, 7.584414, 12.65632, 15.48968, 15.3851, 14.603, 13.72872, 
    12.59349, 10.83363, 9.218384, 8.306968, 7.637958, 7.177593, 6.33272, 
    5.621321,
  5.649923, 6.157523, 11.53938, 15.08162, 15.04088, 14.37391, 13.61662, 
    12.40011, 10.34799, 8.445848, 8.114645, 7.95319, 7.461242, 6.895094, 
    5.935649,
  3.973242, 4.921639, 9.674673, 14.16089, 14.29818, 13.77507, 13.29327, 
    12.29614, 8.465993, 6.195182, 6.8126, 8.296908, 7.963631, 7.447773, 
    6.617007,
  5.839097, 7.767067, 6.047562, 8.16014, 8.389047, 6.858011, 8.918523, 
    8.824747, 7.849889, 4.907332, 4.257459, 4.700275, 4.332245, 3.822458, 
    3.123525,
  8.57812, 7.813663, 7.729199, 9.821604, 8.290367, 6.076345, 7.797724, 
    8.15948, 7.359007, 6.110617, 5.054885, 6.243737, 6.857506, 3.950485, 
    3.143384,
  9.900608, 7.370914, 8.703374, 12.52251, 10.64708, 6.789098, 6.474343, 
    7.229965, 7.674582, 6.851814, 6.458362, 6.531173, 6.5347, 6.245239, 
    4.849757,
  10.4972, 7.538527, 9.588696, 14.31067, 15.01069, 11.05813, 7.145831, 
    5.249508, 4.627479, 5.675888, 6.382882, 6.348921, 6.022473, 5.894065, 
    5.997695,
  9.857825, 7.175072, 9.06354, 14.13899, 14.86155, 13.90774, 12.71368, 
    7.19388, 4.194857, 4.342322, 6.510937, 6.731597, 6.415232, 6.547609, 
    6.578607,
  8.305125, 6.5877, 7.867459, 13.48471, 14.54837, 13.34579, 13.56544, 
    12.67198, 7.794148, 6.374915, 6.18995, 7.289944, 6.682051, 6.120767, 
    5.595904,
  5.672099, 5.25224, 6.219098, 12.86172, 14.40201, 12.93868, 11.71488, 
    9.769508, 8.350676, 9.261846, 9.066932, 7.861595, 7.076093, 6.15863, 
    5.58787,
  3.738698, 4.179608, 4.831912, 12.17375, 14.30728, 12.95924, 12.34227, 
    11.58175, 10.6146, 9.909423, 8.912461, 7.995789, 7.123761, 6.01428, 
    5.319082,
  3.130254, 4.366344, 4.399421, 11.86948, 14.13635, 12.96502, 12.4774, 
    11.53084, 10.33734, 8.777138, 8.348053, 8.068311, 7.26598, 6.141002, 
    5.261745,
  3.652116, 4.310866, 4.322384, 12.66872, 13.48687, 12.11084, 12.26486, 
    11.7888, 8.271675, 6.189666, 6.871573, 8.341354, 7.598471, 6.713354, 
    5.589857,
  8.895617, 11.38966, 8.437229, 8.980242, 5.85453, 4.797215, 7.165349, 
    8.685318, 9.496642, 6.152259, 4.874162, 4.739924, 3.610005, 2.940481, 
    2.718281,
  12.79487, 12.96796, 11.34474, 9.246323, 5.169561, 5.484601, 6.446891, 
    7.884461, 8.797247, 7.950727, 5.817205, 6.381366, 5.921828, 2.993968, 
    2.228096,
  11.50912, 12.07256, 11.53891, 10.7661, 8.332661, 7.602123, 5.812239, 
    6.428265, 8.347151, 8.636318, 7.682037, 6.959749, 5.89752, 4.802031, 
    3.591634,
  10.78272, 11.02136, 11.39592, 12.45963, 13.62328, 11.37059, 7.9446, 
    5.261195, 4.767939, 6.745978, 7.358379, 6.827299, 5.76002, 4.903977, 
    4.677398,
  9.663803, 10.40054, 11.07242, 12.66924, 14.51031, 14.50291, 12.71087, 
    8.289728, 5.069082, 5.230855, 7.314806, 7.401412, 6.655904, 6.010241, 
    5.314946,
  5.4956, 7.731597, 9.98372, 12.24633, 14.15051, 13.64473, 12.47402, 
    11.47059, 8.851384, 8.02397, 6.855247, 8.097767, 7.098215, 6.003314, 
    5.126198,
  2.54684, 4.237545, 7.729001, 11.44271, 13.75696, 12.41875, 9.129221, 
    7.125559, 9.310932, 11.48629, 10.0748, 8.735577, 7.600688, 6.394137, 
    5.689399,
  4.073161, 4.041876, 7.026491, 11.28358, 13.64359, 12.39177, 10.56406, 
    10.03975, 11.10972, 11.0615, 9.562682, 8.575883, 7.554519, 6.400938, 
    5.500429,
  5.368705, 5.658418, 7.867544, 11.95021, 13.60579, 12.06443, 10.71421, 
    10.69934, 11.34084, 9.716097, 8.813335, 8.267971, 7.362853, 6.392867, 
    5.272295,
  5.807045, 6.55253, 9.296298, 12.76416, 13.11293, 11.49898, 11.24824, 
    11.68311, 9.168622, 6.423991, 6.920878, 8.01168, 7.195494, 6.48683, 
    5.480461,
  9.291058, 12.6029, 9.72068, 11.29859, 9.830462, 7.362054, 8.742034, 
    7.910439, 7.81055, 6.245427, 5.82114, 6.334308, 5.197194, 3.533327, 
    2.995494,
  11.67847, 12.56745, 11.64202, 10.31243, 5.870804, 4.919988, 6.371441, 
    6.902138, 7.734049, 7.708408, 6.875756, 8.280399, 7.468118, 3.794744, 
    3.267843,
  9.08332, 10.18539, 10.596, 9.688328, 6.556779, 4.855489, 4.662786, 
    5.437953, 7.717808, 9.073013, 9.047544, 8.824284, 7.244364, 4.534768, 
    3.155366,
  7.839289, 8.524514, 9.525136, 10.26561, 10.41453, 8.062525, 6.287494, 
    5.128244, 4.979869, 6.755024, 8.511065, 7.955365, 6.137851, 3.429316, 
    2.466045,
  7.205176, 7.768897, 8.898479, 10.4172, 11.3647, 11.17158, 10.10961, 
    6.809333, 3.978314, 4.667311, 7.792432, 7.922721, 6.306642, 3.604276, 
    2.234044,
  5.135448, 5.317132, 7.815398, 10.49615, 11.88845, 10.96343, 10.04997, 
    9.58745, 7.125926, 6.965603, 7.141756, 8.548489, 6.697217, 3.627453, 
    2.214212,
  3.720038, 2.995456, 6.83181, 11.45037, 11.87531, 10.42301, 8.164786, 
    6.084878, 7.255379, 10.48711, 10.73178, 9.220748, 7.064221, 4.111246, 
    2.42021,
  4.525662, 4.006391, 8.51537, 12.11833, 11.50779, 10.14535, 8.81671, 
    8.219898, 9.059975, 10.51993, 10.22009, 9.176188, 7.078311, 4.452853, 
    2.974844,
  11.18315, 10.35657, 12.1575, 12.22811, 10.79515, 9.742363, 8.796161, 
    8.866441, 9.581351, 9.558532, 9.443902, 8.78937, 7.111765, 4.914725, 
    3.346168,
  15.72618, 14.60607, 13.19917, 11.69217, 10.55463, 10.35034, 10.64956, 
    10.78821, 8.928448, 6.748058, 7.247637, 8.431788, 6.941093, 5.148037, 
    3.639045,
  8.589997, 11.78567, 10.0555, 12.18091, 10.93116, 8.742011, 10.64785, 
    9.916585, 8.767631, 5.483337, 5.229387, 5.723007, 5.447008, 5.721446, 
    5.715511,
  11.5929, 13.7112, 13.7077, 13.22782, 7.594492, 6.703971, 9.822159, 
    8.844158, 8.311103, 7.037801, 5.685511, 7.407275, 8.260503, 5.675547, 
    5.141064,
  9.134246, 11.14571, 12.67955, 12.8151, 9.315285, 5.681967, 6.687533, 
    6.752685, 6.417387, 6.853599, 7.074884, 7.50953, 8.448064, 8.927131, 
    7.419007,
  7.92367, 8.435283, 9.386366, 10.50418, 12.03665, 8.716913, 4.013165, 
    3.181226, 3.471663, 4.726052, 6.151625, 7.18096, 7.810943, 8.376506, 
    7.987623,
  7.768876, 7.023847, 6.758883, 7.732458, 10.01978, 10.77923, 8.24627, 
    4.712191, 2.912263, 3.305221, 5.742612, 7.766065, 8.578366, 9.026924, 
    9.467457,
  8.026958, 6.629237, 4.766871, 4.721602, 7.286209, 9.039314, 7.932282, 
    7.077328, 5.747453, 5.27871, 5.786669, 8.64974, 8.842858, 8.27484, 7.5942,
  9.521709, 9.884056, 7.862948, 7.938314, 10.39852, 9.393473, 6.712989, 
    5.056853, 6.138112, 7.704525, 8.675035, 9.544795, 8.906872, 7.777997, 
    6.620601,
  9.171968, 10.70298, 11.74608, 11.92285, 10.6961, 8.724646, 7.630558, 
    7.811148, 7.778371, 7.67639, 8.721936, 9.435916, 8.222692, 6.625766, 
    5.230736,
  8.279612, 8.629157, 9.079409, 9.292394, 8.696535, 8.028303, 7.783595, 
    8.094641, 7.934926, 7.464917, 8.389536, 8.553215, 7.236615, 5.42321, 
    4.210852,
  9.51403, 9.460857, 9.243361, 8.917013, 8.542821, 8.141731, 8.344992, 
    8.312265, 6.763889, 5.415628, 6.555961, 7.809352, 6.354362, 4.13155, 
    3.657389,
  4.924578, 8.218732, 7.665888, 10.22308, 9.291537, 8.051071, 10.20482, 
    9.919801, 9.420779, 6.198598, 5.819244, 6.649394, 5.992643, 5.422652, 
    5.311869,
  4.712364, 7.123869, 8.710311, 10.18235, 6.763952, 6.801691, 10.05799, 
    9.172796, 8.810289, 7.581461, 6.409682, 8.067238, 8.446638, 5.423975, 
    4.793713,
  6.018211, 6.621734, 7.272404, 8.267639, 6.977053, 5.637906, 7.290514, 
    8.411089, 8.305216, 8.209365, 8.273726, 7.923851, 8.260628, 7.646031, 
    5.975302,
  7.110886, 8.343338, 8.297446, 7.132611, 7.996524, 7.014221, 3.947145, 
    3.494801, 5.256433, 7.730227, 7.902313, 7.068445, 6.711743, 6.818763, 
    7.054543,
  6.882226, 8.661888, 8.744613, 7.475801, 5.886613, 8.050939, 7.289742, 
    4.132585, 4.068218, 5.472119, 7.814561, 7.538503, 6.865985, 7.391201, 
    9.048898,
  6.253427, 8.661381, 9.426735, 9.349397, 7.296642, 5.802363, 5.80281, 
    4.755908, 4.210639, 4.723291, 6.479745, 8.211772, 7.675992, 7.749981, 
    8.702809,
  4.802395, 7.674612, 9.2999, 10.24239, 10.25261, 8.476569, 5.87923, 
    3.868314, 3.147388, 5.692359, 8.553767, 9.054599, 8.923697, 9.099156, 
    9.845649,
  3.735114, 5.886822, 7.553457, 8.544281, 8.772363, 8.291295, 7.579453, 
    7.283876, 5.980511, 5.638488, 8.120025, 9.492843, 9.794854, 10.18993, 
    10.43624,
  4.103688, 5.058459, 6.402925, 7.305828, 7.569199, 7.382584, 7.3166, 
    7.731902, 7.325851, 7.121349, 8.334328, 9.650839, 10.50718, 10.80243, 
    9.225475,
  5.148306, 5.288192, 6.032767, 6.820711, 6.936125, 6.431073, 6.383383, 
    6.604459, 5.640278, 5.014345, 6.750042, 9.667536, 10.47979, 10.50399, 
    8.6068,
  1.95126, 3.890397, 4.051109, 6.340527, 6.635725, 5.884193, 7.102674, 
    6.331611, 5.718166, 3.907724, 3.707589, 4.440774, 4.510697, 4.802792, 
    5.128998,
  1.769526, 3.281513, 4.447633, 5.645931, 4.275019, 4.691635, 6.945122, 
    6.373693, 6.035481, 5.593698, 4.790101, 5.63553, 6.571523, 4.523042, 
    4.5352,
  2.206552, 4.477715, 4.977884, 5.231035, 4.082056, 3.339027, 4.740393, 
    4.749286, 4.704863, 5.785641, 6.461643, 6.334168, 6.871462, 7.17376, 
    5.92737,
  1.969861, 4.398706, 6.527816, 7.318563, 5.658043, 3.605853, 2.392074, 
    3.187484, 3.720573, 4.900344, 6.06636, 6.188241, 6.313978, 6.724384, 
    7.244533,
  1.766885, 3.409473, 5.979143, 7.531456, 7.716484, 6.451503, 4.047099, 
    2.146026, 3.305344, 4.022179, 5.598476, 6.611527, 6.785377, 7.393089, 
    8.226617,
  2.470508, 2.939265, 5.46442, 7.371833, 7.892899, 7.405473, 5.982249, 
    4.300996, 4.43799, 3.859216, 4.019189, 6.051015, 6.858758, 6.993656, 
    7.319333,
  3.649887, 3.237666, 5.532919, 7.331959, 7.814179, 7.246213, 6.534157, 
    6.159909, 5.902369, 3.881433, 3.854581, 5.718704, 6.918921, 7.358212, 
    7.650434,
  4.196799, 4.030068, 6.416598, 7.516764, 7.732657, 6.993893, 6.082221, 
    5.950402, 5.647569, 4.024989, 3.68268, 5.865267, 7.199618, 7.901174, 
    8.293525,
  4.169679, 5.468691, 7.406497, 7.557376, 7.442039, 6.573332, 5.397388, 
    5.285844, 4.713102, 3.797276, 3.286231, 6.07333, 7.617061, 8.96474, 
    8.74495,
  5.296374, 7.82111, 8.597513, 7.720603, 7.167897, 6.21358, 4.338688, 
    4.059829, 3.152551, 2.286671, 3.198566, 6.610484, 8.616172, 9.653437, 
    8.51845,
  2.605921, 2.152991, 2.667245, 4.733387, 5.964045, 6.086497, 8.830505, 
    8.851597, 6.895988, 4.395713, 4.221075, 4.419935, 3.600956, 3.304041, 
    3.609279,
  3.967503, 3.060782, 4.043332, 6.257998, 5.386803, 6.337051, 9.039639, 
    9.378992, 8.286767, 5.508854, 4.569724, 5.076075, 4.771149, 3.155638, 
    3.102716,
  4.883531, 4.695889, 5.820492, 7.738281, 6.622588, 6.066204, 8.121935, 
    8.857442, 7.501038, 5.633254, 5.301751, 5.028364, 4.227845, 4.383569, 
    3.657127,
  5.051993, 5.955008, 8.491395, 11.17093, 11.52007, 8.760118, 7.145154, 
    6.51173, 5.978065, 5.476351, 5.283985, 4.543087, 3.434781, 3.594624, 
    4.314188,
  5.141493, 7.360495, 10.25823, 13.07317, 14.48495, 13.3618, 9.465333, 
    4.293832, 3.858016, 3.912107, 4.677895, 3.837749, 3.33803, 4.033847, 
    5.15419,
  6.537518, 9.169109, 11.9389, 13.99374, 14.61854, 13.00986, 9.094267, 
    5.639819, 3.797319, 3.758581, 3.287241, 2.518277, 2.402032, 4.338387, 
    4.97391,
  7.878586, 10.62354, 12.73755, 13.73209, 12.687, 10.12236, 7.938677, 
    5.098709, 3.666939, 4.572064, 3.155543, 1.473099, 1.757583, 4.831894, 
    5.528393,
  8.262756, 11.2311, 12.79678, 12.91387, 10.1517, 7.558726, 7.357684, 
    5.419947, 3.784616, 3.817076, 1.943574, 0.9700216, 2.655376, 5.023011, 
    5.88532,
  9.11334, 11.79431, 12.54489, 11.75776, 8.048891, 6.170735, 6.861265, 
    4.905568, 4.232346, 3.060604, 1.275396, 1.914632, 4.01428, 5.865089, 
    6.191621,
  9.620073, 11.26613, 11.43688, 10.61592, 7.250388, 5.604003, 6.091016, 
    3.278339, 3.314796, 2.395619, 1.560881, 3.050135, 4.746294, 6.057144, 
    5.730482,
  3.36732, 2.298503, 4.128647, 7.360623, 8.161851, 8.024634, 11.03662, 
    12.94737, 12.80564, 9.44072, 9.476556, 9.381746, 7.894847, 6.343388, 
    5.755483,
  3.05326, 4.09707, 6.818953, 8.70939, 7.010116, 7.46797, 10.52843, 11.25533, 
    11.40607, 10.35702, 8.728272, 9.287934, 6.870952, 4.606439, 5.24388,
  3.345664, 7.161252, 8.99044, 9.110828, 6.141913, 5.43284, 7.96771, 
    8.841794, 9.769118, 10.03628, 9.240612, 8.441886, 9.568735, 9.221061, 
    7.130671,
  5.735354, 8.31814, 9.355413, 9.501351, 7.326774, 4.098248, 4.029028, 
    6.614467, 10.14433, 10.15284, 9.145062, 9.825917, 8.899934, 7.672088, 
    6.020428,
  7.180729, 7.858589, 8.262321, 8.783969, 7.75483, 6.568194, 4.46289, 
    3.620692, 5.405038, 6.067145, 7.953315, 6.877335, 5.138144, 4.553028, 
    4.597962,
  7.092477, 6.553257, 6.954412, 8.028013, 7.528071, 6.568806, 6.288574, 
    4.847325, 3.785006, 4.761351, 4.66331, 5.18966, 3.216179, 3.274454, 
    4.389734,
  6.538945, 6.017395, 6.542206, 7.480423, 7.250793, 6.50151, 6.302023, 
    5.407474, 5.128536, 5.694758, 5.065716, 3.987578, 2.949985, 4.077959, 
    5.235933,
  5.991771, 6.407711, 7.070031, 7.723953, 7.494708, 6.845462, 6.316929, 
    5.400907, 4.552996, 4.438726, 4.038702, 3.466898, 3.225496, 4.288692, 
    4.79916,
  5.381413, 6.362178, 7.367427, 7.923941, 7.50081, 6.759041, 6.51658, 
    5.525671, 4.060938, 3.658225, 3.424579, 3.083719, 3.485289, 4.12358, 
    4.018316,
  4.759393, 6.104749, 7.458272, 8.288696, 8.233918, 7.360497, 6.770483, 
    6.004455, 3.867804, 3.482753, 3.233229, 3.349771, 3.362241, 3.635033, 
    3.099082,
  4.97754, 5.372701, 3.099575, 3.802004, 4.489738, 5.195583, 7.567156, 
    7.399602, 5.28963, 4.298879, 5.276932, 7.665074, 6.493046, 4.04879, 
    2.420708,
  7.631038, 4.996937, 2.834424, 3.59098, 3.373286, 4.983339, 7.767824, 
    8.191584, 6.044715, 5.225369, 5.015223, 8.278605, 9.412121, 5.016244, 
    2.856391,
  8.248001, 4.964729, 2.694964, 3.296103, 3.160893, 4.147873, 7.206414, 
    7.497314, 4.826772, 4.75615, 4.51346, 6.683093, 8.340954, 7.848657, 
    5.369947,
  7.573234, 4.239823, 2.51434, 3.535111, 4.098195, 4.028389, 5.00175, 
    6.608928, 7.003411, 3.773843, 4.675604, 4.241382, 5.67295, 6.525344, 
    5.556519,
  6.374149, 3.214161, 2.700632, 4.26806, 5.613776, 6.391734, 6.427222, 
    5.082153, 5.782652, 3.384846, 5.294734, 2.86115, 3.176065, 4.254694, 
    4.690302,
  4.808226, 2.295161, 2.865, 4.714081, 6.403734, 7.692542, 8.429973, 
    8.873991, 7.979944, 4.228271, 4.622608, 4.094793, 2.568057, 2.860465, 
    3.575516,
  4.235516, 3.046867, 3.362824, 4.585654, 6.420014, 7.820775, 9.439979, 
    10.25758, 11.64391, 7.378737, 6.221971, 5.429905, 3.94698, 3.492823, 
    3.086294,
  4.096029, 3.128742, 3.654599, 5.323676, 6.706697, 7.586792, 8.970536, 
    10.2316, 11.66951, 9.837398, 7.146096, 6.690623, 6.171566, 5.278289, 
    3.838128,
  3.428097, 2.586069, 3.92366, 5.92962, 6.962903, 7.051828, 8.778952, 
    10.47261, 11.78475, 10.04272, 8.100296, 7.686262, 8.059292, 7.02034, 
    5.354798,
  2.576032, 2.800481, 5.039061, 7.055212, 7.865094, 8.051758, 8.481507, 
    9.964593, 10.07739, 6.96226, 6.988136, 9.160413, 8.72201, 8.604092, 
    7.039433,
  6.461444, 5.995696, 2.963517, 4.262152, 4.536984, 4.63354, 6.520946, 
    3.150526, 1.734185, 2.008384, 4.06732, 5.01922, 4.229353, 4.333174, 
    4.080698,
  8.99523, 5.595871, 3.656477, 3.865836, 3.244337, 4.17437, 7.554466, 
    6.580654, 1.714878, 1.108767, 2.596858, 4.758885, 4.641344, 2.983372, 
    2.734708,
  8.894064, 5.476086, 3.856565, 3.259222, 2.81267, 2.78745, 6.058961, 
    7.136121, 3.611036, 1.703856, 1.8589, 3.082912, 3.943363, 3.73033, 
    2.846953,
  7.897395, 4.995766, 3.736276, 3.370725, 2.442301, 2.162895, 3.124631, 
    5.530218, 7.959625, 3.158257, 2.976697, 2.757921, 3.136174, 3.10453, 
    2.870035,
  6.522305, 4.024882, 2.940112, 2.592863, 2.283457, 3.291406, 3.406497, 
    3.411052, 5.28479, 3.858845, 3.608674, 4.013934, 4.235393, 3.56607, 
    3.283715,
  5.231599, 3.16124, 2.261882, 1.930981, 2.571181, 3.868414, 4.7988, 4.7023, 
    5.197456, 5.51382, 3.828821, 4.204152, 5.642905, 5.344779, 4.388505,
  4.32422, 2.922448, 2.175699, 2.272446, 3.804487, 4.970246, 6.009185, 
    5.950684, 6.962451, 7.84767, 7.176057, 4.634639, 5.499825, 6.631464, 
    6.147568,
  4.561878, 4.037528, 3.933532, 4.607664, 5.934269, 6.544913, 6.680161, 
    6.634634, 7.127656, 7.942959, 7.889876, 5.850307, 5.196702, 6.984777, 
    7.363868,
  5.633444, 5.815431, 6.072745, 6.53737, 7.166964, 7.661928, 8.057818, 
    7.937157, 8.068979, 8.305924, 8.138157, 7.29882, 5.676492, 6.613069, 
    7.28002,
  7.001377, 7.120262, 6.877158, 7.946825, 8.7561, 9.249374, 9.165827, 
    8.424098, 7.76005, 6.300441, 6.731203, 8.020354, 6.941205, 6.011815, 
    7.102108,
  8.065275, 8.646607, 5.933161, 5.357009, 3.889817, 2.772856, 3.312241, 
    3.961234, 4.837741, 3.772869, 3.648563, 3.806012, 3.285856, 3.099118, 
    3.201274,
  10.8015, 9.033883, 6.302083, 4.447338, 2.864153, 2.103127, 2.885189, 
    3.791091, 4.829357, 5.420571, 5.216301, 5.813585, 5.649034, 3.85088, 
    3.672226,
  10.42886, 8.46696, 6.364297, 3.978868, 2.636075, 2.077927, 3.666857, 
    5.011136, 5.5253, 6.304181, 7.217472, 7.717963, 8.10497, 8.278874, 
    6.058067,
  8.917574, 7.344297, 6.054513, 5.043814, 4.670925, 4.157118, 3.679348, 
    5.147419, 6.549631, 6.861212, 7.458726, 8.568681, 9.25921, 9.504897, 
    8.438663,
  7.064256, 5.960095, 5.832644, 6.470734, 7.661632, 8.382626, 7.03648, 
    4.924456, 6.157115, 5.886672, 7.950924, 9.601405, 10.13413, 10.55552, 
    10.91035,
  5.683478, 5.638901, 6.889125, 8.323494, 9.776981, 10.72546, 11.18878, 
    10.76433, 9.935609, 8.288198, 8.049425, 11.47964, 11.74066, 11.8857, 
    11.77859,
  5.888927, 6.983333, 8.765258, 10.17808, 11.60277, 12.56751, 13.4185, 
    13.72743, 13.70856, 13.63859, 13.51841, 13.62643, 13.32716, 12.78143, 
    12.6909,
  7.755212, 9.411577, 11.11612, 12.32632, 13.68209, 14.62486, 15.11186, 
    15.3877, 16.06118, 15.73315, 15.82093, 15.21832, 14.51656, 13.63211, 
    12.99297,
  10.70226, 12.26831, 13.59181, 14.53593, 15.22424, 16.10616, 17.05745, 
    17.41052, 17.45589, 15.64286, 15.55822, 15.61883, 15.02923, 13.63632, 
    11.65026,
  13.39646, 14.65394, 15.8561, 16.3577, 17.20862, 17.74561, 18.69611, 
    16.92273, 15.87807, 10.97716, 11.5425, 15.25607, 14.16348, 11.02382, 
    9.505904,
  4.589754, 7.08382, 5.952003, 6.647703, 5.555925, 4.90057, 7.311667, 
    8.610833, 9.344582, 7.667127, 9.15028, 10.51501, 10.26118, 9.541093, 
    9.827024,
  7.633014, 7.913537, 7.207823, 6.096901, 3.830373, 4.069031, 7.352252, 
    8.664817, 11.04484, 10.74454, 10.18261, 12.20675, 13.0843, 9.831044, 
    10.31079,
  8.524915, 8.453454, 7.694353, 6.701498, 4.812936, 3.518308, 6.933348, 
    9.043306, 11.5895, 13.33203, 13.5577, 14.2273, 14.23368, 14.56336, 
    12.73197,
  8.746974, 8.595675, 8.188046, 7.993624, 8.118217, 6.090369, 5.666656, 
    8.324142, 11.97648, 12.24062, 13.87514, 16.04006, 16.02773, 16.28972, 
    14.59611,
  8.793663, 8.431553, 8.325192, 8.615528, 9.688123, 10.59728, 9.368897, 
    8.193244, 11.00892, 10.29006, 15.15225, 17.38431, 17.48172, 18.01437, 
    18.15504,
  8.750056, 8.482159, 8.733485, 9.446156, 10.67778, 12.1433, 13.48311, 
    14.0825, 14.55972, 12.66253, 12.2297, 17.43657, 18.46261, 19.24906, 
    19.29802,
  8.486227, 8.825687, 9.598787, 10.54722, 11.84281, 13.4142, 15.03031, 
    16.8589, 17.78467, 15.68351, 16.04142, 17.70607, 18.83356, 19.46054, 
    20.01875,
  8.183181, 9.175594, 10.39141, 11.55324, 13.04301, 14.61801, 15.50814, 
    15.90091, 15.61952, 15.154, 16.25766, 17.84289, 18.95739, 19.70515, 20.482,
  8.386169, 9.806472, 11.30004, 12.64402, 13.94754, 14.92912, 15.92788, 
    14.83153, 13.59725, 14.61379, 15.70954, 17.61357, 18.69223, 19.64177, 
    19.41017,
  9.425107, 10.81575, 12.53734, 13.79062, 15.14483, 14.79, 13.31916, 12.312, 
    11.09076, 9.819706, 12.07896, 17.52671, 18.77538, 19.72611, 18.56501,
  4.907539, 6.944307, 6.425174, 8.459392, 7.383606, 6.191475, 8.284791, 
    8.061208, 7.860134, 6.2276, 6.497819, 7.202978, 6.5139, 5.725469, 5.596255,
  7.284283, 8.05917, 7.778505, 7.813025, 4.851676, 4.656235, 8.06778, 
    8.01769, 8.732933, 7.99911, 7.618636, 8.896794, 8.17002, 5.791728, 
    5.977933,
  8.16967, 8.787725, 8.691195, 8.8709, 6.434834, 3.651825, 6.38932, 7.962315, 
    9.498778, 10.02045, 9.741449, 9.420407, 8.59265, 8.63098, 7.024489,
  9.032202, 9.450165, 9.741198, 10.17743, 10.94883, 7.93666, 3.636772, 
    4.804811, 7.095157, 8.716683, 9.426886, 9.285622, 8.24012, 8.203367, 
    7.238749,
  9.695542, 9.650736, 9.874179, 10.1305, 10.83536, 11.767, 9.794992, 
    5.335646, 5.335075, 5.629405, 8.265936, 8.681805, 8.548452, 9.156713, 
    9.693992,
  10.03445, 9.906662, 10.03547, 10.12955, 10.45042, 11.25704, 12.50634, 
    13.04246, 10.26301, 8.831516, 7.895225, 10.61472, 11.02504, 11.19607, 
    11.47012,
  9.756432, 9.752199, 9.928717, 10.01798, 10.40428, 10.86546, 11.73826, 
    12.83747, 13.23845, 13.29863, 12.56344, 11.96219, 11.52672, 11.44749, 
    11.53214,
  8.760397, 8.936779, 9.338573, 9.758771, 10.43108, 11.06172, 11.6159, 
    12.17061, 12.61485, 12.53203, 12.59248, 11.828, 11.69479, 11.51533, 
    11.75812,
  8.04698, 8.006783, 8.317191, 8.549935, 9.252556, 10.074, 11.25757, 
    12.27521, 12.36997, 12.58703, 12.82486, 12.30455, 11.73081, 11.6769, 
    11.39631,
  7.328394, 6.654385, 6.442967, 6.752027, 7.659811, 9.253445, 10.95024, 
    11.63048, 11.00762, 8.800835, 9.969233, 12.59687, 12.28914, 12.06994, 
    11.4049,
  5.632582, 8.013103, 7.070198, 9.111292, 8.102086, 6.310418, 8.084504, 
    7.28156, 6.043377, 4.397289, 4.484409, 5.106802, 4.487449, 4.345492, 
    5.137443,
  8.116549, 8.807858, 8.867144, 9.215082, 5.750497, 4.862683, 7.093439, 
    6.203499, 6.059912, 5.663074, 5.413603, 6.895892, 6.928577, 5.188092, 
    5.719394,
  9.644295, 9.295216, 8.913316, 8.783309, 6.000756, 3.928626, 5.385315, 
    5.49767, 6.077214, 6.764528, 7.287745, 8.040941, 8.477276, 8.783764, 
    6.674435,
  9.657825, 9.454304, 9.464175, 9.277369, 7.961195, 5.725778, 3.380029, 
    3.642488, 5.15096, 6.280447, 6.6518, 6.9691, 6.840179, 6.952892, 6.342839,
  8.97808, 9.258945, 9.363728, 9.035834, 8.55458, 7.697242, 6.486232, 
    3.465809, 3.790431, 4.352829, 5.289487, 5.694154, 6.619588, 7.225214, 
    7.493439,
  9.012897, 9.505297, 9.199256, 8.495121, 7.773428, 6.970999, 7.233263, 
    7.491719, 5.62365, 4.631305, 4.235062, 7.079431, 7.928417, 8.005767, 
    9.032051,
  10.05647, 9.791106, 8.830452, 7.459492, 6.632951, 5.809059, 6.125558, 
    6.498305, 5.710815, 5.480597, 6.518417, 7.537048, 7.490439, 8.235303, 
    9.575067,
  10.43816, 9.096024, 7.564416, 6.442621, 5.630524, 5.399734, 5.292477, 
    4.844778, 4.320035, 5.978598, 6.961492, 6.693306, 7.361582, 8.665261, 
    10.05957,
  9.536826, 8.136032, 6.661068, 5.089463, 4.367864, 4.312202, 4.639758, 
    4.170678, 5.391892, 6.303363, 6.734145, 6.825578, 7.80101, 9.214664, 
    10.24604,
  7.905557, 6.456662, 5.172566, 4.064262, 3.847535, 4.497144, 4.121133, 
    5.08877, 5.565697, 4.598684, 5.642163, 6.910814, 7.740183, 9.324182, 
    9.993925,
  3.966881, 5.757541, 5.624527, 8.527819, 8.726269, 7.955436, 10.16301, 
    10.20953, 8.279534, 4.703174, 4.332859, 4.392266, 3.763209, 3.517688, 
    3.985496,
  5.444806, 6.126239, 7.022631, 8.609432, 6.617291, 6.614872, 9.994211, 
    9.837117, 8.58295, 5.966787, 5.022641, 5.526935, 5.498663, 4.063727, 
    4.250309,
  6.641526, 6.713795, 7.447269, 9.197515, 7.108441, 6.310119, 8.286802, 
    8.665269, 7.744537, 6.86899, 6.358835, 6.114986, 6.499959, 7.104738, 
    5.803327,
  7.390232, 7.638204, 8.787926, 9.758463, 9.904513, 7.081066, 6.503247, 
    6.878013, 6.988294, 6.407273, 6.207407, 6.298368, 6.600472, 7.253205, 
    6.423577,
  7.566547, 7.900764, 8.981761, 9.690468, 10.07508, 9.414853, 7.251514, 
    5.502158, 6.057775, 5.585142, 6.450126, 7.227382, 7.56303, 7.634594, 
    7.172334,
  8.03075, 8.751756, 9.186185, 9.325825, 9.599879, 9.797177, 9.161345, 
    8.380027, 7.241158, 6.247975, 5.580977, 8.179564, 8.405831, 7.589909, 
    7.31732,
  8.786489, 8.996142, 9.077247, 9.062965, 9.477909, 9.775964, 10.12078, 
    10.10261, 8.946314, 8.316951, 8.028964, 8.737837, 7.282291, 7.039179, 
    7.339139,
  9.298402, 9.189827, 9.211653, 9.375534, 9.874307, 10.49462, 10.64458, 
    10.43954, 9.500745, 9.395203, 9.28778, 6.760854, 6.883211, 7.296303, 
    6.280485,
  9.256129, 9.600507, 9.926404, 10.08833, 10.71813, 10.93428, 11.37983, 
    11.06881, 10.47432, 9.774623, 7.130588, 7.445878, 7.428695, 6.047299, 
    6.166179,
  9.41323, 9.954017, 10.62161, 11.30707, 11.88957, 12.16035, 11.99688, 
    11.35092, 9.232738, 5.009841, 6.455523, 8.129824, 5.938131, 5.422133, 
    5.836925,
  4.775323, 6.93188, 5.784063, 7.721228, 7.35574, 6.336759, 9.493462, 
    10.87782, 9.768135, 7.393202, 7.505285, 8.159516, 7.537706, 7.38461, 
    7.503653,
  7.463597, 8.093822, 7.576242, 7.893085, 5.269836, 6.109254, 9.791971, 
    10.70368, 11.53484, 10.08314, 8.549201, 9.645884, 9.991165, 7.840322, 
    8.096815,
  10.14068, 10.06385, 9.341694, 9.168849, 6.510934, 5.788563, 9.642544, 
    10.00339, 10.455, 10.72887, 10.95689, 11.75162, 12.52257, 12.37758, 
    10.06725,
  11.8344, 11.58417, 11.25619, 10.55121, 9.486598, 7.851147, 7.283763, 
    8.892419, 11.00501, 10.60543, 11.64806, 13.61481, 14.23229, 13.40781, 
    9.933846,
  13.06832, 12.51322, 11.87846, 11.35872, 11.24359, 11.01668, 9.330772, 
    7.611208, 9.430731, 9.815365, 13.60762, 15.49498, 15.35206, 13.23065, 
    10.83526,
  13.38029, 12.66196, 11.8567, 11.38459, 11.52344, 11.64766, 11.6597, 
    12.34801, 11.60343, 11.58106, 11.58005, 15.58658, 15.12705, 12.29594, 
    9.953204,
  11.89587, 11.64167, 11.44814, 11.16613, 11.74809, 11.85046, 12.57042, 
    13.56988, 14.7378, 15.13478, 14.98195, 15.51466, 13.27136, 9.871435, 
    7.589566,
  11.12915, 11.43394, 11.55765, 11.64102, 11.88998, 12.44739, 12.97803, 
    13.45803, 14.41286, 14.92225, 14.99733, 14.19674, 9.968064, 7.120341, 
    5.459701,
  12.20708, 12.29741, 12.2916, 11.6102, 12.15119, 12.53138, 13.27058, 
    13.70231, 13.79541, 13.71918, 13.71213, 11.4124, 6.650217, 5.860879, 
    5.192508,
  12.90528, 12.55723, 12.596, 12.44257, 12.40148, 13.10829, 13.57481, 
    13.03213, 10.97064, 8.915184, 9.265345, 6.991678, 6.199343, 5.365197, 
    3.649051,
  7.341906, 10.49476, 8.892182, 10.7143, 9.485789, 7.753011, 11.01424, 
    12.17919, 12.41286, 9.20507, 9.081838, 9.834546, 9.039924, 8.399747, 
    7.876414,
  11.5803, 12.76347, 11.49442, 10.86124, 7.038514, 7.086524, 11.20128, 
    11.89894, 12.74125, 11.23498, 9.684829, 11.342, 10.13175, 7.53705, 
    7.593989,
  13.80291, 14.64935, 14.25878, 12.70125, 9.43778, 7.10761, 10.64758, 
    11.15339, 11.38459, 11.58669, 11.17493, 11.03386, 10.27872, 10.15384, 
    8.816453,
  15.01682, 15.1584, 14.90321, 14.32632, 12.9609, 9.380743, 7.508859, 
    9.401525, 9.64398, 9.053165, 10.05169, 10.97336, 11.13041, 11.51748, 
    8.863223,
  16.13871, 15.70477, 15.05437, 14.34807, 13.63943, 12.41833, 10.36436, 
    7.117217, 7.273443, 6.803825, 9.723221, 11.35951, 11.4981, 11.50883, 
    9.572118,
  15.83627, 15.1221, 14.36612, 13.63805, 12.96855, 12.2749, 11.96371, 
    12.06271, 9.776066, 8.669621, 8.554097, 11.74091, 11.86138, 11.31951, 
    8.111616,
  13.47161, 13.12642, 12.77562, 12.09644, 11.88077, 11.5934, 11.74674, 
    11.66906, 11.95294, 12.04257, 11.83022, 11.90035, 11.53766, 9.93153, 
    6.706125,
  12.42001, 12.37835, 12.33983, 11.89201, 11.7882, 11.93957, 11.68039, 
    11.55552, 11.96778, 12.04927, 12.04346, 11.70715, 11.0304, 8.447457, 
    7.746727,
  14.54957, 14.30994, 14.06657, 13.26523, 13.27674, 12.50485, 12.85668, 
    12.76877, 12.4495, 11.8119, 11.46576, 11.30999, 10.28031, 8.607561, 
    7.818399,
  16.79136, 16.36722, 15.9435, 14.78991, 14.39614, 13.97718, 13.97504, 
    13.49794, 10.76876, 8.643887, 8.777, 10.73292, 9.424251, 9.478948, 
    7.419141,
  8.663574, 12.04714, 10.27772, 13.57296, 12.70426, 9.898085, 12.38502, 
    12.12765, 11.65235, 9.09772, 8.856795, 9.149226, 8.465245, 7.724981, 
    7.526527,
  13.36772, 15.10272, 13.40902, 13.55432, 9.14475, 8.511754, 14.54745, 
    13.89457, 13.42849, 11.86622, 9.889562, 11.17946, 11.40621, 8.055403, 
    7.696053,
  15.30925, 16.36048, 15.97681, 14.87396, 11.23856, 8.43725, 12.3991, 
    12.86554, 12.77742, 12.49117, 11.68031, 11.47792, 11.39529, 10.80559, 
    8.664862,
  16.09891, 16.8919, 16.94312, 16.76452, 15.97914, 11.20575, 8.086926, 
    9.448102, 11.38651, 11.47369, 11.76913, 10.89407, 9.756338, 9.643085, 
    8.04821,
  16.57775, 16.8897, 16.80466, 16.35005, 15.90426, 14.8998, 12.46563, 
    7.889956, 7.235853, 6.654891, 9.846677, 9.818428, 8.697864, 8.889918, 
    8.888384,
  15.55007, 15.7209, 15.7103, 15.46084, 14.92861, 14.31325, 14.06364, 
    14.02854, 9.967444, 7.365764, 6.999464, 9.316428, 9.016885, 9.440075, 
    9.953072,
  12.74086, 12.99337, 13.19962, 13.2697, 13.3265, 13.09557, 12.96424, 
    12.74356, 12.19037, 10.76665, 10.33911, 10.11157, 10.05489, 9.939396, 
    9.867867,
  11.22703, 11.63509, 12.03704, 11.97801, 12.08656, 12.39666, 12.2804, 
    11.95751, 11.73994, 10.68386, 10.49429, 10.18372, 9.915276, 9.686652, 
    9.763459,
  10.75965, 11.16269, 11.48836, 11.37791, 11.39563, 11.43497, 12.1767, 
    12.6884, 12.01979, 10.68419, 10.79193, 10.4448, 10.27741, 10.4497, 9.71771,
  8.830853, 9.364546, 9.805141, 9.711924, 9.617078, 9.724428, 9.806045, 
    9.849158, 9.303368, 8.324406, 8.720638, 11.07602, 10.57308, 10.11204, 
    9.336377,
  7.994765, 11.33155, 9.236082, 12.216, 10.30365, 9.083072, 11.70503, 
    10.99381, 10.43845, 8.678534, 8.428713, 8.997336, 7.769568, 6.69565, 
    6.534934,
  11.87981, 13.54423, 12.65143, 11.88999, 7.414193, 7.639849, 13.22342, 
    11.87672, 11.77137, 11.22798, 9.871661, 11.03488, 10.62575, 7.288893, 
    7.004771,
  11.77174, 13.78466, 14.20521, 14.10404, 9.339788, 7.26328, 11.76514, 
    12.89533, 12.93035, 11.83277, 12.70317, 12.93871, 12.01396, 11.23957, 
    8.552814,
  10.22183, 12.37981, 14.06613, 14.83362, 14.50087, 11.35233, 6.892925, 
    8.75951, 11.228, 12.62028, 13.0998, 13.08751, 12.74861, 11.78372, 9.522237,
  7.057811, 7.770425, 9.691849, 11.69031, 13.18303, 14.97981, 13.01854, 
    8.127806, 7.705493, 7.390484, 11.09801, 11.86355, 10.76197, 9.90717, 
    9.654879,
  5.371058, 4.406931, 4.479873, 5.108244, 6.29831, 8.344103, 11.40439, 
    14.15012, 9.928927, 7.251176, 7.202673, 10.34983, 9.927858, 9.45672, 
    9.342295,
  5.732053, 4.911368, 4.686472, 4.806464, 5.578444, 6.540004, 8.14242, 
    9.950212, 10.73959, 9.54291, 9.72089, 10.10792, 9.940026, 9.718131, 
    9.703918,
  7.359737, 6.670643, 6.33172, 6.441312, 7.07798, 7.532363, 7.475904, 
    7.445293, 8.244545, 7.511616, 8.578312, 9.09361, 9.357041, 9.342032, 
    9.458412,
  8.441084, 8.039426, 7.337409, 6.687409, 6.372502, 5.928829, 5.545047, 
    6.251218, 7.539355, 8.291124, 9.711678, 9.667569, 9.758489, 9.520528, 
    9.104902,
  8.716559, 8.611614, 8.130584, 7.246423, 6.252102, 5.309008, 5.548575, 
    6.036343, 5.791883, 5.529872, 6.149316, 6.439639, 5.332125, 4.580302, 
    4.15126,
  7.926132, 11.53982, 9.966699, 13.00688, 10.85432, 9.50803, 13.50087, 
    12.19413, 11.65613, 8.943577, 8.238787, 9.082815, 7.56053, 6.686445, 
    6.545029,
  11.24237, 13.75457, 13.79372, 13.2685, 7.578278, 8.302008, 14.07668, 
    13.83216, 12.79304, 11.82152, 10.32747, 12.24644, 11.45861, 7.775909, 
    7.078757,
  9.178668, 11.9137, 13.97236, 15.26425, 10.53859, 7.846483, 11.70148, 
    13.14493, 12.98818, 12.20791, 13.14618, 13.32776, 12.9176, 12.10754, 
    8.939709,
  5.808053, 5.919355, 7.481746, 10.12245, 13.36023, 11.47319, 6.728641, 
    7.882558, 10.74176, 11.69564, 12.52108, 13.53196, 12.91938, 12.69916, 
    10.16552,
  4.38201, 3.772671, 4.030073, 4.890412, 6.351172, 11.0052, 11.20362, 
    6.296522, 5.908024, 6.745683, 9.381012, 10.5516, 10.44345, 10.76547, 
    11.10524,
  5.376784, 4.224195, 4.186141, 4.550744, 5.127196, 4.239688, 7.920691, 
    10.55273, 6.844709, 4.256399, 4.911076, 7.425514, 7.977898, 8.701768, 
    9.520775,
  6.234181, 5.285413, 4.343836, 4.151442, 4.419007, 5.003121, 4.217373, 
    4.533627, 4.297369, 3.561443, 4.125385, 4.829304, 5.065878, 5.622617, 
    6.526359,
  6.441652, 6.279205, 5.43468, 4.740715, 4.378609, 4.152784, 3.762094, 
    3.165291, 3.050644, 2.826123, 3.706691, 4.03187, 4.732415, 5.65955, 
    6.566969,
  5.870571, 6.20538, 5.806958, 5.34035, 5.296319, 5.123976, 4.843025, 
    4.932444, 4.839251, 5.189277, 6.347566, 5.120063, 5.821865, 6.908258, 
    8.320672,
  5.207568, 6.121751, 6.142336, 5.774269, 6.035481, 5.858891, 5.007393, 
    4.475603, 4.112211, 3.846956, 4.389255, 4.655527, 4.474283, 4.76727, 
    4.938929,
  6.918136, 10.02486, 8.489274, 10.46282, 8.320137, 7.826704, 10.89137, 
    10.85588, 10.36577, 8.24132, 8.709214, 9.840137, 8.978568, 7.837048, 
    7.91839,
  9.420902, 11.70944, 11.84859, 11.28796, 5.980603, 7.051376, 11.33163, 
    11.58043, 11.36178, 10.61195, 10.16879, 12.48136, 12.52858, 8.361846, 
    7.828475,
  8.591183, 9.906183, 11.53893, 13.06239, 9.169972, 6.882656, 10.17841, 
    11.60633, 12.13202, 12.31451, 13.60725, 14.08297, 14.03851, 13.79228, 
    9.384964,
  7.20944, 6.440169, 7.06363, 8.467301, 10.91241, 10.08443, 6.052303, 
    7.076087, 9.593836, 11.15609, 13.43975, 14.8776, 14.85104, 14.81966, 
    11.53715,
  5.552757, 4.533463, 4.406484, 4.621559, 5.247386, 8.23674, 8.853203, 
    5.542877, 5.686531, 7.008614, 10.60432, 12.54752, 13.32349, 13.47293, 
    14.01616,
  5.423586, 4.495244, 3.780025, 3.327708, 3.072092, 3.68924, 5.687346, 
    7.786209, 5.112791, 3.789542, 4.962769, 7.979461, 8.929288, 10.38687, 
    11.57547,
  5.993237, 5.262032, 4.595596, 4.436851, 4.181571, 4.139256, 4.340569, 
    4.531144, 3.754132, 2.20206, 2.478877, 3.773983, 5.011126, 6.031296, 
    6.724302,
  7.311162, 6.944034, 6.441803, 6.6978, 6.535512, 6.187756, 5.519081, 
    5.111628, 4.492574, 3.371371, 2.671863, 2.171845, 2.753861, 3.437135, 
    3.941323,
  8.22169, 8.014817, 7.533977, 7.699752, 7.269883, 6.809836, 6.167861, 
    5.502224, 4.553516, 3.979915, 3.509241, 1.777504, 2.055371, 2.600999, 
    3.169652,
  7.498715, 7.726908, 7.603349, 7.616731, 7.374992, 6.818921, 6.285107, 
    5.620216, 4.645057, 3.784507, 3.213393, 2.069803, 1.398749, 1.498108, 
    2.529433,
  7.006031, 10.24924, 8.92412, 10.6759, 8.390185, 7.452877, 10.03468, 
    9.057471, 8.533552, 6.06228, 6.639796, 7.776071, 7.299487, 6.63395, 
    7.167916,
  8.599765, 10.83796, 11.8746, 11.75425, 7.188746, 7.377628, 11.05442, 
    10.25516, 9.519897, 8.169953, 7.944502, 9.642612, 9.908898, 6.699843, 
    6.726335,
  7.174895, 8.071877, 10.44559, 12.86479, 10.19774, 7.2323, 9.886349, 
    11.36304, 11.4353, 9.866199, 10.85051, 10.77131, 10.58875, 10.52299, 
    7.586085,
  5.685074, 5.449182, 6.810699, 7.525985, 12.59769, 11.36321, 6.451606, 
    7.359145, 10.54559, 11.43935, 12.39793, 12.35731, 11.10741, 10.8601, 
    9.411854,
  5.36727, 5.914389, 6.486267, 7.365334, 5.545304, 9.761511, 10.23814, 
    6.452518, 6.926855, 8.40978, 12.32577, 13.3127, 12.48339, 12.0299, 
    12.13444,
  5.815313, 6.314986, 6.371386, 7.371893, 8.684986, 5.869844, 5.039331, 
    7.547489, 4.800012, 4.187159, 6.836758, 10.80788, 11.50053, 11.60747, 
    11.66542,
  5.498315, 5.619778, 5.174541, 6.012064, 7.351456, 9.090627, 8.813745, 
    6.479463, 4.234925, 2.86841, 4.47894, 6.773468, 8.399676, 9.389131, 
    10.35398,
  5.129647, 4.214808, 3.386335, 3.812048, 4.490149, 5.295952, 6.003269, 
    6.812887, 7.254392, 6.086573, 3.239693, 3.023862, 3.908889, 5.226842, 
    6.7613,
  5.603343, 3.728987, 2.730119, 2.863148, 3.387181, 4.020356, 4.018888, 
    3.649492, 3.245123, 3.4232, 3.576055, 4.081785, 3.22915, 2.636678, 
    3.155168,
  7.543195, 4.846857, 3.586866, 3.015412, 3.34138, 3.792654, 3.775384, 
    3.142384, 2.389662, 2.369592, 2.086066, 2.319512, 2.630766, 2.456403, 
    1.586817,
  8.41614, 10.80358, 8.690897, 10.70745, 8.582168, 8.060695, 10.63265, 
    9.849052, 9.020896, 6.230458, 5.932719, 6.745738, 6.013844, 5.384382, 
    5.421659,
  11.83375, 11.98555, 10.66483, 10.31169, 5.951675, 6.819415, 10.69208, 
    10.23846, 9.967419, 8.705914, 7.479095, 8.752672, 9.060072, 5.988956, 
    5.845898,
  9.844406, 10.18568, 8.691715, 8.021039, 6.622321, 5.406794, 8.374403, 
    9.852211, 10.04634, 10.05829, 10.42241, 9.811371, 9.467305, 9.162641, 
    6.780938,
  7.469975, 7.414132, 5.446503, 4.41408, 6.518598, 6.361928, 3.9101, 
    5.447662, 7.600817, 10.10319, 11.34346, 10.35735, 9.428762, 9.027519, 
    8.072526,
  9.794755, 9.223598, 5.974895, 3.917845, 3.049935, 4.775267, 5.233277, 
    2.796766, 3.279208, 4.666019, 9.556993, 10.95734, 10.32213, 9.898237, 
    10.19241,
  12.7021, 10.83592, 6.41649, 3.56427, 4.307945, 4.240978, 4.104814, 
    4.587831, 2.967997, 2.904171, 3.627338, 8.060287, 9.790917, 9.790559, 
    9.722826,
  13.3927, 10.52332, 6.167932, 3.077475, 3.339198, 5.597589, 7.288008, 
    7.506471, 6.197301, 5.369491, 4.679679, 5.912416, 8.200921, 9.704959, 
    10.02542,
  12.27549, 8.695733, 4.086173, 3.881066, 4.249318, 4.940921, 5.581526, 
    4.85133, 3.718749, 4.019516, 5.135986, 4.595884, 7.069961, 9.211696, 
    9.72423,
  12.50381, 9.821888, 6.987216, 5.634136, 5.221043, 4.514585, 3.853451, 
    3.077951, 2.219937, 2.780174, 4.969094, 5.995456, 4.413427, 8.127573, 
    8.975019,
  12.84492, 10.72856, 9.350798, 9.352737, 9.376216, 7.334558, 4.821069, 
    2.275774, 1.162336, 1.914391, 3.737747, 6.225011, 5.198403, 6.068448, 
    8.340454,
  6.125191, 9.243629, 8.252221, 11.70309, 10.94531, 9.284458, 11.30307, 
    9.332506, 8.878311, 6.189525, 5.718972, 5.890442, 4.620955, 3.926888, 
    3.609342,
  7.246834, 9.011479, 9.038326, 9.213657, 6.68137, 7.551662, 11.02849, 
    9.94908, 9.673506, 8.639371, 7.167788, 8.121687, 7.966005, 4.727671, 
    3.957521,
  7.166672, 8.826312, 9.248557, 8.594337, 7.045533, 5.294721, 8.566237, 
    10.35103, 9.817625, 9.387334, 9.841292, 9.484324, 9.449425, 8.373607, 
    5.882167,
  6.964635, 8.170289, 8.991039, 9.472919, 9.911841, 6.781621, 3.855163, 
    6.031063, 8.344953, 9.974833, 10.42072, 9.466505, 9.357623, 8.972085, 
    7.489356,
  8.141449, 10.11059, 9.946653, 8.874425, 8.092104, 8.625385, 6.893522, 
    4.600459, 5.010869, 6.192439, 9.594114, 10.02908, 9.61557, 9.972809, 
    10.30792,
  13.22034, 12.38782, 10.53089, 7.983847, 5.072946, 4.506749, 7.306881, 
    8.870315, 5.666564, 4.595253, 4.915902, 7.18577, 8.422196, 9.164972, 
    9.427046,
  14.44245, 12.97699, 10.90955, 7.711246, 5.030205, 4.227388, 5.558386, 
    8.249209, 8.104679, 7.411481, 6.39844, 5.622386, 4.73445, 5.523359, 
    7.178075,
  16.02467, 14.24608, 12.24198, 9.918852, 8.876146, 8.263943, 9.308054, 
    10.6902, 11.06146, 8.681739, 6.119808, 4.961356, 4.808645, 3.97346, 
    4.012646,
  17.06454, 14.88157, 12.39638, 10.42016, 10.15723, 10.98689, 8.268681, 
    9.526078, 10.92635, 9.097545, 6.631729, 4.949448, 4.548931, 4.146641, 
    3.383058,
  14.16861, 12.2336, 10.50686, 9.414855, 9.323755, 10.88393, 12.68971, 
    10.5422, 7.20204, 5.372768, 4.736567, 4.993361, 4.938401, 5.009414, 
    4.318545,
  3.124835, 5.009633, 4.898648, 7.813118, 7.784956, 7.741634, 10.64822, 
    10.55241, 9.869846, 6.63827, 5.496022, 5.530376, 4.231553, 3.363661, 
    3.831719,
  5.025331, 5.033085, 5.486198, 6.386228, 4.804728, 5.853378, 9.461428, 
    10.21963, 9.996264, 8.430034, 6.392724, 7.042452, 6.088778, 3.260238, 
    3.052416,
  4.813605, 6.057136, 6.422193, 6.740529, 5.750445, 4.71711, 6.918292, 
    9.221786, 10.26856, 9.966555, 8.945482, 7.957417, 6.432559, 4.842874, 
    3.058125,
  2.797315, 3.197209, 5.588875, 6.784421, 7.549508, 5.575066, 4.515642, 
    6.010225, 7.913672, 9.253654, 8.977026, 7.966863, 6.327118, 4.78518, 
    3.374217,
  7.769537, 8.899569, 8.053387, 7.200591, 6.205252, 6.505454, 6.365842, 
    4.847955, 4.623837, 6.045368, 8.609871, 8.072249, 6.8497, 5.654285, 
    4.121358,
  12.03768, 11.42532, 10.4558, 9.442932, 7.987475, 6.135656, 5.809166, 
    7.230727, 5.724924, 5.675894, 6.360046, 8.340475, 7.634799, 6.382027, 
    4.73167,
  12.55409, 12.36794, 11.85874, 11.44026, 10.2458, 8.708429, 5.94775, 
    3.723347, 4.812312, 8.586658, 9.432415, 8.867268, 8.133629, 7.241541, 
    5.867773,
  11.67158, 11.83834, 11.46947, 11.27478, 10.24597, 9.137996, 7.955299, 
    6.611323, 5.03154, 4.366658, 8.784206, 9.48259, 8.623542, 7.779967, 
    6.674906,
  9.733024, 9.656174, 9.369434, 8.991346, 8.308368, 7.599203, 7.092296, 
    7.095933, 6.162048, 4.862097, 6.524266, 9.261983, 9.127145, 8.250257, 
    6.830996,
  8.152355, 8.019052, 7.686921, 7.025869, 6.57982, 6.621836, 6.862376, 
    7.10763, 5.544075, 4.115241, 5.56547, 8.929018, 9.186124, 8.688392, 
    7.290181,
  2.753623, 4.602363, 4.707425, 6.618659, 6.404032, 6.146551, 8.755889, 
    9.30365, 9.039429, 7.101398, 7.444187, 8.775519, 8.383475, 7.413267, 
    6.672776,
  5.650109, 5.839239, 5.35974, 5.871241, 4.426733, 5.567955, 8.492505, 
    9.071499, 9.358581, 8.968619, 8.363191, 11.2477, 11.69753, 7.323828, 
    6.242078,
  4.472658, 6.661644, 7.321323, 6.839839, 5.119354, 4.179793, 6.858679, 
    8.964841, 10.07041, 10.51914, 11.10788, 11.53487, 12.07874, 10.65066, 
    7.459824,
  4.635715, 2.532458, 4.270802, 7.841187, 8.543081, 6.021083, 3.702208, 
    5.264395, 7.999933, 10.33012, 10.8878, 11.0138, 10.71832, 9.896152, 
    7.924004,
  10.99875, 10.39365, 7.345465, 3.280034, 7.125709, 9.000741, 6.899289, 
    4.96115, 5.274234, 6.496629, 10.33381, 10.69294, 10.3261, 9.868205, 
    8.779789,
  10.57602, 12.00061, 13.00896, 10.99362, 7.014787, 5.735965, 7.522892, 
    8.452374, 6.216481, 6.34679, 7.740251, 10.88361, 10.40728, 9.399941, 
    7.919319,
  8.648606, 9.614352, 11.3322, 13.12145, 13.61526, 11.7295, 7.367898, 
    5.819263, 7.141265, 9.441898, 10.95653, 10.96432, 10.71584, 9.558194, 
    7.911439,
  7.068779, 7.412221, 8.355783, 9.797224, 10.9417, 11.72305, 11.42307, 
    8.661677, 5.743363, 7.245043, 9.919738, 10.93092, 10.76229, 9.727194, 
    8.39765,
  6.652332, 6.876401, 7.609805, 8.378008, 8.794291, 9.041407, 9.422804, 
    9.648304, 7.433936, 5.504736, 7.951591, 10.55326, 10.59713, 10.0869, 
    8.310847,
  7.75372, 6.885871, 7.012293, 6.712972, 6.667916, 6.967369, 7.215663, 
    7.315251, 6.380817, 4.308013, 4.88621, 9.197021, 10.2743, 10.02819, 
    8.386638,
  2.046262, 1.935232, 1.613695, 3.056677, 3.338199, 3.163897, 4.314057, 
    4.875574, 7.818687, 7.356246, 8.074167, 10.23819, 10.01199, 8.804729, 
    7.703516,
  4.282676, 3.258535, 1.770269, 2.706413, 2.791684, 3.918282, 5.411696, 
    5.596682, 7.418353, 9.244013, 9.171255, 12.52084, 13.10673, 8.613863, 
    7.875501,
  7.646522, 3.830935, 4.847346, 2.840457, 3.038169, 2.989741, 5.536727, 
    6.610081, 8.537676, 10.18043, 11.47501, 12.3732, 12.81522, 12.27248, 
    9.928728,
  11.8749, 6.825361, 4.051771, 5.97823, 4.620021, 3.815391, 3.526927, 
    6.241296, 7.881002, 8.401297, 10.56906, 11.84482, 12.52564, 12.33458, 
    10.61964,
  11.08436, 12.65411, 6.666608, 4.689046, 7.280972, 6.150502, 5.568507, 
    4.586266, 4.657198, 5.662213, 9.924659, 11.79759, 12.46183, 12.19841, 
    11.53347,
  8.090278, 10.99609, 13.06784, 7.078585, 6.113657, 7.887335, 7.460114, 
    7.767378, 6.291453, 6.558193, 7.841592, 11.73588, 11.8552, 10.84852, 
    9.819549,
  7.038412, 8.538788, 11.79374, 12.42898, 7.934934, 7.156164, 6.625026, 
    7.80589, 8.59823, 9.724263, 10.86956, 11.44114, 11.06097, 10.7276, 
    10.06377,
  6.896848, 7.439422, 9.395768, 11.38433, 11.3498, 9.577136, 7.829947, 
    6.238678, 8.683788, 9.641728, 10.06818, 10.94841, 10.82444, 10.40881, 
    10.39563,
  8.52721, 8.200041, 8.565865, 9.670375, 10.73642, 10.75487, 9.150397, 
    6.755408, 5.059507, 8.405321, 9.490151, 10.35012, 10.46752, 10.50189, 
    10.05719,
  8.7249, 8.350951, 7.923244, 7.958899, 8.314026, 8.899194, 8.5003, 6.707024, 
    3.821482, 4.889319, 7.062862, 9.966773, 10.30786, 10.98728, 9.787642,
  5.430339, 5.667033, 4.542571, 7.455359, 8.110503, 6.896481, 8.629191, 
    8.36188, 9.251388, 7.115257, 7.088131, 7.473067, 6.406602, 5.470098, 
    4.811154,
  9.856898, 6.175679, 5.517942, 6.449395, 3.94778, 2.767044, 3.457728, 
    5.488703, 7.862203, 8.920415, 7.804753, 9.848071, 9.761844, 5.435277, 
    4.703709,
  12.45741, 9.679731, 5.795285, 4.438346, 3.61749, 2.505532, 4.071552, 
    5.647927, 8.127137, 9.537881, 9.818081, 9.323881, 9.25399, 8.608319, 
    6.504304,
  12.37016, 12.24374, 8.801517, 6.293118, 5.143125, 4.10913, 3.680037, 
    6.028337, 7.182637, 7.301754, 8.490506, 8.574835, 8.345718, 8.716149, 
    8.104975,
  11.63299, 12.68005, 10.79872, 7.838345, 6.8672, 5.863629, 6.193138, 
    4.937071, 4.588082, 4.679272, 7.535711, 8.447741, 8.777122, 9.406423, 
    9.57737,
  11.20863, 12.88227, 12.47861, 9.645444, 7.680282, 7.108093, 6.196747, 
    6.940438, 6.301047, 6.587919, 6.618929, 9.059555, 9.202303, 8.843834, 
    8.848527,
  10.79904, 12.84641, 13.59628, 12.03315, 9.313472, 8.464104, 8.011597, 
    7.664349, 8.183096, 9.599447, 10.15356, 10.34337, 10.14636, 9.979152, 
    10.61456,
  10.80433, 12.59138, 13.70135, 13.69187, 11.73235, 9.803362, 9.106781, 
    9.261095, 9.379016, 10.04533, 11.11642, 11.66286, 12.38678, 12.40338, 
    12.24391,
  11.14369, 12.60471, 13.4639, 13.7451, 12.86369, 11.08553, 9.937767, 
    9.930904, 9.993778, 10.71029, 11.98598, 13.21297, 13.67093, 13.13074, 
    11.51605,
  10.14607, 11.4706, 12.65016, 13.16134, 12.69377, 11.14238, 9.868936, 
    9.947495, 8.917809, 7.649108, 9.693225, 13.34825, 12.85854, 11.90249, 
    10.71062,
  6.77118, 8.041276, 4.689914, 4.09279, 3.188748, 7.384395, 13.46854, 
    13.25512, 10.82323, 7.021139, 6.722671, 7.392819, 6.624201, 5.689495, 
    4.561367,
  9.561997, 6.718038, 4.978483, 3.685384, 3.35315, 3.554666, 12.64255, 
    14.31952, 11.56209, 9.654725, 7.758338, 9.265641, 9.194431, 5.245401, 
    4.289484,
  10.04604, 7.026825, 4.486609, 3.586159, 3.867593, 4.477468, 9.262283, 
    12.81619, 12.09043, 10.83935, 9.634307, 8.952485, 8.548989, 7.612966, 
    5.714382,
  11.34038, 9.239757, 7.797303, 7.311958, 7.524203, 8.509294, 8.458971, 
    8.766582, 9.364092, 8.561193, 8.471504, 7.755666, 7.182194, 7.241573, 
    6.561892,
  12.33867, 11.02152, 9.923008, 9.833643, 10.49343, 11.80503, 11.5408, 
    8.143855, 5.633473, 4.813231, 7.280922, 7.265155, 6.921313, 6.862079, 
    7.015183,
  12.97737, 12.08481, 11.15347, 10.75266, 11.38174, 11.68812, 11.29314, 
    10.84297, 7.778862, 6.779126, 5.705063, 7.019043, 6.347729, 5.661335, 
    5.187773,
  13.47257, 12.81489, 11.98616, 11.28646, 11.37773, 11.73614, 11.19413, 
    10.08091, 9.282883, 8.983205, 7.73091, 6.550955, 5.533137, 4.390108, 
    4.041677,
  13.83633, 13.21997, 12.52316, 11.90211, 11.18851, 11.10629, 10.8977, 
    10.35418, 8.54961, 7.37377, 6.427352, 5.198428, 4.571035, 4.881497, 
    5.403453,
  13.54289, 13.15103, 12.49966, 11.81767, 10.67932, 10.10196, 9.614981, 
    8.764876, 7.317331, 5.890547, 5.177976, 5.446314, 5.999284, 6.347046, 
    6.019304,
  11.96201, 12.04261, 11.62898, 10.86778, 9.302081, 8.139674, 7.63348, 
    7.644833, 5.674323, 4.182939, 4.702157, 7.015374, 7.577833, 7.385654, 
    7.097704,
  3.324945, 4.661197, 3.58685, 5.18865, 5.990315, 5.035372, 5.03194, 
    4.519783, 4.076797, 2.620807, 2.850103, 4.580425, 5.266807, 5.14102, 
    4.120699,
  7.026899, 6.076353, 5.938957, 5.74843, 4.487033, 4.424012, 6.437444, 
    6.399878, 4.109198, 2.204661, 3.192816, 6.166247, 8.40239, 5.561035, 
    4.333514,
  11.41306, 9.694257, 8.736979, 8.14789, 7.970681, 6.687906, 7.927919, 
    7.867574, 6.589664, 5.802066, 5.810363, 6.641816, 9.637486, 10.01274, 
    6.652562,
  13.13645, 12.72431, 12.16792, 11.52611, 10.92968, 8.586721, 5.288869, 
    6.085059, 8.407784, 8.042767, 7.856328, 7.027654, 8.487322, 10.39392, 
    8.891323,
  11.7069, 12.0062, 11.93356, 11.63192, 10.23944, 8.624166, 7.152623, 
    4.152034, 4.251839, 5.1143, 7.682769, 7.358636, 7.846739, 10.61115, 
    10.73487,
  9.691937, 10.05785, 9.944374, 9.652772, 8.980604, 7.60631, 6.143782, 
    6.27997, 4.688306, 5.323975, 6.055204, 8.206379, 8.162006, 9.787657, 
    9.704897,
  7.962752, 8.15694, 8.041018, 7.807797, 7.718844, 7.713162, 7.011883, 
    6.384545, 6.125504, 7.03317, 7.964237, 8.467962, 8.961399, 9.321864, 
    9.22926,
  6.995246, 7.499608, 7.568061, 7.48751, 7.097023, 6.901573, 6.684433, 6.398, 
    5.729642, 5.762889, 6.294121, 6.923497, 7.442172, 7.677914, 7.426886,
  6.287759, 6.948289, 7.221578, 7.057464, 6.215367, 5.660274, 5.265417, 
    4.775769, 4.002716, 3.66809, 3.942865, 4.523659, 5.186311, 5.70668, 
    5.859753,
  4.817498, 5.224532, 5.583289, 5.383502, 4.875451, 4.341858, 3.76087, 
    3.270866, 2.782217, 2.370946, 2.857739, 3.754956, 4.181449, 4.42557, 
    4.514952,
  4.063093, 5.52918, 4.693204, 5.078868, 4.189802, 3.678061, 5.187124, 
    6.854042, 8.103045, 7.128722, 8.002794, 8.378294, 6.507639, 5.818626, 
    5.292125,
  7.161475, 6.141449, 5.543669, 4.788356, 3.650604, 3.988451, 6.079613, 
    7.067529, 8.247313, 8.584629, 8.108314, 9.598722, 9.12369, 5.460778, 
    4.511392,
  7.537874, 6.420023, 5.83829, 4.819464, 4.400695, 3.357798, 5.48945, 
    6.406963, 7.128817, 8.267559, 8.664932, 8.606221, 8.415209, 6.841357, 
    5.414375,
  7.897155, 7.481236, 7.170998, 6.38531, 5.255733, 4.160327, 2.365238, 
    4.944489, 7.7049, 8.288102, 7.98448, 7.353884, 7.114559, 6.755639, 
    5.396346,
  6.875486, 7.004159, 6.859826, 6.579339, 5.502967, 4.75954, 3.963162, 
    2.762068, 4.313725, 5.297597, 6.946974, 5.945016, 6.013834, 6.624986, 
    5.732248,
  4.375096, 4.703048, 4.668834, 4.614788, 4.616342, 4.920135, 4.862081, 
    5.068837, 4.561892, 5.628444, 5.092865, 4.996941, 4.522886, 6.608604, 
    6.041259,
  2.626914, 2.845414, 2.645634, 2.826238, 3.610639, 4.508487, 4.787837, 
    5.644962, 6.885816, 8.350297, 8.11008, 5.790379, 3.842766, 6.278813, 
    5.934032,
  2.382569, 2.704163, 2.648276, 3.024342, 3.538852, 3.593828, 3.527346, 
    4.001101, 4.871687, 6.847753, 8.030437, 7.251878, 5.104017, 6.214923, 
    5.94204,
  3.327787, 3.900385, 3.509055, 3.362324, 2.780252, 2.523487, 2.344489, 
    2.109015, 2.794287, 4.931823, 6.683977, 7.181183, 5.573553, 5.528216, 
    5.648085,
  3.187274, 3.011022, 2.686061, 1.943461, 1.677308, 1.73945, 2.296683, 
    1.886146, 0.9870979, 2.128285, 3.721301, 5.710023, 5.171721, 4.274569, 
    4.519774,
  2.463506, 4.039179, 4.305976, 6.034028, 5.914042, 5.308556, 7.993198, 
    9.083668, 9.617331, 7.452503, 6.78626, 8.113035, 10.18038, 8.804582, 
    6.976809,
  3.24172, 3.34972, 4.434185, 5.026849, 4.302467, 4.804021, 8.654188, 
    10.08146, 11.39578, 10.60198, 6.739723, 9.48319, 13.82394, 8.872798, 
    6.718905,
  3.476893, 2.771883, 3.080269, 3.622725, 4.21594, 3.969602, 7.70493, 
    9.124776, 10.95845, 11.85746, 8.721631, 9.981004, 14.23397, 13.30076, 
    9.010524,
  4.184581, 3.108205, 2.780439, 3.832949, 5.197693, 5.714309, 4.659194, 
    8.033169, 14.56778, 14.36623, 10.72937, 10.48071, 12.83917, 12.7441, 
    10.75559,
  5.206693, 4.147093, 3.005223, 2.991695, 4.246911, 6.793689, 7.165829, 
    5.642301, 7.977856, 9.081412, 10.48469, 10.88466, 11.97862, 11.92139, 
    12.12517,
  7.617042, 6.904759, 5.647019, 3.840427, 2.639913, 4.71749, 7.562216, 
    8.480468, 6.816887, 7.580768, 7.803361, 10.97612, 10.40281, 9.744331, 
    9.718484,
  8.141341, 7.896224, 7.53949, 6.165953, 3.627471, 2.359604, 5.713424, 
    8.564301, 10.56435, 11.48607, 10.80645, 10.59728, 9.847662, 9.073619, 
    8.565985,
  6.696235, 5.69837, 5.267569, 4.476182, 4.121151, 3.542518, 3.926772, 
    5.899568, 8.090914, 9.884747, 10.1409, 9.662423, 8.986651, 8.236636, 
    7.326674,
  6.468043, 4.681486, 4.142505, 4.538822, 4.835237, 5.192509, 4.413657, 
    4.073026, 5.843755, 8.023082, 8.604777, 8.165546, 7.508235, 6.990059, 
    6.544864,
  8.141651, 5.882261, 5.838133, 5.25644, 5.194846, 5.281798, 5.287919, 
    4.679672, 3.588427, 4.144383, 5.266311, 6.90426, 5.968462, 5.412266, 
    5.368721,
  6.007084, 7.539449, 6.245363, 7.886899, 7.61016, 6.348398, 8.824435, 
    7.864081, 6.327886, 5.150867, 5.163828, 4.594299, 3.951895, 3.942212, 
    3.548551,
  9.836522, 9.147225, 8.603543, 8.969646, 6.423924, 5.879911, 8.444431, 
    7.477467, 6.020135, 6.612463, 6.695105, 7.477695, 7.510789, 4.311496, 
    3.716669,
  9.514306, 9.267067, 8.908349, 9.354999, 7.808288, 6.037019, 6.428018, 
    4.729482, 4.940657, 6.86012, 8.843998, 9.203848, 8.835074, 7.759616, 
    6.027698,
  8.476702, 7.734901, 8.052903, 9.229112, 7.756389, 3.596658, 2.522702, 
    4.254344, 4.953768, 5.486028, 8.88323, 10.29218, 9.581718, 8.247446, 
    7.32965,
  7.467896, 5.677696, 6.920628, 7.651481, 5.602736, 4.270687, 3.864279, 
    2.651498, 3.256828, 3.991648, 8.561984, 10.56033, 10.34031, 8.959089, 
    8.188246,
  7.194434, 5.345214, 7.491236, 8.088925, 5.814638, 5.156504, 4.932249, 
    4.543606, 4.516096, 6.551526, 7.872529, 10.94283, 9.422538, 9.120632, 
    8.095545,
  8.056532, 6.880251, 8.32515, 8.160312, 7.95522, 7.453392, 7.720872, 
    7.94453, 8.7523, 10.83594, 11.43651, 10.88295, 9.436029, 9.563075, 
    8.741739,
  8.704347, 7.604408, 8.50326, 9.76717, 10.44617, 9.912295, 10.15338, 
    10.66499, 10.96731, 11.31661, 11.26324, 10.02467, 9.828753, 9.300145, 
    8.25456,
  9.24428, 8.65496, 10.38088, 12.05016, 11.41801, 10.84824, 10.93837, 
    11.28222, 11.19732, 10.51444, 10.17968, 9.586059, 9.380065, 8.51025, 
    7.093587,
  10.53145, 11.13988, 12.51499, 11.55982, 10.67438, 10.11968, 10.19351, 
    10.52472, 8.25924, 6.292176, 6.348064, 8.100892, 7.39935, 6.330917, 
    5.183959,
  7.650518, 12.20802, 10.84851, 12.98872, 10.74376, 8.124389, 9.968848, 
    9.711125, 9.36817, 6.506998, 6.001859, 6.072195, 4.799609, 4.308477, 
    4.419899,
  5.705524, 8.620122, 10.85404, 12.02848, 7.70952, 6.261999, 9.568454, 
    9.736969, 9.76605, 8.423285, 6.428238, 6.077674, 5.232408, 3.25658, 
    3.141626,
  4.02464, 5.500645, 8.242646, 10.9309, 8.7826, 5.946659, 7.710866, 7.580417, 
    6.450057, 6.838816, 5.931027, 3.28228, 2.887136, 3.976663, 3.600745,
  4.115305, 5.553671, 8.411047, 10.7197, 9.488341, 6.088063, 3.268903, 
    2.810126, 4.11876, 4.847726, 4.54446, 1.981103, 2.106177, 2.800617, 
    3.520234,
  3.516226, 4.370674, 6.028726, 7.415572, 8.021212, 6.022747, 5.286959, 
    4.503026, 3.720922, 3.3567, 3.653085, 2.686882, 2.767017, 2.638469, 
    2.648893,
  7.520443, 7.403225, 7.891272, 8.413143, 7.240082, 5.319914, 5.714954, 
    8.120917, 6.589386, 5.05024, 3.924739, 4.66406, 4.780559, 4.721537, 
    4.349187,
  10.672, 10.43814, 10.10994, 9.653752, 9.072618, 9.51789, 10.21122, 
    9.873931, 8.884652, 7.566541, 6.963684, 6.608361, 6.361864, 5.957064, 
    5.615534,
  12.7837, 13.02895, 12.98156, 12.74645, 12.50359, 12.87629, 12.78964, 
    11.64539, 9.887609, 8.456223, 7.731195, 7.112883, 6.395843, 5.687741, 
    5.005826,
  14.82227, 15.19453, 15.09516, 14.7492, 14.1454, 13.46896, 12.38451, 
    11.0602, 9.130594, 7.959527, 7.293401, 6.979262, 6.418846, 5.809186, 
    5.130359,
  14.85753, 15.07567, 14.81936, 13.98446, 12.83553, 11.38444, 10.03172, 
    9.400653, 6.914542, 5.060616, 5.086132, 6.278331, 5.995584, 5.578815, 
    5.193089,
  3.288126, 6.546033, 8.691699, 12.96469, 11.14573, 8.101997, 9.154812, 
    7.670301, 6.414485, 4.273284, 3.828339, 4.623392, 4.414782, 4.340955, 
    4.970497,
  4.014085, 5.273526, 8.49763, 11.69076, 8.341431, 6.74712, 9.013269, 
    7.882494, 6.320963, 5.35135, 4.537971, 5.993142, 7.07395, 5.076458, 
    5.095068,
  3.47171, 4.107701, 6.975731, 10.46323, 9.305791, 6.351601, 6.437128, 
    6.723073, 5.901901, 5.88487, 6.330989, 6.728478, 7.331079, 7.882483, 
    5.995027,
  3.45053, 4.853343, 7.726731, 10.66658, 12.05624, 8.745826, 5.235968, 
    3.32319, 2.48374, 4.206813, 4.887958, 5.248831, 5.455517, 5.757924, 
    4.958866,
  7.059029, 7.795032, 9.606691, 11.13224, 10.62507, 9.426773, 8.317603, 
    4.153512, 2.935398, 3.154444, 2.616132, 3.289755, 3.827099, 4.056417, 
    3.98061,
  10.50705, 11.01562, 11.40469, 11.42217, 10.22717, 8.006063, 6.468365, 
    5.663372, 3.071362, 1.327618, 1.057067, 2.298086, 3.025126, 3.006505, 
    2.774384,
  11.36248, 11.76425, 11.34451, 10.73006, 9.858697, 8.879578, 6.894938, 
    4.922043, 3.901877, 2.939642, 1.889001, 2.383472, 2.356346, 2.153875, 
    1.807775,
  11.35931, 11.60947, 11.16093, 10.70754, 10.15585, 9.588464, 8.375355, 
    6.75699, 4.86021, 3.644274, 3.114264, 2.963476, 2.654941, 2.233335, 
    1.926197,
  12.44788, 12.50515, 11.86807, 11.06083, 9.929377, 8.755733, 7.055882, 
    5.275887, 3.87925, 3.452933, 3.775861, 3.905756, 3.617913, 3.20663, 
    2.852906,
  12.33415, 11.96827, 10.97019, 9.362766, 7.555505, 6.088203, 4.571867, 
    3.823238, 2.671819, 2.191586, 2.804679, 3.811215, 3.859599, 3.589478, 
    3.266977,
  3.724024, 4.734351, 4.015353, 5.823142, 6.277359, 6.386002, 8.985866, 
    9.473833, 8.178412, 4.811536, 3.302145, 3.265589, 3.067654, 2.941719, 
    2.959477,
  4.866862, 3.690666, 3.547935, 5.72679, 6.00079, 6.168383, 8.71302, 
    8.874709, 6.822147, 5.12965, 3.443239, 3.666867, 4.048068, 3.403849, 
    3.430607,
  5.067159, 4.677657, 4.762616, 7.71773, 8.215933, 6.940046, 6.962729, 
    6.639726, 5.654957, 4.581093, 3.797457, 4.131487, 5.193696, 6.152781, 
    4.613594,
  5.205319, 5.764443, 6.659311, 9.239985, 10.63865, 8.770657, 6.229157, 
    4.052139, 1.593624, 3.160047, 4.18325, 4.917655, 5.46232, 5.457083, 
    4.037433,
  6.616492, 7.204059, 8.434149, 10.26839, 9.8043, 9.172959, 8.169889, 
    4.353103, 2.567197, 3.528427, 2.850871, 3.324821, 3.495812, 3.558246, 
    3.249512,
  8.359628, 8.81375, 9.584289, 10.28391, 9.24628, 7.282617, 6.350183, 
    5.271881, 2.200549, 1.147725, 1.069049, 1.486019, 2.47833, 2.662822, 
    2.62312,
  9.665668, 9.867461, 9.66452, 9.390837, 8.324152, 7.171093, 5.317752, 
    3.463836, 3.451741, 3.223553, 1.940684, 1.989976, 2.09551, 1.985329, 
    1.901598,
  9.620554, 9.291242, 8.393673, 7.871654, 7.212345, 6.71454, 6.177634, 
    5.275591, 3.874201, 2.359642, 2.098184, 2.317351, 2.436782, 2.38147, 
    2.225358,
  9.927986, 9.336452, 8.251928, 7.307794, 6.194212, 5.596499, 5.102601, 
    4.155066, 2.905432, 2.09942, 2.334165, 2.765225, 2.905003, 2.94988, 
    2.899883,
  9.523639, 9.156234, 8.116011, 6.389078, 4.79739, 3.976336, 3.896054, 
    3.626161, 2.555354, 1.258042, 1.307616, 2.460298, 2.988733, 3.032491, 
    3.160733,
  2.377323, 3.324789, 2.654313, 3.131397, 2.223197, 1.82025, 2.785603, 
    3.263569, 4.856977, 5.3222, 5.662945, 6.191155, 5.558879, 4.313589, 
    3.390664,
  2.62938, 1.854817, 1.552319, 2.230764, 2.716184, 3.349885, 4.80113, 
    6.607621, 8.447064, 8.615907, 7.149622, 7.108994, 5.779792, 3.350193, 
    2.985818,
  2.996348, 2.766411, 2.96158, 4.008781, 4.733012, 3.966421, 6.738122, 
    8.900436, 9.816621, 9.100948, 7.113141, 4.888041, 3.293997, 2.91595, 
    2.999497,
  4.003637, 4.239846, 4.845367, 5.714641, 5.99264, 6.030674, 4.950457, 
    6.886593, 7.883101, 5.659951, 4.418493, 2.969966, 2.43499, 2.710471, 
    2.434892,
  5.81096, 6.081522, 6.698955, 7.640128, 6.703606, 6.810206, 7.164852, 
    4.437575, 3.374688, 2.322455, 2.575337, 2.082636, 2.235031, 2.731896, 
    3.529291,
  6.241228, 7.116601, 7.836869, 8.427878, 7.748, 6.218494, 5.089957, 5.34856, 
    3.768525, 2.807863, 2.985573, 2.903576, 3.118748, 3.410064, 4.320805,
  5.909877, 7.047361, 7.480958, 7.760295, 7.615301, 7.461253, 6.36391, 
    5.425925, 5.056397, 4.666674, 3.865915, 3.336189, 3.434301, 3.850242, 
    4.667091,
  5.318964, 6.298123, 6.468415, 6.699001, 7.04322, 7.506001, 7.430766, 
    6.835417, 5.702538, 4.784174, 3.952062, 3.650365, 3.696484, 4.210918, 
    4.743052,
  5.410142, 6.238715, 6.421603, 6.788876, 7.336728, 7.572669, 6.98873, 
    6.082913, 5.257689, 4.600412, 4.20757, 4.158679, 4.251076, 4.565887, 
    4.856019,
  7.004964, 7.543252, 8.011435, 7.608167, 7.39236, 7.191501, 6.568009, 
    5.70717, 4.371089, 3.368517, 3.614686, 4.571617, 4.71652, 4.90143, 
    5.139664,
  2.604736, 3.164532, 3.268926, 4.120303, 4.311902, 4.584155, 5.613937, 
    5.031392, 4.258307, 3.406353, 3.573194, 4.104302, 4.016783, 3.847035, 
    3.079958,
  4.436202, 3.7448, 4.447227, 4.082877, 3.661724, 5.2749, 8.205246, 8.212709, 
    8.189522, 7.209296, 5.461368, 5.571701, 4.926123, 2.940957, 1.98823,
  5.176639, 4.188649, 4.581109, 3.734842, 3.667003, 3.582677, 6.496487, 
    7.911553, 8.261163, 7.789128, 6.71627, 5.600736, 4.683542, 2.593828, 
    1.370219,
  5.750343, 4.974338, 5.054529, 4.472768, 3.731646, 3.306556, 2.502589, 
    5.915532, 9.465473, 8.164799, 6.941185, 6.267991, 6.269579, 5.433208, 
    3.820894,
  6.077724, 5.451712, 5.398916, 5.185925, 4.06176, 3.964228, 3.441005, 
    3.197201, 4.09271, 4.730156, 6.133584, 6.468391, 7.068055, 7.208547, 
    6.926483,
  6.741251, 6.081148, 5.789247, 5.137516, 4.725662, 5.177565, 5.302907, 
    4.810399, 3.065775, 3.811877, 4.384554, 6.292449, 6.833614, 6.965579, 
    7.518078,
  7.546416, 7.170853, 6.315218, 5.352635, 5.377681, 6.396506, 6.852753, 
    6.698181, 6.010795, 6.102026, 5.957236, 6.195266, 6.354801, 6.32725, 
    6.847486,
  8.36742, 7.635324, 6.500051, 6.124116, 6.522049, 6.895284, 6.927755, 
    6.553693, 6.178686, 5.937274, 5.877733, 5.843189, 5.864657, 6.000105, 
    6.433581,
  9.196681, 8.333322, 8.051425, 8.015608, 7.821414, 7.433978, 6.625197, 
    5.998456, 5.840734, 5.654291, 5.705967, 5.723771, 5.749143, 5.626181, 
    5.656345,
  10.59894, 10.62177, 10.64707, 9.359697, 7.526596, 6.503716, 5.683999, 
    5.578397, 4.739279, 3.887856, 4.163688, 5.543253, 5.432811, 5.334173, 
    5.114191,
  6.807353, 9.124041, 7.113951, 8.122395, 6.005073, 4.372156, 4.796605, 
    3.997174, 3.687266, 2.687089, 2.733318, 3.366975, 3.050505, 2.904996, 
    2.983591,
  8.831664, 8.361941, 7.168569, 5.536273, 3.867169, 3.537392, 4.473014, 
    4.369362, 4.197387, 3.903658, 3.274778, 4.115681, 3.92576, 2.66155, 
    2.193841,
  8.072029, 6.77035, 4.964127, 3.032902, 2.550826, 2.128685, 3.096367, 
    3.60364, 3.714895, 4.107339, 4.59217, 4.922691, 4.922778, 3.589652, 
    1.42828,
  6.717324, 5.488729, 4.102933, 2.783672, 1.847437, 2.264378, 1.496587, 
    3.188708, 5.302355, 4.765328, 4.90771, 5.156133, 5.191102, 4.385972, 
    2.659636,
  5.9424, 4.594004, 4.060941, 4.076907, 3.777309, 3.228359, 2.540616, 
    2.228524, 2.560252, 3.196076, 4.252009, 5.033411, 5.483032, 5.481641, 
    4.992775,
  6.335068, 4.723277, 4.26685, 4.19932, 4.341737, 4.770409, 4.400479, 
    2.78123, 1.514744, 2.435818, 3.135594, 4.629334, 5.375052, 5.880297, 
    6.57367,
  7.181074, 5.045915, 4.306807, 4.241221, 4.438647, 4.526045, 4.717887, 
    4.477593, 3.892189, 3.919939, 3.959473, 4.375764, 5.042978, 5.43095, 
    6.088218,
  7.688771, 5.032829, 4.674617, 4.924415, 4.900226, 4.361449, 3.883674, 
    3.449731, 3.4598, 3.739686, 3.766874, 3.848321, 4.163296, 4.508969, 
    4.916742,
  7.671663, 6.150377, 6.692809, 6.165352, 5.613476, 4.685407, 3.675915, 
    2.897419, 2.947943, 3.236629, 3.327361, 3.27059, 3.180697, 3.213784, 
    3.052262,
  8.947272, 8.731135, 8.634392, 6.93815, 5.409757, 4.211857, 3.241178, 
    2.540363, 2.216949, 1.798685, 1.813828, 2.209969, 2.144483, 1.938732, 
    1.757054,
  8.933265, 12.63888, 10.64474, 13.9363, 12.15591, 9.355865, 11.19816, 
    10.089, 8.628136, 5.115265, 3.688205, 2.742298, 2.204127, 1.982841, 
    1.935941,
  10.98292, 11.38388, 11.49973, 11.15157, 7.909095, 6.552531, 8.956481, 
    7.807144, 6.462614, 4.603543, 2.552436, 1.927439, 2.266265, 2.567001, 
    2.683758,
  8.907149, 8.684194, 8.822289, 8.083841, 6.019164, 4.331905, 5.463171, 
    5.598244, 4.871892, 3.527794, 1.920926, 1.869841, 2.652546, 3.239308, 
    2.685951,
  6.213506, 6.554322, 6.714542, 5.664972, 4.70944, 4.610734, 3.128763, 
    3.931854, 3.823419, 2.728544, 2.338439, 2.696074, 2.491395, 1.767868, 
    1.979356,
  4.763286, 5.413214, 5.699361, 5.214414, 3.619991, 3.207037, 4.485005, 
    2.670512, 0.9432118, 1.376331, 2.727388, 3.193958, 2.400407, 1.906397, 
    2.583785,
  4.482621, 4.857017, 4.93811, 4.446016, 3.839671, 3.122361, 2.598891, 
    3.279921, 2.574504, 1.747135, 2.628631, 3.532408, 3.865379, 3.684774, 
    3.382041,
  4.800951, 4.607007, 4.407052, 3.804446, 3.631621, 4.3687, 4.683091, 
    4.462212, 3.677396, 2.95159, 2.77546, 3.343428, 3.531154, 3.084197, 
    2.328977,
  4.945456, 3.955348, 3.934414, 3.23446, 3.473798, 4.631608, 4.991404, 
    4.31945, 3.033527, 2.1451, 2.19438, 2.684177, 3.115558, 3.230621, 3.059644,
  3.716348, 2.692842, 3.942521, 3.734946, 4.14483, 5.034891, 4.877035, 
    3.465399, 2.287026, 1.93058, 2.194803, 2.804352, 3.550802, 4.408499, 
    4.940699,
  5.190265, 5.662534, 5.546874, 4.937419, 4.519971, 4.388822, 3.917203, 
    3.053207, 2.377297, 1.739889, 2.289557, 3.801101, 5.134641, 6.716304, 
    7.874723,
  9.181049, 13.11982, 11.72984, 15.31936, 14.79456, 12.0352, 15.77458, 
    15.53963, 15.13514, 10.10958, 9.10917, 9.21134, 8.770933, 7.786312, 
    5.733503,
  11.00777, 12.98553, 14.50397, 14.92954, 11.90034, 11.91155, 17.22258, 
    16.18213, 15.02888, 12.42273, 9.41427, 9.916623, 9.205894, 5.815994, 
    4.271616,
  8.753013, 10.24861, 12.11851, 12.30142, 9.274858, 7.565269, 11.07024, 
    13.42954, 12.61765, 11.36473, 9.644917, 8.208684, 7.045415, 6.034934, 
    4.62219,
  6.797002, 8.314024, 9.549659, 9.843519, 9.037498, 6.487185, 4.377428, 
    7.755252, 9.232929, 7.278325, 6.06655, 4.852654, 4.542503, 4.470607, 
    4.387825,
  5.70842, 6.582566, 7.510178, 7.888657, 6.914118, 5.644403, 4.900199, 
    3.332385, 2.963447, 2.867899, 3.606115, 2.889714, 2.465987, 2.610399, 
    3.296868,
  5.010841, 5.262913, 6.140001, 5.977821, 5.707853, 4.605525, 3.750579, 
    3.919556, 3.078466, 1.702433, 2.013566, 1.713802, 1.65304, 1.549415, 
    1.885185,
  6.566417, 5.238867, 4.261615, 3.750982, 3.879555, 4.261562, 3.845536, 
    2.986428, 1.79664, 1.483126, 1.80403, 2.161171, 2.243519, 2.171316, 
    1.89843,
  9.305581, 9.294168, 6.827005, 4.588328, 3.053024, 3.112835, 2.632316, 
    2.767666, 3.089704, 4.201698, 5.098217, 5.591687, 5.609611, 5.363031, 
    4.688654,
  6.971587, 8.490836, 5.8252, 4.36876, 4.439495, 3.278146, 2.933362, 
    3.925439, 5.864307, 7.298258, 8.079697, 9.01154, 8.966953, 8.838226, 
    7.590121,
  4.840448, 5.812581, 6.651137, 7.568285, 5.516306, 4.093489, 4.426734, 
    6.198977, 7.198628, 6.172516, 7.896704, 11.91826, 12.38097, 12.46356, 
    11.12653,
  6.714076, 11.56013, 10.68688, 13.00597, 12.69321, 10.22493, 9.857308, 
    7.138762, 7.123812, 5.275975, 5.209972, 6.883826, 7.826876, 7.184661, 
    5.730278,
  7.222783, 10.48148, 12.80395, 13.09474, 9.999922, 11.44134, 15.61011, 
    12.98468, 10.86195, 8.743242, 6.966595, 8.798603, 10.16635, 6.884584, 
    5.635273,
  7.067636, 8.235501, 10.79074, 12.22121, 9.216439, 7.332664, 11.73979, 
    15.15478, 14.44071, 12.23922, 10.61191, 10.15979, 10.30419, 9.609786, 
    7.083537,
  6.750349, 7.837406, 9.041272, 10.00671, 10.34359, 6.484506, 4.329642, 
    10.54856, 14.42114, 12.40777, 11.18395, 10.78628, 10.56819, 9.179466, 
    7.172898,
  5.807842, 6.177511, 6.852155, 6.670012, 7.28719, 7.66071, 5.171988, 
    4.066459, 5.329873, 6.116657, 7.960858, 8.328808, 9.050336, 8.398044, 
    7.089611,
  6.298443, 4.976714, 4.435468, 3.882715, 2.982712, 3.572549, 4.275075, 
    3.75982, 2.048203, 2.043362, 3.586778, 5.260587, 6.30233, 6.749297, 
    6.745426,
  8.363139, 5.94104, 3.54805, 2.579353, 2.397321, 2.07099, 1.523731, 
    2.288153, 2.726691, 2.35889, 2.643382, 3.672399, 4.556922, 5.180971, 
    5.642932,
  7.505007, 5.496239, 4.653592, 3.390452, 3.357453, 4.031478, 4.404677, 
    4.058021, 6.202883, 6.958578, 6.459185, 5.870418, 5.407043, 5.1408, 
    5.349922,
  6.559212, 6.295129, 4.640364, 3.787896, 4.005131, 5.093758, 5.305789, 
    5.283677, 5.70785, 6.545276, 8.631816, 9.164701, 8.356159, 7.472453, 
    6.129193,
  7.920549, 7.411219, 6.486041, 5.106052, 5.087946, 5.736691, 5.519982, 
    4.617361, 3.850082, 3.331241, 4.830999, 9.901758, 10.94197, 10.10206, 
    7.987736,
  4.180389, 6.168169, 5.668745, 8.351419, 8.721951, 7.778723, 8.894515, 
    3.787718, 1.941056, 2.448217, 2.739174, 3.704023, 3.854388, 3.754405, 
    3.095796,
  5.763111, 6.162735, 5.67428, 6.624306, 5.872149, 6.546904, 10.59215, 
    9.521228, 5.833081, 2.697208, 1.61934, 3.976188, 6.0842, 4.086301, 
    3.373453,
  7.071506, 6.040445, 3.908087, 4.200082, 4.587101, 4.217044, 7.424599, 
    10.03207, 10.5731, 9.288918, 6.257605, 3.52582, 3.810812, 5.696108, 
    4.890101,
  8.550479, 7.991414, 4.162094, 2.526881, 3.871739, 3.447041, 2.555683, 
    7.146793, 11.23398, 10.95975, 9.297104, 7.2772, 4.865152, 3.172613, 
    4.647818,
  9.170203, 8.36085, 4.590378, 2.444665, 1.920238, 2.958726, 2.230921, 
    2.622861, 4.48647, 5.734901, 7.170362, 7.018778, 6.389301, 4.70876, 
    3.336484,
  9.113062, 7.32044, 2.924424, 1.702448, 2.011428, 1.110661, 1.565956, 
    1.532612, 0.7297996, 2.500839, 4.047672, 5.680657, 6.035442, 5.62008, 
    4.881455,
  7.8207, 4.648525, 2.985725, 2.268956, 1.616414, 1.996624, 1.498075, 
    0.9579957, 0.7784835, 1.469261, 2.531255, 4.028845, 5.264916, 5.664977, 
    6.515962,
  5.203276, 4.436409, 4.905917, 2.869181, 2.16095, 2.360906, 2.085, 1.676523, 
    1.302011, 1.46636, 1.403993, 2.283638, 3.763879, 4.906043, 6.003836,
  4.46609, 4.859188, 5.186096, 3.119179, 2.131431, 2.02635, 1.646249, 
    1.288973, 1.945724, 2.114513, 1.337048, 2.30304, 3.10746, 4.063775, 
    4.713543,
  4.507638, 4.828298, 4.334645, 2.343944, 2.18489, 2.22384, 1.926804, 
    1.211731, 1.251309, 1.074523, 1.29796, 1.773316, 3.458335, 3.982415, 
    4.208992,
  4.299973, 4.572807, 3.216139, 2.746847, 2.192267, 2.655215, 5.019428, 
    5.766331, 4.517214, 2.09637, 1.403433, 1.239388, 1.972906, 2.800297, 
    2.631286,
  7.750441, 6.449234, 4.483675, 3.530564, 2.296478, 1.928893, 4.139105, 
    5.712608, 6.498797, 5.358572, 3.154016, 2.170493, 1.77562, 0.9898524, 
    1.005877,
  9.556479, 8.456779, 6.097873, 4.506954, 3.415371, 1.688359, 2.081042, 
    3.21687, 5.09072, 6.667306, 6.776878, 5.650879, 3.392694, 2.60707, 
    1.736146,
  10.40697, 10.42517, 8.404405, 5.579846, 4.735682, 3.390818, 1.493101, 
    2.241912, 5.336684, 5.880439, 6.139112, 6.574358, 6.431525, 4.718031, 
    2.759752,
  10.58465, 10.94737, 9.612772, 6.718136, 5.052522, 3.780158, 3.258166, 
    1.80189, 2.196025, 2.648139, 4.288968, 5.351207, 6.078061, 6.28203, 
    4.716318,
  10.33187, 10.82676, 9.823875, 7.187252, 5.505502, 3.860728, 1.999046, 
    1.835453, 2.187688, 1.767677, 2.611942, 4.087735, 5.242029, 5.938504, 
    6.237403,
  9.858362, 10.30295, 9.76491, 7.497544, 5.86605, 4.774475, 3.344147, 
    2.84036, 2.964615, 2.333542, 2.347682, 3.043882, 4.221778, 5.176788, 
    5.850594,
  9.21613, 9.752844, 9.677572, 7.701788, 5.387705, 4.723897, 4.611523, 
    3.733225, 2.956976, 2.226747, 2.095664, 2.406821, 3.521655, 4.746377, 
    5.580483,
  8.698319, 9.329983, 9.479807, 7.7833, 5.277115, 4.854648, 5.133233, 
    4.178118, 3.363662, 2.531107, 2.090187, 2.050376, 3.138815, 4.470817, 
    5.303863,
  8.49652, 9.290187, 9.222922, 6.962132, 5.359644, 5.300233, 5.252917, 
    4.792628, 3.743461, 1.963314, 1.593533, 1.984758, 2.647186, 3.983359, 
    4.975543,
  2.655463, 3.413733, 3.682619, 6.057751, 5.765499, 2.972319, 2.176325, 
    2.229636, 2.957948, 2.222842, 1.611277, 1.417403, 1.408452, 2.106115, 
    1.930278,
  5.037313, 4.153607, 4.854711, 6.774251, 5.321348, 2.717974, 1.823143, 
    2.275056, 3.057496, 3.5418, 3.085677, 3.309287, 2.469192, 1.928035, 
    1.687955,
  6.636138, 6.431565, 6.237018, 7.605649, 6.384414, 3.078604, 1.490473, 
    1.706368, 2.266664, 3.028497, 3.915357, 4.793106, 4.744298, 3.962957, 
    2.917556,
  7.783188, 8.292048, 8.298461, 8.724997, 8.777021, 5.658094, 2.685153, 
    2.146304, 2.279774, 1.679173, 2.880729, 3.604036, 4.30567, 4.545714, 
    4.029346,
  8.492778, 8.924681, 9.224543, 9.588288, 8.777426, 7.363444, 5.993827, 
    2.671385, 1.870795, 1.894027, 2.350773, 2.465878, 3.279184, 3.75984, 
    3.901818,
  9.117317, 9.499712, 9.713428, 10.12562, 9.560122, 7.435246, 5.949619, 
    4.068042, 2.423132, 3.441428, 3.095746, 2.696088, 2.834047, 3.665516, 
    4.499185,
  8.866316, 9.544811, 9.925311, 10.34565, 10.24671, 8.447514, 5.500404, 
    3.186479, 3.724685, 4.91357, 4.517084, 3.181378, 2.700478, 3.717192, 
    5.069798,
  7.075018, 8.455081, 9.559328, 10.28053, 10.28511, 8.921043, 6.610458, 
    5.657071, 5.238514, 4.782473, 4.494323, 3.291362, 2.836208, 4.226069, 
    5.740092,
  5.093663, 6.819864, 8.347121, 9.596598, 9.519036, 8.001059, 7.419577, 
    6.984467, 5.897707, 4.97144, 4.317304, 3.482777, 3.082431, 4.485919, 
    5.881731,
  4.911364, 6.031469, 7.395377, 7.908233, 7.703626, 7.713835, 8.245022, 
    7.835506, 5.295374, 3.534148, 3.537743, 3.774185, 3.280375, 4.349156, 
    5.727548,
  3.213648, 3.131639, 1.819071, 1.52105, 3.13458, 3.775473, 4.201134, 
    3.332879, 4.4622, 3.588292, 3.389316, 3.628006, 2.937365, 2.645608, 
    1.770232,
  3.688361, 2.935173, 2.534641, 3.128959, 3.213398, 3.744381, 4.821379, 
    3.514113, 3.477027, 3.861848, 3.37558, 4.196087, 3.809705, 2.46497, 
    1.420357,
  3.46019, 4.185769, 4.112935, 3.922202, 3.73186, 2.629889, 4.052079, 
    4.410627, 4.414268, 4.471204, 4.661388, 5.054501, 4.349944, 3.503078, 
    2.372346,
  3.802916, 5.717462, 5.603534, 4.601357, 4.18013, 3.265981, 2.547529, 
    4.303767, 5.13151, 4.561037, 5.52612, 5.691565, 5.057652, 3.952034, 
    2.825493,
  3.627936, 6.093613, 6.218638, 5.111734, 3.67424, 3.098307, 4.528083, 
    2.849633, 2.257366, 2.940844, 4.666784, 4.903395, 4.222312, 2.968188, 
    1.840898,
  3.284883, 6.6545, 7.232192, 5.987168, 5.03033, 3.649756, 3.215405, 
    2.978044, 3.644505, 4.276067, 3.810409, 4.426199, 3.357457, 2.666203, 
    2.812813,
  2.8058, 6.958509, 7.656582, 6.466801, 6.090472, 4.865005, 3.325897, 
    2.343074, 5.147399, 6.329541, 5.707022, 4.371098, 3.02133, 3.032267, 
    3.55914,
  3.064147, 7.318744, 8.073634, 6.611314, 6.376267, 5.774895, 4.880862, 
    4.976156, 6.371394, 6.595588, 5.789921, 4.010737, 3.09404, 3.611454, 
    4.231545,
  3.430907, 7.569471, 8.826347, 7.162249, 6.603192, 6.466393, 5.687428, 
    5.70614, 6.415429, 6.219902, 5.253743, 3.697103, 3.26188, 3.97651, 
    4.348477,
  3.543499, 6.672317, 8.730539, 7.164937, 6.099807, 6.485456, 6.75035, 
    6.685686, 5.567986, 4.081356, 3.844059, 3.609652, 3.329228, 4.125678, 
    4.507218,
  5.530205, 6.250065, 4.348656, 5.028918, 3.465563, 3.113167, 4.669001, 
    4.159874, 3.053542, 2.165881, 2.246592, 3.311704, 4.011841, 3.921091, 
    3.050169,
  7.496229, 6.639652, 6.162572, 5.741653, 3.341407, 2.552392, 3.916958, 
    3.622379, 2.638955, 2.581893, 2.580409, 4.142756, 5.568186, 3.466331, 
    2.979677,
  7.065361, 6.448265, 6.710683, 6.460086, 4.060613, 2.181515, 2.866496, 
    3.311291, 3.272834, 3.507001, 3.9653, 4.592401, 5.165792, 5.228354, 
    4.232298,
  6.601122, 7.022759, 7.980389, 6.646387, 4.034545, 2.486001, 1.256644, 
    3.483155, 5.516728, 5.026339, 5.47837, 5.946182, 6.105325, 5.5905, 
    4.489399,
  6.133731, 8.226214, 9.265897, 6.4002, 2.597295, 1.619999, 2.767957, 
    2.196144, 2.065088, 3.254878, 5.371854, 6.271091, 6.350683, 5.74043, 
    4.285623,
  7.587534, 9.924611, 9.43838, 5.767109, 2.925173, 1.288329, 1.320519, 
    3.510117, 4.0756, 3.935264, 4.222139, 5.655923, 5.390379, 4.995909, 
    3.897138,
  9.796251, 10.78021, 9.05715, 5.352292, 3.052191, 2.905793, 4.147434, 
    4.916526, 5.79678, 6.215475, 5.996344, 5.381734, 4.585981, 4.088945, 
    3.392522,
  10.91321, 10.7186, 8.23959, 4.897991, 4.121412, 5.346821, 6.29471, 
    6.645581, 6.933332, 6.632696, 5.719083, 4.606791, 3.883716, 3.659122, 
    3.385519,
  11.08407, 10.25726, 7.473332, 5.732379, 6.331406, 6.832181, 6.519651, 
    6.534908, 6.616066, 5.59047, 4.618542, 3.863083, 3.631714, 3.796288, 
    3.47271,
  10.72166, 9.865647, 7.898799, 6.86658, 6.473637, 6.4201, 6.210479, 
    6.097027, 4.808072, 3.218984, 3.11221, 3.365847, 3.394247, 3.565579, 
    3.545329,
  4.596758, 7.02112, 6.321066, 8.583488, 7.562239, 5.153273, 6.62885, 
    6.338374, 5.428856, 4.032948, 3.921038, 4.498856, 4.344049, 4.164762, 
    3.797297,
  6.850652, 7.587802, 7.619163, 7.542422, 3.696209, 4.091378, 5.576503, 
    5.268101, 4.731496, 3.871149, 3.340271, 4.710061, 6.019967, 4.17311, 
    3.660585,
  7.34382, 6.752494, 6.624101, 5.669584, 5.653619, 4.955882, 4.655605, 
    4.385701, 3.722146, 2.697479, 2.222432, 3.455669, 5.511128, 6.330976, 
    5.380731,
  7.493269, 6.854589, 6.634005, 7.727946, 7.845821, 5.024106, 3.578867, 
    3.875199, 4.157333, 3.028644, 1.491765, 2.339915, 4.595984, 6.045479, 
    6.486456,
  7.568204, 7.88624, 9.152049, 9.383375, 7.926709, 5.580814, 4.554688, 
    2.926377, 1.571719, 1.575846, 2.274393, 2.497187, 5.118585, 6.732787, 
    7.266587,
  9.109754, 9.38274, 9.212757, 8.582067, 7.573466, 6.298562, 5.041969, 
    4.065621, 2.797183, 2.355834, 2.61148, 4.153255, 5.950121, 7.287766, 
    7.521283,
  9.616075, 9.240609, 8.668174, 7.796725, 7.020594, 6.937008, 6.700441, 
    5.974594, 5.257016, 5.051615, 5.17659, 6.219406, 7.424488, 8.384464, 
    8.97604,
  9.218278, 8.968129, 8.574813, 8.124071, 7.723718, 7.590091, 7.194547, 
    6.853125, 6.600998, 6.383423, 6.657809, 7.352658, 7.977158, 8.701903, 
    8.909435,
  8.254478, 8.528157, 8.495124, 8.372562, 8.143888, 7.73815, 7.00154, 
    6.784594, 6.769297, 6.408043, 6.749629, 7.390018, 7.67099, 7.898256, 
    6.787302,
  6.646924, 7.065726, 7.137675, 6.542143, 6.077387, 6.201035, 5.930054, 
    5.81261, 5.102727, 4.006207, 4.624669, 6.530742, 6.547353, 6.357418, 
    5.608847,
  4.007155, 5.212507, 5.177567, 7.215271, 6.579455, 4.389714, 5.370503, 
    5.787821, 5.068422, 3.472503, 3.30725, 3.705398, 3.80897, 4.288052, 
    4.824895,
  5.116595, 4.980296, 5.272219, 7.030739, 5.247229, 4.136146, 5.405674, 
    5.523267, 5.261274, 4.743004, 3.836553, 4.042168, 4.071477, 2.866246, 
    3.819068,
  5.365892, 4.036645, 4.229584, 6.145126, 5.745682, 3.749592, 4.845569, 
    4.911935, 4.454433, 4.74206, 4.610852, 4.172168, 4.050005, 4.65553, 
    5.458092,
  6.866332, 7.43815, 7.417689, 6.704844, 7.601987, 5.881294, 3.287648, 
    4.402752, 6.297812, 5.413006, 4.163486, 2.880849, 3.660437, 4.984319, 
    6.126682,
  7.018579, 7.821485, 8.38773, 7.578844, 7.049031, 7.795364, 5.964621, 
    3.170521, 3.717753, 3.822631, 3.673659, 2.063841, 3.662388, 5.564099, 
    6.71393,
  6.822623, 7.631293, 8.534897, 8.25275, 7.346864, 7.811225, 8.083214, 
    6.447409, 4.757772, 3.989417, 2.395247, 2.48888, 4.297789, 5.793304, 
    6.278193,
  6.38152, 7.224325, 8.207752, 8.809416, 8.530273, 8.174342, 8.317059, 
    8.310685, 7.585647, 6.242518, 4.327268, 4.301663, 5.464783, 6.245535, 
    7.112971,
  5.830729, 6.456906, 7.16512, 8.373369, 9.102818, 8.846511, 8.128154, 
    7.993776, 8.201088, 7.835663, 6.661909, 6.602293, 7.029846, 7.711701, 
    8.42747,
  5.774872, 5.771883, 5.631555, 6.324038, 7.556821, 8.005405, 7.59142, 
    7.664025, 8.04439, 8.296699, 8.058366, 8.086936, 8.264865, 8.349346, 
    7.289204,
  5.987809, 5.355644, 4.446199, 3.745453, 4.82732, 6.337551, 6.847159, 
    6.866543, 6.283371, 5.215593, 5.598852, 7.855842, 7.804135, 7.541958, 
    6.300257,
  4.397202, 4.348351, 3.685079, 4.917318, 5.086413, 4.203467, 5.908451, 
    6.195679, 5.350577, 3.995894, 4.262474, 4.604365, 3.553554, 2.907412, 
    2.558155,
  6.138947, 4.404757, 4.055943, 4.496314, 4.198717, 4.08277, 6.136395, 
    6.610194, 6.33562, 5.261529, 4.26008, 4.500748, 2.860173, 1.974155, 
    2.163019,
  6.350414, 4.131943, 3.741776, 3.870939, 4.200151, 3.509809, 5.647336, 
    6.296444, 5.68375, 5.520862, 5.259545, 4.35856, 3.001687, 2.549492, 
    4.428608,
  7.365188, 6.076111, 6.139303, 4.460297, 5.167321, 4.686858, 3.502344, 
    5.60323, 8.751656, 8.184301, 6.744844, 5.583506, 5.10619, 5.625607, 
    6.435296,
  7.599554, 5.96784, 6.529662, 6.094005, 4.819973, 5.665895, 4.960911, 
    3.405502, 4.937439, 5.581117, 6.81768, 6.765988, 6.845968, 7.414542, 
    7.778358,
  8.253222, 5.801217, 6.313159, 6.499375, 5.525357, 5.164592, 5.766839, 
    5.148915, 3.967426, 4.50115, 4.677162, 7.321852, 8.024026, 8.539442, 
    8.580484,
  8.73038, 6.051154, 5.864623, 6.831719, 5.855355, 5.205044, 5.331966, 
    6.107622, 6.524114, 6.936315, 6.60336, 7.337554, 7.976656, 8.525998, 
    9.07717,
  9.563788, 7.033384, 5.342176, 7.385615, 6.370974, 5.294985, 4.927736, 
    5.211631, 5.980787, 6.539163, 6.78172, 7.041519, 7.434502, 7.959757, 
    8.209147,
  10.44634, 8.086143, 5.03802, 8.079563, 7.519607, 5.663121, 4.636438, 
    4.348542, 5.148601, 5.785421, 6.193146, 6.407738, 6.617872, 6.735303, 
    6.167296,
  10.94412, 8.846152, 5.763844, 7.82883, 9.725867, 6.679091, 4.613615, 
    4.119566, 3.909941, 3.453247, 3.990667, 5.312953, 5.180909, 4.949526, 
    4.504261,
  7.017314, 6.009379, 7.635952, 8.175966, 4.726665, 2.758483, 3.002658, 
    3.54646, 3.760348, 3.095459, 3.409144, 3.983519, 4.019845, 3.400181, 
    2.683553,
  10.5929, 6.593845, 10.63129, 8.389393, 4.097288, 3.164072, 4.323673, 
    4.805409, 5.228672, 3.881326, 2.098542, 2.897654, 4.514848, 3.29515, 
    2.638412,
  10.27293, 6.940237, 11.30731, 8.464349, 4.750302, 2.522837, 4.505389, 
    5.681637, 6.182662, 5.84776, 4.810209, 4.444657, 4.400125, 4.521682, 
    3.553662,
  9.971231, 7.170192, 11.41359, 8.83647, 5.420275, 3.700067, 2.225171, 
    5.516699, 9.897442, 8.92067, 7.134856, 6.104386, 5.207756, 4.203278, 
    3.795086,
  9.964257, 7.883896, 10.8931, 10.61452, 6.698012, 5.379653, 4.320599, 
    3.385959, 5.002897, 5.697402, 6.892425, 6.665791, 6.254649, 5.299433, 
    4.567837,
  10.11054, 9.026964, 10.16592, 12.48347, 9.224872, 7.702087, 6.723919, 
    6.10544, 3.723334, 4.858142, 5.449049, 7.941567, 8.209489, 7.987656, 
    7.73316,
  10.23565, 10.34508, 10.41031, 13.59895, 10.57414, 9.156338, 7.801009, 
    7.422705, 7.495994, 8.225508, 8.028272, 8.728455, 8.854885, 8.778734, 
    8.676483,
  10.39291, 10.91601, 10.68856, 13.80491, 11.32786, 9.812711, 8.284776, 
    7.950888, 7.833326, 8.068604, 8.167875, 8.397985, 8.33637, 8.461627, 
    7.993256,
  10.33517, 10.72343, 10.9563, 14.1122, 12.26036, 10.45848, 8.524474, 
    7.787858, 7.557091, 7.366313, 7.536875, 7.698954, 7.75028, 8.036801, 
    7.741229,
  10.18066, 10.16878, 10.95395, 13.70377, 12.52752, 10.31137, 8.619662, 
    7.590051, 5.877256, 4.754426, 5.285691, 7.503208, 7.404661, 7.767132, 
    7.784039,
  6.735251, 8.593094, 6.013465, 6.656524, 5.788588, 5.206618, 5.580133, 
    2.941958, 1.478409, 1.994853, 2.88095, 3.835838, 4.170156, 4.037362, 
    3.563703,
  9.845153, 8.685614, 7.374119, 5.922732, 4.40455, 4.934627, 7.174548, 
    5.847574, 3.217604, 1.744008, 2.760353, 4.304909, 5.443959, 3.794063, 
    3.428433,
  10.25306, 8.598551, 7.873216, 6.98143, 5.215424, 3.633089, 6.102593, 
    6.48616, 4.983178, 3.019213, 3.13136, 4.249056, 5.251079, 5.586034, 
    4.691283,
  10.02292, 9.255935, 8.896137, 8.479557, 8.347184, 5.829399, 3.224273, 
    6.009656, 8.737659, 5.669368, 2.830338, 3.524357, 5.117895, 5.941002, 
    5.910652,
  10.06864, 9.760349, 9.649944, 9.68277, 9.721323, 9.395734, 7.140353, 
    4.225637, 5.087614, 4.727176, 4.091534, 3.255225, 4.458701, 6.014872, 
    7.369195,
  10.12117, 9.958644, 9.906973, 9.904728, 10.21417, 10.79558, 10.61357, 
    9.025954, 6.006954, 5.775167, 3.851494, 3.652087, 3.973213, 4.928133, 
    6.116441,
  10.07072, 10.15192, 10.1473, 10.28801, 10.63437, 10.88567, 10.9017, 
    11.0077, 11.44601, 11.41365, 8.950985, 5.433736, 4.15829, 4.265644, 
    5.180583,
  10.20623, 10.45019, 10.5681, 10.90765, 11.25677, 11.163, 10.98646, 
    11.27961, 11.78936, 12.53364, 12.19423, 9.361794, 6.112007, 4.87158, 
    4.988081,
  10.42565, 10.72374, 10.87278, 11.0466, 11.12784, 10.94328, 10.95766, 
    11.3565, 11.83988, 12.38731, 13.22483, 12.68684, 9.539623, 7.122937, 
    6.134631,
  10.7664, 10.99806, 10.98173, 10.76848, 10.50628, 10.46523, 10.13439, 
    10.66608, 9.389489, 7.996468, 9.643641, 13.62806, 12.4796, 9.916165, 
    7.694248,
  3.147098, 4.506719, 4.803689, 5.872737, 4.279723, 3.562809, 4.405045, 
    3.463586, 2.279666, 1.883888, 1.804398, 2.814018, 2.970123, 3.106664, 
    3.64239,
  3.600337, 4.009491, 6.37694, 6.675806, 4.443701, 3.692502, 5.256959, 
    4.339206, 2.111879, 2.341742, 1.383815, 2.400036, 3.511693, 2.765628, 
    3.14451,
  5.283635, 4.120203, 5.925281, 7.935366, 6.283111, 3.599502, 5.318992, 
    5.039168, 2.175535, 2.10182, 2.85414, 2.309388, 3.543442, 3.910249, 
    3.698262,
  6.671097, 7.085452, 7.676769, 8.470203, 9.161263, 6.648427, 3.763818, 
    4.909752, 6.232865, 1.794448, 3.014253, 3.239023, 3.658469, 4.600595, 
    4.441005,
  7.334021, 8.115564, 8.454964, 8.476722, 9.135614, 9.538419, 6.943838, 
    3.632034, 4.185579, 2.855028, 1.906628, 4.01066, 4.112788, 4.779595, 
    5.282991,
  7.671347, 8.523319, 8.85862, 9.001515, 9.290334, 9.77247, 9.335911, 
    7.042622, 5.06898, 3.802109, 1.45116, 4.151901, 4.732996, 4.856647, 
    5.412839,
  8.016011, 8.920809, 9.479537, 9.883525, 10.25152, 10.27199, 9.917336, 
    9.290854, 9.017709, 7.466576, 2.401215, 3.510498, 4.633615, 5.139052, 
    5.425382,
  8.080739, 9.138443, 9.9752, 10.75331, 11.08182, 10.97369, 10.4092, 
    9.425683, 9.234733, 9.246675, 6.089331, 2.182959, 4.512594, 5.289927, 
    5.625956,
  8.065344, 8.998033, 9.836545, 10.60917, 10.9677, 11.11761, 11.17597, 
    10.50808, 10.04063, 9.811533, 8.703123, 4.022555, 3.16284, 5.394681, 
    5.881886,
  7.768325, 8.628949, 9.336848, 10.02389, 10.5492, 11.08869, 11.30782, 
    11.12834, 8.949922, 6.616657, 6.68038, 7.405001, 2.958947, 4.261409, 
    5.757795,
  2.863268, 3.500072, 3.324294, 3.64834, 2.21959, 1.985795, 3.16348, 
    3.676548, 3.354009, 3.006743, 3.149232, 3.289993, 2.927173, 2.542456, 
    2.563128,
  2.188134, 2.052257, 3.99236, 4.410567, 2.820272, 2.558352, 3.828746, 
    4.141441, 3.696092, 3.321012, 3.256749, 3.479881, 3.457672, 2.702554, 
    2.815333,
  3.318106, 2.265729, 3.003447, 4.913236, 4.359295, 2.992944, 4.319507, 
    3.97901, 2.825653, 2.385048, 3.500928, 3.329794, 3.503647, 4.052084, 
    3.646657,
  5.23635, 4.588008, 4.616124, 4.995283, 6.020556, 4.952785, 3.213931, 
    4.148595, 5.496555, 2.947039, 2.358164, 2.857767, 3.056464, 3.91417, 
    3.395072,
  6.322681, 6.42601, 6.163143, 5.857523, 6.08138, 6.702093, 5.313141, 
    2.92154, 3.630798, 3.391545, 2.479411, 2.357944, 2.051855, 3.632978, 
    3.932232,
  6.993645, 7.262748, 7.259206, 7.104339, 7.125558, 7.489276, 6.862209, 
    4.749669, 4.354042, 3.721075, 1.950926, 2.125671, 1.200917, 3.153314, 
    4.776194,
  7.371143, 7.819649, 8.312229, 8.760053, 8.971271, 8.602974, 8.007187, 
    6.857643, 6.425264, 5.089179, 1.251872, 2.215588, 1.127777, 2.770377, 
    4.798377,
  7.404276, 8.14269, 8.951765, 9.792616, 10.20751, 9.861816, 8.982486, 
    7.671893, 7.249698, 6.502784, 2.976, 1.749632, 1.782964, 2.745982, 
    4.665901,
  7.357185, 7.915068, 8.591231, 9.332996, 9.790495, 10.08805, 10.19658, 
    9.66558, 9.10239, 8.302744, 5.989112, 1.396327, 2.467186, 2.916835, 
    4.229303,
  7.074299, 7.277792, 7.48632, 7.786295, 8.498025, 9.62723, 10.49227, 
    10.67502, 8.909922, 6.88395, 5.896163, 3.741861, 1.89032, 3.055609, 
    3.966806,
  5.137158, 6.365047, 4.707055, 5.01077, 4.281831, 3.216679, 2.936878, 
    2.35254, 2.161019, 2.249683, 2.839856, 3.677411, 3.540861, 3.200533, 
    2.7742,
  5.233267, 4.855487, 5.086246, 4.099685, 2.806047, 2.481276, 2.963236, 
    2.641284, 2.712123, 3.171139, 3.639381, 4.765402, 5.33513, 3.443403, 
    2.959581,
  4.328739, 2.721827, 4.080815, 4.449905, 3.564614, 2.416791, 3.341309, 
    2.939027, 2.398381, 3.060131, 4.074055, 4.831275, 5.787648, 6.081452, 
    4.269075,
  4.269543, 3.961187, 4.153632, 4.199409, 5.376405, 3.899087, 2.638022, 
    3.629593, 4.276242, 3.03948, 2.753759, 3.408386, 4.542792, 5.457705, 
    5.333923,
  4.603538, 4.682399, 4.736611, 4.117258, 4.694311, 5.424877, 3.902256, 
    2.674179, 3.301537, 3.381633, 3.233692, 2.820757, 3.53933, 4.339622, 
    5.664928,
  3.952327, 4.299052, 4.650633, 4.705749, 5.145071, 5.742414, 5.377385, 
    3.94045, 3.683973, 3.503963, 2.672848, 2.50108, 2.553194, 3.322163, 
    4.525619,
  3.320659, 4.008035, 4.623409, 5.383753, 6.14418, 6.055136, 6.190962, 
    5.670473, 5.241075, 4.605243, 3.293227, 2.152986, 2.117156, 3.150353, 
    4.610837,
  2.995064, 3.823109, 4.775092, 5.664287, 6.385307, 6.408453, 6.65487, 
    6.105189, 5.639097, 5.269191, 4.285251, 3.010025, 3.019356, 4.107893, 
    5.284472,
  2.612879, 3.232167, 4.212482, 5.075799, 5.768156, 6.415647, 7.239879, 
    7.22192, 6.749896, 6.029038, 5.627769, 4.51883, 3.658047, 4.286097, 
    5.043276,
  2.72939, 3.143926, 4.311642, 5.283004, 6.288626, 6.978086, 7.469135, 
    7.928956, 6.624732, 4.796696, 4.923618, 5.732574, 4.264913, 4.175828, 
    4.5286,
  3.768456, 4.621556, 3.378977, 3.269908, 2.310895, 2.13436, 3.195608, 
    3.693029, 3.643469, 3.378, 3.852706, 4.242917, 4.168421, 4.359154, 
    4.204696,
  2.600227, 2.53545, 2.866326, 3.120301, 2.764094, 3.197452, 4.72927, 
    4.981407, 4.978683, 4.22099, 3.457133, 3.703867, 3.640863, 2.786051, 
    2.984635,
  3.491566, 4.149375, 4.830566, 5.830877, 4.894716, 3.731752, 5.207658, 
    5.764956, 5.583993, 5.784593, 5.819061, 5.560789, 5.244434, 4.826178, 
    3.420279,
  4.922343, 6.101369, 7.080131, 7.426317, 8.547017, 7.302141, 5.381006, 
    5.306284, 7.23508, 7.611067, 7.475981, 7.192229, 6.704388, 6.476033, 
    5.7402,
  6.323097, 8.002919, 8.860147, 8.267013, 9.50502, 9.415774, 8.610518, 
    5.869024, 6.139829, 6.370485, 8.37359, 9.190074, 7.948299, 7.827123, 
    8.077088,
  8.956412, 9.948202, 9.384739, 8.391082, 9.618307, 10.27569, 10.90193, 
    10.69389, 9.00298, 7.137362, 6.74073, 9.319983, 8.810594, 8.542075, 
    8.372696,
  10.63777, 9.821877, 8.805327, 8.929187, 9.903095, 9.532039, 10.24756, 
    11.05608, 10.39455, 10.08818, 9.748589, 10.13, 9.633837, 8.942726, 
    8.371419,
  10.14092, 8.636889, 8.772447, 9.358495, 9.734528, 9.287442, 9.409169, 
    10.25744, 10.64065, 10.83538, 10.71886, 10.49794, 9.796032, 9.192084, 
    8.593546,
  8.477361, 8.1551, 8.916659, 9.266773, 9.245569, 9.1369, 9.978216, 11.21163, 
    11.39443, 10.82667, 10.52868, 10.09307, 10.05104, 9.512473, 8.381189,
  7.119902, 7.764457, 8.729387, 8.769807, 9.111691, 9.376992, 10.24539, 
    11.1869, 9.919512, 7.434291, 7.98271, 10.34896, 9.526193, 9.462411, 
    8.137463,
  3.349769, 4.781948, 4.717046, 5.013167, 3.261989, 2.457854, 3.671098, 
    4.209255, 4.3258, 3.576613, 3.602702, 4.256979, 3.584373, 2.944923, 
    2.806767,
  5.760389, 6.737896, 7.62235, 7.819958, 4.909075, 4.325331, 6.775561, 
    7.347939, 7.739737, 7.250622, 6.356989, 7.639456, 7.541894, 5.026417, 
    4.633189,
  8.281878, 8.610403, 10.01808, 10.16963, 6.40217, 4.395743, 5.415417, 
    6.689916, 7.469416, 7.880731, 8.462403, 9.33154, 10.23667, 10.53653, 
    7.301083,
  10.66541, 12.48549, 12.74699, 10.03253, 6.095386, 4.233013, 3.669071, 
    4.487644, 5.296177, 6.166537, 7.858568, 8.825026, 9.484912, 10.72883, 
    9.481247,
  12.37977, 13.99111, 12.72311, 6.185439, 5.253111, 4.966657, 4.742967, 
    3.806627, 4.555583, 5.132082, 7.390146, 8.832026, 8.841529, 9.601233, 
    11.49835,
  13.6906, 12.94321, 7.447946, 4.816825, 6.414325, 7.45016, 7.093992, 
    6.180014, 5.254102, 5.017708, 5.874152, 9.637832, 10.05476, 10.55991, 
    11.01712,
  12.9959, 8.698565, 5.31636, 6.240417, 7.628657, 5.924661, 5.745175, 
    6.349652, 7.157805, 8.426644, 9.544491, 10.83799, 11.82892, 11.95403, 
    11.78069,
  9.257873, 6.737713, 6.618832, 7.399226, 6.71425, 6.698296, 6.203581, 
    6.696828, 8.678884, 10.15802, 10.89472, 11.41223, 11.9355, 11.6193, 
    11.49109,
  7.692203, 7.296361, 6.88837, 6.502803, 6.612267, 5.939624, 7.215243, 
    9.500479, 10.82331, 11.54622, 11.15829, 10.40753, 9.86008, 9.696324, 
    9.089722,
  7.550208, 7.178907, 6.732379, 6.408842, 5.961302, 6.695157, 8.769803, 
    10.40981, 9.940824, 8.105594, 8.260255, 9.357061, 7.23542, 6.962642, 
    6.685326,
  3.381097, 5.654964, 6.567787, 9.298553, 9.583117, 7.233143, 7.301142, 
    5.416293, 4.925996, 3.710887, 3.49655, 3.454714, 2.38713, 2.163035, 
    2.307427,
  6.311053, 7.807475, 9.369683, 10.60509, 7.618958, 4.857646, 4.57462, 
    5.916036, 6.676645, 6.109573, 5.686225, 6.546392, 5.956516, 2.99464, 
    2.02417,
  8.943481, 9.336801, 10.85186, 11.84486, 6.266838, 2.941783, 4.966224, 
    5.168726, 5.327308, 6.461246, 7.389677, 7.836381, 7.723239, 6.880043, 
    4.36256,
  10.4014, 12.14177, 13.19997, 7.780651, 3.143768, 3.005662, 3.227947, 
    4.81672, 5.314606, 6.62155, 7.94249, 8.147317, 8.030183, 8.036681, 
    6.443399,
  11.20665, 12.60025, 9.636737, 4.194529, 5.549096, 4.158841, 3.17538, 
    3.065865, 4.498383, 5.635445, 7.897432, 8.305407, 7.847022, 8.197412, 
    8.676125,
  11.22621, 8.6589, 3.404835, 6.244145, 3.896364, 3.975118, 4.778515, 
    4.432303, 5.131704, 5.257406, 5.230126, 7.274816, 7.125096, 7.375922, 
    7.997086,
  7.596602, 3.164748, 5.119858, 2.559513, 3.639392, 3.247909, 5.36969, 
    6.934583, 7.439285, 7.136899, 6.762051, 6.816481, 6.960735, 7.268905, 
    7.922257,
  3.911257, 4.881298, 2.650887, 3.160273, 4.145364, 4.762133, 6.239089, 
    7.390624, 7.816797, 7.374683, 6.853887, 7.083786, 7.96844, 8.509641, 
    9.403666,
  6.452739, 4.044165, 3.170352, 3.628217, 4.683999, 6.195495, 7.920039, 
    8.785092, 8.255791, 7.401836, 6.569639, 7.192877, 8.812731, 9.52625, 
    8.968075,
  6.842703, 4.555626, 4.043464, 4.400224, 5.577618, 7.412194, 8.397295, 
    8.393729, 6.649351, 4.708823, 5.622563, 8.018125, 8.554915, 8.471377, 
    6.446541,
  4.877141, 6.097232, 5.26614, 6.321538, 6.279653, 5.822381, 8.285276, 
    6.905836, 4.762, 2.6403, 3.095186, 4.04387, 4.708833, 4.868396, 4.734977,
  7.524161, 7.491811, 7.396045, 7.681952, 5.045675, 4.749011, 6.357161, 
    4.619868, 2.878788, 2.92235, 3.790129, 5.210786, 6.148961, 4.922032, 
    5.360183,
  8.352903, 8.326014, 8.277662, 8.831391, 6.553121, 4.317513, 3.984531, 
    3.349994, 3.18241, 4.176192, 5.579005, 6.581509, 7.144022, 7.480835, 
    6.418639,
  8.025884, 9.111281, 9.704985, 9.341156, 7.699974, 5.22292, 2.379769, 
    2.522862, 3.469652, 4.617725, 6.160417, 7.330284, 7.71543, 8.112208, 
    6.710906,
  7.917638, 8.778609, 9.501494, 7.393722, 6.286183, 5.371848, 4.764415, 
    2.863457, 4.05484, 4.642933, 6.465098, 8.010402, 8.14242, 8.682849, 
    8.617391,
  8.192232, 8.730947, 8.03092, 6.850433, 5.970149, 5.019116, 4.834066, 
    5.218452, 5.019958, 4.698425, 5.417342, 8.489943, 8.868702, 8.937844, 
    8.790593,
  8.716963, 8.483632, 7.5194, 5.802631, 4.882894, 3.017133, 2.786722, 
    3.835255, 5.658218, 7.106773, 7.976122, 8.568663, 8.527312, 8.509609, 
    8.702507,
  9.174378, 8.057794, 7.344306, 5.772896, 4.660107, 3.839241, 3.408458, 
    4.690281, 6.78792, 7.406372, 7.036882, 7.200563, 7.750978, 8.29135, 
    8.990889,
  6.897754, 8.452795, 7.913337, 5.86986, 4.546245, 3.956599, 4.473063, 
    6.178144, 7.10669, 6.646144, 5.68856, 6.77549, 8.029216, 8.907675, 
    8.929192,
  7.330835, 7.723237, 7.000081, 6.152135, 4.359185, 3.78284, 4.488925, 
    6.136101, 5.670326, 4.192778, 5.025443, 7.133782, 8.040771, 9.142536, 
    8.789962,
  3.716071, 5.88463, 6.006604, 7.98495, 7.587369, 6.341441, 7.766815, 
    8.160785, 7.568537, 5.459877, 5.131597, 5.426785, 4.532355, 4.094138, 
    4.253998,
  5.24329, 6.412721, 7.369294, 8.018457, 5.774964, 4.754699, 7.756246, 
    8.103565, 8.005587, 7.239934, 5.941856, 6.528536, 6.597935, 4.59907, 
    4.348785,
  5.656244, 6.76145, 7.709749, 8.668441, 6.937169, 4.480491, 5.817256, 
    7.782506, 7.883132, 7.793018, 7.550595, 7.469329, 7.802547, 7.847431, 
    6.075355,
  5.904345, 7.450434, 8.942603, 9.935773, 10.24259, 7.482007, 4.291843, 
    4.370042, 6.020327, 8.112254, 8.448177, 8.363579, 7.996899, 8.147392, 
    7.199672,
  6.319826, 7.343106, 9.046626, 10.19127, 9.96945, 10.18134, 8.086107, 
    5.243581, 4.730884, 5.333842, 7.142734, 8.094687, 7.8167, 8.396537, 8.4989,
  6.492655, 6.775328, 8.21066, 9.540665, 10.04251, 9.723605, 10.32377, 
    9.899494, 6.612349, 3.826364, 3.82108, 6.068512, 6.364768, 6.796319, 
    7.46663,
  6.280407, 6.182994, 7.055225, 8.337295, 9.552208, 8.950044, 8.520253, 
    7.938957, 6.567246, 5.341694, 4.685809, 4.815875, 5.575642, 6.268142, 
    7.153998,
  5.427825, 5.324474, 5.915055, 7.121586, 8.398583, 7.697282, 7.515631, 
    6.843037, 5.143019, 4.380856, 4.503246, 4.97539, 5.474617, 6.517367, 
    8.539714,
  4.394516, 4.936242, 6.133009, 6.89051, 5.829907, 5.811954, 5.841555, 
    5.109279, 4.780968, 4.643316, 4.348553, 4.559, 6.019354, 8.162159, 
    9.677949,
  5.036506, 4.503013, 5.017933, 5.610029, 7.127327, 8.795297, 8.461867, 
    6.657609, 4.764401, 3.197883, 3.087732, 5.199017, 7.351007, 9.645195, 
    10.66413,
  5.279352, 7.398857, 6.188842, 8.062771, 7.384412, 6.053782, 7.648091, 
    8.288631, 8.20425, 6.49378, 6.804005, 8.064036, 7.63795, 7.05282, 6.772824,
  7.058001, 7.279212, 6.978424, 7.205485, 4.98578, 4.810221, 7.089266, 
    7.989904, 8.432391, 8.030289, 7.813762, 10.40615, 11.04038, 7.5378, 
    6.811099,
  6.494901, 5.353679, 5.699671, 6.06222, 5.026644, 4.067032, 4.666127, 
    6.030793, 7.697678, 8.366125, 8.606699, 10.12122, 11.47316, 10.60749, 
    7.66106,
  4.743029, 4.357486, 4.618295, 4.268599, 5.514885, 4.864006, 3.808489, 
    3.50191, 4.481721, 6.749999, 7.757684, 8.557752, 9.801394, 9.77701, 
    8.704462,
  3.808903, 3.942549, 3.423982, 3.490527, 4.009559, 5.299709, 5.992938, 
    4.41227, 2.82022, 3.897577, 6.652672, 7.689423, 8.315649, 9.381671, 
    10.69269,
  3.627918, 3.506987, 3.407693, 4.574921, 5.373312, 4.836806, 5.28457, 
    5.400009, 3.719802, 3.323335, 4.021486, 6.168681, 6.922062, 7.753381, 
    8.537244,
  4.698017, 4.154902, 4.503836, 5.863219, 6.716462, 6.398791, 5.475893, 
    4.459192, 4.093088, 4.260278, 4.475525, 4.340611, 3.771081, 3.58563, 
    3.553741,
  7.107863, 6.678009, 7.067274, 7.847039, 8.120215, 7.597869, 6.986395, 
    6.708508, 6.030072, 5.49147, 5.231965, 5.354787, 5.267434, 4.21556, 
    3.204587,
  9.936207, 9.538785, 9.461057, 9.49991, 9.224304, 8.845977, 8.577232, 
    8.59208, 8.706805, 8.615043, 8.193873, 7.180003, 5.174729, 3.652605, 
    3.261007,
  12.3043, 12.28582, 12.03778, 11.63656, 11.5283, 11.31019, 10.84826, 
    9.92223, 7.297513, 4.674092, 3.763805, 3.100143, 2.440162, 3.252425, 
    4.187578,
  6.218492, 8.260777, 7.567139, 10.05772, 9.331735, 7.956689, 10.04462, 
    10.36215, 9.886511, 6.80656, 5.966089, 6.206025, 4.847787, 4.316322, 
    4.269813,
  7.809103, 7.865151, 8.184283, 8.143619, 5.783537, 5.858934, 8.822469, 
    8.97148, 9.19402, 8.262157, 6.883191, 7.565322, 7.105604, 4.392684, 
    3.985159,
  8.104725, 7.068769, 6.936589, 6.905678, 5.111057, 4.487309, 6.026703, 
    6.670161, 6.462053, 7.014635, 7.159947, 6.657639, 6.806518, 6.189365, 
    4.763966,
  8.672322, 8.627823, 8.313741, 7.513737, 6.265177, 4.175173, 2.601961, 
    2.880095, 3.523701, 4.352267, 4.794472, 5.240045, 5.388599, 5.55148, 
    5.094715,
  9.136581, 9.135276, 9.152264, 8.647245, 8.171873, 6.483603, 4.242887, 
    2.361805, 2.102326, 2.239404, 2.76441, 3.162105, 3.471588, 4.040023, 
    4.841073,
  9.686349, 9.550535, 9.597262, 9.625074, 9.831469, 9.835409, 8.103793, 
    5.556935, 3.866637, 4.102674, 3.528312, 3.835112, 3.773268, 3.792274, 
    3.807334,
  9.788415, 9.762583, 9.8189, 10.12546, 10.50639, 10.78176, 10.80564, 
    10.32678, 9.85638, 9.656783, 9.128321, 8.752936, 8.135353, 7.325096, 
    6.461607,
  9.362477, 9.463734, 9.440029, 9.835176, 10.26302, 10.35559, 10.7943, 
    11.41951, 11.74155, 11.84751, 11.76143, 11.71607, 11.13553, 10.22344, 
    8.659704,
  8.695656, 8.449901, 7.894839, 7.623851, 7.91382, 8.273017, 8.725917, 
    9.532962, 9.831021, 9.316591, 8.962348, 8.676834, 8.06601, 7.225804, 
    5.845362,
  7.745787, 7.385979, 6.532128, 5.638867, 5.17563, 5.312193, 5.952312, 
    6.681969, 5.852228, 4.433482, 4.475496, 5.452068, 4.765945, 4.064925, 
    3.359379,
  2.730413, 4.298683, 4.452045, 6.290372, 6.833196, 6.636867, 8.539001, 
    9.283224, 8.920192, 7.171221, 8.035291, 8.92959, 8.18732, 7.723514, 
    7.607666,
  4.852492, 5.539942, 5.751392, 6.126348, 4.997643, 5.675241, 7.74816, 
    7.965709, 7.489945, 6.486352, 6.510343, 8.239676, 8.470304, 5.994435, 
    6.23617,
  7.478673, 6.252262, 5.831138, 5.713232, 4.794509, 4.870783, 7.029787, 
    6.773781, 5.414629, 5.624399, 6.198441, 6.811258, 7.305794, 7.550668, 
    6.175549,
  9.200929, 8.515507, 7.408032, 5.999131, 6.067992, 4.882903, 4.283884, 
    5.16574, 6.669788, 7.36276, 7.033288, 6.536077, 6.507965, 6.739386, 
    5.75983,
  10.21765, 9.162952, 7.95601, 6.241696, 6.041399, 5.712588, 4.481283, 
    2.848784, 4.439811, 5.795312, 7.51135, 7.447412, 6.749879, 6.244253, 
    5.848955,
  10.70724, 9.855535, 8.617102, 6.838993, 5.672985, 5.112078, 4.484664, 
    3.893818, 4.069847, 5.112128, 5.90446, 8.513177, 8.45834, 7.750915, 
    6.644266,
  10.69885, 10.30833, 9.058816, 5.969345, 6.84469, 4.891295, 3.90883, 
    4.625544, 6.074009, 7.38951, 8.170013, 8.576854, 8.77139, 8.739826, 
    8.261137,
  8.795982, 8.002669, 7.107451, 9.702911, 7.618424, 4.334849, 3.221849, 
    4.033188, 5.177459, 6.051948, 6.589668, 6.957914, 7.165312, 7.642409, 
    7.707292,
  8.148254, 8.37419, 11.77126, 12.32016, 7.767972, 4.243204, 3.340025, 
    4.170277, 5.036476, 5.578979, 5.758654, 5.902825, 5.982474, 6.492385, 
    6.54647,
  10.34008, 10.7223, 12.8397, 12.09335, 7.377153, 4.666506, 4.281938, 
    4.918084, 4.718578, 3.825527, 4.108209, 5.324973, 5.384952, 5.992739, 
    6.072619,
  2.023928, 3.256519, 3.667361, 5.161232, 5.158569, 4.398436, 5.937185, 
    6.433596, 6.398063, 5.082932, 5.166198, 5.826021, 5.516366, 5.21405, 
    5.270184,
  3.166847, 3.83606, 4.603246, 5.483035, 4.362402, 3.823222, 5.559821, 
    6.116671, 6.608421, 6.079669, 5.441498, 6.71223, 7.100056, 5.103991, 
    5.148989,
  4.861131, 4.962968, 5.345423, 5.83863, 4.70127, 3.551538, 4.440444, 
    5.991869, 6.200151, 5.771774, 6.118149, 6.795235, 7.298179, 7.175822, 
    6.022288,
  6.756408, 6.619703, 6.751022, 6.565979, 6.258886, 5.232737, 3.533093, 
    3.842737, 5.264035, 5.784602, 5.816951, 6.017201, 6.348107, 6.534168, 
    5.345121,
  6.755268, 7.083167, 7.726489, 7.699749, 7.188234, 6.805088, 4.581202, 
    3.138113, 3.27585, 3.684333, 4.703134, 5.243156, 5.256104, 5.81257, 
    6.067114,
  8.061091, 9.050199, 9.547561, 9.150732, 8.368183, 8.031854, 8.091585, 
    6.029166, 3.152646, 2.405059, 2.838741, 4.443328, 4.651592, 4.983613, 
    5.633725,
  11.79048, 12.35993, 12.62966, 12.96398, 12.93331, 11.88955, 8.587932, 
    5.930949, 3.718925, 3.321434, 3.943575, 4.029003, 3.835489, 4.26249, 
    5.053755,
  14.26106, 13.83113, 13.11605, 12.12137, 9.659561, 6.984595, 4.841742, 
    3.951305, 4.506318, 5.025992, 5.00833, 4.809124, 4.77358, 5.261751, 
    5.551317,
  13.21972, 12.3126, 10.64938, 8.721289, 6.595242, 5.387743, 5.311005, 
    5.931079, 6.518827, 6.493073, 6.552054, 6.84, 6.600441, 6.406583, 5.865828,
  10.04868, 9.035789, 7.652828, 6.198454, 5.610036, 5.912658, 6.556132, 
    7.657242, 7.044956, 5.603863, 6.329926, 8.364647, 7.545133, 6.93834, 
    6.078799,
  6.699501, 10.02985, 10.77024, 13.8799, 10.94565, 8.231762, 10.85701, 
    11.13067, 10.56882, 8.019631, 7.483054, 8.359339, 7.682897, 6.700788, 
    5.595259,
  9.108404, 10.6878, 12.8321, 14.14556, 11.57475, 10.28595, 12.21335, 
    11.41225, 10.90746, 9.569546, 7.971438, 9.216963, 9.035531, 6.058027, 
    5.371757,
  8.806067, 9.91919, 11.68054, 12.4943, 10.03939, 8.771832, 11.78661, 
    12.80958, 11.93629, 11.3143, 9.941688, 8.800355, 7.957819, 7.051359, 
    5.821899,
  7.575396, 9.172131, 10.39032, 10.70961, 9.904722, 7.073596, 6.504238, 
    10.318, 12.60715, 10.63876, 10.32425, 9.163946, 8.117757, 6.863415, 
    5.276506,
  7.511653, 8.579481, 9.441186, 9.639093, 8.818645, 7.371912, 5.735042, 
    5.232053, 5.06747, 5.369792, 7.609172, 7.194927, 6.354584, 5.43537, 
    4.787763,
  8.245001, 8.684514, 9.33623, 9.825264, 9.878939, 9.097858, 6.941346, 
    6.491057, 4.342207, 3.092962, 3.615374, 5.15697, 5.439825, 5.507167, 
    5.197381,
  5.93326, 6.184446, 6.419726, 6.566968, 6.747757, 7.159425, 6.955881, 
    5.283577, 3.306625, 3.943858, 4.885287, 5.929276, 6.801542, 7.440961, 
    7.615554,
  4.102269, 3.894984, 3.535352, 2.982111, 2.260982, 1.84542, 1.931828, 
    2.914172, 4.525929, 6.013017, 7.30837, 8.498918, 9.773647, 10.74596, 
    10.78892,
  5.320076, 4.987888, 4.688984, 4.301133, 4.352338, 5.328163, 6.081006, 
    6.833988, 7.777022, 8.740318, 10.25389, 11.52255, 12.39547, 12.74073, 
    11.85894,
  8.040432, 7.843603, 7.739113, 6.400361, 7.144625, 8.457851, 8.817469, 
    9.466858, 8.639012, 7.281658, 8.77114, 12.18526, 12.33147, 12.18993, 
    10.9528,
  6.926449, 12.27375, 14.04768, 17.96508, 9.362514, 3.356735, 5.343076, 
    7.448446, 9.015299, 8.289425, 8.311369, 8.829939, 8.247941, 6.688984, 
    5.311761,
  8.596939, 12.1743, 16.25671, 18.50144, 11.39791, 4.98357, 3.913612, 
    7.978913, 9.77195, 10.09135, 8.705906, 10.73315, 10.14178, 6.321767, 
    5.682052,
  9.099792, 11.0954, 14.37413, 17.16403, 12.70991, 6.802546, 5.493988, 
    7.349094, 10.76904, 11.2327, 10.7521, 10.84692, 10.34538, 9.583691, 
    7.940386,
  7.741561, 9.997177, 12.90167, 15.62731, 16.30569, 9.575233, 4.299725, 
    7.817464, 9.917912, 9.139556, 10.34698, 10.02863, 9.514692, 9.456431, 
    9.120317,
  6.010683, 7.303818, 9.979209, 12.3689, 15.63619, 15.48942, 8.922228, 
    5.622292, 5.28204, 5.660793, 8.984491, 9.61538, 9.760948, 10.09733, 
    10.2128,
  5.092283, 5.173232, 6.619413, 8.014247, 11.25803, 14.97628, 14.61213, 
    9.057079, 6.04258, 6.272152, 6.780329, 9.600322, 9.906316, 10.07637, 
    9.809115,
  6.263931, 5.266447, 4.287856, 3.072221, 5.067585, 8.921745, 11.89199, 
    12.16628, 10.36584, 9.853608, 9.269517, 9.802654, 9.842295, 10.21947, 
    10.33379,
  9.07042, 8.788432, 7.91859, 5.14671, 3.100112, 3.38141, 6.022742, 8.545395, 
    9.130862, 8.856745, 9.129297, 9.363003, 9.646588, 10.42999, 10.76287,
  12.21105, 12.98921, 12.61707, 10.6317, 8.688389, 6.734744, 4.574211, 
    5.245054, 6.781189, 7.255335, 7.603944, 8.594125, 9.373068, 9.874765, 
    9.678651,
  8.262482, 7.45354, 7.245455, 8.417222, 10.34507, 11.57305, 9.011393, 
    6.629673, 5.455518, 4.53375, 5.650297, 8.01076, 8.623528, 8.95739, 
    7.847092,
  3.7614, 5.416264, 5.879829, 9.602655, 12.44172, 8.079916, 4.446569, 
    2.795774, 3.231327, 3.23276, 4.533813, 5.333292, 4.998843, 4.228204, 
    3.913955,
  6.048334, 6.485603, 7.018987, 9.420158, 8.987215, 5.381797, 2.881387, 
    3.521544, 3.102229, 4.585931, 5.298749, 6.19052, 5.883113, 3.798962, 
    3.725809,
  6.629481, 6.224563, 6.413977, 8.188482, 7.747436, 4.658936, 2.034494, 
    3.138722, 4.557278, 6.389605, 6.748473, 6.000259, 5.694283, 5.623442, 
    4.990471,
  7.659088, 6.401256, 6.362383, 6.468809, 9.097452, 5.963131, 1.648032, 
    3.71556, 5.145907, 6.342779, 6.41697, 5.752365, 6.066769, 5.996162, 
    5.337361,
  8.782578, 6.66251, 5.545297, 4.44093, 7.604704, 9.118731, 3.160414, 
    4.82861, 4.172633, 4.090621, 5.51255, 5.828027, 6.240751, 6.074116, 
    6.311269,
  9.413311, 7.8647, 5.50071, 3.239861, 4.892034, 8.816462, 5.020744, 5.50523, 
    5.247863, 4.792101, 4.302744, 6.517119, 6.489888, 6.641144, 7.664474,
  9.860023, 9.180005, 7.182028, 3.848681, 2.325056, 5.488831, 6.253259, 
    5.23977, 6.819709, 7.058067, 6.511698, 7.116712, 7.198833, 8.228992, 
    9.9012,
  10.6469, 10.28075, 9.208417, 6.170085, 3.271909, 1.823803, 4.940078, 
    5.555861, 6.402454, 6.952536, 7.14187, 7.724471, 8.128371, 9.602488, 
    11.29666,
  10.63143, 10.24185, 9.453642, 6.605247, 4.818685, 4.099123, 3.379204, 
    4.998713, 5.536707, 5.604992, 6.944857, 8.109056, 8.921733, 10.44555, 
    10.55841,
  11.24035, 11.62121, 9.971588, 7.323823, 3.3014, 5.962692, 4.495204, 
    4.253775, 4.18349, 3.386153, 4.840205, 8.154481, 9.41072, 10.69779, 
    10.29821,
  5.954861, 7.372508, 5.443836, 6.301877, 4.24969, 2.896143, 3.248931, 
    2.206113, 2.902217, 1.342932, 1.352409, 2.735332, 3.69835, 4.085977, 
    3.836759,
  9.082234, 8.806593, 8.151716, 6.308257, 3.429083, 2.451253, 1.833603, 
    2.285528, 1.887809, 0.7843283, 1.379102, 3.229883, 5.193675, 3.861139, 
    3.729956,
  11.37474, 10.23582, 8.60186, 7.049553, 3.740357, 2.025737, 0.9158511, 
    1.341452, 1.466837, 1.237742, 2.514571, 3.913942, 5.348858, 5.920148, 
    5.73176,
  11.59492, 12.17432, 10.35664, 7.977229, 5.625549, 2.839925, 0.8107606, 
    0.9113466, 0.9526374, 2.089209, 3.840278, 4.721329, 5.72604, 6.577114, 
    6.630123,
  11.23475, 12.57381, 11.30675, 8.169507, 6.066802, 4.330575, 2.912696, 
    2.468521, 1.521814, 2.079396, 4.715918, 5.488698, 6.252747, 6.558113, 
    6.623132,
  11.18716, 12.51977, 11.91346, 8.710414, 6.467676, 5.599241, 2.921767, 
    3.727603, 2.809539, 3.416971, 4.150976, 6.275698, 5.920831, 5.761989, 
    7.523404,
  11.46542, 12.69534, 12.12515, 9.752422, 6.572253, 4.026724, 1.64241, 
    2.289578, 3.577638, 5.804459, 6.155358, 6.371515, 6.493234, 8.981426, 
    12.30402,
  11.71815, 13.1515, 12.67315, 11.31354, 7.330547, 2.84264, 1.400873, 
    3.714786, 4.645341, 6.557366, 6.876244, 7.438605, 9.667562, 13.3706, 
    13.91578,
  11.55522, 13.26301, 12.95784, 12.34397, 8.102937, 2.382027, 2.632094, 
    4.387681, 5.687434, 7.004736, 7.700405, 9.947825, 13.05869, 14.11721, 
    12.32745,
  10.3841, 11.9312, 12.47033, 12.80395, 8.852984, 3.893921, 3.938221, 
    5.270272, 5.381377, 5.207002, 7.162687, 12.10789, 13.43116, 12.87607, 
    11.32223,
  4.900963, 5.308014, 4.703533, 6.703769, 8.183158, 4.331439, 2.412306, 
    4.179758, 5.214477, 4.178637, 4.607205, 5.100274, 5.809648, 6.793358, 
    7.069689,
  7.057414, 5.426917, 5.021613, 5.793402, 6.064347, 3.771308, 2.565938, 
    3.662931, 4.894256, 4.381749, 3.938743, 5.43741, 7.576514, 6.191633, 
    7.196302,
  10.53851, 7.996851, 4.904456, 4.545931, 5.000851, 3.978018, 3.125626, 
    3.182744, 3.903961, 3.969655, 4.509861, 6.027673, 8.084514, 9.300667, 
    8.558343,
  11.18979, 10.61083, 8.42439, 5.586777, 6.047787, 4.809714, 2.466869, 
    3.159467, 5.532567, 5.193178, 5.35416, 6.90018, 8.979195, 10.38759, 
    10.0731,
  11.1211, 11.15661, 9.524488, 6.117795, 6.069551, 6.661215, 3.526954, 
    2.066236, 3.222182, 3.721336, 6.313526, 8.463223, 10.09519, 11.28714, 
    11.77997,
  10.80879, 11.38789, 10.42063, 7.451927, 6.334538, 6.41457, 5.76625, 
    4.440547, 4.017562, 4.85898, 5.912575, 9.965575, 11.2414, 12.49363, 
    13.09037,
  10.12915, 11.3519, 11.47967, 9.687855, 6.435893, 5.235565, 5.962829, 
    6.921439, 7.39897, 8.002995, 9.372372, 11.064, 12.38991, 13.16741, 
    13.25343,
  9.120262, 10.65645, 11.62754, 11.34165, 7.913357, 4.93718, 5.625947, 
    6.997928, 7.450372, 9.189251, 10.39232, 11.77244, 12.35902, 12.16436, 
    11.09466,
  8.169032, 9.579942, 10.64473, 11.54723, 9.201951, 5.04329, 5.051394, 
    6.379103, 8.181237, 8.760863, 9.934697, 11.24998, 11.0233, 10.22029, 
    8.876083,
  6.70822, 8.220192, 8.916462, 10.41554, 10.68534, 6.281641, 4.24401, 
    6.009867, 6.619737, 6.060287, 7.436767, 10.08617, 9.59558, 9.066276, 
    8.097672,
  4.15569, 5.220757, 5.832652, 8.278697, 6.893951, 5.3102, 7.052245, 
    8.118551, 8.3042, 6.244497, 6.43747, 6.909864, 4.447735, 2.800673, 
    1.860646,
  5.50771, 4.766739, 6.52172, 8.202251, 5.451418, 4.543163, 7.311135, 
    8.548594, 9.066199, 9.018328, 8.286896, 10.45642, 9.662517, 4.818551, 
    3.481284,
  6.830308, 5.624654, 6.360645, 8.096553, 5.68866, 3.87663, 5.522971, 
    7.877743, 9.081367, 10.27754, 11.14838, 12.71248, 13.39935, 11.71467, 
    8.276373,
  6.234872, 6.495163, 6.910457, 7.722161, 8.006001, 4.835666, 2.848227, 
    6.071673, 10.83496, 10.73334, 10.74005, 11.8617, 13.56396, 14.03915, 
    11.81215,
  5.450272, 5.82921, 5.776482, 5.787095, 7.039165, 7.757727, 4.50403, 
    3.316483, 4.963561, 6.045592, 8.990299, 10.29601, 11.55749, 12.59676, 
    12.67436,
  5.023657, 5.412645, 5.235502, 4.964688, 5.357789, 6.562976, 6.615752, 
    5.263433, 3.36465, 4.198753, 5.383499, 8.500986, 9.271973, 9.795913, 
    10.4387,
  4.707724, 5.248526, 5.508842, 4.834965, 4.626709, 5.153038, 5.286741, 
    5.662423, 5.908147, 6.206519, 6.238449, 6.844602, 7.322115, 7.494636, 
    7.651744,
  4.536314, 4.974341, 5.816924, 5.552305, 4.667476, 4.607123, 4.688547, 
    5.026202, 5.015625, 5.201132, 5.161439, 5.257002, 5.472457, 5.754834, 
    5.782894,
  4.866104, 5.031948, 5.625663, 5.835775, 4.995297, 4.283738, 4.746807, 
    4.552235, 4.203468, 3.906923, 3.898513, 4.001139, 4.154923, 4.624987, 
    4.811815,
  5.565936, 5.375542, 5.541885, 5.801471, 6.177599, 4.870497, 5.301524, 
    5.100564, 3.65181, 2.606859, 2.706017, 3.395961, 3.461683, 4.024002, 
    4.609127,
  4.488751, 6.087145, 5.533736, 7.433467, 6.801384, 5.956373, 8.154728, 
    8.722865, 8.854111, 6.971456, 6.915949, 7.270044, 5.288756, 3.84597, 
    2.041229,
  6.533156, 7.610296, 7.450725, 7.546472, 5.605305, 5.321685, 8.024883, 
    8.439001, 9.11004, 8.287993, 7.384586, 8.113754, 7.475264, 4.172941, 
    3.269105,
  6.977688, 7.961829, 8.195388, 7.943889, 5.915702, 5.24248, 7.329676, 
    8.113153, 8.125317, 8.056179, 8.165917, 8.205976, 7.707887, 6.288254, 
    4.178811,
  7.466661, 8.208101, 8.781422, 8.264216, 8.325502, 6.933171, 5.72655, 
    6.122144, 8.107431, 8.933128, 7.906032, 7.471612, 7.082344, 6.122005, 
    5.141019,
  8.141976, 8.473555, 9.035369, 8.408813, 9.414382, 9.856582, 8.482275, 
    5.897025, 6.188719, 6.343122, 7.704875, 7.33339, 6.632485, 5.517546, 
    5.365922,
  8.628342, 8.975595, 9.466785, 9.126837, 10.795, 12.02234, 12.14174, 
    12.02358, 9.543623, 7.095761, 6.389116, 7.71306, 6.698452, 5.328975, 
    4.305028,
  8.680593, 9.390144, 10.12327, 10.55982, 11.63668, 12.81289, 14.44653, 
    14.34187, 12.54002, 10.41873, 9.01278, 8.465728, 7.381705, 5.892504, 
    4.588767,
  8.857987, 9.610674, 10.49378, 11.22656, 12.44649, 13.58879, 14.83804, 
    15.00222, 13.02052, 10.53973, 9.209797, 9.073251, 8.296965, 6.515563, 
    4.985296,
  9.001642, 9.588625, 10.60221, 11.15771, 12.63092, 14.42981, 15.80052, 
    15.23647, 12.48432, 9.480052, 8.834542, 10.13869, 9.271288, 7.081638, 
    5.42928,
  8.438832, 9.094535, 10.24549, 10.68488, 12.79954, 15.30346, 16.55298, 
    14.65277, 10.13862, 6.464263, 7.552165, 10.57434, 9.018094, 6.990366, 
    5.480607,
  5.593488, 8.06286, 7.353003, 10.02815, 9.664703, 8.488304, 11.71885, 
    12.03023, 9.85885, 6.680262, 6.775606, 7.043602, 6.218967, 6.278816, 
    6.732489,
  8.172467, 8.538612, 9.196442, 10.2011, 8.038859, 8.284203, 12.21061, 
    13.30608, 12.0552, 8.497497, 6.280676, 6.756769, 7.155055, 5.556152, 
    5.909313,
  9.105819, 9.768388, 10.42836, 11.17774, 8.558034, 8.027821, 12.03327, 
    12.72849, 11.12329, 8.781956, 6.567148, 5.809264, 6.811903, 7.622413, 
    6.961539,
  8.965528, 10.04455, 11.28572, 12.16544, 12.30103, 9.669764, 8.60815, 
    11.43507, 13.54197, 9.441135, 6.70147, 5.04102, 5.259702, 6.987663, 
    8.056849,
  8.196916, 9.244289, 10.6824, 11.58403, 13.43045, 14.40753, 11.44786, 
    8.791684, 9.049562, 7.57456, 6.886267, 5.440176, 6.237312, 9.353239, 
    8.910859,
  7.407897, 8.559823, 9.975427, 11.39822, 13.56163, 15.05717, 15.34212, 
    13.34404, 8.886059, 6.991748, 5.594456, 6.578373, 9.016994, 10.57764, 
    8.530391,
  6.538937, 7.634353, 9.026264, 10.9165, 12.68798, 13.7793, 14.85872, 
    14.74787, 12.86884, 9.700654, 8.186818, 8.098665, 10.01342, 10.32489, 
    8.777458,
  5.787495, 6.809218, 8.118066, 9.884195, 11.67432, 12.70376, 13.63718, 
    13.78044, 12.78725, 10.70888, 7.977609, 8.710603, 9.749504, 9.157674, 
    8.061359,
  5.269555, 5.966418, 6.853259, 8.160256, 10.01572, 11.22683, 12.4088, 
    13.0089, 12.94326, 11.55725, 9.557902, 9.103176, 8.690768, 7.166345, 
    5.649909,
  4.977449, 5.340729, 6.205247, 7.293159, 9.122457, 10.01307, 10.69036, 
    11.07357, 9.85561, 7.936159, 7.320745, 8.521041, 7.118302, 5.625388, 
    4.025198,
  4.05439, 5.499039, 5.651557, 8.831993, 8.212473, 6.287442, 8.886549, 
    9.25975, 8.508864, 5.991523, 4.548458, 3.372696, 2.609318, 2.76133, 
    2.321473,
  5.643249, 6.315533, 6.924856, 8.465354, 6.519024, 5.843796, 9.188891, 
    9.960848, 9.774113, 8.122522, 5.549376, 4.816123, 3.481185, 2.288177, 
    1.782069,
  7.10793, 7.606851, 7.857297, 8.224813, 6.102499, 5.582763, 7.926403, 
    8.412895, 8.960748, 9.00797, 8.263024, 6.767416, 5.285684, 3.752728, 
    2.147972,
  7.641052, 8.206672, 8.647191, 8.327172, 8.016385, 6.209985, 5.370532, 
    6.72393, 9.714854, 10.12437, 9.313501, 8.36861, 6.934584, 5.40928, 
    3.621052,
  8.471297, 8.514209, 8.808757, 7.995518, 8.377095, 8.354856, 6.939215, 
    5.029393, 5.855522, 6.799616, 8.34349, 8.235311, 7.533815, 6.459296, 
    5.038871,
  9.421611, 9.02944, 8.87307, 8.359725, 8.910513, 8.904449, 9.017295, 
    8.905935, 7.194924, 6.012856, 5.699669, 7.285141, 6.700143, 6.026933, 
    5.4383,
  10.15445, 9.719569, 9.563461, 9.061027, 9.276185, 9.192432, 9.300815, 
    9.402899, 9.202537, 8.452343, 7.947373, 7.117301, 5.888076, 5.142167, 
    4.486298,
  10.80046, 10.35692, 9.833623, 9.575286, 10.14684, 9.872824, 9.430689, 
    9.196363, 9.071821, 8.736063, 8.310905, 7.046378, 5.461505, 4.314538, 
    3.453932,
  11.57847, 11.30082, 10.58282, 10.18393, 10.61803, 10.48992, 10.08308, 
    9.659781, 9.078125, 8.085342, 8.039546, 7.273574, 5.488567, 4.250993, 
    3.259363,
  12.09172, 11.57831, 10.83687, 10.64499, 10.69644, 10.58293, 10.2215, 
    9.640037, 7.929002, 5.526898, 5.922418, 7.167124, 5.446254, 4.178081, 
    3.46633,
  7.876667, 10.51197, 8.807687, 10.17775, 8.795548, 6.714339, 8.529855, 
    9.469645, 9.228305, 7.822615, 8.514099, 8.636744, 6.99633, 5.515326, 
    4.507407,
  11.35686, 12.06196, 11.50532, 10.1993, 5.83861, 4.948026, 7.908394, 
    8.273156, 7.99271, 8.555492, 9.073599, 10.9148, 10.26999, 6.548621, 
    5.012214,
  11.36891, 11.41677, 11.23619, 10.42671, 6.02451, 4.494877, 6.181764, 
    7.330166, 7.256877, 8.011367, 9.732965, 11.47789, 12.26941, 10.9426, 
    7.218622,
  11.98131, 11.79725, 11.37602, 10.54894, 8.764813, 5.473118, 4.416515, 
    4.996928, 6.140122, 7.414011, 9.207355, 10.81819, 11.92515, 11.2763, 
    8.365538,
  12.21201, 11.6743, 11.30488, 10.36834, 9.421535, 8.048417, 6.095859, 
    4.319929, 4.738457, 5.230673, 8.00718, 10.0831, 11.24082, 11.75906, 
    10.53156,
  12.15128, 11.38709, 10.73851, 10.21424, 9.45735, 9.190211, 8.581426, 
    7.563458, 6.27125, 5.638865, 5.970404, 9.458275, 10.32862, 10.7194, 
    9.964663,
  11.70484, 10.92586, 10.22726, 9.756738, 9.354618, 9.187424, 9.354053, 
    9.626579, 9.429798, 9.054906, 8.720992, 8.838733, 8.521822, 10.48119, 
    9.859196,
  11.24429, 10.45224, 9.626987, 9.235958, 9.175964, 9.312007, 9.186576, 
    9.557216, 10.17597, 10.57995, 9.589372, 8.504317, 11.70327, 12.10366, 
    9.23213,
  10.89376, 9.908236, 8.933686, 8.487325, 8.622918, 8.95496, 9.398642, 
    9.882589, 10.51005, 10.62039, 9.434822, 12.06434, 13.90866, 11.18946, 
    7.548073,
  10.32333, 9.212391, 8.353323, 8.862226, 9.199131, 8.993453, 8.984384, 
    9.182862, 8.47204, 6.977021, 7.921102, 12.17805, 10.95012, 8.179531, 
    5.545743,
  6.471545, 8.354462, 7.033316, 8.322896, 6.837212, 4.690313, 5.833926, 
    5.816845, 5.012103, 4.214959, 5.074752, 5.933212, 6.838181, 7.580469, 
    7.718194,
  9.209978, 8.81733, 8.591742, 7.584839, 4.965464, 4.200938, 5.852379, 
    6.105105, 5.823089, 5.156921, 4.993867, 6.163682, 7.285954, 6.869452, 
    7.424492,
  9.402581, 8.637018, 8.054487, 6.757031, 4.509642, 3.92842, 5.496034, 
    5.151974, 4.958455, 6.046637, 6.677182, 6.199225, 6.840617, 9.146613, 
    8.264415,
  9.526074, 8.771851, 8.060595, 6.571509, 5.373141, 4.288056, 3.694878, 
    4.768753, 6.574939, 8.006137, 8.507703, 7.075112, 5.796536, 7.444214, 
    8.59991,
  9.911901, 8.679172, 7.986476, 6.350246, 5.637116, 5.712099, 4.76186, 
    3.332533, 4.708402, 6.586174, 9.202026, 8.32281, 5.863571, 6.210266, 
    9.682719,
  10.30013, 9.026123, 7.889543, 6.733202, 6.244021, 6.051563, 6.182519, 
    5.311611, 4.439581, 4.981909, 6.236722, 8.791049, 6.647761, 3.911378, 
    5.104253,
  10.49735, 9.531001, 8.390411, 7.412739, 6.818542, 6.319212, 6.40119, 
    6.141756, 6.156184, 6.946125, 8.543134, 9.534191, 8.572868, 7.609184, 
    8.585183,
  11.0606, 10.19154, 9.228089, 8.228224, 7.308575, 6.694461, 6.594733, 
    6.440218, 5.85102, 6.04248, 7.033429, 8.285522, 9.901028, 10.95464, 
    10.80439,
  11.3715, 10.73739, 9.759086, 8.708261, 7.616619, 7.087141, 7.076797, 
    6.9388, 6.374691, 5.542613, 5.470099, 5.744291, 5.992554, 6.365892, 
    6.123429,
  10.95901, 10.48842, 10.15837, 9.588516, 7.976598, 7.287607, 7.783485, 
    7.875065, 6.896825, 5.089215, 4.323542, 5.1778, 4.482603, 4.221744, 
    3.855775,
  8.886944, 11.23397, 9.044133, 8.287483, 4.11628, 2.845541, 3.89294, 
    4.779144, 4.444775, 2.942602, 2.477704, 2.983084, 2.58762, 1.783648, 
    3.506462,
  12.56162, 12.52314, 11.71357, 9.033828, 3.708484, 2.588165, 4.354779, 
    4.866256, 5.002882, 4.213793, 3.619086, 3.956537, 3.215575, 1.888296, 
    2.531859,
  12.64713, 11.96731, 11.21366, 9.674581, 4.89374, 2.714203, 3.548989, 
    5.146468, 5.656065, 5.235523, 5.323958, 5.427471, 4.596286, 3.938587, 
    3.116015,
  13.10595, 12.53059, 11.56991, 10.04478, 7.428977, 4.370364, 2.482666, 
    2.389452, 4.191025, 6.367186, 6.550302, 6.176183, 5.222133, 4.345975, 
    4.154614,
  13.76225, 12.50482, 11.24753, 9.760297, 8.153539, 6.516434, 4.637578, 
    3.064593, 3.296997, 4.299376, 5.708221, 6.362148, 5.457904, 4.326061, 
    5.431409,
  14.37421, 12.31032, 10.68272, 9.351507, 8.254795, 7.351451, 6.544735, 
    6.396448, 4.789531, 3.485084, 3.552557, 5.476594, 5.523129, 4.766326, 
    4.498114,
  14.67574, 12.56475, 10.38744, 8.737782, 8.247668, 7.472528, 6.721631, 
    6.458539, 6.107975, 6.035869, 5.728198, 5.190442, 5.213181, 5.124749, 
    3.406827,
  14.73722, 12.56262, 9.692386, 8.171042, 8.359533, 7.773421, 6.710371, 
    6.434093, 6.810291, 7.352857, 7.357646, 6.488923, 5.256828, 4.586759, 
    4.026456,
  14.7042, 11.99566, 8.381892, 6.735209, 7.277021, 7.52939, 7.24344, 
    7.086017, 7.231136, 7.827792, 8.736023, 8.77392, 7.282205, 5.692508, 
    4.119646,
  13.10729, 10.66675, 6.90357, 5.699414, 6.750176, 7.415307, 7.480627, 
    7.407702, 6.489807, 5.566195, 6.979995, 9.7927, 8.659669, 7.253363, 
    5.335776,
  8.735644, 10.40433, 7.405, 8.908333, 7.258971, 4.754297, 5.262037, 
    5.105028, 5.234237, 4.551244, 4.204492, 3.595767, 2.525035, 1.923848, 
    1.682624,
  12.02994, 10.71605, 8.755972, 8.29305, 5.928795, 5.021801, 6.508492, 
    5.939787, 5.725978, 5.330823, 5.157833, 6.111233, 4.813625, 2.419232, 
    1.363088,
  11.50717, 10.22494, 8.676508, 7.48851, 6.210741, 5.366949, 6.670069, 
    6.156997, 6.170626, 6.580809, 6.639017, 7.100982, 7.643258, 5.689656, 
    2.952108,
  11.46724, 10.40241, 8.786702, 7.396243, 7.685075, 6.057148, 5.018999, 
    4.97524, 6.751382, 7.988094, 8.184909, 7.93961, 8.139157, 8.479893, 
    6.232254,
  11.671, 9.830035, 8.394338, 6.874412, 7.882476, 8.252765, 6.418165, 4.4721, 
    4.927631, 5.918146, 7.597567, 7.983165, 7.549824, 8.042828, 9.345209,
  11.78092, 9.768629, 7.882009, 6.917819, 8.163097, 8.51563, 7.89732, 
    6.130666, 4.361438, 4.902651, 5.124476, 6.967165, 7.32582, 6.98919, 
    7.667581,
  11.10363, 9.64821, 7.662778, 7.101743, 7.970222, 8.271297, 7.969742, 
    7.757124, 7.191893, 7.274165, 7.555294, 7.614722, 7.340298, 7.316772, 
    6.47155,
  10.48746, 9.351181, 7.708759, 7.461562, 8.023391, 8.139438, 7.661125, 
    7.34929, 7.346257, 7.52963, 8.037963, 8.56827, 8.322143, 7.637168, 
    6.725583,
  9.743064, 8.521679, 7.234226, 7.126099, 7.326521, 8.153402, 8.045933, 
    7.668775, 7.249084, 7.237519, 7.523588, 8.164729, 8.592405, 8.148974, 
    6.795491,
  8.514677, 7.10219, 6.431729, 6.778811, 7.510027, 8.326104, 8.19096, 
    8.02453, 6.719144, 4.883125, 5.325156, 7.469192, 7.969676, 8.308082, 
    7.116552,
  4.895745, 6.619992, 6.856863, 8.606681, 7.089405, 6.22975, 8.424249, 
    9.214838, 10.15913, 8.027913, 7.632987, 7.492661, 4.841619, 2.975988, 
    1.980081,
  7.04321, 6.728611, 8.133873, 8.431044, 5.698224, 5.186177, 8.077895, 
    8.893528, 10.03564, 10.38888, 9.247399, 9.462342, 7.881031, 4.11244, 
    2.656034,
  7.801558, 7.639779, 8.250813, 8.168321, 6.354294, 4.878517, 6.645821, 
    6.815059, 7.716058, 9.852848, 11.24086, 11.10969, 8.99471, 7.607923, 
    4.33582,
  7.982491, 7.794591, 7.729874, 7.09739, 7.726202, 5.639592, 4.536414, 
    6.004493, 8.43394, 8.878334, 9.625147, 10.59704, 10.09329, 8.291101, 
    6.243723,
  8.100611, 7.727673, 7.345656, 6.141373, 6.795271, 6.728909, 5.673229, 
    4.120403, 5.228672, 6.410332, 8.001139, 8.639421, 9.446372, 8.976495, 
    7.156723,
  8.595629, 8.020708, 7.385828, 6.71996, 7.242015, 6.355734, 6.798099, 
    6.344288, 5.431177, 5.034659, 4.890437, 6.919161, 7.861528, 9.302105, 
    7.718401,
  9.144824, 8.435331, 7.563068, 7.229502, 7.492734, 6.901594, 7.385154, 
    7.515635, 7.119051, 6.513867, 6.299146, 6.182454, 6.536656, 7.795881, 
    9.870391,
  9.701232, 9.103498, 8.285733, 7.628793, 8.133608, 7.963315, 7.711889, 
    7.26615, 6.722321, 5.88064, 5.554147, 5.234489, 5.438498, 6.872614, 
    9.477059,
  10.03615, 9.359219, 8.551148, 7.107073, 7.465578, 8.574001, 8.705123, 
    8.193077, 6.726885, 5.235723, 4.611546, 4.463654, 4.291228, 5.830158, 
    8.056696,
  9.924532, 9.0684, 8.654039, 7.557353, 7.867325, 9.289444, 9.185931, 
    8.41406, 5.934314, 3.373283, 3.433856, 3.979964, 3.195274, 4.600444, 
    7.048283,
  6.943941, 9.45974, 8.265703, 10.31325, 8.576743, 6.090276, 7.888267, 
    6.427649, 4.57967, 3.08284, 3.894108, 6.299458, 6.90445, 5.709614, 
    3.366674,
  11.0456, 10.24206, 9.575996, 8.902641, 5.487318, 5.145285, 8.006429, 
    6.663682, 5.074492, 3.547152, 2.490617, 5.209481, 7.092147, 5.008973, 
    4.21649,
  12.27701, 11.29246, 9.815669, 7.320168, 5.241891, 4.045168, 6.065686, 
    6.59969, 5.958681, 4.488541, 3.029002, 2.84817, 5.563114, 6.504182, 
    5.657956,
  12.43608, 11.44182, 9.524088, 6.375175, 5.756579, 4.331347, 3.903757, 
    4.169518, 4.98556, 5.510732, 4.630979, 2.324742, 3.166033, 5.74716, 
    6.535131,
  12.23096, 11.18995, 9.054278, 5.294122, 4.680415, 4.274677, 5.317487, 
    4.064439, 3.699226, 4.144971, 5.40584, 4.124956, 1.940109, 4.026444, 
    7.023339,
  12.24718, 11.26856, 8.990433, 5.431946, 4.181664, 2.432795, 3.850813, 
    5.787661, 4.302445, 3.391382, 4.134708, 5.304479, 3.131647, 2.454464, 
    5.850441,
  12.32659, 11.57489, 9.564316, 6.566139, 4.096422, 2.284784, 2.507053, 
    3.959004, 4.323151, 4.345227, 5.589909, 6.10781, 4.268013, 1.927874, 
    4.621753,
  12.41912, 12.02537, 10.58258, 8.057496, 5.811327, 3.580263, 4.092482, 
    4.430723, 4.392878, 3.934225, 5.113002, 6.407794, 4.866919, 1.954516, 
    4.152006,
  12.21307, 11.9075, 10.90142, 8.502921, 6.533328, 4.927823, 4.691582, 
    4.814841, 4.196366, 3.594224, 4.854043, 6.482013, 5.073493, 2.026823, 
    3.65446,
  11.67108, 11.33895, 11.38265, 10.04674, 8.083236, 6.342342, 4.495068, 
    4.129875, 3.698045, 2.963322, 4.07108, 6.478892, 4.651683, 1.874066, 
    3.597867,
  6.235058, 7.310905, 6.322994, 8.187187, 8.648587, 7.031651, 6.724217, 
    8.183472, 8.773394, 6.102549, 3.747475, 2.805973, 3.668271, 3.562579, 
    3.068126,
  11.10532, 9.420387, 8.206757, 8.221266, 6.00788, 3.621668, 3.828984, 
    8.286696, 9.937363, 7.573442, 4.176386, 3.173924, 4.217481, 3.361649, 
    3.121175,
  12.1377, 11.25266, 10.23205, 7.492525, 4.116024, 2.899827, 5.704461, 
    10.42644, 11.13022, 7.786112, 4.788429, 3.158921, 4.824502, 4.890994, 
    3.702994,
  12.37492, 11.48817, 9.805054, 6.103563, 5.480298, 3.901076, 5.759575, 
    8.637135, 7.95506, 6.062168, 4.377696, 3.07881, 4.804433, 4.750496, 
    3.881448,
  12.4789, 11.39116, 9.183859, 4.951307, 4.113454, 3.886304, 6.623165, 
    6.529733, 4.252656, 4.134331, 4.129059, 3.395496, 4.693578, 4.883433, 
    3.901873,
  12.59293, 11.82133, 9.792376, 6.07578, 3.671856, 3.42732, 5.193328, 
    8.966925, 6.062925, 4.971031, 3.578078, 4.069685, 4.409632, 5.009241, 
    4.361728,
  12.58959, 12.60588, 11.40217, 8.448568, 5.102826, 4.122042, 5.187008, 
    8.251019, 8.061745, 7.293776, 5.937484, 5.035676, 4.607326, 4.907867, 
    5.497127,
  12.26801, 13.1051, 12.99335, 11.47725, 8.531289, 7.438081, 9.511434, 
    9.879354, 8.728963, 7.552365, 6.387392, 5.674956, 5.0727, 5.228567, 
    5.906221,
  10.8958, 12.09889, 12.28382, 12.00942, 11.01879, 10.00051, 9.82144, 
    9.092261, 7.788741, 6.813842, 6.331918, 6.249318, 5.655723, 5.537612, 
    5.319595,
  7.923519, 9.590316, 10.43369, 10.57411, 10.16294, 9.341429, 8.353385, 
    7.968114, 5.99972, 4.429864, 4.850245, 6.5389, 5.900251, 5.826276, 
    5.253123,
  5.1829, 5.561595, 5.411452, 9.047524, 10.58254, 7.267153, 7.084814, 
    6.204123, 5.429786, 3.580496, 7.186674, 8.852221, 8.070936, 6.214831, 
    4.179255,
  8.722227, 7.078452, 7.125458, 9.215744, 7.991054, 5.863528, 3.530707, 
    6.452127, 6.007947, 6.294598, 8.150336, 9.639408, 9.191658, 5.131351, 
    3.750796,
  8.848653, 8.399355, 9.380424, 9.748466, 8.230823, 6.312757, 6.295262, 
    6.664488, 7.484307, 8.322175, 9.513011, 8.73648, 7.533957, 6.433614, 
    4.592819,
  8.241585, 8.027596, 8.960412, 9.949958, 10.99567, 8.207698, 5.804432, 
    8.760221, 10.0094, 8.827831, 8.263949, 6.25483, 5.898805, 5.947799, 
    5.101046,
  7.662321, 7.184024, 7.90002, 8.65556, 10.38734, 10.48519, 7.373779, 
    5.015408, 5.36179, 5.069868, 5.053619, 4.01431, 4.741367, 5.384888, 
    5.963712,
  7.518757, 6.884744, 7.232691, 8.182008, 9.273029, 9.709245, 9.204886, 
    6.734554, 3.100603, 2.420022, 2.155753, 3.516844, 4.203985, 5.267178, 
    5.899731,
  7.827893, 7.661288, 7.449476, 7.648603, 8.08998, 8.003314, 7.721817, 
    6.689058, 4.945522, 3.094506, 3.157206, 3.894297, 4.18539, 5.918336, 
    6.327093,
  7.482641, 8.09177, 7.933784, 7.506267, 7.501739, 7.397828, 6.797164, 
    5.63697, 4.443689, 4.313993, 4.155162, 3.732513, 4.876189, 6.324624, 
    6.301627,
  6.563354, 7.403, 7.353052, 7.014168, 6.762234, 7.141145, 6.969525, 6.33912, 
    5.495527, 4.935384, 4.18118, 4.774114, 5.900884, 5.866412, 4.83525,
  4.857814, 5.868044, 6.107352, 6.404912, 6.380527, 7.046111, 7.408241, 
    7.521377, 6.060873, 4.63544, 4.822312, 6.437052, 5.897691, 5.106303, 
    3.478458,
  2.536837, 2.958106, 4.334505, 9.825414, 11.70893, 10.22899, 13.24324, 
    11.39979, 7.549855, 4.713545, 4.337368, 5.279008, 7.018151, 9.472269, 
    9.110688,
  3.229115, 3.598338, 5.543311, 9.347168, 8.411202, 8.729715, 13.83974, 
    14.43968, 11.86727, 10.85622, 8.453197, 10.08899, 12.92663, 9.077103, 
    8.139907,
  4.057111, 4.604789, 7.34861, 9.231394, 8.07529, 6.820337, 11.07372, 
    15.35523, 16.2486, 15.96297, 15.96411, 16.46889, 14.10901, 11.26587, 
    8.613203,
  4.889728, 5.19251, 6.982358, 8.666441, 10.29051, 7.635639, 5.681685, 
    10.98351, 16.86323, 15.65166, 14.31086, 14.11877, 13.32953, 11.21517, 
    8.115137,
  5.734564, 5.52082, 6.299926, 7.032328, 8.972573, 9.904155, 7.028701, 
    5.327661, 7.248883, 8.35474, 10.46104, 10.58777, 10.40375, 10.22351, 
    8.837163,
  6.8184, 6.286572, 6.621483, 7.042805, 7.57173, 7.785417, 7.521772, 
    4.981303, 2.792164, 3.452803, 4.513565, 7.202951, 7.655639, 7.496092, 
    7.389325,
  7.329075, 7.403028, 7.612999, 7.606234, 7.196562, 6.355442, 4.981586, 
    4.136737, 3.685344, 3.382688, 3.345666, 4.284927, 4.954238, 4.900643, 
    5.132349,
  6.683897, 7.548498, 8.226637, 8.490789, 7.984772, 7.063184, 5.225284, 
    3.615729, 2.915323, 2.117281, 2.170902, 2.665555, 3.056998, 3.500978, 
    3.899722,
  5.809824, 6.717765, 7.467141, 8.34832, 8.727608, 8.294522, 6.685644, 
    3.893833, 3.244611, 3.503972, 3.74928, 3.758724, 3.685271, 3.51516, 
    3.494512,
  4.129466, 5.069407, 6.225089, 7.44302, 9.139974, 10.61569, 9.898829, 
    7.044361, 2.9695, 1.421431, 2.033344, 2.881837, 3.231454, 3.169063, 
    3.064118,
  2.970157, 5.221294, 5.853499, 8.900648, 8.718477, 7.359936, 10.8585, 
    12.64284, 13.04369, 9.837622, 5.904964, 3.931762, 3.623036, 4.55709, 
    4.276134,
  5.15133, 5.40995, 6.540275, 8.229134, 6.661727, 6.478346, 10.01539, 
    11.44299, 12.33919, 12.71007, 9.819398, 4.320601, 3.939177, 3.556392, 
    4.049606,
  6.427784, 6.814312, 7.30449, 7.571208, 6.080245, 5.741426, 9.006838, 
    9.229313, 9.37404, 11.88493, 13.99657, 8.974895, 3.864969, 5.305141, 
    4.96908,
  6.495484, 6.813895, 7.22067, 6.925536, 7.429324, 6.044141, 6.121865, 
    7.86651, 9.985341, 10.48855, 12.73729, 13.71039, 5.59446, 6.285543, 
    6.042218,
  6.154293, 6.505091, 7.011546, 6.204633, 7.556765, 8.111288, 6.76138, 
    5.248099, 6.122297, 6.78222, 9.676294, 11.55824, 9.80412, 6.003584, 
    6.861887,
  5.62944, 6.411924, 7.180392, 7.277688, 8.032253, 8.673295, 8.376656, 
    7.515834, 5.955343, 4.635493, 5.027839, 8.875822, 9.428161, 6.764446, 
    6.939703,
  5.645917, 6.850403, 7.557318, 7.343288, 7.730765, 8.591178, 9.377913, 
    9.209237, 7.160835, 5.044592, 4.840361, 6.573628, 7.729285, 6.839534, 
    6.109477,
  6.65989, 7.709863, 7.695125, 6.881804, 7.189578, 8.283884, 9.183159, 
    8.906203, 6.871612, 4.447245, 3.475779, 4.514612, 5.870365, 6.069664, 
    5.009976,
  8.240059, 8.058333, 6.434917, 5.593608, 6.124615, 7.222778, 9.189708, 
    9.310699, 7.496634, 4.291308, 2.433782, 2.89624, 4.270532, 4.774659, 
    4.343502,
  8.684676, 6.694614, 4.588715, 5.026778, 5.020778, 6.410869, 8.89188, 
    9.454918, 6.872541, 3.188787, 1.442309, 1.670923, 3.032173, 3.743527, 
    3.560758,
  6.173068, 8.79357, 7.616009, 8.803557, 7.916435, 6.851763, 9.055634, 
    8.361834, 7.268116, 6.066, 6.571813, 5.267171, 5.077105, 6.519026, 
    5.646587,
  9.396643, 9.272593, 8.396758, 8.051475, 5.948367, 5.80017, 7.934275, 
    7.105532, 7.054904, 6.604858, 6.535429, 5.593249, 5.162566, 5.511367, 
    5.884459,
  9.301391, 8.736396, 7.901792, 7.400696, 5.44284, 5.181551, 5.818656, 
    5.901892, 5.258086, 6.349253, 7.552786, 5.904832, 4.244686, 6.127415, 
    5.903894,
  8.295926, 7.937299, 8.06512, 7.742296, 8.04239, 4.933505, 3.149324, 
    4.60916, 5.694965, 7.177332, 7.795706, 6.266413, 3.839393, 4.485296, 
    4.575484,
  7.345765, 7.233984, 8.147886, 8.205422, 8.558248, 5.239046, 3.374207, 
    2.480207, 4.113805, 5.425122, 7.320457, 7.012825, 4.12765, 3.217965, 
    2.985607,
  7.594079, 7.174893, 8.195435, 8.777102, 7.870663, 5.077738, 3.82998, 
    2.800831, 4.317341, 4.537219, 4.58999, 7.070213, 5.245402, 4.725518, 
    4.424105,
  7.663872, 7.69953, 8.42201, 7.922668, 5.873648, 4.800638, 3.667835, 
    4.647137, 5.38702, 5.459397, 5.720231, 6.827714, 6.6297, 4.885561, 
    4.794777,
  7.266692, 7.128932, 7.022614, 5.966534, 5.21353, 3.992558, 4.378045, 
    4.775366, 4.664177, 4.396028, 4.841867, 6.396028, 6.80131, 5.594558, 
    4.659537,
  5.835435, 4.894664, 4.317317, 4.069386, 3.76658, 3.720051, 5.888488, 
    6.018336, 4.646605, 3.480286, 4.167299, 6.180474, 6.686422, 5.492376, 
    4.3649,
  3.599001, 2.847361, 3.03203, 2.766639, 2.281169, 3.680812, 6.456867, 
    6.609024, 4.043956, 2.173705, 2.860455, 5.512537, 6.466372, 5.191157, 
    4.188747,
  3.563003, 6.094785, 6.079535, 7.614806, 6.803026, 4.910349, 5.467535, 
    3.63619, 2.995455, 2.16147, 1.957035, 3.973509, 4.665431, 5.032099, 
    5.697142,
  5.401812, 6.192305, 6.491637, 6.5568, 4.610427, 3.905142, 4.872532, 
    3.758277, 3.413956, 1.449859, 2.705306, 5.44357, 6.101377, 4.330386, 
    5.148079,
  5.089451, 5.517632, 6.016797, 5.730915, 4.406908, 3.524543, 4.164386, 
    4.291429, 2.527256, 1.908211, 4.41643, 6.385076, 6.991206, 6.972763, 
    5.503929,
  4.240266, 4.861509, 5.301196, 5.286963, 5.722898, 4.197026, 2.998682, 
    3.620545, 3.499388, 3.282726, 4.62465, 6.775009, 8.157595, 7.769153, 
    5.413695,
  3.685334, 3.800832, 4.332503, 4.270061, 5.265198, 5.792593, 4.049283, 
    2.31338, 3.200153, 3.654185, 5.512053, 7.482768, 8.788976, 8.344231, 
    6.335365,
  3.421201, 3.839141, 4.013798, 3.588358, 4.313582, 5.323528, 5.585064, 
    4.451697, 4.399086, 3.965338, 4.54741, 7.310833, 8.864064, 8.568578, 
    4.921539,
  3.257926, 4.00542, 3.719097, 3.365191, 3.617946, 4.699202, 6.560009, 
    6.674537, 5.875875, 5.377859, 6.271244, 7.415389, 8.665141, 7.29654, 
    3.559526,
  3.036424, 4.083029, 3.698086, 3.349074, 3.246821, 3.92893, 6.734908, 
    6.996368, 6.293121, 5.728782, 6.647537, 7.255539, 7.609257, 5.821623, 
    3.32221,
  3.642215, 4.509266, 4.171875, 3.633387, 2.939147, 3.36152, 6.903512, 
    7.873394, 6.866573, 6.339449, 6.980642, 7.138917, 6.771601, 5.117175, 
    3.891386,
  3.769895, 4.283587, 4.880465, 3.614789, 3.493482, 3.047562, 6.711556, 
    7.816908, 6.349886, 4.593127, 5.222155, 7.092693, 6.649602, 6.013025, 
    5.246552,
  2.371078, 3.733912, 4.346071, 5.979611, 5.337307, 4.309295, 5.382964, 
    5.942914, 5.225554, 3.554037, 3.07011, 3.302032, 3.33289, 3.462025, 
    4.054954,
  3.917878, 4.501789, 5.557296, 6.41396, 4.505875, 3.722063, 5.009765, 
    5.812255, 6.099825, 5.113291, 4.16575, 4.988424, 5.520399, 4.223361, 
    4.967197,
  4.242023, 5.838534, 6.597249, 6.389236, 4.047633, 3.093813, 4.26631, 
    4.965369, 4.955429, 5.49917, 5.700253, 6.180643, 7.262824, 8.366376, 
    7.709289,
  4.545258, 5.907902, 7.204455, 6.739122, 4.945326, 3.443665, 3.109119, 
    5.222024, 6.671719, 6.836798, 6.864665, 6.974563, 7.787764, 8.846927, 
    8.425855,
  4.289573, 5.857435, 7.693781, 7.009717, 5.448933, 3.882871, 2.821952, 
    3.55083, 5.533477, 6.467901, 8.031562, 7.936364, 8.308175, 8.684485, 
    9.080086,
  3.686425, 5.239581, 7.319218, 6.631006, 5.386438, 3.506557, 3.885471, 
    5.77241, 6.341922, 5.97755, 5.901773, 8.259695, 9.08991, 9.288792, 
    9.543114,
  3.030431, 4.75871, 6.603245, 5.492865, 5.258877, 3.381004, 5.39825, 
    7.580389, 7.783244, 7.797855, 8.439961, 9.138906, 9.669049, 9.507186, 
    9.983739,
  2.403503, 4.291116, 6.033339, 4.94511, 5.023834, 4.08532, 5.707613, 
    6.990878, 7.3129, 8.106365, 9.067719, 10.34414, 10.49541, 9.98974, 9.16099,
  2.360564, 3.596058, 4.608272, 4.738157, 5.196245, 4.808421, 6.260164, 
    7.137155, 7.133554, 7.88319, 9.65163, 11.53139, 11.79491, 11.28159, 
    10.22308,
  2.090449, 3.308274, 3.556895, 4.269173, 4.771663, 5.414181, 6.38715, 
    6.674364, 5.79044, 5.315067, 7.449688, 11.95324, 13.40151, 13.76692, 
    12.58605,
  3.025732, 4.388057, 4.43587, 6.158565, 6.068995, 4.720215, 4.802524, 
    4.532814, 5.112736, 4.784064, 5.313695, 5.677998, 4.857633, 3.786477, 
    3.463165,
  4.054319, 4.579547, 4.951855, 5.696508, 4.016025, 3.455048, 4.934821, 
    5.565336, 6.414419, 6.040285, 5.830867, 6.936924, 6.629276, 4.466505, 
    4.107855,
  3.99631, 4.03504, 4.583746, 5.262984, 3.924638, 3.005702, 4.733467, 
    5.968775, 5.798495, 7.031874, 7.954549, 8.154655, 7.660956, 7.082125, 
    5.832409,
  3.661305, 3.742556, 3.936947, 4.838178, 4.750074, 3.335555, 3.275144, 
    5.989672, 8.782182, 9.599318, 9.838425, 9.715942, 9.049025, 8.442188, 
    7.372284,
  2.903829, 3.336305, 2.903111, 3.840565, 4.125857, 4.823015, 3.981586, 
    3.894682, 6.202528, 8.322724, 11.12763, 11.12986, 10.17741, 9.283412, 
    8.885693,
  2.476856, 3.387957, 2.498515, 3.010643, 3.188865, 4.432409, 5.05173, 
    5.183895, 5.384218, 6.671309, 7.959475, 11.70122, 11.19615, 9.183167, 
    8.111078,
  2.800711, 3.902774, 2.481814, 2.693743, 2.802465, 3.996251, 5.169369, 
    7.271048, 9.004292, 10.6216, 12.13321, 12.79301, 11.90475, 9.684036, 
    6.712837,
  3.588108, 4.856163, 2.984513, 2.700518, 2.822259, 3.745628, 4.608013, 
    6.637572, 8.961761, 10.8448, 12.60944, 13.827, 13.20813, 11.39629, 7.36959,
  4.168775, 6.163915, 3.951787, 2.822731, 2.927082, 3.573743, 4.373223, 
    6.526174, 8.928462, 10.49414, 12.39498, 14.24655, 14.25113, 12.59605, 
    8.742614,
  4.523974, 7.502968, 5.530034, 3.4005, 3.168113, 3.824087, 4.088194, 
    5.99678, 6.928421, 6.311909, 8.069599, 13.61909, 14.85162, 13.68565, 
    9.90566,
  2.738188, 3.195323, 2.331898, 2.141834, 2.071858, 2.730647, 3.888318, 
    4.679889, 4.888758, 4.447911, 4.918025, 5.197059, 5.182657, 4.410162, 
    3.612194,
  4.304594, 3.149089, 2.736037, 2.306079, 2.02647, 2.770616, 4.15032, 
    5.094849, 5.765584, 5.457147, 5.227314, 6.845007, 6.220621, 4.234007, 
    4.082566,
  6.127538, 4.767773, 3.867992, 3.143522, 2.51317, 2.602523, 4.20604, 
    4.601324, 4.700732, 5.757039, 6.756876, 7.681459, 7.97559, 7.355861, 
    5.40379,
  6.994355, 6.244806, 4.939726, 4.32364, 3.976697, 3.063454, 3.225912, 
    4.915287, 6.313287, 6.49879, 7.287323, 8.606178, 9.019066, 8.890355, 
    6.45751,
  6.908587, 6.626612, 5.950408, 5.707299, 5.521937, 4.976511, 4.513053, 
    3.766098, 5.466892, 6.490436, 8.257224, 9.559442, 9.756136, 9.6872, 
    8.87927,
  5.915751, 5.97374, 5.949955, 6.388134, 6.758645, 6.782135, 7.02362, 
    7.633542, 7.616799, 7.325448, 6.668839, 9.744223, 10.40841, 10.3769, 
    10.03035,
  5.342714, 5.599019, 5.865134, 6.249621, 7.039826, 7.477186, 8.35737, 
    9.454986, 10.16669, 9.855739, 9.629251, 9.840277, 10.13583, 10.90863, 
    10.48546,
  4.460449, 5.200938, 5.940015, 6.589127, 7.645421, 8.503873, 9.437004, 
    9.72862, 9.990608, 9.831098, 9.603707, 9.250658, 9.825191, 11.19703, 
    10.85965,
  3.786772, 5.119436, 6.315629, 7.29679, 8.493991, 9.194346, 9.826562, 
    9.837547, 9.260954, 8.654163, 8.120065, 8.453798, 9.667005, 10.95417, 
    10.74997,
  3.904502, 5.437088, 7.099237, 8.511621, 9.24276, 9.741487, 9.275127, 
    8.365623, 6.901584, 5.247199, 5.190687, 7.463872, 8.782491, 10.63332, 
    10.37282,
  6.013389, 8.476631, 7.351713, 8.51762, 6.855712, 5.114303, 6.876598, 
    6.935609, 6.517407, 4.859675, 4.435352, 4.0676, 3.253159, 2.73225, 
    2.248256,
  8.568719, 9.08208, 8.472037, 7.805806, 4.487135, 3.876714, 6.387099, 
    7.153781, 7.877005, 6.5421, 5.551101, 5.671068, 5.181068, 3.572262, 
    3.096732,
  7.852459, 7.505268, 7.199591, 6.214971, 4.626069, 3.23074, 5.07914, 
    6.984967, 8.363592, 8.600634, 8.405166, 7.8968, 7.777942, 7.727328, 
    5.552744,
  5.96244, 5.009434, 5.342766, 5.415858, 6.192833, 5.753703, 3.891165, 
    5.152351, 7.305247, 8.017715, 8.602505, 9.020227, 9.16131, 9.501766, 
    8.203864,
  3.876865, 3.456378, 4.320911, 5.027984, 5.84309, 7.285038, 7.286936, 
    5.138441, 5.826635, 5.72197, 8.052115, 9.754173, 10.08442, 10.29293, 
    10.88973,
  3.196308, 3.539397, 4.200294, 5.128266, 6.357978, 7.887444, 9.266786, 
    9.952949, 8.456707, 7.391763, 7.327, 11.00797, 11.57, 11.21959, 11.22333,
  4.225796, 4.666916, 5.160499, 6.192811, 7.671842, 8.869426, 9.181289, 
    9.094543, 9.279971, 9.877098, 10.22251, 10.3864, 10.09944, 9.653162, 
    9.858718,
  5.150714, 5.214503, 6.114443, 7.501764, 9.21305, 9.017083, 8.210098, 
    8.424918, 8.883891, 8.749671, 8.093721, 7.947623, 7.876478, 7.913996, 
    8.179378,
  5.163098, 5.643075, 6.726101, 8.787704, 9.19486, 7.99867, 8.028957, 
    8.364094, 7.886926, 6.864199, 6.963026, 8.432964, 8.74322, 8.49611, 
    8.041276,
  5.039153, 5.961956, 7.953098, 9.680032, 8.387856, 7.625395, 7.243993, 
    7.254753, 6.565723, 5.668063, 7.163712, 9.870276, 8.610125, 7.34805, 
    6.512046,
  3.305653, 5.05236, 4.749658, 5.65913, 4.55979, 2.855164, 3.221373, 
    3.820244, 4.592036, 4.082492, 4.708769, 5.142577, 4.018793, 2.747689, 
    1.807998,
  5.370856, 5.805265, 5.716407, 4.880281, 2.806634, 2.581192, 3.941802, 
    4.850187, 6.1299, 6.362546, 6.244666, 7.18303, 6.952245, 4.258943, 
    3.233962,
  5.647549, 5.66663, 5.803102, 5.134507, 3.800853, 3.322821, 4.679233, 
    5.675139, 7.177587, 8.327398, 8.357808, 8.067593, 7.184076, 6.497176, 
    5.167887,
  5.083356, 5.431839, 6.173975, 6.68945, 6.695181, 5.039047, 4.006532, 
    4.684326, 6.635523, 7.582614, 7.436769, 6.415322, 5.003994, 4.699182, 
    3.708219,
  4.80651, 5.644809, 6.70753, 7.682263, 8.15573, 7.645029, 5.869618, 
    4.376675, 4.826858, 4.615758, 5.474711, 5.071968, 4.83328, 5.198473, 
    5.050274,
  4.839664, 6.023246, 6.896644, 7.765746, 8.088558, 8.147244, 7.48588, 
    5.480357, 3.655433, 3.656464, 3.532534, 4.402289, 4.405489, 4.604714, 
    5.087126,
  4.8221, 6.096343, 6.850808, 7.426653, 7.42874, 7.520417, 7.458199, 7.11461, 
    6.196774, 5.146813, 4.727796, 4.992702, 5.498092, 5.894016, 6.301614,
  4.645754, 5.75221, 6.432049, 6.950935, 7.135554, 7.225884, 7.115294, 
    6.729686, 6.40091, 6.179178, 6.139582, 6.434231, 7.024384, 7.411829, 
    7.509202,
  4.204123, 5.031547, 5.441083, 5.499443, 5.934556, 6.409206, 7.316316, 
    8.281115, 8.026512, 7.776756, 7.298759, 7.522512, 7.727033, 7.697262, 
    7.452783,
  3.708739, 4.266459, 4.275677, 4.348142, 4.803854, 6.135077, 7.940722, 
    8.551419, 7.861922, 6.113187, 6.496526, 8.237024, 7.675691, 7.386023, 
    6.761296,
  4.875767, 6.705606, 6.537482, 7.55252, 6.533724, 6.108841, 8.098567, 
    8.424724, 8.388987, 6.78152, 6.470866, 6.488017, 5.118647, 3.497231, 
    2.079739,
  6.399883, 7.047006, 7.97135, 7.884996, 5.497053, 5.254477, 7.859136, 
    8.599193, 8.935516, 8.340075, 7.392375, 8.327549, 7.177797, 4.139429, 
    3.219544,
  5.467566, 6.085273, 7.439791, 7.546352, 5.718279, 4.397051, 6.344525, 
    6.502168, 6.904, 8.013335, 8.331477, 8.805305, 8.33415, 7.086587, 5.038761,
  4.452192, 5.11412, 5.969694, 6.674297, 6.805243, 4.620148, 4.045507, 
    5.434025, 7.35536, 8.057937, 7.619534, 7.400272, 7.049309, 7.538748, 
    7.064248,
  3.758631, 4.320332, 4.77523, 4.965263, 5.68956, 6.403242, 4.952189, 
    3.693469, 4.965292, 5.747033, 7.083959, 6.831014, 5.671044, 5.122609, 
    5.897942,
  3.615899, 4.018199, 4.114876, 4.358974, 5.254575, 5.418808, 6.127492, 
    5.891308, 5.175908, 4.88869, 4.385783, 6.197071, 5.981263, 4.305419, 
    3.439274,
  3.771403, 4.067837, 3.753364, 3.725339, 4.726554, 4.862643, 6.060981, 
    7.145675, 7.411194, 7.125555, 6.551996, 6.369521, 6.328894, 5.095326, 
    3.143737,
  4.581096, 4.603666, 3.908756, 3.731379, 4.941289, 4.72991, 5.873226, 
    6.527219, 6.892147, 6.764876, 6.553473, 6.676883, 6.616212, 5.718946, 
    4.019164,
  5.490472, 4.828572, 3.811445, 3.949807, 5.051956, 4.468046, 5.750257, 
    6.887949, 7.484652, 7.699315, 7.136168, 7.119806, 6.631167, 5.915597, 
    4.389459,
  5.958161, 4.983526, 4.665157, 4.949707, 5.093077, 4.384046, 5.23619, 
    6.147687, 6.28604, 5.252695, 5.480661, 6.862422, 6.145115, 5.778605, 
    4.578306,
  3.733363, 4.818157, 4.773763, 6.63829, 6.693108, 5.663667, 6.9752, 
    6.861635, 5.952466, 4.597996, 4.801058, 5.300307, 5.261598, 5.284022, 
    5.06571,
  6.08744, 6.563444, 6.861777, 7.862533, 5.887674, 5.116416, 7.163911, 
    7.008981, 6.771699, 5.679075, 4.752075, 5.388735, 5.263871, 4.190175, 
    4.704868,
  6.682047, 7.530148, 8.000917, 8.54917, 6.139652, 4.847384, 6.356835, 
    6.545888, 6.584699, 6.230224, 5.868853, 5.617915, 5.185561, 4.962646, 
    4.579366,
  6.727475, 7.677144, 8.464869, 8.757381, 8.636769, 6.419299, 4.825965, 
    4.793852, 5.972663, 6.573406, 6.139932, 5.564846, 5.178267, 4.966974, 
    3.858509,
  6.786624, 7.345289, 8.593844, 8.773232, 9.256378, 8.872663, 7.155409, 
    4.565448, 4.462164, 4.955766, 5.86217, 5.431387, 5.068362, 5.011137, 
    3.837514,
  6.502294, 7.126547, 7.825589, 8.268197, 9.097902, 9.414172, 9.657617, 
    8.592108, 5.475013, 4.502418, 3.98997, 4.8932, 4.903728, 4.93289, 4.103454,
  6.150062, 6.50293, 6.896884, 7.690698, 8.936546, 8.892022, 9.205179, 
    6.764947, 7.341681, 6.154454, 5.140564, 4.553709, 4.565471, 4.774426, 
    4.313322,
  5.553789, 5.940236, 6.619542, 8.137755, 8.524985, 8.346354, 7.32806, 
    6.48807, 7.43379, 5.543706, 4.356491, 3.935123, 4.090319, 4.676242, 
    4.239934,
  4.696618, 5.410566, 6.786629, 8.151649, 7.950442, 7.73058, 6.89434, 
    6.718284, 5.805406, 3.824841, 2.630821, 3.139716, 3.676525, 4.214162, 
    4.149008,
  4.38447, 5.455795, 7.541557, 8.526927, 8.115942, 6.992361, 6.652779, 
    6.77158, 4.11432, 2.157371, 2.122083, 3.533182, 3.633554, 3.708782, 
    3.747138,
  5.030089, 7.635671, 7.774604, 10.16202, 10.01009, 8.572594, 10.86845, 
    10.97728, 9.396014, 7.053697, 7.363592, 7.344725, 5.811811, 3.813246, 
    2.795027,
  7.179128, 8.078465, 8.931463, 9.841882, 6.359516, 5.585195, 8.913718, 
    9.682654, 8.411827, 6.694199, 6.963369, 8.794448, 8.247634, 4.122684, 
    2.425483,
  6.769485, 7.245292, 8.044274, 7.966333, 5.40472, 4.11964, 6.780901, 
    8.304779, 8.118555, 7.917843, 7.982601, 8.424147, 9.420941, 6.100912, 
    2.553313,
  6.029788, 6.27525, 6.884396, 7.050125, 7.019897, 4.972373, 4.347962, 
    5.977822, 8.107106, 8.682367, 7.693871, 9.538383, 9.383108, 5.823813, 
    2.460596,
  5.614812, 5.643327, 6.310213, 6.823706, 7.658781, 7.600739, 5.617341, 
    4.456107, 5.672052, 5.423202, 8.131817, 10.04403, 8.530675, 5.766497, 
    3.405086,
  5.228539, 5.468494, 5.989915, 6.563969, 7.540301, 8.445187, 8.299379, 
    6.596585, 4.143837, 4.844713, 5.369114, 7.912459, 6.415279, 4.89425, 
    3.782947,
  4.640005, 5.395734, 6.09379, 6.556326, 7.050149, 7.668324, 7.590041, 
    7.990458, 7.497478, 6.609601, 6.041046, 5.059379, 4.339145, 4.120275, 
    3.628431,
  4.345908, 5.788942, 6.424648, 6.901217, 7.124533, 7.08396, 7.113769, 
    7.010029, 6.098073, 5.056329, 3.863583, 2.301799, 2.396056, 3.376446, 
    3.723785,
  5.022658, 6.325091, 6.892479, 7.312233, 7.097653, 6.876248, 6.789196, 
    6.274011, 5.341651, 4.298645, 2.88321, 1.495157, 1.229415, 2.423969, 
    3.933072,
  5.708282, 6.846152, 7.434091, 7.155832, 6.825329, 6.731318, 6.509235, 
    5.873706, 4.755548, 3.118381, 2.399424, 2.0544, 1.678319, 2.092455, 
    3.303101,
  5.130231, 7.97189, 7.380106, 8.137959, 7.02, 7.058786, 9.851826, 10.30065, 
    9.893672, 7.351881, 5.913312, 5.738534, 5.653381, 6.334366, 6.491904,
  6.671037, 8.119482, 9.211805, 8.937675, 5.343812, 5.437273, 9.05003, 
    10.38978, 11.4205, 11.14455, 8.47059, 5.321965, 5.931521, 5.792884, 
    5.864251,
  6.04506, 7.510176, 9.145753, 9.350968, 6.437632, 4.493182, 6.71223, 
    8.250513, 10.11246, 12.84807, 12.35769, 6.914056, 3.972776, 8.457891, 
    7.19174,
  5.623781, 6.838472, 8.212439, 9.230722, 9.02387, 5.906301, 4.191795, 
    6.835984, 11.44586, 13.91238, 13.76886, 10.74642, 7.299641, 8.897576, 
    7.395188,
  5.577715, 6.394, 7.376988, 8.084586, 8.928741, 9.048074, 6.503115, 
    4.732984, 6.546689, 8.491673, 12.19593, 12.8794, 10.93448, 9.594442, 
    8.342923,
  5.586995, 6.118831, 6.90625, 7.619422, 8.20715, 8.478246, 8.57516, 
    7.349016, 4.870141, 4.953914, 6.590765, 10.25544, 10.54532, 10.02623, 
    9.189168,
  5.528462, 6.231934, 6.597878, 7.208973, 7.519813, 8.00359, 7.949673, 
    7.77517, 7.150998, 6.61497, 6.678656, 7.538726, 8.028619, 7.974745, 
    7.636354,
  5.695416, 6.45804, 6.630692, 7.017244, 7.170176, 7.829386, 7.878131, 
    7.148263, 6.340178, 5.477149, 5.013443, 4.689868, 4.811741, 4.91616, 
    5.443671,
  5.851654, 6.319296, 6.284603, 6.393928, 6.793781, 7.454206, 8.002739, 
    7.619155, 6.492896, 5.395409, 4.258661, 3.262049, 2.886217, 2.824627, 
    3.217334,
  5.671166, 5.976677, 6.202265, 6.33356, 6.718823, 7.415916, 8.103863, 
    7.523731, 5.616453, 3.505224, 2.718977, 1.938182, 1.407222, 1.79409, 
    2.236202,
  4.5341, 7.208234, 7.183094, 9.025417, 7.364671, 4.923476, 6.31092, 
    6.987154, 6.652081, 6.365095, 7.472379, 8.156704, 6.66619, 5.30304, 
    4.857944,
  7.90764, 8.444409, 8.224494, 8.366421, 5.391117, 4.624192, 6.623808, 
    7.545889, 7.631449, 7.965908, 8.704692, 9.50306, 8.325081, 5.775013, 
    5.772517,
  8.891034, 9.696839, 9.377176, 7.691337, 5.036367, 4.440203, 6.653004, 
    6.970291, 6.771475, 9.429745, 11.91769, 11.23562, 6.940794, 7.423498, 
    7.194506,
  9.034582, 9.953355, 9.726498, 8.296339, 6.434102, 4.459606, 4.641893, 
    6.052167, 8.274145, 10.52204, 12.74341, 13.47892, 7.947633, 5.122508, 
    7.576662,
  8.988174, 9.687409, 9.697818, 8.563704, 7.294005, 6.249416, 4.8921, 
    3.661159, 5.160456, 7.287263, 10.91483, 13.2899, 12.27116, 6.947807, 
    8.018232,
  8.920984, 9.702572, 9.612028, 8.897494, 7.537151, 6.957684, 6.224391, 
    4.617913, 3.615482, 4.623783, 6.536967, 10.62537, 12.41144, 11.61342, 
    8.599333,
  8.690052, 9.501457, 9.50941, 8.773963, 7.3983, 7.115569, 6.560286, 
    5.827798, 5.552845, 6.787846, 8.301649, 9.181737, 9.785406, 9.806163, 
    8.714789,
  8.508806, 9.449655, 9.370408, 8.584322, 7.44838, 7.079735, 6.463001, 
    5.379172, 4.887107, 6.227301, 7.327082, 8.350623, 8.851926, 8.620948, 
    7.414143,
  7.995178, 8.794388, 8.418941, 7.709094, 7.104321, 6.913029, 6.84712, 
    6.326967, 5.588855, 6.072583, 6.998302, 7.681789, 8.399003, 9.029461, 
    8.241613,
  7.199745, 7.747315, 7.449536, 7.515871, 7.561385, 7.526321, 6.877102, 
    6.530638, 5.282618, 4.018661, 4.443635, 6.715124, 7.926753, 9.002356, 
    9.516198,
  3.730302, 4.757496, 4.283849, 6.54504, 5.674945, 4.359392, 5.461015, 
    5.621859, 4.954644, 4.515191, 5.289076, 5.68545, 6.020315, 6.175553, 
    4.479539,
  5.512421, 4.653363, 4.671892, 5.845747, 4.497976, 4.227147, 6.070745, 
    6.685225, 6.490904, 5.757453, 5.376036, 6.751932, 6.377026, 4.509506, 
    3.988867,
  6.354535, 4.867756, 4.957156, 5.250803, 4.400102, 3.824648, 5.705739, 
    6.244249, 5.780544, 6.374912, 6.847538, 7.216319, 6.259607, 5.17572, 
    4.111101,
  6.371094, 4.969573, 4.821468, 5.219038, 5.473013, 4.045871, 3.852405, 
    6.071121, 8.869392, 9.078269, 8.339254, 7.738572, 6.632608, 4.128643, 
    4.760738,
  6.001711, 4.762549, 4.462961, 4.734615, 5.367531, 6.015384, 4.499115, 
    3.941221, 5.854828, 7.241122, 9.204986, 8.4298, 7.072002, 4.204996, 
    4.176437,
  5.518331, 4.827742, 4.385458, 4.736217, 5.378916, 6.267951, 6.260535, 
    5.754508, 5.353556, 6.244409, 6.979955, 8.99021, 7.252298, 6.168036, 
    3.35749,
  5.123486, 4.898668, 4.323793, 4.507054, 5.123462, 6.104509, 6.70234, 
    7.84323, 8.693141, 10.03622, 11.70744, 11.05829, 7.343699, 6.263604, 
    5.300653,
  5.039083, 4.905472, 4.07759, 4.181283, 4.977445, 6.048189, 6.718656, 
    7.778111, 9.077327, 10.59054, 12.74727, 13.3128, 9.608854, 6.420431, 
    6.477169,
  5.283459, 4.812665, 3.812891, 3.586328, 4.436064, 5.83083, 6.958193, 
    8.574875, 9.92205, 11.28725, 13.38912, 14.8712, 13.44241, 7.139483, 
    6.712635,
  5.649896, 4.695731, 3.456741, 3.153157, 4.240089, 5.701818, 6.992538, 
    8.349966, 8.466695, 7.468859, 9.785301, 14.87202, 15.55883, 12.39998, 
    5.989007,
  5.667792, 9.861054, 5.697868, 3.104542, 2.36109, 3.979468, 6.8244, 
    7.898607, 6.477004, 4.958436, 5.332841, 6.280069, 7.224287, 8.088655, 
    5.932729,
  11.67533, 11.32482, 6.350156, 2.995663, 2.749736, 4.372473, 7.461507, 
    8.766291, 8.179262, 5.785412, 5.17468, 6.527222, 6.717733, 6.270746, 
    6.587019,
  12.53416, 9.883056, 6.434718, 4.091528, 3.587837, 4.055944, 7.573145, 
    8.454372, 7.46233, 6.894836, 6.042554, 5.821153, 5.268262, 6.696894, 
    7.308098,
  10.39168, 7.902397, 5.667711, 4.709157, 5.290252, 4.405002, 5.536764, 
    8.09978, 10.55021, 10.16939, 7.481745, 5.154327, 3.715286, 4.030991, 
    6.641348,
  7.962404, 6.172441, 4.731473, 4.511693, 5.531099, 7.28868, 6.503393, 
    5.396419, 7.16376, 8.446284, 8.985214, 5.200574, 2.89623, 1.86402, 
    5.601025,
  6.151836, 5.152081, 4.385026, 4.685975, 5.993515, 7.656744, 8.803703, 
    8.043556, 6.84602, 7.557886, 6.678556, 5.256769, 2.852347, 3.171849, 
    3.686076,
  5.032794, 4.477167, 4.126705, 4.454681, 5.866613, 7.782741, 9.328668, 
    10.36868, 11.55599, 13.01055, 12.29922, 7.372914, 2.61134, 3.820991, 
    3.589998,
  4.622408, 4.125598, 3.684206, 4.035153, 5.723168, 7.959082, 9.299107, 
    9.952121, 11.34257, 13.21475, 13.5335, 10.11238, 4.013336, 3.812772, 
    3.810479,
  4.447771, 4.030855, 3.008189, 2.989768, 4.814374, 6.957612, 8.948109, 
    10.54067, 11.63918, 12.80642, 13.56216, 12.00141, 6.369207, 2.167198, 
    3.937557,
  4.531761, 3.798745, 2.137663, 2.17039, 3.916909, 5.965846, 8.164853, 
    9.566855, 9.235287, 7.738825, 9.378585, 12.53969, 9.800224, 3.036503, 
    3.279793,
  6.25659, 8.118848, 4.933078, 4.458513, 3.524905, 3.371009, 4.695673, 
    5.515089, 5.627332, 5.105206, 5.537499, 5.675204, 5.384732, 5.535329, 
    6.525201,
  8.9073, 7.533527, 5.791392, 4.925858, 3.780656, 3.760345, 5.394253, 
    6.444239, 7.2481, 5.844193, 5.091877, 5.253482, 4.545837, 3.870698, 
    6.395146,
  7.439638, 6.691087, 6.541468, 6.106449, 4.752018, 3.848323, 6.076629, 
    6.536151, 6.589988, 6.811646, 5.611067, 4.201701, 3.350573, 5.155102, 
    7.427216,
  5.473611, 5.666299, 6.128872, 6.549283, 6.662408, 4.916386, 4.353755, 
    6.406621, 9.172581, 9.305777, 7.055681, 4.628247, 3.990281, 6.183089, 
    7.431144,
  3.967417, 4.657702, 5.67417, 6.537142, 7.159868, 7.44057, 5.472585, 
    4.419492, 6.042244, 7.061566, 7.179514, 5.467759, 4.592757, 6.835124, 
    8.971112,
  2.714394, 3.382589, 4.817349, 6.395445, 7.05924, 7.464474, 7.460787, 
    6.542287, 5.724651, 6.143534, 5.130737, 5.606728, 5.49366, 6.967605, 
    8.911205,
  2.174047, 2.012469, 3.381052, 5.323845, 6.572313, 7.234046, 7.831201, 
    8.232909, 9.292439, 10.16656, 9.026736, 6.331042, 5.422461, 6.734677, 
    8.324047,
  2.434264, 1.52505, 1.735249, 3.649235, 5.648885, 6.837098, 7.522994, 
    7.448736, 8.687477, 10.36223, 10.16249, 7.826664, 5.495412, 6.44179, 
    7.878479,
  3.117228, 2.342123, 1.3238, 1.975197, 3.811753, 5.451927, 7.019375, 
    8.167681, 9.331037, 10.41964, 10.70622, 9.475924, 6.775011, 5.855091, 
    7.072472,
  4.174861, 3.473053, 2.395637, 1.808032, 2.39321, 3.733289, 5.80163, 
    7.382049, 7.61621, 6.626839, 7.347349, 10.03318, 8.213078, 5.677425, 
    5.73209,
  2.125355, 3.230781, 3.920905, 5.232425, 4.216912, 3.0979, 3.911947, 
    4.335047, 4.473898, 4.09817, 4.49556, 4.143344, 3.48183, 3.491853, 
    4.173389,
  2.335519, 2.452754, 4.403342, 5.753551, 3.955862, 3.45841, 4.878748, 
    5.377684, 5.758962, 5.669002, 5.217556, 4.886556, 4.190024, 3.172047, 
    3.635123,
  2.356157, 2.99439, 4.473212, 5.684221, 4.348107, 3.38418, 5.133716, 
    5.227089, 5.205696, 6.563324, 7.117524, 5.765512, 4.698816, 4.968129, 
    5.169871,
  2.311784, 2.447637, 3.878616, 4.957731, 5.363504, 3.886806, 3.659201, 
    4.990788, 7.124381, 8.476176, 8.643362, 7.148588, 5.623805, 5.472908, 
    5.662197,
  2.863462, 1.760832, 3.167349, 4.447094, 5.187026, 5.62389, 4.497539, 
    3.623218, 4.965151, 6.758267, 8.81552, 8.037886, 6.502162, 6.221369, 
    6.695365,
  4.000605, 1.6463, 2.338907, 3.9185, 4.7776, 5.516834, 5.857795, 5.269103, 
    4.904205, 5.527175, 6.218498, 8.096229, 7.38201, 6.978347, 6.62879,
  5.073925, 2.08899, 1.34218, 2.781772, 4.262426, 5.386111, 6.206185, 
    6.637655, 7.279332, 8.699484, 9.734892, 9.334773, 8.16348, 7.712053, 
    5.363132,
  5.895756, 2.894951, 1.439346, 1.639037, 3.82917, 5.263067, 6.245866, 
    6.497888, 7.114894, 8.901579, 10.34737, 10.32066, 9.206928, 8.409966, 
    5.216876,
  6.10259, 3.702544, 3.23012, 1.769029, 2.284001, 4.704071, 6.318354, 
    7.232965, 8.04355, 9.377636, 10.80651, 11.22301, 10.04259, 8.60707, 
    6.182712,
  5.716303, 3.224146, 3.627928, 2.126851, 1.583851, 3.693083, 5.596639, 
    7.133415, 7.203068, 6.342897, 8.138962, 11.47777, 10.6041, 8.655468, 
    6.758204,
  2.32044, 2.451323, 3.148127, 4.333826, 3.655387, 3.040212, 4.079263, 
    4.615154, 4.572065, 4.217107, 5.243555, 6.120952, 5.166992, 3.5121, 
    2.571395,
  3.151183, 1.901879, 3.472002, 4.537079, 3.402725, 3.193837, 4.612344, 
    5.216824, 5.028565, 5.130198, 5.881779, 7.469724, 6.693174, 3.503727, 
    2.907155,
  3.675436, 1.780593, 3.28487, 4.465673, 3.66827, 3.10533, 4.628488, 
    4.628105, 4.028625, 5.563977, 7.486359, 8.418316, 7.667295, 5.834404, 
    3.894398,
  5.085946, 2.241526, 3.227722, 4.174583, 4.66134, 3.694804, 3.50003, 
    4.455936, 5.764039, 7.007546, 8.354527, 9.375966, 8.687266, 6.486197, 
    4.385917,
  5.367703, 2.648633, 2.940411, 3.719416, 4.440848, 5.160017, 4.337641, 
    3.387756, 4.495162, 6.014611, 8.725371, 10.15076, 9.232433, 6.986163, 
    5.489381,
  5.09637, 2.789088, 2.731289, 3.493684, 4.304685, 5.178081, 5.406551, 
    4.95525, 4.549355, 5.261946, 6.561006, 10.25466, 9.183216, 7.057552, 
    5.443787,
  4.28381, 2.80754, 2.385401, 2.875907, 4.108588, 5.205338, 5.837595, 
    6.510145, 7.229435, 8.204713, 9.682145, 10.93926, 9.019213, 7.066102, 
    3.698006,
  3.731261, 2.893796, 2.262275, 2.622382, 4.171014, 5.24008, 5.90797, 
    6.461941, 7.29931, 8.623436, 10.4288, 11.42694, 8.773616, 6.140867, 
    2.673638,
  3.392414, 2.755495, 2.016932, 2.48623, 3.936367, 4.84507, 5.580381, 
    6.904922, 8.177739, 9.327064, 11.1384, 11.53825, 8.334092, 5.03837, 
    3.350187,
  3.09043, 3.409309, 3.313175, 3.564689, 4.057131, 4.115321, 4.480311, 
    6.029708, 6.787979, 6.073861, 8.429012, 10.88835, 7.793093, 4.670509, 
    3.621922,
  1.686502, 2.671853, 3.132903, 4.162825, 3.817627, 3.217187, 4.238862, 
    4.33733, 3.386983, 3.03137, 3.569714, 4.104347, 4.433851, 4.082917, 
    3.649033,
  1.996451, 3.301788, 4.103914, 4.582201, 3.509156, 3.253317, 4.618452, 
    4.633446, 4.223876, 3.96082, 4.044078, 4.991011, 5.639368, 3.676991, 
    3.676436,
  2.430599, 4.335355, 4.833547, 5.03932, 3.833424, 3.497406, 4.59195, 
    4.568292, 4.131503, 4.633475, 5.128411, 6.012105, 6.417562, 5.847018, 
    4.469928,
  3.586803, 5.496468, 6.12054, 6.037518, 5.85377, 4.809917, 4.039382, 
    4.257452, 4.434238, 4.756636, 5.749473, 6.815754, 7.071306, 6.517533, 
    4.832188,
  5.165553, 6.688153, 7.074007, 6.860399, 6.840921, 6.668228, 5.808839, 
    4.17771, 4.141627, 4.528879, 6.388993, 7.523285, 7.654592, 6.815706, 
    5.555126,
  6.512869, 7.781093, 7.483294, 7.00736, 7.112057, 7.374579, 7.552542, 
    7.697651, 6.332778, 5.289978, 5.228106, 7.863252, 7.933676, 6.608442, 
    5.728251,
  7.564444, 8.368467, 8.082239, 7.452971, 7.756711, 7.88951, 8.124894, 
    7.937937, 7.855288, 7.441941, 7.128023, 7.953763, 7.854709, 6.25037, 
    5.379701,
  8.185482, 8.998043, 8.527885, 8.118625, 8.431298, 8.199074, 7.406078, 
    5.947275, 5.047627, 5.693646, 6.563309, 7.862001, 7.692132, 6.17195, 
    4.977793,
  8.660125, 9.116856, 8.293658, 8.12087, 8.589615, 7.915985, 6.262572, 
    3.967452, 3.483189, 4.021519, 6.062839, 7.919308, 7.698816, 5.915386, 
    4.452616,
  8.956388, 8.707696, 8.301989, 8.477445, 8.521746, 7.135811, 4.800728, 
    3.029349, 2.760858, 3.604353, 5.941803, 8.776789, 7.16144, 5.590346, 
    4.369606,
  3.685625, 5.285949, 5.268285, 7.122995, 6.911534, 6.360572, 8.136237, 
    8.160883, 7.560526, 5.268076, 4.257013, 3.57776, 2.411347, 1.571649, 
    1.954484,
  5.569728, 6.97339, 7.682635, 8.502868, 6.249047, 6.38006, 9.557194, 
    9.477779, 9.007659, 7.517758, 5.788081, 5.465451, 4.197347, 1.793829, 
    1.23737,
  6.543299, 8.160968, 8.546268, 8.590949, 5.932563, 5.309897, 7.608562, 
    9.28642, 9.581846, 9.260018, 8.411839, 7.333502, 5.897762, 3.792913, 
    1.632691,
  7.495176, 7.905906, 7.766999, 7.285642, 6.596558, 4.726171, 4.300434, 
    5.447289, 6.958665, 8.800714, 10.04432, 9.011317, 7.168379, 5.153117, 
    2.72073,
  7.696424, 7.338217, 7.35524, 6.887368, 6.314342, 5.466665, 4.490171, 
    3.183173, 3.708358, 4.271169, 7.902797, 10.09885, 8.573471, 6.523205, 
    4.119341,
  7.323919, 7.182924, 7.511789, 7.486452, 7.170782, 6.87372, 6.400703, 
    6.625677, 5.530377, 3.687713, 4.366167, 9.199336, 9.459157, 7.168706, 
    5.008132,
  7.220008, 7.463075, 7.875081, 7.809114, 8.043963, 7.252795, 7.00747, 
    6.74099, 6.129685, 6.177238, 6.46285, 8.662836, 9.570481, 7.690621, 
    5.732122,
  7.581317, 7.802509, 8.038416, 8.383687, 8.983486, 8.033381, 6.173992, 
    5.225332, 3.771315, 4.054854, 6.553249, 8.654038, 9.764725, 8.320726, 
    6.362292,
  7.903901, 7.978513, 8.069279, 8.697926, 9.518082, 8.657922, 6.195903, 
    4.502319, 3.772699, 2.455355, 5.942789, 8.802641, 9.626422, 8.520728, 
    6.353417,
  8.046511, 8.179563, 8.413036, 9.828894, 11.23152, 10.32402, 7.35103, 
    3.710347, 5.140011, 3.669491, 4.991907, 9.299438, 9.560884, 8.4501, 
    6.527164,
  3.096293, 3.590151, 3.20848, 3.2931, 2.716099, 2.312509, 3.460509, 
    4.388363, 5.676505, 4.747056, 4.524399, 4.52176, 3.562664, 2.277769, 
    1.19646,
  4.879488, 4.912076, 5.276945, 5.246616, 3.377175, 2.941529, 3.727559, 
    3.902761, 5.661718, 6.600757, 5.565567, 5.851747, 5.481241, 2.870084, 
    1.184529,
  5.767039, 6.588507, 6.365032, 5.861879, 4.521881, 3.665358, 3.859909, 
    3.185731, 3.970684, 6.675342, 7.669799, 7.203724, 6.552987, 4.928332, 
    1.962119,
  6.844092, 7.309398, 6.975689, 5.261694, 4.955563, 4.602893, 3.209767, 
    2.580037, 2.578793, 4.051567, 7.2169, 8.050968, 7.610229, 5.930317, 
    2.746667,
  7.471982, 7.08797, 5.930838, 3.398798, 3.247629, 4.747588, 5.550014, 
    3.917758, 3.10026, 2.443743, 5.047457, 8.139416, 8.67029, 7.418575, 
    2.78936,
  7.696493, 6.711078, 4.421993, 3.218823, 3.889377, 4.905604, 6.116199, 
    7.890728, 5.814229, 3.229293, 3.1053, 7.705014, 9.637033, 7.887837, 
    3.423576,
  7.674646, 6.446871, 4.397213, 4.019292, 5.431439, 6.307226, 5.577468, 
    6.146436, 7.246934, 6.045132, 4.240312, 7.360747, 10.5637, 8.493814, 
    4.920674,
  7.735454, 6.749447, 5.128788, 5.423997, 6.871085, 6.547233, 4.802649, 
    4.55101, 7.487153, 7.751974, 5.181873, 7.706087, 11.52739, 9.044061, 
    5.910525,
  7.93223, 7.105894, 5.81003, 6.429674, 6.684157, 4.63504, 3.627173, 
    4.213782, 8.4547, 8.226187, 6.007089, 9.377515, 12.30903, 9.170903, 
    5.849138,
  7.884896, 7.527554, 6.61494, 7.021079, 6.534059, 4.568059, 3.853379, 
    6.724612, 8.493989, 5.420573, 5.815576, 11.309, 11.5772, 8.507961, 
    5.001537,
  4.159345, 6.325218, 5.957095, 7.427367, 6.433836, 4.455762, 3.95559, 
    1.892727, 1.578059, 2.837821, 3.648263, 4.268304, 3.978059, 3.201962, 
    2.710592,
  4.730346, 5.545348, 6.039441, 7.055407, 5.572299, 5.549993, 7.172269, 
    4.494085, 2.642428, 3.492016, 4.090087, 5.333202, 5.245983, 3.153945, 
    2.781082,
  4.229478, 4.55782, 4.73049, 5.067556, 4.449118, 4.468998, 6.631915, 
    7.221831, 4.773491, 4.245323, 5.10422, 5.959546, 5.533237, 4.374974, 
    3.470243,
  5.168655, 4.786511, 4.046414, 2.208763, 1.976752, 2.312826, 3.132133, 
    5.205232, 5.353807, 4.888149, 5.529302, 6.095989, 5.870831, 4.660262, 
    3.72726,
  5.668899, 4.279093, 2.807587, 0.9932436, 1.385936, 1.999543, 2.549249, 
    4.445842, 4.15548, 3.837293, 6.033859, 6.366197, 6.087077, 5.493418, 
    3.27793,
  5.828238, 4.028072, 1.778339, 1.964105, 2.331012, 1.218768, 1.845479, 
    5.475215, 5.434137, 4.963375, 5.308749, 7.054428, 6.712421, 5.293649, 
    2.924316,
  5.646012, 4.042382, 2.354627, 1.92731, 3.276054, 1.843713, 1.815829, 
    4.257364, 7.059637, 7.423542, 7.633446, 7.485266, 6.790578, 4.931045, 
    3.256842,
  5.701716, 4.69024, 3.373283, 1.955613, 2.623174, 2.99686, 3.340391, 
    6.462562, 7.77048, 7.906186, 7.778518, 7.685353, 6.451999, 4.632257, 
    3.135002,
  6.205777, 5.720439, 4.044811, 2.775805, 2.649217, 4.218502, 5.455263, 
    7.273319, 8.10288, 8.027838, 7.358194, 7.618468, 6.273396, 4.749903, 
    2.235447,
  6.157211, 6.260479, 5.096251, 4.581851, 4.672826, 5.423843, 6.929907, 
    8.564953, 7.646699, 5.79556, 5.740782, 7.837328, 5.664469, 3.430748, 
    1.640009,
  1.394028, 2.083516, 3.014941, 4.637712, 4.312543, 4.02556, 4.90425, 
    3.837334, 2.406496, 1.918372, 1.299302, 3.113515, 3.828556, 4.516675, 
    5.796059,
  2.608343, 3.842876, 4.401703, 4.575889, 2.827214, 3.162676, 5.147645, 
    4.694308, 2.830601, 2.467092, 1.963205, 3.403646, 4.546727, 3.911058, 
    4.851293,
  3.793535, 4.496412, 4.230668, 3.920918, 2.689933, 2.46387, 4.395526, 
    5.795762, 3.948998, 3.738288, 3.429211, 3.960479, 4.946692, 5.202467, 
    4.916282,
  5.081136, 5.251092, 4.787831, 3.519516, 2.434941, 1.945242, 2.669945, 
    4.166281, 3.952251, 4.304899, 4.634457, 4.347811, 4.648079, 5.082017, 
    5.259093,
  5.654206, 5.278713, 4.037992, 2.720253, 1.819125, 1.674675, 3.118108, 
    3.999199, 3.454686, 3.628148, 5.431635, 4.995209, 4.703285, 5.086613, 
    5.594097,
  5.918975, 4.600214, 2.873176, 1.662995, 3.456665, 2.840858, 1.858785, 
    3.768227, 5.173142, 5.301276, 5.046317, 5.912242, 5.216738, 5.333846, 
    5.630382,
  5.694351, 3.33107, 1.969775, 0.9521869, 3.878565, 3.796572, 1.722267, 
    2.236254, 7.20991, 8.370402, 7.965342, 6.767531, 5.880556, 5.489139, 
    6.127582,
  5.362928, 3.553457, 1.488382, 0.920377, 3.068726, 3.387201, 1.744073, 
    4.705158, 8.399533, 8.766111, 8.083426, 7.107541, 5.391289, 5.198467, 
    5.823062,
  5.801253, 4.994324, 3.111048, 2.920056, 3.867157, 2.804313, 3.014788, 
    6.847915, 9.228541, 8.696585, 8.173409, 6.911164, 5.181894, 5.137623, 
    4.971517,
  6.107138, 6.109696, 5.319133, 4.87165, 4.408502, 4.180257, 6.441334, 
    9.377023, 8.391569, 6.039836, 6.087082, 6.822254, 4.990656, 4.892703, 
    3.631882,
  1.307616, 1.548155, 1.726615, 2.506641, 2.750428, 3.06134, 4.525491, 
    4.85814, 4.541306, 3.441434, 2.57088, 3.212562, 4.333379, 5.54595, 
    6.226547,
  2.254493, 2.856043, 3.735721, 4.055254, 3.031619, 3.551241, 5.437887, 
    4.842277, 4.160699, 2.99284, 2.32666, 3.702293, 5.462535, 5.389098, 
    4.685044,
  2.546785, 3.880473, 4.429324, 4.663224, 3.526691, 3.023165, 3.794998, 
    3.314914, 3.091317, 2.417681, 2.165053, 4.768085, 6.676984, 6.819794, 
    3.704982,
  4.194179, 5.625927, 5.665509, 4.802332, 3.932188, 2.695571, 1.603502, 
    2.080487, 2.688578, 2.204077, 2.571255, 5.237847, 6.557226, 4.718843, 
    4.642734,
  5.732358, 5.635215, 4.572282, 2.48978, 2.403485, 2.523633, 2.525719, 
    2.269091, 2.114722, 1.974374, 3.23862, 5.15098, 4.424369, 4.185804, 
    6.344978,
  5.466173, 4.028532, 1.967994, 1.248399, 1.442161, 1.087922, 2.104369, 
    2.461188, 2.57864, 2.484668, 2.677894, 3.687773, 4.020281, 6.710579, 
    8.427588,
  4.584195, 2.688093, 1.462678, 1.449944, 1.688515, 1.800887, 1.564142, 
    3.800876, 5.021909, 4.333836, 3.923548, 5.108872, 7.895837, 9.602176, 
    10.12197,
  3.537305, 2.535074, 1.658272, 1.768196, 2.381169, 1.923571, 4.005203, 
    6.86781, 6.941155, 5.820214, 6.825029, 8.642351, 10.13863, 10.68263, 
    10.3035,
  3.753837, 3.125594, 2.765312, 3.312557, 3.456764, 3.754842, 6.328453, 
    8.469604, 7.986617, 7.015053, 8.237969, 9.145607, 9.49337, 9.352166, 
    8.398838,
  4.154312, 3.866297, 3.466787, 3.6934, 4.087505, 5.541384, 8.012986, 
    8.980663, 6.881265, 5.212565, 6.233058, 8.3337, 8.284302, 8.039257, 
    7.518186,
  4.139874, 5.313426, 4.647046, 5.20763, 4.424725, 3.470677, 4.597951, 
    5.213777, 5.387692, 3.952996, 3.502793, 3.844421, 3.514037, 3.084018, 
    2.847853,
  6.250857, 4.899128, 3.862625, 3.675088, 2.541308, 3.101267, 5.595132, 
    6.362526, 6.74505, 6.052496, 4.907429, 5.104503, 4.963714, 3.299234, 
    3.164437,
  4.375514, 2.987448, 2.565776, 3.415045, 2.730384, 2.975693, 3.958723, 
    4.960949, 5.418814, 5.012949, 4.875903, 4.908935, 5.017354, 4.881989, 
    4.373243,
  2.659741, 3.499525, 4.454097, 2.997904, 2.183897, 2.244921, 2.474054, 
    2.0145, 3.091057, 4.260273, 4.553153, 4.408583, 4.600162, 5.289343, 
    5.197583,
  3.797436, 4.562211, 3.476512, 1.174137, 1.385342, 3.43711, 3.420933, 
    1.96999, 2.308197, 2.448706, 3.996102, 4.795374, 5.308631, 5.70824, 
    5.640424,
  4.183165, 3.319977, 2.283719, 2.131538, 3.608833, 4.496775, 4.560292, 
    4.32713, 3.049601, 2.042998, 2.675695, 4.80942, 5.253915, 5.150731, 
    5.609466,
  3.348148, 2.370839, 3.007194, 3.647566, 4.464292, 4.219961, 3.186455, 
    2.936748, 3.772895, 4.75186, 4.508108, 4.164834, 4.74053, 5.560352, 
    5.945594,
  2.650772, 3.141231, 3.632376, 3.81172, 3.616614, 2.679405, 2.847957, 
    3.527498, 4.993868, 4.024334, 4.593348, 5.660214, 6.442445, 7.300256, 
    7.418613,
  3.170064, 3.639104, 3.641628, 4.085973, 3.809037, 4.253114, 4.380724, 
    3.900522, 3.277719, 5.63123, 6.939974, 8.103263, 8.69158, 8.426462, 
    7.355602,
  3.619398, 4.320367, 4.635872, 5.80089, 5.964645, 5.202258, 3.618671, 
    4.290895, 5.969665, 5.7955, 7.375075, 9.66654, 9.070355, 8.408607, 
    7.626259,
  6.951286, 8.211737, 5.704196, 6.329492, 5.453324, 3.819982, 4.398412, 
    4.489924, 4.57489, 3.641351, 3.130688, 2.485161, 1.836937, 2.073669, 
    2.240334,
  9.84689, 8.67444, 7.502655, 7.246634, 4.560812, 3.488399, 4.659251, 
    5.029404, 5.674293, 5.254243, 4.317807, 4.328439, 3.293462, 2.145339, 
    1.819131,
  9.877298, 8.865843, 8.163866, 6.943089, 4.383836, 3.100825, 3.368508, 
    3.812658, 4.38136, 4.855301, 4.534564, 4.514787, 4.672301, 3.883861, 
    2.632234,
  10.05776, 9.378069, 7.773365, 5.223779, 3.943919, 3.263061, 2.431302, 
    2.569374, 2.75157, 3.661907, 3.838027, 3.575348, 4.341745, 4.452459, 
    3.388782,
  9.698224, 7.777601, 5.952264, 4.167098, 3.706305, 4.387686, 4.350475, 
    2.595648, 2.623408, 2.43118, 2.96562, 2.897088, 3.640482, 4.52602, 
    4.002055,
  7.342583, 5.56784, 4.465336, 3.929983, 4.612629, 5.775061, 5.832896, 
    5.464408, 3.725378, 1.796152, 1.340501, 2.008973, 2.644294, 4.206679, 
    4.223235,
  5.667292, 4.395339, 4.042178, 4.391224, 5.91449, 6.098384, 5.03345, 
    4.182375, 3.619712, 2.323955, 1.472562, 1.915254, 2.900473, 3.84163, 
    4.180788,
  4.582212, 3.811191, 4.054387, 5.398933, 6.865443, 5.36956, 3.696454, 
    3.063359, 2.872461, 3.015983, 2.291061, 2.253057, 2.87734, 3.293851, 
    3.500862,
  3.35346, 4.195244, 4.747879, 6.680311, 5.686555, 3.580704, 3.776984, 
    3.205806, 3.043994, 3.399115, 3.197488, 2.755806, 2.793803, 3.274516, 
    3.523529,
  3.236859, 5.031218, 5.470143, 5.700101, 3.346754, 2.510483, 3.152459, 
    3.620443, 3.062619, 2.393375, 2.358036, 3.263083, 3.431242, 3.659453, 
    3.557984,
  7.514862, 9.824857, 7.352287, 9.732175, 9.116546, 7.762655, 9.671262, 
    10.36912, 9.989787, 7.091558, 6.575269, 6.608792, 5.796978, 4.293056, 
    3.233154,
  9.408909, 9.960472, 9.423143, 9.617181, 7.241876, 6.088988, 8.511043, 
    8.82201, 8.829655, 7.877429, 6.9923, 7.508587, 6.447099, 3.848763, 
    2.690461,
  9.175187, 9.317482, 9.373819, 9.850688, 7.549833, 5.641829, 5.189419, 
    7.031215, 8.741411, 9.350488, 8.587681, 7.171042, 5.451472, 4.253849, 
    3.031888,
  8.355904, 7.974255, 8.014946, 8.286335, 9.400252, 8.913497, 7.729734, 
    7.637066, 8.524625, 7.705036, 7.217003, 5.587894, 4.475292, 3.906973, 
    2.78859,
  6.810507, 8.006995, 10.30529, 12.19847, 11.84694, 11.31988, 9.359244, 
    6.516198, 5.072853, 4.43798, 5.056102, 4.756609, 4.254679, 3.985486, 
    3.300311,
  13.77484, 15.60547, 15.85187, 14.57053, 12.64516, 9.984213, 8.497131, 
    7.956007, 5.556458, 3.788006, 2.722496, 3.449403, 3.771075, 3.953672, 
    3.57748,
  14.49807, 14.79557, 13.58054, 11.87516, 10.31538, 9.050317, 8.005454, 
    7.198815, 6.200141, 4.624697, 2.533278, 2.155015, 3.55767, 4.362513, 
    3.957042,
  11.67555, 11.45954, 10.25152, 8.806629, 7.972268, 8.21123, 7.752204, 
    7.097328, 5.630671, 4.14741, 2.474146, 3.22913, 4.057134, 4.567956, 
    3.229941,
  8.337463, 8.072527, 7.082008, 6.586489, 6.905415, 6.989456, 6.636785, 
    5.810079, 4.629476, 3.674651, 3.048393, 3.632855, 3.80624, 3.399897, 
    1.6633,
  6.177373, 6.250618, 6.046633, 6.241143, 6.655776, 6.447309, 5.681068, 
    4.462315, 2.982006, 2.160694, 2.430608, 3.292431, 2.970126, 2.146874, 
    1.677321,
  5.72097, 10.89071, 11.26874, 15.27674, 14.31086, 10.81108, 12.19015, 
    12.22087, 11.18716, 7.934265, 7.88931, 8.050259, 7.173957, 6.369071, 
    6.263559,
  9.690592, 13.63069, 15.44635, 15.39377, 9.788487, 7.212472, 9.4973, 
    8.996441, 8.412619, 6.651915, 6.308527, 8.016592, 9.010255, 6.860663, 
    6.852462,
  11.72889, 13.79374, 13.78776, 12.32623, 7.385254, 4.321255, 3.328522, 
    4.447197, 4.643109, 3.702495, 3.36844, 4.757918, 7.612993, 9.871095, 
    8.799854,
  11.15307, 11.80562, 10.63273, 8.633683, 6.392814, 5.980621, 5.864886, 
    8.366776, 12.32363, 10.30205, 8.520135, 7.30755, 7.8245, 9.773837, 
    9.711141,
  9.015068, 9.373736, 9.390231, 11.17124, 12.72466, 11.65646, 8.813233, 
    6.165233, 6.672567, 7.352176, 9.855824, 10.70678, 11.54361, 12.09495, 
    11.35522,
  7.318593, 9.485225, 11.71869, 13.13711, 13.77845, 13.35336, 12.16605, 
    10.63297, 7.024369, 6.347711, 7.383781, 11.59708, 12.29952, 11.98062, 
    10.76521,
  6.090907, 8.251379, 10.12903, 11.19832, 11.50421, 11.21734, 10.77845, 
    10.19812, 9.026281, 8.671287, 8.947016, 9.888791, 10.3839, 10.1306, 
    8.845942,
  5.387882, 7.032693, 8.060462, 9.03459, 9.425648, 9.410253, 8.57325, 
    7.780239, 7.230688, 7.323253, 7.371324, 7.681136, 8.00717, 7.528951, 
    5.876077,
  5.08206, 5.622021, 5.860687, 6.653298, 7.107471, 7.415601, 7.293123, 
    6.954009, 6.455627, 6.122911, 6.412472, 6.67721, 6.553191, 5.346625, 
    3.731801,
  4.942921, 4.468466, 4.352119, 4.788554, 4.988835, 5.088184, 5.412005, 
    5.374502, 4.925735, 4.14259, 4.81939, 6.279142, 5.51935, 4.296762, 
    3.108459,
  5.968748, 7.305185, 6.826405, 8.830269, 7.691085, 4.883582, 5.743217, 
    6.006975, 6.24793, 5.933007, 7.219185, 8.473219, 8.254594, 6.990866, 
    6.003627,
  9.402742, 9.064221, 9.209753, 8.636412, 5.359462, 3.983577, 5.64474, 
    6.29171, 7.039519, 7.25579, 7.834287, 10.1854, 10.5866, 6.911164, 5.732992,
  10.70665, 9.669326, 9.110277, 8.385256, 5.296729, 3.568028, 4.613772, 
    5.229323, 6.62752, 9.007415, 10.79869, 11.32183, 11.12162, 9.845507, 
    6.596533,
  9.420182, 9.450794, 8.943141, 7.784721, 5.971469, 3.897571, 2.976371, 
    3.98045, 6.577118, 9.289709, 11.98551, 12.96907, 11.97711, 8.446168, 
    5.831782,
  11.11313, 9.57101, 8.309858, 6.461749, 4.895535, 4.266561, 3.764251, 
    3.107172, 4.681276, 6.915855, 12.05986, 14.01602, 13.39773, 6.518683, 
    5.243539,
  9.872309, 8.276926, 6.628011, 4.648084, 3.675263, 3.4346, 3.775557, 
    4.275279, 4.494422, 5.552221, 8.226834, 13.42265, 12.94719, 7.978747, 
    6.009706,
  7.097744, 6.102508, 4.480974, 2.928091, 2.659295, 2.921102, 3.707906, 
    4.83317, 5.625301, 7.096753, 9.685291, 11.7921, 10.49352, 9.065828, 
    9.562233,
  4.910827, 4.046904, 2.329307, 1.937584, 2.649029, 3.678136, 4.12321, 
    3.965254, 4.713819, 6.101606, 8.621233, 9.556819, 7.905096, 8.173949, 
    9.130311,
  3.836426, 2.339122, 1.195289, 2.049139, 3.142101, 3.985626, 4.299569, 
    3.845134, 3.968306, 5.002132, 7.044197, 7.642647, 6.123227, 6.386483, 
    7.497486,
  3.710315, 1.460558, 1.313709, 3.113223, 3.675033, 3.635947, 3.577955, 
    3.194839, 2.763613, 2.986612, 4.582068, 5.789166, 5.144267, 6.013829, 
    7.31798,
  9.729269, 13.91445, 12.36124, 15.94815, 13.65107, 9.850479, 11.41197, 
    11.41109, 10.06169, 7.158137, 6.590545, 6.146424, 5.447438, 5.097923, 
    5.27506,
  13.80319, 14.62388, 14.76513, 14.65693, 9.583276, 8.053489, 10.27617, 
    9.722125, 9.830834, 9.041741, 7.202137, 6.99773, 6.579993, 5.197864, 
    5.998962,
  13.14289, 13.64367, 13.33733, 12.95388, 10.20772, 8.623502, 9.552092, 
    11.65163, 11.70341, 9.241956, 7.184424, 6.70882, 7.372483, 9.027465, 
    8.68983,
  11.88571, 12.61122, 12.79486, 14.04561, 14.32402, 11.84466, 9.822556, 
    9.903992, 9.594731, 6.979484, 5.739778, 5.916625, 8.254464, 11.86062, 
    9.865947,
  10.77784, 12.59689, 13.95132, 14.88981, 14.28466, 12.59759, 9.097857, 
    5.987504, 4.590039, 3.60315, 4.351129, 6.276352, 10.08206, 12.2605, 
    7.300433,
  7.859733, 9.739417, 11.01322, 11.57216, 11.11636, 10.14733, 8.01201, 
    6.379817, 4.062398, 3.071515, 3.562857, 7.569849, 10.68195, 8.620585, 
    2.657441,
  5.296824, 6.470161, 7.50641, 7.613502, 7.53929, 7.075568, 5.723751, 
    4.913461, 3.842487, 3.500398, 5.598119, 7.849634, 8.121148, 5.760394, 
    3.970906,
  3.649451, 4.326989, 4.439634, 4.434964, 4.086006, 3.661545, 2.910617, 
    2.284777, 2.316835, 3.836531, 6.596104, 6.424726, 4.818917, 4.816568, 
    5.437138,
  3.214106, 3.241839, 3.014367, 2.848742, 2.256917, 1.6956, 1.901392, 
    1.580946, 2.277437, 4.459561, 6.206844, 4.503366, 3.59966, 4.779689, 
    5.755674,
  3.674176, 3.337338, 4.051155, 4.282445, 2.497905, 0.8963051, 0.9493821, 
    1.247668, 1.602904, 3.057186, 3.586511, 4.014008, 4.618836, 5.860037, 
    6.37162,
  4.566665, 5.73957, 4.776226, 9.004472, 10.62949, 9.920549, 13.0732, 
    13.46873, 11.38326, 7.308867, 5.808895, 8.269007, 10.13635, 9.050732, 
    7.210649,
  5.181449, 4.960437, 5.793924, 8.138896, 7.324691, 8.116054, 12.03615, 
    13.628, 12.8276, 10.70754, 9.945755, 12.19077, 11.72508, 7.203209, 
    5.532135,
  3.687866, 4.302346, 6.281939, 6.758329, 5.990911, 6.174798, 9.586873, 
    12.36067, 13.75897, 14.12669, 12.97893, 11.62341, 9.81438, 7.241813, 
    4.75776,
  3.57527, 4.261025, 6.032994, 5.734393, 6.822223, 5.847518, 5.281719, 
    8.708241, 13.06174, 12.35113, 10.52275, 8.411185, 6.099341, 4.020996, 
    3.45955,
  2.830256, 4.576725, 5.392044, 4.590339, 5.54865, 7.155675, 6.09657, 
    4.756941, 6.205981, 6.726479, 7.294, 5.880918, 3.95004, 2.963044, 3.145937,
  2.647658, 4.473223, 5.388419, 4.654811, 4.684464, 5.487415, 6.417318, 
    6.33904, 5.023706, 5.082079, 4.446656, 5.104445, 4.643462, 4.18486, 
    3.20596,
  2.702453, 4.005078, 5.803762, 5.976366, 5.01317, 4.09611, 4.562609, 
    5.834845, 7.110698, 7.252642, 6.13462, 5.00996, 4.513259, 4.019812, 
    4.551898,
  4.373045, 4.598917, 4.959938, 5.913389, 5.528434, 3.620597, 3.339463, 
    4.213918, 5.734076, 6.256017, 5.872817, 4.907413, 4.321795, 4.137877, 
    4.301745,
  5.0772, 4.412389, 4.051963, 5.335083, 5.539722, 3.9024, 2.606283, 2.986233, 
    4.918272, 5.525475, 5.072638, 4.719071, 4.449382, 4.470676, 4.361481,
  5.004166, 4.227044, 4.08257, 4.879226, 5.53793, 4.053899, 1.745789, 
    2.248958, 3.613988, 3.1782, 3.100884, 4.132089, 4.264055, 4.537349, 
    4.861667,
  2.578507, 3.231148, 2.561214, 4.925063, 5.086739, 2.323211, 4.025913, 
    6.487714, 8.278476, 7.449491, 7.180476, 7.46607, 7.135643, 6.302011, 
    5.44591,
  3.127608, 2.576297, 3.763133, 6.755276, 3.463165, 1.953717, 3.570992, 
    6.327447, 8.233388, 8.446393, 7.191055, 7.810575, 7.725171, 5.5847, 
    4.703831,
  3.768252, 3.876154, 6.302528, 6.109921, 2.517555, 1.693289, 3.756073, 
    5.298323, 6.92299, 8.837653, 8.930089, 7.944199, 7.548165, 7.383819, 
    5.481002,
  4.416405, 3.767884, 6.1043, 5.30712, 2.075357, 1.518629, 2.746898, 4.86742, 
    7.584758, 9.453128, 9.537274, 8.304862, 7.212005, 7.082396, 6.231048,
  4.486826, 3.137636, 4.852022, 4.799227, 3.033293, 1.559057, 2.593517, 
    2.990312, 4.765488, 6.403527, 8.613939, 7.902403, 6.944304, 6.742039, 
    6.546172,
  4.131157, 2.591176, 3.456842, 4.986271, 5.963345, 4.942424, 3.449689, 
    3.960803, 4.743459, 5.43875, 5.696213, 7.005308, 6.51423, 6.393756, 
    6.113472,
  3.390166, 3.603733, 3.839919, 4.936548, 6.081288, 6.192308, 4.423817, 
    3.517274, 6.008022, 7.42472, 7.760346, 7.058645, 6.262535, 6.419023, 
    5.870562,
  4.221092, 4.023413, 3.796343, 4.203461, 4.328714, 4.227703, 3.398725, 
    2.213709, 5.199077, 6.716758, 7.182174, 6.875724, 6.414193, 6.501583, 
    6.018156,
  4.524578, 4.364417, 3.964788, 3.79196, 2.668521, 4.240485, 4.480431, 
    2.290784, 4.747807, 6.01435, 6.493346, 6.50914, 6.365624, 6.673023, 
    6.215126,
  3.918012, 4.401687, 5.248535, 4.708655, 2.918736, 4.881489, 4.38554, 
    2.81492, 4.046171, 3.8797, 4.54807, 5.795297, 6.073484, 6.587388, 6.432084,
  6.084434, 8.068972, 7.148673, 9.391942, 7.63821, 4.500289, 3.958337, 
    3.901067, 4.587611, 5.030398, 6.142195, 6.770978, 5.903592, 4.924731, 
    4.509196,
  8.897402, 9.185845, 8.788509, 7.688766, 4.508142, 3.044667, 3.935743, 
    4.755202, 5.461016, 6.721138, 7.178289, 8.049959, 6.893485, 4.252796, 
    4.222587,
  9.776675, 9.475314, 8.15909, 5.832149, 3.321048, 2.3534, 3.575788, 
    4.193601, 4.412805, 7.137453, 9.176482, 8.838119, 7.165286, 5.842621, 
    4.733214,
  10.20061, 8.993945, 7.06308, 5.003005, 3.287555, 2.532403, 2.743251, 
    4.096309, 6.094682, 8.389143, 9.720734, 9.169725, 7.474607, 5.959756, 
    4.74121,
  9.630903, 7.618942, 5.382354, 3.422093, 2.354905, 3.138715, 3.713633, 
    3.413299, 4.675117, 6.331336, 9.042299, 8.821304, 7.585643, 6.355388, 
    5.603274,
  8.655436, 6.713774, 5.138793, 3.822802, 3.212048, 3.653519, 4.258744, 
    4.908537, 4.583368, 5.405103, 5.854782, 7.807315, 7.466548, 6.513604, 
    5.973603,
  8.139923, 7.02319, 6.195512, 5.8312, 5.426626, 5.067983, 5.010443, 
    5.900962, 6.118107, 7.22398, 7.674193, 7.48475, 7.054881, 6.797509, 
    6.750087,
  7.877615, 6.70252, 5.81726, 5.806335, 6.25481, 6.54376, 6.484674, 6.28363, 
    6.482932, 6.614762, 7.081485, 7.113154, 6.778552, 7.166646, 7.507485,
  7.425463, 6.194591, 5.142911, 5.270324, 6.013222, 6.565032, 6.526864, 
    6.728936, 6.841133, 6.61425, 6.861776, 6.88857, 6.504981, 7.3982, 7.377754,
  6.940652, 5.653308, 4.70545, 4.932364, 5.783169, 6.461397, 6.947235, 
    6.901775, 5.91229, 4.4483, 5.134927, 6.628623, 6.37788, 7.082258, 7.506353,
  7.443436, 8.830438, 5.396954, 4.750201, 3.270135, 2.818722, 3.909804, 
    4.881592, 5.520867, 5.115001, 5.798831, 6.164289, 5.122076, 3.939429, 
    3.399234,
  9.663918, 8.03284, 5.744534, 4.088457, 2.95023, 3.086249, 4.765794, 
    6.275388, 6.886387, 6.683034, 6.503424, 7.234287, 6.170165, 3.923161, 
    3.877316,
  8.937181, 6.808421, 5.370986, 4.837787, 3.702304, 3.262977, 5.176557, 
    5.564097, 5.552172, 6.78358, 8.149739, 7.822779, 6.793291, 6.016077, 
    5.126537,
  8.163181, 5.841264, 4.579003, 4.999186, 5.202277, 4.297071, 4.106473, 
    5.341384, 6.452888, 7.322016, 8.555694, 8.318347, 7.280718, 6.941268, 
    5.870325,
  7.479594, 4.904557, 3.850221, 4.556492, 5.276158, 6.032076, 5.238713, 
    3.868681, 4.857858, 6.067864, 8.293118, 8.437496, 7.780133, 7.704091, 
    7.375225,
  6.823903, 4.489832, 3.903683, 4.835734, 5.756822, 6.461123, 6.268765, 
    5.607107, 5.317203, 5.453798, 5.896907, 8.065314, 8.13402, 8.008396, 
    7.517764,
  6.649617, 4.540398, 3.912299, 4.838732, 6.160708, 6.957278, 7.027182, 
    7.011385, 7.186962, 7.482113, 8.161801, 8.538381, 8.160316, 7.997959, 
    7.327442,
  6.393133, 4.094501, 3.748367, 5.254678, 6.565691, 7.298712, 7.04408, 
    6.821303, 7.046202, 7.482174, 8.351067, 8.612493, 8.2096, 8.078849, 
    7.500876,
  5.885612, 3.516909, 3.436052, 5.16285, 6.680999, 7.516103, 7.304945, 
    7.294888, 7.433271, 7.648993, 8.230218, 8.667066, 8.335119, 8.150845, 
    7.238098,
  5.108588, 3.051543, 3.693625, 5.343654, 7.063961, 7.827036, 7.559279, 
    7.18174, 6.177115, 5.010316, 5.803638, 8.050215, 8.089046, 8.082212, 
    7.257362,
  4.652858, 5.687837, 3.892633, 4.096245, 3.675138, 3.24162, 4.678705, 
    5.744971, 5.276903, 4.323086, 4.893898, 5.643377, 5.921574, 5.314015, 
    4.437138,
  6.011617, 5.013546, 4.544637, 4.702092, 3.766623, 3.673494, 5.227595, 
    6.01695, 5.768956, 5.090009, 5.547692, 7.361078, 7.274546, 4.791304, 
    4.430137,
  5.446683, 4.104946, 4.402699, 5.234233, 4.175748, 3.863304, 5.813213, 
    5.324454, 4.412287, 5.4448, 7.457614, 8.258209, 7.389779, 6.097433, 
    4.668443,
  4.457997, 3.34329, 4.170568, 5.36531, 5.64071, 4.757866, 4.328369, 
    4.986431, 5.348096, 6.41604, 8.25492, 8.641547, 7.259491, 5.765297, 
    3.846611,
  3.530918, 2.958135, 4.400486, 5.608913, 6.418237, 6.280226, 5.076686, 
    3.546366, 4.447924, 5.863933, 8.596588, 8.541612, 6.638381, 5.41921, 
    4.349879,
  2.787829, 2.984489, 4.745108, 5.926569, 6.918806, 7.172493, 6.188945, 
    5.642689, 5.606257, 5.836391, 6.104379, 7.430709, 6.224082, 5.600541, 
    4.826008,
  2.327468, 3.119877, 4.951993, 6.005224, 7.194591, 7.651114, 7.514721, 
    7.446488, 7.367102, 7.451462, 7.540776, 6.785213, 5.937396, 6.010017, 
    5.424652,
  2.182599, 3.577334, 5.192337, 6.309313, 7.555552, 8.149636, 8.00158, 
    7.446622, 7.209827, 7.236029, 6.870722, 6.257405, 6.022545, 6.182257, 
    5.924354,
  2.468798, 4.096445, 5.090364, 6.066605, 7.470377, 8.350773, 8.612132, 
    8.162002, 7.480428, 6.857183, 6.294489, 5.977381, 5.75667, 6.037643, 
    5.84421,
  3.022678, 4.767258, 5.239201, 6.251131, 7.942361, 9.236679, 9.010199, 
    8.126148, 6.243183, 4.582788, 4.488494, 5.363643, 4.94983, 5.093126, 
    5.081191,
  3.510148, 3.568302, 2.806002, 4.886309, 5.043803, 4.324579, 5.466763, 
    6.211999, 5.265723, 3.81323, 3.734246, 3.765343, 3.623667, 3.105183, 
    2.425612,
  3.904027, 2.215195, 3.969098, 5.617564, 4.754234, 4.642085, 6.253866, 
    6.969957, 6.709616, 5.323512, 4.465867, 5.032444, 4.597116, 2.766902, 
    2.213319,
  2.657267, 2.096815, 4.741139, 6.218047, 4.965067, 4.791895, 7.098656, 
    6.999095, 6.56335, 6.15366, 5.988784, 6.003641, 5.31697, 4.338974, 
    2.918247,
  1.773443, 3.034988, 5.810017, 7.084332, 6.979499, 5.810116, 5.895841, 
    6.718745, 6.409164, 5.609342, 6.29279, 6.615903, 5.940412, 5.032027, 
    3.600158,
  1.667097, 4.263512, 6.921751, 7.377625, 7.999217, 8.027457, 6.860871, 
    5.492474, 5.540708, 5.209855, 6.528203, 7.233687, 6.519502, 5.743093, 
    4.945245,
  2.289981, 5.625086, 7.433821, 7.515643, 8.547606, 9.227502, 8.853489, 
    8.215578, 7.09355, 5.932242, 5.237381, 7.287799, 6.775018, 6.200098, 
    5.735801,
  3.296724, 6.371831, 7.230726, 7.425498, 8.513923, 9.400626, 9.962536, 
    9.552691, 8.247339, 7.005391, 6.31759, 6.48488, 6.379492, 6.306053, 
    6.155266,
  4.285204, 6.680775, 6.899928, 7.274683, 8.444448, 9.577949, 9.683411, 
    8.892779, 7.758016, 6.5441, 5.460681, 4.642043, 5.152205, 5.817284, 
    5.711402,
  5.298802, 6.598237, 5.905826, 6.692853, 8.098804, 9.300637, 9.475121, 
    9.125298, 7.778394, 6.037069, 4.555848, 3.276026, 3.289892, 4.267163, 
    4.80992,
  5.998925, 6.348254, 5.722981, 6.502735, 8.331654, 9.399215, 9.178941, 
    8.398985, 6.491601, 4.378747, 3.75394, 3.484225, 2.570668, 3.409486, 
    4.56056,
  3.961302, 3.938841, 1.829641, 4.699436, 5.891311, 5.200517, 6.694751, 
    7.049599, 6.163695, 4.568396, 4.229771, 4.079998, 3.293356, 2.255652, 
    1.060518,
  4.229977, 1.618651, 3.739586, 5.982693, 4.848755, 4.617608, 6.582582, 
    7.193106, 6.483713, 5.011147, 4.416325, 5.23716, 5.153856, 2.976444, 
    1.465423,
  2.775343, 2.231209, 5.220922, 5.918705, 4.368438, 4.428874, 6.048573, 
    6.471203, 5.894968, 4.564513, 4.280564, 5.206669, 6.387516, 5.509103, 
    2.988375,
  1.580218, 3.912913, 5.778943, 5.992256, 5.935798, 4.810228, 4.883358, 
    5.141255, 4.69748, 3.433193, 3.453153, 4.411375, 6.200716, 6.391632, 
    4.521099,
  1.811112, 4.622564, 5.565541, 5.945582, 7.150774, 6.784921, 5.486651, 
    4.167355, 3.729585, 2.996564, 3.397436, 4.070026, 6.063494, 7.200484, 
    6.282054,
  2.713555, 4.369704, 5.260134, 6.656686, 8.15206, 8.389306, 7.372664, 
    6.355908, 4.89603, 3.593253, 2.724032, 3.681464, 5.650462, 7.344178, 
    6.978189,
  3.133896, 4.079565, 5.329723, 7.428953, 8.923047, 8.948499, 8.393973, 
    7.00301, 5.895844, 4.757103, 3.384584, 3.168375, 5.46642, 7.440119, 
    7.587461,
  3.533773, 4.252082, 5.793657, 8.117177, 9.650985, 9.636585, 8.652927, 
    6.373183, 5.77106, 4.928487, 3.313741, 3.154536, 5.261129, 7.28497, 
    7.668458,
  3.573808, 3.954098, 5.501093, 8.180192, 9.947165, 10.16742, 9.327611, 
    7.2477, 5.756925, 5.121824, 3.532803, 3.54726, 5.374897, 7.187072, 
    7.789378,
  3.998962, 3.810606, 5.52222, 8.659118, 10.82462, 11.13792, 10.27442, 
    8.24513, 5.253314, 4.084838, 3.766505, 4.627475, 6.010468, 7.320277, 
    7.452598,
  4.593127, 5.074707, 2.829183, 3.132869, 3.529236, 3.273968, 4.066905, 
    3.635206, 3.582778, 3.031706, 3.436708, 3.918738, 3.376921, 2.220147, 
    1.807525,
  4.498754, 3.221072, 3.589457, 4.204761, 3.767017, 3.6548, 4.80493, 
    3.969554, 3.450287, 3.345849, 3.471351, 5.06222, 5.182308, 2.747345, 
    2.018504,
  3.032837, 3.294162, 4.384931, 5.314302, 4.478287, 4.144092, 4.083385, 
    3.87234, 3.631629, 3.751463, 4.271932, 5.895147, 6.059231, 4.322983, 
    2.739554,
  2.558171, 4.093118, 5.507698, 6.825188, 6.984971, 4.779856, 2.739717, 
    2.454788, 3.162791, 3.513704, 4.749067, 6.236986, 6.512786, 5.009397, 
    3.172538,
  2.782366, 4.510483, 6.428663, 7.508706, 8.055825, 5.857471, 3.00889, 
    2.584203, 2.635954, 2.77189, 5.345867, 6.559332, 7.024455, 5.780061, 
    4.02284,
  2.910197, 4.855429, 6.905313, 7.832013, 8.01616, 6.834067, 3.534248, 
    4.073774, 4.432196, 4.521874, 4.601462, 6.743392, 7.141952, 6.117825, 
    4.666445,
  3.274265, 5.305025, 6.869614, 7.855854, 7.984631, 7.089448, 5.770415, 
    4.831483, 6.657166, 6.610988, 6.302245, 7.137002, 7.444102, 6.716065, 
    5.443997,
  3.94106, 5.793549, 6.707504, 7.750443, 8.13084, 7.847519, 6.955901, 
    6.612029, 6.856847, 6.315151, 6.494046, 7.421209, 7.583839, 7.03123, 
    5.85858,
  4.553251, 5.828889, 6.401479, 7.339746, 7.756388, 7.778035, 7.255027, 
    6.620713, 6.167236, 5.627468, 6.346132, 7.734414, 7.794248, 7.138212, 
    5.852251,
  4.873408, 5.644233, 6.600768, 7.687816, 7.825012, 7.374688, 6.755183, 
    5.911225, 4.62433, 4.15536, 5.422693, 8.122777, 7.692417, 6.969933, 
    5.612424,
  2.112349, 1.938897, 1.765726, 3.007736, 3.607843, 3.383726, 3.611677, 
    3.124149, 2.323736, 2.529611, 3.153374, 2.56186, 1.154825, 1.660343, 
    3.134291,
  2.431624, 2.215174, 2.644233, 3.530991, 3.187398, 2.594927, 3.118295, 
    2.937578, 3.073661, 3.252403, 3.464662, 3.323867, 1.620951, 1.718469, 
    3.213398,
  2.929339, 2.28373, 2.808897, 3.442934, 2.92259, 2.292918, 1.253935, 
    2.495476, 3.680459, 4.25955, 4.613438, 3.831308, 2.004441, 2.945107, 
    3.559594,
  2.716973, 2.317202, 3.038785, 3.718026, 3.317595, 1.421009, 1.214193, 
    3.20164, 3.645521, 4.195246, 5.136121, 3.951216, 2.658972, 3.700219, 
    3.581654,
  3.203964, 3.193929, 3.749726, 4.000719, 3.304827, 1.494517, 2.019152, 
    2.985132, 2.949565, 3.444325, 4.869134, 3.51046, 3.16042, 3.6133, 3.604018,
  4.215957, 4.178389, 4.380737, 4.73728, 4.605488, 3.905914, 3.469256, 
    4.518987, 4.673696, 4.869235, 3.699721, 4.00953, 3.691201, 3.976868, 
    5.136459,
  5.293286, 5.105473, 4.723985, 5.308014, 5.684165, 6.054245, 6.177609, 
    6.432252, 7.134417, 6.768421, 5.680859, 5.13605, 5.160396, 6.101845, 
    7.085255,
  6.180939, 5.533978, 4.757706, 5.41505, 5.864539, 6.366319, 6.953441, 
    7.460179, 7.660124, 7.539793, 7.157724, 6.987378, 7.139089, 7.300676, 
    7.262776,
  6.645617, 5.55127, 4.867862, 5.394397, 6.046981, 6.633699, 7.160275, 
    7.644794, 7.972369, 7.876359, 7.823992, 7.867248, 7.747328, 7.659399, 
    6.848152,
  6.783386, 5.864025, 5.347458, 5.271443, 5.666945, 6.363478, 7.155316, 
    7.350777, 6.694509, 5.625304, 6.275286, 8.093423, 8.02153, 8.098676, 
    7.518355,
  5.323083, 6.547487, 5.45559, 5.773393, 4.494079, 3.247134, 3.727078, 
    3.38602, 1.75193, 0.4886339, 2.01238, 2.210936, 1.030248, 2.52713, 
    4.144566,
  8.345502, 7.513963, 5.910537, 4.555771, 2.687877, 2.226647, 3.644198, 
    3.457841, 2.489383, 1.120707, 1.519376, 1.480535, 1.29069, 2.536952, 
    4.44015,
  9.225501, 7.107168, 5.01255, 3.309081, 2.239658, 1.339236, 1.905803, 
    3.369461, 3.041189, 2.290324, 2.03644, 1.76213, 1.869601, 4.149532, 
    5.430993,
  8.716697, 6.133072, 3.624037, 2.211602, 2.323681, 1.456449, 0.9135218, 
    2.475263, 2.673128, 2.495208, 2.69638, 2.222168, 3.483416, 5.957811, 
    5.33309,
  7.802373, 5.197698, 2.733415, 1.621115, 1.725087, 2.182214, 1.578119, 
    1.877507, 2.085502, 1.929093, 2.625328, 2.593348, 4.748963, 6.040844, 
    4.535234,
  7.083781, 4.963465, 3.171259, 2.200475, 1.734929, 1.778754, 1.953367, 
    2.165243, 2.282483, 2.014568, 1.345366, 2.905423, 4.803412, 4.01893, 
    2.503887,
  6.672111, 5.107272, 3.578007, 2.925256, 2.974498, 3.277131, 3.269618, 
    2.453985, 1.912932, 2.082134, 2.76304, 3.444835, 3.222574, 2.305282, 
    3.39055,
  6.313592, 5.131826, 3.769, 3.315205, 3.236792, 3.044706, 2.912228, 
    2.444618, 2.155585, 2.42624, 2.993462, 3.111759, 2.5107, 3.674245, 
    5.255366,
  6.613481, 5.810369, 4.977878, 4.545085, 4.115565, 3.528343, 3.35208, 
    3.157401, 3.158082, 3.301092, 3.54069, 3.554394, 4.45442, 5.541081, 
    5.997453,
  7.168694, 6.748442, 6.243951, 5.765567, 5.314854, 4.573498, 4.395575, 
    3.969903, 3.410305, 2.950871, 3.758171, 5.870842, 6.393638, 6.925784, 
    7.378078,
  4.492879, 6.433449, 7.76363, 11.72882, 11.37677, 8.596026, 9.78044, 
    8.486322, 5.825492, 3.542471, 2.935062, 2.703412, 2.132231, 2.76632, 
    3.964048,
  7.25491, 9.197427, 10.8113, 13.05062, 9.334537, 7.148826, 8.657099, 
    7.445328, 4.729696, 2.768892, 1.851113, 1.929201, 2.750225, 3.308379, 
    5.005332,
  9.133286, 10.37429, 11.49125, 11.67111, 8.263697, 6.10818, 6.297534, 
    5.880544, 4.005445, 2.244102, 1.028944, 2.146568, 3.810201, 6.089744, 
    6.558998,
  10.80422, 10.92151, 10.69419, 9.583282, 8.033422, 6.225557, 4.681412, 
    3.753198, 2.82775, 2.396253, 2.491693, 3.454337, 5.575734, 8.039979, 
    6.239913,
  10.9298, 9.879169, 8.806252, 7.58128, 6.060916, 5.558741, 5.312748, 
    3.451055, 2.170838, 2.142968, 2.676457, 4.133526, 6.447542, 8.393238, 
    5.89833,
  9.60912, 8.315928, 6.860953, 5.413033, 5.005381, 4.45375, 4.302803, 
    3.793687, 2.180811, 1.483281, 1.451653, 4.567258, 7.31517, 6.585628, 
    3.365438,
  7.406801, 6.300727, 4.731768, 3.215047, 3.587983, 4.155447, 3.711793, 
    2.847689, 2.703008, 1.982354, 2.494646, 5.964189, 6.285355, 3.166959, 
    3.56909,
  4.813438, 3.777536, 2.545421, 2.09554, 2.730744, 3.716673, 4.465297, 
    4.513498, 3.074902, 1.642556, 4.473336, 5.8209, 3.281438, 3.014512, 
    5.099977,
  3.12783, 2.373512, 2.308245, 2.251225, 2.797329, 3.538068, 4.328125, 
    4.173468, 2.396126, 3.037446, 4.732606, 3.090226, 2.614494, 4.889056, 
    6.427299,
  2.844944, 2.6435, 2.811254, 2.899779, 3.174659, 3.664759, 4.474132, 
    3.830334, 2.577326, 2.490495, 2.144869, 2.316149, 4.677498, 6.607718, 
    8.245794,
  3.350342, 5.208306, 6.038963, 8.616463, 8.686428, 8.7562, 12.02026, 
    11.78938, 10.21155, 7.068875, 5.923479, 4.519629, 2.785463, 1.654064, 
    1.48364,
  5.3555, 7.510163, 9.335673, 11.29968, 9.899303, 9.979164, 12.57156, 
    11.65946, 9.93343, 7.819829, 5.194863, 3.840545, 2.149468, 1.291052, 
    2.044202,
  6.043754, 8.786137, 11.02838, 13.63931, 11.7241, 10.39064, 10.38643, 
    10.4472, 9.45225, 6.848524, 3.904366, 2.180785, 2.402987, 4.099425, 
    3.779627,
  7.582534, 10.77722, 12.95332, 13.91485, 13.88465, 11.52383, 8.989481, 
    7.405899, 5.563577, 2.973212, 1.481692, 2.611008, 4.956118, 6.281328, 
    4.583825,
  9.399341, 11.84604, 13.312, 13.48678, 12.35805, 11.5807, 9.717013, 
    5.986004, 2.646849, 1.27721, 1.314972, 4.460739, 6.437719, 6.547581, 
    4.211971,
  10.85648, 12.65913, 13.33466, 13.27221, 12.25133, 9.212277, 6.898428, 
    6.391608, 3.825391, 2.255361, 2.226424, 6.236782, 6.470547, 4.483719, 
    1.901668,
  11.71817, 13.01267, 13.22054, 12.7942, 11.27023, 9.183258, 7.193345, 
    6.416307, 5.320942, 3.260052, 4.776575, 6.157645, 4.704956, 2.911617, 
    3.046642,
  11.7401, 12.48563, 12.17059, 11.39424, 10.24799, 9.05962, 8.061252, 6.9768, 
    4.076562, 3.067142, 5.769854, 5.26148, 3.317932, 3.028853, 3.943807,
  10.64422, 11.24398, 10.80005, 10.00642, 9.313128, 8.498592, 7.070443, 
    4.675784, 2.478216, 4.377243, 5.805562, 4.131948, 2.710633, 3.102617, 
    4.122482,
  9.296144, 9.909732, 9.565985, 8.769542, 8.302839, 7.68655, 5.994524, 
    3.138779, 2.053572, 3.458204, 3.645, 2.623274, 3.120944, 4.449511, 
    6.079962,
  5.307834, 7.689221, 7.622944, 9.7141, 8.68327, 7.380922, 9.327675, 
    10.15812, 9.891477, 8.08188, 7.439319, 6.788157, 5.105536, 3.205649, 
    1.69473,
  5.611659, 7.56321, 9.22979, 10.10778, 8.226689, 7.674519, 9.963756, 
    10.82749, 10.81592, 9.580626, 7.658125, 7.511306, 5.391117, 2.318782, 
    1.142509,
  5.429908, 7.922499, 9.628836, 11.59921, 9.594709, 9.251943, 9.762693, 
    11.10141, 11.57088, 10.15805, 8.61991, 6.21192, 3.881357, 2.844165, 
    2.097631,
  7.768142, 9.288099, 9.966231, 11.23137, 11.35087, 11.46286, 10.1517, 
    9.455685, 8.641166, 6.929673, 5.737508, 4.211576, 3.863485, 4.763323, 
    4.456717,
  8.752702, 9.784859, 10.36541, 11.71821, 12.05754, 11.72865, 10.18772, 
    7.656278, 4.667713, 3.585036, 4.174286, 4.538383, 5.643821, 6.604434, 
    6.9301,
  9.59452, 10.52079, 10.773, 12.48745, 12.13482, 9.108303, 7.285314, 
    8.210038, 6.301459, 3.836416, 2.390356, 4.6243, 5.885256, 4.945672, 
    4.600136,
  10.02547, 11.35627, 12.34851, 12.92678, 12.12183, 10.40443, 9.057784, 
    8.124415, 6.617699, 3.035604, 2.574009, 3.151957, 2.805465, 1.854979, 
    2.43291,
  11.29556, 12.68254, 12.9415, 12.74332, 11.71804, 10.57476, 9.650527, 
    7.645362, 4.509909, 2.370878, 1.807746, 1.807232, 1.990548, 2.168762, 
    2.539461,
  12.91545, 13.71483, 13.38867, 12.56792, 11.47421, 9.834125, 7.635831, 
    5.533505, 4.10456, 3.548961, 3.344698, 2.853104, 2.432015, 2.437912, 
    2.866537,
  13.95029, 14.13318, 13.29822, 12.03456, 10.32614, 8.354545, 6.305112, 
    4.951518, 3.538447, 2.610122, 2.714729, 3.32082, 3.021569, 3.684152, 
    4.939462,
  7.526241, 7.237547, 4.913599, 3.717779, 4.881094, 4.999369, 5.297647, 
    4.777257, 5.927516, 6.466885, 7.492273, 8.225288, 7.706977, 5.316778, 
    3.641923,
  10.49711, 9.152086, 7.659022, 5.21232, 3.660429, 3.583177, 4.731077, 
    5.248475, 5.314406, 6.421004, 7.767774, 9.471597, 9.949802, 5.421128, 
    3.854753,
  8.408777, 8.981205, 8.058387, 6.840285, 4.497072, 2.910816, 2.926933, 
    4.303191, 5.419873, 7.577154, 9.452744, 9.979228, 9.779704, 7.319693, 
    5.187578,
  8.334959, 8.723668, 8.020819, 7.08527, 5.888256, 4.187221, 2.952271, 
    4.458419, 5.933664, 5.969016, 9.507608, 10.72703, 9.22171, 7.135568, 
    5.136609,
  9.621422, 8.907662, 8.206658, 7.200862, 6.004178, 5.434869, 5.187474, 
    4.377917, 3.655417, 4.096328, 8.672186, 10.30171, 8.913139, 7.125668, 
    5.653861,
  11.07155, 9.748174, 8.56524, 7.343872, 6.000964, 5.070413, 5.016436, 
    6.618071, 6.239886, 6.766042, 6.933266, 9.174501, 7.758317, 6.386684, 
    5.192681,
  11.42555, 10.55178, 9.491512, 8.499122, 7.986619, 7.880147, 8.305653, 
    9.156181, 10.26504, 9.869476, 8.982243, 7.327109, 5.544071, 4.290128, 
    3.710449,
  11.92553, 11.81993, 11.26685, 11.04438, 11.1989, 11.55454, 11.74076, 
    11.36943, 10.16096, 8.390798, 6.462622, 4.369446, 3.246639, 2.380667, 
    2.091633,
  11.96248, 12.18665, 12.01363, 11.97761, 11.73215, 11.22076, 10.24617, 
    9.023, 7.407491, 5.753458, 4.044907, 3.276837, 2.917262, 1.851512, 
    1.195624,
  11.50305, 11.76998, 11.78285, 11.25272, 10.46975, 9.729711, 8.643811, 
    7.310935, 5.198575, 3.480392, 3.444107, 4.661504, 4.302035, 3.258085, 
    2.805991,
  2.775185, 2.917824, 1.746094, 2.980581, 5.625031, 5.513534, 7.09855, 
    7.635716, 7.122707, 5.290862, 5.582362, 5.909791, 6.439266, 5.463192, 
    3.993279,
  5.283486, 3.888653, 2.087459, 3.269582, 4.289331, 5.305911, 7.657098, 
    7.789406, 7.909644, 7.392296, 6.806741, 7.574872, 8.478504, 5.611314, 
    5.121096,
  5.553885, 4.30358, 3.835726, 5.100145, 4.684995, 5.183946, 6.594779, 
    7.320766, 8.085533, 8.609184, 8.70574, 8.567899, 8.700787, 8.671327, 
    6.94019,
  5.488324, 4.842212, 4.946596, 5.928045, 6.545852, 5.510627, 5.21764, 
    5.897007, 6.834455, 7.679961, 9.209903, 9.566014, 9.291985, 9.03583, 
    7.329372,
  5.362506, 4.960872, 5.028304, 5.274485, 5.544338, 7.001375, 5.900908, 
    5.005644, 4.132093, 4.765216, 8.547848, 10.16649, 10.53114, 9.630301, 
    7.731281,
  5.255696, 5.200638, 5.220131, 5.081663, 4.868718, 5.731453, 6.00887, 
    4.752025, 4.232653, 5.604672, 7.213036, 10.74067, 10.57784, 9.220948, 
    7.041637,
  5.762497, 6.125134, 6.05367, 6.334447, 6.536511, 6.609125, 6.704527, 
    6.584285, 7.490578, 9.144408, 10.31174, 11.23734, 10.50544, 8.979618, 
    7.222423,
  7.868483, 8.690602, 8.761815, 9.624242, 10.41031, 10.4961, 10.42792, 
    10.56252, 10.68561, 10.94197, 10.95002, 10.67942, 9.49915, 8.061516, 
    6.639201,
  10.26575, 10.68256, 11.03351, 11.87033, 12.45729, 12.77293, 12.67363, 
    12.1485, 11.56225, 10.61618, 9.979596, 9.405378, 8.292573, 6.856054, 
    5.544287,
  10.56089, 10.61128, 10.98563, 11.06623, 11.25851, 11.35075, 11.32848, 
    10.91902, 8.958592, 6.682334, 6.698585, 7.867575, 6.573941, 5.267165, 
    4.123254,
  3.474753, 4.03143, 3.61297, 4.792715, 4.522716, 3.701345, 4.296802, 
    5.308021, 5.976187, 3.147759, 1.533848, 2.516747, 4.161571, 4.225686, 
    3.292921,
  6.068634, 6.142813, 5.692944, 5.527792, 3.549018, 3.501865, 4.929893, 
    5.438673, 6.058026, 4.142796, 1.442838, 2.664692, 5.2005, 4.064755, 
    3.833578,
  7.607922, 7.637062, 7.458606, 7.411335, 5.559192, 4.101174, 4.206063, 
    5.633392, 6.764155, 5.194894, 2.338679, 2.716835, 4.377849, 5.963567, 
    5.901174,
  8.81743, 8.713732, 8.180127, 8.840391, 10.11609, 7.330832, 4.866857, 
    4.457161, 5.576282, 4.670491, 3.037865, 2.787762, 4.038094, 6.049178, 
    6.69073,
  10.35898, 9.84794, 8.794621, 7.714772, 10.6164, 11.21926, 9.345628, 
    6.765659, 4.485798, 3.19539, 3.672823, 3.478301, 4.557477, 7.062501, 
    9.156579,
  11.62296, 11.15017, 9.368301, 4.892226, 9.188533, 12.13107, 11.08555, 
    9.318898, 6.086436, 4.301757, 3.350479, 4.44818, 5.385212, 7.165557, 
    8.21145,
  12.52827, 12.45267, 9.601436, 5.149517, 8.509732, 11.91973, 10.20848, 
    7.908988, 7.060442, 6.351167, 5.486054, 5.70435, 6.413223, 7.563715, 
    8.043307,
  12.96172, 13.46305, 11.47878, 8.597486, 10.17907, 11.18448, 9.688319, 
    8.886436, 7.793475, 6.538233, 5.887767, 6.460299, 7.090076, 8.111259, 
    8.338476,
  12.59676, 13.68254, 12.92204, 11.73626, 11.65816, 11.19165, 9.675533, 
    8.464055, 7.507902, 6.600886, 6.50205, 7.328193, 8.064488, 8.816447, 
    8.544014,
  11.35092, 13.34006, 14.06527, 13.11353, 11.84958, 10.89121, 9.806964, 
    8.713435, 6.831774, 5.023928, 5.552676, 8.229177, 8.6334, 8.820601, 
    7.682074,
  3.401387, 4.799524, 4.998209, 6.078526, 5.66992, 4.647433, 5.394286, 
    5.041995, 4.496493, 3.719604, 2.720994, 2.499259, 2.566438, 2.869145, 
    3.320728,
  6.023068, 7.245213, 7.604006, 7.687506, 4.74919, 4.038935, 5.459596, 
    4.806417, 4.821895, 4.230046, 2.23188, 2.709743, 3.970801, 3.321084, 
    3.973204,
  7.291216, 8.892542, 8.967738, 8.243851, 5.659421, 4.175705, 3.968385, 
    3.966854, 4.185298, 4.115258, 2.124917, 2.641604, 4.525533, 5.477861, 
    6.610081,
  8.944961, 9.966869, 9.834556, 8.9939, 8.546962, 6.012475, 3.395938, 
    1.705111, 2.641578, 2.639133, 1.630827, 2.882981, 4.676459, 6.273156, 
    7.536399,
  10.50753, 10.64167, 10.37319, 9.196906, 8.716568, 8.842624, 6.916265, 
    3.754986, 2.162327, 1.709227, 1.882211, 3.263948, 5.726909, 7.984727, 
    9.745482,
  10.94326, 10.70656, 9.610979, 8.509042, 8.210636, 8.889717, 8.902181, 
    6.590706, 3.745441, 2.553494, 1.751889, 4.125323, 7.079236, 8.360414, 
    8.421423,
  10.9354, 10.42124, 7.964578, 6.266479, 7.181136, 8.60927, 8.203122, 
    5.25493, 4.187626, 3.781818, 3.039828, 5.865248, 7.525175, 8.315766, 
    8.487534,
  10.57152, 9.63395, 5.814607, 2.792288, 6.995783, 9.056296, 8.712554, 
    6.754275, 5.431685, 4.096931, 4.446428, 6.635538, 7.53808, 8.418462, 
    8.991082,
  10.25154, 9.54628, 6.980147, 6.535919, 9.024757, 9.564078, 8.338859, 
    6.484004, 5.737754, 4.848068, 5.348483, 6.889003, 7.924553, 9.142179, 
    9.436306,
  9.27603, 9.409713, 9.300041, 9.21309, 9.251458, 8.930807, 7.924055, 
    7.139286, 5.321671, 3.727863, 4.328834, 6.857671, 8.261016, 9.399374, 
    8.371819,
  3.006135, 4.124927, 3.927167, 5.014788, 4.867869, 4.740211, 6.50417, 
    6.965465, 6.875519, 5.337157, 5.605123, 5.746657, 4.917598, 4.230541, 
    3.955782,
  3.519307, 4.0101, 4.527236, 5.289698, 3.879048, 4.286747, 7.163624, 
    7.425045, 7.560474, 6.754385, 6.128335, 6.518106, 5.7101, 3.889907, 
    3.899985,
  2.880117, 3.733949, 5.278544, 6.434294, 5.325291, 4.597637, 5.824998, 
    7.099271, 7.338202, 6.970058, 6.856325, 6.515921, 5.860122, 5.290824, 
    4.135547,
  4.955483, 7.262222, 8.642375, 9.233256, 9.509992, 7.329875, 4.692343, 
    3.856311, 5.313264, 5.996239, 5.702863, 5.185871, 4.759024, 4.388706, 
    4.027902,
  8.882757, 9.896937, 10.36273, 10.24376, 10.17361, 10.00041, 7.982892, 
    4.641161, 3.179333, 2.839556, 3.228874, 3.740078, 3.482846, 4.308908, 
    5.62497,
  10.05221, 10.00775, 9.586461, 9.440598, 9.446986, 9.484324, 9.901513, 
    8.893309, 4.272437, 2.597857, 2.84728, 4.253334, 4.096179, 5.899557, 
    6.333845,
  9.309406, 8.486599, 7.797218, 7.053235, 7.272843, 7.616357, 7.826637, 
    7.328125, 5.71084, 5.384355, 5.826317, 4.815242, 6.363375, 7.066927, 
    8.355978,
  7.70793, 7.470363, 5.633401, 3.642552, 3.818337, 5.482789, 6.309928, 
    6.140309, 5.447157, 5.578964, 4.697579, 6.202789, 7.736673, 8.950753, 
    10.57773,
  7.013495, 6.398411, 5.26811, 4.039137, 4.213778, 5.327099, 5.640692, 
    4.369602, 3.605803, 3.595146, 5.538477, 8.392316, 9.809714, 11.18912, 
    10.84591,
  6.065263, 6.260602, 6.054527, 5.466807, 4.979349, 4.873323, 4.182468, 
    3.052818, 2.438024, 3.288848, 6.758769, 10.36036, 10.71399, 10.83041, 
    9.498553,
  4.771297, 5.949106, 5.023509, 6.229692, 5.449824, 4.035744, 5.012703, 
    4.628866, 3.813023, 2.893858, 2.82701, 2.773844, 3.60579, 5.645966, 
    7.049871,
  6.757607, 6.791123, 6.209363, 6.189419, 4.560802, 3.596622, 4.863028, 
    4.686846, 4.255019, 3.765617, 2.78407, 3.077784, 5.096293, 5.588117, 
    7.706246,
  7.650397, 7.089321, 5.870754, 5.525173, 4.86857, 3.644294, 3.756277, 
    5.081248, 5.348271, 4.457025, 3.44089, 4.22905, 6.102228, 7.587686, 
    8.150611,
  7.952559, 6.06117, 5.626781, 5.469392, 5.68918, 5.008163, 3.657321, 
    3.124814, 4.282526, 4.57151, 4.282172, 3.970725, 4.565882, 6.756877, 
    6.686429,
  5.407135, 5.529634, 5.854462, 5.981646, 6.046612, 6.716352, 6.582891, 
    4.765185, 3.114243, 2.752347, 3.145581, 1.897676, 2.411053, 5.718931, 
    5.903516,
  4.664464, 4.8297, 5.366481, 5.856351, 6.425826, 6.927681, 8.215537, 
    8.86484, 5.270947, 3.002533, 2.44902, 2.46829, 2.399898, 4.939703, 
    4.703473,
  5.351723, 4.886478, 5.206175, 5.956482, 6.73502, 7.082877, 7.439281, 
    7.771141, 6.7937, 5.499582, 4.87675, 3.715677, 1.741023, 3.540948, 
    5.372167,
  5.445718, 5.405824, 5.626616, 6.256125, 6.592615, 6.874523, 7.275496, 
    8.053418, 8.352966, 6.994541, 5.895192, 4.14114, 1.775428, 3.206836, 
    6.805009,
  6.080042, 6.42066, 6.407734, 6.309405, 5.47905, 5.430425, 6.60751, 
    7.614252, 8.203394, 7.689709, 6.755205, 4.499308, 2.806082, 5.298325, 
    7.330272,
  6.889575, 7.500194, 6.26756, 4.844078, 3.857524, 4.526871, 6.228007, 
    7.719975, 7.361559, 5.608391, 5.159583, 4.906621, 4.632962, 7.199097, 
    8.112029,
  8.764199, 7.877611, 3.822595, 6.283848, 6.7219, 7.304638, 11.16217, 
    10.94514, 9.575599, 8.034684, 7.199025, 5.285167, 3.382046, 3.426749, 
    3.535747,
  11.09461, 7.344759, 5.278272, 7.617711, 6.763711, 7.394744, 10.34596, 
    10.68228, 10.42392, 9.744804, 7.116471, 5.4765, 4.108067, 2.740862, 
    3.131847,
  11.55522, 7.387227, 5.737859, 8.224138, 7.91221, 7.439523, 7.953716, 
    9.52312, 10.98675, 9.61219, 6.706225, 4.53324, 3.87944, 3.923696, 3.331713,
  13.95558, 8.540824, 5.74445, 8.3228, 9.248665, 8.835874, 8.230157, 
    8.266933, 8.645768, 6.557708, 5.270415, 3.559714, 3.500555, 4.19592, 
    3.542605,
  13.78609, 11.08038, 5.937087, 8.553916, 8.92709, 9.68792, 10.15031, 
    8.102933, 4.677975, 3.215854, 4.056982, 3.150974, 3.295597, 4.016831, 
    4.453091,
  10.70099, 11.17075, 7.400594, 8.373795, 8.566898, 8.252116, 8.334518, 
    8.139454, 5.852145, 4.594676, 3.669826, 3.87785, 3.53408, 4.359591, 
    5.513425,
  6.511325, 8.523251, 7.165061, 7.074338, 7.486809, 7.515647, 6.658889, 
    6.399565, 7.071671, 6.789527, 5.755173, 4.300159, 4.09647, 5.549392, 
    6.638815,
  3.05358, 5.153729, 5.663061, 5.855079, 6.63325, 7.132846, 7.279863, 
    7.49727, 7.583908, 6.752384, 5.65288, 4.425648, 4.613679, 5.595643, 
    5.959683,
  2.464071, 3.039056, 4.455592, 5.464352, 6.191049, 6.844649, 6.970182, 
    6.994821, 7.271744, 6.26518, 5.340816, 4.75932, 4.806981, 4.995825, 
    4.843226,
  3.597784, 3.944723, 4.817676, 5.82425, 6.345942, 6.919253, 7.383012, 
    7.608333, 6.376141, 4.334155, 4.166292, 5.222756, 4.974719, 5.256585, 
    5.723138,
  6.341107, 10.83976, 8.823115, 8.45902, 6.418128, 5.029895, 8.196727, 
    10.25821, 10.51389, 8.505161, 8.62526, 8.035576, 6.744782, 5.339475, 
    3.804637,
  8.181557, 10.53881, 9.140781, 7.629435, 7.155796, 7.540196, 10.86221, 
    10.97253, 10.91008, 9.448105, 8.784444, 8.567597, 7.219652, 3.960924, 
    2.651301,
  7.495365, 10.00955, 7.287779, 6.17613, 6.74229, 6.471496, 9.245654, 
    10.93628, 11.83895, 10.6849, 9.28597, 8.008835, 6.425981, 4.450497, 
    3.078124,
  7.042449, 9.210582, 5.427816, 5.182, 7.255434, 6.085771, 6.787819, 
    9.385942, 10.59398, 8.583773, 8.145993, 7.170505, 6.341466, 5.249379, 
    4.17452,
  6.544911, 7.827337, 3.895379, 4.754435, 6.48583, 6.094203, 5.155256, 
    5.562873, 4.656131, 4.46014, 6.416672, 6.716185, 6.606447, 6.119861, 
    5.711893,
  6.064644, 6.82529, 3.312964, 4.356499, 5.873203, 4.8548, 4.45834, 6.34875, 
    6.056769, 4.926392, 4.923239, 6.847845, 6.498847, 6.422534, 6.095851,
  5.48048, 6.190969, 3.048249, 4.740534, 6.230367, 5.760315, 6.464291, 
    7.865478, 7.731878, 7.204741, 7.013679, 6.785767, 6.148965, 5.487364, 
    5.142855,
  4.501649, 5.534325, 3.030907, 5.187149, 7.428945, 7.269705, 8.378889, 
    9.425632, 8.847477, 7.961762, 6.956933, 6.220843, 5.152202, 4.328479, 
    3.843132,
  3.320643, 4.420231, 3.143526, 5.021569, 8.350395, 8.55103, 9.314709, 
    9.098018, 8.541685, 7.377637, 6.201391, 5.211763, 4.265819, 3.73057, 
    3.515331,
  2.11459, 3.172889, 3.814344, 4.669136, 8.963868, 9.932427, 10.45922, 
    9.417968, 7.040546, 4.769721, 4.464002, 4.746527, 4.236407, 4.254245, 
    4.433413,
  4.895441, 5.457362, 4.031568, 4.493909, 3.857341, 3.617407, 5.290527, 
    5.984023, 6.37107, 5.144282, 5.409388, 5.639904, 5.631036, 5.592321, 
    5.372873,
  8.102873, 7.298892, 5.954859, 5.377881, 4.063879, 4.190941, 6.227142, 
    6.444605, 6.539688, 5.88177, 6.027861, 6.581379, 6.318485, 4.006005, 
    3.662915,
  9.121426, 8.567737, 7.455547, 6.736969, 5.518513, 4.586431, 5.630278, 
    6.667044, 6.962353, 6.561688, 6.562931, 6.822064, 6.514612, 5.091942, 
    3.339982,
  10.98028, 10.25864, 8.935369, 8.235326, 7.877962, 6.551228, 5.26802, 
    5.207098, 5.47281, 5.237845, 6.260062, 6.594309, 6.208323, 5.437226, 
    4.132678,
  12.33615, 11.14355, 10.11714, 9.42401, 8.550694, 8.181841, 6.777822, 
    4.605456, 3.437151, 3.667571, 5.783823, 6.136298, 5.606153, 5.140803, 
    4.397835,
  12.36541, 11.39334, 10.79798, 10.13558, 9.339741, 7.896911, 6.313283, 
    5.731121, 5.243187, 5.344291, 4.600097, 5.599951, 4.403528, 3.585338, 
    2.895682,
  11.13799, 10.48782, 10.51179, 10.64107, 9.75931, 8.128725, 6.452934, 
    5.876254, 7.308482, 7.705529, 6.22604, 4.935259, 3.044804, 2.082412, 
    2.440267,
  10.26757, 9.168105, 8.163693, 9.404113, 9.871246, 8.931346, 8.622907, 
    8.781632, 8.913465, 8.094223, 6.12072, 4.054743, 2.287678, 1.963428, 
    2.455557,
  8.219985, 7.811659, 6.362936, 7.928233, 10.07164, 9.425247, 9.13597, 
    9.001863, 9.037432, 7.344121, 5.119528, 3.284714, 2.222678, 2.597287, 
    2.76496,
  5.468838, 6.100594, 4.881977, 7.096457, 9.525796, 9.74007, 9.873559, 
    9.686917, 7.647559, 4.871364, 3.827992, 3.247207, 2.481851, 3.314687, 
    3.656773,
  4.856919, 5.958483, 5.300701, 5.3798, 3.783406, 2.76229, 3.330795, 
    3.144691, 3.382277, 2.92728, 3.252316, 3.177695, 2.984639, 2.936482, 
    3.097259,
  6.451963, 5.960823, 5.993693, 5.053934, 3.156441, 2.644112, 3.909877, 
    4.016714, 4.257825, 3.954369, 4.310053, 4.560706, 4.006134, 2.129683, 
    1.725881,
  5.880063, 5.197948, 4.845639, 4.381755, 3.0066, 2.523216, 3.56987, 
    4.446575, 5.119485, 5.123972, 5.747009, 5.815612, 4.426738, 3.252071, 
    2.241172,
  4.473745, 4.154109, 4.345843, 4.675807, 4.20635, 3.647499, 3.448128, 
    3.735668, 4.478722, 5.01586, 5.904694, 6.210719, 5.162748, 4.021371, 
    3.07535,
  3.681, 4.737454, 6.289669, 6.7519, 6.910068, 6.755624, 6.123393, 4.313725, 
    3.988552, 3.810951, 6.034224, 6.642538, 6.113847, 5.009855, 3.736877,
  5.908927, 7.572368, 8.816413, 9.374795, 9.498336, 9.725106, 9.605769, 
    9.472946, 6.600896, 5.38523, 5.160168, 7.16326, 6.667161, 5.208774, 
    2.838696,
  8.179172, 9.731719, 10.82516, 11.30585, 11.5391, 10.96843, 11.1731, 
    9.927972, 9.069762, 9.173327, 8.463593, 7.938223, 6.968513, 4.792111, 
    2.549035,
  9.874085, 11.24985, 12.29174, 12.82271, 12.90779, 12.52697, 12.52957, 
    11.13676, 10.71719, 10.27648, 9.23417, 8.477435, 6.964707, 4.462785, 
    2.284553,
  10.45598, 12.26689, 12.51635, 13.77858, 13.29644, 13.64802, 13.08269, 
    11.76047, 11.20545, 10.47052, 9.786209, 8.750044, 6.731177, 4.37383, 
    2.644032,
  9.567395, 11.08139, 12.63369, 11.75156, 10.70997, 10.87275, 12.05752, 
    12.47425, 10.39009, 8.150321, 8.087931, 8.692059, 6.059055, 4.573244, 
    3.363755,
  5.095816, 6.669696, 5.48365, 6.68114, 5.581913, 4.654222, 5.635038, 
    3.970187, 2.822906, 2.001362, 2.228679, 3.22207, 4.087158, 3.421025, 
    1.853695,
  8.901944, 9.727968, 9.809859, 9.247342, 7.05416, 6.200647, 7.113941, 
    5.616723, 4.290644, 3.560037, 3.459509, 3.277899, 4.367136, 3.672973, 
    2.651763,
  11.78589, 11.55759, 10.52633, 8.44801, 5.23056, 3.177397, 3.389716, 
    2.685423, 2.528389, 3.13956, 3.811212, 4.419418, 4.641477, 5.053554, 
    3.96506,
  10.46747, 9.758495, 8.286391, 6.506525, 4.470928, 2.521685, 1.607154, 
    2.395563, 1.769274, 2.3436, 3.154191, 4.202782, 5.124385, 5.318207, 
    4.902085,
  6.842549, 5.531592, 4.41431, 3.797505, 3.521644, 3.275235, 3.379689, 
    2.056691, 1.650301, 1.720141, 2.980837, 3.81841, 5.237499, 5.746255, 
    6.176231,
  3.300912, 3.601396, 3.945282, 4.438937, 5.157836, 6.108057, 7.313029, 
    8.219937, 5.837998, 3.944988, 3.160258, 3.476887, 4.337955, 4.928586, 
    5.687095,
  3.242043, 4.048459, 4.761926, 5.840171, 7.247582, 8.481062, 9.871485, 
    10.74615, 9.831508, 8.355762, 6.278503, 3.880922, 3.668633, 4.827628, 
    6.072401,
  3.911315, 5.446394, 6.135077, 7.336526, 8.893971, 10.16903, 11.4873, 
    11.54181, 11.05684, 9.739491, 7.462476, 4.661253, 4.179734, 5.949833, 
    6.592796,
  5.195327, 6.331345, 6.641488, 7.809633, 9.533514, 9.836067, 9.924506, 
    8.603547, 8.11933, 8.395448, 7.311809, 5.270021, 5.671714, 7.478117, 
    6.129735,
  6.311141, 6.944431, 5.892725, 7.344551, 8.087946, 6.213342, 4.960057, 
    5.310446, 5.996823, 5.383107, 5.033202, 6.466913, 7.701811, 7.604761, 
    5.347944,
  7.028694, 10.64195, 10.9291, 13.6614, 12.8978, 10.70429, 12.70907, 
    12.19083, 10.7371, 7.842993, 6.593657, 5.661095, 5.091051, 5.297849, 
    5.72447,
  8.438213, 9.715081, 11.39983, 12.54454, 9.745272, 9.310986, 11.43436, 
    11.52899, 11.41173, 9.789445, 8.594566, 7.940831, 6.157727, 4.074429, 
    4.760899,
  9.922235, 10.57897, 10.56689, 10.66299, 9.072794, 7.591312, 8.048326, 
    8.605666, 9.230232, 9.94186, 9.779834, 8.507111, 6.609456, 4.493724, 
    4.9933,
  10.27023, 12.52916, 13.92043, 13.91512, 11.66969, 8.380016, 6.751686, 
    7.427485, 8.613161, 7.274038, 7.999055, 7.497152, 6.626199, 4.741838, 
    5.314224,
  8.085166, 9.484995, 11.09851, 11.95785, 11.88345, 10.24445, 6.833245, 
    5.152062, 5.458782, 5.811602, 7.727582, 7.004285, 6.429543, 5.479308, 
    5.140218,
  6.490534, 7.455637, 8.094666, 8.434374, 8.293175, 8.207557, 6.920693, 
    5.35784, 5.165458, 5.099389, 5.2632, 6.002999, 5.170694, 5.234885, 
    3.917954,
  5.395487, 5.991727, 6.291533, 6.897727, 6.625959, 5.662983, 5.361573, 
    5.884772, 5.825631, 6.869003, 6.617472, 5.23145, 3.809045, 4.177136, 
    4.775024,
  4.411446, 4.622979, 5.089219, 6.005301, 6.175967, 5.611557, 4.310242, 
    3.889102, 4.910666, 6.230625, 6.164032, 4.668979, 3.36277, 4.515412, 
    7.741251,
  3.661052, 3.461867, 4.132383, 5.367166, 6.022191, 6.083495, 5.300116, 
    4.208152, 3.47782, 4.474551, 5.445365, 4.920897, 4.594382, 6.796452, 
    7.656184,
  2.901376, 3.045726, 3.959919, 5.247986, 6.168332, 6.725642, 6.698537, 
    6.159797, 5.082872, 4.436319, 4.938486, 5.820471, 6.154412, 6.999577, 
    6.457168,
  7.213525, 8.368214, 6.207285, 6.471536, 5.5265, 4.581683, 6.073585, 
    7.916316, 8.55278, 8.180918, 9.709243, 11.18131, 11.15084, 10.22952, 
    9.208579,
  7.307653, 6.52938, 5.935091, 5.336448, 4.287819, 4.468304, 6.595137, 
    9.020411, 9.658677, 8.901062, 10.11771, 13.23498, 13.93829, 9.81917, 
    8.734571,
  4.684958, 4.507169, 4.727111, 4.960705, 4.333033, 4.535334, 7.3329, 
    7.996437, 7.485653, 8.423338, 11.0934, 13.37947, 12.56797, 11.07544, 
    7.594855,
  2.932611, 3.030916, 3.380894, 4.791726, 4.949446, 4.889506, 5.850035, 
    6.493715, 7.623352, 9.80025, 11.23213, 11.24865, 9.681664, 7.990447, 
    5.289001,
  2.690071, 2.496079, 3.280641, 4.539895, 5.309381, 5.712247, 5.144096, 
    4.00531, 5.819771, 8.496035, 11.65303, 10.00358, 7.316319, 6.457363, 
    6.53884,
  3.156308, 2.413141, 2.971916, 4.058523, 5.391058, 5.619038, 4.602715, 
    4.415654, 5.303369, 6.669967, 6.907678, 8.885803, 9.823861, 9.852771, 
    9.708825,
  2.921088, 1.852051, 2.363204, 4.268739, 5.102563, 4.28224, 3.598276, 
    4.626799, 6.172086, 7.391205, 6.815008, 7.633138, 9.537362, 10.88069, 
    11.48498,
  1.54109, 1.457306, 2.604942, 4.058218, 4.219053, 3.476736, 2.761937, 
    3.501129, 5.00721, 5.951344, 5.783169, 6.582488, 8.441476, 9.743121, 
    10.08804,
  1.882925, 1.757863, 2.513991, 3.426818, 3.472221, 3.193777, 2.985902, 
    3.457291, 4.342843, 5.15292, 5.270474, 5.882341, 7.142393, 7.977903, 
    8.18788,
  3.150651, 2.271961, 2.949041, 3.585849, 3.778373, 3.69475, 3.436255, 
    3.128183, 3.178876, 3.022184, 3.502244, 5.391356, 6.07242, 7.026118, 
    7.804147,
  4.849519, 6.697682, 6.247329, 7.844195, 6.757779, 7.331517, 9.636107, 
    9.473237, 7.62007, 5.230213, 4.574164, 4.151122, 4.067165, 4.657979, 
    5.489256,
  12.03947, 7.935115, 9.070918, 8.839728, 6.868136, 6.909606, 8.512488, 
    8.693694, 7.63705, 6.16502, 5.101448, 5.163026, 4.885547, 4.304946, 
    5.594584,
  14.53053, 12.98183, 10.20273, 9.444815, 7.832664, 7.142177, 7.293772, 
    7.86096, 7.616495, 6.173853, 5.316803, 4.740098, 4.764718, 5.787791, 
    5.796064,
  12.29752, 13.03901, 12.15689, 10.06677, 8.650727, 7.275253, 6.502321, 
    6.204388, 5.800838, 4.506689, 4.690324, 4.136286, 5.081362, 6.041972, 
    4.721054,
  9.298114, 10.3285, 10.64142, 9.63623, 7.985795, 6.528892, 6.297173, 
    4.724793, 3.268876, 3.17347, 3.890576, 3.406426, 4.683069, 5.669099, 
    5.173812,
  6.72336, 7.784155, 7.937356, 7.329429, 6.82881, 6.000018, 4.71829, 
    4.506767, 3.74256, 3.263551, 2.363359, 2.445959, 3.971004, 4.437923, 
    4.595152,
  5.255044, 6.349622, 5.882463, 5.37505, 5.283039, 5.14339, 4.823349, 
    4.542672, 4.195524, 3.793675, 2.53326, 1.956472, 2.882977, 3.28725, 
    3.975866,
  4.721154, 4.806427, 3.912508, 3.955722, 3.989755, 4.011432, 3.786649, 
    3.39777, 3.173409, 3.367092, 2.346022, 2.070395, 2.601384, 2.541119, 
    3.085972,
  4.264127, 3.196545, 2.383366, 2.449608, 2.538494, 2.868284, 2.68791, 
    2.142464, 2.258997, 2.740186, 2.425166, 2.078836, 2.275029, 2.387333, 
    2.83533,
  2.689933, 1.713213, 1.657744, 1.532416, 1.649835, 1.847466, 1.9799, 
    1.759528, 1.355135, 1.077939, 1.166522, 1.705947, 2.335178, 3.272196, 
    4.617418,
  5.446392, 5.238118, 4.416406, 3.869411, 2.867603, 2.750278, 4.995563, 
    7.253987, 7.080687, 5.707461, 6.019893, 6.922927, 6.521385, 4.517231, 
    2.42585,
  8.829627, 6.592779, 5.556293, 4.693962, 2.401077, 1.823459, 3.460289, 
    5.753863, 6.991104, 6.460632, 6.761354, 8.549068, 8.443936, 4.585291, 
    2.597812,
  9.535536, 8.930303, 5.797768, 4.726174, 3.317416, 2.805788, 1.857745, 
    3.369798, 6.886041, 8.264245, 8.651887, 9.490877, 8.820193, 5.758525, 
    3.37664,
  9.73194, 10.08341, 8.793593, 4.719197, 4.636816, 4.817885, 3.926577, 
    3.613769, 3.868354, 6.807208, 8.917513, 9.317327, 8.037491, 5.502522, 
    3.351651,
  9.491121, 10.43446, 10.52185, 8.492375, 4.807645, 5.720863, 7.133018, 
    6.056583, 4.13975, 4.658035, 8.554315, 9.571018, 8.278092, 5.993183, 
    3.86116,
  8.807062, 9.713847, 10.75879, 10.16564, 7.986231, 4.80788, 6.920769, 
    9.270761, 7.414253, 7.182706, 7.321981, 9.657363, 8.283387, 6.187466, 
    4.500975,
  7.775854, 8.743905, 9.739348, 10.18149, 9.5331, 7.578257, 5.524167, 
    7.100517, 9.44803, 10.21691, 10.17731, 9.770988, 8.110232, 6.351974, 
    5.027245,
  6.24199, 7.432822, 8.577971, 9.462882, 9.655067, 8.552699, 7.395772, 
    9.170116, 10.94244, 10.94289, 10.52888, 9.482881, 7.523209, 6.123614, 
    4.842787,
  4.160594, 5.611945, 6.947287, 8.292248, 9.189067, 9.034992, 8.640772, 
    9.760755, 10.94089, 10.72233, 9.881694, 8.29712, 6.532421, 5.407978, 
    4.359436,
  1.912566, 3.561745, 5.399423, 6.883632, 8.22743, 8.955896, 9.462241, 
    9.786531, 8.645732, 6.79964, 6.434638, 6.793284, 5.560605, 4.897193, 
    4.556606,
  6.894981, 8.477451, 7.408788, 7.191946, 5.275501, 2.574337, 4.469018, 
    5.878564, 5.647833, 4.325972, 4.390372, 4.272595, 4.502282, 4.380605, 
    4.487089,
  8.951414, 9.161383, 9.77741, 8.445866, 5.092245, 3.742932, 3.769081, 
    3.734448, 4.863478, 4.206432, 4.356809, 5.540048, 6.025453, 4.739902, 
    4.915941,
  8.198508, 8.672601, 9.080655, 8.928103, 6.283056, 3.591544, 3.952872, 
    2.739358, 3.864243, 4.376059, 4.41196, 5.341108, 6.678141, 6.772247, 
    6.353806,
  7.292546, 7.775356, 8.177082, 8.49297, 7.509329, 4.384715, 2.931775, 
    4.090069, 4.119691, 2.66319, 3.831117, 4.485607, 5.563385, 6.456314, 
    6.880931,
  5.668055, 6.55447, 7.273026, 7.498227, 6.913019, 5.644059, 3.719604, 
    2.202728, 2.70635, 2.020335, 3.007312, 3.784902, 5.012343, 6.931277, 
    8.580631,
  4.166437, 5.169961, 6.304863, 6.972683, 6.809396, 5.933918, 5.161427, 
    5.305657, 3.904666, 2.427546, 2.062012, 2.934891, 4.165476, 6.710786, 
    8.372405,
  4.273325, 4.379354, 5.402464, 6.57966, 7.024457, 6.448889, 6.382019, 
    6.453076, 5.943045, 5.575696, 4.61981, 3.646059, 4.691202, 6.697053, 
    8.548772,
  4.769485, 4.067357, 5.178155, 6.496868, 6.996431, 6.849244, 6.663252, 
    7.170614, 7.788753, 7.571014, 6.569674, 6.292196, 6.946683, 7.959548, 
    9.354668,
  3.942078, 3.425509, 4.633104, 5.811302, 6.56644, 6.897014, 7.2482, 
    6.673256, 6.983768, 7.253531, 8.14058, 8.952731, 9.252007, 9.921359, 
    9.98681,
  3.08034, 2.620667, 4.021649, 5.393831, 6.443192, 7.305288, 8.045398, 
    7.11769, 5.854347, 5.303143, 6.875795, 10.10259, 10.491, 11.10038, 
    10.08122,
  13.13416, 13.22418, 8.946644, 8.746314, 7.269735, 6.040694, 7.814629, 
    8.381728, 7.554328, 5.681574, 5.028837, 4.255634, 4.155594, 3.3015, 
    3.68283,
  17.06646, 16.42697, 13.03458, 9.449042, 6.431849, 5.799402, 7.160745, 
    7.291222, 6.429863, 4.964789, 4.733939, 5.222225, 5.205321, 3.457781, 
    3.556006,
  15.16313, 16.4949, 15.82368, 12.00936, 7.808858, 5.422373, 5.7002, 
    7.435496, 8.045794, 6.637553, 5.095074, 4.613773, 5.013182, 4.290956, 
    4.055051,
  12.62999, 14.17358, 15.19056, 14.49618, 10.79091, 6.275465, 5.194381, 
    7.217674, 9.435438, 7.306308, 6.129875, 4.278567, 3.264741, 3.17085, 
    4.112574,
  9.07763, 10.81748, 12.49263, 13.32673, 12.32681, 9.335169, 6.825334, 
    5.803777, 3.969116, 3.984956, 5.954625, 5.091694, 3.623789, 3.022007, 
    4.492898,
  5.695218, 6.761245, 8.778517, 10.42833, 11.20617, 10.84186, 9.18921, 
    7.177787, 4.582901, 3.814633, 3.96455, 5.47993, 4.307748, 3.224613, 
    3.437693,
  4.233797, 3.418757, 4.253102, 6.537618, 8.188684, 9.083473, 9.186789, 
    8.605873, 7.502001, 6.084728, 5.307794, 4.825275, 4.152715, 3.609135, 
    3.285234,
  4.88066, 2.951183, 2.628366, 3.154004, 4.689366, 5.853837, 6.445164, 
    6.653204, 6.393076, 5.941787, 5.628731, 5.035728, 4.167665, 3.665191, 
    3.608237,
  5.391673, 3.975232, 3.108789, 2.872565, 2.53288, 3.500651, 4.462963, 
    5.415377, 5.759231, 5.317258, 4.875828, 4.777114, 4.748961, 4.404317, 
    3.842753,
  4.690629, 4.181886, 4.049606, 4.03226, 3.596185, 2.926877, 3.215047, 
    3.884419, 3.974143, 3.313015, 3.89499, 5.284369, 5.465339, 5.464512, 
    5.110958,
  8.82373, 4.502766, 6.782233, 7.112494, 4.024956, 3.360124, 6.900246, 
    8.948024, 8.700441, 7.721816, 7.282036, 6.5457, 6.164057, 4.63747, 
    3.912602,
  15.23502, 5.500703, 6.366843, 6.857337, 3.796307, 2.920209, 6.036795, 
    8.295141, 8.429219, 7.26784, 7.253067, 7.649803, 7.455578, 4.67877, 
    3.934631,
  17.06556, 10.31511, 4.947399, 4.952072, 3.62499, 3.715375, 3.805992, 
    6.266484, 8.585501, 8.499972, 8.299003, 8.466105, 7.914664, 6.51083, 
    4.687759,
  16.74542, 14.73749, 7.795951, 3.981294, 3.782686, 4.936934, 5.463252, 
    5.080249, 4.954477, 5.776124, 7.665699, 7.893254, 7.179914, 5.941054, 
    4.688737,
  15.22263, 15.94014, 13.20772, 7.4376, 3.575706, 5.870448, 8.185777, 
    7.784316, 3.846896, 2.754889, 6.243372, 7.437523, 6.921732, 6.024578, 
    5.585401,
  12.38815, 14.60624, 15.24258, 12.35792, 6.899786, 4.784735, 7.511741, 
    8.843608, 6.395909, 4.797386, 5.127626, 7.436916, 7.252568, 6.175236, 
    4.974196,
  10.33969, 12.0183, 13.62376, 14.20562, 11.84437, 6.987851, 5.783485, 
    6.272863, 6.939361, 7.615171, 7.968435, 8.116656, 7.739203, 6.944548, 
    5.695306,
  8.484245, 9.190569, 10.72125, 12.69333, 13.43422, 10.8542, 7.366512, 
    7.937701, 8.285395, 8.400275, 8.533827, 8.449413, 8.012759, 7.424284, 
    6.345759,
  6.744414, 6.040021, 6.832954, 9.098031, 11.69339, 12.2778, 10.0245, 
    8.269794, 8.296827, 8.26159, 8.525517, 8.526464, 8.006399, 7.475688, 
    6.250872,
  5.048091, 3.947186, 3.939659, 5.257596, 8.014087, 10.16755, 10.64253, 
    9.12299, 6.915665, 5.478219, 6.151503, 7.790438, 7.134297, 6.560935, 
    5.363628,
  9.155606, 7.062159, 5.457249, 7.744963, 5.40996, 2.902866, 1.851812, 
    5.693299, 3.32926, 5.293374, 7.38138, 7.128666, 6.889565, 5.653759, 
    5.612637,
  13.03429, 7.447168, 3.962338, 7.71385, 5.565305, 3.138498, 2.749649, 
    4.599032, 4.087406, 3.999299, 7.799711, 8.344926, 7.814964, 5.378044, 
    4.849393,
  13.07407, 9.109155, 2.23417, 6.885345, 5.854567, 3.074416, 2.148866, 
    3.134564, 3.072026, 6.52974, 9.236265, 9.166161, 8.133965, 6.434314, 
    4.341554,
  13.07491, 10.90151, 3.298849, 5.430676, 6.086651, 4.751099, 2.359554, 
    1.86496, 3.972288, 5.366837, 8.86335, 8.893727, 7.961802, 6.30617, 
    4.412956,
  12.67781, 12.26396, 7.638721, 2.591517, 5.584771, 5.358903, 4.740006, 
    3.669361, 2.703204, 2.950822, 7.690864, 8.546163, 7.9704, 6.484456, 
    4.951147,
  10.64942, 12.47238, 10.56213, 4.754796, 3.966083, 5.873827, 6.291904, 
    6.330359, 3.907019, 3.620124, 5.26643, 8.39141, 8.022913, 6.668335, 
    5.052404,
  9.561071, 11.68722, 11.50898, 9.213329, 3.578922, 5.842888, 6.918415, 
    5.754853, 4.870613, 5.390426, 7.137321, 8.603675, 8.377584, 7.2376, 
    5.702349,
  8.024294, 10.24938, 11.02248, 11.18165, 8.934473, 3.878348, 7.542635, 
    8.161186, 7.438506, 6.466627, 6.645336, 8.093866, 8.356019, 7.591771, 
    6.252765,
  5.91396, 7.799906, 9.296934, 11.01853, 11.6371, 7.518558, 5.612966, 
    8.278048, 7.853463, 6.636777, 6.402252, 7.395855, 7.998558, 7.718518, 
    6.586434,
  3.881672, 5.077774, 6.857814, 9.522912, 12.1377, 12.05439, 6.258943, 
    7.195383, 7.176999, 5.268175, 5.142565, 7.10473, 7.443623, 7.689149, 
    6.916959,
  5.164035, 7.932854, 7.006207, 8.409231, 7.152252, 5.168714, 5.020635, 
    5.35068, 6.304421, 4.922925, 4.765639, 4.675841, 4.71022, 4.507028, 
    4.885571,
  7.776678, 8.927336, 8.155127, 7.927776, 5.564947, 4.229182, 4.897328, 
    5.435915, 6.352144, 4.989834, 5.147924, 5.281723, 5.367083, 4.179287, 
    4.340236,
  8.571608, 9.326718, 7.55374, 6.754242, 5.206567, 3.384226, 3.497126, 
    5.409825, 5.170029, 5.708859, 5.629691, 5.936276, 5.705239, 4.802189, 
    3.657056,
  8.823874, 9.159299, 6.795011, 5.529991, 5.270615, 4.367245, 2.356508, 
    2.350541, 3.333331, 5.068872, 6.133062, 6.08517, 5.315892, 4.894925, 
    3.829165,
  8.437321, 9.221612, 6.923173, 4.229639, 4.059733, 3.644211, 2.933925, 
    2.674262, 2.552289, 2.792619, 6.577591, 6.069457, 5.118259, 5.074435, 
    5.048997,
  7.080398, 9.091602, 7.683642, 3.61771, 3.455913, 3.167454, 3.29459, 
    4.122608, 3.784014, 4.34095, 5.018593, 6.277502, 5.246156, 4.99191, 
    5.416875,
  5.808038, 8.713177, 8.437987, 4.253547, 2.306669, 2.497292, 2.786858, 
    4.236498, 4.92165, 7.300268, 7.761946, 7.090953, 5.784944, 5.254837, 
    5.260636,
  4.88026, 7.984374, 9.057528, 6.440904, 2.577509, 2.415875, 2.920164, 
    3.402395, 5.11643, 7.312286, 7.804193, 7.256716, 6.224021, 5.397762, 
    4.714524,
  3.89826, 6.296294, 8.597513, 8.642954, 5.016088, 2.770928, 2.33588, 
    3.408221, 4.326931, 6.477668, 7.031742, 6.982741, 6.405489, 5.611956, 
    4.480409,
  3.120549, 4.259376, 6.966366, 9.706118, 9.299993, 5.747087, 2.859148, 
    3.084452, 4.410027, 4.308087, 4.893874, 6.457248, 6.123126, 5.773396, 
    4.826194,
  2.208369, 2.613814, 2.531166, 4.468501, 4.687168, 3.841121, 4.91228, 
    5.891494, 5.7616, 5.317498, 6.396518, 4.635158, 2.873797, 4.465592, 
    4.835207,
  3.746592, 3.840329, 3.223744, 4.283708, 3.905568, 3.565547, 4.974542, 
    5.810862, 6.101556, 5.582231, 6.118119, 4.286261, 3.770484, 4.392477, 
    5.000389,
  3.966678, 4.02202, 3.943467, 4.148715, 3.560373, 3.311895, 4.269326, 
    4.49086, 4.682515, 5.364942, 5.755418, 2.915123, 4.348617, 5.820222, 
    5.246014,
  3.812805, 4.048143, 4.121704, 4.560594, 4.725406, 4.577282, 3.679518, 
    4.197295, 4.546856, 4.970923, 4.395502, 2.046375, 4.533478, 6.275774, 
    5.53631,
  4.013972, 3.946543, 4.581974, 5.698781, 6.118657, 6.278297, 5.629612, 
    3.14497, 3.163141, 3.515553, 3.876245, 2.137939, 4.31838, 6.830602, 
    6.860566,
  4.001795, 4.091582, 5.840725, 6.979544, 7.348427, 7.345922, 7.053062, 
    6.793381, 4.295692, 3.021831, 2.906549, 2.07416, 3.906929, 6.809902, 
    6.972611,
  4.537658, 5.682896, 7.09245, 7.692375, 7.907038, 7.528639, 7.368187, 
    6.341737, 5.178372, 4.03298, 3.751572, 2.150457, 4.360098, 6.866338, 
    7.226377,
  6.041417, 6.974679, 7.594732, 7.581002, 7.406912, 7.457977, 7.441743, 
    7.487858, 6.753515, 4.76974, 3.651074, 2.538024, 4.978662, 7.195449, 
    7.078366,
  7.029872, 6.689198, 6.543024, 7.349446, 6.455606, 7.249287, 7.837016, 
    7.502401, 6.709147, 5.019769, 4.214327, 3.253537, 5.622864, 7.59697, 
    6.878005,
  7.22835, 5.732898, 5.366126, 7.89891, 7.251448, 6.150222, 7.93618, 
    8.183071, 6.432843, 3.863955, 3.405776, 3.814185, 5.949995, 7.700608, 
    6.633212,
  3.734597, 4.571475, 4.052641, 5.193661, 5.197143, 5.556209, 7.808095, 
    8.620811, 8.43556, 6.726915, 6.296112, 5.254887, 4.780618, 5.002146, 
    5.651872,
  4.773776, 4.326461, 2.80522, 3.256109, 3.237171, 3.805671, 6.005261, 
    7.783999, 8.994744, 8.812435, 7.419776, 5.718769, 5.408138, 4.003829, 
    4.605845,
  4.735138, 5.110541, 3.013344, 1.461923, 2.162066, 2.409953, 4.075742, 
    4.804381, 6.760654, 9.581813, 10.13194, 6.908973, 5.488644, 4.635751, 
    3.546661,
  3.161077, 4.528432, 4.38562, 2.988048, 1.416, 1.669374, 2.087781, 3.86212, 
    5.859931, 8.663264, 10.37311, 7.881028, 5.01109, 4.720503, 3.563085,
  1.534946, 2.26097, 4.231514, 4.618116, 3.898331, 2.89699, 2.562579, 
    1.816852, 3.071601, 5.058673, 8.538294, 8.901331, 5.068403, 4.608878, 
    4.495711,
  2.704643, 3.461367, 4.519759, 5.448011, 5.959195, 6.087643, 5.295117, 
    4.124422, 2.869802, 2.790856, 4.802467, 8.296811, 5.190074, 4.481622, 
    4.464855,
  5.111732, 5.028253, 5.612343, 6.238102, 7.012059, 7.582553, 7.46891, 
    6.496912, 4.838844, 3.617757, 4.266809, 6.367482, 5.143775, 4.17275, 
    4.392303,
  5.141289, 5.237875, 6.022956, 6.950103, 7.65423, 8.150665, 8.349325, 
    8.408996, 7.504627, 5.810707, 4.23905, 4.395581, 4.349041, 3.846516, 
    4.210544,
  5.45635, 6.064852, 6.604811, 7.450222, 7.991413, 8.314653, 8.670855, 
    8.763239, 8.277762, 7.202728, 5.659241, 3.967233, 3.373574, 3.738333, 
    4.005767,
  6.41678, 7.372137, 7.649807, 7.935794, 7.995557, 8.299212, 8.868142, 
    9.012712, 7.858825, 5.936742, 5.02608, 4.676367, 3.10219, 3.878608, 
    3.998158 ;

 sftlf =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 ts =
  261.4232, 272.5475, 265.6495, 272.4573, 269.0145, 261.5891, 265.9818, 
    266.0406, 265.0528, 248.9288, 251.1606, 254.6861, 246.4969, 248.7467, 
    236.9789,
  273.9857, 274.3366, 273.8667, 273.251, 262.0461, 259.3752, 268.0388, 
    267.6493, 267.2528, 261.5524, 253.6797, 261.9098, 261.2255, 243.566, 
    237.404,
  274.549, 274.3253, 274.1998, 273.7679, 266.4384, 246.4558, 265.5848, 
    268.087, 269.0542, 265.7857, 264.2489, 264.5054, 263.9605, 262.2203, 
    252.6757,
  275.2407, 274.548, 274.3043, 273.9989, 273.6055, 266.5992, 241.8416, 
    259.9698, 270.1733, 266.5981, 265.2796, 265.0668, 264.6185, 263.4366, 
    258.1172,
  275.598, 274.8677, 274.3722, 274.0643, 273.6554, 273.1092, 268.7558, 
    240.5218, 245.7056, 254.8214, 264.954, 265.1902, 264.7043, 264.1416, 
    263.6872,
  275.8509, 275.1342, 274.492, 274.0281, 273.6563, 273.1708, 272.5679, 
    271.3146, 262.1692, 259.521, 257.3068, 265.1455, 264.8419, 264.7994, 
    264.5615,
  276.2159, 275.3926, 274.6307, 274.0139, 273.5748, 273.1279, 272.6599, 
    272.2452, 271.8737, 271.8689, 269.0397, 265.0277, 264.8685, 264.9608, 
    264.8604,
  276.4522, 275.5732, 274.7629, 274.0305, 273.4726, 273.0077, 272.5783, 
    272.2553, 271.9786, 271.9466, 270.1411, 265.6964, 265.1457, 265.4391, 
    265.4749,
  276.076, 275.4014, 274.6709, 273.9366, 273.3167, 272.8689, 272.4659, 
    272.192, 272.1202, 271.609, 270.9261, 266.1559, 265.1629, 265.1784, 
    264.4437,
  275.1428, 274.4504, 274.0824, 273.6014, 273.04, 272.6216, 272.3374, 
    271.7111, 269.3892, 261.0533, 264.7556, 266.5723, 265.1909, 265.252, 
    264.9557,
  260.9113, 272.2013, 264.2051, 272.1252, 264.4835, 258.6393, 260.5332, 
    260.2623, 259.5305, 251.6197, 253.2786, 255.6495, 252.4703, 252.1744, 
    246.4348,
  273.7076, 274.2257, 273.8093, 273.0449, 260.6055, 256.1472, 261.8936, 
    261.2067, 260.5548, 258.2043, 254.7179, 258.2436, 257.6117, 247.8571, 
    244.5694,
  274.3864, 274.1931, 274.1149, 273.6838, 265.6578, 243.3604, 261.3607, 
    262.2855, 262.1299, 260.058, 259.6718, 259.3856, 258.4526, 257.9774, 
    251.9971,
  275.0886, 274.4305, 274.1885, 273.8976, 273.556, 266.2726, 244.3935, 
    259.4481, 263.0703, 260.6169, 260.1694, 259.7016, 258.9276, 257.6768, 
    254.7654,
  275.4106, 274.7136, 274.2326, 273.9288, 273.5631, 272.934, 268.6429, 
    247.075, 247.5125, 255.497, 260.1198, 259.8994, 259.2355, 258.479, 
    258.1149,
  275.7095, 274.9878, 274.3295, 273.8784, 273.5259, 273.0885, 272.3579, 
    271.2177, 264.4097, 262.9635, 257.2044, 260.3738, 259.7642, 259.4067, 
    259.0878,
  276.0925, 275.2771, 274.483, 273.8482, 273.4282, 273.0031, 272.5526, 
    272.0751, 271.6267, 271.6322, 265.3049, 260.7178, 260.1572, 259.9277, 
    259.4501,
  276.3787, 275.4912, 274.6779, 273.9168, 273.352, 272.8666, 272.4411, 
    272.1112, 271.8094, 271.6971, 267.1726, 261.1601, 260.6808, 260.5198, 
    259.9947,
  276.0173, 275.3458, 274.6049, 273.8161, 273.1679, 272.6839, 272.3007, 
    272.0397, 271.9105, 271.4145, 268.4091, 261.677, 261.1417, 260.8136, 
    259.8739,
  275.0603, 274.3744, 273.9991, 273.4661, 272.8647, 272.4332, 272.1444, 
    271.5997, 269.7004, 263.2733, 264.592, 262.1345, 261.5235, 261.2768, 
    260.2748,
  266.9581, 272.4611, 263.8467, 271.8894, 264.7606, 259.7199, 261.139, 
    261.0038, 260.9916, 252.8575, 252.7801, 252.9339, 250.2005, 251.7315, 
    246.3572,
  273.6947, 274.1797, 273.7932, 272.927, 259.5136, 257.1024, 262.884, 
    262.2315, 262.2334, 259.1941, 254.1138, 255.872, 257.2929, 248.7141, 
    245.2556,
  274.3526, 274.1608, 274.0523, 273.6401, 266.582, 248.0284, 262.4416, 
    263.3374, 263.0574, 260.3058, 258.2545, 257.4529, 257.6061, 259.5309, 
    253.6783,
  275.0125, 274.373, 274.1254, 273.8594, 273.5971, 267.4239, 245.8319, 
    260.0533, 262.7541, 260.4036, 258.7846, 258.2536, 258.2664, 257.8349, 
    257.0465,
  275.3269, 274.6401, 274.1682, 273.8805, 273.5484, 273.0114, 269.2608, 
    247.2702, 251.175, 257.9452, 259.4659, 259.2844, 258.9626, 258.5599, 
    258.5129,
  275.6413, 274.9382, 274.2602, 273.8158, 273.4867, 273.0997, 272.5183, 
    271.2987, 265.9336, 265.646, 259.8548, 259.8284, 259.3519, 259.224, 
    258.9186,
  276.0531, 275.2315, 274.4219, 273.7866, 273.3915, 272.988, 272.5378, 
    272.0823, 271.6559, 271.479, 263.5905, 260.5712, 259.7262, 259.902, 
    259.7477,
  276.3444, 275.4417, 274.6267, 273.8831, 273.3414, 272.8773, 272.4042, 
    272.0865, 271.7866, 271.591, 264.9236, 261.0053, 260.3088, 260.7182, 
    259.5829,
  275.9795, 275.3147, 274.5796, 273.79, 273.1452, 272.6529, 272.2452, 
    271.9998, 271.8486, 271.2299, 265.9212, 261.2701, 260.9381, 260.4531, 
    258.7062,
  274.9955, 274.3195, 273.9604, 273.4071, 272.7852, 272.3469, 272.0625, 
    271.5429, 270.0785, 265.6929, 264.393, 261.4113, 261.4474, 260.308, 
    259.8017,
  268.2433, 272.5414, 266.413, 271.8187, 265.5292, 260.7764, 261.9235, 
    259.2482, 257.4232, 248.1523, 248.8481, 248.7672, 244.2604, 245.6659, 
    235.9377,
  273.5627, 274.1088, 273.7657, 272.8929, 258.7083, 256.8725, 264.2878, 
    262.0244, 259.8647, 256.2357, 250.5677, 252.3837, 254.0294, 242.0861, 
    236.8434,
  274.2689, 274.1042, 274.0269, 273.6133, 265.3709, 247.7682, 263.1978, 
    263.3817, 261.8015, 258.4598, 255.8, 253.3345, 253.3334, 256.3084, 
    249.8748,
  274.9724, 274.3317, 274.0931, 273.8428, 273.5976, 267.2036, 250.9528, 
    260.1742, 260.8491, 257.7421, 254.9741, 253.549, 253.8431, 254.812, 
    254.4188,
  275.2951, 274.616, 274.1387, 273.8532, 273.5339, 273.027, 269.6444, 
    251.7839, 252.139, 253.649, 254.3732, 254.2474, 254.99, 256.2798, 256.8486,
  275.6046, 274.9187, 274.2285, 273.7925, 273.4683, 273.1018, 272.5204, 
    271.0408, 263.5948, 262.9958, 255.6959, 255.4267, 256.0606, 256.9972, 
    256.0624,
  276.0326, 275.2077, 274.4032, 273.7736, 273.3885, 272.9814, 272.5187, 
    272.0536, 271.5334, 271.1066, 260.8328, 256.9967, 257.3243, 257.1219, 
    256.8154,
  276.3285, 275.412, 274.5975, 273.8758, 273.3459, 272.8961, 272.3749, 
    272.0553, 271.7337, 271.1598, 261.2251, 258.3658, 257.711, 257.518, 257.2,
  275.9539, 275.2995, 274.5721, 273.7888, 273.1504, 272.6853, 272.2274, 
    271.9639, 271.7912, 270.9352, 262.8768, 259.299, 258.0822, 258.2564, 
    257.5042,
  274.935, 274.2646, 273.935, 273.3792, 272.7463, 272.3162, 272.04, 271.4784, 
    270.1179, 264.9203, 261.7554, 259.5533, 259.2415, 258.597, 259.1073,
  267.4596, 272.5972, 268.3535, 271.8336, 265.3606, 262.1751, 261.6399, 
    256.3508, 254.6736, 246.9529, 244.2722, 246.7943, 241.833, 243.1037, 
    234.2209,
  273.4676, 274.0057, 273.7329, 272.7888, 262.9688, 261.3247, 260.2725, 
    257.2383, 255.5462, 253.543, 247.2299, 252.2016, 255.3134, 239.4828, 
    232.8709,
  274.2053, 274.0147, 273.9927, 273.5595, 268.4596, 255.294, 260.3916, 
    258.8813, 256.6668, 254.9126, 254.6928, 253.7459, 255.1882, 257.3857, 
    247.0334,
  274.9181, 274.2754, 274.055, 273.8246, 273.5725, 268.175, 252.2421, 
    257.2417, 257.3658, 255.7791, 254.2335, 253.9239, 255.095, 255.6094, 
    252.3885,
  275.2532, 274.5909, 274.1123, 273.8397, 273.516, 273.1097, 268.9947, 
    248.4467, 246.8338, 251.4336, 253.6988, 254.6718, 255.7691, 256.8853, 
    258.1474,
  275.56, 274.8989, 274.2181, 273.7846, 273.4538, 273.094, 272.5924, 
    270.4323, 261.851, 260.6966, 255.0816, 255.4867, 256.4041, 257.5228, 
    257.7222,
  275.9943, 275.196, 274.4126, 273.7645, 273.3781, 272.9613, 272.5406, 
    272.0344, 270.9618, 270.5199, 260.7969, 256.4236, 256.9974, 257.8633, 
    258.1747,
  276.3141, 275.4146, 274.5933, 273.8651, 273.3329, 272.8994, 272.37, 
    272.0236, 271.6773, 270.6799, 259.509, 257.1565, 257.7242, 258.3683, 
    258.352,
  275.9433, 275.3134, 274.5847, 273.7634, 273.1164, 272.7312, 272.2384, 
    271.9082, 271.7235, 270.5957, 260.6623, 257.8233, 258.2107, 258.8047, 
    258.9296,
  274.9331, 274.2496, 273.9149, 273.3295, 272.726, 272.335, 272.0378, 
    271.4134, 269.8429, 263.5536, 259.6741, 258.383, 258.7697, 259.8268, 
    261.6818,
  263.9435, 272.2047, 266.3773, 271.6471, 263.2143, 260.9157, 261.723, 
    257.9201, 255.3701, 244.3055, 240.6227, 247.4505, 243.9388, 245.6341, 
    237.3573,
  273.3396, 273.8849, 273.6863, 272.8015, 262.4869, 261.1938, 261.6315, 
    257.4351, 254.8957, 252.3257, 244.3177, 254.1342, 257.2939, 240.5549, 
    236.5019,
  274.1534, 273.9449, 273.9348, 273.4992, 268.8662, 257.4631, 259.9808, 
    257.7526, 255.0571, 255.3475, 255.1752, 255.8233, 257.6718, 258.153, 
    247.5691,
  274.8667, 274.2186, 273.9969, 273.8016, 273.5594, 268.4082, 252.6995, 
    254.7995, 255.4984, 254.9664, 254.6343, 255.5012, 256.9476, 257.287, 
    253.1065,
  275.1965, 274.5468, 274.0687, 273.8174, 273.5121, 273.1667, 268.3338, 
    246.3331, 242.5652, 248.5963, 253.6851, 255.833, 257.4677, 258.3761, 
    259.1075,
  275.502, 274.8462, 274.1916, 273.7732, 273.4538, 273.0958, 272.6004, 
    269.7813, 260.9453, 258.4045, 253.2261, 256.8468, 258.0024, 259.3187, 
    259.8003,
  275.9421, 275.1591, 274.3956, 273.7387, 273.3783, 272.9633, 272.5465, 
    271.9915, 270.2461, 269.3599, 261.2072, 257.9833, 258.5791, 259.6784, 
    260.682,
  276.2698, 275.3829, 274.5671, 273.8432, 273.344, 272.9125, 272.3591, 
    271.9674, 271.6112, 270.4501, 259.9236, 258.4246, 258.8052, 260.5119, 
    261.1411,
  275.9336, 275.3066, 274.5935, 273.7749, 273.1505, 272.7556, 272.2344, 
    271.8367, 271.6638, 270.3604, 260.4205, 258.6363, 259.6832, 261.2455, 
    261.9372,
  275.0149, 274.2575, 273.9263, 273.3412, 272.737, 272.339, 272.0338, 
    271.3848, 269.6542, 263.8236, 260.0703, 258.8664, 259.8386, 261.6104, 
    263.7567,
  261.1124, 271.8733, 264.5701, 270.7391, 257.687, 255.2397, 258.0868, 
    256.3057, 256.2793, 247.3473, 248.9675, 252.6294, 246.2282, 246.373, 
    240.419,
  273.1369, 273.7495, 273.605, 272.7885, 257.3758, 256.3075, 259.363, 
    257.1053, 256.443, 255.9084, 251.2973, 257.7324, 257.6642, 242.5402, 
    238.7871,
  274.1075, 273.884, 273.9063, 273.474, 266.3386, 253.5141, 258.2889, 
    257.5391, 256.8131, 257.5833, 257.5655, 258.5088, 259.106, 257.8298, 
    249.6864,
  274.8271, 274.1964, 273.9559, 273.7639, 273.4939, 267.7504, 253.0625, 
    252.3206, 256.235, 256.6241, 256.9484, 258.1416, 258.8394, 257.7557, 
    253.7147,
  275.146, 274.4969, 274.0324, 273.7665, 273.4544, 273.1153, 268.1027, 
    246.1869, 239.9875, 249.3446, 256.2171, 258.3426, 258.9175, 259.8886, 
    258.9174,
  275.5153, 274.7827, 274.1498, 273.7227, 273.4118, 273.0777, 272.5275, 
    270.0615, 259.7371, 257.1087, 253.2428, 258.6251, 260.1042, 260.7333, 
    259.7813,
  275.9653, 275.1094, 274.3459, 273.6947, 273.3437, 272.9526, 272.5456, 
    271.957, 270.1925, 268.6031, 262.1385, 259.0749, 260.4636, 260.9416, 
    260.596,
  276.2911, 275.3461, 274.5255, 273.8016, 273.3205, 272.9165, 272.3547, 
    271.9429, 271.555, 270.5832, 260.5206, 259.231, 260.5456, 261.6005, 
    261.3397,
  275.9615, 275.3074, 274.6109, 273.8112, 273.1952, 272.7687, 272.2258, 
    271.8155, 271.6118, 270.2993, 260.4783, 259.2056, 260.4858, 262.3375, 
    262.2982,
  275.0998, 274.2589, 273.9467, 273.388, 272.7543, 272.322, 272.0186, 
    271.4573, 270.0175, 263.6717, 260.1099, 259.4453, 260.5099, 262.3698, 
    263.1304,
  261.7363, 271.4237, 263.3221, 268.8239, 256.9417, 252.0104, 257.9299, 
    257.2326, 256.9525, 247.4311, 245.0631, 246.8502, 242.126, 243.3412, 
    237.716,
  273.0098, 273.6548, 273.5107, 272.5155, 254.5597, 249.4205, 258.5711, 
    258.3406, 257.7094, 256.1109, 248.7267, 254.0993, 254.4664, 240.2621, 
    236.7513,
  274.1129, 273.8542, 273.8855, 273.4256, 265.4718, 248.39, 256.1584, 
    258.8839, 258.6175, 258.2431, 256.9497, 256.6734, 256.3073, 255.8174, 
    249.2625,
  274.7974, 274.1876, 273.9321, 273.7369, 273.4415, 266.8122, 242.5681, 
    253.8942, 258.6292, 258.2465, 257.4656, 256.7981, 256.5521, 255.8676, 
    252.9954,
  275.1128, 274.474, 274.0123, 273.7248, 273.4187, 273.0749, 267.4781, 
    244.0155, 244.8339, 252.6437, 257.6479, 257.8631, 257.0428, 256.7134, 
    256.826,
  275.4903, 274.7397, 274.114, 273.6739, 273.3856, 273.0449, 272.429, 
    269.8653, 260.9554, 259.0914, 254.7075, 258.5045, 257.83, 258.235, 
    257.7079,
  275.9751, 275.1031, 274.3023, 273.6597, 273.3044, 272.9131, 272.4978, 
    271.8685, 269.9613, 268.0117, 261.843, 259.5562, 258.8282, 258.73, 
    258.1916,
  276.3077, 275.3453, 274.504, 273.7691, 273.285, 272.8698, 272.2964, 
    271.8938, 271.4991, 270.1426, 260.9374, 260.3817, 260.0012, 259.4552, 
    258.351,
  275.9885, 275.3087, 274.6245, 273.8289, 273.2027, 272.7344, 272.142, 
    271.7415, 271.5593, 269.5054, 260.5508, 260.5426, 260.4678, 259.9895, 
    259.1409,
  275.1982, 274.2737, 273.9579, 273.4156, 272.7361, 272.2618, 271.9321, 
    271.3716, 269.8225, 263.5882, 261.1229, 260.5834, 260.8812, 261.0603, 
    261.5252,
  263.0708, 270.7419, 261.5298, 265.5985, 256.0223, 253.1685, 254.4779, 
    253.0471, 252.969, 242.0873, 241.0491, 244.5164, 240.7443, 243.4241, 
    236.8141,
  272.8782, 273.54, 273.2657, 271.8618, 254.4479, 252.033, 256.17, 254.4057, 
    253.5008, 251.6497, 243.2083, 252.1838, 253.9379, 236.9551, 234.5235,
  274.0759, 273.799, 273.8455, 273.3594, 264.5103, 246.7874, 255.8831, 
    255.8812, 254.6382, 254.1717, 254.0794, 254.5702, 255.29, 255.3371, 
    247.4625,
  274.7646, 274.1438, 273.8929, 273.6977, 273.3279, 266.3121, 246.9043, 
    253.1799, 254.7043, 253.9121, 253.5221, 254.0724, 255.1887, 255.4147, 
    252.7348,
  275.0877, 274.4268, 273.9696, 273.6865, 273.3756, 272.9689, 267.2433, 
    246.9314, 243.9406, 248.9307, 253.6532, 254.7244, 255.7782, 256.3349, 
    256.9955,
  275.468, 274.7034, 274.072, 273.6322, 273.3365, 272.9896, 272.1694, 
    269.0132, 260.1767, 256.9154, 253.396, 255.632, 256.0714, 256.6968, 
    257.1712,
  275.9957, 275.0956, 274.2582, 273.6196, 273.2612, 272.8442, 272.4146, 
    271.655, 268.6841, 264.8691, 259.078, 256.8132, 256.3311, 257.0309, 
    257.7691,
  276.3198, 275.3277, 274.4662, 273.7328, 273.2353, 272.7945, 272.2167, 
    271.8291, 271.3987, 268.8894, 258.9529, 257.6884, 256.7748, 257.3061, 
    257.6007,
  275.993, 275.2983, 274.6071, 273.7831, 273.1396, 272.659, 272.0416, 
    271.6628, 271.4876, 268.8007, 259.3813, 258.451, 257.6712, 257.6299, 
    257.0624,
  275.2492, 274.2621, 273.9238, 273.3662, 272.6459, 272.1527, 271.8124, 
    271.2362, 269.3967, 262.8392, 261.3418, 259.9736, 258.3296, 258.3919, 
    258.1836,
  258.7344, 269.1049, 258.2493, 261.9556, 254.0632, 250.942, 254.3486, 
    254.0804, 255.3644, 248.1058, 247.487, 250.4166, 246.2, 245.6898, 239.1406,
  272.4656, 273.3843, 272.8066, 270.6246, 251.1052, 248.064, 254.774, 
    254.721, 254.4761, 254.3661, 248.7949, 254.9108, 256.253, 245.1077, 
    242.799,
  273.9827, 273.7234, 273.771, 273.2513, 262.1109, 244.6616, 252.6146, 
    254.808, 254.5642, 254.6463, 254.4886, 255.4542, 256.9922, 257.9901, 
    252.517,
  274.7054, 274.0907, 273.8301, 273.642, 273.1999, 264.5095, 245.567, 
    249.7584, 253.7267, 253.45, 253.6119, 254.6466, 256.465, 257.7623, 
    256.6761,
  275.041, 274.3675, 273.9087, 273.6406, 273.3306, 272.8951, 266.6671, 
    242.3952, 240.0457, 246.8207, 252.8125, 254.711, 256.5843, 258.0399, 
    259.662,
  275.4219, 274.6673, 274.0138, 273.5827, 273.3003, 272.9508, 272.045, 
    269.0595, 257.0401, 253.2696, 250.0012, 255.2472, 256.5043, 258.2053, 
    259.4999,
  276.0062, 275.0853, 274.2246, 273.5873, 273.2279, 272.7715, 272.3635, 
    271.5877, 268.7217, 264.4316, 258.795, 256.1262, 256.8917, 258.4243, 
    260.0999,
  276.3353, 275.3192, 274.4251, 273.7073, 273.2012, 272.7146, 272.1321, 
    271.7705, 271.2605, 268.3074, 257.8518, 256.8062, 257.2178, 258.4415, 
    259.7106,
  276.0136, 275.2884, 274.5872, 273.7401, 273.0653, 272.5688, 271.9345, 
    271.5723, 271.3958, 267.882, 257.9074, 257.4628, 256.9693, 258.4042, 
    259.3104,
  275.3009, 274.2386, 273.8794, 273.2974, 272.5501, 272.0278, 271.6898, 
    271.1641, 268.8966, 261.3301, 260.6493, 258.2077, 256.7633, 257.79, 
    259.0513,
  256.0547, 267.5735, 255.5841, 261.2415, 255.1591, 250.2682, 254.9458, 
    255.2014, 256.9654, 252.2241, 251.9227, 253.5082, 248.1113, 247.7612, 
    241.5481,
  272.0666, 273.2245, 272.7478, 269.8798, 249.7635, 247.5349, 254.8302, 
    255.5184, 256.0513, 257.2657, 254.3952, 258.3767, 258.4517, 243.4737, 
    242.8945,
  273.9179, 273.6344, 273.7255, 273.1617, 260.5818, 244.1057, 252.132, 
    255.6209, 256.7296, 257.4854, 258.4975, 259.9125, 260.458, 260.5782, 
    256.382,
  274.6455, 274.044, 273.788, 273.6263, 273.274, 264.1954, 244.4649, 
    251.0762, 255.7589, 256.9673, 258.6336, 260.0292, 260.9445, 261.266, 
    260.2172,
  274.9929, 274.3179, 273.8784, 273.6287, 273.3345, 272.9153, 267.0238, 
    244.3012, 247.6882, 253.8584, 258.83, 260.1953, 261.0816, 260.8702, 
    261.8288,
  275.3694, 274.6462, 273.9997, 273.5833, 273.2849, 272.9394, 272.0663, 
    268.8506, 256.9297, 255.2601, 257.3967, 260.3128, 260.6381, 260.7121, 
    261.4378,
  275.9828, 275.0732, 274.2289, 273.5674, 273.2015, 272.7139, 272.3181, 
    271.304, 268.0767, 264.0417, 260.4763, 261.2055, 261.7663, 260.6693, 
    261.1686,
  276.3317, 275.3253, 274.4116, 273.6974, 273.1785, 272.6189, 272.0475, 
    271.6994, 271.0421, 266.6947, 259.746, 261.0594, 261.7307, 261.064, 
    261.1573,
  276.0236, 275.2959, 274.6054, 273.7143, 272.9988, 272.4687, 271.8117, 
    271.4673, 271.1575, 265.9151, 258.6565, 260.4384, 261.1664, 261.7325, 
    261.6529,
  275.3553, 274.2736, 273.9008, 273.2834, 272.5017, 271.919, 271.5616, 
    271.0046, 268.8804, 262.5709, 258.5878, 260.2164, 260.6185, 261.581, 
    262.1179,
  254.9844, 266.7078, 256.2479, 261.7444, 256.8997, 251.0382, 256.961, 
    258.4613, 259.8134, 253.2231, 253.7732, 256.701, 253.6305, 253.5282, 
    249.7036,
  271.4563, 273.086, 272.8708, 270.2336, 254.3277, 249.2959, 256.7924, 
    258.0692, 258.6342, 258.9026, 255.5981, 259.9731, 260.6905, 250.9922, 
    251.5643,
  273.8395, 273.5293, 273.7067, 273.1008, 261.8173, 249.184, 253.0892, 
    258.1307, 258.9257, 258.9058, 258.5948, 259.636, 260.4421, 260.6278, 
    258.9453,
  274.5888, 274, 273.756, 273.6044, 273.2786, 264.463, 244.6446, 251.8942, 
    257.5504, 257.7927, 258.0379, 258.5286, 259.4493, 259.9791, 259.8974,
  274.9623, 274.2723, 273.8523, 273.6089, 273.307, 272.8636, 266.6365, 
    244.461, 249.6289, 251.0372, 256.6053, 257.6006, 258.4891, 258.8051, 
    259.7604,
  275.3355, 274.6484, 273.9874, 273.5603, 273.2319, 272.867, 271.8957, 
    267.7462, 256.429, 255.0652, 256.5939, 257.1265, 257.6491, 258.0772, 
    258.979,
  275.9623, 275.0689, 274.2415, 273.5623, 273.1661, 272.5992, 272.2316, 
    270.7809, 266.6182, 263.8119, 258.3108, 257.6032, 257.5847, 257.7484, 
    258.2825,
  276.334, 275.3205, 274.4169, 273.7029, 273.1769, 272.5452, 271.9664, 
    271.6275, 270.5271, 265.6189, 257.8878, 257.7196, 257.7774, 257.8984, 
    258.213,
  276.0262, 275.3021, 274.6427, 273.7456, 273.0204, 272.4655, 271.7491, 
    271.3806, 270.9822, 265.1923, 257.9356, 257.4417, 257.4038, 258.1793, 
    258.9951,
  275.3715, 274.2681, 273.8803, 273.2968, 272.5431, 271.9644, 271.5353, 
    271.0184, 269.1597, 261.439, 258.8222, 258.4683, 257.0549, 257.9058, 
    259.3874,
  255.3133, 265.6208, 259.5375, 262.4636, 257.5513, 252.0197, 259.1443, 
    257.6997, 257.4532, 252.3165, 252.3258, 255.4952, 254.5423, 254.8708, 
    250.6309,
  270.3796, 272.7484, 272.7814, 269.9684, 254.146, 250.6026, 256.8045, 
    259.3344, 256.7977, 256.3917, 254.5661, 257.0272, 258.3889, 252.7138, 
    251.3291,
  273.7852, 273.3992, 273.635, 272.9759, 264.7735, 252.148, 254.6519, 
    256.5119, 256.1799, 256.117, 255.9141, 257.2132, 258.5168, 259.0701, 
    257.8647,
  274.5171, 273.9458, 273.6912, 273.5402, 273.2387, 267.1989, 250.8799, 
    251.1846, 255.1062, 255.3668, 255.5533, 256.5909, 257.8994, 258.9374, 
    258.9826,
  274.8929, 274.2115, 273.7839, 273.5614, 273.2582, 272.7612, 268.1661, 
    245.0708, 245.2993, 252.5891, 256.1136, 256.2057, 256.7911, 257.7514, 
    259.3914,
  275.2686, 274.6214, 273.9446, 273.5193, 273.1681, 272.7621, 271.791, 
    267.5242, 256.7053, 253.2679, 254.829, 256.7251, 256.5588, 257.0464, 
    258.537,
  275.9199, 275.0461, 274.2226, 273.5508, 273.119, 272.5074, 272.2066, 
    270.8007, 267.2951, 262.9399, 258.9227, 258.3706, 257.3155, 256.4828, 
    257.8602,
  276.3246, 275.2837, 274.3971, 273.6827, 273.1523, 272.4875, 271.94, 
    271.6324, 270.5158, 266.3707, 261.1541, 259.8624, 258.463, 256.9846, 
    257.6781,
  276.0309, 275.3107, 274.6389, 273.6954, 272.9686, 272.441, 271.7638, 
    271.3987, 271.1348, 267.8981, 263.859, 261.4677, 259.5493, 257.9658, 
    259.2708,
  275.4294, 274.2887, 273.821, 273.2244, 272.485, 271.9181, 271.5509, 
    271.1154, 269.4875, 267.7783, 266.9395, 263.7391, 260.8296, 258.8926, 
    258.2512,
  257.8484, 262.9321, 258.2532, 258.6942, 257.5598, 256.1154, 258.4031, 
    257.8722, 254.9996, 251.904, 252.8035, 253.4739, 252.8228, 254.2226, 
    248.4757,
  269.8528, 272.3668, 272.1473, 268.2592, 255.3764, 254.4165, 258.5296, 
    259.3849, 255.8515, 253.9002, 252.8162, 256.7096, 258.0749, 251.2712, 
    250.8299,
  273.8242, 273.3284, 273.5565, 272.8175, 265.7813, 248.0203, 258.3732, 
    259.0348, 255.828, 254.8096, 255.7894, 258.8674, 259.8073, 259.1673, 
    257.6708,
  274.4552, 273.896, 273.6314, 273.4874, 273.1468, 267.6811, 253.9932, 
    254.3598, 256.5142, 255.2372, 255.9678, 259.959, 259.9866, 260.0898, 
    258.7133,
  274.8072, 274.1448, 273.7352, 273.5175, 273.2256, 272.6704, 269.0146, 
    256.439, 253.5935, 256.5647, 256.8487, 261.2872, 260.8449, 260.3583, 
    259.472,
  275.1932, 274.581, 273.908, 273.4819, 273.1196, 272.6393, 271.7257, 
    268.472, 263.8436, 260.5077, 259.1074, 262.6526, 262.6084, 261.3609, 
    260.7387,
  275.8719, 275.0561, 274.1823, 273.5023, 273.0554, 272.4315, 272.1454, 
    270.9206, 268.2538, 266.9952, 264.7383, 264.5096, 264.4232, 263.1309, 
    261.619,
  276.2607, 275.2393, 274.3685, 273.6564, 273.123, 272.4442, 271.8976, 
    271.6105, 270.5653, 267.9244, 266.7465, 266.1372, 265.6398, 264.384, 
    263.3113,
  275.9695, 275.2695, 274.6404, 273.6423, 272.8834, 272.3953, 271.7643, 
    271.3493, 271.018, 267.4733, 266.1728, 266.0613, 266.3351, 265.3022, 
    264.5887,
  275.3896, 274.2384, 273.7788, 273.1583, 272.4116, 271.8451, 271.522, 
    271.0857, 269.4509, 266.9691, 268.8282, 267.8737, 267.0375, 266.2297, 
    265.3116,
  259.8051, 262.1688, 259.4472, 258.6809, 255.6031, 253.335, 255.7259, 
    255.1952, 255.5512, 250.886, 250.8684, 254.0594, 254.0474, 256.6777, 
    249.4466,
  269.7392, 271.3168, 270.6687, 264.8833, 254.5056, 252.6844, 256.8243, 
    257.1283, 256.8672, 256.3022, 253.4411, 257.0636, 260.2488, 259.0181, 
    251.002,
  273.9132, 273.4326, 273.5182, 272.3384, 263.1278, 248.8943, 255.1485, 
    258.5269, 259.3969, 258.5767, 258.5746, 261.4783, 262.6459, 263.8695, 
    256.2332,
  274.4861, 273.9047, 273.5846, 273.4464, 272.9479, 265.5757, 249.5002, 
    254.8813, 260.7254, 262.5602, 261.5485, 263.8246, 264.4998, 264.5926, 
    259.1998,
  274.7736, 274.1234, 273.6849, 273.4635, 273.1832, 272.5741, 267.4618, 
    252.7394, 256.3778, 262.2302, 263.9773, 264.8841, 265.2112, 265.1161, 
    261.8595,
  275.1326, 274.5336, 273.8748, 273.4467, 273.0793, 272.5741, 271.5771, 
    267.6047, 263.2307, 264.8909, 264.3774, 265.602, 265.736, 265.448, 
    264.0216,
  275.8089, 275.075, 274.1571, 273.467, 273.012, 272.3793, 272.0926, 
    270.9685, 268.496, 267.795, 266.7874, 266.321, 266.1225, 265.4735, 264.829,
  276.2372, 275.2337, 274.3397, 273.6215, 273.0972, 272.3881, 271.8414, 
    271.5706, 270.3883, 265.8582, 264.7303, 265.7419, 266.5438, 266.4671, 
    265.0345,
  275.9367, 275.2625, 274.662, 273.5799, 272.7669, 272.3225, 271.7168, 
    271.231, 270.8013, 266.7975, 265.5283, 266.9633, 267.1128, 267.0129, 
    266.6698,
  275.348, 274.2106, 273.7214, 273.0666, 272.3137, 271.7346, 271.4595, 
    270.9091, 268.9311, 265.4422, 267.7896, 268.0709, 267.8289, 267.8049, 
    267.7654,
  257.7408, 260.0534, 257.1849, 257.1173, 254.1974, 251.1339, 253.6207, 
    254.5422, 256.2919, 257.2204, 256.066, 256.5437, 250.8286, 247.9422, 
    239.5541,
  269.9369, 269.9408, 269.2879, 261.4961, 253.0112, 249.7826, 254.943, 
    255.5426, 257.7307, 260.4174, 259.8125, 260.7949, 260.2144, 249.5608, 
    245.9465,
  273.9305, 273.3701, 273.456, 271.3721, 262.0311, 245.5097, 253.4762, 
    256.0917, 259.5244, 262.7686, 264.1909, 264.8886, 264.1262, 261.6875, 
    254.5158,
  274.5044, 273.8914, 273.5399, 273.4133, 272.6728, 264.6778, 247.4635, 
    253.2871, 259.1862, 264.3049, 264.6717, 265.3629, 265.506, 264.7501, 
    259.6867,
  274.7625, 274.0936, 273.6428, 273.4323, 273.1629, 272.4818, 267.0288, 
    247.6311, 253.4996, 261.8378, 264.8713, 265.419, 265.5477, 265.6792, 
    263.021,
  275.0899, 274.5039, 273.8474, 273.4293, 273.0679, 272.5971, 271.417, 
    266.8936, 259.108, 263.3022, 263.9113, 265.64, 265.5958, 263.4796, 
    265.2494,
  275.7655, 275.0854, 274.142, 273.4499, 273.005, 272.395, 272.0625, 
    270.6679, 267.8633, 265.43, 266.1409, 265.9814, 265.6881, 264.4514, 
    266.1855,
  276.2305, 275.2447, 274.3293, 273.618, 273.0891, 272.3822, 271.8036, 
    271.5392, 269.9291, 264.6161, 265.006, 265.9821, 266.2925, 266.4375, 
    266.8127,
  275.9325, 275.2645, 274.7031, 273.5467, 272.6991, 272.2752, 271.6626, 
    270.9646, 270.4804, 266.213, 262.5095, 262.3091, 265.9637, 265.8518, 
    266.869,
  275.3578, 274.2258, 273.6504, 272.9764, 272.2437, 271.6275, 271.3204, 
    270.675, 268.5437, 262.2607, 264.8125, 263.7725, 263.7009, 266.0242, 
    266.8346,
  255.4913, 258.4057, 254.9804, 256.2148, 252.7913, 249.6349, 256.9388, 
    258.9534, 261.0703, 260.2957, 260.2229, 261.9276, 260.5851, 259.0136, 
    250.4834,
  269.3956, 268.6115, 268.3885, 259.5112, 248.369, 246.7717, 254.6773, 
    258.3635, 260.6009, 262.2577, 261.1853, 263.2956, 263.89, 259.396, 
    251.0966,
  273.8749, 273.2404, 273.3706, 270.585, 260.53, 239.7695, 252.648, 255.6781, 
    259.4355, 261.8608, 262.7415, 263.7034, 264.638, 262.953, 256.0867,
  274.4667, 273.8389, 273.4886, 273.3974, 272.7339, 264.2141, 247.0208, 
    253.0855, 257.242, 261.2064, 262.3086, 263.5543, 264.6618, 263.6299, 
    258.0237,
  274.7085, 274.0462, 273.6031, 273.4174, 273.1544, 272.4672, 267.5945, 
    248.3837, 244.4841, 256.056, 261.5176, 262.288, 264.4021, 264.0652, 
    261.124,
  275.0496, 274.4895, 273.8286, 273.4103, 273.0544, 272.6043, 271.5776, 
    267.4005, 260.6358, 257.6543, 257.631, 261.8921, 263.8722, 264.2943, 
    262.3595,
  275.7498, 275.1176, 274.1256, 273.4279, 272.9846, 272.3968, 272.0557, 
    270.8692, 267.7672, 263.5724, 261.6072, 261.6573, 263.817, 264.5846, 
    263.5871,
  276.2297, 275.2646, 274.3403, 273.6097, 273.0684, 272.3772, 271.7845, 
    271.5191, 269.7391, 265.1537, 261.8109, 261.5683, 262.4059, 263.8673, 
    264.6624,
  275.9505, 275.2633, 274.7433, 273.4926, 272.6369, 272.2443, 271.6693, 
    270.8749, 270.4726, 266.8119, 262.8987, 261.5976, 260.7947, 260.8566, 
    265.2458,
  275.3916, 274.2032, 273.4849, 272.8431, 272.1842, 271.5215, 271.1727, 
    270.7617, 269.0523, 265.3802, 266.1292, 263.2765, 260.2289, 259.8576, 
    264.7091,
  256.3999, 260.2122, 257.7697, 257.7547, 254.0236, 250.4558, 255.4427, 
    256.0873, 256.7245, 249.7368, 250.5279, 250.6935, 242.5144, 239.2376, 
    232.677,
  269.8129, 269.1241, 268.978, 261.6635, 246.9639, 247.5541, 256.0057, 
    257.4374, 258.0507, 254.9801, 251.8942, 254.7084, 250.269, 235.7221, 
    231.2793,
  273.863, 273.1712, 273.3541, 270.9569, 260.4221, 245.3307, 255.5185, 
    258.5309, 259.3324, 258.0014, 256.3949, 255.8771, 251.7251, 248.3212, 
    240.5035,
  274.4283, 273.8021, 273.453, 273.3936, 272.9745, 266.2814, 252.6779, 
    258.4551, 260.2054, 259.0168, 256.7413, 256.7397, 252.9282, 249.3103, 
    245.5215,
  274.6831, 274.0278, 273.5776, 273.4177, 273.1613, 272.5593, 269.0302, 
    253.895, 256.4208, 257.1531, 257.2198, 256.2703, 254.5514, 251.0252, 
    250.2293,
  275.0233, 274.4883, 273.8141, 273.4017, 273.0447, 272.5921, 271.7986, 
    268.7964, 263.2321, 260.7208, 256.8461, 256.8776, 256.1172, 252.4184, 
    251.4064,
  275.7327, 275.1438, 274.1218, 273.4101, 272.9698, 272.3792, 272.0386, 
    271.1184, 268.4152, 264.9672, 261.5956, 258.2572, 259.0488, 254.5694, 
    252.586,
  276.2053, 275.2741, 274.3437, 273.5945, 273.0442, 272.3465, 271.7448, 
    271.487, 269.6131, 265.7553, 262.4025, 259.8885, 260.5084, 257.2082, 
    254.388,
  275.9474, 275.2489, 274.7729, 273.414, 272.5318, 272.1577, 271.5998, 
    270.6494, 270.5451, 266.502, 262.8755, 261.3647, 258.9998, 260.5729, 
    256.0471,
  275.4208, 274.1606, 273.2431, 272.6469, 272.0695, 271.2407, 270.5667, 
    270.1634, 268.4155, 264.597, 265.6621, 262.9386, 259.9089, 258.4049, 
    260.6532,
  259.765, 261.2604, 254.5857, 258.3969, 256.2451, 254.3397, 258.1888, 
    257.3545, 252.6005, 240.3658, 238.1652, 240.4409, 237.0461, 240.0196, 
    238.3978,
  270.1086, 269.5253, 268.7261, 262.0442, 253.6621, 253.9248, 260.1737, 
    260.6653, 255.9677, 249.692, 242.4517, 247.2364, 247.8545, 236.8153, 
    238.1164,
  273.7943, 273.0945, 273.3292, 270.9405, 261.7723, 252.53, 260.6912, 
    262.3778, 259.8159, 254.4771, 251.2998, 249.7056, 248.9686, 248.9385, 
    246.263,
  274.3969, 273.7846, 273.4286, 273.361, 273.0148, 268.0624, 258.457, 
    261.3614, 260.0614, 256.6569, 252.387, 250.6059, 249.6981, 249.6912, 
    249.0191,
  274.6638, 274.0318, 273.5482, 273.405, 273.1481, 272.5963, 269.6706, 
    259.8327, 257.6483, 255.683, 253.904, 251.7775, 250.2782, 250.4131, 
    251.584,
  275.0144, 274.4876, 273.8128, 273.3782, 273.0254, 272.5782, 271.8358, 
    268.4071, 260.7597, 258.2345, 255.0059, 253.4947, 251.2734, 250.733, 
    251.9906,
  275.7466, 275.1935, 274.1363, 273.3914, 272.947, 272.3426, 271.9915, 
    270.9395, 267.0555, 262.5739, 259.4057, 255.106, 252.8938, 251.694, 
    252.325,
  276.1856, 275.2856, 274.3539, 273.5707, 272.9977, 272.2794, 271.6616, 
    271.4023, 268.799, 265.0356, 260.3691, 257.2482, 255.2074, 253.1591, 
    252.9545,
  275.9142, 275.2336, 274.7815, 273.3258, 272.3955, 272.004, 271.4297, 
    270.0335, 270.3896, 267.3374, 264.0775, 261.3741, 258.7661, 256.4271, 
    252.8472,
  275.3447, 274.1028, 273.0961, 272.4668, 271.938, 270.9314, 269.786, 
    269.8009, 267.3459, 262.9824, 265.3964, 263.382, 261.3765, 258.2724, 
    255.0062,
  257.1618, 260.1322, 255.7452, 259.7032, 258.47, 258.9236, 261.5641, 
    260.6756, 256.7481, 254.0261, 251.5913, 250.4711, 244.506, 246.055, 
    243.8724,
  269.0121, 268.8453, 268.7527, 262.9405, 257.0565, 258.1103, 262.215, 
    260.795, 258.5734, 259.2452, 255.0893, 254.9616, 250.9405, 243.2707, 
    243.7855,
  273.6679, 272.9898, 273.2352, 271.3289, 264.1736, 256.7648, 261.9223, 
    261.385, 260.028, 259.3921, 259.4135, 256.497, 252.3278, 252.5511, 250.963,
  274.3492, 273.729, 273.377, 273.3178, 273.0088, 268.2652, 255.3313, 
    260.2639, 260.6092, 259.5465, 259.1792, 257.1452, 253.1092, 253.3548, 
    252.7137,
  274.6209, 273.9923, 273.4908, 273.374, 273.1312, 272.5627, 269.5948, 
    262.0695, 261.4711, 258.2891, 258.7147, 256.7664, 254.414, 253.7513, 
    254.9216,
  274.9905, 274.4518, 273.7841, 273.3468, 273.0012, 272.5346, 271.7939, 
    268.4343, 262.7001, 263.283, 260.3106, 258.8006, 255.4392, 254.0135, 
    255.3004,
  275.717, 275.2013, 274.141, 273.3602, 272.9126, 272.2973, 271.9579, 
    270.928, 268.1529, 265.0478, 263.4847, 259.8573, 256.8588, 253.8092, 
    255.0793,
  276.1672, 275.2779, 274.3417, 273.5353, 272.9347, 272.2413, 271.6227, 
    271.2839, 268.8209, 265.9385, 263.1435, 260.5706, 258.4793, 255.4518, 
    255.0401,
  275.8836, 275.2153, 274.772, 273.2664, 272.3131, 271.9322, 271.3247, 
    269.6071, 269.7917, 266.2745, 262.7999, 261.1917, 259.2701, 258.4158, 
    254.4539,
  275.2849, 274.1093, 273.1631, 272.4637, 271.9373, 270.5397, 269.1557, 
    269.4005, 268.3123, 262.6289, 263.759, 262.5549, 260.0944, 261.4789, 
    254.432,
  258.5455, 260.0048, 257.9618, 258.3116, 256.456, 256.6202, 258.1718, 
    258.7594, 258.8764, 257.8605, 257.0996, 256.5689, 254.7032, 250.6881, 
    245.2284,
  267.7038, 267.4616, 268.3911, 262.4344, 255.7056, 256.3724, 259.9209, 
    260.1223, 260.2967, 259.7435, 258.3181, 258.9698, 257.8702, 249.021, 
    243.3015,
  273.5511, 272.9118, 273.1674, 271.3489, 264.4506, 255.1225, 261.4525, 
    261.3624, 261.2821, 260.7027, 260.6651, 260.2331, 258.9054, 256.1511, 
    248.1142,
  274.2895, 273.6789, 273.3191, 273.2758, 272.9517, 267.7283, 255.4467, 
    260.7475, 261.863, 261.7559, 261.4262, 261.16, 260.1241, 257.2688, 
    250.0364,
  274.5691, 273.9396, 273.4363, 273.3292, 273.1275, 272.5593, 269.6757, 
    258.5706, 261.4299, 260.9512, 262.0744, 261.3398, 259.8461, 257.4077, 
    252.7568,
  274.9619, 274.4014, 273.7498, 273.3208, 272.9897, 272.5237, 271.8645, 
    268.9284, 264.2185, 262.4013, 261.7179, 262.1866, 260.5555, 258.1072, 
    254.1449,
  275.6987, 275.1789, 274.1142, 273.3354, 272.9136, 272.3357, 272.019, 
    271.1593, 269.0353, 265.9861, 264.47, 263.4713, 261.579, 258.0096, 254.659,
  276.202, 275.251, 274.3218, 273.5177, 272.9291, 272.3442, 271.6817, 
    271.2896, 269.445, 266.5284, 264.8203, 263.8855, 262.3618, 258.6783, 
    253.9778,
  275.9111, 275.2562, 274.7729, 273.3042, 272.3711, 272.0134, 271.4651, 
    269.7815, 269.3014, 266.9438, 265.3837, 264.8672, 262.7949, 258.6864, 
    253.2752,
  275.2826, 274.1603, 273.2781, 272.5515, 272.0021, 270.9426, 269.1411, 
    268.913, 268.5025, 266.7578, 267.8131, 266.135, 263.4007, 259.2018, 
    253.2122,
  257.2408, 259.2545, 257.7996, 257.7455, 255.5109, 255.7518, 256.7701, 
    255.9015, 255.4782, 254.3918, 254.8634, 254.8193, 254.7322, 255.4051, 
    251.251,
  266.0839, 266.3321, 267.7519, 261.9953, 254.1998, 255.8492, 258.5388, 
    257.4074, 257.1887, 256.7464, 258.168, 259.5324, 259.1149, 256.3187, 
    250.3964,
  273.5185, 272.8719, 273.1445, 271.5328, 263.2332, 258.2949, 261.029, 
    260.1366, 260.0413, 260.6573, 261.8568, 262.5756, 261.75, 260.5084, 
    252.3062,
  274.2519, 273.6601, 273.3004, 273.2778, 272.9305, 267.4917, 256.3882, 
    261.8626, 263.8237, 264.4254, 265.7059, 265.1502, 264.2549, 262.3358, 
    252.3319,
  274.5382, 273.9296, 273.4319, 273.3287, 273.1759, 272.6329, 270.1475, 
    262.4747, 263.2605, 266.809, 267.9079, 265.5099, 264.9532, 262.7173, 
    252.6517,
  274.9944, 274.3956, 273.7484, 273.3305, 273.0586, 272.638, 272.133, 
    270.4645, 268.2478, 268.3206, 266.8927, 264.536, 264.8539, 262.8098, 
    251.8761,
  275.6975, 275.1724, 274.0934, 273.3505, 272.9596, 272.4801, 272.1797, 
    271.6091, 270.6943, 268.6085, 264.7259, 264.1185, 265.0194, 261.2762, 
    251.1647,
  276.2596, 275.2292, 274.3107, 273.5246, 272.9436, 272.4702, 271.7656, 
    271.4477, 269.9432, 266.0569, 262.5257, 265.0721, 265.3208, 259.3888, 
    249.682,
  275.9636, 275.2982, 274.7947, 273.3591, 272.434, 272.0595, 271.5509, 
    270.6318, 269.4323, 266.4699, 262.5348, 265.6458, 264.1146, 256.2823, 
    246.7563,
  275.2642, 274.2906, 273.4614, 272.6441, 272.0522, 271.161, 270.0121, 
    269.2784, 268.0649, 263.283, 266.812, 266.8287, 262.2794, 253.8378, 
    247.8748,
  255.2176, 257.2505, 255.0183, 254.3205, 251.4027, 252.1358, 253.9391, 
    252.3714, 251.745, 249.4204, 250.1017, 251.9785, 252.122, 255.0968, 
    257.0967,
  263.9683, 264.6019, 264.802, 259.4423, 250.2698, 254.5575, 256.5143, 
    253.899, 253.3924, 252.5178, 252.047, 255.0724, 256.6092, 257.9641, 
    257.9482,
  273.5501, 272.668, 273.0653, 271.2196, 259.7646, 250.7071, 259.0922, 
    256.4021, 255.0151, 254.6192, 255.327, 257.0214, 259.5905, 261.2477, 
    255.9668,
  274.2795, 273.7451, 273.381, 273.3422, 272.7873, 265.0733, 252.9165, 
    257.9372, 258.2026, 257.0858, 257.6763, 259.6982, 261.215, 262.2988, 
    253.8214,
  274.5779, 273.9961, 273.558, 273.3848, 273.213, 272.6584, 268.9424, 
    254.5214, 254.8228, 259.2424, 260.9365, 261.5836, 262.4968, 262.0359, 
    254.4305,
  275.1104, 274.4443, 273.7893, 273.3686, 273.1443, 272.7885, 272.3354, 
    269.2272, 261.0244, 259.6162, 260.6879, 262.4651, 263.5399, 260.584, 
    251.8785,
  275.7755, 275.2254, 274.1018, 273.3737, 273.0326, 272.6858, 272.3557, 
    271.7706, 269.5887, 263.5669, 262.39, 263.1355, 262.8331, 257.916, 251.451,
  276.3286, 275.2251, 274.3158, 273.5371, 272.9827, 272.6343, 271.9421, 
    271.6789, 270.1666, 265.8268, 263.8296, 263.6819, 262.7558, 255.6921, 
    249.2518,
  276.0054, 275.3188, 274.8228, 273.4669, 272.5674, 272.1721, 271.7829, 
    271.1333, 270.2589, 267.7849, 265.0698, 264.5752, 261.6354, 253.4746, 
    246.7913,
  275.2088, 274.307, 273.5334, 272.7013, 272.1494, 271.5162, 271.0345, 
    270.7685, 270.2915, 268.5139, 267.4306, 265.2571, 260.4205, 252.065, 
    248.028,
  257.5839, 259.4006, 255.1185, 254.4659, 250.3105, 250.8833, 253.7178, 
    250.7767, 249.3303, 243.7212, 244.0152, 246.4687, 243.1907, 244.7571, 
    240.8385,
  263.3293, 264.3548, 262.5408, 257.2349, 249.1114, 254.1671, 255.6238, 
    251.8483, 250.8727, 248.5475, 246.6271, 249.869, 249.5187, 244.2839, 
    238.0291,
  273.4686, 271.8941, 272.2135, 269.3552, 256.0433, 248.266, 258.1459, 
    254.0362, 252.0791, 250.3408, 250.5912, 250.1963, 250.3256, 250.8261, 
    245.7233,
  274.2995, 273.7518, 273.3999, 273.3279, 271.6852, 262.1872, 249.7182, 
    256.0474, 255.2117, 252.8592, 251.8204, 251.4317, 251.669, 253.0149, 
    250.4192,
  274.559, 273.9901, 273.5477, 273.3637, 273.1767, 272.4173, 267.4933, 
    250.194, 251.0845, 255.3389, 255.8887, 254.2383, 252.949, 254.6861, 
    253.2577,
  275.1367, 274.416, 273.7405, 273.3247, 273.1206, 272.7885, 272.3514, 
    268.842, 259.1638, 256.53, 256.3115, 256.4973, 254.9452, 255.1307, 
    253.0535,
  275.8188, 275.2771, 274.0569, 273.3147, 273.0007, 272.734, 272.4352, 
    271.9037, 270.0084, 262.5981, 259.3196, 257.3875, 256.1146, 255.7249, 
    252.7049,
  276.3302, 275.2278, 274.2772, 273.455, 272.9102, 272.6602, 272.0147, 
    271.8365, 270.3573, 264.2873, 261.5746, 259.5772, 257.1716, 255.4298, 
    251.9996,
  276.0013, 275.3087, 274.8162, 273.3798, 272.4781, 272.1068, 271.7961, 
    271.3369, 269.9147, 266.7169, 263.4074, 261.3708, 257.6349, 255.9137, 
    250.0415,
  275.1629, 274.271, 273.4054, 272.3837, 272.0106, 271.1245, 269.3828, 
    269.4795, 269.6342, 268.5923, 266.7255, 263.2189, 259.2096, 256.0294, 
    251.2969,
  257.9846, 260.2383, 257.4946, 256.8639, 252.9679, 253.5941, 256.3068, 
    251.6525, 250.5468, 244.3374, 243.1411, 243.8471, 238.097, 238.2909, 
    233.1817,
  263.0524, 264.2772, 262.2477, 257.7983, 251.4593, 256.1444, 256.3396, 
    252.2338, 251.3289, 249.2435, 246.2572, 248.9768, 247.508, 235.9785, 
    231.9022,
  273.139, 270.9613, 270.6339, 265.8912, 257.5349, 250.4442, 256.7338, 
    253.1002, 251.952, 250.6457, 251.6358, 249.5214, 247.4429, 246.0038, 
    238.8611,
  274.2741, 273.7215, 273.3588, 273.1169, 270.0858, 262.3517, 250.0483, 
    253.5003, 253.089, 251.4441, 251.06, 250.2439, 248.7409, 247.9058, 
    244.3198,
  274.5521, 273.9572, 273.5092, 273.3179, 273.0782, 271.7834, 267.068, 
    248.8077, 248.2294, 251.9908, 253.1551, 252.5349, 250.4329, 250.8084, 
    249.7747,
  275.1724, 274.3629, 273.6976, 273.2752, 273.0797, 272.7534, 272.2237, 
    267.9279, 258.7344, 255.0169, 254.9373, 254.7903, 251.9631, 251.3439, 
    249.3944,
  275.822, 275.3112, 274.0594, 273.2678, 272.9647, 272.7124, 272.4189, 
    271.8678, 269.5392, 261.1646, 257.4056, 255.2584, 253.2736, 252.0195, 
    250.1723,
  276.2973, 275.2265, 274.2392, 273.4134, 272.8535, 272.637, 272.001, 
    271.8039, 269.8463, 261.7938, 257.2992, 255.5166, 254.2171, 251.9277, 
    249.5964,
  276.0026, 275.3013, 274.8289, 273.3494, 272.445, 272.0746, 271.7484, 
    271.3371, 268.8109, 261.9336, 258.0487, 256.8496, 254.838, 252.235, 
    248.7702,
  275.1239, 274.254, 273.3891, 272.4114, 271.9694, 271.0024, 268.9856, 
    268.2802, 266.3049, 261.657, 262.5665, 259.1699, 256.281, 253.3983, 
    250.6303,
  257.3974, 259.3055, 257.3921, 256.4687, 252.0229, 251.6227, 254.4621, 
    249.3326, 249.6694, 242.1081, 239.8974, 242.3671, 238.8073, 239.1202, 
    235.7393,
  263.3317, 264.0448, 263.2162, 256.9912, 250.936, 253.2241, 252.6225, 
    250.0126, 249.5572, 248.5078, 243.8342, 247.9144, 247.6811, 235.7902, 
    232.946,
  271.9964, 269.7082, 269.2904, 262.5642, 257.5266, 247.2527, 251.8458, 
    250.6836, 250.5468, 249.8687, 250.7668, 247.9116, 246.6388, 245.8637, 
    238.5804,
  274.246, 273.6585, 273.2713, 272.1198, 268.8778, 260.9869, 246.0151, 
    250.3982, 250.8472, 249.7423, 249.1476, 247.7763, 246.9193, 246.4116, 
    244.3435,
  274.5376, 273.9007, 273.4701, 273.2679, 272.7692, 270.64, 266.1456, 
    246.3027, 242.8291, 246.5489, 250.3294, 249.9253, 248.3321, 248.7202, 
    249.1043,
  275.1648, 274.2884, 273.6589, 273.2292, 273.0457, 272.7052, 271.7821, 
    266.9371, 258.361, 254.0828, 251.0541, 252.6142, 249.7502, 248.9411, 
    247.9025,
  275.797, 275.2505, 274.0341, 273.2294, 272.9352, 272.6911, 272.3976, 
    271.6802, 268.8371, 261.4758, 256.8692, 253.6195, 251.0448, 249.7973, 
    248.1467,
  276.3008, 275.2379, 274.21, 273.404, 272.832, 272.6361, 272.0127, 271.7712, 
    269.3201, 260.7247, 255.89, 253.2117, 252.0289, 249.7044, 247.701,
  276.0572, 275.3099, 274.8426, 273.3829, 272.4914, 272.0625, 271.75, 
    271.4413, 268.8755, 259.7021, 255.8278, 254.2458, 252.8054, 250.1986, 
    247.3439,
  275.1562, 274.2844, 273.4535, 272.5233, 272.043, 271.2617, 269.6443, 
    268.6699, 263.6026, 257.913, 259.5656, 256.199, 253.541, 251.5326, 
    249.6402,
  257.4521, 258.2274, 255.5104, 254.7123, 250.2363, 248.9707, 251.9292, 
    248.8988, 251.291, 244.469, 242.8387, 245.1734, 241.8293, 240.945, 
    237.0543,
  264.8885, 262.763, 262.1396, 254.8195, 249.2115, 248.2616, 250.1127, 
    249.3316, 249.5894, 251.0685, 245.8151, 249.1857, 250.0144, 239.0983, 
    236.0677,
  271.2649, 267.9334, 267.567, 259.0616, 256.8001, 243.297, 249.1681, 
    250.2745, 250.4766, 250.1766, 250.7491, 249.2624, 249.3917, 248.9642, 
    242.5973,
  274.1644, 273.4067, 272.972, 269.957, 267.7047, 259.6415, 243.9872, 
    249.0561, 250.2373, 249.3274, 249.0091, 248.7189, 249.0112, 249.4817, 
    248.1353,
  274.5092, 273.8067, 273.3994, 273.1853, 272.2384, 269.596, 265.9099, 
    243.4655, 239.4586, 245.3037, 249.818, 250.3722, 249.7821, 250.4848, 
    251.9268,
  275.0787, 274.214, 273.6041, 273.1562, 272.9766, 272.5529, 271.0225, 
    265.8235, 257.0087, 253.0668, 249.454, 252.0919, 250.5391, 250.4632, 
    251.2423,
  275.713, 275.0955, 273.9364, 273.1538, 272.8747, 272.6291, 272.3139, 
    271.134, 267.6054, 260.1685, 255.0851, 252.7498, 251.4361, 250.8238, 
    250.4841,
  276.2202, 275.1645, 274.1198, 273.3406, 272.765, 272.5799, 271.9516, 
    271.6836, 267.1855, 258.6861, 254.3005, 252.9212, 252.3999, 250.5809, 
    250.7149,
  276.0113, 275.2356, 274.7756, 273.3801, 272.4804, 271.9947, 271.692, 
    271.0983, 267.2644, 256.8272, 254.8345, 254.4334, 253.9112, 251.8138, 
    250.9388,
  275.1264, 274.2669, 273.5304, 272.5751, 272.0034, 271.0981, 269.2435, 
    267.8434, 259.5915, 253.5431, 257.7595, 255.6172, 254.4427, 253.6789, 
    252.1361,
  256.2746, 257.5533, 254.0743, 254.9568, 250.8271, 249.1298, 251.8147, 
    250.1349, 252.3763, 244.7259, 241.9314, 244.5828, 242.2917, 242.1575, 
    238.6417,
  265.054, 262.0869, 261.3595, 255.3523, 248.651, 247.1106, 250.8935, 
    250.9965, 251.1021, 253.0903, 247.8186, 251.8668, 253.4694, 243.2242, 
    241.2866,
  271.3152, 266.9032, 267.0373, 259.5907, 257.9151, 241.4212, 249.6796, 
    251.8373, 252.9228, 253.3464, 253.8209, 253.7143, 254.4439, 254.2383, 
    248.552,
  274.0993, 273.1487, 272.6738, 269.1543, 268.3638, 260.375, 240.7971, 
    250.9343, 253.2367, 253.4199, 253.562, 254.1458, 254.7355, 255.0873, 
    253.5862,
  274.4668, 273.7447, 273.3539, 273.1531, 272.321, 269.9882, 266.3231, 
    243.634, 245.4554, 252.5764, 254.3455, 255.4681, 255.229, 255.9684, 
    256.5717,
  274.9944, 274.1907, 273.5665, 273.1268, 272.9574, 272.4264, 270.6579, 
    265.8049, 258.7833, 257.02, 253.8152, 255.7851, 256.42, 256.5999, 257.9458,
  275.6849, 275.0205, 273.8943, 273.1256, 272.8561, 272.6041, 272.2311, 
    270.769, 266.8594, 260.3363, 256.8398, 256.088, 256.3405, 256.7915, 
    257.7694,
  276.1913, 275.1321, 274.0812, 273.3196, 272.7349, 272.5338, 271.8901, 
    271.5464, 265.468, 259.079, 256.8101, 255.6787, 255.7464, 255.9022, 
    257.4897,
  275.9829, 275.2013, 274.7446, 273.3934, 272.4686, 271.9475, 271.6088, 
    270.394, 266.1137, 258.4798, 257.7256, 256.8001, 255.1494, 255.1968, 
    256.5917,
  275.1001, 274.2632, 273.6003, 272.5879, 271.9432, 270.8187, 268.7047, 
    267.6531, 259.6153, 255.7826, 259.0283, 256.8707, 254.954, 254.2061, 
    255.8466,
  254.1161, 257.9501, 253.0348, 254.8094, 250.5652, 247.839, 250.2364, 
    249.129, 250.9357, 242.0159, 240.1481, 243.6634, 242.5377, 244.2217, 
    241.0517,
  265.1042, 262.2183, 260.5763, 255.6806, 248.6924, 246.5492, 251.4139, 
    251.1435, 250.7698, 251.0127, 245.2794, 249.9681, 251.3574, 241.6057, 
    239.0264,
  271.7818, 267.5018, 267.8704, 260.4503, 258.1057, 240.187, 251.2689, 
    254.0592, 253.8924, 253.5131, 252.8562, 251.8599, 251.6858, 251.1175, 
    245.2935,
  274.0724, 273.2577, 272.7676, 269.7541, 268.8676, 262.2003, 245.613, 
    252.815, 255.0368, 254.1364, 252.8099, 252.19, 251.8052, 252.5608, 
    250.1825,
  274.4107, 273.7129, 273.3458, 273.1797, 272.7254, 270.4934, 267.4274, 
    249.3441, 249.0307, 251.8792, 253.8612, 253.1291, 253.183, 255.3174, 
    253.3496,
  274.9336, 274.1894, 273.5632, 273.1249, 272.9749, 272.4213, 270.5567, 
    266.1417, 260.6613, 257.541, 254.3233, 256.1063, 256.3432, 255.3706, 
    253.6412,
  275.6716, 275.0376, 273.888, 273.1171, 272.8534, 272.5955, 272.1342, 
    270.6456, 266.2964, 262.1576, 260.3064, 258.0371, 257.35, 255.5912, 
    254.1984,
  276.1874, 275.1228, 274.0721, 273.3124, 272.6979, 272.5018, 271.8423, 
    271.1288, 264.438, 261.2134, 260.152, 259.9408, 259.1609, 259.412, 260.107,
  275.9585, 275.1785, 274.7184, 273.3971, 272.4479, 271.9045, 271.4261, 
    269.5452, 265.0253, 260.9955, 260.4804, 260.2276, 259.2066, 257.6466, 
    256.9321,
  275.0826, 274.2427, 273.6453, 272.5838, 271.9053, 270.2486, 268.4061, 
    267.0065, 262.0448, 259.5826, 260.3714, 257.7854, 257.1207, 256.1399, 
    257.0607,
  253.1099, 256.1921, 252.171, 254.0396, 250.2621, 249.2637, 252.8562, 
    253.4417, 255.8459, 252.224, 251.0199, 251.1218, 247.0618, 247.0502, 
    242.6216,
  263.3271, 260.6336, 258.9454, 255.0649, 248.5797, 247.366, 252.4522, 
    253.5781, 254.0506, 256.0924, 252.3246, 254.2985, 254.4421, 245.9573, 
    242.1832,
  271.4276, 266.4766, 266.817, 259.2923, 256.5161, 241.8642, 251.0937, 
    253.6473, 254.463, 255.0117, 255.2888, 254.2202, 254.3996, 252.785, 
    247.402,
  274.0431, 273.1837, 272.5995, 268.3494, 267.3824, 259.7665, 243.5015, 
    250.6545, 253.5056, 253.7616, 253.6221, 253.3419, 253.5508, 252.6574, 
    250.6391,
  274.3841, 273.6919, 273.3, 273.1218, 272.6639, 269.6481, 266.2161, 245.497, 
    243.5335, 250.6455, 254.1523, 254.4897, 254.506, 254.2551, 253.1869,
  274.9441, 274.2058, 273.5624, 273.0866, 272.9543, 272.2946, 269.9509, 
    264.8732, 259.0874, 257.1989, 253.9452, 256.0368, 255.8408, 254.6507, 
    254.0274,
  275.7346, 275.1613, 273.924, 273.109, 272.8218, 272.5489, 271.9723, 
    269.9324, 265.1796, 260.0078, 258.4264, 256.6062, 255.9302, 253.8126, 
    253.6113,
  276.249, 275.171, 274.099, 273.2876, 272.651, 272.4335, 271.7762, 270.9297, 
    263.5533, 259.6612, 258.3961, 257.4798, 257.0883, 255.6969, 254.6959,
  275.9928, 275.2042, 274.7374, 273.3633, 272.4213, 271.8487, 271.3405, 
    269.4715, 263.724, 260.2927, 259.5827, 259.312, 257.7398, 254.7487, 
    253.6403,
  275.0726, 274.2224, 273.6266, 272.4986, 271.8418, 270.0565, 268.9704, 
    267.7858, 262.6658, 260.8493, 261.3207, 259.0689, 255.3562, 253.4216, 
    254.1455,
  251.4681, 255.7788, 250.8235, 254.8812, 249.7813, 250.9408, 256.4041, 
    255.3145, 255.069, 248.6559, 248.187, 248.157, 244.3119, 242.4046, 
    238.4978,
  260.8959, 260.1083, 259.3758, 255.5512, 247.1116, 249.34, 256.1734, 
    256.0118, 255.1262, 254.5261, 247.6773, 250.6775, 250.2852, 241.0845, 
    240.1223,
  270.4635, 266.5772, 267.1268, 260.5518, 258.6562, 248.7139, 255.0821, 
    256.8192, 256.1246, 254.4206, 253.0108, 251.3809, 250.8321, 250.3852, 
    245.5341,
  273.9788, 273.1358, 272.6374, 268.8552, 267.6557, 261.8646, 249.5057, 
    253.8112, 253.0882, 252.6526, 251.3931, 250.2177, 249.8697, 249.6259, 
    249.7967,
  274.3799, 273.6537, 273.2578, 273.0742, 272.5873, 269.4557, 266.6178, 
    247.6555, 245.8061, 249.2591, 251.0592, 250.2711, 250.1853, 250.8262, 
    251.2147,
  274.9768, 274.1867, 273.5465, 273.0521, 272.9328, 272.1469, 269.5549, 
    264.6026, 259.8364, 257.2274, 251.7672, 251.4923, 250.9796, 251.0322, 
    251.4568,
  275.7752, 275.2395, 273.9755, 273.0966, 272.7901, 272.4908, 271.8429, 
    268.9964, 263.7325, 257.7569, 254.8433, 252.6791, 251.7225, 250.9346, 
    251.3348,
  276.2927, 275.2279, 274.1313, 273.246, 272.5981, 272.3619, 271.7059, 
    270.7208, 262.2509, 257.2063, 254.6604, 253.3227, 252.1593, 251.1425, 
    251.4176,
  276.0703, 275.24, 274.7689, 273.3117, 272.3831, 271.7628, 271.2152, 
    268.7807, 261.1973, 256.8266, 255.0476, 254.0198, 252.1987, 251.2677, 
    251.8877,
  275.1141, 274.2129, 273.5556, 272.3948, 271.7679, 270.033, 269.0065, 
    266.9785, 259.6298, 258.101, 257.166, 254.5811, 252.6616, 252.0983, 
    252.671,
  248.9198, 255.3319, 251.2292, 255.9121, 253.6618, 253.3477, 254.9478, 
    253.1472, 254.1902, 248.2948, 245.7835, 246.2175, 243.3771, 241.5579, 
    237.0471,
  259.5123, 259.3848, 258.7333, 256.0197, 249.0624, 250.4051, 254.1403, 
    253.078, 252.772, 253.1079, 248.7374, 250.1749, 250.8346, 240.4587, 
    238.0164,
  269.5685, 267.1025, 267.2154, 261.3081, 256.1218, 244.5208, 251.4761, 
    252.6851, 253.1365, 253.5631, 253, 250.5443, 250.566, 250.8917, 244.8284,
  273.8984, 273.1169, 272.7786, 269.5369, 267.7686, 260.3098, 243.9233, 
    249.3667, 252.0858, 252.356, 251.1642, 248.6685, 248.8862, 248.7862, 
    249.4867,
  274.3961, 273.5835, 273.192, 273.0051, 272.6305, 269.5181, 266.1531, 
    243.3089, 241.7229, 247.7632, 249.813, 248.5959, 248.8314, 249.764, 
    250.909,
  275.0541, 274.1627, 273.5388, 273.0184, 272.9129, 272.1521, 269.5251, 
    263.7668, 257.4698, 255.6619, 250.0385, 249.3747, 249.2716, 249.7533, 
    250.5287,
  275.8438, 275.2972, 274.0477, 273.077, 272.7588, 272.4412, 271.8243, 
    267.9873, 261.6664, 255.2629, 252.6296, 250.5163, 249.9587, 249.7338, 
    250.4733,
  276.3104, 275.3196, 274.1892, 273.2077, 272.5406, 272.3162, 271.6502, 
    270.795, 261.209, 254.0663, 251.8837, 250.9335, 250.3645, 249.6588, 
    250.1877,
  276.1419, 275.2851, 274.7917, 273.2291, 272.3141, 271.6714, 271.1694, 
    268.8577, 259.1045, 253.0279, 251.3775, 251.2904, 250.5268, 249.8486, 
    250.7094,
  275.152, 274.1856, 273.3727, 272.2148, 271.5926, 270.041, 269.1037, 
    266.9337, 258.2263, 253.8731, 254.4631, 252.2057, 251.2635, 251.1693, 
    251.5549,
  250.9916, 254.9588, 251.2384, 256.8748, 253.5828, 251.6057, 252.3947, 
    249.8441, 249.0851, 240.8763, 239.7119, 244.9798, 244.341, 239.6141, 
    233.8912,
  258.253, 258.3376, 258.4221, 257.1427, 249.6232, 247.341, 251.1536, 
    250.7276, 248.7654, 248.5828, 243.0863, 249.2433, 252.0812, 237.962, 
    234.0253,
  268.7014, 266.9093, 266.3731, 261.1729, 257.4292, 243.1647, 248.0502, 
    250.2701, 249.6869, 249.5782, 249.2242, 250.0524, 251.8389, 250.3592, 
    243.3525,
  273.8438, 273.0887, 272.8058, 269.9133, 267.6759, 261.1727, 242.5165, 
    248.2352, 251.0977, 249.7037, 248.0465, 247.7475, 249.1666, 250.4836, 
    248.0103,
  274.3906, 273.5419, 273.1373, 272.9281, 272.6264, 269.9988, 265.5868, 
    243.4818, 241.9013, 248.7223, 248.0305, 247.5223, 248.4883, 249.8371, 
    249.9851,
  275.0467, 274.127, 273.5189, 272.981, 272.8809, 272.1895, 269.6862, 
    263.2824, 257.5309, 256.4718, 251.145, 248.8263, 248.4202, 248.6481, 
    248.9314,
  275.8218, 275.232, 274.0206, 273.0493, 272.7299, 272.3868, 271.8955, 
    267.9938, 263.0237, 257.4594, 253.6852, 249.7434, 248.9394, 248.4084, 
    248.7997,
  276.2523, 275.2907, 274.1722, 273.1698, 272.4984, 272.2493, 271.5903, 
    271.002, 263.7486, 256.3093, 252.82, 250.3744, 249.1239, 248.1884, 248.328,
  276.1106, 275.265, 274.744, 273.1786, 272.2488, 271.5043, 271.1202, 
    269.2352, 260.7984, 254.7581, 252.7836, 251.3666, 249.6111, 248.3539, 
    248.6759,
  275.1497, 274.1418, 273.2144, 272.0735, 271.3949, 269.5202, 268.821, 
    267.3398, 259.9612, 256.3078, 256.308, 252.3901, 250.4729, 249.9325, 
    249.4377,
  256.2216, 255.8438, 253.5358, 254.5523, 252.7565, 249.1104, 248.1023, 
    247.9798, 247.9537, 239.2133, 238.2341, 242.1687, 239.3678, 237.4415, 
    231.7962,
  259.3495, 258.6533, 257.4804, 256.1133, 251.515, 246.8957, 247.9223, 
    247.7342, 246.838, 246.755, 242.0114, 248.6534, 249.663, 235.6185, 232.252,
  267.0787, 266.2352, 263.4526, 259.435, 255.3161, 242.5214, 246.9189, 
    247.5124, 247.108, 248.2099, 248.9582, 250.0945, 251.0307, 248.8377, 
    242.1992,
  273.8237, 272.7597, 272.2201, 268.1805, 264.5037, 256.4087, 241.7403, 
    245.5747, 246.8666, 247.1748, 247.2468, 248.5026, 251.2439, 249.7354, 
    246.6447,
  274.3411, 273.5347, 273.1399, 272.9276, 272.4421, 268.2218, 263.3477, 
    242.3742, 239.8401, 245.0989, 247.0635, 248.0223, 250.5528, 251.7527, 
    249.1626,
  274.9766, 274.0958, 273.492, 272.9774, 272.8546, 272.0922, 269.0747, 
    262.6012, 256.4459, 255.3415, 251.1415, 248.9799, 248.9644, 249.9489, 
    248.7636,
  275.7298, 275.0738, 273.9169, 273.0197, 272.728, 272.371, 271.9065, 
    267.516, 263.7223, 258.4695, 253.9239, 249.6044, 249.0255, 249.2159, 
    248.6393,
  276.1982, 275.1733, 274.084, 273.1797, 272.5744, 272.2977, 271.5504, 
    270.9574, 265.6963, 260.7762, 254.7693, 250.578, 249.0831, 248.088, 
    247.7999,
  276.0409, 275.2072, 274.6552, 273.3866, 272.3855, 271.4953, 270.8924, 
    268.8925, 262.5913, 261.1925, 259.0763, 254.776, 250.3772, 247.9753, 
    247.1773,
  275.12, 274.1942, 273.5717, 272.4172, 271.5469, 269.3432, 268.1049, 
    266.0171, 261.1167, 260.644, 262.4797, 259.1064, 255.1835, 251.3601, 
    248.3136,
  264.2712, 262.4092, 258.0812, 253.6475, 249.5433, 246.9764, 247.9901, 
    248.125, 248.66, 239.6874, 238.0395, 240.2962, 237.0039, 236.7011, 
    230.6905,
  265.7346, 264.0482, 260.6443, 254.4781, 248.5598, 245.5392, 246.9679, 
    247.5795, 247.5703, 246.7787, 241.8177, 246.7174, 246.5787, 234.5442, 
    231.2742,
  270.0378, 268.4935, 263.5876, 257.2388, 253.2885, 242.2089, 245.8106, 
    247.2767, 247.515, 248.4281, 248.4841, 248.4159, 248.3168, 246.7545, 
    241.2826,
  273.8704, 273.061, 271.52, 265.7963, 260.7081, 255.4077, 241.7094, 
    244.6169, 246.5392, 247.7237, 247.5567, 248.0138, 248.2952, 247.4673, 
    245.0144,
  274.325, 273.5225, 273.128, 272.7355, 270.9522, 265.9546, 262.3366, 
    242.0899, 239.7778, 244.5512, 247.4326, 248.5104, 248.5712, 248.6752, 
    247.6759,
  274.9778, 274.0892, 273.4594, 272.9564, 272.8117, 271.8737, 267.7545, 
    261.1922, 255.3836, 254.8468, 250.798, 249.7592, 248.8509, 248.7054, 
    247.486,
  275.764, 275.0428, 273.8655, 272.9903, 272.7156, 272.3963, 271.7026, 
    265.2187, 260.4065, 256.8994, 253.6048, 249.8972, 249.3965, 248.6379, 
    247.8431,
  276.2041, 275.1299, 274.0563, 273.1906, 272.6376, 272.4221, 271.6294, 
    270.4015, 262.9222, 255.6949, 252.5627, 250.2223, 249.5748, 248.1504, 
    247.6404,
  276.0355, 275.1832, 274.6097, 273.5705, 272.618, 271.6865, 271.0397, 
    268.9676, 259.5729, 255.0842, 253.29, 251.299, 249.767, 247.9862, 246.6318,
  275.1302, 274.1876, 273.7263, 272.8222, 271.9072, 269.9682, 267.9725, 
    264.0702, 257.8773, 255.9524, 258.1293, 254.9928, 252.1638, 249.5937, 
    247.5457,
  264.8376, 266.6855, 266.2374, 261.1334, 254.4167, 249.4921, 250.007, 
    248.7418, 247.2183, 238.2913, 237.6193, 239.0633, 235.6888, 235.6104, 
    231.1857,
  266.8638, 268.3983, 267.4174, 260.4619, 250.9598, 247.8916, 248.0402, 
    247.519, 246.1313, 244.8852, 240.7733, 244.7794, 244.346, 233.2941, 
    230.4253,
  271.0384, 269.8776, 268.2294, 261.2747, 254.8114, 243.3681, 246.1768, 
    247.1348, 246.7383, 246.3795, 245.9865, 245.6228, 245.4221, 244.1422, 
    239.0371,
  273.8917, 273.3023, 272.2925, 266.5638, 261.6694, 256.4609, 241.696, 
    244.52, 245.8308, 246.1315, 245.0354, 245.042, 244.8213, 244.5234, 
    243.1342,
  274.341, 273.5213, 273.1414, 272.4619, 268.6402, 264.8018, 261.6974, 
    240.8943, 237.8516, 242.8212, 244.7879, 245.4069, 245.3941, 245.5959, 
    245.6923,
  275.0287, 274.1216, 273.4573, 272.9691, 272.7603, 271.4397, 267.0188, 
    260.2139, 254.317, 254.306, 248.7426, 247.0641, 246.176, 245.8655, 
    245.4709,
  275.8333, 275.1405, 273.8792, 273.008, 272.7065, 272.395, 271.2053, 
    263.0855, 257.8555, 255.4659, 251.7533, 247.7025, 247.0538, 246.1781, 
    246.0484,
  276.2359, 275.1218, 274.0517, 273.2187, 272.6535, 272.4647, 271.7157, 
    269.3546, 260.3687, 253.4185, 250.428, 248.2521, 247.5569, 246.5829, 
    246.2887,
  276.0851, 275.226, 274.6212, 273.5784, 272.7204, 271.7506, 271.4021, 
    269.4075, 257.3737, 251.9681, 250.1451, 249.0115, 248.2686, 246.9071, 
    245.9997,
  275.1794, 274.1555, 273.6474, 272.9306, 272.0193, 270.6844, 268.1062, 
    262.9472, 254.0783, 251.9884, 254.1052, 250.5337, 249.5056, 248.4081, 
    246.6353,
  263.8649, 264.5756, 264.1212, 264.0512, 260.8704, 257.2018, 255.6522, 
    252.511, 248.7819, 239.5549, 238.5541, 239.5162, 235.3382, 235.1175, 
    231.3656,
  265.1851, 265.245, 264.8302, 264.1109, 259.8521, 254.9155, 252.9822, 
    250.1265, 247.3721, 245.4428, 241.5154, 245.0121, 244.7108, 232.2352, 
    229.1841,
  271.2666, 269.7313, 267.5161, 265.3408, 261.975, 250.8986, 249.4168, 
    248.7629, 246.7803, 246.3294, 246.107, 245.8245, 245.3283, 243.9384, 
    238.1039,
  273.867, 273.36, 272.557, 269.4612, 266.1053, 260.0972, 245.8576, 244.843, 
    245.5413, 245.392, 245.5036, 244.9079, 244.2091, 243.6959, 241.9912,
  274.4067, 273.5294, 273.1265, 272.7211, 269.0633, 265.5799, 262.9719, 
    242.564, 238.9225, 242.4482, 244.6405, 244.8008, 244.2866, 244.1396, 
    244.1299,
  275.1111, 274.1438, 273.4511, 272.9801, 272.7119, 271.0701, 267.4582, 
    261.1193, 254.5889, 253.799, 248.2499, 246.0312, 245.0869, 243.6823, 
    243.3546,
  275.9305, 275.2438, 273.9271, 273.0054, 272.7346, 272.4095, 271.037, 
    263.08, 256.7528, 255.4013, 251.3748, 246.533, 245.5281, 243.746, 243.1948,
  276.2755, 275.1885, 274.0504, 273.1809, 272.6893, 272.5022, 271.7405, 
    268.6928, 258.1267, 251.5373, 248.6592, 246.5094, 245.4748, 243.7554, 
    243.219,
  276.1713, 275.3016, 274.6462, 273.5558, 272.7823, 271.7881, 271.5359, 
    269.2523, 254.7341, 249.272, 247.3541, 246.2238, 245.4281, 243.993, 
    243.0918,
  275.277, 274.1682, 273.5616, 272.9324, 272.062, 271.104, 268.588, 260.9873, 
    250.4657, 248.7352, 250.6692, 247.0278, 246.6107, 245.5358, 244.4229,
  264.9955, 265.2259, 264.1137, 263.3201, 261.7794, 260.7383, 261.0329, 
    258.404, 255.7749, 248.2613, 244.2262, 243.0608, 236.9497, 236.0605, 
    235.226,
  267.2143, 266.0282, 264.9137, 263.5848, 261.4948, 260.1719, 259.2984, 
    257.0688, 254.0924, 250.9866, 246.2688, 247.2402, 245.7505, 233.046, 
    232.3322,
  271.8588, 269.9702, 267.8288, 264.2735, 262.334, 256.4315, 256.3895, 
    255.7337, 252.3498, 250.6424, 249.1399, 248.1996, 246.7401, 244.6214, 
    238.5482,
  273.8374, 273.3841, 272.6489, 269.5504, 266.206, 263.713, 251.0067, 
    249.4351, 249.3361, 249.0392, 248.0875, 246.4161, 245.5191, 244.1981, 
    241.7343,
  274.4969, 273.504, 273.0948, 272.8323, 268.6993, 267.2382, 264.4823, 
    245.3517, 242.3009, 245.5678, 246.6161, 245.9769, 245.2654, 244.806, 
    244.7643,
  275.2175, 274.1355, 273.4511, 272.9596, 272.6024, 270.835, 267.8789, 
    262.4724, 257.5152, 255.7381, 250.5105, 247.261, 245.8129, 244.071, 
    243.4138,
  276.0266, 275.3433, 274.004, 272.9834, 272.7181, 272.384, 270.8119, 
    264.898, 260.9588, 258.3773, 253.8029, 247.5505, 245.8867, 243.5254, 
    242.8596,
  276.3087, 275.3611, 274.0876, 273.1459, 272.6923, 272.5045, 271.7059, 
    268.8931, 260.0093, 252.8994, 250.0553, 247.1663, 245.4886, 243.119, 
    242.2569,
  276.2038, 275.3493, 274.6462, 273.5443, 272.7915, 271.7788, 271.5334, 
    269.0077, 255.1479, 249.8213, 247.6924, 246.5629, 244.8571, 243.0098, 
    241.8183,
  275.2642, 274.2666, 273.7536, 272.9352, 272.0454, 271.2556, 268.954, 
    260.0207, 249.9538, 248.5914, 250.5425, 247.1413, 245.6896, 244.2763, 
    243.1654,
  263.5825, 264.3999, 262.9669, 262.4062, 260.4833, 259.3706, 260.1083, 
    259.0638, 258.4248, 253.3089, 252.4293, 252.5663, 248.2325, 246.5484, 
    243.7915,
  267.3286, 264.9192, 263.6924, 262.0604, 259.7216, 259.0504, 259.2169, 
    258.1284, 257.5, 257.1385, 254.9183, 255.8457, 253.0741, 243.071, 240.6434,
  272.2733, 270.6076, 268.5581, 265.2131, 262.462, 257.4176, 257.9413, 
    257.3614, 255.7427, 255.8909, 256.1127, 254.7558, 252.1089, 248.9265, 
    244.0969,
  273.8353, 273.4185, 272.8547, 270.8642, 267.5674, 264.331, 253.5382, 
    252.8448, 252.295, 253.3237, 253.554, 252.5275, 250.5606, 247.6469, 
    244.6033,
  274.5991, 273.4813, 273.0566, 272.8658, 270.8212, 269.2035, 266.1864, 
    253.6379, 250.9117, 250.0441, 251.7993, 251.5095, 249.3261, 247.2984, 
    245.2198,
  275.3148, 274.1438, 273.4411, 272.9208, 272.7094, 271.5736, 268.5692, 
    264.4291, 259.9037, 259.0979, 254.2649, 251.0666, 248.7276, 245.9033, 
    243.8956,
  276.0823, 275.3646, 274.0669, 272.9529, 272.7083, 272.3662, 270.7464, 
    264.5563, 260.6283, 260.9341, 257.0399, 250.9648, 247.8986, 244.9726, 
    243.1361,
  276.2759, 275.3832, 274.0843, 273.0824, 272.6681, 272.4615, 271.5698, 
    267.9058, 259.1176, 255.0396, 252.9162, 249.1947, 247.1914, 243.8483, 
    242.6329,
  276.1533, 275.31, 274.6003, 273.4838, 272.7516, 271.6961, 271.2931, 
    267.6764, 254.9886, 250.8088, 249.3108, 247.9535, 245.6317, 243.4237, 
    242.5557,
  275.1654, 274.2593, 273.7552, 272.8694, 271.9716, 271.1754, 269.0087, 
    260.5956, 250.3057, 248.6398, 250.6495, 247.3095, 246.092, 244.2492, 
    244.4112,
  263.8031, 265.2842, 263.5369, 262.303, 259.5475, 256.9249, 257.624, 
    255.3058, 253.4595, 246.4843, 246.8529, 249.7597, 247.2273, 246.686, 
    244.7404,
  269.4368, 268.1623, 266.9151, 264.9341, 261.2884, 259.7237, 257.8944, 
    255.0329, 253.4016, 252.0505, 250.7067, 253.717, 253.0289, 245.5247, 
    244.2104,
  272.3623, 271.0725, 269.4193, 267.8227, 264.6574, 258.9158, 259.0899, 
    257.5557, 255.0888, 253.8287, 254.2215, 254.4885, 254.1036, 253.0023, 
    248.3423,
  273.8203, 273.4078, 272.9094, 271.4865, 268.7131, 265.3005, 257.2347, 
    255.3661, 254.8028, 254.869, 254.3204, 254.0276, 253.3793, 252.6512, 
    249.8041,
  274.624, 273.4536, 273.0197, 272.795, 271.4158, 270.0712, 266.4003, 
    254.8598, 252.0357, 254.8757, 254.8812, 254.593, 253.6512, 252.4273, 
    250.8394,
  275.2762, 274.093, 273.4393, 272.8941, 272.6173, 271.9505, 269.0592, 
    266.264, 263.4205, 262.8775, 258.4525, 256.1432, 254.4029, 251.202, 
    248.5834,
  276.009, 275.2168, 273.9904, 272.9178, 272.6826, 272.3512, 270.8353, 
    265.511, 263.3983, 264.068, 260.5847, 256.5061, 253.8201, 249.9697, 
    247.874,
  276.2372, 275.3018, 274.0043, 273.0042, 272.6408, 272.4206, 271.3439, 
    267.3368, 259.9227, 258.4836, 256.8915, 254.6512, 252.3237, 248.5743, 
    246.6039,
  276.1558, 275.3061, 274.5764, 273.425, 272.6686, 271.5267, 270.7758, 
    265.9448, 254.701, 253.6314, 253.486, 252.5813, 249.8839, 246.7316, 
    244.3254,
  275.1599, 274.2403, 273.6919, 272.7567, 271.8, 270.6489, 267.9908, 260.307, 
    250.7682, 249.219, 252.7812, 250.5016, 248.8779, 246.6514, 244.8548,
  267.1424, 267.9669, 265.3858, 266.6588, 264.9429, 263.1674, 263.1456, 
    261.1554, 258.0447, 249.1245, 248.8381, 252.0096, 249.1107, 248.789, 
    246.9653,
  267.4896, 265.251, 263.6689, 265.7778, 264.2351, 263.9926, 263.2695, 
    261.5181, 259.613, 254.9712, 253.2319, 255.0115, 253.2441, 245.5741, 
    245.156,
  272.221, 270.7922, 267.0637, 263.6399, 263.7311, 260.9674, 261.9909, 
    261.8249, 260.479, 258.3517, 256.8728, 255.6349, 253.0218, 251.2462, 
    247.6648,
  273.7779, 273.3471, 272.8748, 270.1732, 265.0824, 263.5508, 257.3059, 
    257.479, 257.1919, 256.7188, 255.3191, 253.265, 252.8122, 251.8867, 
    249.4706,
  274.6696, 273.4064, 272.9418, 272.7224, 270.0966, 268.7296, 265.1359, 
    249.7842, 253.9555, 254.853, 256.1656, 254.9329, 253.3023, 252.5966, 
    251.3092,
  275.3244, 274.0476, 273.3791, 272.838, 272.5544, 271.637, 268.0198, 
    264.3112, 260.7745, 261.9682, 258.6468, 256.4109, 254.6471, 252.4419, 
    250.721,
  276.0431, 275.1699, 273.946, 272.8661, 272.6189, 272.2878, 270.6479, 
    263.8739, 261.0585, 262.6249, 260.8775, 256.6653, 254.6033, 252.4144, 
    250.4467,
  276.2457, 275.3409, 274.0368, 272.9942, 272.6259, 272.3626, 270.9984, 
    265.94, 258.2297, 257.0221, 257.4212, 256.0852, 254.5398, 251.6431, 
    249.4879,
  276.2083, 275.3754, 274.6222, 273.4154, 272.6047, 271.3571, 270.5294, 
    264.9535, 254.7088, 253.1449, 255.3978, 255.2109, 253.5037, 250.1208, 
    247.0838,
  275.2138, 274.2533, 273.6327, 272.6792, 271.6836, 270.4805, 268.0692, 
    262.2862, 251.2436, 246.6118, 253.7504, 254.664, 252.854, 249.5261, 
    248.0045,
  262.1857, 263.5632, 257.3104, 262.0073, 259.6715, 259.4481, 262.0602, 
    261.5788, 260.7632, 255.9426, 255.6046, 255.4745, 252.4488, 251.924, 
    249.8085,
  263.2982, 261.2001, 259.7246, 260.2074, 257.6928, 259.5024, 261.3029, 
    260.9213, 260.7875, 258.5679, 257.1983, 257.9873, 257.4361, 250.7382, 
    248.8446,
  272.0396, 270.5219, 266.617, 263.1595, 260.2078, 257.9544, 260.8681, 
    261.2595, 260.7289, 258.3516, 258.0365, 258.0299, 256.0835, 254.7561, 
    251.3174,
  273.706, 273.3096, 272.8968, 270.9175, 267.6271, 266.1137, 261.4441, 
    259.5063, 258.9954, 257.6004, 254.9595, 254.0759, 253.9671, 253.5073, 
    252.2706,
  274.7224, 273.369, 272.9245, 272.7319, 271.5612, 270.9571, 268.831, 
    260.6085, 255.3098, 253.8217, 254.4495, 254.2315, 252.8436, 254.4976, 
    253.0728,
  275.4049, 274.06, 273.4034, 272.8716, 272.6756, 272.1504, 270.1937, 
    266.9146, 261.5025, 259.469, 255.1971, 254.6185, 253.8182, 252.7414, 
    251.4984,
  276.1184, 275.1522, 273.9608, 272.9046, 272.668, 272.3263, 271.3326, 
    265.7506, 262.3054, 261.8685, 255.8277, 252.5963, 253.648, 253.0656, 
    251.39,
  276.2591, 275.3644, 274.0893, 273.0665, 272.6857, 272.3806, 271.0129, 
    266.9547, 261.26, 257.8759, 252.4971, 250.5327, 252.7698, 251.8198, 
    250.353,
  276.2415, 275.3969, 274.6282, 273.4016, 272.5833, 271.1956, 270.4702, 
    265.5824, 259.4849, 255.3893, 250.6094, 250.4415, 251.4694, 250.5604, 
    248.6974,
  275.2505, 274.2539, 273.6232, 272.6347, 271.5634, 270.155, 267.5437, 
    261.975, 256.8417, 249.8201, 248.0475, 250.7348, 251.7596, 250.44, 
    249.3105,
  258.4344, 260.9731, 257.2294, 260.4416, 259.7751, 260.0849, 261.7463, 
    261.1169, 261.334, 260.0338, 261.1302, 261.9497, 260.5061, 259.0499, 
    254.7351,
  262.2694, 263.4084, 262.0828, 261.5349, 260.1939, 261.5663, 261.8733, 
    261.069, 260.5547, 260.3381, 261.4746, 262.8926, 261.9741, 256.0568, 
    253.4842,
  271.8927, 270.835, 268.9024, 265.9787, 262.0673, 257.4507, 261.7218, 
    261.7706, 260.7203, 258.9812, 260.5033, 261.4428, 259.9645, 258.1269, 
    254.513,
  273.652, 273.376, 272.9453, 271.8251, 266.8979, 260.5696, 255.3078, 
    257.6251, 258.5, 257.0389, 257.6931, 258.0309, 257.7903, 257.6828, 256.103,
  274.7381, 273.3647, 272.954, 272.7441, 271.8675, 270.2811, 261.6538, 
    254.0173, 254.7205, 253.8758, 254.8311, 255.2373, 256.17, 257.851, 
    257.3705,
  275.3899, 274.0854, 273.4175, 272.855, 272.6898, 272.1112, 267.9173, 
    263.7554, 259.8426, 257.746, 252.8675, 255.5897, 257.4579, 257.7432, 
    254.8511,
  276.1306, 275.1176, 273.8907, 272.8391, 272.6297, 272.2529, 271.0593, 
    263.7872, 260.0479, 258.0887, 253.4827, 252.7997, 256.3466, 253.9359, 
    252.0447,
  276.2624, 275.3151, 274.0388, 273.0327, 272.6656, 272.3394, 270.6542, 
    266.2478, 259.4254, 256.1223, 251.6298, 251.0361, 250.0601, 249.4072, 
    248.4128,
  276.2375, 275.3737, 274.599, 273.3581, 272.5342, 271.1265, 270.3139, 
    265.976, 258.5338, 253.4728, 250.9926, 248.723, 248.3202, 247.5968, 
    247.4788,
  275.2787, 274.2278, 273.4866, 272.4801, 271.5398, 270.2581, 268.1623, 
    263.8378, 258.6569, 252.456, 248.2429, 248.7706, 247.8689, 247.8456, 
    247.5572,
  259.7058, 261.1056, 257.6552, 258.4177, 256.6455, 257.4155, 259.9093, 
    257.7872, 256.2256, 250.515, 252.9295, 255.707, 252.831, 251.6681, 
    247.7207,
  264.9595, 262.088, 258.8499, 258.6729, 255.6329, 258.9966, 260.4536, 
    259.1279, 257.493, 253.325, 252.6293, 255.7331, 254.5401, 247.491, 244.846,
  271.8166, 269.8803, 267.4335, 264.0962, 259.7693, 256.2852, 262.9379, 
    261.3481, 260.0744, 254.4971, 254.9585, 255.2066, 254.4194, 252.9465, 
    248.9747,
  273.6327, 273.3631, 272.9474, 271.623, 267.6553, 263.5656, 261.6033, 
    260.8553, 260.8186, 256.374, 253.9565, 256.0721, 254.8823, 252.445, 
    250.7816,
  274.7569, 273.3445, 272.9324, 272.7119, 272.0568, 271.1628, 267.9552, 
    261.8599, 260.2993, 258.4151, 254.4944, 255.7552, 254.8231, 253.5162, 
    256.3385,
  275.3894, 274.1261, 273.4017, 272.8449, 272.675, 272.2033, 270.7759, 
    268.4927, 266.8408, 263.631, 255.0236, 256.1459, 253.5707, 252.0308, 
    249.6893,
  276.153, 275.1748, 273.8932, 272.8134, 272.6456, 272.2764, 271.6909, 
    269.7314, 268.2711, 266.0963, 259.1581, 254.0547, 254.1403, 248.7711, 
    247.1146,
  276.279, 275.3289, 274.0587, 273.0063, 272.702, 272.3687, 271.2124, 
    270.3751, 268.7959, 266.8877, 262.062, 255.4505, 252.973, 250.8143, 245.61,
  276.2724, 275.404, 274.6096, 273.3022, 272.5128, 271.2377, 271.1745, 
    270.0761, 269.0455, 267.4041, 263.4937, 257.7619, 253.5397, 248.6838, 
    245.7953,
  275.3858, 274.2307, 273.2744, 272.2604, 271.4167, 270.1598, 270.1835, 
    269.6389, 269.3486, 267.7412, 264.9632, 260.0364, 255.1981, 250.6978, 
    247.614,
  260.9863, 262.0452, 263.2642, 266.5576, 265.7618, 265.8605, 266.7978, 
    264.6841, 258.6557, 244.744, 248.8865, 251.6571, 247.3335, 244.3564, 
    242.5595,
  263.595, 264.3477, 266.6391, 266.852, 265.2227, 266.2051, 266.7898, 
    263.9554, 262.2278, 253.2445, 247.3214, 253.2531, 252.5754, 241.5202, 
    239.4204,
  271.359, 270.061, 270.0178, 268.2882, 265.8099, 263.278, 266.666, 265.7747, 
    265.673, 260.6617, 254.9426, 253.2158, 252.502, 253.4588, 249.4222,
  273.5819, 273.3376, 272.98, 271.7115, 269.2344, 267.087, 263.3783, 260.826, 
    266.4007, 264.6834, 259.5202, 255.3742, 251.2305, 251.3448, 253.1336,
  274.7737, 273.3474, 272.9063, 272.665, 272.0522, 271.2673, 268.3827, 
    263.4547, 264.4885, 266.3118, 262.734, 259.9228, 253.3173, 250.21, 
    251.9469,
  275.432, 274.2046, 273.4082, 272.8088, 272.6144, 272.1255, 270.6111, 
    268.6709, 267.2524, 267.6553, 264.9007, 263.0606, 258.7032, 252.9309, 
    249.8867,
  276.2002, 275.255, 274.0056, 272.8334, 272.6253, 272.2354, 271.6659, 
    269.3645, 268.3967, 267.3821, 266.9257, 263.8937, 261.5626, 256.2022, 
    250.999,
  276.3054, 275.3981, 274.188, 273.0528, 272.7045, 272.3165, 271.1436, 
    270.1968, 268.6414, 267.1378, 267.1686, 264.747, 262.9213, 258.9468, 
    253.635,
  276.3152, 275.466, 274.6428, 273.1729, 272.4177, 271.3076, 271.0369, 
    269.9436, 268.874, 268.1526, 267.6236, 265.1062, 263.9045, 260.9231, 
    255.9344,
  275.5091, 274.2908, 273.1305, 272.1653, 271.5407, 270.7185, 269.3578, 
    267.8631, 268.9192, 267.3148, 267.593, 266.3282, 264.1617, 261.5593, 
    258.1965,
  265.5417, 265.4822, 264.6469, 264.7645, 264.4337, 264.3524, 265.0551, 
    262.9978, 261.6739, 251.9585, 247.3303, 249.1224, 241.347, 242.0529, 
    241.3186,
  266.8918, 266.3261, 265.6113, 264.0049, 262.3565, 263.8398, 262.5971, 
    264.3973, 263.5671, 261.3013, 253.8942, 253.5723, 252.6275, 246.198, 
    242.8944,
  270.8498, 268.9745, 268.4733, 266.3998, 264.3658, 259.0244, 264.7567, 
    264.6234, 264.4154, 263.4218, 261.7052, 259.6595, 257.1063, 255.339, 
    250.5651,
  273.5719, 273.2484, 272.9484, 271.1633, 268.0238, 265.1742, 262.3501, 
    260.4583, 261.4829, 261.6714, 262.1048, 261.8765, 260.9571, 258.9045, 
    257.0824,
  274.7731, 273.3401, 272.871, 272.6008, 271.9781, 271.1168, 268.2034, 
    263.1129, 263.2772, 262.8518, 264.2169, 264.4014, 263.5137, 261.5324, 
    259.5701,
  275.4534, 274.2699, 273.4118, 272.7578, 272.565, 272.0803, 270.7373, 
    268.8297, 268.2267, 267.2323, 267.0002, 265.1614, 265.2484, 264.0807, 
    262.1324,
  276.2383, 275.3224, 274.0752, 272.8417, 272.6178, 272.2448, 271.7803, 
    270.1337, 269.4219, 268.5459, 267.5476, 266.1848, 265.8065, 265.2248, 
    264.0784,
  276.3238, 275.437, 274.2599, 273.1117, 272.7306, 272.3671, 271.4263, 
    271.0301, 270.3116, 269.7208, 269.3173, 267.3823, 266.7105, 266.16, 
    264.6792,
  276.2864, 275.4757, 274.6458, 273.188, 272.4611, 271.5988, 271.5252, 
    271.2316, 270.878, 270.442, 269.9639, 269.0146, 268.1187, 266.1773, 
    264.9194,
  275.4557, 274.3524, 273.5168, 272.3551, 271.7944, 271.4575, 271.4531, 
    270.9008, 271.2465, 270.7271, 270.57, 269.8804, 269.0902, 267.3554, 
    264.7454,
  266.2019, 263.4551, 259.8967, 257.9187, 254.3646, 254.9731, 257.5441, 
    258.0667, 258.8882, 257.9193, 259.4132, 260.1769, 259.3808, 258.9901, 
    259.9278,
  266.4654, 264.0808, 261.0669, 257.8975, 253.6301, 254.6518, 259.3762, 
    259.5687, 259.9939, 259.6373, 260.2663, 262.6188, 263.416, 262.0981, 
    261.5356,
  270.0049, 266.7931, 265.1737, 260.9676, 256.8026, 251.021, 259.209, 
    259.8879, 261.9698, 262.6302, 263.6709, 265.3318, 266.2931, 266.1531, 
    265.4285,
  273.5241, 273.0314, 272.7849, 270.1512, 264.8652, 259.46, 258.7143, 
    261.7816, 265.3589, 266.7007, 267.5973, 268.3289, 267.8181, 267.016, 
    266.085,
  274.7281, 273.3, 272.8342, 272.559, 272.0383, 271.0736, 268.2714, 265.0007, 
    266.4371, 268.1554, 269.8581, 269.3293, 267.917, 266.8658, 266.187,
  275.41, 274.2622, 273.3911, 272.7339, 272.5928, 272.1649, 271.4304, 
    269.5733, 270.1509, 270.5824, 270.3494, 268.2851, 267.0772, 266.325, 
    265.4037,
  276.2063, 275.2868, 274.0099, 272.8233, 272.6158, 272.3272, 271.9939, 
    271.3703, 271.5391, 270.9609, 268.3848, 266.7185, 265.8391, 264.9578, 
    264.2464,
  276.3009, 275.3725, 274.1819, 273.0979, 272.7378, 272.5067, 271.8294, 
    271.5897, 271.4664, 268.6506, 266.2915, 264.8777, 264.3805, 263.3425, 
    263.1761,
  276.226, 275.4112, 274.5942, 273.2854, 272.5484, 271.8077, 271.8352, 
    271.613, 269.4336, 267.0228, 265.4129, 263.2037, 262.2, 261.584, 261.7984,
  275.3311, 274.2928, 273.7339, 272.648, 271.9489, 271.7436, 271.5464, 
    268.4556, 266.6268, 262.6353, 264.5779, 262.0088, 260.7061, 260.2259, 
    260.1727,
  266.3993, 264.8229, 262.4151, 259.9966, 256.153, 254.4873, 256.1296, 
    252.8419, 251.5787, 249.7008, 251.9059, 255.6396, 257.6511, 259.7136, 
    256.879,
  267.5602, 266.8361, 263.6435, 260.4395, 255.8454, 254.9569, 256.748, 
    253.8224, 253.4495, 252.624, 254.2252, 258.9751, 261.2792, 257.8906, 
    254.7111,
  270.5204, 268.4767, 267.2751, 263.8799, 258.508, 254.4162, 258.8419, 
    257.946, 257.1099, 256.2344, 258.0056, 260.7807, 261.1384, 258.5388, 
    255.1245,
  273.5143, 273.0942, 272.782, 270.6721, 265.863, 259.8291, 256.4024, 
    257.2772, 258.5237, 258.5493, 261.1462, 262.3574, 260.6917, 259.1396, 
    256.3559,
  274.6588, 273.2776, 272.8321, 272.5482, 272.022, 270.6782, 265.8167, 
    259.1491, 257.7156, 263.2297, 266.0291, 263.7159, 261.8839, 260.6471, 
    259.106,
  275.326, 274.2516, 273.3813, 272.7247, 272.5802, 272.1651, 271.4685, 
    267.5372, 265.2751, 266.7055, 267.0455, 264.8725, 263.5034, 261.5472, 
    258.9412,
  276.1107, 275.2331, 273.9805, 272.8108, 272.6063, 272.3226, 272.0306, 
    270.7838, 268.6712, 268.3344, 267.3353, 265.2457, 263.4985, 261.2653, 
    258.4838,
  276.2505, 275.3093, 274.1365, 273.0864, 272.7051, 272.5425, 271.8624, 
    271.1024, 268.9734, 268.1652, 267.2315, 264.8053, 263.0564, 260.3278, 
    258.1669,
  276.1819, 275.382, 274.5517, 273.2547, 272.5038, 271.7691, 271.4991, 
    270.4236, 269.3712, 268.9623, 268.14, 264.9631, 262.5455, 259.6313, 
    257.8102,
  275.3102, 274.2921, 273.7039, 272.3697, 271.2725, 270.8069, 270.2346, 
    269.3723, 269.4732, 267.6749, 268.1039, 264.4904, 261.4473, 258.6849, 
    256.5536,
  267.2129, 266.4179, 266.3036, 266.3236, 264.761, 263.5384, 263.1969, 
    259.9304, 256.9395, 250.5798, 249.7067, 251.5012, 248.9693, 247.6992, 
    246.303,
  266.9453, 266.8938, 266.7766, 266.4668, 264.8014, 263.5108, 263.9352, 
    260.4788, 257.9661, 255.7283, 254.0449, 254.9085, 253.7298, 249.2047, 
    249.0615,
  270.9435, 269.5103, 268.6579, 267.6676, 266.2557, 262.1836, 264.6854, 
    263.1667, 258.6942, 257.8922, 258.057, 257.9426, 257.4608, 258.2432, 
    257.3627,
  273.5515, 273.2763, 272.8959, 271.5415, 269.2726, 265.6631, 262.1785, 
    262.2612, 261.1139, 260.687, 260.8093, 260.4912, 261.3536, 260.1084, 
    256.9872,
  274.5965, 273.2674, 272.8303, 272.5389, 272.0511, 271.101, 268.0919, 
    261.5843, 261.7336, 263.4556, 264.8994, 263.8416, 262.6569, 258.5551, 
    257.0297,
  275.2921, 274.2962, 273.3766, 272.7104, 272.5596, 272.1391, 271.5977, 
    269.4355, 266.737, 265.6916, 266.932, 265.336, 260.8862, 257.6148, 
    256.3272,
  276.0676, 275.2208, 273.9787, 272.7985, 272.5878, 272.2915, 272.0157, 
    270.8759, 266.318, 267.2131, 265.7785, 261.515, 257.9507, 256.1929, 
    254.9878,
  276.2493, 275.2842, 274.1346, 273.0748, 272.6664, 272.5336, 271.8361, 
    271.0826, 268.5772, 266.6296, 261.4157, 257.4402, 255.7207, 254.058, 
    253.3753,
  276.1764, 275.3983, 274.5351, 273.1638, 272.4228, 271.7492, 271.3893, 
    270.6244, 268.5959, 265.8481, 263.1521, 256.2294, 253.8288, 252.4151, 
    252.138,
  275.3494, 274.2855, 273.5663, 272.1728, 271.0564, 270.4362, 269.7793, 
    267.9533, 265.9419, 260.6219, 262.2389, 255.8159, 252.5187, 251.137, 
    250.2212,
  262.8116, 263.7238, 263.5239, 266.1033, 265.8125, 267.4249, 268.3117, 
    268.0323, 266.8921, 263.9668, 261.3156, 260.0544, 256.2135, 253.7088, 
    249.8924,
  264.7351, 265.0204, 267.162, 268.6396, 267.9943, 269.3922, 269.869, 
    268.8982, 267.2636, 263.9164, 262.7429, 261.8089, 259.7289, 253.9366, 
    251.9368,
  270.9826, 269.8822, 269.9982, 270.8331, 270.4888, 269.6832, 270.0133, 
    269.3829, 267.2505, 264.7677, 264.0781, 262.8909, 261.853, 260.557, 
    257.5813,
  273.5363, 273.3615, 272.9518, 272.1184, 271.9132, 271.4777, 269.7739, 
    268.7077, 266.9694, 265.6714, 264.1934, 263.3131, 263.3385, 262.3562, 
    260.9053,
  274.5902, 273.3163, 272.8701, 272.57, 272.1448, 271.8206, 271.2935, 
    267.836, 266.7484, 265.9029, 266.8708, 266.4944, 265.3385, 263.6912, 
    262.0641,
  275.3409, 274.3767, 273.4104, 272.7408, 272.5854, 272.1484, 271.7305, 
    270.6253, 269.6273, 268.6986, 267.7667, 267.2269, 266.1969, 264.4545, 
    261.5033,
  276.0729, 275.2582, 274.0258, 272.8474, 272.6298, 272.3105, 272.0412, 
    271.2921, 268.3111, 267.1225, 266.311, 266.8275, 265.0633, 262.7144, 
    257.6987,
  276.2778, 275.3125, 274.1872, 273.1209, 272.6943, 272.56, 271.8442, 
    271.3427, 269.3281, 268.3778, 267.9535, 266.2452, 264.2059, 258.5146, 
    253.6002,
  276.1947, 275.4501, 274.5703, 273.1221, 272.4275, 271.7879, 271.6434, 
    270.7175, 269.5258, 269.1759, 268.848, 264.6074, 258.74, 253.177, 251.7335,
  275.3944, 274.3257, 273.5646, 272.3135, 271.6842, 271.115, 270.2506, 
    269.4171, 269.8113, 268.0223, 266.8225, 259.7879, 253.1116, 249.9035, 
    248.0187,
  259.617, 261.6701, 261.6107, 263.0143, 262.7346, 264.7657, 266.5186, 
    266.7595, 265.798, 265.0623, 264.5154, 265.0399, 263.615, 264.5858, 
    263.6672,
  263.7336, 263.8291, 263.4698, 263.0299, 263.3061, 267.0608, 267.1713, 
    266.0974, 265.534, 264.3478, 264.3748, 264.8581, 265.3761, 265.4543, 
    265.2933,
  271.1048, 269.2915, 268.0737, 266.0732, 267.8657, 266.5052, 268.9042, 
    266.4183, 265.3549, 264.8282, 265.6929, 266.6711, 268.4174, 268.3392, 
    267.3625,
  273.4943, 273.3468, 272.9321, 271.6769, 269.6162, 269.8442, 268.3898, 
    267.8751, 267.0023, 266.6609, 267.658, 268.9568, 269.277, 268.867, 
    265.9005,
  274.5499, 273.3209, 272.846, 272.5464, 272.1554, 271.5721, 270.7778, 
    267.7699, 267.7715, 269.2151, 270.2438, 269.9932, 269.7901, 268.9272, 
    265.4212,
  275.3075, 274.335, 273.383, 272.7162, 272.5805, 272.1526, 271.7642, 
    270.8733, 270.1254, 270.5622, 270.054, 269.8269, 269.7856, 268.3693, 
    262.8107,
  276.0091, 275.23, 274.0327, 272.8455, 272.6339, 272.3208, 272.0685, 
    271.5686, 270.5842, 269.5874, 269.2609, 269.4967, 269.6941, 266.2338, 
    259.1068,
  276.2553, 275.3116, 274.1872, 273.1247, 272.6977, 272.5955, 271.8853, 
    271.5477, 270.5142, 269.5946, 269.1627, 270.0543, 268.5354, 261.1888, 
    254.0797,
  276.1785, 275.4548, 274.582, 273.1174, 272.4399, 271.8055, 271.7159, 
    271.027, 270.2369, 270.0018, 270.5858, 269.8649, 264.4836, 254.758, 
    250.7329,
  275.3685, 274.3427, 273.612, 272.3361, 271.7043, 271.3492, 270.6894, 
    269.6766, 269.7783, 269.4792, 270.5466, 267.5731, 257.4786, 250.6939, 
    247.3719,
  258.4252, 260.031, 259.2716, 259.615, 257.2449, 257.3978, 260.6736, 
    260.7722, 262.5562, 263.235, 264.0945, 264.9583, 264.7411, 265.1204, 
    265.3149,
  263.2697, 262.9278, 260.8537, 259.3682, 258.0883, 262.9023, 264.9879, 
    264.3543, 265.3988, 265.6366, 265.8434, 266.0692, 265.2705, 265.0094, 
    266.2041,
  271.6316, 269.8479, 267.6798, 265.4147, 266.7875, 265.343, 268.2636, 
    267.6609, 266.8917, 266.172, 265.3649, 265.5666, 266.7293, 268.3651, 
    269.1781,
  273.5672, 273.3848, 272.9128, 272.0577, 269.8145, 268.2768, 266.6955, 
    269.1433, 267.2819, 264.6721, 265.9717, 267.3679, 268.8501, 269.6667, 
    269.4095,
  274.4646, 273.2972, 272.8665, 272.5358, 272.2183, 271.2994, 270.1184, 
    266.3055, 266.9165, 268.241, 269.7182, 269.3956, 269.9538, 269.928, 
    269.2636,
  275.2054, 274.2393, 273.3726, 272.7032, 272.5961, 272.1695, 271.7753, 
    270.6137, 269.5846, 270.0434, 270.3066, 270.2265, 270.1563, 270.0305, 
    268.2637,
  275.9168, 275.1581, 273.9846, 272.8251, 272.6231, 272.3247, 272.0775, 
    271.6254, 271.0108, 270.6276, 270.5758, 270.4575, 270.2506, 269.756, 
    266.062,
  276.2155, 275.2754, 274.1617, 273.1299, 272.6911, 272.6228, 271.9098, 
    271.6327, 271.2587, 270.8666, 270.6863, 270.5782, 270.3973, 268.6475, 
    264.1252,
  276.1247, 275.4267, 274.5904, 273.1517, 272.4518, 271.8257, 271.7972, 
    271.5036, 271.3151, 271.2498, 271.2787, 270.742, 270.0799, 267.0079, 
    261.7885,
  275.2435, 274.3284, 273.6839, 272.4246, 271.8298, 271.6006, 271.3786, 
    271.1015, 271.3025, 271.5259, 271.402, 270.8646, 269.0205, 265.0959, 
    259.4162,
  257.5888, 259.249, 258.6602, 259.5597, 257.4293, 257.5934, 258.9878, 
    257.3445, 257.7643, 257.8221, 259.6331, 260.3739, 260.8979, 262.1771, 
    262.7328,
  263.003, 261.355, 259.1487, 258.0856, 255.8516, 260.89, 262.8879, 261.4229, 
    261.0563, 261.4636, 262.2603, 263.2755, 263.8958, 263.5149, 264.3643,
  272.0959, 270.6219, 267.6503, 264.2244, 260.5131, 260.5348, 267.2551, 
    265.2237, 264.1271, 263.8455, 263.8938, 264.6171, 265.3148, 265.8885, 
    266.3225,
  273.6465, 273.4414, 272.9228, 272.3669, 268.9817, 264.5754, 263.5533, 
    268.1522, 267.1821, 266.1211, 265.4735, 264.8074, 265.9664, 266.4769, 
    266.7333,
  274.3867, 273.3031, 272.9027, 272.56, 272.2984, 271.0958, 269.2155, 
    264.7191, 265.6899, 266.723, 268.381, 265.9598, 266.2354, 267.2864, 
    266.4668,
  275.1317, 274.1917, 273.3565, 272.7092, 272.6118, 272.1967, 271.77, 
    269.9078, 267.3834, 267.9051, 268.062, 266.7773, 266.9095, 267.6568, 
    268.0326,
  275.8184, 275.0723, 273.9062, 272.7942, 272.5995, 272.3145, 272.0641, 
    271.6178, 270.1506, 268.0752, 267.6865, 267.412, 268.019, 268.2186, 
    268.5048,
  276.1429, 275.1862, 274.0844, 273.0858, 272.6561, 272.6176, 271.8957, 
    271.6, 270.5037, 268.6958, 268.0318, 267.7694, 267.7599, 267.8638, 
    268.5667,
  276.0309, 275.336, 274.5472, 273.2074, 272.4568, 271.8196, 271.7946, 
    271.3665, 270.2293, 269.7611, 270.05, 268.5174, 268.6187, 268.6992, 
    268.6146,
  275.0351, 274.1876, 273.6457, 272.469, 271.3294, 270.8208, 270.5136, 
    270.366, 270.5427, 270.418, 270.8947, 270.3648, 269.7429, 269.3161, 
    268.9783,
  257.0275, 258.5514, 258.3503, 259.259, 255.6421, 256.0599, 257.1558, 
    254.5353, 252.4643, 252.0817, 252.9886, 253.4942, 252.2196, 251.8752, 
    251.4125,
  262.1255, 259.1576, 257.566, 256.2385, 254.1121, 259.2172, 260.8375, 
    257.0621, 254.3383, 253.3211, 254.0905, 255.0885, 254.3876, 252.3958, 
    253.3374,
  272.3159, 270.1377, 266.5883, 261.3094, 255.0662, 253.5243, 265.3074, 
    261.4197, 258.0418, 255.3024, 256.1754, 256.3998, 255.5538, 255.6169, 
    256.1923,
  273.6753, 273.4559, 272.9145, 272.3814, 267.5505, 259.4362, 257.2731, 
    265.8293, 263.6035, 260.6438, 259.4542, 260.1441, 260.2647, 260.9674, 
    261.1835,
  274.3521, 273.2971, 272.8977, 272.552, 272.3235, 270.1896, 266.0356, 
    260.2221, 261.281, 263.6058, 265.4756, 264.2286, 263.8584, 263.9111, 
    263.8571,
  275.1205, 274.1603, 273.3127, 272.6843, 272.5912, 272.2212, 271.7672, 
    269.5705, 263.9951, 264.2016, 264.8233, 265.9051, 265.9119, 265.8243, 
    265.6363,
  275.7404, 274.9904, 273.8264, 272.7334, 272.5503, 272.2773, 272.0437, 
    271.6192, 270.1424, 266.6673, 267.1958, 267.15, 266.9965, 266.7928, 
    266.4106,
  276.0725, 275.0794, 273.957, 272.9725, 272.5621, 272.5634, 271.8296, 
    271.5604, 269.8047, 264.8181, 265.9496, 266.0219, 266.5884, 266.7796, 
    266.6035,
  275.9512, 275.2238, 274.426, 273.0844, 272.3155, 271.6818, 271.6352, 
    270.6942, 267.557, 266.058, 268.524, 266.6438, 266.5421, 266.1188, 
    266.0224,
  274.8577, 273.7884, 273.189, 271.87, 269.8705, 267.3199, 263.3215, 
    260.2935, 263.9553, 264.7719, 267.8375, 267.3782, 265.3396, 265.6891, 
    266.1124,
  259.4874, 260.3489, 260.0607, 260.6207, 258.1136, 258.5215, 259.4492, 
    256.8496, 255.2615, 253.5978, 253.1339, 254.1424, 251.9299, 251.2668, 
    249.3127,
  264.7248, 261.2207, 259.3977, 258.1694, 255.9321, 260.6499, 261.5324, 
    258.4799, 255.8772, 255.0491, 255.4855, 256.032, 254.2177, 250.5154, 
    249.41,
  272.4667, 270.4749, 268.138, 262.7576, 257.7968, 255.8427, 264.501, 
    261.0665, 258.1753, 255.5597, 257.062, 255.9462, 254.6749, 252.8855, 
    251.1701,
  273.6537, 273.4246, 272.8888, 272.3383, 268.2645, 259.7957, 256.8864, 
    264.7908, 262.5665, 259.186, 257.9304, 257.5959, 255.7485, 255.1727, 
    253.3602,
  274.3622, 273.2783, 272.8531, 272.4986, 272.2487, 270.1461, 264.6422, 
    257.5705, 257.4815, 261.8367, 263.127, 260.0357, 257.8585, 255.9205, 
    254.2217,
  275.1409, 274.105, 273.2689, 272.6026, 272.5196, 272.1566, 271.6476, 
    268.0887, 262.0287, 259.6765, 261.6192, 262.3015, 262.5296, 262.2085, 
    261.5618,
  275.698, 274.9491, 273.7824, 272.6652, 272.5047, 272.2097, 271.9857, 
    271.5054, 269.9667, 266.1613, 264.7666, 264.5708, 264.0037, 263.5516, 
    263.4481,
  276.0386, 275.052, 273.8991, 272.8975, 272.4805, 272.4989, 271.7092, 
    271.3397, 268.252, 257.5721, 255.6352, 255.2609, 254.7744, 255.546, 
    255.9279,
  275.934, 275.1852, 274.4012, 273.0115, 272.2, 271.4745, 271.109, 269.5703, 
    264.6599, 261.1567, 264.9253, 255.1681, 253.7155, 253.0368, 253.9736,
  274.8053, 273.6943, 273.0626, 271.4397, 269.6807, 266.937, 261.257, 
    256.1098, 256.5564, 254.3773, 259.8407, 255.1988, 254.2038, 254.1245, 
    254.6224,
  259.5141, 261.1654, 260.3459, 261.2226, 258.3525, 259.1678, 260.1729, 
    258.8778, 257.5536, 255.5845, 255.6648, 256.19, 255.2811, 254.5789, 
    254.0363,
  266.2959, 264.1576, 261.4086, 259.7472, 256.5803, 261.6212, 262.9001, 
    259.8714, 258.1398, 257.2781, 257.8931, 257.9286, 256.5502, 253.8343, 
    253.7548,
  272.4223, 270.8537, 269.3261, 264.7105, 259.261, 257.2164, 265.0692, 
    262.4646, 260.332, 258.4662, 259.1959, 258.3904, 257.0011, 256.2332, 
    254.9445,
  273.6013, 273.3645, 272.8461, 272.1501, 268.0407, 260.9975, 257.7769, 
    265.1198, 263.6368, 260.6077, 260.5152, 259.7986, 258.459, 257.4841, 
    256.2206,
  274.4149, 273.2639, 272.8206, 272.4537, 272.1214, 269.8008, 265.3878, 
    259.2801, 260.284, 261.6211, 263.3521, 261.1851, 259.941, 258.5201, 
    257.692,
  275.1878, 274.0824, 273.2814, 272.547, 272.4554, 272.0885, 271.4568, 
    267.9007, 262.8261, 259.4322, 259.3258, 259.6316, 259.3914, 259.4344, 
    259.1372,
  275.7049, 274.961, 273.7905, 272.6389, 272.4855, 272.1635, 271.9305, 
    271.2973, 268.5481, 263.746, 261.4055, 260.8976, 261.3166, 260.4219, 
    258.4448,
  276.0548, 275.0782, 273.8936, 272.8578, 272.4012, 272.4135, 271.5116, 
    270.8107, 265.8189, 257.0833, 255.9784, 255.7599, 255.5085, 255.414, 
    254.4553,
  275.9485, 275.1709, 274.3975, 272.9061, 271.9755, 270.6125, 269.6284, 
    266.6776, 260.9843, 257.6153, 261.037, 251.4124, 251.9077, 250.9417, 
    250.0473,
  274.632, 273.3607, 272.6549, 270.164, 266.9894, 262.7599, 257.1188, 
    254.2197, 254.1043, 250.0492, 254.0388, 248.9429, 248.4425, 247.8214, 
    249.9206,
  260.796, 262.1544, 261.339, 261.3478, 258.1153, 257.1975, 259.3176, 
    257.425, 256.2739, 252.904, 254.3954, 255.1884, 252.9041, 251.3217, 
    250.406,
  266.4415, 264.3941, 262.2983, 259.9831, 258.5806, 262.2366, 262.5268, 
    258.3563, 255.8292, 254.1635, 255.9089, 257.3057, 255.8261, 251.7323, 
    251.7868,
  272.4471, 271.0953, 269.3868, 264.4872, 259.996, 257.3217, 264.6871, 
    261.4247, 258.3856, 254.4494, 256.9997, 256.9497, 255.4738, 254.8703, 
    253.2303,
  273.5941, 273.324, 272.8766, 271.9834, 268.0404, 261.2384, 258.039, 
    264.0443, 261.5656, 258.0464, 257.4809, 257.0085, 255.6166, 255.978, 
    255.1336,
  274.4369, 273.2235, 272.7759, 272.4095, 272.0542, 269.2909, 263.8752, 
    258.4258, 258.6143, 260.5052, 261.3456, 259.229, 257.4156, 256.4163, 
    255.4666,
  275.1595, 274.0287, 273.2364, 272.4724, 272.3992, 272.0071, 271.1864, 
    266.8506, 261.7724, 260.2104, 260.009, 259.4098, 258.5063, 257.5388, 
    256.2419,
  275.6602, 274.8771, 273.7101, 272.5669, 272.4286, 272.1033, 271.841, 
    270.6686, 266.4048, 261.8921, 260.0746, 259.0655, 258.9893, 258.2548, 
    257.6782,
  276.0289, 275.0295, 273.812, 272.7524, 272.2843, 272.2841, 270.9515, 
    269.4313, 260.9182, 255.7156, 255.9309, 256.4408, 256.9569, 256.6931, 
    256.4802,
  275.9472, 275.1302, 274.3533, 272.8402, 271.6504, 269.5731, 267.7792, 
    263.7655, 258.727, 255.7405, 257.1746, 251.2243, 250.9033, 251.2355, 
    252.024,
  274.7241, 273.4572, 272.4626, 269.4321, 266.0283, 261.0604, 256.0958, 
    253.3719, 252.2496, 248.136, 249.9594, 246.4073, 245.8501, 246.269, 
    248.3954,
  263.4989, 263.3398, 261.8231, 262.0274, 257.8688, 257.768, 258.7488, 
    256.4366, 255.8676, 252.6535, 253.2039, 253.7838, 249.4416, 248.0734, 
    245.8754,
  267.0827, 265.2071, 262.6913, 261.4232, 258.1365, 262.2015, 262.1362, 
    257.9399, 255.8908, 255.0891, 255.3784, 256.7192, 254.3219, 248.5182, 
    247.119,
  272.451, 270.9428, 268.8775, 263.3363, 261.0733, 258.4611, 264.5856, 
    261.3639, 258.0557, 255.0207, 257.904, 257.5777, 254.8938, 253.3579, 
    250.2575,
  273.5721, 273.2602, 272.8488, 271.4796, 267.2533, 262.3413, 258.5616, 
    263.2534, 261.552, 257.9155, 257.1779, 257.2753, 256.2173, 255.1175, 
    253.2411,
  274.4532, 273.1983, 272.7422, 272.3593, 271.8151, 268.1916, 264.1394, 
    258.3539, 255.9982, 259.3603, 260.9657, 258.2466, 257.5142, 256.5136, 
    254.437,
  275.1302, 273.9904, 273.1782, 272.4166, 272.3326, 271.9218, 270.5302, 
    265.0579, 257.7693, 255.862, 257.7806, 259.0048, 257.4879, 256.7572, 
    255.048,
  275.6414, 274.8176, 273.6585, 272.5386, 272.4031, 272.0599, 271.7022, 
    269.0381, 261.4911, 257.058, 257.2979, 256.6916, 257.0245, 256.4543, 
    255.8543,
  276.0158, 275.0313, 273.826, 272.7086, 272.2079, 272.1991, 270.4782, 
    268.2808, 258.4894, 252.9574, 252.0259, 254.1499, 256.9509, 256.2738, 
    255.87,
  275.9268, 275.0923, 274.3467, 272.751, 271.4554, 269.2531, 267.6261, 
    263.0736, 257.4825, 253.4946, 252.7164, 250.3784, 253.2791, 256.0321, 
    255.667,
  274.6565, 273.2935, 272.0197, 267.4762, 263.4888, 259.2328, 256.3286, 
    254.0592, 250.5184, 245.1722, 246.7389, 246.3779, 249.8736, 254.8152, 
    255.6954,
  266.3373, 266.6425, 265.4037, 264.2509, 260.6729, 259.5548, 260.6503, 
    257.1045, 257.9081, 255.2384, 255.9423, 256.2124, 252.0522, 249.1591, 
    245.8963,
  267.6804, 266.0492, 264.7731, 263.1618, 260.0432, 262.8686, 262.5864, 
    258.7665, 257.8704, 258.2169, 257.9663, 258.9186, 256.5894, 250.0502, 
    246.9382,
  272.5032, 270.5911, 267.9276, 263.9613, 260.9688, 257.9801, 263.8073, 
    261.2767, 258.46, 256.3954, 260.5186, 259.8492, 257.3042, 254.9141, 
    251.2141,
  273.5465, 273.2479, 272.8142, 270.6438, 264.8434, 260.1135, 256.3771, 
    261.8282, 260.6446, 257.8536, 257.6528, 257.7697, 257.5439, 256.4236, 
    254.116,
  274.4283, 273.152, 272.7228, 272.3288, 271.5332, 266.6365, 261.261, 
    256.9066, 257.0092, 258.378, 259.4753, 257.3059, 256.701, 257.0841, 
    255.8604,
  275.035, 273.9162, 273.1339, 272.3675, 272.2874, 271.85, 269.7927, 
    263.5756, 257.7074, 256.2779, 256.4518, 258.0962, 256.7837, 255.6284, 
    254.8566,
  275.5836, 274.743, 273.6097, 272.5254, 272.3928, 272.052, 271.638, 
    269.2792, 262.3379, 258.3854, 254.7232, 252.61, 253.5411, 253.7796, 
    253.8195,
  275.9731, 274.9892, 273.7829, 272.6283, 272.1349, 272.1322, 270.4541, 
    268.8469, 261.652, 255.8991, 252.0229, 250.4379, 248.7828, 248.5379, 
    249.281,
  275.8317, 274.9607, 274.2412, 272.6729, 269.8435, 266.8328, 267.0011, 
    265.2455, 261.0796, 256.8586, 252.3722, 248.3927, 246.4949, 245.0852, 
    245.5809,
  274.4431, 273.0766, 271.6979, 264.4708, 258.8762, 254.5939, 255.3477, 
    258.2135, 256.2619, 251.9028, 248.3932, 245.6276, 243.7844, 243.8903, 
    245.026,
  259.6546, 264.9276, 264.2466, 265.5115, 264.1454, 264.2561, 264.4707, 
    261.4751, 259.446, 255.9729, 254.1493, 252.4697, 247.8217, 247.4662, 
    247.7153,
  264.8755, 263.8149, 263.9841, 263.7193, 261.7851, 265.3572, 265.6127, 
    262.0249, 259.9664, 257.5606, 256.4327, 256.7001, 253.0992, 245.4035, 
    246.8122,
  272.469, 269.9156, 266.3132, 263.6126, 262.8212, 262.0798, 265.5292, 
    262.9896, 260.275, 258.5355, 259.9726, 258.1978, 252.7228, 250.5692, 
    248.3544,
  273.5057, 273.1756, 272.7606, 269.967, 265.6669, 262.8953, 260.6978, 
    262.5699, 260.7898, 258.136, 258.0731, 257.9555, 254.1638, 251.6912, 
    250.392,
  274.409, 273.0872, 272.6934, 272.2938, 271.1168, 266.7941, 262.5673, 
    256.7285, 255.7958, 257.4186, 257.4048, 256.8331, 255.4982, 254.0803, 
    250.6472,
  274.9618, 273.8338, 273.0737, 272.3082, 272.2294, 271.7341, 269.3999, 
    263.884, 259.5428, 258.0414, 256.6685, 256.7931, 257.0326, 256.5155, 
    252.1673,
  275.5247, 274.6684, 273.5151, 272.4604, 272.3508, 271.9934, 271.4946, 
    269.6836, 263.1716, 260.1623, 257.2824, 256.0438, 256.1754, 257.0407, 
    255.7919,
  275.9181, 274.8673, 273.6506, 272.5306, 272.0869, 271.8896, 269.5124, 268, 
    260.2725, 257.3715, 258.1045, 256.7015, 255.955, 255.922, 256.1066,
  275.7473, 274.8805, 274.1679, 272.6003, 267.7961, 264.0921, 262.4177, 
    259.2763, 255.2571, 254.4377, 259.0869, 257.6639, 255.9386, 254.9637, 
    254.1311,
  274.3489, 272.8357, 271.1656, 263.102, 256.7216, 252.5395, 251.4574, 
    252.7435, 252.1, 251.2443, 257.1728, 256.6649, 255.3224, 254.421, 254.3555,
  259.0945, 261.7176, 258.9331, 262.3412, 261.8521, 262.5234, 262.6436, 
    260.2773, 257.3482, 257.041, 256.6996, 257.4236, 256.8247, 256.4772, 
    255.4115,
  265.2934, 263.4417, 261.0409, 259.8875, 260.6419, 263.1209, 263.1836, 
    261.7594, 259.2524, 258.7539, 259.0265, 260.3337, 259.308, 254.7429, 
    254.2553,
  272.4167, 269.8807, 265.8751, 261.4167, 259.0481, 257.2587, 263.5735, 
    263.1762, 262.0529, 260.0014, 261.5132, 260.3712, 258.5004, 257.4, 
    254.1973,
  273.4343, 273.1357, 272.7513, 269.899, 263.7296, 261.4178, 259.0708, 
    263.3231, 262.9146, 260.6553, 260.218, 260.1214, 258.2664, 256.8474, 
    254.6212,
  274.3583, 273.0148, 272.653, 272.2453, 270.728, 266.1226, 263.6588, 
    259.9963, 259.432, 259.8407, 260.5202, 259.2833, 257.3143, 255.7999, 
    253.2124,
  274.9075, 273.7422, 272.9986, 272.2528, 272.1962, 271.5849, 269.2563, 
    265.2867, 262.5337, 261.9067, 261.0812, 259.9161, 257.447, 254.9089, 
    252.6388,
  275.4474, 274.6067, 273.422, 272.3856, 272.3193, 271.9774, 271.3371, 
    269.2808, 264.934, 263.2789, 261.3665, 258.8653, 256.4193, 253.6407, 
    251.3281,
  275.9022, 274.809, 273.5488, 272.4389, 272.015, 271.5105, 269.048, 
    267.7071, 262.5303, 261.208, 259.9829, 258.2953, 255.9328, 253.0441, 
    250.7436,
  275.7697, 274.8874, 274.1478, 272.3553, 265.9788, 262.7239, 260.7225, 
    258.1875, 258.263, 259.1595, 259.0065, 257.4693, 254.0737, 252.5938, 
    250.7098,
  274.4087, 272.7931, 270.7038, 262.239, 254.8331, 251.3761, 250.83, 
    253.1998, 252.335, 251.7654, 256.6029, 255.243, 253.5665, 252.1842, 
    251.9873,
  260.9606, 262.8603, 258.3127, 261.6676, 260.7036, 259.9873, 261.2365, 
    258.9669, 257.36, 255.2707, 255.8925, 258.5995, 258.1948, 257.9652, 
    256.757,
  264.6526, 260.6516, 260.0658, 259.1856, 259.3103, 260.9724, 261.3217, 
    258.7744, 256.3209, 257.9471, 257.7755, 260.0176, 260.4053, 256.2386, 
    255.4127,
  272.3986, 269.658, 263.5257, 258.1619, 259.087, 254.0184, 260.8974, 
    259.729, 258.052, 258.4626, 260.1295, 259.1953, 257.9809, 258.2353, 
    256.4302,
  273.4419, 273.1059, 272.6872, 269.0225, 260.6221, 258.9212, 255.6619, 
    259.0991, 259.149, 258.627, 258.8623, 258.8174, 257.1274, 256.8612, 
    257.5804,
  274.2583, 272.9374, 272.5954, 272.1971, 270.053, 263.7521, 261.378, 
    252.5448, 254.0732, 257.8159, 258.8599, 258.3541, 257.197, 256.9545, 
    257.3455,
  274.8955, 273.6689, 272.9213, 272.1703, 272.1243, 271.3398, 267.7314, 
    263.1039, 260.5124, 260.1078, 260.486, 259.4975, 257.8861, 256.3441, 
    255.7797,
  275.4387, 274.586, 273.3499, 272.3192, 272.2856, 271.944, 271.0313, 
    268.408, 262.9805, 261.9948, 260.7957, 259.0431, 257.1534, 256.3462, 
    256.4766,
  275.9161, 274.84, 273.504, 272.3657, 271.9363, 271.21, 269.6521, 267.5331, 
    262.0314, 259.8676, 258.1794, 259.0099, 257.7666, 256.2876, 256.603,
  275.8079, 274.8988, 274.1242, 271.8025, 264.4283, 262.6924, 262.5566, 
    261.9547, 260.2159, 259.2316, 257.8687, 258.8469, 257.8843, 256.7358, 
    255.6939,
  274.3128, 272.4663, 270.0839, 260.8147, 253.5571, 251.5975, 253.5323, 
    258.6498, 257.4313, 256.3954, 258.2589, 259.132, 258.1289, 257.4677, 
    255.5081,
  261.2717, 264.5676, 260.6876, 263.2983, 261.8976, 260.7939, 261.8486, 
    260.5477, 260.0972, 255.8938, 255.7107, 257.2783, 254.4798, 253.1226, 
    251.6639,
  265.7742, 263.8473, 263.278, 262.4718, 260.2881, 260.3821, 261.6, 259.564, 
    257.4244, 258.5975, 256.6797, 259.2792, 259.5356, 252.0677, 251.0388,
  272.5482, 269.6129, 265.8564, 262.913, 259.6905, 254.0734, 259.6464, 
    258.2969, 256.9793, 257.9147, 259.2509, 257.6773, 257.57, 258.4203, 
    254.245,
  273.5387, 273.2374, 272.7584, 269.6805, 261.6739, 258.382, 249.8297, 
    255.6758, 256.8596, 256.8397, 256.7679, 256.9963, 256.5424, 257.267, 
    257.715,
  274.1925, 272.911, 272.5804, 272.1921, 269.5605, 262.3202, 259.7466, 
    250.2382, 251.6672, 254.6542, 255.8534, 256.7717, 256.6819, 257.3284, 
    257.799,
  274.889, 273.6796, 272.873, 272.1162, 272.0984, 271.0356, 265.657, 
    261.7879, 259.9172, 260.7445, 259.1383, 258.0194, 257.2548, 255.7809, 
    254.5856,
  275.4377, 274.5333, 273.3108, 272.2846, 272.2694, 271.901, 270.8713, 
    266.8925, 262.7972, 263.0443, 260.9611, 258.4757, 256.9581, 254.8793, 
    251.9201,
  275.8897, 274.824, 273.4521, 272.3115, 271.9436, 271.1049, 269.8938, 
    267.1785, 261.3029, 259.9351, 258.1941, 257.3925, 255.4134, 251.7253, 
    249.5168,
  275.7778, 274.8695, 274.0464, 270.7808, 265.4904, 265.4991, 264.756, 
    262.5588, 260.1392, 258.0334, 256.2738, 255.2406, 252.5972, 250.9111, 
    250.2373,
  273.88, 271.6243, 268.8763, 260.8651, 258.1988, 259.6879, 260.439, 
    261.2766, 257.7355, 255.9399, 254.9156, 253.7023, 252.683, 251.2689, 
    251.8006,
  262.5247, 265.3215, 264.0033, 263.6715, 261.1655, 262.3289, 261.5924, 
    258.8268, 258.0913, 255.6035, 257.1654, 257.8587, 255.9759, 253.9682, 
    251.5872,
  267.9325, 265.1882, 262.283, 258.512, 255.204, 260.4875, 261.8193, 
    259.2246, 257.3886, 258.3657, 257.3211, 259.3318, 259.3208, 252.621, 
    250.6082,
  272.6463, 269.7642, 264.2969, 258.0283, 255.9374, 256.6867, 260.8687, 
    258.7915, 258.0287, 258.3514, 258.318, 258.0706, 257.5064, 256.8036, 
    252.7099,
  273.6204, 273.316, 272.8128, 268.3945, 260.1014, 260.2931, 255.1379, 
    257.1521, 257.6877, 256.8416, 256.6536, 256.4699, 255.9438, 258.0504, 
    257.324,
  274.1849, 272.9116, 272.553, 272.1347, 267.8576, 262.1682, 261.7852, 
    252.0535, 252.7283, 252.8775, 255.1835, 255.6422, 255.978, 257.1462, 
    258.4099,
  274.8694, 273.6807, 272.8124, 272.072, 272.0358, 269.9138, 262.9032, 
    260.7653, 259.2113, 259.101, 256.2122, 256.3201, 256.4484, 256.4096, 
    256.2154,
  275.3845, 274.4982, 273.2769, 272.2395, 272.2294, 271.7175, 270.1694, 
    264.5754, 260.8708, 261.9622, 259.7814, 256.2812, 255.6936, 254.463, 
    253.5089,
  275.8536, 274.7817, 273.4017, 272.1639, 272.0915, 270.8967, 269.6075, 
    266.0023, 258.5046, 256.8418, 256.0322, 254.9635, 252.9176, 252.2755, 
    250.8825,
  275.7164, 274.8325, 273.9695, 270.1853, 266.1866, 265.6422, 264.1836, 
    260.7319, 256.8492, 253.3286, 251.732, 253.5362, 252.4417, 250.5995, 
    249.5925,
  272.9717, 270.6259, 268.4306, 262.2444, 258.8739, 257.6407, 257.7254, 
    259.5548, 254.9359, 251.2984, 249.935, 251.6096, 250.7295, 248.5688, 
    249.015,
  259.0594, 260.4117, 256.5064, 259.3853, 255.6192, 255.2365, 257.9043, 
    257.3987, 256.7132, 249.1468, 249.985, 258.6036, 257.0949, 255.3027, 
    258.5386,
  265.8105, 260.4805, 258.4048, 257.0361, 255.6887, 257.7407, 259.4408, 
    257.2072, 252.19, 258.4021, 254.4046, 261.0996, 260.9005, 255.0895, 
    255.2845,
  272.4719, 268.3197, 262.7958, 259.9695, 260.6637, 255.7227, 257.11, 
    255.4373, 254.5572, 256.2429, 258.8556, 259.094, 259.6381, 258.973, 
    256.574,
  273.678, 273.329, 272.6145, 267.1205, 261.2271, 260.644, 251.2829, 
    251.5423, 253.8609, 254.4169, 255.328, 256.6206, 257.6886, 258.6017, 
    258.343,
  274.1769, 272.8907, 272.5331, 271.8012, 265.3416, 262.2036, 261.7845, 
    245.2659, 250.6481, 253.75, 255.0135, 255.5452, 256.0429, 258.6951, 
    258.7129,
  274.847, 273.6166, 272.7477, 272.0458, 271.7437, 268.1479, 262.1685, 
    261.3177, 257.2503, 259.4851, 256.3829, 256.3642, 257.2078, 257.1763, 
    255.9777,
  275.3337, 274.4773, 273.251, 272.1839, 272.187, 271.4533, 269.4818, 
    262.5121, 260.2741, 260.1836, 257.0792, 255.895, 256.1493, 255.8867, 
    254.5617,
  275.8365, 274.7977, 273.3876, 272.1609, 272.2885, 271.0657, 269.7089, 
    265.1411, 257.8497, 255.8587, 254.188, 254.4342, 253.1372, 252.8829, 
    251.042,
  275.7376, 274.8404, 274.0199, 270.6672, 266.7466, 265.8002, 264.3968, 
    258.6823, 254.2146, 250.8972, 249.2766, 250.0955, 249.9244, 249.9766, 
    250.39,
  273.1393, 271.4408, 269.3667, 261.9268, 258.8546, 255.3834, 255.6484, 
    256.2596, 251.246, 247.2048, 247.6308, 249.9058, 250.3784, 249.8964, 
    251.3905,
  258.9599, 260.0194, 256.5262, 256.9224, 253.9537, 253.6313, 256.356, 
    256.8848, 257.4827, 256.0832, 256.148, 260.0696, 259.2657, 258.1195, 
    256.4995,
  264.9008, 261.3712, 258.7211, 256.75, 254.0102, 252.5405, 254.9353, 
    254.8919, 255.3674, 258.742, 256.8945, 260.5026, 260.9635, 256.7428, 
    255.0182,
  272.05, 267.0549, 261.3986, 257.7141, 257.156, 247.5238, 254.4672, 
    255.5285, 255.8209, 255.0048, 257.6074, 257.9246, 259.3516, 259.4714, 
    257.6481,
  273.642, 273.286, 272.1061, 265.8249, 259.8408, 258.3354, 247.1387, 
    248.1539, 251.1411, 252.5932, 253.7141, 256.8236, 256.3668, 257.6071, 
    258.7881,
  274.2054, 272.8127, 272.4681, 271.2745, 263.9833, 262.1783, 262.4992, 
    249.6394, 250.7398, 250.6826, 252.4495, 253.1317, 255.0602, 256.5207, 
    258.2218,
  274.9118, 273.6019, 272.7146, 271.9808, 271.4387, 267.4413, 260.7271, 
    262.0122, 256.6493, 257.5114, 251.5296, 254.9934, 254.683, 256.3849, 
    256.2454,
  275.4428, 274.5507, 273.3087, 272.1409, 272.1616, 271.3582, 268.914, 
    261.1883, 257.4868, 255.5284, 252.6996, 254.758, 255.3109, 256.8565, 
    255.893,
  275.8838, 274.9374, 273.4919, 272.1892, 272.3526, 271.3571, 269.5038, 
    263.1196, 253.7773, 251.5656, 250.5007, 253.8295, 256.6502, 256.7982, 
    254.4882,
  275.8409, 274.9171, 274.0556, 270.9475, 267.0159, 264.7074, 263.0365, 
    256.8624, 252.2203, 250.3148, 248.7681, 249.6612, 253.8672, 254.7075, 
    254.2638,
  273.6508, 271.8488, 269.6584, 260.2981, 257.9695, 252.3379, 251.9772, 
    252.8453, 250.8786, 248.6201, 245.886, 248.3718, 248.5586, 252.0001, 
    252.7183,
  257.1446, 259.8371, 256.472, 258.1072, 256.7612, 255.3257, 255.8961, 
    255.3389, 257.2112, 257.0406, 257.7213, 258.4482, 255.4362, 253.9836, 
    255.2035,
  262.6311, 259.3404, 258.0506, 256.59, 255.8876, 252.231, 255.9941, 
    255.0231, 256.2417, 258.4708, 258.4205, 260.4415, 258.996, 252.8269, 
    252.5828,
  271.9044, 266.2172, 260.8501, 256.4602, 255.3535, 250.1969, 255.7203, 
    255.0676, 255.6481, 257.5635, 259.2833, 260.4654, 259.0002, 257.7046, 
    254.9254,
  273.5775, 273.2525, 272.1338, 265.6521, 258.9377, 259.4004, 253.2591, 
    252.1529, 254.9308, 256.4738, 258.3133, 259.1388, 258.0907, 256.905, 
    257.2379,
  274.2552, 272.7465, 272.4361, 271.1952, 262.9105, 261.9305, 260.9454, 
    250.2016, 251.4174, 255.7072, 256.7426, 256.7979, 256.755, 256.5886, 
    257.7593,
  275.0107, 273.6719, 272.7164, 271.9538, 271.4179, 267.495, 260.3697, 
    259.3002, 256.954, 257.1604, 255.5405, 255.8947, 255.19, 254.8338, 
    255.6999,
  275.6084, 274.6599, 273.3994, 272.0979, 272.1537, 271.4995, 268.7219, 
    260.5423, 256.8301, 255.1909, 255.3875, 255.2905, 254.2491, 254.1177, 
    253.7637,
  275.9572, 275.0901, 273.6525, 272.1901, 272.404, 271.4424, 269.0344, 
    262.2911, 254.5494, 254.0838, 253.8384, 254.7876, 254.1602, 253.5144, 
    252.8084,
  275.9471, 275.0639, 274.0921, 271.2745, 267.3645, 264.0931, 261.2242, 
    255.3647, 252.6819, 252.4753, 251.4452, 251.6873, 253.7288, 252.5448, 
    253.6608,
  274.2874, 272.6759, 270.9753, 263.2744, 259.2817, 256.0779, 254.7262, 
    253.5685, 249.8499, 250.1688, 246.6412, 248.9318, 248.9178, 250.7645, 
    252.7841,
  256.4814, 259.0824, 258.8637, 259.3612, 258.7901, 257.1351, 257.6859, 
    256.9637, 257.5657, 254.8968, 251.9905, 252.1908, 251.8174, 253.3633, 
    254.6246,
  262.6754, 259.5424, 258.9857, 258.2303, 258.0347, 255.9005, 258.4064, 
    257.5533, 257.0442, 257.7173, 254.8237, 255.8172, 257.079, 253.6592, 
    253.7438,
  272.1181, 266.4084, 262.6973, 260.0224, 260.4764, 256.9932, 259.537, 
    257.6502, 256.931, 257.7569, 256.9421, 255.7321, 256.2546, 258.6968, 
    257.5111,
  273.5425, 273.2211, 272.3739, 267.8637, 263.79, 263.2154, 253.5292, 
    255.966, 257.2495, 257.2685, 257.5031, 256.1235, 255.321, 256.8092, 
    259.2628,
  274.2444, 272.6998, 272.4279, 271.693, 265.7359, 262.1342, 260.6368, 
    249.4179, 250.5785, 256.0619, 256.0281, 254.8234, 254.7785, 256.6601, 
    259.1776,
  274.9966, 273.7105, 272.6857, 271.954, 271.5196, 266.9668, 260.524, 
    259.6876, 257.4058, 257.6918, 254.9334, 254.1119, 254.4414, 257.824, 
    257.983,
  275.6129, 274.6842, 273.4223, 272.0561, 272.1027, 271.4176, 268.1345, 
    260.813, 257.9145, 256.2324, 254.8945, 253.776, 254.6176, 257.274, 
    257.3297,
  275.9547, 275.1259, 273.7426, 272.2003, 272.3894, 271.1861, 268.015, 
    260.0216, 256.0698, 254.5016, 253.1042, 252.701, 256.0143, 256.6788, 
    255.0426,
  275.9288, 275.1532, 274.104, 270.8204, 265.0641, 262.6425, 259.7726, 
    255.8024, 254.3739, 252.8994, 252.371, 253.3189, 254.8789, 255.2393, 
    254.2823,
  274.2549, 272.6413, 270.5107, 259.5549, 256.2605, 254.2355, 253.5109, 
    254.2597, 251.6226, 249.9514, 249.2967, 251.5032, 252.3875, 251.7078, 
    251.8233,
  259.8631, 259.602, 258.4859, 256.981, 255.1913, 254.8802, 256.0842, 
    254.4879, 254.2674, 252.8407, 253.3438, 254.9569, 254.5797, 254.4415, 
    252.0469,
  263.8566, 260.6142, 259.3263, 257.3401, 255.6616, 256.2578, 257.2292, 
    255.8933, 255.5175, 257.1531, 256.5771, 257.6141, 259.4334, 253.0672, 
    249.8941,
  272.3206, 266.0375, 262.1095, 258.7659, 257.8625, 253.4015, 257.288, 
    257.3012, 256.8036, 259.0737, 257.9599, 255.8654, 258.6742, 259.5486, 
    253.9097,
  273.4812, 273.1827, 272.3833, 267.7995, 260.8354, 260.1324, 252.3211, 
    255.2179, 257.2099, 256.7222, 254.533, 252.8897, 257.0544, 256.7781, 
    255.0688,
  274.2465, 272.6699, 272.4097, 271.7752, 264.0296, 261.1687, 262.4978, 
    251.405, 251.5724, 249.5391, 249.1008, 253.4269, 256.0222, 256.0371, 
    255.8701,
  274.993, 273.6976, 272.5882, 271.8618, 271.0445, 266.5657, 261.524, 
    260.7713, 256.5405, 255.3032, 250.9687, 255.3428, 255.2436, 254.7302, 
    253.5748,
  275.5454, 274.6288, 273.3394, 271.9743, 272.043, 271.2237, 266.5217, 
    259.2718, 256.3603, 255.3078, 255.3063, 254.1115, 253.2457, 251.0795, 
    249.7432,
  275.8632, 274.9762, 273.5842, 272.2313, 272.255, 270.872, 267.7474, 
    259.6271, 255.1342, 253.8901, 253.3951, 252.6469, 251.0128, 249.2363, 
    247.0558,
  275.7563, 274.9614, 273.9787, 270.161, 266.1605, 263.9921, 260.8808, 
    256.7937, 253.7067, 252.7358, 252.3033, 252.1562, 251.0187, 250.0936, 
    249.964,
  273.9895, 272.5174, 268.8995, 258.4139, 257.166, 255.2672, 254.8063, 
    256.4702, 253.2797, 251.9247, 251.1666, 251.9891, 252.3035, 250.0768, 
    251.2854,
  260.5865, 261.4242, 259.8529, 259.0652, 255.7873, 254.3885, 255.6098, 
    252.9617, 251.0067, 244.9999, 245.461, 247.6796, 245.1874, 245.865, 
    245.3301,
  263.9491, 262.6833, 261.0201, 259.0295, 256.2479, 256.4225, 256.0026, 
    253.5887, 251.9271, 251.2301, 249.7422, 252.8901, 253.4716, 248.3926, 
    248.1439,
  272.2503, 266.8392, 262.1855, 259.8428, 258.2526, 253.2572, 255.3209, 
    253.6996, 251.8295, 252.8725, 253.6181, 254.3464, 256.2003, 257.9372, 
    256.4128,
  273.3944, 273.1481, 271.8246, 266.1934, 259.6409, 259.5916, 251.039, 
    250.9521, 250.7959, 250.7762, 253.1276, 254.5056, 256.8004, 257.717, 
    257.6982,
  274.2358, 272.6151, 272.3757, 271.5047, 261.8523, 259.7968, 260.5553, 
    246.8982, 244.5823, 246.5923, 247.9577, 252.0274, 254.9527, 255.4305, 
    255.6064,
  274.9578, 273.5982, 272.5143, 271.704, 269.4482, 264.4995, 259.2184, 
    260.4949, 254.5621, 255.5688, 248.7714, 251.8553, 252.5246, 251.9902, 
    252.8714,
  275.4601, 274.5579, 273.2831, 271.9399, 272.0033, 270.9772, 264.5993, 
    258.6888, 254.0675, 252.968, 251.8916, 251.0802, 250.2119, 248.8351, 
    249.5666,
  275.8039, 274.8903, 273.5141, 272.2777, 272.2301, 270.8215, 267.5418, 
    257.9006, 252.8826, 250.1703, 248.5898, 248.5047, 247.5258, 246.0618, 
    247.0848,
  275.6418, 274.8291, 273.9008, 271.2233, 268.3838, 265.7605, 260.8128, 
    254.1147, 250.5007, 247.278, 246.4794, 246.5153, 245.8995, 245.7696, 
    245.6443,
  274.1826, 272.9869, 268.9546, 259.1511, 256.8239, 255.0137, 252.9646, 
    253.8003, 248.813, 243.114, 242.3684, 245.9263, 245.792, 245.4556, 
    246.0951,
  259.1696, 261.4662, 261.0815, 260.4169, 256.8549, 255.6836, 256.9158, 
    254.0131, 250.6825, 244.6628, 243.9519, 245.1392, 241.6819, 242.8457, 
    241.4035,
  261.3535, 261.1794, 261.1136, 259.4754, 255.4894, 255.8396, 256.2176, 
    253.1357, 249.1865, 248.5485, 245.8464, 250.5472, 250.8295, 245.1293, 
    245.4049,
  272.0183, 265.3487, 261.3056, 259.0875, 258.1468, 252.0065, 254.501, 
    251.8907, 248.4331, 249.2781, 250.5135, 251.3488, 253.3715, 255.2322, 
    253.9019,
  273.3377, 273.0671, 271.0493, 264.3133, 259.8882, 259.478, 247.7511, 
    248.4393, 247.2389, 246.8423, 249.7892, 251.864, 254.2399, 256.3497, 
    255.948,
  274.2337, 272.5775, 272.3442, 271.0133, 260.7134, 259.6979, 260.4322, 
    245.0948, 240.3021, 245.533, 246.5, 249.6616, 253.8384, 254.113, 254.8605,
  274.9122, 273.4661, 272.4675, 271.3942, 267.8546, 262.6721, 258.631, 
    259.9866, 252.6227, 250.7954, 245.7722, 249.6659, 251.32, 251.0645, 
    251.3873,
  275.3685, 274.4726, 273.2278, 271.8915, 271.9428, 270.5418, 263.0861, 
    256.1115, 251.3916, 249.6348, 249.3356, 249.0358, 248.8915, 247.2036, 
    249.0522,
  275.7612, 274.8595, 273.5012, 272.2733, 272.2286, 270.8979, 267.3734, 
    258.8097, 251.1186, 248.7982, 248.3058, 247.8905, 247.6025, 246.6543, 
    248.1839,
  275.6089, 274.7833, 273.8626, 271.7433, 269.8098, 266.9825, 262.041, 
    253.3018, 249.3477, 246.6534, 245.8897, 246.667, 246.5597, 247.4449, 
    247.5611,
  274.2987, 273.1945, 269.0548, 259.9994, 257.5954, 254.8839, 254.85, 
    251.7941, 247.7038, 241.8185, 240.4769, 244.8396, 245.0281, 244.8661, 
    245.8154,
  259.6088, 260.9905, 259.6631, 257.8233, 255.611, 252.1186, 257.6465, 
    257.0772, 255.9929, 251.918, 250.8458, 250.7971, 246.7553, 245.083, 
    241.0278,
  262.6853, 258.0966, 258.6836, 257.1794, 250.9131, 253.916, 256.8338, 
    255.7285, 254.4804, 254.1733, 251.0314, 251.5514, 250.1384, 240.8517, 
    241.1037,
  271.6891, 264.9216, 259.5443, 256.8665, 256.338, 249.7398, 253.5977, 
    253.4476, 252.7958, 252.8168, 251.4341, 249.6924, 249.8046, 250.6667, 
    250.1256,
  273.2829, 273.0212, 270.635, 262.7473, 258.1106, 259.2571, 246.6338, 
    249.453, 249.2251, 246.7339, 248.4753, 249.1982, 251.0084, 252.8573, 
    253.9211,
  274.2401, 272.5414, 272.2993, 270.0197, 257.627, 259.2943, 259.9664, 
    243.0191, 237.6842, 242.4251, 246.5981, 248.7687, 251.1508, 252.266, 
    254.6588,
  274.936, 273.362, 272.4206, 270.8512, 266.031, 259.8691, 258.0673, 259.646, 
    251.7865, 249.5233, 245.7467, 247.5714, 249.7271, 250.5896, 253.2414,
  275.3643, 274.4428, 273.2061, 271.8224, 271.86, 269.8387, 261.5082, 
    255.4035, 251.1901, 249.6301, 247.9676, 247.225, 247.0747, 248.2503, 
    250.5793,
  275.7715, 274.8869, 273.5242, 272.2494, 272.2341, 270.8599, 266.8486, 
    255.7146, 250.4577, 248.4094, 247.1726, 246.8611, 246.3801, 247.2377, 
    248.9243,
  275.6484, 274.8181, 273.8485, 271.9599, 269.7841, 266.5344, 260.8394, 
    252.7945, 249.9576, 247.611, 247.0508, 247.2189, 247.5155, 247.9093, 
    248.7333,
  274.3793, 273.2914, 269.4502, 262.4212, 258.1624, 255.9212, 255.4554, 
    251.3522, 248.2344, 243.4877, 244.3643, 247.0987, 247.5022, 246.981, 
    248.0615,
  260.4787, 261.7389, 259.4434, 255.556, 251.5312, 250.2576, 254.183, 
    254.7769, 255.8515, 250.6791, 249.0646, 250.8064, 249.675, 245.858, 
    242.1237,
  262.486, 258.3177, 256.7177, 253.7328, 249.0538, 249.3065, 252.0676, 
    252.6048, 253.6681, 254.9178, 250.4764, 251.3992, 251.1046, 239.66, 
    236.286,
  271.0037, 263.5158, 257.1821, 254.2061, 253.5033, 243.0643, 248.4238, 
    250.2092, 251.239, 253.3275, 253.1838, 251.8484, 251.6767, 250.3146, 
    246.6385,
  273.2122, 272.8782, 270.0196, 261.8691, 255.3249, 257.3934, 240.6842, 
    247.0974, 249.6743, 250.1421, 252.5315, 252.719, 253.3748, 252.7577, 
    249.8791,
  274.2428, 272.5255, 272.2618, 268.878, 254.8212, 257.7577, 259.744, 
    240.067, 240.9039, 247.1503, 249.7, 250.9679, 252.0523, 251.7513, 251.2891,
  274.9935, 273.327, 272.3704, 270.3055, 264.8222, 258.3596, 257.4606, 
    258.9108, 252.3751, 251.1552, 248.2931, 249.9489, 250.7002, 250.2424, 
    250.4941,
  275.4125, 274.4478, 273.1986, 271.7609, 271.7667, 269.2777, 258.9603, 
    253.5866, 251.3524, 249.7925, 248.8026, 248.6323, 248.8477, 247.8548, 
    249.0576,
  275.7748, 274.9108, 273.5736, 272.2078, 272.2317, 270.7525, 265.3923, 
    253.8451, 250.2482, 248.3009, 247.8321, 247.5563, 247.5401, 248.0578, 
    249.2243,
  275.6651, 274.8554, 273.8367, 271.9459, 269.6838, 265.1043, 256.8426, 
    251.9609, 249.3303, 247.2109, 246.8884, 247.0326, 247.3419, 247.7156, 
    249.2783,
  274.4764, 273.4926, 269.2017, 260.4489, 255.0113, 252.9314, 251.9942, 
    251.6419, 248.0887, 244.5391, 244.1308, 246.8575, 246.5381, 246.1583, 
    247.4584,
  259.43, 259.0674, 255.6512, 254.7086, 250.8981, 248.1916, 250.6408, 
    250.0411, 251.0863, 244.8849, 243.8487, 246.4203, 244.926, 242.3899, 
    239.8359,
  259.941, 257.1175, 255.6418, 252.4523, 247.2508, 244.4439, 247.5073, 
    247.9252, 248.6007, 250.8872, 245.5333, 249.0529, 249.4653, 237.7634, 
    235.1716,
  269.3198, 261.1945, 255.8955, 253.5664, 251.7647, 239.8668, 244.437, 
    246.3327, 246.4212, 248.7357, 249.5554, 249.4342, 249.7957, 248.466, 
    241.947,
  273.0931, 272.5113, 269.6005, 262.3768, 256.8117, 256.6157, 238.9997, 
    244.118, 247.1406, 245.9697, 247.9007, 248.8513, 249.6482, 248.8516, 
    245.5701,
  274.1941, 272.5106, 272.258, 269.0538, 255.0724, 259.498, 259.0038, 
    238.4008, 240.2622, 244.9521, 246.4517, 247.4182, 249.461, 249.4277, 
    249.9759,
  275.006, 273.3341, 272.2811, 270.0905, 264.8024, 258.3817, 257.4925, 
    258.2664, 252.1586, 250.8656, 246.1339, 247.1986, 248.5393, 249.2088, 
    249.9837,
  275.4402, 274.4828, 273.2253, 271.7039, 271.7394, 268.6773, 258.3528, 
    254.228, 252.2166, 250.4369, 248.5505, 246.9264, 246.1739, 245.8215, 
    247.4581,
  275.7629, 274.9315, 273.6607, 272.1855, 272.2288, 270.7128, 264.3574, 
    253.9148, 251.1255, 249.2879, 247.7287, 246.4572, 244.907, 244.6938, 
    246.2852,
  275.6541, 274.8816, 273.8463, 271.9684, 269.5645, 265.0477, 256.7905, 
    252.7229, 250.2499, 246.772, 245.7189, 245.0279, 244.2809, 244.149, 
    244.7063,
  274.5017, 273.5526, 269.2547, 259.1728, 254.0471, 252.7112, 252.6865, 
    252.2477, 247.5596, 242.2125, 240.5472, 243.9599, 242.8866, 242.5169, 
    243.7603,
  258.1907, 258.8572, 256.3211, 256.3411, 254.7811, 252.9251, 253.1042, 
    252.4525, 252.678, 246.7261, 244.6268, 244.9948, 241.3746, 239.8895, 
    235.9352,
  258.5123, 257.1925, 256.2868, 254.3613, 252.0598, 247.2206, 249.7383, 
    249.7144, 249.5625, 250.1578, 243.9541, 247.0221, 247.6603, 237.2442, 
    235.5956,
  267.7568, 258.9985, 256.3255, 254.6778, 253.7638, 242.1491, 245.4062, 
    247.1383, 246.6226, 247.7644, 247.7554, 247.6464, 248.5591, 248.3302, 
    241.9048,
  272.9007, 272.2509, 268.5122, 259.7621, 256.1412, 256.1417, 239.727, 
    243.6596, 245.2052, 244.0032, 245.6695, 247.1856, 248.6483, 248.9703, 
    245.6466,
  274.1699, 272.4995, 272.2889, 268.5241, 254.555, 258.3133, 258.0126, 
    239.1371, 237.1562, 241.128, 243.9848, 246.1634, 248.4506, 248.9447, 
    249.0916,
  275.0352, 273.3286, 272.1402, 269.5504, 264.0786, 256.6103, 258.4141, 
    258.1757, 250.0672, 246.4512, 242.1488, 245.1972, 247.0725, 247.761, 
    247.9451,
  275.4847, 274.5575, 273.2603, 271.6219, 271.6607, 267.8269, 258.3606, 
    253.6946, 249.3132, 246.9578, 244.9672, 244.3293, 244.1843, 244.4803, 
    245.1619,
  275.7812, 274.9828, 273.7733, 272.2065, 272.2206, 270.5521, 263.4162, 
    252.7909, 248.5755, 245.2345, 243.6667, 242.9806, 241.9991, 242.8808, 
    245.1833,
  275.6859, 274.9523, 273.8826, 271.894, 269.4733, 265.0724, 257.09, 
    251.2084, 247.34, 243.5492, 242.6883, 242.4181, 242.4361, 243.8966, 
    245.6364,
  274.5453, 273.5621, 269.5274, 260.6513, 257.1375, 255.075, 252.8393, 
    250.2941, 245.4331, 239.503, 239.3989, 243.4092, 243.8689, 245.283, 
    247.1755,
  258.8004, 259.1078, 256.8472, 257.411, 258.3888, 256.613, 256.8646, 
    257.1333, 258.7336, 255.4659, 253.773, 254.0701, 251.723, 250.4962, 
    246.875,
  259.409, 258.6281, 257.847, 258.2368, 257.3169, 253.2266, 254.5882, 
    254.9165, 255.9276, 256.4686, 252.4887, 253.248, 252.9126, 245.2023, 
    242.5052,
  266.8798, 260.2284, 258.7259, 258.8072, 258.4747, 248.5589, 250.6363, 
    251.8451, 252.2074, 253.1056, 252.2798, 251.3003, 251.4602, 250.6313, 
    245.1383,
  272.7533, 272.4661, 267.744, 260.0857, 258.1843, 258.3276, 245.1137, 
    247.8513, 248.0655, 247.4878, 248.5539, 248.9895, 249.8479, 249.5839, 
    246.6244,
  274.1421, 272.4673, 272.3308, 266.7253, 255.8648, 256.8748, 258.3817, 
    239.6915, 236.8975, 242.1297, 244.9446, 247.5254, 248.2108, 248.2407, 
    248.6624,
  275.0616, 273.3067, 271.9774, 268.5518, 262.6186, 255.8023, 258.0801, 
    257.9146, 249.2823, 245.4091, 241.6819, 244.4211, 245.4341, 246.347, 
    246.6989,
  275.518, 274.5852, 273.2843, 271.5101, 271.4725, 267.1614, 257.7515, 
    252.0389, 247.3236, 245.9536, 244.5235, 243.2775, 243.2804, 243.9831, 
    244.1166,
  275.7961, 274.9697, 273.8119, 272.2352, 272.1394, 270.4814, 261.7361, 
    251.0146, 247.6323, 246.057, 244.7638, 244.1455, 243.0312, 242.8265, 
    244.4766,
  275.7237, 275.0088, 273.9028, 271.8769, 269.4856, 264.8893, 256.1817, 
    251.5233, 249.5602, 248.8624, 248.4287, 248.2074, 247.3742, 247.7602, 
    247.0798,
  274.6536, 273.6475, 270.3719, 263.0328, 257.5746, 254.9988, 253.5034, 
    252.9224, 251.9377, 249.9093, 251.0732, 251.8335, 250.3188, 250.0193, 
    249.4837,
  259.6781, 260.6625, 258.83, 258.9066, 260.173, 258.3745, 260.6538, 
    261.8452, 263.7401, 260.904, 260.9009, 262.8369, 261.6283, 260.2476, 
    257.3708,
  259.592, 260.7215, 260.1227, 261.8474, 260.0248, 255.4794, 256.7141, 
    259.6638, 261.6363, 262.9886, 260.1108, 262.096, 262.3113, 256.9912, 
    254.4223,
  266.4127, 262.7101, 261.3254, 262.7239, 261.6755, 252.9832, 254.2203, 
    255.1156, 257.5823, 259.7875, 260.1452, 260.1577, 260.3246, 260.0181, 
    255.7889,
  272.8208, 272.808, 268.7046, 262.2997, 261.9383, 261.7914, 250.0261, 
    252.033, 251.9096, 254.1541, 256.2878, 256.6939, 257.1088, 256.3901, 
    254.6369,
  274.121, 272.4713, 272.4021, 266.6713, 259.8199, 260.5043, 261.3893, 
    243.9802, 241.0144, 247.6457, 251.1571, 252.9212, 254.4314, 254.2656, 
    253.6877,
  275.1059, 273.3383, 271.9311, 268.6966, 262.6949, 258.39, 259.0488, 
    258.6301, 249.6194, 246.5628, 244.8225, 247.601, 250.5598, 251.2695, 
    251.3522,
  275.5497, 274.614, 273.3408, 271.5339, 271.5219, 267.657, 258.0262, 
    253.2361, 248.8948, 247.2242, 244.8407, 244.7483, 245.9493, 247.3173, 
    248.0689,
  275.7971, 274.9461, 273.8324, 272.2658, 272.0612, 270.8011, 263.165, 
    254.8827, 255.1941, 251.0238, 247.2492, 245.2798, 243.7906, 243.448, 
    247.6083,
  275.7317, 274.9977, 273.8853, 271.5831, 269.1044, 264.7765, 258.6472, 
    255.9743, 254.3759, 253.6851, 252.3282, 249.8186, 247.0997, 246.2874, 
    246.2421,
  274.7303, 273.7089, 269.5036, 262.622, 259.8992, 258.3505, 256.9821, 
    255.3775, 252.0756, 249.197, 253.3465, 253.8645, 250.7313, 249.3187, 
    248.1377,
  259.5938, 263.5518, 258.9337, 259.3853, 262.0176, 257.8409, 258.6132, 
    260.4178, 262.1269, 258.2808, 257.8349, 263.5099, 260.3489, 261.0625, 
    257.5914,
  261.1052, 262.9237, 260.3318, 261.9106, 261.3174, 255.6868, 256.492, 
    259.1756, 262.9087, 263.5103, 259.7782, 263.8396, 264.1777, 260.4861, 
    257.7878,
  267.3782, 265.3337, 261.7117, 262.8511, 262.4826, 253.5352, 254.7867, 
    255.9019, 257.5066, 260.7038, 262.4824, 262.8291, 263.4555, 263.4121, 
    259.8583,
  273.0147, 273.0616, 270.1289, 262.2192, 263.6103, 262.9471, 249.5713, 
    253.1927, 253.7963, 254.2548, 258.2271, 260.8243, 261.9709, 261.7815, 
    260.4412,
  274.1268, 272.5185, 272.6017, 266.9779, 261.6205, 263.1075, 262.3784, 
    243.3296, 243.8206, 249.031, 251.3436, 255.9242, 258.882, 260.4222, 
    260.6281,
  275.072, 273.422, 271.9735, 268.8012, 265.6946, 264.5045, 262.4502, 
    260.2638, 251.4242, 247.7519, 245.7257, 249.0498, 252.8492, 256.7229, 
    258.7005,
  275.5351, 274.6837, 273.4427, 271.5466, 271.5645, 269.1668, 262.1134, 
    257.4688, 255.6942, 251.4269, 246.4602, 245.4711, 246.9328, 249.5406, 
    254.1833,
  275.8289, 274.9994, 273.874, 272.2881, 271.9821, 270.9241, 263.6721, 
    256.9346, 256.6613, 255.4934, 252.2045, 245.2322, 243.7567, 244.7115, 
    248.5964,
  275.7318, 275.0174, 273.8571, 271.2771, 268.0079, 262.3917, 256.2407, 
    252.72, 251.7468, 250.8457, 248.8431, 249.3437, 246.7396, 244.3615, 
    244.5607,
  274.7761, 273.7292, 270.0489, 262.9868, 257.6908, 253.7775, 252.7635, 
    251.8601, 249.879, 247.709, 249.109, 248.9283, 246.471, 244.0277, 243.7136,
  260.6398, 261.2549, 259.6977, 257.6264, 257.1772, 250.1156, 251.7934, 
    255.6342, 260.2357, 260.028, 257.1023, 260.4227, 259.4512, 255.4312, 
    254.0698,
  262.1429, 261.3932, 260.3196, 261.3967, 259.019, 247.26, 250.3139, 
    251.9923, 257.0998, 259.6954, 260.3753, 264.377, 264.8841, 258.5468, 
    255.7169,
  267.4194, 263.7004, 262.2266, 262.6028, 261.934, 250.7954, 248.5342, 
    249.8963, 251.6787, 253.9176, 256.925, 259.7121, 262.4601, 263.516, 
    261.6289,
  273.008, 272.9493, 270.1448, 263.9321, 263.4439, 262.232, 248.4958, 
    249.1505, 250.3648, 249.8622, 251.6972, 255.4436, 257.7211, 258.5811, 
    258.1513,
  274.1067, 272.5584, 272.7067, 268.096, 262.8687, 263.9033, 262.7494, 
    244.3853, 241.5215, 246.7003, 247.7769, 250.2171, 253.6694, 255.7412, 
    257.377,
  275.0268, 273.4484, 271.9856, 269.5355, 265.5479, 263.2354, 263.7091, 
    262.3289, 253.7701, 248.9159, 244.1622, 246.923, 248.916, 251.5704, 
    254.4405,
  275.5017, 274.681, 273.4585, 271.5561, 271.4033, 268.7962, 262.3599, 
    258.656, 255.7488, 254.362, 247.9169, 245.4005, 245.8439, 247.0103, 
    250.1438,
  275.8221, 274.9937, 273.8809, 272.2979, 271.9348, 271.0087, 263.4387, 
    257.3928, 254.7284, 255.2172, 252.0139, 245.4328, 243.6728, 244.5862, 
    247.2084,
  275.7133, 275.0349, 273.8633, 271.5786, 269.1722, 265.153, 259.4631, 
    255.4399, 254.2249, 252.0711, 250.9737, 246.5248, 243.5224, 243.663, 
    245.3651,
  274.8387, 273.8339, 271.3484, 265.7158, 261.1992, 259.1758, 257.2859, 
    255.999, 252.5266, 251.2, 252.9408, 247.7918, 242.9536, 242.627, 243.8527,
  260.4153, 260.601, 259.5498, 260.2839, 259.2316, 252.535, 251.0961, 
    252.3159, 258.5429, 260.6726, 260.3444, 262.0056, 260.5826, 252.6794, 
    251.8049,
  265.1947, 261.2311, 261.0304, 261.6637, 260.0303, 251.1383, 250.3828, 
    250.1261, 253.2506, 257.8323, 259.9854, 263.5287, 262.9988, 258.9315, 
    254.0759,
  268.1478, 264.4604, 262.1292, 263.4637, 262.509, 253.8992, 249.5099, 
    248.7114, 249.8901, 251.7717, 253.5881, 256.4331, 258.1589, 259.7172, 
    255.7322,
  273.0378, 272.7518, 270.1215, 265.3316, 264.4427, 262.7045, 253.2398, 
    248.4379, 249.2431, 248.7281, 250.7711, 252.0187, 252.7576, 252.9495, 
    251.9332,
  274.1052, 272.6221, 272.7359, 269.2259, 264.6198, 264.2521, 263.4354, 
    255.6407, 253.5568, 246.5816, 247.2484, 249.0677, 250.5176, 250.896, 
    251.547,
  275.0144, 273.4684, 272.1119, 270.2728, 266.5842, 264.3688, 264.0709, 
    263.3047, 256.0044, 251.2623, 245.9175, 246.5076, 247.4837, 248.6922, 
    250.0664,
  275.4741, 274.6529, 273.4396, 271.5092, 271.1707, 268.9217, 263.7617, 
    260.2627, 256.6051, 252.9223, 248.8759, 246.5434, 245.2127, 245.7212, 
    248.7094,
  275.8087, 274.9757, 273.8539, 272.3075, 272.1031, 271.1729, 265.3426, 
    259.4661, 254.8416, 252.5024, 249.3709, 247.882, 243.3445, 244.3581, 
    248.4043,
  275.6962, 275.0258, 273.9124, 271.9695, 270.7615, 267.8021, 263.4123, 
    258.0514, 253.6098, 252.157, 248.7492, 248.4699, 242.5574, 243.9671, 
    247.8237,
  274.8717, 273.8909, 271.99, 268.372, 266.1717, 265.1483, 261.6178, 
    256.2777, 251.9432, 249.8121, 249.6235, 246.6727, 242.1373, 242.9602, 
    246.311,
  266.5439, 264.6774, 261.337, 260.9308, 256.513, 255.1918, 256.9372, 
    258.7992, 261.8239, 260.2247, 259.9045, 260.6326, 259.5923, 256.1285, 
    253.0727,
  266.9889, 265.159, 261.4611, 260.2429, 255.1287, 252.3137, 256.1183, 
    257.8327, 260.0284, 262.0286, 261.2427, 262.7991, 262.4353, 249.8884, 
    251.8482,
  270.0323, 267.4024, 263.9798, 263.037, 259.8144, 250.1751, 253.6763, 
    255.5292, 257.5544, 258.4493, 259.4359, 259.8552, 258.2026, 257.1497, 
    248.0327,
  273.0482, 272.6327, 270.0876, 264.6514, 262.2987, 261.6577, 250.9744, 
    253.4012, 254.3809, 255.2259, 256.186, 254.9761, 254.0509, 252.1127, 
    248.9071,
  274.128, 272.656, 272.7462, 269.0863, 262.0106, 262.8805, 262.1261, 
    249.5895, 249.0818, 250.7515, 252.4255, 252.6962, 252.1749, 250.8078, 
    250.4683,
  275.0578, 273.5025, 272.1226, 269.9714, 264.8948, 262.35, 263.021, 
    262.9366, 258.717, 254.5793, 250.1348, 249.7417, 248.7573, 248.2378, 
    249.0487,
  275.516, 274.6724, 273.427, 271.3319, 270.4788, 268.2745, 262.624, 
    261.2745, 258.175, 254.7393, 251.5823, 248.7775, 246.2613, 245.759, 
    248.3423,
  275.8459, 274.9921, 273.8447, 272.2765, 272.1154, 271.1838, 264.627, 
    259.6599, 256.1375, 253.008, 250.1934, 247.8025, 243.6658, 244.7509, 
    248.5396,
  275.7488, 275.0577, 273.9308, 272.111, 271.3296, 268.3214, 263.2994, 
    259.0208, 254.562, 251.4305, 248.8299, 245.7105, 242.6738, 244.4734, 
    247.7997,
  275.0108, 273.9426, 272.0958, 267.2232, 263.5083, 264.3096, 262.2171, 
    257.2631, 252.3113, 249.3486, 247.3087, 244.7651, 242.198, 243.7429, 
    246.9771,
  267.3691, 266.361, 265.5461, 264.2054, 258.0256, 251.0632, 254.8842, 
    256.9943, 258.8, 255.9777, 256.5318, 256.9198, 255.2807, 253.2158, 
    248.8688,
  267.837, 267.0732, 266.2478, 263.1862, 255.6834, 248.874, 252.0004, 
    255.5001, 258.419, 259.8636, 258.8098, 259.8577, 259.148, 250.9849, 
    249.1748,
  269.6921, 267.663, 266.2772, 263.5048, 259.3261, 247.1438, 250.3279, 
    254.0302, 257.9332, 260.3087, 261.0014, 260.3502, 259.6114, 258.5676, 
    253.2354,
  272.9974, 272.4644, 270.4538, 264.7583, 261.5797, 260.3322, 249.1026, 
    253.2249, 256.6364, 258.8332, 259.2859, 258.679, 257.8383, 256.3087, 
    252.6238,
  274.1426, 272.6883, 272.7962, 268.8646, 258.6025, 261.1599, 262.8043, 
    248.6703, 249.7007, 255.0258, 256.2654, 256.0794, 255.6705, 254.4866, 
    252.8358,
  275.0849, 273.5493, 272.1193, 270.0241, 260.8665, 258.0605, 262.4564, 
    262.839, 259.1288, 257.0618, 254.0331, 253.6838, 253.2978, 252.6119, 
    251.1418,
  275.5274, 274.6919, 273.406, 271.2036, 269.6307, 266.9979, 261.6427, 
    260.0454, 257.2792, 255.9866, 253.7069, 252.2474, 250.7722, 249.6792, 
    249.2866,
  275.8454, 274.9804, 273.7867, 272.2245, 272.0728, 270.8065, 261.5439, 
    257.9783, 255.1763, 253.761, 251.6278, 250.1426, 246.8863, 246.707, 
    248.2023,
  275.7414, 275.0467, 273.91, 272.046, 271.1954, 266.6958, 259.3856, 
    256.5177, 253.0379, 250.596, 248.946, 247.3875, 244.3337, 245.5576, 
    247.0123,
  275.0955, 273.9959, 272.0558, 265.1299, 259.5369, 259.7523, 257.3287, 
    254.6597, 251.1216, 247.9411, 246.2887, 246.0441, 243.1948, 244.2306, 
    246.0378,
  269.5026, 268.8225, 268.4525, 267.941, 266.9363, 264.939, 263.0189, 
    261.3358, 260.1566, 256.2009, 255.1867, 255.674, 254.4336, 254.2958, 
    251.218,
  269.4416, 269.1334, 268.6007, 267.583, 265.3025, 259.6059, 258.5428, 
    257.0888, 257.4237, 256.7875, 255.9731, 258.0602, 258.1295, 252.0875, 
    250.2323,
  270.1181, 268.8595, 267.5454, 266.503, 264.1872, 255.7367, 256.7991, 
    257.4971, 256.025, 256.1873, 257.1875, 258.0943, 258.7675, 259.1112, 
    255.3946,
  273.0111, 272.584, 270.3035, 266.0015, 264.0949, 260.9439, 251.7346, 
    254.1112, 253.1488, 254.0225, 255.9218, 257.536, 258.749, 258.7556, 
    256.1418,
  274.1392, 272.6956, 272.7742, 267.9512, 262.8317, 262.8606, 262.3989, 
    249.0466, 245.021, 252.5457, 255.3719, 257.4911, 258.5023, 258.4144, 
    256.9712,
  275.0396, 273.4754, 272.1024, 269.2672, 264.6027, 260.7212, 261.8297, 
    261.1631, 257.7299, 255.9142, 255.1288, 256.8021, 257.464, 257.2066, 
    256.4873,
  275.443, 274.5836, 273.3282, 270.9185, 269.7782, 266.0115, 259.7465, 
    258.8434, 257.1168, 256.9518, 256.4355, 256.4403, 256.1546, 255.7399, 
    255.3491,
  275.7605, 274.8918, 273.7112, 272.156, 272.0025, 269.6756, 259.3861, 
    256.9862, 255.9384, 255.5662, 255.409, 255.1291, 254.2037, 254.2401, 
    253.8466,
  275.6409, 274.9759, 273.8524, 271.9621, 270.4688, 264.7497, 257.4765, 
    255.5483, 254.1536, 253.6612, 253.3495, 253.11, 251.9488, 251.8578, 
    250.2944,
  274.9916, 273.9548, 271.4405, 261.5417, 256.1399, 257.1428, 255.8391, 
    254.2792, 252.4126, 250.8542, 250.3618, 250.8586, 249.2874, 248.3464, 
    247.9785,
  264.3358, 262.3791, 260.4057, 260.3383, 261.5548, 257.0281, 255.8687, 
    257.3257, 258.4814, 257.8019, 257.7218, 259.1094, 258.9014, 259.6219, 
    258.3502,
  264.0065, 262.346, 260.1769, 260.3132, 259.4236, 255.9386, 254.1843, 
    252.6494, 254.3076, 256.1425, 255.2288, 257.9478, 257.0878, 251.7597, 
    255.0326,
  268.2289, 262.3528, 259.8756, 260.3922, 260.7096, 252.476, 253.5418, 
    253.2438, 253.8622, 255.2157, 256.7593, 257.9617, 258.3131, 258.8868, 
    257.3067,
  272.9469, 272.4271, 268.9489, 262.6563, 262.2708, 260.6881, 249.5482, 
    251.0373, 253.2644, 254.7963, 256.2881, 258.3123, 258.6568, 259.0453, 
    257.8289,
  274.1102, 272.6678, 272.7306, 266.6061, 261.1039, 261.4104, 260.8491, 
    244.3804, 246.0229, 253.487, 256.06, 257.1478, 258.8604, 259.0278, 
    258.1323,
  275.0084, 273.4359, 272.061, 268.5543, 262.7639, 259.9985, 260.3384, 
    259.7118, 256.8571, 256.7462, 255.3529, 256.811, 257.9611, 257.879, 
    256.8889,
  275.4133, 274.54, 273.2697, 270.7678, 269.6962, 264.1729, 258.1872, 
    257.2684, 256.8877, 257.683, 257.3987, 257.2904, 257.2272, 256.9031, 
    256.5619,
  275.739, 274.8636, 273.6464, 272.0772, 271.9624, 268.0775, 256.876, 
    255.5133, 255.1342, 256.0605, 256.721, 256.9626, 256.35, 256.0801, 
    256.0102,
  275.6364, 274.96, 273.8119, 271.6809, 268.8613, 261.0751, 255.5925, 
    254.6906, 254.0922, 253.8924, 254.4501, 254.7406, 254.2417, 254.0659, 
    252.7429,
  275.0131, 273.9332, 271.0094, 260.4691, 253.9536, 253.6024, 254.0386, 
    253.8486, 252.6492, 251.027, 251.1238, 252.3503, 251.9409, 251.5846, 
    250.7054,
  267.1716, 263.2942, 259.3987, 257.3455, 256.7599, 252.7489, 252.6857, 
    252.4543, 254.868, 254.0029, 255.545, 257.0833, 256.6121, 255.2825, 
    254.4698,
  268.1913, 263.5404, 260.9297, 257.3423, 255.8974, 250.3767, 252.6434, 
    251.5736, 253.7766, 256.117, 256.025, 258.8506, 258.9989, 251.741, 
    253.5859,
  270.0583, 264.5409, 262.3533, 258.4672, 258.7979, 248.0598, 251.7263, 
    254.1367, 255.5419, 257.1696, 258.2154, 259.3288, 259.4422, 258.6344, 
    259.8053,
  272.932, 272.6781, 270.1263, 260.7535, 261.7522, 258.0241, 247.101, 
    251.5848, 255.0218, 257.3139, 258.8138, 259.3371, 259.3143, 258.938, 
    258.7901,
  274.1384, 272.6972, 272.7773, 265.9466, 259.0055, 259.056, 258.5872, 
    243.5465, 249.3925, 256.1855, 258.2049, 258.5667, 259.0164, 258.2988, 
    258.5195,
  275.037, 273.4773, 272.0882, 268.7695, 262.4637, 258.4942, 258.4707, 
    256.4102, 255.0306, 257.1088, 256.0365, 257.6021, 258.3383, 257.8684, 
    257.4309,
  275.4385, 274.5774, 273.2784, 271.0444, 270.4068, 263.9914, 256.5424, 
    253.7547, 253.5344, 254.8996, 254.7464, 255.7945, 256.3602, 256.1641, 
    256.1165,
  275.7588, 274.9169, 273.6664, 272.0618, 271.9692, 267.4458, 255.0897, 
    252.6698, 251.6754, 252.1864, 252.6291, 253.2476, 253.1422, 253.5259, 
    253.5817,
  275.6654, 274.9988, 273.8475, 271.8841, 269.5391, 260.3301, 254.4426, 
    251.9079, 250.4831, 249.4986, 249.894, 250.3921, 250.7157, 250.9065, 
    250.6274,
  275.0444, 273.9981, 272.2333, 268.946, 262.4441, 255.0748, 253.1642, 
    252.1897, 249.1738, 245.5689, 246.1705, 248.742, 248.6233, 248.9569, 
    249.7081,
  272.4455, 270.3125, 265.7239, 259.7213, 253.9937, 249.8455, 248.7894, 
    250.1204, 256.0867, 254.8494, 256.2732, 257.5027, 255.0526, 253.2183, 
    248.9969,
  272.3829, 269.9299, 265.1559, 258.0833, 252.4408, 248.6283, 249.6878, 
    250.1663, 254.0297, 255.9905, 255.8476, 259.4399, 258.9755, 250.444, 
    244.9212,
  272.0077, 269.8389, 264.9496, 259.2435, 256.74, 247.0605, 249.059, 
    251.4552, 255.0717, 256.583, 257.1792, 257.4774, 256.7822, 255.8604, 
    252.8981,
  273.008, 272.6795, 269.5547, 261.4797, 260.404, 257.0796, 245.0016, 
    250.7092, 253.6911, 256.1076, 257.3882, 257.006, 256.6591, 256.643, 
    257.4054,
  274.2119, 272.7737, 272.8297, 265.9432, 260.0587, 260.1339, 258.7277, 
    244.6128, 250.1244, 253.5623, 255.9939, 257.0775, 258.2823, 258.5537, 
    259.0059,
  275.0881, 273.5443, 272.0823, 268.4543, 262.3859, 259.1873, 259.5145, 
    256.5919, 252.6753, 255.2285, 253.7388, 255.9878, 257.2658, 257.2346, 
    257.6181,
  275.4813, 274.6636, 273.2794, 270.5536, 269.5861, 262.9922, 257.6154, 
    253.5372, 252.1793, 252.7576, 252.5227, 254.3957, 255.2343, 255.7778, 
    256.4871,
  275.7869, 274.9526, 273.7076, 272.0658, 271.9691, 266.9494, 256.194, 
    253.1174, 250.8574, 250.1529, 250.4453, 251.6504, 252.3253, 253.9848, 
    254.4858,
  275.6729, 275.0151, 273.9025, 272.2638, 270.91, 262.2312, 255.1084, 
    252.549, 250.1745, 248.8179, 249.175, 250.1351, 250.8532, 252.4242, 
    253.601,
  274.9923, 273.9767, 272.1117, 267.7691, 261.6054, 256.7401, 254.2479, 
    252.9773, 250.3322, 247.1016, 247.3678, 250.134, 251.1359, 252.5, 253.6561,
  260.9599, 257.9031, 255.2676, 254.6004, 253.4953, 252.7623, 253.9178, 
    248.7867, 251.1697, 248.1497, 249.8076, 252.8124, 251.5941, 249.4843, 
    247.1681,
  261.722, 258.1299, 256.9372, 255.0309, 253.9311, 252.1835, 254.2723, 
    250.8476, 251.2057, 250.5767, 249.6655, 253.5649, 253.9952, 245.436, 
    244.2781,
  268.6425, 260.4238, 258.58, 258.5208, 257.882, 248.4196, 252.7691, 
    253.4775, 255.3015, 253.944, 253.5725, 254.1452, 253.5882, 252.9955, 
    250.125,
  272.8957, 271.3744, 266.6506, 260.2231, 261.587, 259.681, 250.2144, 
    253.6121, 255.3785, 256.6731, 257.6458, 256.6579, 255.319, 254.6923, 
    252.6794,
  274.1315, 272.6917, 272.4397, 264.5256, 261.213, 261.373, 260.8783, 
    246.9533, 250.4477, 255.2516, 257.1027, 258.727, 259.0191, 257.8202, 
    256.4374,
  274.9734, 273.393, 271.8238, 266.9809, 262.1273, 259.7936, 259.7504, 
    258.3078, 256.0253, 256.7451, 255.3314, 256.9402, 258.2315, 258.3076, 
    257.7332,
  275.3852, 274.5092, 273.125, 270.018, 269.0494, 261.5229, 258.2785, 
    256.7127, 256.0091, 256.1512, 256.5267, 256.4804, 257.0273, 257.6273, 
    258.0382,
  275.6936, 274.8172, 273.6031, 272.0057, 271.7979, 264.8845, 257.8197, 
    256.4568, 255.4641, 255.3941, 256.2202, 257.2891, 256.5432, 257.34, 
    257.7262,
  275.5786, 274.8906, 273.8834, 272.3489, 269.9733, 261.6926, 257.9075, 
    256.5609, 255.6988, 255.3686, 255.1569, 256.869, 257.5673, 257.7591, 
    258.7493,
  274.8896, 273.9593, 272.0927, 265.5419, 260.0628, 258.836, 257.1022, 
    257.6334, 255.5409, 253.9203, 253.7389, 255.354, 257.1969, 258.2813, 
    259.1978,
  260.6612, 259.5373, 259.8752, 259.5754, 254.0597, 250.5457, 250.7972, 
    250.3324, 250.8753, 245.8155, 245.5979, 249.4847, 250.2693, 250.6588, 
    250.3581,
  261.2411, 258.5789, 259.7155, 259.0103, 255.3057, 250.5965, 251.9609, 
    250.7394, 252.251, 249.9273, 246.2463, 250.9682, 254.6788, 246.9767, 
    247.6035,
  268.6479, 261.9407, 260.0821, 260.4779, 259.7817, 248.6604, 251.5799, 
    252.5113, 254.0201, 253.5255, 251.8744, 251.7866, 253.2551, 255.1533, 
    253.0041,
  272.8059, 271.686, 267.4766, 261.5757, 261.7722, 259.2473, 248.9751, 
    251.4926, 253.855, 253.6722, 254.8825, 253.2098, 252.5109, 254.4255, 
    253.6125,
  274.0961, 272.6627, 272.0824, 264.1687, 260.8606, 260.1237, 259.4547, 
    245.3231, 248.5216, 251.9686, 253.0046, 253.6294, 253.0698, 253.3279, 
    254.3201,
  274.9075, 273.3331, 271.5778, 266.7773, 263.068, 259.1603, 258.1293, 
    256.1891, 255.1426, 255.4307, 250.1993, 253.2074, 254.6785, 253.0503, 
    253.1036,
  275.3388, 274.443, 272.9879, 269.8426, 269.0577, 260.5249, 257.2573, 
    254.5074, 254.7758, 256.5207, 254.4164, 253.5552, 252.4124, 252.1367, 
    252.2051,
  275.639, 274.7419, 273.5096, 271.9862, 271.2229, 262.3202, 256.7672, 
    253.6895, 252.4698, 254.4166, 256.7665, 254.9229, 252.7404, 253.6735, 
    252.0789,
  275.5239, 274.8087, 273.8095, 272.0161, 266.0287, 258.2513, 256.7906, 
    254.2093, 252.5905, 253.4249, 254.2792, 257.0511, 255.8735, 254.4439, 
    253.9805,
  274.8053, 273.8088, 270.764, 260.3401, 254.8441, 254.9814, 254.3687, 
    257.1588, 254.0696, 251.356, 251.3942, 254.5425, 257.2469, 257.457, 
    256.0044,
  260.8344, 257.6029, 257.4727, 256.989, 252.5001, 249.8268, 249.5446, 
    251.1424, 251.8709, 249.826, 249.4869, 249.8641, 247.2825, 247.159, 
    246.6594,
  259.584, 257.1951, 259.2419, 258.5055, 254.995, 247.1465, 247.6621, 
    249.1485, 250.4962, 252.3519, 250.3378, 251.7066, 253.1434, 246.2754, 
    246.0483,
  267.9873, 258.7915, 256.3967, 258.5504, 258.7138, 246.9976, 247.9688, 
    249.2204, 250.0447, 250.4697, 251.5202, 251.9137, 252.4694, 253.841, 
    251.1201,
  272.7105, 271.1733, 266.0932, 257.7874, 260.1746, 256.6748, 245.4408, 
    249.0706, 251.0269, 253.6126, 253.6361, 252.9898, 252.7616, 254.2621, 
    252.8959,
  274.0734, 272.6405, 271.6358, 261.8291, 258.5529, 258.5706, 256.6526, 
    240.5637, 243.9038, 253.634, 253.5334, 252.3525, 252.373, 253.9891, 
    256.085,
  274.8615, 273.2952, 271.1035, 264.6456, 261.0267, 257.9079, 257.0345, 
    253.6899, 253.2227, 254.8023, 252.1051, 251.7582, 251.533, 253.9937, 
    255.5658,
  275.3037, 274.3824, 272.8051, 268.7818, 268.0089, 258.2939, 256.0163, 
    253.4427, 254.2536, 255.5894, 254.1889, 251.4771, 250.0098, 251.2697, 
    254.5042,
  275.5945, 274.6768, 273.3913, 271.9253, 269.9676, 258.4855, 255.3257, 
    253.7575, 253.785, 255.0414, 254.9641, 251.8834, 250.1987, 250.8887, 
    252.8329,
  275.4858, 274.7327, 273.7351, 270.9006, 261.1939, 254.0381, 253.8663, 
    253.9347, 253.9142, 255.2009, 254.9249, 253.143, 249.9451, 250.4862, 
    252.238,
  274.7397, 273.5959, 268.8953, 256.5496, 251.6212, 251.2423, 251.5301, 
    257.8227, 255.7282, 253.1616, 252.9024, 254.4777, 252.5429, 250.3473, 
    251.0837,
  257.9643, 256.359, 254.4302, 253.3769, 252.8536, 249.7096, 249.1526, 
    248.2792, 249.2503, 246.8241, 251.0113, 251.8082, 248.4862, 247.7899, 
    246.8901,
  257.239, 255.2402, 255.1535, 253.5363, 251.9892, 244.9232, 246.315, 
    247.3459, 248.2895, 250.9505, 251.7511, 253.5495, 253.918, 249.4822, 
    245.4434,
  265.3192, 255.3743, 255.4823, 255.8508, 255.3383, 243.9139, 246.1498, 
    246.4402, 246.9222, 249.1234, 251.9475, 252.8347, 252.7713, 252.3591, 
    248.9868,
  272.4302, 269.8875, 263.6051, 255.5347, 259.5165, 255.4169, 242.1294, 
    247.936, 249.2374, 250.8473, 252.5708, 253.6593, 253.6528, 253.7711, 
    251.9993,
  274.0398, 272.6067, 271.1606, 259.1046, 256.7083, 257.5324, 255.756, 
    239.0868, 242.7602, 253.8003, 254.8163, 253.5419, 252.9224, 253.3984, 
    254.386,
  274.8412, 273.2698, 270.6057, 263.1634, 259.7527, 256.633, 256.2057, 
    254.6437, 252.9848, 253.4457, 251.0191, 251.444, 251.7208, 252.4838, 
    253.2255,
  275.3129, 274.3712, 272.6871, 268.5099, 267.5318, 256.687, 253.9724, 
    252.9766, 252.977, 252.6774, 250.6256, 249.1362, 249.0186, 250.2803, 
    252.3838,
  275.6018, 274.6898, 273.3539, 271.8842, 269.1413, 256.8921, 253.1555, 
    252.2554, 251.2979, 250.6353, 249.5744, 248.8998, 248.2547, 250.378, 
    252.379,
  275.5175, 274.733, 273.7512, 270.5943, 261.1125, 254.7148, 252.7405, 
    252.4203, 251.4375, 250.5155, 248.8315, 249.1976, 248.7023, 251.0126, 
    252.3804,
  274.7895, 273.6048, 269.4061, 259.8495, 255.0423, 253.8687, 252.8767, 
    258.796, 254.8568, 248.3091, 245.4107, 248.0434, 248.8167, 251.0091, 
    252.069,
  255.8112, 253.9482, 252.1409, 252.0758, 249.7414, 245.9064, 246.9535, 
    247.6462, 248.3606, 245.8712, 248.4586, 251.3006, 249.8592, 250.5214, 
    251.0263,
  255.4733, 254.2256, 253.4666, 252.9279, 250.5595, 246.31, 248.1742, 
    248.6521, 249.7864, 249.805, 249.3891, 251.8441, 252.9238, 248.6076, 
    248.4859,
  264.5616, 256.9147, 255.8119, 257.0121, 256.6557, 248.4927, 249.3361, 
    249.1053, 249.2971, 249.907, 251.1833, 252.4292, 252.5819, 252.4088, 
    249.9982,
  272.3496, 269.9356, 265.4708, 259.5405, 261.3406, 258.4985, 251.289, 
    251.6786, 251.2949, 251.8883, 252.7626, 253.0576, 252.686, 252.4112, 
    250.581,
  274.0518, 272.6389, 271.9215, 263.5452, 262.331, 261.7618, 259.6518, 
    248.6517, 248.4271, 253.7717, 255.6631, 254.8245, 254.066, 254.0023, 
    253.7146,
  274.8823, 273.3126, 271.2852, 266.6805, 265.2756, 262.7704, 260.6389, 
    257.9575, 255.2596, 253.9191, 253.6432, 254.5516, 254.2392, 254.1185, 
    253.9785,
  275.3447, 274.4152, 272.8989, 269.8413, 269.5443, 263.157, 259.2749, 
    257.2768, 254.7863, 253.5305, 252.223, 252.4481, 253.3504, 253.3448, 
    253.819,
  275.6213, 274.7337, 273.3808, 271.9268, 270.3308, 262.5194, 258.1492, 
    255.7892, 253.6167, 252.1815, 251.3221, 250.5125, 250.6998, 252.0049, 
    252.8006,
  275.5439, 274.7465, 273.7694, 271.0026, 264.4467, 259.6198, 256.6027, 
    255.1492, 253.4284, 251.7658, 250.2079, 249.3562, 249.691, 250.9269, 
    251.3881,
  274.8233, 273.4397, 270.3768, 263.996, 260.3374, 257.3997, 254.6297, 
    257.4389, 254.9517, 250.0983, 248.5207, 248.7762, 248.2898, 249.5376, 
    250.1806,
  258.7963, 258.4424, 258.7744, 258.8214, 256.5471, 251.9182, 251.421, 
    250.0732, 249.6226, 245.7924, 246.9855, 248.3146, 246.1128, 247.1131, 
    245.2956,
  260.0986, 259.6239, 259.9375, 260.234, 257.425, 255.6631, 256.2794, 
    256.328, 254.1612, 253.4212, 253.2394, 253.5903, 252.6714, 248.5679, 
    247.1252,
  267.5082, 263.3466, 263.951, 265.5009, 262.9861, 261.469, 258.7087, 
    255.9414, 254.8333, 254.279, 253.7061, 254.9831, 253.8475, 252.7435, 
    251.1005,
  272.6729, 271.9062, 270.5418, 268.3108, 266.7047, 263.5661, 256.4066, 
    255.5265, 255.6537, 255.5367, 255.7432, 254.7532, 254.1599, 255.1386, 
    254.1912,
  274.0219, 272.6967, 272.7393, 268.8305, 266.0013, 263.7417, 261.2047, 
    250.926, 250.6951, 255.5913, 256.8593, 255.4624, 254.8844, 254.7421, 
    254.8843,
  274.8271, 273.368, 271.8315, 268.684, 266.3513, 262.5391, 261.0933, 
    257.6909, 253.7658, 250.1006, 252.2336, 253.2371, 253.4536, 253.9198, 
    254.3815,
  275.3047, 274.4081, 272.9798, 270.3276, 269.8531, 262.2134, 257.9666, 
    255.0224, 252.8186, 249.9873, 249.2574, 249.7389, 250.6322, 251.209, 
    252.2886,
  275.6078, 274.7161, 273.346, 271.9153, 269.8503, 258.5659, 252.9126, 
    250.5643, 249.9861, 249.1653, 249.0951, 249.2446, 249.6214, 249.6911, 
    250.6584,
  275.5302, 274.7365, 273.7358, 270.187, 260.7695, 254.5117, 251.1045, 
    250.9918, 251.4072, 251.9189, 250.0421, 248.9606, 248.8004, 249.1503, 
    249.1496,
  274.7581, 273.0882, 269.3007, 259.4597, 254.5565, 251.5212, 249.9803, 
    254.4348, 254.0123, 249.6079, 249.5217, 248.62, 246.4905, 247.0586, 
    247.9381,
  259.1216, 257.5306, 257.9857, 258.6227, 261.6372, 262.1972, 265.5913, 
    262.4041, 259.5857, 254.7055, 255.8359, 255.4968, 251.6699, 250.2198, 
    248.1423,
  259.2369, 258.7725, 259.0841, 260.6042, 261.8218, 260.8578, 265.2902, 
    260.3276, 259.739, 258.308, 258.2841, 259.5206, 258.728, 255.7382, 254.736,
  268.0066, 262.6867, 263.1107, 265.3153, 266.4744, 263.8415, 259.7612, 
    257.9323, 256.1799, 255.5114, 255.4023, 257.2383, 257.1549, 257.1472, 
    255.3228,
  272.8485, 272.6227, 271.6309, 268.4015, 266.5385, 262.1584, 252.2568, 
    253.8526, 253.9313, 253.5916, 254.6716, 254.7788, 255.1294, 255.913, 
    256.6478,
  274.0129, 272.7959, 272.887, 267.1522, 261.3809, 259.671, 257.4654, 
    247.555, 249.3093, 253.5344, 255.827, 254.7755, 254.2419, 254.7574, 
    256.081,
  274.8333, 273.3862, 271.7548, 266.4233, 262.4336, 255.339, 253.2961, 
    251.7136, 250.1312, 247.9436, 250.3282, 252.7641, 252.8152, 253.2641, 
    253.8721,
  275.3148, 274.4349, 272.9177, 269.6022, 268.7963, 255.0677, 250.8396, 
    249.7113, 248.8768, 248.1793, 248.1181, 248.8481, 249.2964, 249.2899, 
    249.5176,
  275.6248, 274.7191, 273.3468, 271.8697, 268.7473, 254.6362, 250.9795, 
    250.2059, 249.937, 249.2942, 248.6291, 248.7723, 248.4946, 248.2899, 
    248.8996,
  275.5365, 274.7294, 273.6751, 269.1196, 257.2006, 252.9794, 251.593, 
    251.9549, 252.4173, 252.4267, 248.9592, 247.4444, 248.5814, 249.4444, 
    248.7545,
  274.751, 272.6334, 267.6136, 256.0881, 252.6248, 252.1895, 251.7416, 
    255.1297, 255.1219, 249.2632, 248.8019, 247.1893, 247.9169, 249.5996, 
    247.7515,
  262.4104, 261.0229, 259.4676, 258.6266, 257.7945, 257.6598, 260.3863, 
    261.252, 260.2466, 255.7185, 253.0901, 250.92, 248.6836, 249.4995, 
    248.6963,
  262.7704, 261.5593, 260.292, 259.5471, 257.6307, 257.742, 259.9851, 
    258.453, 253.7752, 251.7405, 249.9082, 250.4205, 250.2093, 248.4793, 
    248.8636,
  268.8803, 263.7057, 261.9597, 261.5456, 261.7857, 259.2908, 258.2792, 
    255.4653, 251.8292, 251.3409, 250.9917, 250.7628, 250.8018, 250.2575, 
    249.7058,
  272.8828, 272.7766, 271.7002, 267.0188, 265.1195, 263.6876, 253.8304, 
    252.4568, 251.0893, 251.0664, 251.8647, 251.5507, 250.9413, 250.5944, 
    249.4793,
  274.0205, 272.83, 272.9242, 267.5908, 264.5459, 263.317, 258.731, 247.9903, 
    246.1197, 251.0813, 253.2518, 251.6353, 250.585, 250.6566, 250.7793,
  274.8338, 273.3404, 271.8057, 268.3794, 265.4282, 261.0051, 258.3695, 
    253.3687, 249.7478, 247.2105, 247.9314, 250.4727, 250.6619, 250.4483, 
    250.0412,
  275.332, 274.4733, 272.9844, 270.1606, 269.6948, 260.915, 254.3125, 
    250.6249, 249.9948, 249.3969, 250.8187, 250.851, 250.7431, 249.8194, 
    249.325,
  275.654, 274.7784, 273.4254, 271.9008, 269.721, 256.4568, 252.2749, 
    250.4474, 251.1293, 250.8879, 250.9124, 250.3441, 249.0898, 248.1821, 
    249.1798,
  275.6115, 274.7719, 273.6811, 269.9735, 260.0558, 254.3722, 252.1894, 
    252.1999, 253.4983, 252.9817, 248.9648, 247.446, 247.4494, 248.6012, 
    249.1032,
  274.854, 273.3583, 269.1545, 260.1382, 254.2358, 252.3631, 250.9503, 
    254.3257, 255.3372, 248.7723, 247.3183, 244.7065, 245.7459, 249.2017, 
    249.3094,
  264.5597, 263.5631, 262.5639, 261.7055, 259.9709, 259.2642, 259.4214, 
    258.5158, 258.2756, 257.705, 258.4965, 259.0467, 257.6158, 257.1524, 
    254.8467,
  264.6449, 263.3595, 262.5901, 260.7199, 259.1959, 259.0776, 259.6169, 
    258.6995, 258.3653, 258.6444, 257.848, 257.3604, 256.3411, 254.5927, 
    253.3005,
  268.8559, 264.3456, 262.4004, 261.5307, 260.9439, 256.7001, 259.071, 
    259.6631, 258.6336, 258.8668, 258.31, 257.5345, 256.5147, 255.3845, 
    254.4662,
  272.882, 272.451, 270.9302, 265.3814, 261.9087, 262.316, 256.0069, 
    258.9497, 259.6732, 259.425, 259.0225, 258.1902, 256.9239, 255.3506, 
    254.2507,
  274.0646, 272.8646, 272.9351, 267.9417, 262.6097, 262.8721, 261.7906, 
    256.1867, 256.4406, 258.8711, 260.2286, 258.7583, 256.8262, 255.4349, 
    254.2083,
  274.8525, 273.3274, 271.9633, 268.9623, 265.4322, 262.7557, 262.3697, 
    260.7576, 259.8803, 256.7237, 255.4726, 256.1982, 254.7438, 253.4625, 
    252.3048,
  275.3399, 274.4544, 273.0287, 270.3381, 269.6726, 264.4842, 262.6479, 
    261.0073, 258.5481, 255.8596, 254.5514, 253.4045, 253.0745, 250.8174, 
    249.5535,
  275.6346, 274.7586, 273.4129, 271.9176, 271.2283, 265.6425, 263.3476, 
    260.5003, 257.607, 254.7849, 253.6898, 252.2646, 249.8235, 248.7476, 
    248.9613,
  275.6441, 274.7978, 273.7301, 271.4501, 267.8158, 265.4121, 263.2662, 
    259.5625, 257.4221, 255.0138, 251.0081, 248.614, 247.6004, 246.9927, 
    247.4872,
  274.9017, 273.6321, 271.1395, 267.5251, 265.3915, 262.3197, 259.565, 
    258.0498, 256.4901, 248.8311, 244.1672, 244.3395, 244.589, 246.2788, 
    247.9898,
  265.2407, 264.655, 264.241, 263.4622, 262.3985, 261.3045, 261.1509, 
    261.8748, 260.889, 258.5152, 258.6937, 259.2385, 257.0804, 257.3098, 
    256.1159,
  265.8554, 265.4879, 265.1444, 263.7401, 262.3611, 261.5816, 260.8547, 
    260.6625, 260.6155, 260.0595, 259.5453, 259.9607, 258.8253, 256.1897, 
    255.6126,
  269.5488, 265.511, 264.7527, 264.9228, 264.1034, 260.4671, 261.1271, 
    260.4164, 260.6535, 259.6844, 259.1986, 258.8715, 258.311, 257.5377, 
    256.8464,
  272.8311, 272.342, 271.1923, 267.148, 265.0611, 264.0728, 257.884, 
    260.0178, 260.3773, 259.5041, 259.0091, 258.757, 258.3327, 257.3204, 
    257.3863,
  274.1109, 272.9225, 272.9753, 268.5276, 264.0911, 264.3839, 262.5997, 
    256.2508, 255.9038, 258.1102, 260.3705, 259.5936, 258.4316, 257.6749, 
    257.6768,
  274.9167, 273.416, 272.0124, 268.7128, 264.7787, 263.2885, 262.5927, 
    260.185, 257.8189, 255.7437, 256.5744, 257.8457, 257.4153, 257.6111, 
    257.5686,
  275.4204, 274.5158, 273.0392, 269.9416, 268.4223, 263.1436, 261.1203, 
    259.2512, 257.0551, 256.5127, 256.0602, 255.3411, 255.7601, 255.3629, 
    256.1335,
  275.6591, 274.794, 273.3772, 271.8714, 271.0383, 262.8331, 260.675, 
    259.137, 257.1339, 255.966, 255.4472, 256.2641, 255.6097, 254.0623, 
    253.8522,
  275.6313, 274.8133, 273.7004, 271.1104, 265.7036, 262.5968, 261.0765, 
    259.6352, 257.5172, 255.3708, 251.4986, 250.2571, 249.7628, 247.4077, 
    245.2555,
  274.8259, 273.4722, 269.4967, 262.8073, 260.3853, 258.5766, 256.8068, 
    257.1457, 253.0178, 246.4415, 243.1129, 243.0754, 242.4653, 242.8893, 
    243.6976,
  266.6662, 265.8494, 266.7137, 266.0796, 264.5416, 263.9706, 264.7679, 
    265.0001, 264.6272, 263.026, 262.164, 262.5446, 260.8984, 260.0053, 
    259.036,
  266.7181, 267.0807, 266.7684, 264.7794, 263.6586, 264.028, 263.735, 
    262.7918, 264.3935, 263.8695, 263.1497, 263.1228, 262.519, 258.9758, 
    257.2568,
  270.4225, 267.1086, 265.6111, 264.5765, 263.9777, 262.0739, 263.573, 
    263.3231, 262.46, 262.7432, 261.8461, 260.4107, 259.96, 259.2355, 258.4691,
  272.8213, 272.598, 271.3565, 266.1214, 264.1214, 264.1099, 259.5803, 
    262.3239, 261.2523, 260.6715, 259.6963, 259.7014, 259.2991, 259.8675, 
    258.9178,
  274.0953, 272.8992, 272.942, 266.2263, 262.4672, 263.5448, 263.4403, 
    255.926, 257.4993, 259.826, 260.855, 259.9257, 259.0993, 258.6923, 
    258.8838,
  274.845, 273.3827, 271.8083, 266.2119, 261.6289, 260.3186, 261.1981, 
    261.049, 260.3691, 259.7314, 259.4423, 259.9179, 259.6001, 259.3685, 
    258.5893,
  275.3443, 274.4104, 272.8641, 267.7722, 265.0426, 257.7712, 257.502, 
    258.1472, 258.5263, 258.4823, 258.2683, 258.1768, 258.2601, 257.8526, 
    258.1138,
  275.5777, 274.6741, 273.2542, 271.7759, 268.2446, 256.3762, 255.2922, 
    254.1641, 254.293, 253.7989, 253.6747, 254.0224, 253.9143, 254.1076, 
    254.2897,
  275.4993, 274.6783, 273.5836, 268.9317, 257.3884, 253.9603, 252.8754, 
    252.0845, 250.427, 248.5673, 246.4964, 247.2046, 247.4878, 247.3605, 
    246.3638,
  274.6461, 273.1447, 267.3923, 255.5079, 251.0011, 250.0111, 250.6884, 
    254.0674, 249.8515, 244.5471, 243.043, 244.005, 243.7451, 243.9005, 
    243.304,
  262.8457, 260.9058, 261.7915, 260.8709, 258.848, 258.6263, 259.3712, 
    258.6811, 259.2944, 259.7358, 260.9621, 262.2207, 262.0786, 261.9429, 
    261.5314,
  262.6438, 262.1123, 261.6675, 260.4267, 257.0616, 257.5588, 257.1198, 
    256.7075, 256.9452, 258.4185, 260.5415, 262.2247, 262.3345, 260.4638, 
    260.4189,
  270.2337, 264.4969, 261.838, 260.5218, 257.7277, 253.261, 256.0173, 
    255.6254, 256.387, 258.2184, 259.8706, 260.6726, 260.3238, 260.3566, 
    259.8286,
  272.8689, 272.7013, 271.3868, 264.7553, 259.555, 257.3508, 249.741, 
    253.5951, 256.5064, 256.6988, 257.8372, 258.1749, 258.6573, 258.9029, 
    258.966,
  274.1049, 272.873, 272.9084, 265.9138, 260.1693, 258.4537, 257.2456, 
    245.6997, 249.5348, 255.0329, 256.6074, 256.0188, 255.7166, 256.3931, 
    257.5929,
  274.8058, 273.3521, 271.8102, 266.684, 260.8587, 256.7111, 255.6729, 
    253.8008, 252.5063, 252.5381, 251.814, 253.4299, 253.7896, 254.9016, 
    256.0229,
  275.3073, 274.3656, 272.871, 268.6702, 264.5992, 255.3721, 252.5674, 
    252.248, 251.3647, 251.3456, 250.9316, 250.6158, 251.0038, 251.973, 
    253.6138,
  275.5743, 274.6795, 273.2563, 271.763, 266.9468, 253.4585, 250.9479, 
    249.9024, 249.8878, 249.6348, 249.0453, 249.4285, 247.9811, 249.3885, 
    250.7191,
  275.5232, 274.702, 273.6381, 269.6367, 257.5933, 252.2829, 250.9904, 
    250.8368, 250.3498, 249.1511, 247.5337, 247.7917, 245.999, 246.7149, 
    247.9374,
  274.6352, 273.3915, 269.7022, 259.8926, 252.4566, 250.6643, 251.2744, 
    253.3939, 251.1248, 246.9896, 245.6607, 245.7503, 244.1011, 244.8359, 
    245.2243,
  264.8893, 263.8517, 263.0027, 262.5679, 261.2498, 261.4761, 263.0127, 
    260.7621, 259.2281, 257.5973, 256.8898, 256.5677, 254.5369, 253.6516, 
    253.097,
  262.6357, 262.1246, 262.3506, 262.264, 261.3349, 262.11, 261.0873, 
    259.8036, 258.7809, 256.8547, 256.3398, 257.1352, 255.6349, 253.1065, 
    251.7918,
  270.0504, 266.0499, 262.3899, 262.046, 260.109, 257.2448, 258.6647, 
    258.042, 256.2415, 257.3542, 258.067, 257.4006, 256.2868, 254.3527, 
    252.4332,
  272.9554, 272.7169, 271.502, 266.3748, 261.0115, 260.4518, 257.5938, 
    258.5398, 259.4582, 258.135, 257.0754, 255.1962, 254.3393, 252.9578, 
    250.9723,
  274.1466, 272.8748, 272.9607, 268.1123, 263.7215, 265.0367, 264.6922, 
    254.2625, 248.722, 252.3008, 254.005, 252.3304, 251.8183, 250.9123, 
    250.7083,
  274.836, 273.3611, 271.926, 266.7899, 262.9958, 260.7258, 257.9347, 
    254.6561, 250.5364, 247.3195, 247.4725, 249.1021, 249.5267, 249.3947, 
    249.3484,
  275.2837, 274.3084, 272.5962, 264.6499, 260.5052, 254.9001, 252.6735, 
    249.9007, 247.6824, 246.9909, 247.0486, 247.4215, 247.4364, 247.0243, 
    247.8922,
  275.5087, 274.5955, 273.1731, 271.2973, 263.8176, 252.627, 249.8555, 
    247.5482, 247.3495, 247.307, 246.4454, 246.651, 245.1919, 245.7591, 
    247.0466,
  275.424, 274.5644, 273.5081, 267.9715, 254.8753, 250.7261, 249.0011, 
    248.3969, 248.1172, 246.7942, 245.1685, 245.1669, 244.6513, 244.8006, 
    245.7554,
  274.4088, 273.2493, 266.8887, 253.4785, 249.6702, 248.9576, 248.7456, 
    251.6105, 249.3391, 245.6894, 244.8634, 244.8186, 244.0981, 244.038, 
    244.3133,
  266.2425, 265.6275, 264.7428, 264.7109, 266.1557, 266.9893, 267.4908, 
    266.3989, 265.7478, 265.047, 264.7604, 264.7415, 263.2065, 262.3463, 
    260.6259,
  265.6638, 264.9796, 264.5334, 264.5434, 264.3059, 264.2355, 264.738, 
    264.7026, 264.6047, 264.7791, 263.7532, 264.342, 263.4007, 261.1355, 
    259.8646,
  270.2657, 266.1344, 264.4563, 263.7309, 263.0385, 259.9138, 261.4659, 
    261.7562, 262.0367, 263.4814, 263.9907, 263.1946, 262.6186, 262.2739, 
    260.6829,
  272.953, 272.617, 271.103, 265.7383, 262.2428, 262.1606, 259.6958, 
    260.6643, 260.884, 260.6547, 259.8384, 258.0534, 257.4886, 256.2997, 
    253.9946,
  274.1727, 272.8688, 272.9378, 266.7178, 261.8473, 263.3929, 264.1403, 
    255.8383, 253.0513, 253.9181, 255.2915, 253.5012, 252.4738, 251.6478, 
    250.4848,
  274.7953, 273.2926, 271.372, 262.5304, 259.0561, 257.3907, 258.2021, 
    257.3609, 252.4987, 249.0594, 248.3752, 249.5541, 249.0108, 248.4874, 
    247.555,
  275.2055, 274.1847, 271.6212, 261.0301, 258.1143, 253.8371, 252.5278, 
    251.1236, 248.4673, 248.1802, 247.3058, 247.0436, 247.4748, 247.5179, 
    247.4379,
  275.4654, 274.5112, 273.0882, 271.0057, 262.6296, 251.8745, 249.1712, 
    247.9184, 248.0765, 248.0498, 247.1755, 247.4229, 247.4781, 248.1214, 
    248.5841,
  275.4224, 274.5074, 273.5287, 269.2848, 258.017, 253.7244, 251.8431, 
    251.0189, 250.4655, 250.2706, 250.1235, 249.6905, 249.4557, 249.5574, 
    249.0586,
  274.3942, 273.3874, 269.2917, 259.7312, 256.0674, 254.53, 252.8325, 
    253.2884, 253.3216, 252.8206, 253.8773, 252.5094, 251.7712, 252.1113, 
    251.5562,
  264.6592, 262.6892, 262.9083, 264.006, 267.8942, 268.6088, 269.4053, 
    268.5178, 269.3113, 268.2831, 267.9532, 268.4333, 267.6087, 266.375, 
    266.124,
  263.661, 262.606, 262.8318, 264.1349, 265.5603, 267.5012, 268.0684, 
    268.4359, 269.0964, 268.7143, 268.0823, 268.1158, 267.3751, 265.0943, 
    264.5744,
  269.8364, 265.2261, 263.9928, 264.1202, 264.0514, 262.6792, 266.6181, 
    268.29, 268.9378, 268.807, 268.3284, 267.3642, 266.7735, 266.2789, 
    264.6499,
  272.9149, 272.666, 271.0306, 264.1982, 263.524, 264.8367, 263.2237, 
    265.8152, 267.323, 267.621, 267.662, 266.552, 266.1389, 264.868, 263.7723,
  274.1511, 272.8314, 272.5522, 263.2281, 261.5776, 263.2891, 265.4301, 
    261.1682, 260.0291, 265.1084, 266.2554, 265.1356, 264.5935, 263.6693, 
    262.8305,
  274.8324, 273.3003, 270.8427, 261.2659, 260.44, 260.5416, 261.9134, 
    263.3997, 262.4417, 263.0284, 263.2255, 263.0153, 262.7855, 261.8768, 
    260.538,
  275.2611, 274.2339, 271.7979, 263.3034, 261.1882, 258.8136, 258.7995, 
    259.5434, 260.7817, 261.2379, 260.5677, 260.4464, 260.1405, 259.6061, 
    257.9314,
  275.4991, 274.5634, 273.1455, 271.2862, 264.7582, 255.3759, 255.0181, 
    255.739, 256.2597, 257.7843, 258.203, 257.9756, 257.4809, 257.0959, 
    255.851,
  275.4832, 274.5391, 273.6133, 271.1758, 264.7645, 257.5627, 254.1616, 
    254.0769, 254.5583, 254.9308, 255.4182, 255.5841, 255.2631, 254.2342, 
    253.0265,
  274.3776, 273.4853, 272.048, 269.2463, 266.7564, 260.8561, 254.7614, 
    252.6691, 252.5695, 252.0809, 254.6939, 253.9027, 253.4246, 253.608, 
    252.6586,
  260.9147, 259.0072, 258.2674, 261.5195, 265.3336, 265.364, 264.3879, 
    262.19, 260.9261, 264.9815, 261.8655, 265.5195, 265.4269, 264.2748, 
    263.0304,
  262.608, 261.5587, 261.0428, 263.9178, 264.7466, 264.3844, 264.5199, 
    260.6625, 264.9725, 263.9795, 263.2829, 267.2099, 267.1518, 266.4273, 
    262.8465,
  270.6693, 266.3844, 264.3458, 264.8049, 263.502, 264.3238, 265.9572, 
    262.5645, 267.6724, 267.8365, 268.0863, 267.8283, 268.4877, 268.1825, 
    266.0997,
  272.916, 272.7374, 272.155, 266.0941, 263.937, 266.0278, 263.9316, 
    264.5284, 268.1406, 267.998, 267.9897, 267.0894, 267.2645, 266.7527, 
    264.6231,
  274.192, 272.8549, 272.7159, 264.2975, 263.218, 265.8365, 268.1992, 
    265.6404, 265.1392, 267.081, 267.7453, 265.94, 266.1771, 264.7171, 
    264.1661,
  274.8706, 273.3582, 271.4435, 264.257, 264.0308, 264.3765, 265.46, 
    266.4154, 266.3282, 266.34, 266.1547, 266.6581, 265.0673, 262.5366, 
    262.0996,
  275.3018, 274.2596, 272.4755, 267.8691, 265.4504, 263.3114, 265.2173, 
    264.6583, 265.9794, 266.7751, 265.8256, 266.195, 264.2882, 262.6982, 
    260.8703,
  275.4898, 274.5724, 273.1647, 271.6111, 267.0751, 262.0934, 261.7244, 
    262.1704, 264.6186, 265.5384, 265.4191, 265.9117, 264.0492, 261.9456, 
    259.4933,
  275.4741, 274.5065, 273.6378, 271.603, 268.2873, 265.4649, 259.8762, 
    262.4438, 263.0357, 263.7751, 265.3735, 265.549, 263.5808, 260.6349, 
    258.2123,
  274.0003, 272.3876, 269.2792, 266.2061, 268.4, 265.8689, 261.0811, 
    259.8312, 261.5498, 262.2865, 264.0797, 265.009, 262.8974, 260.0839, 
    258.7976,
  263.4403, 261.6751, 260.0878, 261.6962, 261.4827, 258.8357, 261.894, 
    262.5667, 262.6957, 264.527, 261.6078, 263.2551, 263.0839, 262.6795, 
    260.8434,
  264.6704, 263.7505, 263.0406, 261.813, 262.1452, 258.5176, 260.2926, 
    261.6534, 264.4206, 259.2783, 262.2247, 263.9424, 264.7364, 263.6223, 
    258.6528,
  271.02, 267.4683, 264.1356, 263.4605, 261.9326, 258.9397, 258.2966, 
    257.6553, 261.7146, 261.4873, 265.8653, 265.813, 265.442, 264.6101, 
    262.8092,
  273.0164, 272.78, 272.1509, 265.9778, 262.9641, 262.3266, 260.3213, 
    259.9283, 266.0942, 265.5008, 261.2643, 263.102, 264.8386, 265.8542, 
    265.2893,
  274.0905, 272.8073, 272.6193, 264.2244, 263.1494, 263.9582, 264.8078, 
    262.3922, 258.2354, 259.9085, 263.1689, 265.4453, 266.0268, 266.2816, 
    266.0745,
  274.7198, 273.2893, 271.2037, 264.496, 263.8439, 264.3376, 264.5679, 
    263.7266, 262.028, 264.2225, 260.9034, 265.0578, 266.0891, 265.9528, 
    263.8976,
  275.1939, 274.1296, 272.3307, 266.0507, 265.8204, 262.9761, 266.9414, 
    259.7493, 263.4819, 266.2628, 264.12, 264.6342, 265.3777, 263.8763, 
    258.5986,
  275.4001, 274.3998, 273.0263, 271.5958, 268.1662, 261.9098, 261.1832, 
    263.9034, 263.6337, 265.7884, 263.6854, 264.2231, 262.652, 257.8365, 
    253.0533,
  275.3804, 274.3777, 273.4512, 269.7448, 266.8981, 264.6774, 261.0375, 
    262.2039, 265.108, 264.5529, 263.3402, 262.7267, 257.9383, 253.8831, 
    252.1246,
  272.8926, 270.1717, 264.8889, 258.5331, 264.0257, 266.0149, 262.947, 
    264.6832, 263.5311, 263.3327, 262.3007, 259.1952, 255.4152, 253.3392, 
    252.8145,
  262.2574, 259.122, 256.9444, 257.7267, 261.6333, 262.2524, 260.897, 
    263.0356, 264.0122, 262.5397, 262.3483, 264.2555, 262.9067, 262.5276, 
    260.9782,
  263.5565, 260.048, 258.4686, 258.7066, 261.457, 260.8197, 262.2704, 
    263.1588, 263.1105, 262.9351, 261.9463, 264.5318, 264.5899, 260.4211, 
    258.8407,
  271.1882, 266.779, 261.6777, 259.7309, 259.1165, 260.2081, 259.7581, 
    260.6952, 257.143, 258.6623, 263.6471, 264.6555, 263.4528, 262.6112, 
    258.8833,
  273.0678, 272.8069, 272.2226, 263.5295, 260.5089, 261.616, 259.3052, 
    257.8394, 260.4238, 261.7011, 262.0603, 263.1744, 262.2415, 260.7239, 
    259.2201,
  274.028, 272.7515, 272.4825, 264.0121, 261.6508, 262.5047, 263.9442, 
    254.3123, 257.3996, 258.6238, 261.9427, 262.3348, 261.1125, 259.933, 
    258.4822,
  274.6693, 273.2456, 271.2025, 265.9889, 264.9541, 263.2461, 263.8572, 
    264.2258, 260.4338, 262.226, 260.0468, 261.4121, 259.8539, 257.9486, 
    256.0091,
  275.1227, 274.0446, 272.4166, 268.5388, 266.6567, 262.1749, 262.2153, 
    261.4163, 261.4292, 261.2323, 261.3437, 260.1652, 257.5839, 254.3658, 
    252.5477,
  275.3884, 274.3077, 272.8871, 271.6535, 268.9276, 262.2477, 260.0104, 
    260.9319, 259.5046, 260.7841, 259.0962, 256.1029, 253.243, 251.1884, 
    250.3297,
  275.3771, 274.3611, 273.172, 267.855, 264.8043, 263.4726, 259.5654, 
    259.4268, 261.6162, 258.1969, 254.9376, 252.7378, 250.7929, 250.3593, 
    250.3265,
  272.0804, 268.8717, 264.1064, 259.5811, 260.3958, 260.5273, 259.8206, 
    259.4169, 259.6479, 255.9136, 252.4089, 250.6224, 250.1293, 250.1175, 
    251.0812,
  264.1294, 260.8277, 259.5364, 262.2245, 261.4364, 259.1692, 257.8833, 
    260.0049, 260.7996, 259.5551, 259.3129, 260.856, 259.7747, 259.4532, 
    256.8244,
  265.6437, 262.2114, 261.7124, 262.1073, 260.7208, 256.0506, 256.8264, 
    258.7039, 258.1333, 259.2393, 258.1902, 260.7535, 261.595, 257.7089, 
    256.6306,
  271.6338, 268.193, 264.3646, 263.9204, 259.5689, 256.217, 254.5643, 
    257.3425, 256.7497, 257.5531, 257.9575, 259.2551, 260.5034, 261.0331, 
    258.9101,
  273.1191, 272.8336, 272.2304, 265.1183, 261.768, 259.9296, 251.6279, 
    254.5663, 255.7788, 255.7529, 255.4341, 256.1852, 257.6634, 258.6843, 
    259.6507,
  274.0688, 272.7872, 272.1478, 263.5208, 261.4596, 260.8348, 259.1836, 
    250.4274, 251.1048, 253.7672, 254.4035, 254.0018, 255.045, 255.8868, 
    257.5467,
  274.745, 273.2213, 271.0786, 266.4108, 264.2371, 260.4811, 259.4242, 
    259.1529, 255.4264, 256.0633, 252.7401, 253.1986, 252.7377, 253.1399, 
    254.5533,
  275.1872, 274.0844, 272.3992, 268.921, 265.1073, 259.4433, 255.5806, 
    254.3462, 254.3544, 253.4508, 252.0291, 251.7782, 251.6211, 251.211, 
    251.6167,
  275.5311, 274.4417, 272.8774, 271.5728, 268.263, 260.1887, 254.937, 
    252.6169, 251.1551, 250.8244, 249.9281, 250.0934, 249.9526, 250.1673, 
    249.9767,
  275.5401, 274.5079, 273.2482, 267.8585, 265.78, 263.5751, 255.8397, 
    252.7878, 250.5011, 248.9311, 248.2468, 248.8721, 248.5975, 249.2635, 
    249.8258,
  273.3187, 270.725, 266.4364, 262.8655, 262.6288, 262.1324, 256.9604, 
    254.386, 250.9953, 248.0397, 247.5218, 248.0659, 247.5214, 248.0967, 
    250.0058,
  270.4998, 266.5532, 263.4181, 263.7397, 261.9478, 258.9768, 257.3646, 
    256.4405, 256.1381, 255.6144, 255.2911, 257.6304, 255.6956, 255.7138, 
    255.4378,
  270.0447, 268.7886, 265.5664, 264.2931, 263.6129, 259.9294, 258.5184, 
    257.26, 256.704, 257.2002, 255.4273, 257.0789, 258.4174, 253.2897, 
    251.8337,
  272.0103, 270.798, 268.1245, 265.9231, 262.9731, 258.4762, 258.5525, 
    257.1342, 256.8359, 256.4509, 256.2523, 256.5207, 257.8075, 258.0726, 
    254.4865,
  273.1538, 272.8438, 272.414, 267.5108, 264.3133, 261.6074, 256.3464, 
    256.5428, 256.556, 256.0302, 255.6134, 255.1932, 255.974, 256.5534, 
    256.1791,
  274.173, 272.8095, 272.6024, 267.225, 264.6982, 262.4662, 260.6491, 
    252.6187, 251.3512, 255.4453, 255.5965, 254.8803, 254.5554, 254.8256, 
    256.4388,
  274.8683, 273.2365, 271.5502, 267.7016, 265.9932, 262.8187, 260.7298, 
    260.4902, 258.3291, 257.6855, 255.6397, 255.0722, 253.7192, 253.6135, 
    254.2335,
  275.3321, 274.1848, 272.6091, 269.4967, 265.7559, 261.8174, 260.0536, 
    259.2116, 258.5271, 257.9521, 255.7379, 255.0225, 253.4652, 252.3368, 
    253.1728,
  275.6438, 274.6377, 272.9908, 271.403, 266.9213, 260.855, 259.6012, 
    259.7151, 258.7914, 257.7456, 256.9133, 255.2727, 253.0551, 251.4269, 
    251.4857,
  275.6646, 274.6519, 273.3444, 266.9493, 261.9846, 259.3488, 259.1582, 
    260.1435, 259.5427, 258.3826, 257.1898, 255.8298, 253.0983, 251.403, 
    251.5346,
  273.7804, 271.249, 266.9095, 261.6762, 259.0417, 257.5297, 258.3316, 
    260.545, 260.6545, 258.5092, 257.6422, 255.6738, 252.5806, 251.4009, 
    251.3493,
  267.9629, 266.7784, 264.3719, 262.9966, 262.0818, 261.0293, 260.9873, 
    259.9811, 259.2471, 257.4353, 258.1735, 257.4659, 256.0557, 256.5949, 
    256.5068,
  268.0361, 266.8944, 264.1995, 262.3293, 261.3262, 259.0677, 259.5964, 
    259.0942, 257.8063, 257.9761, 255.2951, 256.5823, 257.6806, 255.394, 
    255.1049,
  271.9591, 269.9478, 266.6343, 262.2608, 259.4817, 257.3662, 258.901, 
    258.9432, 257.4883, 255.836, 255.8942, 256.818, 257.6245, 258.9578, 
    258.0712,
  273.1695, 272.856, 272.2545, 264.0477, 259.5402, 258.2601, 255.6287, 
    258.2789, 258.3665, 256.8822, 255.8669, 258.1512, 257.7426, 259.5071, 
    259.8441,
  274.1543, 272.7725, 271.9755, 262.4258, 260.2187, 259.2371, 258.493, 
    254.5225, 255.8629, 258.4485, 256.4085, 257.5789, 259.6024, 259.2866, 
    259.9688,
  274.8459, 273.2219, 270.6342, 262.4244, 261.7557, 260.6333, 259.5399, 
    259.7467, 259.7678, 259.26, 256.4224, 257.6994, 258.6422, 258.4415, 
    258.838,
  275.3422, 274.1572, 272.4617, 267.6754, 262.1852, 258.726, 259.4122, 
    259.3132, 258.9949, 258.1938, 256.8098, 256.8762, 256.9193, 256.6671, 
    255.9908,
  275.6406, 274.6266, 272.9155, 270.3514, 263.9144, 257.4711, 257.6954, 
    258.2103, 258.285, 258.2113, 255.1082, 256.3618, 255.4036, 254.3594, 
    254.0961,
  275.6718, 274.6534, 272.8435, 263.3535, 258.7525, 256.5816, 257.0243, 
    257.4457, 257.5882, 256.8704, 255.8356, 255.0105, 253.5452, 252.0606, 
    250.598,
  273.7513, 270.5625, 264.8357, 258.9409, 257.3997, 255.9411, 255.6714, 
    258.3981, 257.6754, 254.2409, 252.9433, 252.9975, 251.5294, 251.0046, 
    250.2126,
  266.2712, 264.5087, 262.0914, 260.7996, 261.0186, 258.2716, 257.2083, 
    256.969, 256.4764, 255.2878, 257.9663, 257.2467, 252.9974, 251.7706, 
    252.0722,
  267.0563, 266.4961, 264.3817, 262.6199, 262.3684, 259.2404, 259.2311, 
    258.4168, 257.8736, 257.2688, 254.677, 258.1101, 257.5477, 254.7076, 
    249.2683,
  271.9562, 270.4456, 268.5072, 265.0697, 262.3902, 258.9822, 260.8631, 
    259.9731, 259.1624, 257.391, 256.8906, 256.8954, 258.3883, 260.282, 
    254.7839,
  273.1615, 272.8456, 272.3747, 267.7554, 264.6897, 261.7737, 258.3517, 
    260.1555, 260.1322, 258.0615, 256.8111, 258.0725, 258.6368, 257.7196, 
    257.4978,
  274.161, 272.7655, 272.5156, 268.1001, 266.5025, 264.369, 261.3547, 
    255.7824, 256.3053, 259.0883, 256.8965, 255.9015, 256.803, 257.6907, 
    258.4803,
  274.8779, 273.3115, 271.7025, 269.4092, 268.885, 266.8217, 263.7952, 
    261.5648, 259.8686, 258.3352, 255.7048, 254.9542, 254.5043, 255.0961, 
    256.493,
  275.4174, 274.2625, 272.6596, 271.0648, 269.5866, 267.2784, 265.2447, 
    263.1816, 260.8658, 258.8808, 256.7211, 255.4382, 253.9815, 253.2546, 
    253.6265,
  275.7305, 274.7298, 273.0547, 271.6508, 270.7144, 268.4345, 266.1554, 
    264.5533, 262.3191, 260, 257.0186, 254.8783, 253.4573, 252.0645, 251.3608,
  275.7221, 274.7558, 273.4745, 271.9347, 270.9664, 269.3673, 267.4919, 
    265.9638, 264.044, 261.1582, 257.6751, 254.9928, 252.8305, 251.5773, 
    250.3658,
  274.2288, 273.1234, 272.3574, 271.9905, 271.1446, 269.8258, 268.1918, 
    267.1057, 265.4977, 261.1622, 257.4845, 254.8365, 251.8508, 250.0934, 
    251.0638,
  271.6324, 271.3039, 271.283, 271.4643, 271.2443, 270.4384, 269.6855, 
    267.9865, 265.4085, 261.6975, 261.7135, 261.02, 258.3385, 256.9769, 
    254.787,
  271.4671, 271.773, 271.8091, 272.0527, 272.0757, 271.2844, 270.5646, 
    269.6203, 267.9942, 264.9157, 262.7686, 262.1148, 261.2005, 258.4181, 
    255.39,
  272.2341, 271.8208, 271.7916, 272.1471, 272.3684, 271.0335, 270.909, 
    270.7761, 269.3991, 267.7673, 265.4146, 263.5037, 262.1815, 261.678, 
    260.1594,
  273.2578, 272.9193, 272.6422, 271.6818, 272.0329, 272.0127, 270.5396, 
    270.0525, 269.3518, 268.2069, 266.1874, 264.5212, 262.9262, 261.7917, 
    260.9164,
  274.1844, 272.8031, 272.8385, 271.0718, 271.3206, 271.4247, 271.302, 
    268.5738, 268.052, 269.701, 268.8488, 266.4608, 264.0062, 262.2094, 
    261.4095,
  274.8939, 273.3645, 271.9652, 270.4288, 270.712, 270.143, 270.1467, 
    270.1898, 270.049, 269.8733, 268.9166, 267.3048, 264.6393, 262.4395, 
    260.9646,
  275.393, 274.2977, 272.7029, 271.0853, 270.0209, 268.6955, 268.3815, 
    269.0722, 269.1212, 269.2562, 268.5125, 266.7482, 263.8146, 261.4726, 
    259.9552,
  275.7032, 274.7193, 273.0913, 271.127, 269.1124, 267.6096, 267.0103, 
    267.5292, 267.0915, 267.8106, 267.6212, 265.4853, 262.2576, 259.6841, 
    258.1754,
  275.6298, 274.7214, 273.2202, 268.1247, 265.7203, 265.6557, 265.1318, 
    265.2751, 265.5482, 265.6293, 264.6335, 262.1096, 259.0554, 257.3088, 
    255.5467,
  273.787, 271.9317, 269.1145, 266.3591, 263.8807, 263.2921, 262.4915, 
    263.4159, 263.1162, 261.0164, 259.9555, 257.1571, 255.3248, 253.6367, 
    251.6045,
  272.4596, 271.5997, 270.9995, 269.776, 267.6528, 266.0602, 265.7303, 
    265.1786, 268.8505, 268.7142, 268.9482, 268.1056, 264.3124, 261.489, 
    258.7935,
  272.2067, 271.8253, 271.1846, 269.6165, 266.5595, 264.0741, 264.0075, 
    262.7773, 263.5245, 266.0105, 267.0964, 268.2112, 266.6131, 262.1943, 
    259.7005,
  272.2659, 271.7318, 271.3937, 269.8713, 267.1731, 261.9691, 263.643, 
    261.8192, 262.6575, 265.6709, 266.9338, 267.9755, 267.8977, 266.0953, 
    262.4933,
  273.3202, 272.9538, 272.6368, 270.2154, 267.5792, 264.3812, 258.6301, 
    260.8528, 260.5041, 262.6954, 265.3351, 267.1226, 268.0351, 267.5221, 
    264.4298,
  274.1886, 272.8131, 272.8404, 269.968, 267.9786, 264.8994, 261.9405, 
    254.677, 257.067, 261.2842, 263.9611, 266.1966, 267.7681, 268.4279, 
    267.1399,
  274.9258, 273.354, 272.0211, 270.5083, 269.8557, 266.1922, 262.7203, 
    260.9218, 257.5494, 258.5655, 260.7787, 265.07, 266.8274, 267.8171, 
    265.782,
  275.4129, 274.338, 272.7156, 271.3125, 270.1924, 267.181, 263.8548, 
    261.2921, 258.5669, 256.954, 258.7262, 262.0004, 265.2544, 264.6584, 
    262.6757,
  275.7471, 274.7563, 273.1063, 271.623, 270.6003, 267.8008, 264.9394, 
    262.1764, 258.4287, 256.01, 257.9823, 257.2654, 258.8003, 259.2201, 
    258.6352,
  275.657, 274.7653, 273.4201, 271.7288, 270.0248, 267.9163, 265.176, 
    262.7052, 259.8239, 256.764, 255.5548, 256.9433, 255.102, 254.6893, 
    254.6283,
  274.1996, 273.3162, 272.48, 271.6348, 270.1624, 268.329, 265.9933, 
    264.0922, 261.7431, 257.3102, 254.461, 253.676, 252.7961, 252.2189, 
    252.1092,
  273.0796, 272.4509, 272.3637, 272.6858, 272.3289, 269.3365, 267.5626, 
    264.7215, 263.2098, 263.5432, 259.2875, 264.0744, 265.5887, 265.2071, 
    263.8026,
  272.6207, 272.2422, 272.0025, 272.2403, 272.3311, 270.3112, 268.0573, 
    264.6255, 261.4969, 260.8024, 261.6063, 264.4177, 265.6373, 264.1667, 
    262.3287,
  272.3326, 271.8331, 271.7316, 271.7566, 272.2755, 269.9303, 268.1984, 
    265.6429, 262.5739, 261.6035, 261.9782, 264.0118, 264.3506, 265.9223, 
    265.127,
  273.396, 273.011, 272.702, 271.4425, 271.7963, 271.8256, 268.1864, 
    265.8034, 263.8527, 262.7866, 262.6552, 261.3846, 262.4756, 264.565, 
    266.232,
  274.2325, 272.8451, 272.8869, 271.1067, 271.0972, 271.5826, 270.6469, 
    264.5916, 262.0725, 265.0544, 263.495, 262.0026, 262.9316, 264.6392, 
    266.1054,
  274.985, 273.3604, 272.0753, 270.8485, 270.8016, 270.7479, 270.7433, 
    269.5173, 267.0618, 264.2132, 262.5278, 262.2552, 261.844, 263.0703, 
    265.5786,
  275.4245, 274.3872, 272.7511, 271.2065, 270.4366, 269.6999, 269.9692, 
    269.6717, 268.2071, 265.648, 263.0215, 261.7811, 261.4033, 262.0831, 
    263.2088,
  275.7647, 274.7894, 273.1557, 271.0914, 269.3202, 268.0394, 268.4532, 
    268.969, 268.1479, 265.8555, 263.546, 261.9513, 260.7975, 259.9633, 
    261.4048,
  275.6445, 274.7802, 273.1397, 268.8, 266.2719, 266.2634, 266.7113, 
    267.0662, 266.5314, 265.0356, 263.0746, 261.7151, 260.8687, 259.4434, 
    258.4847,
  274.099, 272.6836, 270.9059, 267.8355, 264.8507, 264.4795, 264.5747, 
    264.7752, 264.782, 262.9632, 261.9831, 261.4899, 260.2283, 259.4645, 
    257.8573,
  273.004, 272.0264, 271.4937, 269.9207, 268.2594, 268.5684, 268.5517, 
    270.6173, 269.5021, 267.0661, 263.0072, 263.2569, 260.485, 264.2976, 
    265.6456,
  272.3794, 271.941, 270.9648, 269.2264, 265.8105, 264.9597, 266.7562, 
    268.7094, 269.4276, 267.7461, 265.8391, 264.8265, 262.6133, 260.46, 
    264.3622,
  272.4045, 271.8245, 271.3887, 268.797, 266.1307, 264.4929, 265.7836, 
    267.2866, 268.2964, 267.5254, 266.5516, 266.0961, 264.5383, 261.8435, 
    262.2845,
  273.4717, 273.0598, 272.6906, 268.5329, 265.3898, 264.968, 263.7174, 
    264.0534, 265.5497, 266.1781, 265.7224, 266.1321, 265.6078, 264.1588, 
    263.868,
  274.2237, 272.8575, 272.778, 267.7458, 264.7918, 263.4092, 263.9094, 
    261.0913, 261.3076, 264.644, 265.4136, 265.5833, 266.1309, 265.3413, 
    264.0559,
  274.9709, 273.3263, 271.9881, 268.3059, 266.6886, 261.2718, 261.7898, 
    262.03, 261.7839, 262.0044, 261.4289, 262.6393, 264.1204, 265.3431, 
    264.5633,
  275.3778, 274.369, 272.7284, 270.7158, 266.4495, 260.5146, 259.2389, 
    258.7979, 258.1723, 258.0004, 257.8876, 259.5547, 261.0368, 262.7711, 
    264.1546,
  275.7262, 274.7593, 273.1377, 269.5965, 264.082, 258.7634, 257.5067, 
    256.725, 256.0228, 255.2883, 255.1617, 256.3995, 258.4186, 260.4736, 
    262.8987,
  275.5856, 274.7518, 272.457, 263.994, 258.3517, 258.0456, 256.7824, 
    255.8443, 254.2678, 254.4369, 253.3744, 253.4497, 255.0105, 258.099, 
    260.7413,
  273.5169, 270.9178, 266.8714, 261.3337, 258.0386, 256.2104, 254.8168, 
    255.9016, 254.9674, 252.026, 250.8954, 251.6782, 252.3655, 255.1006, 
    258.3778,
  265.5678, 261.2939, 259.0284, 258.8555, 258.0294, 257.3604, 256.2166, 
    256.9847, 258.1767, 258.3463, 260.1208, 263.4817, 263.9135, 263.4058, 
    261.8929,
  269.1344, 264.3975, 259.8787, 258.3176, 257.5347, 254.3686, 254.5078, 
    255.2615, 255.8919, 256.2273, 256.8349, 261.2032, 262.8769, 261.4939, 
    260.8553,
  272.4056, 271.7608, 268.8876, 259.6206, 257.0319, 252.65, 254.8095, 
    253.3602, 253.1218, 253.5682, 254.4135, 257.3488, 260.5376, 262.9039, 
    263.3429,
  273.4739, 273.0233, 272.3392, 260.632, 257.5777, 255.3913, 250.6642, 
    253.1943, 253.4314, 252.9157, 252.6831, 254.4972, 257.6464, 260.8633, 
    263.1727,
  274.1773, 272.8236, 272.1996, 261.7539, 259.7793, 255.826, 254.1027, 
    247.5111, 249.5138, 254.4805, 253.283, 252.417, 254.0196, 257.6427, 
    262.4366,
  274.9459, 273.249, 271.6603, 265.4315, 264.3839, 256.2694, 254.138, 
    252.9567, 251.0756, 249.0057, 248.4575, 250.2777, 251.7903, 254.2785, 
    259.2756,
  275.338, 274.3228, 272.668, 269.5275, 264.2435, 256.6111, 254.4645, 
    253.3644, 252.4006, 250.3571, 249.0071, 249.1053, 250.7305, 251.8982, 
    256.057,
  275.6901, 274.7267, 273.105, 268.2637, 262.9548, 257.1605, 255.2429, 
    253.9747, 252.7978, 251.1538, 249.4908, 248.5315, 248.9864, 250.3547, 
    254.6932,
  275.5666, 274.7173, 271.7454, 262.2274, 258.405, 257.6218, 255.2342, 
    254.3321, 253.3785, 252.6337, 249.5316, 247.8519, 247.4977, 249.342, 
    253.6859,
  272.9431, 269.3895, 265.9796, 260.463, 258.0209, 257.1842, 254.9016, 
    255.5695, 255.3539, 250.9301, 248.4639, 247.0012, 246.2669, 248.0546, 
    251.9288,
  266.5688, 264.3759, 262.9661, 262.4084, 262.3802, 260.717, 257.763, 
    253.2284, 251.8416, 249.4835, 248.675, 251.1443, 255.7877, 260.1599, 
    263.098,
  269.8012, 267.2689, 264.6406, 263.2304, 262.6072, 260.2711, 256.7721, 
    253.4718, 252.4776, 251.7141, 248.7118, 250.6686, 253.1672, 254.3337, 
    258.8436,
  272.4227, 271.8224, 270.1371, 264.3048, 263.6396, 258.7159, 258.2115, 
    255.2329, 254.3358, 252.0855, 251.5608, 251.115, 252.4333, 255.3546, 
    258.371,
  273.5376, 273.0475, 272.445, 264.6822, 263.4133, 260.7733, 256.8062, 
    257.1905, 256.0132, 254.8274, 253.3506, 251.4114, 251.5405, 253.0319, 
    256.8259,
  274.1474, 272.8101, 272.3431, 263.5808, 263.2704, 262.51, 258.9848, 
    253.9577, 252.1067, 255.7744, 255.118, 251.841, 250.461, 251.4373, 
    254.4015,
  274.8999, 273.2306, 271.7749, 266.5141, 265.5345, 261.0495, 259.7552, 
    257.3482, 254.306, 251.4759, 251.4423, 251.5459, 249.832, 250.2114, 
    252.8791,
  275.2861, 274.2714, 272.6561, 269.2343, 264.7709, 258.4262, 258.0215, 
    256.5746, 255.2008, 252.4767, 252.5463, 251.7982, 250.4508, 249.2041, 
    251.5761,
  275.6322, 274.6635, 272.9759, 266.9547, 261.9042, 256.995, 255.8746, 
    255.7481, 254.5948, 253.241, 251.6864, 251.5872, 250.2834, 248.6053, 
    251.4656,
  275.4982, 274.4951, 269.9597, 260.5195, 257.5942, 255.7898, 255.4685, 
    255.7378, 254.6769, 252.7353, 250.8628, 250.8603, 249.19, 248.5074, 
    250.9494,
  271.8731, 266.8202, 263.2427, 258.5284, 256.5452, 255.6449, 254.8209, 
    256.4328, 255.4832, 252.1666, 250.186, 250.2325, 248.034, 247.4687, 249.57,
  265.4331, 262.2225, 260.3449, 259.5638, 259.9959, 262.0825, 263.1051, 
    261.2889, 258.8951, 256.7518, 254.8659, 251.6491, 252.6794, 257.5345, 
    261.9726,
  269.2459, 265.9123, 261.96, 259.7552, 261.0584, 262.9616, 261.8701, 
    259.2767, 257.7762, 256.0988, 252.763, 251.6375, 254.3012, 257.0725, 
    260.9395,
  272.4391, 271.8495, 269.9358, 261.2413, 262.1333, 259.6032, 260.5458, 
    257.8774, 255.8885, 253.9258, 252.7342, 251.9541, 255.0867, 259.2569, 
    262.304,
  273.561, 273.0447, 272.3597, 261.894, 261.3588, 260.7733, 255.6193, 
    256.1195, 254.6065, 253.5188, 252.4182, 251.945, 255.7908, 258.97, 
    261.6917,
  274.04, 272.7445, 272.024, 259.9817, 260.4264, 260.3793, 259.1977, 
    252.1492, 249.112, 253.1942, 253.0557, 252.1623, 254.8533, 257.9612, 
    260.5667,
  274.7899, 273.1429, 271.6326, 264.264, 262.6223, 258.1986, 259.5781, 
    258.7417, 254.7974, 252.9281, 251.0202, 252.3539, 253.6606, 257.0692, 
    259.6796,
  275.1676, 274.1366, 272.5185, 267.1819, 262.7788, 257.8483, 259.2163, 
    257.8886, 255.6894, 253.7244, 253.731, 253.291, 254.1976, 257.1319, 
    260.0213,
  275.5217, 274.507, 272.2615, 265.5664, 261.6176, 258.9225, 258.0486, 
    256.3205, 254.0208, 253.9545, 253.2143, 253.5253, 254.7215, 256.8365, 
    259.9364,
  275.4052, 274.057, 267.4467, 259.9704, 259.0703, 257.8808, 257.229, 
    254.8125, 252.9152, 252.3891, 251.9412, 252.6357, 253.7778, 256.4659, 
    258.9464,
  270.7278, 265.0205, 261.0887, 258.1487, 256.9404, 256.5794, 255.1591, 
    255.5409, 253.0135, 250.8527, 250.8045, 251.7281, 252.5118, 255.6784, 
    259.4039,
  262.9224, 259.2565, 257.5345, 256.2971, 257.3144, 257.0507, 256.0577, 
    254.9044, 258.5677, 262.8305, 263.6501, 262.225, 259.9098, 258.6584, 
    255.4809,
  268.8197, 264.9309, 259.774, 256.9202, 258.1595, 257.9413, 258.8973, 
    257.1017, 259.9859, 263.1914, 262.7778, 261.2563, 260.1078, 255.8154, 
    254.6879,
  272.4308, 271.7027, 268.7384, 258.4503, 258.3854, 256.1313, 258.8834, 
    258.569, 260.3019, 262.1667, 261.3251, 260.3324, 259.2499, 257.546, 
    256.4169,
  273.5548, 273.0569, 272.0215, 260.1152, 258.7231, 259.0836, 255.3081, 
    257.9124, 259.3454, 260.264, 258.5654, 258.2762, 259.1197, 257.7669, 
    257.819,
  273.983, 272.7293, 271.5421, 259.5219, 258.7583, 258.8642, 260.0253, 
    251.9449, 251.1087, 257.928, 257.6068, 254.3563, 256.7789, 258.9779, 
    258.8822,
  274.7801, 273.1134, 271.3786, 263.9816, 260.8477, 256.9506, 256.8019, 
    257.5837, 253.2749, 252.6988, 251.5481, 253.5641, 259.2676, 260.3279, 
    259.9906,
  275.1242, 274.08, 272.2512, 266.3872, 261.0217, 255.6577, 254.4093, 
    253.9016, 253.0359, 251.0117, 251.8646, 256.6381, 261.9817, 263.1532, 
    262.6781,
  275.5082, 274.4698, 271.3953, 265.2824, 260.1777, 256.0002, 253.8365, 
    252.6324, 251.338, 252.3239, 255.6312, 260.7573, 262.9539, 263.4315, 
    264.1967,
  275.4556, 274.1914, 266.7271, 260.7746, 257.6503, 256.1703, 254.9207, 
    254.059, 253.645, 255.0576, 258.7574, 262.4013, 262.8734, 262.5997, 
    263.3366,
  271.1384, 265.5701, 261.3153, 258.764, 256.5055, 255.8689, 255.4621, 
    257.0471, 257.2872, 257.2576, 258.8794, 261.2069, 261.496, 262.8839, 
    264.1061,
  264.8289, 258.7737, 256.663, 256.4896, 258.6392, 259.7493, 261.3888, 
    261.796, 262.3678, 261.7625, 261.8768, 262.93, 263.2613, 263.4202, 
    262.5866,
  269.2398, 263.1942, 259.3157, 257.7899, 258.9247, 259.3901, 261.9821, 
    262.1827, 263.1653, 264.191, 264.6466, 265.6638, 265.7126, 263.0924, 
    262.8982,
  272.5125, 271.553, 267.7844, 258.9467, 258.4926, 257.4811, 261.0891, 
    261.5987, 261.773, 262.217, 262.5659, 263.3565, 263.9716, 264.6484, 
    263.773,
  273.5276, 273.0583, 271.5497, 259.9957, 259.1816, 260.1873, 259.254, 
    260.9856, 260.3329, 260.3678, 260.2019, 260.6254, 261.6362, 262.3808, 
    262.6377,
  274.0425, 272.7548, 271.0006, 259.771, 259.5549, 259.8556, 261.6273, 
    256.5574, 255.9823, 259.9211, 259.3234, 258.0045, 258.6094, 259.8763, 
    261.0697,
  274.8515, 273.0818, 271.0179, 263.7743, 261.7552, 258.8523, 259.2209, 
    259.717, 256.3279, 257.2573, 256.9336, 257.7666, 257.8685, 257.6317, 
    258.702,
  275.1523, 274.0702, 271.9162, 266.1227, 261.6807, 259.2796, 258.1819, 
    258.0301, 257.2612, 255.4872, 256.2351, 257.617, 258.4142, 256.8228, 
    259.0505,
  275.5241, 274.5176, 270.9398, 264.5112, 260.7328, 259.2429, 258.062, 
    259.88, 259.3404, 257.8473, 258.0567, 256.772, 256.4615, 259.9711, 
    261.5803,
  275.5351, 274.3012, 265.7678, 260.3455, 258.4181, 257.7898, 259.1076, 
    258.8696, 261.0014, 260.3498, 260.6391, 260.5095, 260.7881, 259.6796, 
    263.0858,
  271.3733, 265.7154, 260.5654, 258.2099, 258.1538, 258.4989, 259.959, 
    263.3842, 262.5783, 262.9738, 263.718, 264.0334, 263.4646, 263.1224, 
    263.3861,
  263.1146, 260.264, 259.1088, 259.3197, 260.9997, 258.463, 257.3599, 
    257.3499, 259.2878, 261.4538, 262.6483, 260.2083, 254.2193, 256.3394, 
    255.2554,
  268.3987, 263.8734, 261.3997, 260.3949, 261.0691, 258.036, 257.6557, 
    257.2346, 258.1402, 261.1021, 261.6917, 263.6595, 260.9525, 253.9549, 
    254.3364,
  272.4818, 271.5287, 268.5902, 261.3509, 258.9988, 256.499, 258.0798, 
    257.6437, 258.0279, 258.7343, 260.1754, 263.3601, 262.302, 259.3235, 
    256.9428,
  273.4603, 273.0267, 271.6052, 262.3531, 260.0797, 259.1687, 256.3397, 
    257.0371, 258.1252, 258.2524, 258.58, 261.5667, 264.6292, 262.7887, 
    258.6578,
  274.0781, 272.7362, 271.2475, 262.2071, 261.6562, 260.8194, 260.4108, 
    256.3673, 256.6302, 259.6693, 259.0844, 259.6458, 262.8114, 263.9437, 
    261.7684,
  274.8983, 273.0894, 271.1735, 266.2833, 263.5358, 260.8676, 260.4786, 
    261.793, 261.3839, 260.4308, 258.7155, 258.9676, 260.9755, 263.0161, 
    263.808,
  275.2755, 274.1144, 272.0805, 267.5629, 262.8002, 260.7024, 260.1451, 
    261.7377, 262.7223, 261.6907, 259.5614, 259.2019, 260.6072, 263.1434, 
    264.4569,
  275.6122, 274.629, 271.5901, 266.0526, 262.408, 259.6975, 259.4246, 
    262.0988, 263.8627, 263.6167, 261.1852, 260.1938, 260.6135, 262.6165, 
    264.0642,
  275.6644, 274.4819, 269.3436, 264.3114, 261.0353, 258.5242, 258.8655, 
    261.617, 264.0198, 264.4742, 263.1576, 262.0676, 261.8641, 262.5905, 
    262.0606,
  273.0327, 269.8184, 266.2553, 263.1768, 260.8419, 257.6458, 258.1565, 
    262.2934, 264.163, 264.4337, 264.2425, 263.4423, 263.4478, 263.7328, 
    263.4362,
  266.2335, 265.3088, 265.3501, 264.1474, 263.0832, 263.0704, 262.2311, 
    260.1571, 258.354, 259.5608, 260.2862, 258.4133, 257.9007, 258.2858, 
    258.7175,
  269.8418, 268.3527, 266.4094, 265.5476, 265.528, 264.3502, 263.5409, 
    260.5603, 257.338, 260.6025, 260.9934, 259.6624, 259.9886, 256.428, 
    257.218,
  272.5475, 271.7992, 270.4461, 266.9377, 265.3478, 264.4486, 264.7978, 
    261.8543, 257.7495, 261.8857, 261.5217, 261.653, 258.9273, 259.5449, 
    258.0392,
  273.5401, 273.0859, 272.3465, 268.7768, 267.8928, 267.1648, 263.6712, 
    259.1834, 256.8013, 260.9504, 262.3183, 262.5904, 261.6672, 259.7401, 
    257.1674,
  274.1934, 272.832, 272.3981, 269.6283, 268.85, 266.3746, 264.5766, 253.167, 
    253.9677, 260.4031, 262.7324, 263.0007, 264.3415, 260.8756, 259.7398,
  275.0196, 273.2922, 271.8673, 270.3536, 268.7023, 264.881, 259.7509, 
    257.7041, 256.2721, 260.8896, 262.0851, 262.6838, 264.4594, 262.9882, 
    262.5041,
  275.4374, 274.2528, 272.5655, 269.9424, 266.7156, 261.9562, 258.7858, 
    259.6694, 260.5366, 263.2982, 262.8729, 262.7226, 263.8015, 265.321, 
    264.6647,
  275.7069, 274.7485, 272.5807, 268.1159, 264.2169, 259.0583, 259.1005, 
    260.5234, 261.9431, 263.8412, 263.1612, 262.3615, 263.244, 264.4362, 
    265.2776,
  275.741, 274.5941, 270.9568, 265.1685, 261.201, 257.5909, 259.0809, 
    260.4842, 263.6831, 264.9462, 263.7114, 262.5851, 262.6853, 263.3829, 
    263.8184,
  273.5663, 271.5825, 269.5353, 264.439, 262.3588, 256.4705, 258.7192, 
    262.7761, 264.5321, 264.1199, 263.4034, 262.9695, 263.7485, 263.8239, 
    264.114,
  268.8901, 268.4638, 269.2775, 268.1565, 267.933, 268.5788, 268.7025, 
    268.937, 267.0258, 261.5115, 257.4364, 261.0507, 260.4634, 259.5105, 
    259.1546,
  270.96, 270.4647, 268.8625, 267.3304, 265.8146, 266.4774, 268.0849, 
    267.4554, 264.7491, 258.9729, 257.3407, 262.418, 261.2827, 258.9667, 
    258.7477,
  272.6295, 271.9315, 270.4437, 265.3108, 264.0425, 262.2029, 264.232, 
    263.6559, 258.7183, 257.341, 260.6284, 262.3046, 262.2148, 262.7856, 
    261.6454,
  273.6205, 273.1252, 272.3066, 264.4813, 262.6042, 261.9077, 258.6115, 
    259.5579, 256.6727, 257.9183, 258.9472, 262.2851, 263.0403, 263.2287, 
    261.6672,
  274.3681, 272.9029, 272.241, 263.7742, 262.5876, 259.8319, 260.2379, 
    254.1767, 252.4258, 258.5881, 262.5816, 262.5267, 263.3041, 262.7521, 
    263.7011,
  275.2757, 273.4576, 271.7143, 266.4415, 264.3562, 260.433, 259.8563, 
    260.2646, 259.4381, 258.9598, 262.4027, 261.0113, 263.0511, 263.1483, 
    263.0412,
  275.6413, 274.4007, 272.5144, 268.2284, 264.8783, 260.554, 259.6168, 
    260.9137, 261.7873, 262.9791, 263.2071, 261.7805, 263.9822, 263.4146, 
    262.4637,
  275.89, 274.8363, 272.5361, 268.4245, 265.6317, 260.1191, 259.4145, 
    261.4793, 263.3357, 264.0297, 264.0866, 262.8179, 264.4952, 263.6563, 
    262.8438,
  275.9028, 274.642, 271.3777, 268.4379, 266.3928, 261.5309, 259.271, 
    261.9998, 263.668, 265.0199, 264.5289, 263.9141, 265.0889, 265.1643, 
    265.1969,
  273.8026, 271.9905, 270.1974, 269.3488, 266.8406, 260.7952, 258.889, 
    264.0885, 265.0849, 264.559, 265.0276, 265.5339, 265.8744, 265.5094, 
    263.1521,
  268.0151, 263.5781, 263.569, 262.0294, 260.3197, 260.8073, 258.8292, 
    261.6501, 262.1783, 262.2623, 261.9235, 263.1261, 262.4112, 261.5862, 
    260.7566,
  270.8189, 267.2523, 266.0076, 264.2726, 262.6527, 260.2202, 259.0439, 
    257.0197, 259.5187, 261.325, 261.5841, 262.7516, 261.9612, 259.2154, 
    259.5318,
  272.7271, 271.9615, 270.6349, 266.249, 264.5664, 261.0312, 258.6096, 
    258.8748, 260.6553, 260.3941, 261.1312, 263.3781, 263.0649, 262.7276, 
    261.9609,
  273.6041, 273.1164, 272.4977, 267.8557, 267.787, 265.3095, 259.1901, 
    257.1638, 260.7358, 262.2207, 263.0271, 263.9658, 264.0046, 264.5041, 
    264.2512,
  274.5017, 272.9302, 272.635, 269.0119, 268.9951, 266.7992, 261.428, 
    257.4167, 259.2246, 264.0095, 264.5773, 263.9256, 264.1704, 264.1535, 
    264.5631,
  275.4318, 273.5728, 271.9635, 270.7944, 269.0336, 266.0402, 262.4764, 
    262.8418, 263.0513, 263.9798, 263.7081, 262.9694, 264.097, 263.592, 
    263.8536,
  275.8579, 274.5467, 272.6559, 270.9945, 267.3816, 263.7236, 261.4832, 
    263.1921, 264.3811, 264.0122, 263.364, 263.1368, 263.8627, 263.9275, 
    264.3161,
  276.1682, 274.9383, 272.5764, 270.1592, 265.2383, 262.4072, 261.6497, 
    264.2484, 263.8245, 263.6548, 262.8225, 263.6528, 264.1755, 264.837, 
    264.7079,
  276.1449, 274.7163, 270.5421, 268.2893, 262.3456, 260.0002, 261.901, 
    264.7497, 264.177, 263.0822, 262.8664, 263.4496, 263.7949, 264.9561, 
    265.7466,
  273.9952, 271.7804, 268.3294, 266.9213, 260.0687, 260.1709, 262.1488, 
    266.2551, 264.9153, 262.4313, 261.955, 262.4365, 263.252, 263.8178, 
    265.1867,
  268.8049, 269.2992, 270.374, 268.1164, 264.8791, 264.3607, 260.6353, 
    261.0582, 261.9038, 262.6039, 261.9936, 262.2327, 262.7127, 260.7356, 
    259.1028,
  270.752, 271.3704, 270.3431, 266.8257, 265.1938, 261.4177, 261.522, 
    258.997, 259.1765, 259.7603, 261.535, 262.8053, 263.2652, 262.0092, 
    260.7644,
  273.0499, 272.1148, 271.119, 267.2068, 263.9258, 262.2752, 260.2226, 
    260.8321, 260.3318, 261.9243, 262.153, 262.8177, 262.8541, 261.9548, 
    261.2101,
  273.7527, 273.2203, 272.5393, 268.0625, 263.5852, 261.7308, 257.4505, 
    260.4218, 261.6065, 262.0932, 262.0652, 262.4898, 262.5879, 262.4839, 
    262.8531,
  274.6702, 273.0783, 272.5764, 267.2412, 263.0924, 261.6039, 261.2313, 
    256.3255, 258.2193, 262.6198, 262.8761, 262.0706, 262.7409, 263.0235, 
    262.511,
  275.5861, 273.7318, 271.8719, 268.6719, 265.5439, 261.0524, 260.256, 
    260.3522, 258.363, 259.4599, 260.913, 262.7525, 263.8529, 263.517, 
    263.7181,
  276.0208, 274.7154, 272.647, 268.8574, 264.7274, 261.5854, 260.1239, 
    259.8841, 259.3007, 259.8466, 260.541, 262.399, 263.7126, 264.4538, 
    264.2459,
  276.336, 275.0804, 271.8783, 267.771, 263.5989, 263.6424, 259.9038, 
    259.3161, 259.8558, 260.2026, 260.5179, 262.1296, 263.3557, 264.8025, 
    264.7692,
  276.2958, 274.7961, 268.6644, 263.7905, 264.1859, 261.843, 259.4965, 
    260.1853, 260.7975, 261.3574, 260.6244, 261.1093, 262.7014, 264.2739, 
    266.1928,
  274.2028, 271.8036, 268.1715, 264.7654, 263.8296, 263.9572, 259.9808, 
    263.6527, 262.8519, 259.7837, 258.7492, 260.4033, 262.0036, 263.7052, 
    266.084,
  266.4561, 263.6903, 263.5316, 259.1304, 256.8217, 256.1964, 255.6992, 
    256.5832, 257.1176, 258.2731, 258.3896, 257.4938, 261.1264, 261.6558, 
    260.4976,
  269.8577, 266.5051, 264.8519, 260.5692, 258.7721, 256.8833, 256.5014, 
    257.4395, 258.1725, 258.0072, 256.8766, 258.3768, 259.3255, 259.9591, 
    258.6166,
  273.0758, 272.1792, 270.2165, 262.9545, 259.9817, 257.1015, 258.326, 
    258.1076, 258.2448, 259.0738, 258.4446, 258.7269, 261.1876, 261.5503, 
    261.1173,
  273.7996, 273.2103, 272.548, 267.6256, 262.8508, 260.7581, 257.8915, 
    259.22, 259.6093, 259.8973, 259.587, 259.7084, 261.2458, 261.7147, 
    260.6337,
  274.847, 273.1186, 272.7277, 269.1567, 265.3321, 263.032, 262.6948, 
    257.2541, 256.9512, 261.9893, 261.5236, 260.5399, 261.039, 260.5942, 
    261.1083,
  275.6441, 273.8902, 272.0184, 270.1394, 268.4817, 265.5133, 263.4565, 
    261.7495, 260.5858, 260.5135, 260.6574, 260.7994, 261.6146, 260.2866, 
    261.212,
  276.0604, 274.8609, 272.828, 270.3348, 268.5364, 266.4335, 264.3955, 
    263.4956, 262.7094, 261.9785, 261.8114, 261.1382, 260.5323, 260.9964, 
    262.234,
  276.4178, 275.2261, 272.8334, 270.637, 269.1281, 267.8113, 266.6405, 
    265.2837, 264.4927, 263.9774, 263.0631, 261.0887, 260.0408, 261.775, 
    263.2029,
  276.3911, 274.9021, 271.9648, 270.3473, 269.2841, 268.691, 267.6947, 
    266.8912, 266.1795, 265.4388, 263.798, 261.5365, 260.8476, 261.1989, 
    264.4763,
  274.4162, 272.4772, 272.1696, 271.7711, 270.4003, 269.868, 268.7457, 
    268.9641, 268.173, 265.9432, 262.7835, 260.7303, 259.0099, 260.7282, 
    263.3207,
  269.8727, 268.5649, 267.9281, 266.5438, 265.9112, 263.684, 261.8983, 
    260.1941, 260.9402, 260.4754, 260.8047, 258.1201, 257.7158, 257.2498, 
    254.6543,
  271.5341, 270.4908, 268.8662, 267.0675, 264.8542, 265.1109, 262.4364, 
    262.8596, 263.0436, 261.3319, 261.9402, 260.2869, 259.5766, 258.5959, 
    256.9376,
  273.0973, 272.2392, 271.1962, 267.8636, 268.0918, 265.8503, 266.7121, 
    265.8436, 265.2841, 264.7328, 264.3252, 263.1898, 262.7854, 261.9732, 
    260.7137,
  274.0305, 273.5017, 272.8547, 270.4381, 270.4108, 267.718, 266.2221, 
    267.6121, 266.6548, 266.541, 265.6187, 264.518, 264.3247, 263.9092, 
    262.4887,
  275.272, 273.4773, 273.1245, 271.8449, 271.6366, 271.2803, 270.324, 
    267.0752, 266.6609, 269.0688, 269.3027, 268.5516, 267.5426, 266.2367, 
    264.6087,
  276.007, 274.3227, 272.2825, 271.7551, 272.0305, 272.2816, 272.0238, 
    271.661, 271.3405, 270.9919, 270.1831, 269.2503, 268.7173, 267.8275, 
    266.8737,
  276.1671, 275.018, 273.0276, 271.9352, 272.228, 272.4637, 272.3287, 
    271.7841, 270.5282, 269.1877, 267.9594, 267.6552, 267.9081, 267.6689, 
    267.5416,
  276.5387, 275.3982, 273.2429, 272.2297, 272.5628, 272.3734, 271.3137, 
    269.4334, 267.4341, 266.5861, 266.2515, 266.7782, 266.4589, 266.6982, 
    266.8648,
  276.5015, 275.0326, 272.257, 272.3339, 271.7246, 270.1196, 268.0467, 
    266.3218, 265.832, 266.0918, 263.9911, 264.5287, 264.8301, 265.1568, 
    266.0056,
  274.6008, 272.4524, 272.0253, 271.4086, 269.77, 266.7341, 264.2835, 
    264.8855, 265.8923, 263.5471, 262.5258, 262.7922, 263.244, 263.9996, 
    264.9387,
  270.9253, 270.5065, 271.9164, 270.9489, 270.9445, 270.7528, 270.0503, 
    267.5896, 266.4431, 265.5953, 266.3155, 266.9157, 266.0329, 266.1896, 
    264.7422,
  271.9331, 271.7192, 271.4276, 271.584, 271.895, 271.7949, 270.2732, 
    268.9719, 267.7522, 267.1535, 267.4799, 267.919, 267.8406, 265.9691, 
    264.7925,
  273.3456, 272.5092, 272.0634, 271.3611, 271.9271, 269.7272, 270.098, 
    269.068, 267.6406, 268.0923, 268.488, 269.3552, 269.6833, 269.3674, 
    267.2403,
  274.4014, 273.7803, 273.0589, 270.963, 270.5981, 269.0258, 267.3157, 
    266.2904, 266.5419, 267.5785, 267.48, 268.4877, 268.8654, 268.9314, 
    268.0008,
  275.5062, 273.6254, 273.1808, 269.738, 268.4117, 267.9043, 267.1362, 
    263.4624, 264.3498, 265.1588, 264.4232, 264.0804, 263.9866, 264.1329, 
    265.3847,
  276.13, 274.4628, 272.3086, 269.4733, 267.0543, 265.0099, 265.2602, 
    265.724, 264.9664, 261.5561, 259.5618, 258.9318, 258.7169, 258.2762, 
    260.5711,
  276.2597, 275.0915, 273.061, 269.2642, 264.6833, 262.2605, 261.1669, 
    262.1145, 261.7284, 260.8074, 259.3954, 258.0195, 259.495, 258.6454, 
    258.9049,
  276.5587, 275.423, 272.515, 266.7552, 263.1996, 260.401, 259.2958, 
    259.8438, 260.9807, 261.5216, 261.1758, 261.3332, 261.6049, 262.3866, 
    262.625,
  276.4572, 275.0598, 268.8943, 262.6138, 262.08, 259.617, 259.3647, 
    261.0354, 261.8871, 263.1044, 262.0089, 261.2786, 262.0398, 262.5584, 
    263.3888,
  274.6488, 271.3924, 265.7441, 261.7276, 259.9581, 259.1736, 259.877, 
    261.9281, 264.581, 263.0174, 262.06, 261.285, 261.347, 262.1295, 262.6349,
  269.6098, 267.2549, 265.8859, 265.0887, 264.9182, 265.0069, 262.3267, 
    261.8599, 261.8057, 262.8011, 263.3201, 263.92, 265.0497, 266.9301, 
    268.1846,
  271.03, 269.0084, 264.7434, 263.6618, 264.202, 261.428, 260.1796, 260.2935, 
    260.4298, 260.743, 262.0165, 263.2536, 264.1035, 264.7493, 266.9508,
  273.2937, 272.4319, 269.6185, 261.9285, 260.8518, 258.1308, 259.2657, 
    259.8246, 260.7263, 259.6605, 259.5195, 260.9547, 261.7948, 262.9034, 
    266.1181,
  274.2296, 273.4535, 272.441, 264.5188, 261.4399, 258.9763, 256.6291, 
    257.8973, 259.5027, 260.6846, 259.437, 259.269, 258.9733, 260.9862, 
    263.0801,
  275.3383, 273.3536, 272.8976, 266.0101, 262.5095, 261.9274, 259.5865, 
    255.2617, 258.1665, 261.2965, 260.3644, 259.1129, 258.5021, 257.923, 
    258.5507,
  275.9845, 274.2517, 272.2033, 268.0975, 264.4207, 260.3002, 261.2596, 
    261.8785, 262.0281, 259.9901, 258.5669, 258.8119, 260.0464, 257.9776, 
    257.1875,
  276.2264, 275.0598, 273.0247, 269.275, 264.2771, 259.5628, 260.2867, 
    261.6735, 261.5176, 261.2639, 260.2981, 259.6159, 261.4287, 261.0594, 
    260.0461,
  276.4981, 275.3796, 272.7624, 268.0583, 265.1882, 260.8246, 259.7333, 
    261.6094, 262.0145, 261.6018, 261.4417, 260.8649, 261.578, 263.0412, 
    263.2825,
  276.3736, 275.0536, 270.7118, 265.2556, 265.6958, 261.4448, 260.7157, 
    262.5144, 262.9457, 264.2457, 262.0702, 261.8386, 260.543, 261.3727, 
    263.111,
  274.6648, 272.2844, 269.9437, 266.8659, 266.3659, 263.3453, 260.8845, 
    263.1591, 265.3369, 263.2495, 261.6785, 261.306, 259.6376, 260.9609, 
    262.2558,
  270.1974, 267.5602, 265.9548, 264.2289, 263.745, 264.0562, 261.4032, 259.6, 
    259.1188, 259.5853, 260.499, 256.9057, 258.0073, 260.8028, 262.3888,
  271.4098, 270.1723, 268.3004, 266.4016, 265.7592, 264.2221, 262.9418, 
    261.6569, 260.4185, 259.2197, 258.3453, 255.9025, 256.3632, 260.3447, 
    259.1605,
  273.2987, 272.4475, 271.3328, 268.3561, 266.7898, 264.7089, 263.9614, 
    263.2425, 262.4029, 260.7947, 259.4619, 257.6064, 257.0912, 260.5232, 
    259.3202,
  274.2433, 273.4408, 272.7499, 270.6495, 269.2776, 266.9896, 263.4305, 
    262.8374, 262.508, 261.3975, 260.7985, 258.0229, 257.4337, 260.9445, 
    258.9424,
  275.3916, 273.3957, 273.0349, 271.5221, 270.6405, 269.4526, 267.3129, 
    261.6013, 260.1178, 262.77, 260.8045, 258.2594, 257.9397, 260.932, 
    260.7392,
  276.0151, 274.3625, 272.2856, 271.6753, 271.6738, 270.3537, 268.6582, 
    266.1435, 263.7418, 262.4059, 260.666, 257.9389, 257.8023, 258.1259, 
    262.0804,
  276.2876, 275.1555, 273.139, 271.8995, 272.0364, 270.5778, 269.1029, 
    266.7183, 263.5498, 261.2238, 260.5076, 259.2125, 257.8161, 259.3421, 
    261.4219,
  276.5567, 275.4414, 273.2881, 272.3442, 272.1614, 270.7754, 268.5409, 
    266.2709, 263.3936, 262.0982, 261.218, 259.1313, 258.3589, 260.9554, 
    261.4475,
  276.4352, 275.1185, 272.3918, 272.6656, 271.8818, 269.8889, 268.8719, 
    266.3733, 264.2707, 263.727, 259.3694, 258.2647, 257.6277, 258.9957, 
    263.0751,
  274.7655, 272.6353, 272.3732, 272.2305, 271.1396, 269.5807, 268.5169, 
    266.6411, 265.485, 261.1137, 257.6363, 257.741, 257.0908, 258.0859, 
    262.6339,
  272.1523, 271.6287, 271.4777, 270.5608, 270.1147, 269.9312, 269.7804, 
    269.999, 269.0876, 267.1027, 266.3655, 264.1939, 262.4728, 260.4831, 
    256.4771,
  272.4018, 272.0091, 271.921, 271.6706, 271.1989, 270.6863, 269.9544, 
    269.9766, 269.5648, 268.0387, 266.6731, 264.7352, 262.074, 260.3093, 
    256.8995,
  273.3425, 272.5175, 272.0703, 271.5187, 271.0445, 270.3918, 270.5931, 
    269.291, 268.2653, 266.4808, 265.3161, 264.3144, 261.6154, 261.4086, 
    260.5372,
  274.3496, 273.5178, 272.874, 271.0964, 270.4589, 270.3824, 268.0799, 
    266.8364, 266.1535, 266.2273, 265.0447, 262.7448, 260.8574, 261.0807, 
    260.8249,
  275.5326, 273.5194, 273.133, 270.4698, 269.4457, 269.0678, 267.2264, 
    263.0932, 262.9693, 265.0221, 263.0884, 261.5777, 261.0462, 260.3647, 
    261.7446,
  276.1602, 274.5607, 272.3818, 270.4669, 269.0772, 267.5316, 266.4312, 
    265.3909, 264.1025, 263.313, 261.9937, 260.7484, 260.4492, 259.9546, 
    259.3484,
  276.4449, 275.2501, 273.1839, 270.3569, 268.1302, 266.3639, 264.4115, 
    263.4532, 262.6596, 258.9906, 259.295, 260.3698, 260.2442, 260.1409, 
    259.5583,
  276.6981, 275.5049, 272.863, 268.9397, 266.5988, 265.0292, 264.3437, 
    263.2432, 261.7765, 259.6185, 258.3843, 259.0811, 260.7023, 260.7834, 
    261.3021,
  276.508, 275.1635, 270.4813, 266.744, 264.8945, 264.1686, 263.997, 
    263.5369, 262.4691, 261.3225, 258.2686, 257.8777, 257.7486, 258.7682, 
    261.6939,
  274.8829, 271.9314, 268.5009, 264.9784, 262.7971, 261.3602, 261.2598, 
    262.9247, 262.8396, 258.878, 255.5392, 256.0227, 256.1838, 257.4395, 
    260.1292,
  269.5051, 268.1059, 267.3565, 266.9397, 266.0316, 262.4323, 260.3944, 
    261.361, 262.9755, 264.4471, 265.9392, 266.8486, 267.0934, 267.0272, 
    265.1378,
  271.0931, 269.091, 266.1112, 265.8511, 264.2396, 260.3205, 259.3066, 
    259.9741, 261.0396, 263.3625, 265.22, 268.6173, 268.0582, 265.935, 
    264.3163,
  273.3271, 272.5207, 269.9554, 264.3074, 262.0367, 259.3747, 259.3127, 
    259.5242, 260.5631, 262.426, 264.6282, 267.562, 268.5357, 266.4742, 
    264.3423,
  274.331, 273.4635, 272.529, 264.8364, 261.1385, 260.1491, 256.8887, 
    258.4472, 259.3379, 260.9735, 263.0661, 265.2903, 265.826, 264.7052, 
    264.0735,
  275.5419, 273.4728, 272.9754, 265.6255, 263.0822, 262.393, 261.9702, 
    256.6145, 257.4059, 260.7223, 261.9488, 263.3376, 264.0967, 264.3766, 
    265.1255,
  276.1256, 274.506, 272.316, 268.0687, 264.0393, 262.0141, 262.0501, 
    261.7455, 259.8527, 259.4023, 260.0432, 261.6573, 262.9441, 263.1103, 
    262.6212,
  276.382, 275.1766, 273.0737, 267.7167, 262.8705, 262.1982, 261.6562, 
    261.7761, 261.5649, 258.8212, 259.3755, 260.8793, 260.8922, 261.2673, 
    261.0488,
  276.6285, 275.3931, 272.0586, 265.0505, 262.2982, 261.845, 261.5594, 
    261.4554, 261.6329, 259.2107, 258.3681, 260.1113, 261.2592, 260.9469, 
    261.9716,
  276.3788, 275.0165, 268.712, 263.6773, 262.1866, 261.4532, 261.6602, 
    262.359, 262.4405, 261.6199, 259.4873, 258.7909, 259.308, 260.2032, 
    260.4716,
  274.7679, 271.4593, 267.4296, 264.2202, 262.3181, 260.9695, 261.2511, 
    263.0027, 263.1078, 259.8488, 257.0806, 255.7541, 259.1035, 259.3323, 
    259.5542,
  268.028, 266.6659, 265.758, 264.8412, 263.8542, 259.8628, 257.9849, 
    256.1796, 256.2798, 258.8544, 260.565, 262.6745, 264.0864, 265.7603, 
    265.6105,
  270.771, 269.2477, 266.6789, 265.6491, 262.7686, 259.183, 258.5045, 
    257.408, 256.9409, 257.1967, 260.4981, 263.8016, 265.8886, 265.512, 
    264.5629,
  273.2285, 272.4962, 270.3327, 265.4567, 261.7835, 259.7703, 258.7298, 
    259.3191, 258.1253, 259.0081, 260.9038, 264.7625, 267.8219, 266.5963, 
    266.5073,
  274.2089, 273.417, 272.5163, 266.4609, 262.3689, 259.4349, 255.9573, 
    258.6032, 259.658, 260.5763, 261.1157, 264.2661, 267.4395, 267.7329, 
    267.2565,
  275.3551, 273.3427, 272.9527, 267.1544, 263.5914, 260.4765, 259.116, 
    254.9106, 256.8423, 261.0681, 260.9647, 262.7475, 265.1513, 267.1701, 
    267.3148,
  275.8906, 274.3433, 272.2598, 268.5656, 264.0144, 262.2791, 259.8135, 
    258.9074, 258.532, 259.7544, 260.0228, 261.062, 262.6543, 264.206, 265.478,
  276.1552, 275.0192, 272.9073, 267.7273, 263.9389, 262.7235, 259.9364, 
    260.034, 259.019, 258.9343, 259.8365, 260.6182, 261.588, 262.4317, 
    263.0743,
  276.4403, 275.2474, 271.7517, 266.1157, 263.8492, 262.6984, 260.9828, 
    260.8095, 260.2646, 259.83, 259.091, 259.7057, 261.3448, 262.2174, 
    263.4175,
  276.2156, 274.8855, 269.0988, 265.1841, 263.1546, 261.7012, 261.8171, 
    262.5351, 262.0041, 261.0075, 261.1092, 260.3994, 260.5001, 261.9657, 
    263.2637,
  274.6413, 271.6412, 267.2182, 264.8372, 262.9915, 261.8633, 261.4153, 
    263.7704, 263.7079, 260.7894, 259.5749, 260.4605, 261.0264, 261.5694, 
    262.9966,
  271.4783, 268.1287, 262.7965, 263.9868, 263.1554, 261.5782, 256.8496, 
    257.5137, 257.0859, 259.9352, 260.3451, 260.3897, 262.5233, 265.0368, 
    267.4225,
  271.9494, 269.4334, 264.1994, 263.2518, 262.9188, 259.7314, 257.5251, 
    258.1071, 258.1442, 257.3359, 259.2657, 262.6576, 263.8713, 264.3252, 
    265.4596,
  273.21, 272.563, 269.8335, 262.9477, 261.0205, 259.5255, 258.2751, 
    259.7805, 260.4313, 259.3082, 258.8208, 263.4076, 264.5181, 265.2086, 
    265.4718,
  274.1873, 273.4948, 272.5374, 265.2333, 261.6894, 258.0001, 257.0509, 
    259.9503, 261.0231, 261.6496, 260.722, 262.0511, 263.3761, 264.1001, 
    263.658,
  275.2324, 273.3194, 272.9534, 266.2266, 262.8588, 261.177, 258.2224, 
    256.4277, 257.54, 262.2218, 262.4999, 262.5162, 263.043, 265.1509, 
    267.3752,
  275.7518, 274.2651, 272.2456, 267.7186, 264.1224, 263.0877, 260.8698, 
    260.6413, 260.9499, 261.3937, 262.0377, 263.4374, 263.3935, 262.4393, 
    266.8405,
  276.0443, 274.9311, 272.6459, 266.3681, 263.5759, 263.3376, 262.4766, 
    262.3139, 261.7428, 261.5142, 262.3717, 263.7599, 265.1243, 264.007, 
    264.5121,
  276.3566, 275.1519, 270.9434, 264.294, 263.1133, 263.0827, 263.0107, 
    263.0621, 262.6502, 261.8529, 262.3731, 263.9811, 265.6158, 266.6118, 
    265.552,
  276.1412, 274.8317, 267.9231, 263.543, 262.6761, 262.9754, 263.518, 
    264.1303, 263.3796, 262.9366, 262.8099, 263.8694, 265.762, 267.2462, 
    267.437,
  274.6133, 271.3893, 264.8996, 264.4876, 263.2014, 263.2248, 263.8013, 
    265.7306, 265.0331, 262.9732, 262.5448, 263.5616, 265.3101, 267.3247, 
    268.6712,
  271.4696, 266.7993, 263.4125, 260.4735, 258.193, 257.77, 259.8994, 
    261.0974, 260.9506, 261.9272, 262.2903, 261.4519, 261.8548, 264.9428, 
    268.4324,
  270.7713, 267.0736, 262.5889, 259.7926, 259.369, 258.2012, 261.4723, 
    261.3105, 261.1668, 258.4611, 261.4572, 263.8253, 261.9623, 263.496, 
    266.8607,
  273.0701, 272.401, 268.3355, 262.941, 260.1972, 257.9664, 261.7821, 
    263.3157, 263.6435, 262.4954, 260.4164, 264.5666, 263.2967, 264.1236, 
    267.3006,
  274.0765, 273.3964, 272.3536, 265.328, 262.983, 260.178, 260.3229, 
    263.3932, 264.112, 264.4972, 262.932, 265.5431, 264.863, 261.3011, 
    266.6824,
  275.144, 273.2745, 272.8625, 266.3102, 263.7951, 263.0723, 262.6951, 
    259.3091, 260.7466, 265.1404, 265.2663, 266.8264, 265.9714, 261.1193, 
    265.9534,
  275.6791, 274.2105, 272.2214, 267.4861, 264.401, 263.1364, 262.983, 
    262.7726, 262.8983, 264.2027, 265.6567, 268.042, 267.3279, 264.8899, 
    265.1295,
  275.9918, 274.9279, 272.5992, 266.2591, 264.1157, 263.0954, 262.6894, 
    262.6668, 262.9219, 264.2067, 265.8171, 268.1017, 268.4717, 265.9439, 
    262.8603,
  276.3154, 275.179, 270.7427, 264.88, 264.0987, 263.6399, 262.7816, 
    261.8838, 262.1713, 263.7204, 265.5941, 266.695, 268.7001, 266.3709, 
    265.6323,
  276.1299, 274.7948, 266.9728, 263.9668, 264.2198, 262.5651, 262.2561, 
    262.9548, 262.8721, 264.166, 264.9226, 266.3335, 267.5389, 267.4844, 
    266.2669,
  274.6561, 271.4349, 263.985, 264.8459, 264.2575, 261.1354, 261.8661, 
    265.0412, 264.5537, 262.9551, 263.7319, 264.9743, 266.9847, 269.4731, 
    266.2866,
  267.6889, 265.4979, 262.8187, 259.5331, 258.9016, 257.5718, 259.0409, 
    260.6849, 262.8654, 264.3479, 265.8406, 265.977, 265.0783, 265.3708, 
    265.0965,
  268.4966, 265.2973, 262.4754, 260.9275, 260.5718, 259.5097, 261.2776, 
    263.5266, 264.1745, 261.8396, 266.3795, 267.0039, 266.5627, 264.4444, 
    264.9511,
  272.9338, 272.1741, 267.8148, 263.1199, 261.4907, 259.0813, 262.5807, 
    264.0272, 264.855, 265.7033, 266.2684, 267.4274, 267.0509, 265.5106, 
    266.4871,
  273.9908, 273.3442, 272.0104, 264.2664, 261.968, 261.2291, 260.1473, 
    263.3598, 265.2732, 266.5471, 266.7809, 267.0042, 266.6406, 265.1432, 
    268.125,
  275.0867, 273.2537, 272.6678, 265.6078, 263.3241, 262.3207, 261.1555, 
    260.7399, 262.8376, 267.203, 267.012, 266.7259, 266.3916, 265.8622, 
    268.9469,
  275.6424, 274.2311, 272.1625, 267.077, 263.6447, 262.0585, 261.4558, 
    262.4967, 264.5939, 265.9796, 266.9209, 267.2187, 266.5299, 266.2938, 
    268.6138,
  276.0287, 275.0382, 272.552, 265.907, 263.8153, 262.1466, 262.361, 262.753, 
    264.2497, 265.7147, 266.5656, 267.9231, 266.9526, 266.5347, 267.9124,
  276.3563, 275.3497, 270.0749, 262.7552, 263.6837, 262.4562, 262.7281, 
    262.7386, 263.1528, 264.7963, 265.8856, 267.5252, 267.9726, 267.0819, 
    267.5954,
  276.1853, 274.8603, 267.0324, 262.0805, 261.628, 262.1007, 262.7054, 
    264.8644, 264.9212, 265.7844, 265.0223, 267.0526, 268.3684, 267.8946, 
    266.9802,
  274.7419, 271.9193, 264.4446, 263.538, 261.4478, 261.5509, 261.9868, 
    266.5074, 266.5958, 264.9047, 262.9894, 265.008, 268.2803, 268.889, 
    267.1617,
  265.9352, 264.885, 260.8197, 261.8116, 259.8789, 259.5086, 260.9569, 
    264.8745, 266.2406, 266.0179, 267.5265, 267.473, 266.9507, 266.886, 
    266.3991,
  267.3902, 264.1004, 263.5823, 263.4414, 263.1088, 259.8885, 260.0909, 
    265.1693, 265.8154, 266.6323, 267.7541, 267.7484, 267.3734, 265.8266, 
    265.5318,
  273.0801, 272.26, 268.1657, 264.5055, 262.5232, 260.7003, 260.5763, 
    262.6329, 265.7709, 267.067, 267.8818, 267.9761, 267.5054, 267.2245, 
    266.5968,
  274.1683, 273.3963, 271.9833, 265.0835, 262.8214, 259.7456, 260.418, 
    261.8947, 265.1702, 266.7219, 267.5093, 268.5039, 268.2288, 268.123, 
    268.2792,
  275.2217, 273.4887, 272.6898, 266.5461, 263.7119, 263.1427, 264.1329, 
    261.4425, 262.8503, 267.044, 267.3408, 268.688, 268.4353, 268.5865, 
    269.0891,
  275.6927, 274.5, 272.3213, 267.2824, 264.2249, 263.445, 264.3786, 264.8481, 
    265.1762, 265.8015, 266.8319, 268.588, 268.8216, 268.6556, 269.4568,
  276.0323, 275.2397, 272.7559, 264.4365, 264.4673, 263.6328, 264.3119, 
    264.8475, 265.1744, 265.5746, 266.3743, 268.3701, 268.9461, 268.8948, 
    269.393,
  276.3364, 275.5027, 269.9498, 261.4952, 264.7697, 263.3679, 264.3939, 
    264.9358, 264.9394, 264.9695, 265.6225, 267.8546, 268.8905, 269.099, 
    269.2867,
  276.1885, 274.9609, 267.8936, 261.5996, 262.7845, 263.5123, 264.2685, 
    265.5844, 265.7014, 265.6377, 264.9127, 266.9787, 268.8245, 269.0482, 
    269.3448,
  274.7858, 272.1466, 266.3962, 261.9667, 264.0264, 263.4332, 262.739, 
    267.0561, 266.8182, 264.6313, 263.8057, 265.6083, 268.4757, 269.0343, 
    268.9771,
  265.9851, 266.472, 264.5549, 264.0268, 263.3854, 263.3695, 264.4742, 
    264.9229, 265.1423, 266.1425, 266.4668, 267.7731, 268.5002, 268.4709, 
    268.5283,
  268.7484, 267.5735, 266.2137, 264.6276, 263.6782, 263.8359, 263.5358, 
    261.5053, 261.2948, 265.382, 266.0616, 267.0094, 268.5481, 268.2126, 
    268.6777,
  273.1102, 272.4328, 268.7001, 265.3652, 263.8457, 262.2669, 261.3794, 
    260.6583, 263.1209, 265.5205, 265.4854, 266.8509, 268.2921, 269.1848, 
    269.4328,
  274.0768, 273.5421, 272.102, 266.1142, 264.5405, 263.5346, 261.8224, 
    260.0342, 261.5923, 264.6129, 264.9137, 266.1507, 268.2419, 268.4521, 
    269.0042,
  275.2074, 273.7119, 272.752, 267.0502, 264.5534, 264.4906, 264.6395, 
    260.3174, 261.2818, 264.5934, 264.6399, 266.0887, 268.1861, 268.0993, 
    268.9227,
  275.7106, 274.7584, 272.5411, 267.3983, 264.1589, 264.0444, 264.7148, 
    264.498, 263.2153, 263.3588, 264.093, 266.0651, 268.1575, 268.6272, 
    269.4679,
  276.0203, 275.3816, 272.9072, 265.4131, 264.3009, 263.903, 264.7569, 
    264.3997, 263.7044, 263.3703, 264.1387, 266.0562, 268.3097, 269.0006, 
    268.2497,
  276.3282, 275.6121, 270.9212, 264.4743, 263.9803, 263.6474, 264.6256, 
    264.6408, 263.846, 263.3562, 263.7624, 266.267, 268.1666, 267.6378, 
    268.6803,
  276.2494, 275.0401, 268.5915, 266.6253, 265.0323, 263.3053, 263.878, 
    265.3197, 265.0379, 264.5654, 264.0628, 266.3172, 267.9745, 265.8385, 
    266.6004,
  274.943, 272.4952, 270.0247, 268.133, 266.9393, 262.9637, 262.8952, 
    267.1182, 266.2815, 263.726, 263.4766, 266.1468, 267.0918, 265.3766, 
    266.3591,
  266.0878, 266.9652, 265.8599, 265.2761, 264.8363, 263.5026, 264.703, 
    264.1629, 261.037, 263.7296, 263.8911, 263.9071, 264.3846, 266.1194, 
    265.9503,
  268.1299, 268.6582, 267.5973, 266.2438, 265.3646, 264.3645, 264.1171, 
    259.65, 259.1276, 261.1484, 262.5344, 263.4656, 262.7519, 265.0578, 
    265.3004,
  273.294, 272.4554, 270.1468, 267.8695, 265.0755, 263.8847, 262.4608, 
    262.5647, 260.7649, 264.0856, 261.5309, 263.9857, 264.6962, 266.0276, 
    266.0379,
  274.2226, 273.4975, 272.2813, 268.877, 267.257, 266.0681, 262.9014, 
    261.8741, 261.6951, 262.2955, 263.3483, 263.5416, 264.7176, 266.2274, 
    266.9352,
  275.2611, 273.6862, 272.8485, 269.8291, 267.7642, 266.9699, 265.4835, 
    261.4258, 260.9226, 263.4912, 263.543, 262.9526, 264.8799, 265.4148, 
    265.0898,
  275.7232, 274.7236, 272.5422, 270.1376, 267.7785, 266.7209, 266.7497, 
    265.5487, 264.1141, 263.3677, 263.344, 263.3253, 264.7383, 264.2668, 
    264.9719,
  276.0005, 275.3205, 273.1002, 269.6455, 267.5745, 266.1884, 266.723, 
    266.6931, 265.6562, 263.81, 262.7174, 262.742, 265.4444, 265.0497, 
    265.3271,
  276.2945, 275.5107, 272.0744, 268.8888, 266.8612, 265.9693, 266.3073, 
    267.6841, 266.6554, 264.458, 262.8877, 263.6742, 265.8317, 266.4676, 
    267.4597,
  276.19, 274.8499, 270.2898, 268.2415, 267.6444, 266.6683, 266.2923, 
    267.538, 266.4385, 264.5871, 262.1739, 263.8049, 266.0192, 266.8087, 
    267.8838,
  274.8445, 272.4244, 269.4471, 268.4465, 267.0297, 265.5144, 265.3472, 
    267.6974, 266.0848, 264.6312, 263.0553, 265.7377, 266.0639, 267.7549, 
    268.5748,
  269.027, 267.1266, 267.0247, 266.4413, 266.5377, 266.5615, 264.8747, 
    264.4294, 265.1523, 265.1786, 265.5197, 264.6809, 263.9294, 264.6996, 
    265.7882,
  269.9394, 268.113, 269.1479, 268.6023, 268.3999, 268.3617, 266.5638, 
    265.7433, 264.6785, 264.1452, 263.4711, 263.2673, 261.3029, 263.3143, 
    264.2969,
  273.2441, 272.5256, 270.8027, 269.1957, 269.4117, 267.9137, 269.2457, 
    268.433, 267.2784, 265.885, 264.2276, 263.3907, 261.7024, 263.9764, 
    264.8506,
  274.1443, 273.4016, 272.5301, 269.4092, 267.7433, 268.3305, 266.6024, 
    268.053, 267.4202, 267.5742, 266.8989, 264.916, 262.4088, 263.9249, 
    264.192,
  275.2104, 273.4814, 272.9681, 269.0366, 266.5403, 266.4694, 266.4815, 
    263.498, 261.876, 266.3236, 266.9393, 265.8241, 263.2234, 263.0157, 
    262.3776,
  275.6427, 274.5303, 272.445, 267.6086, 265.4618, 265.171, 265.162, 
    265.3666, 263.8805, 264.0894, 265.8147, 266.2559, 264.3705, 262.1598, 
    262.8284,
  275.9202, 275.1571, 272.4092, 265.5617, 264.8799, 264.6089, 264.4187, 
    265.0418, 265.0556, 264.1787, 266.9161, 266.1798, 264.1657, 262.4758, 
    263.953,
  276.2014, 275.3347, 270.1581, 265.2217, 264.9811, 265.7005, 265.3211, 
    266.3278, 267.5693, 266.1593, 266.7514, 265.4686, 264.2019, 264.3636, 
    265.6627,
  276.0427, 274.6601, 268.2453, 265.4019, 265.7719, 266.5732, 267.0214, 
    267.2705, 266.8523, 265.3125, 266.3134, 264.7878, 263.9326, 265.1577, 
    265.7994,
  274.6943, 272.0785, 267.5938, 266.2057, 266.0983, 266.7067, 267.2534, 
    268.8813, 267.6928, 267.0648, 265.5466, 265.4875, 264.5957, 265.3199, 
    266.2518,
  269.4489, 265.2569, 268.1471, 264.4727, 263.4208, 262.7209, 264.0256, 
    265.8222, 264.745, 263.7023, 264.7202, 265.0408, 263.6896, 264.0993, 
    265.2648,
  270.8424, 268.0491, 268.4863, 267.3737, 267.5227, 267.8258, 267.6867, 
    267.3871, 266.4941, 264.6984, 264.6364, 265.4154, 264.3742, 262.94, 
    264.5643,
  273.3492, 272.6498, 270.6476, 267.5085, 267.1341, 266.5075, 266.4227, 
    265.7945, 267.8838, 267.2892, 265.175, 265.7868, 264.1986, 264.6605, 
    264.9041,
  274.2081, 273.4681, 272.6268, 269.3467, 267.6891, 267.6427, 264.7621, 
    265.0414, 262.5645, 267.5735, 266.0037, 266.5376, 265.7781, 265.1966, 
    264.6599,
  275.24, 273.5273, 273.0512, 270.2582, 267.5251, 267.1124, 266.1407, 
    262.2803, 261.1843, 263.3401, 268.1315, 267.2535, 266.0527, 266.0523, 
    260.7703,
  275.6469, 274.5444, 272.5388, 269.4497, 266.9262, 265.2602, 266.2268, 
    265.2986, 263.2422, 261.655, 267.6552, 268.3003, 266.7401, 263.2075, 
    262.6539,
  275.9051, 275.131, 272.3499, 267.9796, 265.6071, 265.7041, 266.5403, 
    267.4463, 265.8405, 262.1049, 265.3679, 268.5029, 266.8488, 263.2363, 
    265.3297,
  276.1891, 275.2916, 270.3396, 267.0365, 268.055, 267.4232, 267.5024, 
    268.4432, 265.8495, 265.757, 265.1773, 267.6952, 266.2593, 263.6686, 
    266.2512,
  276.0058, 274.5733, 268.7167, 266.8898, 266.7612, 266.2412, 269.4051, 
    269.2053, 266.868, 266.0885, 264.6752, 267.4344, 265.1618, 264.2442, 
    266.2081,
  274.5829, 271.8715, 267.8812, 267.59, 267.5442, 268.6977, 269.1682, 
    268.9185, 266.7501, 265.9442, 265.9725, 267.1462, 263.8532, 264.2299, 
    265.4101,
  270.6638, 268.5655, 269.8188, 269.8256, 268.2213, 265.4424, 266.2448, 
    266.7244, 266.5526, 268.011, 266.7093, 263.7506, 263.6189, 263.2601, 
    265.926,
  270.6129, 269.2926, 268.7251, 269.8061, 270.1979, 269.3672, 267.0266, 
    266.9186, 266.3718, 268.5387, 267.3775, 265.4645, 262.8099, 260.7007, 
    263.5393,
  273.6299, 272.9586, 271.4042, 271.2552, 271.2815, 269.6047, 268.6595, 
    267.973, 266.6434, 268.3918, 266.8051, 265.8178, 264.8555, 262.0302, 
    263.6427,
  274.4342, 273.6646, 272.8761, 269.6446, 269.339, 271.4948, 268.8481, 
    268.6308, 265.7898, 266.9693, 266.6771, 265.3239, 265.6053, 262.0525, 
    262.8098,
  275.3828, 273.7416, 273.2492, 270.0667, 266.9813, 267.6239, 266.0987, 
    265.7102, 263.581, 265.0302, 267.3139, 265.4375, 264.4674, 263.1295, 
    261.7831,
  275.7224, 274.704, 272.9172, 270.4276, 267.5866, 262.584, 267.1401, 
    266.7884, 265.321, 264.8338, 266.9456, 266.1032, 265.9863, 262.3311, 
    263.3857,
  275.9686, 275.2713, 272.4344, 268.7932, 267.8793, 262.6231, 266.651, 
    266.0469, 265.6782, 264.9936, 266.6337, 265.9061, 265.5525, 262.7793, 
    266.8637,
  276.2415, 275.3788, 270.8451, 268.1075, 268.7581, 265.649, 264.5673, 
    266.8313, 265.0021, 265.5121, 266.4567, 266.078, 264.305, 264.7341, 
    268.2462,
  276.0445, 274.5604, 268.4894, 269.0024, 268.5667, 266.5256, 267.3226, 
    267.4321, 266.2485, 265.6863, 265.1386, 265.6165, 263.4591, 267.1392, 
    268.5049,
  274.5568, 271.6647, 267.008, 268.5209, 267.4164, 267.278, 267.4061, 
    268.0737, 266.124, 265.7252, 265.5764, 266.3123, 263.4999, 267.0368, 
    268.5699,
  272.9221, 267.877, 267.4823, 267.8111, 268.8097, 267.8058, 266.3609, 
    268.1106, 267.7713, 269.5461, 267.4031, 263.5233, 265.7729, 267.0743, 
    269.4999,
  271.4517, 269.4409, 267.9539, 270.0539, 270.6339, 268.5485, 268.1581, 
    268.0783, 265.8504, 265.5888, 269.1061, 264.1056, 265.5918, 266.3349, 
    268.9795,
  273.9622, 273.1935, 271.4157, 269.2137, 269.089, 268.3493, 268.7021, 
    268.1528, 265.6997, 266.6655, 267.4261, 264.4278, 266.2431, 266.182, 
    268.3719,
  274.6399, 273.8395, 273.0579, 269.4849, 267.787, 269.0446, 268.4252, 
    269.3797, 265.915, 267.4804, 266.1617, 264.3623, 264.9435, 265.4589, 
    267.2664,
  275.5047, 273.9148, 273.469, 270.0468, 269.2166, 268.9691, 270.0488, 
    266.7235, 265.9366, 266.6954, 265.7986, 266.4614, 265.2254, 265.1115, 
    266.3893,
  275.8059, 274.8563, 273.2699, 269.7749, 267.4436, 264.8679, 269.1909, 
    270.1249, 267.5419, 266.6576, 267.6915, 266.5751, 265.9706, 264.5457, 
    266.463,
  276.0212, 275.431, 272.4353, 270.1275, 267.0606, 265.2237, 268.6883, 
    269.5787, 268.0154, 266.2921, 267.5727, 266.562, 266.5725, 266.1383, 
    267.8199,
  276.2792, 275.5171, 271.314, 266.5129, 267.9331, 265.2817, 265.0943, 
    268.3397, 267.279, 265.3813, 266.2953, 266.2701, 265.2068, 266.5693, 
    268.5743,
  276.0838, 274.5556, 267.3016, 266.3599, 266.3057, 265.4512, 267.4411, 
    268.4511, 267.7339, 265.1056, 266.3445, 265.9539, 264.5012, 267.0351, 
    268.3853,
  274.5694, 271.7184, 267.374, 267.4566, 266.7913, 267.4092, 268.0235, 
    268.5784, 267.0208, 265.5111, 266.1913, 266.0124, 264.4534, 267.299, 
    268.0939,
  273.4731, 268.1487, 267.3972, 269.6488, 268.9683, 269.1721, 270.0068, 
    270.6644, 270.7656, 270.3799, 269.3828, 267.6674, 267.2619, 267.0279, 
    268.6591,
  271.1006, 269.3916, 268.3063, 268.7599, 271.8575, 271.6331, 270.9995, 
    270.6165, 269.5974, 268.1322, 269.8849, 267.426, 266.7699, 267.4848, 
    269.892,
  274.5657, 273.5961, 271.8085, 268.179, 271.4786, 268.6595, 268.6287, 
    267.3809, 269.6393, 267.8876, 269.1332, 266.9082, 266.4498, 268.1242, 
    271.3295,
  274.8933, 273.9949, 273.2122, 270.3311, 266.9455, 268.5154, 270.116, 
    266.3372, 268.0435, 265.1484, 263.1735, 263.7421, 267.5229, 269.8027, 
    271.4174,
  275.5854, 274.0267, 273.6472, 270.6031, 269.7424, 270.6123, 270.4946, 
    264.9835, 262.8425, 267.4494, 265.0206, 266.5862, 269.4066, 270.4836, 
    270.5422,
  275.869, 275.0226, 273.7133, 269.1425, 270.4141, 269.3468, 268.459, 
    266.2868, 266.432, 266.3555, 267.4465, 268.4417, 270.0555, 270.4699, 
    270.5209,
  276.1021, 275.6511, 272.6648, 268.246, 268.8544, 269.3573, 270.4591, 
    266.8658, 266.5529, 266.776, 268.4394, 269.4614, 269.8225, 270.1223, 
    269.9571,
  276.39, 275.7343, 271.1808, 264.5091, 268.9099, 267.808, 269.2736, 
    268.4235, 266.5366, 267.2351, 268.8649, 269.4948, 269.5745, 269.4264, 
    269.2157,
  276.2007, 274.6503, 268.3327, 268.2819, 268.7418, 267.8437, 269.1478, 
    268.2152, 267.0836, 266.8839, 268.2402, 268.9331, 268.8831, 268.9276, 
    268.5653,
  274.6642, 271.7563, 267.0447, 267.9838, 268.4926, 268.5821, 268.6456, 
    268.2563, 267.1022, 267.3036, 267.8028, 268.1047, 268.3476, 268.1669, 
    268.1615,
  272.6473, 270.232, 268.8002, 271.177, 270.1617, 270.7248, 271.2828, 
    271.3394, 270.637, 270.5875, 270.2822, 270.7537, 270.4771, 270.0037, 
    269.3128,
  272.1346, 269.3157, 268.706, 270.6793, 271.1613, 271.6906, 271.4935, 
    270.8832, 269.9333, 270.4035, 269.4164, 270.9996, 270.7712, 269.6713, 
    269.2214,
  274.4532, 273.9581, 272.2756, 270.0095, 270.4467, 267.6527, 267.1029, 
    267.9774, 268.5237, 268.0404, 268.6517, 270.5034, 269.1752, 267.6377, 
    267.2145,
  275.3692, 274.4745, 273.4796, 270.0052, 265.3225, 266.9691, 266.6849, 
    265.3246, 268.1259, 269.8515, 269.0458, 268.454, 266.619, 266.7353, 
    267.7269,
  275.9023, 274.2761, 273.9803, 270.5222, 264.6571, 269.2817, 268.8394, 
    266.218, 264.4141, 265.632, 266.9968, 266.2204, 266.0435, 266.264, 
    269.9039,
  276.0576, 275.3156, 274.233, 269.1822, 266.718, 267.6759, 267.8882, 
    265.7199, 267.0527, 264.1212, 264.3336, 265.9418, 267.1639, 269.6585, 
    270.2956,
  276.313, 276.0401, 273.0672, 267.9919, 267.0029, 267.2992, 267.8776, 
    264.8752, 267.8618, 268.6632, 269.1774, 269.9811, 270.1019, 270.3398, 
    269.8647,
  276.6882, 275.9587, 270.7992, 266.5908, 267.6351, 267.7262, 267.2949, 
    266.33, 266.2534, 269.4848, 269.9368, 270.0414, 270.1089, 269.3933, 
    268.9639,
  276.4058, 274.653, 268.286, 268.9464, 268.965, 268.6227, 268.1424, 
    267.7723, 268.3616, 270.1459, 270.0925, 269.0177, 268.9739, 268.7476, 
    269.1761,
  274.7991, 271.9609, 268.3804, 268.6206, 268.3787, 268.4066, 268.3177, 
    268.5802, 269.8524, 269.7111, 269.3554, 268.6, 268.6688, 269.0477, 
    269.7583,
  274.4339, 272.1394, 271.68, 271.4691, 270.962, 269.8457, 268.9516, 
    268.5057, 267.5307, 268.4105, 270.6135, 268.33, 268.2534, 269.0453, 
    270.0334,
  272.3277, 270.8148, 270.5168, 271.3683, 270.8246, 271.4018, 269.3964, 
    268.3405, 267.1782, 267.6859, 269.5643, 268.7959, 267.2201, 269.5142, 
    267.9661,
  274.1299, 273.8724, 272.6491, 270.8758, 270.5477, 267.4453, 266.7316, 
    266.3992, 265.9341, 266.5083, 266.9558, 268.6107, 267.5745, 266.3505, 
    268.082,
  275.1544, 274.4158, 273.6088, 271.5437, 268.464, 268.0702, 264.379, 
    263.8116, 263.5464, 267.3777, 269.3415, 268.8735, 268.9823, 268.2769, 
    268.3715,
  275.8847, 274.4927, 274.2518, 271.4622, 266.0967, 266.4146, 265.4852, 
    264.7472, 262.2778, 266.4828, 269.0989, 269.2877, 270.0872, 267.3518, 
    267.1282,
  276.2243, 275.5777, 274.3176, 269.501, 265.572, 266.4094, 266.9859, 
    265.9974, 265.2463, 264.7664, 265.3293, 266.1313, 267.6996, 268.466, 
    269.6288,
  276.5531, 276.1909, 272.507, 267.0213, 265.9757, 267.1717, 267.1117, 
    266.529, 268.387, 266.7154, 269.547, 269.5259, 269.4589, 268.9221, 
    269.8483,
  276.899, 276.0442, 269.5274, 265.8671, 266.9332, 267.1381, 265.7169, 
    266.7844, 263.9851, 265.104, 267.1664, 268.8856, 269.659, 269.6458, 
    269.763,
  276.5717, 274.6494, 267.8175, 267.1764, 268.472, 265.8087, 264.6033, 
    264.6275, 268.362, 268.1854, 265.2947, 267.8985, 269.4174, 269.6028, 
    269.718,
  274.8551, 271.8864, 267.9578, 268.6208, 267.187, 268.8713, 267.3215, 
    268.1926, 269.4051, 269.1695, 266.7812, 269.5479, 269.6132, 269.5696, 
    269.9175,
  277.8656, 272.8303, 272.89, 272.9839, 273.0418, 272.691, 272.1966, 
    271.6826, 271.0173, 270.8149, 271.1079, 270.4245, 270.6152, 270.0578, 
    270.3928,
  272.7811, 272.8274, 272.9152, 273.0723, 272.9742, 272.4456, 271.8974, 
    271.5485, 270.9491, 269.8548, 270.2163, 269.4138, 268.5699, 269.7602, 
    268.8499,
  273.8852, 273.439, 272.8838, 272.8058, 272.4842, 271.6419, 270.5131, 
    269.894, 269.597, 268.5269, 268.139, 267.9932, 267.9578, 266.5793, 268.464,
  274.8787, 274.111, 273.3336, 272.5545, 271.8828, 271.0042, 267.3845, 
    267.8862, 267.815, 267.3771, 267.4724, 266.5267, 269.7398, 270.368, 
    267.4349,
  275.6814, 274.0036, 273.5945, 271.8785, 269.9375, 268.6939, 267.8434, 
    265.9618, 264.8687, 267.2596, 266.4984, 267.5964, 268.9157, 269.8187, 
    270.1369,
  275.6996, 274.7312, 273.173, 270.3527, 268.5087, 267.3436, 266.3906, 
    266.4072, 266.6837, 265.4058, 265.3401, 264.5211, 269.4492, 269.7728, 
    269.3949,
  276.0081, 275.4105, 272.4195, 268.0346, 266.8408, 266.3272, 265.6366, 
    265.6507, 267.7355, 268.439, 269.1674, 267.6862, 268.6392, 269.1161, 
    269.1693,
  276.416, 275.7113, 270.3046, 266.782, 266.2291, 268.4746, 266.3022, 
    267.6482, 267.0696, 268.3069, 267.3934, 267.0586, 268.062, 269.732, 
    270.1526,
  276.3662, 274.6511, 268.6423, 267.607, 269.2767, 267.0476, 266.7238, 
    267.7598, 268.4757, 268.7751, 267.2112, 269.2377, 269.651, 269.9272, 
    270.2083,
  274.8631, 272.1831, 269.2994, 269.4275, 268.2194, 268.696, 268.5045, 
    268.6829, 268.7461, 269.1656, 267.4014, 269.0327, 269.3639, 269.3569, 
    269.9317,
  275.5893, 271.8321, 271.5572, 272.0122, 272.2462, 272.3168, 272.3054, 
    272.4585, 272.6675, 272.837, 272.9664, 272.9773, 273.0798, 272.785, 
    272.4225,
  272.4711, 272.121, 272.0113, 272.1887, 272.4698, 272.5488, 272.5502, 
    272.6473, 272.7574, 272.8967, 272.9857, 272.9984, 272.7923, 272.3509, 
    271.8189,
  273.7861, 273.3622, 272.6157, 272.1126, 272.4621, 272.4096, 272.3235, 
    271.449, 271.6229, 272.0627, 272.3517, 272.4957, 272.1996, 271.7953, 
    271.375,
  274.821, 274.0681, 273.3397, 272.1519, 271.502, 271.4738, 268.9185, 
    269.0903, 269.5712, 270.4318, 270.8996, 271.2606, 271.2558, 270.7787, 
    270.4042,
  275.5162, 273.8838, 273.4938, 270.406, 269.1204, 268.9252, 269.0441, 
    266.5298, 265.4501, 269.413, 269.6456, 269.7326, 269.9092, 269.9792, 
    270.0497,
  275.5381, 274.3419, 272.5472, 268.5449, 267.1972, 266.8246, 266.8403, 
    268.0059, 268.5621, 268.7495, 268.9378, 268.8768, 269.056, 269.2071, 
    269.2274,
  275.8123, 274.9837, 271.3886, 266.9377, 266.2051, 265.7568, 265.4357, 
    265.6228, 266.502, 268.1898, 268.5648, 268.4823, 268.5316, 268.5434, 
    268.5766,
  276.2377, 275.4029, 269.8911, 267.5688, 266.5166, 266.4653, 265.7935, 
    265.6398, 265.5619, 266.3442, 267.4659, 267.7416, 268.0506, 268.3695, 
    268.3607,
  276.2261, 274.5503, 269.0369, 268.3045, 267.9481, 267.834, 266.5588, 
    266.8072, 266.6967, 266.4478, 266.7031, 267.2795, 267.5851, 267.6299, 
    269.5934,
  274.8497, 272.47, 269.4732, 268.7723, 267.9708, 267.9772, 268.1444, 266.61, 
    266.632, 266.7685, 267.1041, 267.8816, 268.0633, 268.8677, 269.8582,
  275.1505, 272.2234, 271.5662, 270.4087, 271.3055, 270.941, 270.7544, 
    266.7937, 266.4386, 267.3123, 269.3043, 270.0685, 270.8922, 271.4802, 
    272.1526,
  272.4484, 271.9355, 271.299, 270.0883, 270.4642, 271.2475, 270.3102, 
    265.8422, 265.6718, 266.347, 268.4371, 270.1438, 270.4912, 271.2237, 
    272.1786,
  273.6659, 273.2979, 272.5398, 269.9136, 269.1084, 269.7325, 269.9647, 
    265.0145, 264.998, 265.816, 267.2059, 269.2965, 270.8048, 271.7087, 
    272.4626,
  274.7532, 274.0355, 273.3506, 270.8522, 267.6688, 269.0504, 266.6783, 
    264.8118, 265.028, 266.0605, 266.7236, 268.5218, 270.7477, 271.9237, 
    272.4912,
  275.4332, 273.8318, 273.4971, 269.2151, 266.4536, 265.1775, 269.7617, 
    265.645, 265.183, 266.9105, 266.9958, 268.0268, 270.4883, 271.9358, 
    272.6301,
  275.5296, 274.2998, 272.5528, 267.5771, 265.3777, 264.6291, 269.5013, 
    269.4568, 268.9615, 267.6675, 266.3625, 268.4978, 269.8728, 270.9886, 
    271.9796,
  275.8187, 274.9866, 271.8236, 268.4653, 265.439, 265.6949, 264.4511, 
    268.1559, 267.753, 266.4417, 265.5403, 268.4888, 269.5587, 270.1146, 
    270.7583,
  276.2529, 275.4455, 270.8577, 269.1948, 268.0547, 267.4534, 264.4361, 
    264.5682, 267.0166, 264.6558, 266.1269, 268.6241, 269.6069, 269.927, 
    270.1992,
  276.3358, 274.6036, 269.8661, 269.0381, 268.4709, 268.2362, 265.4065, 
    264.857, 264.5726, 264.5085, 265.7734, 268.88, 269.7539, 270.1382, 
    270.4075,
  274.9014, 272.6025, 269.9039, 269.2976, 268.9356, 266.2763, 266.692, 
    265.355, 264.4954, 264.9313, 266.8832, 269.2698, 270.1127, 270.3943, 
    270.6928,
  273.762, 271.5305, 271.2699, 271.8176, 271.9525, 271.8871, 271.8578, 
    271.0617, 269.9031, 269.9068, 269.8172, 268.6317, 267.7192, 266.0183, 
    265.0982,
  272.1912, 271.7954, 271.6451, 271.6977, 272.0429, 271.9491, 271.5884, 
    269.903, 268.7236, 268.4675, 269.0451, 267.8057, 265.0626, 264.2186, 
    264.7812,
  273.5456, 273.1957, 272.5397, 271.3954, 271.4949, 270.4321, 270.1658, 
    268.6023, 267.9025, 267.3172, 267.2219, 266.7988, 264.6609, 264.6769, 
    267.7532,
  274.6894, 273.9798, 273.2523, 271.397, 270.2062, 269.9834, 266.9648, 
    267.9521, 267.5594, 266.9604, 266.0739, 264.5042, 264.7688, 268.1364, 
    270.2362,
  275.2002, 273.6436, 273.2956, 269.5797, 268.7982, 268.5663, 269.2522, 
    265.463, 265.2094, 266.8381, 264.9402, 263.8223, 267.028, 270.4048, 
    272.167,
  275.4449, 274.1661, 272.2422, 268.2664, 267.5356, 267.6837, 268.4409, 
    268.881, 268.1951, 268.6669, 267.5353, 266.74, 269.728, 271.5522, 272.7938,
  275.8504, 274.9544, 271.1903, 267.3621, 267.4731, 267.811, 267.4293, 
    267.6843, 268.3787, 268.5569, 264.9007, 269.3815, 270.8946, 271.9558, 
    272.7876,
  276.3896, 275.4053, 269.8579, 268.3763, 268.2954, 268.1841, 266.6398, 
    264.7443, 268.5661, 264.4819, 266.9087, 270.7022, 271.176, 271.2412, 
    271.6643,
  276.5786, 274.5882, 269.5614, 269.4304, 269.6003, 269.5045, 269.0498, 
    263.9268, 263.9753, 266.0303, 269.5542, 271.2842, 270.844, 270.8749, 
    271.0834,
  275.0961, 272.7882, 270.6124, 269.3846, 270.112, 263.8595, 264.0766, 
    264.7361, 264.4154, 268.0384, 270.1413, 271.1196, 270.2555, 270.389, 
    270.5244,
  276.5512, 272.1715, 271.5729, 269.5234, 267.5974, 267.2228, 267.8537, 
    269.2151, 270.6751, 271.5167, 271.9098, 270.8034, 269.8889, 269.2818, 
    269.8195,
  272.4972, 272.0956, 271.4135, 268.9095, 266.8508, 267.0207, 267.4083, 
    268.2339, 269.6221, 270.1749, 270.0099, 269.331, 268.8456, 268.0186, 
    268.1021,
  273.5631, 273.3004, 272.5722, 268.2912, 266.104, 266.7851, 266.9005, 
    267.3434, 267.9495, 268.4698, 268.088, 267.8439, 267.1292, 266.8252, 
    268.0637,
  274.6907, 274.0492, 273.3475, 269.4129, 266.307, 268.2648, 266.7614, 
    267.0693, 267.1999, 267.9817, 268.4915, 268.0585, 267.4772, 267.8209, 
    270.853,
  275.3121, 273.6663, 273.4922, 268.0374, 266.608, 268.4642, 269.1729, 
    264.9891, 264.5889, 268.6315, 269.097, 269.7816, 270.9787, 271.9656, 
    272.3401,
  275.8661, 274.2515, 272.5975, 269.8765, 268.7792, 268.21, 267.8275, 
    268.5118, 268.4276, 269.6013, 270.1952, 271.0052, 272.24, 272.4796, 
    272.4789,
  276.4026, 275.0954, 272.5062, 270.3637, 269.7987, 269.1871, 268.4157, 
    268.2054, 268.5651, 269.7479, 270.6083, 271.7834, 272.5621, 272.6642, 
    272.7155,
  276.6949, 275.544, 272.1703, 271.0489, 270.5502, 270.0022, 269.1448, 
    268.6662, 268.5625, 268.9802, 270.9115, 271.873, 272.5521, 272.7444, 
    272.6251,
  276.6805, 274.7268, 270.7006, 270.4897, 270.9471, 270.4856, 269.8089, 
    265.8671, 267.6941, 269.9864, 270.8708, 271.3343, 271.663, 271.6545, 
    271.6708,
  275.1983, 272.909, 270.5266, 269.2862, 270.0642, 269.666, 267.9685, 
    265.9159, 269.2648, 270.5777, 270.5334, 270.5213, 270.5316, 270.899, 
    271.1752,
  278.927, 272.8116, 272.7104, 271.0758, 268.1495, 265.0035, 262.3561, 
    264.3937, 269.1754, 270.9044, 271.8872, 272.0394, 271.8209, 271.6017, 
    271.8227,
  273.0515, 272.7296, 272.139, 270.2454, 268.1453, 264.9627, 262.3462, 
    264.4752, 267.3019, 270.968, 272.0481, 272.0872, 271.4164, 271.2793, 
    271.9814,
  274.109, 273.7713, 272.7294, 269.4062, 266.581, 264.9511, 263.3729, 
    264.2441, 266.9268, 270.6189, 271.8304, 272.3534, 272.1276, 271.9911, 
    272.1153,
  275.1367, 274.5688, 273.3708, 270.821, 264.8977, 267.031, 265.8045, 
    264.7083, 266.6883, 269.6341, 271.4214, 272.326, 272.3564, 272.2473, 
    272.0433,
  275.7537, 274.2461, 273.5739, 269.8896, 266.9943, 269.1828, 269.773, 
    265.5474, 265.1526, 269.3229, 271.148, 272.091, 272.2128, 271.9621, 
    271.8864,
  276.3818, 274.7505, 273.0456, 271.0264, 269.7906, 269.3942, 269.5671, 
    269.5847, 267.846, 269.7581, 271.1459, 272.0304, 271.8391, 271.3733, 
    271.5179,
  276.8919, 275.3756, 273.0018, 271.8182, 270.8156, 270.4456, 270.3979, 
    270.0469, 267.2477, 269.6995, 270.7205, 271.567, 271.4698, 271.2706, 
    271.3098,
  277.1143, 275.8942, 271.5266, 271.1609, 270.2186, 271.885, 271.3875, 
    270.1624, 269.2777, 269.4495, 270.4487, 271.1289, 271.1994, 270.9227, 
    271.0659,
  276.867, 274.8521, 269.9768, 269.805, 271.6829, 271.7041, 270.7324, 
    267.4147, 269.2628, 269.4674, 270.3926, 270.8857, 270.9721, 270.8238, 
    271.2493,
  275.3699, 273.0612, 270.2385, 269.7219, 269.6066, 270.5213, 269.5112, 
    267.3339, 269.6216, 269.9421, 270.5972, 270.7669, 270.9951, 271.0727, 
    271.3567,
  275.3833, 272.3206, 271.3403, 269.0782, 266.6301, 264.7541, 262.8832, 
    263.1219, 266.1242, 270.0351, 271.4331, 271.7574, 271.7838, 271.7358, 
    271.5295,
  272.8431, 272.453, 271.487, 268.7591, 267.4744, 265.1384, 263.2982, 
    264.0806, 264.1912, 269.7346, 270.8028, 271.4578, 271.8766, 270.9266, 
    270.7777,
  273.8986, 273.5408, 272.7378, 269.2107, 267.7163, 265.9895, 265.7228, 
    268.2157, 265.0523, 269.5168, 270.5897, 271.4443, 271.8142, 271.2961, 
    271.3374,
  274.9657, 274.3672, 273.4338, 270.5984, 266.1196, 268.2334, 267.8021, 
    266.859, 266.3434, 269.408, 270.6033, 271.2486, 271.7665, 271.6777, 
    271.6759,
  275.5002, 274.0798, 273.6761, 271.041, 267.4668, 270.0043, 270.6091, 
    266.9914, 265.7662, 269.3344, 270.4952, 271.171, 271.9427, 271.9797, 
    272.1283,
  275.9968, 274.6931, 273.1505, 271.6095, 271.4576, 270.8253, 269.1385, 
    269.8135, 268.9324, 269.9105, 270.9362, 271.4192, 272.128, 272.1892, 
    272.3571,
  276.4839, 275.3339, 272.4948, 269.6249, 269.5814, 270.4591, 270.5129, 
    269.956, 268.6684, 270.068, 270.2363, 271.0722, 272.1338, 272.2655, 
    272.3932,
  276.9158, 275.8029, 271.2945, 269.9065, 269.9247, 269.6691, 269.4481, 
    269.1246, 270.1285, 269.9684, 270.9434, 271.5443, 272.2038, 272.3597, 
    272.4257,
  276.7469, 274.7768, 270.7913, 270.05, 269.7533, 269.3943, 268.637, 
    269.2438, 270.3038, 270.4142, 271.0215, 271.6631, 272.306, 272.4198, 
    272.1785,
  275.3684, 273.2361, 270.939, 269.9786, 269.3785, 268.3658, 268.6353, 
    269.7092, 270.275, 270.6971, 271.2189, 271.9981, 272.4346, 272.5326, 
    272.2263,
  273.7144, 271.0298, 269.6036, 267.8382, 268.5753, 267.4148, 266.7014, 
    267.0469, 268.8743, 270.241, 271.2254, 272.0122, 272.2278, 272.1431, 
    272.2593,
  272.2625, 271.8749, 271.1211, 269.5236, 269.8896, 269.6927, 268.3398, 
    268.9199, 268.2212, 270.2498, 271.2013, 271.95, 271.9478, 271.7224, 
    271.9041,
  273.7815, 273.4599, 272.7976, 270.1497, 269.1106, 268.2764, 269.7012, 
    269.8997, 269.7715, 270.315, 271.0903, 271.7264, 271.9709, 271.6924, 
    271.8185,
  274.8811, 274.3274, 273.4699, 271.3036, 269.2344, 269.8163, 267.8147, 
    268.2304, 269.3271, 270.2125, 270.4994, 271.5726, 271.4542, 271.6265, 
    271.9681,
  275.4123, 274.0129, 273.7428, 270.2868, 269.131, 269.3332, 270.0277, 
    266.6031, 266.3297, 270.3292, 270.7358, 271.2619, 271.616, 272.0668, 
    272.1635,
  275.7862, 274.5873, 273.1523, 269.7998, 269.3148, 269.4463, 269.5557, 
    269.4028, 269.731, 270.4582, 271.4642, 271.2358, 271.8497, 272.2334, 
    272.4591,
  276.1872, 275.2466, 272.17, 269.3525, 269.3346, 269.4789, 269.4449, 
    269.5028, 269.8919, 270.6342, 271.0081, 271.7663, 272.2661, 272.4982, 
    272.5532,
  276.6614, 275.6668, 271.0373, 269.6252, 269.5198, 269.3463, 269.3189, 
    269.4396, 270.1044, 270.4665, 271.0621, 271.9464, 272.366, 272.4883, 
    272.4187,
  276.575, 274.7312, 270.1038, 269.7024, 269.5532, 269.2429, 268.8631, 
    269.3409, 270.1456, 270.6302, 270.8801, 271.9844, 272.4412, 272.3327, 
    272.1308,
  275.3669, 273.2621, 270.9169, 269.9096, 269.4939, 268.9758, 268.9175, 
    269.5233, 270.215, 270.4886, 271.0621, 271.8967, 272.2929, 272.4593, 
    272.2092,
  273.3308, 271.487, 270.5279, 269.6464, 270.2054, 270.045, 269.3924, 
    269.4818, 269.9434, 270.2455, 270.771, 270.8609, 271.4082, 271.985, 
    272.0325,
  272.1537, 271.9752, 271.4077, 270.2057, 270.3762, 270.2957, 269.5151, 
    269.5545, 270.2301, 270.4509, 270.6439, 271.0532, 271.4648, 271.3586, 
    272.0831,
  273.819, 273.5212, 272.8695, 270.6857, 269.727, 267.977, 269.3131, 
    269.8872, 269.9229, 270.1701, 270.5473, 271.2096, 271.7362, 272.0247, 
    272.4285,
  274.912, 274.4008, 273.513, 271.2032, 269.1872, 269.6835, 267.5082, 
    269.0685, 269.4438, 270.211, 270.3931, 271.7437, 272.2156, 272.2602, 
    272.6761,
  275.5275, 274.1454, 273.7714, 270.155, 269.366, 268.9596, 269.5091, 
    265.8454, 266.2209, 270.2259, 270.9342, 272.1339, 272.3896, 272.3279, 
    272.4705,
  275.8692, 274.6662, 273.1161, 269.6966, 269.4583, 269.0003, 268.7694, 
    268.9815, 269.4395, 270.1195, 271.8403, 272.6375, 272.6569, 272.3318, 
    272.2664,
  276.2604, 275.3228, 272.2017, 269.4066, 269.541, 269.0797, 268.5882, 
    269.1415, 269.9712, 270.7151, 272.175, 272.7792, 272.4824, 272.3796, 
    272.3005,
  276.7117, 275.6948, 271.1494, 269.8669, 269.563, 269.0505, 268.9032, 
    269.5211, 270.4821, 271.2383, 272.3691, 272.7385, 272.5884, 272.3536, 
    271.9713,
  276.6557, 274.6809, 270.915, 270.136, 269.4811, 269.1004, 269.3184, 
    270.0352, 270.6825, 271.5418, 272.3676, 272.7133, 272.6323, 272.3444, 
    271.9878,
  275.4164, 273.3827, 271.4815, 270.4404, 269.5462, 269.1598, 269.5481, 
    270.5272, 271.1843, 272.1785, 272.6064, 272.7635, 272.6631, 272.5354, 
    272.022,
  273.5918, 271.7981, 271.2368, 270.2858, 269.3383, 270.2611, 269.4415, 
    269.9101, 270.4402, 270.8337, 271.4204, 271.8644, 272.3478, 272.5089, 
    272.7188,
  272.2839, 272.1509, 271.8029, 270.6485, 270.6492, 270.4213, 269.6626, 
    269.1962, 269.3944, 270.6344, 271.1501, 271.7079, 271.9324, 272.0403, 
    272.5643,
  274.1119, 273.7001, 272.9109, 271.0956, 270.3653, 268.5046, 269.8594, 
    269.7796, 269.8728, 270.3611, 270.9614, 271.3737, 271.7244, 272.0738, 
    272.5176,
  275.1376, 274.5998, 273.5279, 271.7332, 270.2946, 270.1516, 268.2752, 
    270.3208, 270.3233, 270.2581, 270.5764, 271.0091, 271.644, 272.0106, 
    272.2392,
  275.7815, 274.2678, 273.7472, 271.2972, 270.4469, 270.4388, 270.5818, 
    267.3527, 267.5096, 270.961, 270.7129, 270.6855, 271.507, 271.8939, 
    272.3008,
  276.1597, 274.7252, 273.0523, 271.3425, 270.7645, 270.7014, 270.9983, 
    270.9943, 270.9917, 270.9275, 271.0586, 271.0316, 271.4124, 271.8627, 
    272.164,
  276.4036, 275.334, 272.6505, 271.254, 271.1017, 271.4003, 271.4066, 
    271.4681, 271.3019, 271.4446, 271.5077, 271.4564, 271.7267, 271.9247, 
    272.0721,
  276.7382, 275.6374, 272.0694, 271.2808, 271.2799, 271.7096, 271.6335, 
    271.6497, 271.4974, 271.6255, 271.7952, 272.0478, 271.8627, 271.8974, 
    272.0743,
  276.6384, 274.5873, 271.7231, 271.7765, 271.5466, 271.9051, 271.7246, 
    271.7398, 271.6376, 271.7249, 272.4535, 272.6836, 271.0881, 271.3143, 
    272.1602,
  275.3812, 273.3088, 271.9477, 271.8173, 271.369, 271.9941, 271.8873, 
    271.8426, 271.9343, 272.2762, 272.7239, 272.8661, 272.6469, 272.2613, 
    272.282,
  274.7122, 271.7315, 271.6263, 271.4357, 271.3569, 271.4718, 271.3738, 
    271.5663, 271.5238, 271.9127, 272.25, 271.4272, 272.0383, 272.1853, 
    272.391,
  272.297, 272.4356, 272.0596, 271.5904, 271.8047, 271.7503, 271.6432, 
    271.7302, 271.8127, 272.0122, 272.4442, 272.0048, 271.5378, 271.4138, 
    272.3882,
  274.3512, 273.8821, 272.9392, 271.8701, 271.8521, 270.253, 271.7299, 
    271.6983, 272.1945, 271.9517, 272.0514, 272.1605, 271.7773, 271.4384, 
    272.2021,
  275.4589, 274.6691, 273.537, 272.2429, 271.8202, 272.2137, 270.5879, 
    271.2826, 272.1501, 272.1926, 272.1532, 272.2932, 271.9014, 271.3117, 
    271.7074,
  275.9272, 274.3089, 273.7394, 271.9931, 271.9054, 272.2025, 272.084, 
    269.7947, 269.5282, 272.2159, 272.3795, 272.2236, 271.9036, 271.2705, 
    271.356,
  276.3037, 274.7787, 273.0155, 271.821, 272.0901, 272.5052, 272.5758, 
    272.6023, 272.7373, 272.6843, 272.8665, 272.1999, 272.0653, 271.4436, 
    271.4514,
  276.46, 275.3594, 272.5444, 272.0232, 272.3142, 272.5957, 272.6, 272.5552, 
    272.6457, 272.6266, 272.9109, 272.2036, 272.1649, 271.3109, 271.2212,
  276.7669, 275.586, 272.164, 272.1334, 272.3317, 272.4658, 272.4929, 
    272.5411, 272.6205, 272.7834, 272.8757, 272.8203, 272.1086, 271.266, 
    271.2532,
  276.6749, 274.5862, 272.0718, 272.2994, 272.4413, 272.5751, 272.4338, 
    272.2388, 272.2019, 272.2777, 272.4577, 272.7386, 272.0263, 271.2483, 
    271.5434,
  275.4984, 273.4508, 272.27, 272.3134, 272.4707, 272.5727, 272.5603, 
    272.1315, 272.187, 272.6108, 272.7775, 272.7505, 272.1582, 271.1736, 
    271.5721,
  274.4668, 271.9319, 271.9815, 271.8844, 271.8225, 272.0663, 271.8944, 
    271.9319, 271.7784, 272.1227, 272.7431, 272.0119, 272.2377, 270.0109, 
    271.0262,
  272.2483, 272.5574, 272.3236, 271.4666, 272.2567, 272.3631, 272.1391, 
    271.8692, 271.9373, 272.1653, 271.6108, 271.0013, 272.0526, 272.013, 
    271.4776,
  274.3677, 273.9583, 272.9971, 272.0935, 272.4992, 270.9192, 271.9911, 
    271.7021, 271.5429, 272.2046, 271.2195, 272.3347, 272.1592, 272.2355, 
    272.2296,
  275.4656, 274.697, 273.5617, 272.4029, 272.3747, 272.6295, 271.0738, 
    271.8503, 271.1947, 271.9982, 271.9283, 272.4565, 271.8269, 271.2751, 
    270.7661,
  276.0187, 274.3875, 273.7568, 272.1609, 272.5348, 272.8335, 272.8633, 
    270.0983, 269.8134, 271.7498, 272.6111, 272.4376, 271.8571, 270.8661, 
    269.6723,
  276.3781, 274.843, 273.0133, 272.175, 272.6387, 272.8927, 272.9708, 
    272.3428, 271.6495, 272.5558, 272.8165, 272.1946, 271.6625, 271.2523, 
    270.5023,
  276.503, 275.3891, 272.803, 272.3716, 272.6475, 272.8564, 272.6691, 
    271.7435, 272.0041, 272.7715, 272.505, 272.1409, 271.9148, 271.848, 
    270.8079,
  276.8059, 275.5299, 272.4691, 272.4482, 272.5594, 272.6574, 272.6797, 
    272.6554, 272.7177, 272.8002, 272.6048, 272.1607, 271.7863, 271.8178, 
    271.3204,
  276.6926, 274.5329, 272.212, 272.5407, 272.5888, 272.4499, 272.4806, 
    272.3743, 272.3908, 272.5013, 272.5489, 272.0662, 271.8489, 271.6957, 
    271.8071,
  275.5024, 273.6176, 272.3721, 272.5637, 272.6921, 272.6518, 272.5955, 
    272.1217, 272.3035, 272.7761, 272.6603, 272.178, 271.7561, 271.7014, 
    271.9761,
  274.4258, 272.4156, 272.4321, 272.1924, 271.5922, 271.0398, 272.0684, 
    272.3885, 271.3759, 271.8194, 272.5172, 272.2759, 272.3842, 270.1573, 
    272.5066,
  272.5284, 272.7429, 272.5063, 271.9134, 272.3523, 272.332, 272.2586, 
    272.458, 272.2133, 271.9763, 271.8495, 271.9925, 269.0498, 272.1218, 
    272.6149,
  274.5649, 274.1163, 273.1067, 272.1454, 271.4941, 272.2979, 272.3047, 
    272.614, 272.2346, 272.0578, 271.4378, 271.8378, 268.5228, 270.5839, 
    272.7371,
  275.5524, 274.8285, 273.6525, 272.5849, 272.1844, 272.3978, 272.1593, 
    272.5404, 272.0917, 272.1859, 271.6606, 272.0126, 272.3323, 272.2101, 
    272.6306,
  276.1417, 274.5678, 273.8545, 272.4723, 272.7508, 271.8766, 272.5734, 
    270.1094, 268.8986, 272.2484, 271.7609, 272.2213, 271.0667, 271.9666, 
    272.4401,
  276.43, 274.9373, 273.093, 272.3871, 272.5573, 272.4391, 272.3475, 
    271.0193, 271.1815, 272.0706, 272.1811, 272.2702, 272.5017, 272.0201, 
    272.4929,
  276.519, 275.4382, 272.8747, 272.3998, 272.3613, 272.2902, 271.0108, 
    270.7042, 271.915, 272.2903, 272.4738, 272.6267, 272.6174, 272.3167, 
    272.5417,
  276.7738, 275.5287, 272.5016, 271.7754, 272.1198, 272.2076, 272.3785, 
    272.2482, 272.157, 272.3491, 272.3336, 272.3991, 272.4627, 272.1455, 
    272.4018,
  276.6234, 274.5508, 272.0637, 271.9744, 272.1431, 272.2776, 272.0598, 
    272.1049, 272.2612, 272.2665, 272.3094, 272.3144, 272.3914, 272.442, 
    272.363,
  275.5194, 273.7306, 272.3019, 272.3651, 272.5296, 272.5525, 272.4778, 
    272.0336, 272.1721, 272.4855, 272.5762, 272.338, 272.3203, 272.3188, 
    272.2831,
  277.0735, 272.727, 273.1712, 272.1984, 271.7218, 271.8544, 271.9337, 
    271.9602, 271.9896, 269.5778, 273.252, 271.8145, 271.972, 270.0745, 
    272.4409,
  272.5638, 272.8018, 272.7068, 271.9363, 272.2245, 272.047, 271.7841, 
    272.1074, 271.5534, 271.9695, 272.3726, 272.2826, 267.2344, 271.7552, 
    272.1725,
  274.3676, 274.1567, 273.2983, 272.0465, 272.0185, 272.1003, 271.9296, 
    271.9276, 272.0277, 272.3734, 272.3822, 272.061, 267.1994, 268.6813, 
    272.3692,
  275.2785, 274.8431, 273.8421, 272.6578, 272.1516, 272.5518, 270.0955, 
    272.7745, 272.2686, 271.4318, 272.2987, 271.9897, 268.6005, 270.1673, 
    272.7712,
  276.0078, 274.7242, 274.1344, 272.4105, 272.3761, 272.3108, 272.1942, 
    271.0721, 270.0917, 270.1694, 272.1742, 270.0349, 269.3889, 271.7406, 
    272.945,
  276.296, 275.0078, 273.2466, 272.1957, 271.2124, 271.672, 271.7, 270.2493, 
    270.0671, 269.3256, 269.531, 268.841, 271.114, 272.8136, 272.9349,
  276.4341, 275.4872, 272.696, 272.0736, 272.1591, 272.026, 271.5656, 
    271.9542, 269.5306, 268.9164, 271.92, 272.287, 272.7072, 272.9321, 
    272.9347,
  276.7214, 275.6316, 272.0933, 270.1238, 271.5458, 271.7886, 272.0316, 
    272.0155, 271.6487, 272.4747, 272.1664, 272.7379, 272.8345, 272.8238, 
    272.7758,
  276.6109, 274.6237, 271.9164, 271.8097, 271.8565, 272.0219, 272.2375, 
    272.2772, 272.3954, 272.442, 272.8232, 272.8621, 272.795, 272.6775, 
    272.4989,
  275.6119, 273.9186, 272.1729, 271.618, 272.1661, 272.3418, 271.6628, 
    272.0129, 272.4145, 272.7879, 272.9887, 272.8972, 272.7003, 272.6081, 
    272.3857,
  279.2921, 273.0654, 275.1376, 272.3711, 271.9095, 271.4294, 270.481, 
    270.2238, 270.607, 272.1327, 272.8759, 272.4117, 268.6522, 272.3218, 
    272.455,
  272.7846, 272.8493, 272.7125, 271.9518, 272.0634, 271.6748, 271.5138, 
    271.3443, 271.5718, 270.0969, 269.4746, 268.2523, 268.1786, 271.8232, 
    271.9871,
  274.2144, 273.9681, 273.2253, 272.0292, 271.9846, 270.5249, 271.2299, 
    271.3232, 271.5114, 272.1094, 272.1601, 269.0616, 270.9968, 270.6539, 
    272.5541,
  275.0371, 274.5853, 273.7112, 272.655, 272.0382, 272.0502, 269.7779, 
    271.5265, 271.8387, 271.9564, 269.2071, 270.3598, 271.1068, 271.7093, 
    272.9404,
  275.7684, 274.587, 274.0681, 272.3478, 272.0056, 272.1623, 271.5018, 
    269.8302, 268.4066, 269.4719, 272.2094, 271.5437, 271.2026, 272.5851, 
    273.0232,
  276.1263, 274.9661, 273.3407, 271.903, 271.3043, 272.0956, 272.0589, 
    269.8793, 268.6453, 268.1036, 271.9527, 271.3412, 271.8897, 272.9001, 
    272.9307,
  276.3665, 275.5082, 272.6547, 271.5701, 271.8422, 271.8012, 271.6276, 
    269.5694, 268.2587, 270.4555, 271.8867, 271.8722, 272.7583, 272.8805, 
    272.8986,
  276.7386, 275.7705, 271.7685, 270.9903, 271.657, 271.9482, 272.3183, 
    270.3429, 272.0212, 272.2048, 271.9132, 272.6908, 272.7892, 272.8007, 
    272.797,
  276.9352, 275.022, 272.1631, 271.8477, 272.0211, 271.4298, 271.7767, 
    271.1498, 272.2219, 272.2357, 272.6898, 272.8379, 272.7682, 272.6977, 
    272.5469,
  275.9021, 274.0768, 272.3626, 272.2512, 272.0376, 271.6791, 271.6883, 
    271.3885, 271.2455, 272.1794, 272.9336, 272.8743, 272.7, 272.6037, 
    272.4067,
  281.0798, 273.3346, 276.3502, 272.9138, 272.801, 272.5612, 272.2028, 
    271.9379, 271.4286, 272.0497, 273.3256, 272.4377, 271.928, 272.2927, 
    272.3906,
  273.1426, 272.8526, 272.7195, 272.4477, 272.6991, 272.9136, 272.6664, 
    271.6313, 271.0453, 271.308, 271.2848, 270.766, 271.8136, 271.9052, 
    272.0809,
  274.4266, 274.0204, 273.2068, 272.2733, 272.2191, 271.8762, 272.2286, 
    272.0732, 271.5824, 271.2978, 271.6193, 271.6276, 272.0638, 271.502, 
    272.4303,
  275.0935, 274.4594, 273.5877, 272.9034, 272.1747, 271.8902, 270.1898, 
    271.1822, 271.1901, 271.791, 267.9552, 271.9294, 271.7853, 272.3953, 
    273.0195,
  275.6687, 274.3661, 273.8726, 272.6602, 272.4024, 271.5466, 270.7581, 
    268.4214, 268.3351, 268.1869, 269.4278, 272.371, 272.7121, 272.9846, 
    273.0477,
  275.9384, 274.7592, 273.2486, 272.0719, 272.0392, 271.0492, 270.5219, 
    269.9257, 269.1542, 268.6175, 272.2696, 272.4257, 272.9116, 272.9321, 
    272.9241,
  276.2048, 275.381, 272.8139, 271.8035, 271.5701, 271.2513, 270.9123, 
    270.1803, 269.6833, 270.993, 272.2652, 272.8535, 272.8545, 272.8249, 
    272.8588,
  276.6299, 275.6384, 272.1959, 271.42, 271.2153, 271.0409, 270.7611, 
    269.232, 269.5349, 270.5751, 272.7263, 272.8418, 272.7319, 272.7746, 
    272.772,
  276.7951, 274.8651, 271.994, 271.2895, 271.1425, 270.9088, 270.782, 
    268.4269, 269.6533, 270.3046, 272.7629, 272.7985, 272.7376, 272.7011, 
    272.5926,
  275.9264, 274.1504, 272.3235, 271.3852, 271.145, 271.0929, 271.2024, 
    270.5662, 270.1899, 272.0131, 272.8849, 272.8237, 272.6739, 272.5832, 
    272.3945,
  277.8991, 273.1069, 275.5708, 272.9222, 273.029, 273.0853, 273.0492, 
    272.9716, 272.5315, 272.8619, 273.9372, 272.5132, 271.6312, 271.8383, 
    269.768,
  273.3475, 272.8076, 272.691, 272.666, 272.9539, 273.1514, 273.1287, 
    273.028, 272.705, 272.6463, 272.512, 271.9106, 270.3636, 271.4787, 
    271.9661,
  274.6679, 274.1666, 273.3174, 272.4746, 272.5083, 273.0948, 273.0476, 
    272.9848, 272.6778, 272.1324, 271.8062, 270.8068, 269.6624, 269.6518, 
    272.5835,
  275.2489, 274.5229, 273.6543, 273.1573, 272.5576, 272.524, 271.763, 
    271.9835, 271.9382, 272.0021, 269.8152, 270.0072, 271.525, 272.1935, 
    272.5663,
  275.7661, 274.3861, 273.8619, 273.0683, 272.89, 272.5235, 272.0963, 270.51, 
    268.7574, 270.3612, 271.6615, 271.7431, 271.9834, 272.4135, 272.808,
  275.9515, 274.7054, 273.2581, 272.7395, 272.6709, 272.4151, 271.7825, 
    271.485, 270.5977, 270.3099, 270.5246, 271.7699, 272.6423, 272.8604, 
    272.9357,
  276.1542, 275.2837, 273.1174, 272.3448, 271.6505, 270.4502, 270.3256, 
    270.2154, 270.9191, 271.2927, 272.4911, 272.8016, 272.8086, 272.7843, 
    272.8018,
  276.5249, 275.5829, 272.7491, 271.3941, 270.417, 270.0576, 270.6729, 
    271.176, 271.5983, 272.734, 272.8913, 272.8276, 272.7061, 272.7234, 
    272.7321,
  276.4942, 274.7875, 271.868, 270.6833, 270.6877, 270.7954, 270.8096, 
    271.2916, 272.2262, 272.8326, 272.8411, 272.7813, 272.716, 272.6816, 
    272.6596,
  275.6644, 274.1575, 272.4275, 270.6809, 270.7332, 270.8526, 270.7393, 
    271.8517, 272.593, 272.8926, 272.9146, 272.8212, 272.6488, 272.5425, 
    272.4556,
  277.7828, 273.1527, 275.4878, 272.846, 272.9696, 272.9088, 272.8842, 
    272.9868, 272.811, 272.9741, 274.0854, 273.4173, 272.5867, 273.0333, 
    273.158,
  273.2221, 272.8796, 272.6443, 272.6255, 273.0276, 272.1937, 272.7875, 
    273.002, 272.9466, 272.8177, 273.1302, 272.9083, 272.5749, 272.4183, 
    273.1138,
  274.6933, 274.2636, 273.4304, 272.4031, 272.4019, 271.9291, 271.4, 
    272.5993, 273.0682, 273.0158, 273.0226, 272.9933, 272.4303, 271.9814, 
    272.6761,
  275.3332, 274.6135, 273.7448, 273.1471, 272.4315, 271.8675, 273.1117, 
    273.097, 273.0981, 273.0709, 272.9648, 272.7351, 273.0039, 272.8641, 
    272.1894,
  275.8112, 274.4711, 273.9347, 273.1057, 272.8338, 271.3833, 271.6093, 
    272.9498, 272.4329, 273.0237, 272.906, 272.7675, 272.4881, 272.465, 
    272.4711,
  275.8856, 274.6912, 273.3439, 272.8376, 272.9033, 272.9221, 272.766, 
    272.4359, 272.3342, 272.4524, 272.4857, 272.4353, 272.6545, 272.5673, 
    272.4832,
  276.1193, 275.2519, 273.1787, 272.7205, 272.7289, 272.6387, 272.5887, 
    272.2421, 271.7978, 271.995, 272.4953, 272.6031, 272.4797, 272.3462, 
    272.6329,
  276.4918, 275.5627, 272.73, 272.0061, 272.2573, 272.3907, 272.049, 
    272.0118, 272.2792, 272.3817, 272.5047, 272.2974, 272.5074, 272.5747, 
    272.6729,
  276.4348, 274.8174, 272.3163, 272.1685, 272.4272, 272.5089, 272.2614, 
    272.2186, 272.6398, 272.6988, 272.4167, 272.5615, 272.6916, 272.6754, 
    272.8126,
  275.5827, 274.2703, 272.7865, 272.2589, 272.5127, 272.7721, 272.7359, 
    272.6017, 272.8416, 272.9023, 272.9414, 272.8103, 272.6104, 272.5066, 
    272.6718,
  277.4021, 273.0647, 275.8088, 272.823, 272.7101, 273.3692, 272.6576, 
    272.2553, 271.941, 272.5287, 274.1871, 273.7255, 273.0603, 273.2315, 
    273.0784,
  273.445, 272.9901, 272.9433, 272.4861, 272.9212, 272.9924, 273.0627, 
    272.4652, 271.9956, 272.1986, 273.2295, 273.256, 272.7017, 273.1024, 
    273.1595,
  274.7505, 274.4369, 273.5911, 272.316, 272.7459, 273.1086, 272.9753, 
    272.6111, 272.5028, 272.2973, 272.9789, 272.9726, 272.4888, 272.9411, 
    272.8829,
  275.4625, 274.8104, 273.9588, 273.1245, 272.4501, 272.761, 273.1321, 
    272.915, 272.8983, 273.0021, 273.0584, 272.9344, 272.3086, 273.081, 
    273.0071,
  275.9711, 274.7036, 274.1456, 273.0805, 272.7794, 272.6691, 272.5842, 
    273.0706, 273.1285, 273.1061, 273.0892, 272.7496, 273.0761, 273.0612, 
    272.9442,
  276.0323, 274.873, 273.6024, 272.7302, 272.8456, 272.8945, 272.8206, 
    272.5979, 272.6898, 272.7289, 272.9308, 273.0039, 273.0339, 272.9994, 
    272.9381,
  276.2404, 275.3758, 273.3112, 272.6609, 272.7873, 272.8338, 272.8238, 
    272.8143, 272.7414, 272.725, 272.8071, 272.9216, 272.8449, 272.5976, 
    272.6013,
  276.5096, 275.5707, 273.0471, 272.5883, 272.7658, 272.8007, 272.751, 
    272.7764, 272.8171, 272.8481, 272.822, 272.7342, 272.474, 272.3075, 
    272.4168,
  276.4127, 274.8355, 272.6691, 272.5972, 272.7044, 272.7174, 272.7737, 
    272.7426, 272.8037, 272.8919, 272.7285, 272.6547, 272.4804, 272.5145, 
    272.823,
  275.5783, 274.386, 273.0343, 272.7216, 272.7153, 272.6933, 272.5856, 
    272.5482, 272.8649, 272.9501, 272.9656, 272.6807, 272.4924, 272.4302, 
    273.0064,
  277.2542, 273.2037, 275.2691, 272.7369, 273.0398, 274.2664, 272.9626, 
    272.8249, 272.8492, 272.6248, 273.5771, 273.8486, 273.1631, 273.4089, 
    273.1104,
  273.6978, 273.0707, 273.1883, 272.5714, 273.0929, 273.0623, 272.9841, 
    272.9325, 272.6129, 271.9143, 272.8668, 273.3677, 273.1268, 273.1564, 
    273.1217,
  274.8447, 274.5327, 273.6365, 272.353, 272.7766, 273.1314, 272.8767, 
    272.9215, 272.9863, 271.7072, 272.6241, 273.1066, 273.0761, 273.041, 
    273.0093,
  275.5036, 274.8442, 273.93, 273.0784, 272.4908, 272.7628, 273.1284, 
    272.7821, 272.963, 271.8375, 272.9416, 273.0641, 273.0405, 273.0267, 
    272.937,
  275.9319, 274.6711, 274.09, 272.9492, 272.7429, 272.5886, 272.5948, 
    273.0682, 273.0952, 272.2314, 272.9502, 273.0001, 273.0296, 272.9889, 
    272.9217,
  275.9513, 274.7829, 273.5116, 272.496, 272.7339, 272.8282, 272.7489, 
    272.5316, 272.7245, 272.6127, 272.8316, 272.9506, 272.9952, 272.9198, 
    272.8761,
  276.1307, 275.2816, 273.1681, 272.4247, 272.6209, 272.8189, 272.8529, 
    272.8196, 272.6949, 272.2738, 272.5677, 272.4549, 272.8898, 272.879, 
    272.8387,
  276.4535, 275.4979, 272.8231, 272.5292, 272.6913, 272.8146, 272.7635, 
    272.7711, 272.7271, 272.2181, 272.3928, 272.4781, 272.7491, 272.6274, 
    272.5867,
  276.3761, 274.7826, 272.4377, 272.5608, 272.799, 272.8341, 272.837, 
    272.4727, 272.1699, 272.2858, 272.9111, 272.6713, 272.7205, 272.7143, 
    272.8349,
  275.5514, 274.3994, 272.6319, 272.312, 272.6501, 272.7461, 272.5612, 
    272.3851, 272.3369, 272.5802, 272.4791, 272.8258, 272.6639, 272.5967, 
    272.907,
  277.4802, 273.3079, 274.6265, 272.4947, 273.1168, 273.7265, 272.8964, 
    272.8244, 272.9382, 273.0951, 274.3402, 273.9676, 273.1925, 273.5111, 
    273.1595,
  273.915, 273.1826, 273.1902, 272.4579, 273.1128, 272.938, 272.817, 
    272.8632, 272.7965, 272.9353, 273.5921, 273.2923, 273.1387, 273.157, 
    273.1595,
  274.8413, 274.5139, 273.6596, 272.3453, 272.7713, 273.0143, 272.9969, 
    272.9724, 272.9601, 272.785, 272.7415, 272.6659, 273.0553, 273.0226, 
    273.0585,
  275.4706, 274.8197, 273.9208, 273.1015, 272.5033, 272.7753, 272.9747, 
    272.6016, 272.9257, 272.4629, 272.6159, 272.9087, 273.0262, 272.9855, 
    272.9185,
  275.8342, 274.5969, 274.0807, 272.898, 272.7464, 272.553, 272.5983, 
    272.7128, 273.0953, 272.3319, 272.5447, 272.933, 272.9819, 272.9765, 
    272.9128,
  275.8658, 274.7346, 273.5164, 272.4359, 272.7037, 272.8217, 272.7531, 
    272.541, 272.3674, 272.1202, 272.9011, 272.937, 272.955, 272.9754, 
    272.9793,
  276.0348, 275.2382, 273.103, 272.1606, 272.5728, 272.7998, 272.8558, 
    272.7643, 271.9809, 272.1727, 272.7115, 272.8909, 272.8838, 272.7773, 
    272.6944,
  276.392, 275.4448, 272.6805, 272.3296, 272.6084, 272.7957, 272.7573, 
    272.5606, 272.3255, 272.5717, 272.8432, 272.8212, 272.7564, 272.5768, 
    272.557,
  276.336, 274.7246, 272.5617, 272.7061, 272.795, 272.8309, 272.8216, 
    272.5915, 272.6632, 272.6546, 272.9295, 272.8112, 272.7093, 272.6767, 
    272.8014,
  275.5083, 274.3917, 273.0925, 272.9531, 272.8946, 272.8318, 272.5859, 
    272.4994, 272.6011, 272.9684, 272.9345, 272.8433, 272.6612, 272.6067, 
    272.8925,
  280.3813, 273.7885, 276.4903, 272.5037, 273.3355, 274.5049, 272.9293, 
    272.9308, 273.0469, 273.1404, 274.4956, 274.1579, 273.2041, 273.4029, 
    272.824,
  274.576, 273.6268, 273.5016, 272.4511, 273.3767, 273.5597, 272.8662, 
    272.9422, 272.9235, 273.0238, 273.8923, 273.4922, 273.122, 273.1362, 
    273.1595,
  275.4418, 274.8763, 273.8126, 272.4193, 272.7764, 273.0738, 272.653, 
    272.9181, 272.915, 272.6344, 272.6562, 273.0386, 273.0414, 273.0492, 
    273.0617,
  275.731, 274.9634, 273.9892, 273.2466, 272.4023, 272.819, 273.0736, 
    272.9562, 272.5934, 272.6713, 272.756, 272.8794, 272.8958, 272.7773, 
    272.7809,
  275.872, 274.6136, 274.0875, 272.7894, 272.6944, 272.5857, 272.6722, 
    272.275, 272.5851, 272.8806, 272.5735, 272.8578, 272.9271, 272.7789, 
    272.8436,
  275.8758, 274.7018, 273.519, 272.2215, 272.5929, 272.7717, 272.738, 
    272.6267, 272.8607, 272.7037, 272.845, 272.8747, 272.8314, 272.864, 
    272.8925,
  276.0302, 275.2448, 273.0443, 271.7744, 272.241, 272.6579, 272.7971, 
    272.813, 272.7108, 272.5293, 272.718, 272.8138, 272.805, 272.6768, 
    272.6924,
  276.3979, 275.4312, 272.5934, 271.9436, 272.4569, 272.6853, 272.7233, 
    272.7248, 272.7477, 272.8389, 272.7622, 272.8004, 272.75, 272.5945, 
    272.5528,
  276.3563, 274.6372, 272.5097, 272.6238, 272.7221, 272.809, 272.7938, 
    272.8388, 272.899, 272.9583, 272.9235, 272.8179, 272.7026, 272.6507, 
    272.7908,
  275.5302, 274.3795, 273.0237, 272.9474, 272.9131, 272.8484, 272.6184, 
    272.5673, 272.8413, 272.9647, 272.9297, 272.8608, 272.6626, 272.6367, 
    272.8543,
  280.078, 274.1122, 277.5517, 272.5692, 273.4569, 275.3118, 272.9023, 
    272.9136, 273.1768, 276.2174, 277.0322, 275.7378, 272.7825, 274.5161, 
    273.7459,
  274.7283, 273.9249, 273.8417, 272.6297, 274.7914, 275.6909, 272.8419, 
    272.9003, 272.924, 273.6738, 274.3851, 272.9101, 272.6662, 272.8321, 
    272.9258,
  275.489, 275.0865, 274.0002, 272.6064, 272.8672, 273.1119, 272.5892, 
    272.6012, 272.3997, 272.0231, 271.6277, 271.8057, 272.8223, 273.0052, 
    273.0929,
  275.9742, 275.3848, 274.372, 273.683, 272.3734, 272.9255, 273.1015, 
    272.2021, 271.6153, 271.2524, 271.37, 271.5874, 272.7317, 272.9219, 
    272.8236,
  276.3105, 275.0096, 274.3311, 272.8315, 272.558, 272.313, 272.6356, 
    273.0327, 272.8911, 271.2309, 271.3636, 271.4492, 272.6209, 272.9058, 
    272.2903,
  276.0833, 274.9633, 273.6479, 272.1928, 272.412, 272.6398, 272.435, 
    272.6408, 272.6153, 272.0232, 271.6056, 272.6942, 272.5508, 272.7904, 
    272.5298,
  276.2142, 275.379, 273.0298, 271.8017, 271.9811, 272.6111, 272.7655, 
    272.8099, 272.6896, 271.9633, 272.7072, 272.8153, 272.8314, 272.7111, 
    272.453,
  276.5185, 275.5131, 272.6931, 272.1204, 272.3964, 272.6396, 272.711, 
    272.6646, 272.7788, 272.6955, 272.8071, 272.7976, 272.7253, 272.4609, 
    272.2885,
  276.4568, 274.5331, 272.5327, 272.6771, 272.7172, 272.7653, 272.757, 
    272.8034, 272.9181, 272.9831, 272.9245, 272.737, 272.6461, 272.4698, 
    272.4923,
  275.6086, 274.3764, 272.9533, 272.942, 272.9215, 272.8577, 272.6456, 
    272.6225, 272.9206, 272.9917, 272.881, 272.8165, 272.6483, 272.4889, 
    272.7927,
  277.4829, 274.2249, 277.2755, 272.5737, 273.4837, 275.2364, 272.8642, 
    272.8835, 273.1975, 278.3717, 278.6306, 277.0446, 275.0968, 275.3087, 
    275.1062,
  274.4363, 274.1322, 274.0418, 272.7277, 275.695, 275.7222, 272.8767, 
    272.9234, 272.9286, 274.0445, 276.7812, 273.6413, 272.9386, 273.0575, 
    273.1595,
  275.2946, 275.1934, 274.1448, 272.7014, 273.1462, 273.1445, 272.9479, 
    272.9193, 272.9348, 272.7709, 272.5849, 272.3712, 272.5362, 273.0432, 
    273.1065,
  275.8025, 275.3954, 274.3638, 273.7, 272.2982, 273.0214, 273.1211, 
    272.9458, 272.7035, 272.1809, 272.0075, 272.178, 272.5666, 272.9752, 
    272.9933,
  275.9692, 274.8612, 274.3534, 272.9249, 272.5624, 272.5762, 272.8052, 
    273.1239, 272.6092, 271.9975, 271.8853, 272.1943, 272.646, 272.8148, 
    272.8149,
  276.0424, 274.865, 273.6835, 272.2896, 272.3535, 272.685, 272.6832, 
    272.6293, 272.9033, 272.3338, 272.1591, 272.2976, 272.6448, 272.6128, 
    272.5585,
  276.4406, 275.4367, 273.0027, 271.8257, 271.7776, 272.5694, 272.7685, 
    272.8046, 272.4621, 272.1461, 272.2277, 272.4528, 272.4236, 272.1998, 
    272.0982,
  277.0899, 275.7034, 272.7076, 271.9608, 272.1703, 272.6476, 272.7015, 
    272.6422, 272.2882, 272.5457, 272.2952, 272.2819, 272.2343, 271.9282, 
    271.9103,
  276.8578, 274.6836, 272.54, 272.7134, 272.7159, 272.752, 272.7597, 
    272.7967, 272.8453, 272.8974, 272.5079, 272.3206, 272.1169, 271.9037, 
    272.0006,
  275.7964, 274.4902, 272.9314, 272.9239, 272.9103, 272.877, 272.7079, 
    272.7043, 272.9775, 273.0024, 272.6445, 272.3292, 272.1283, 271.8421, 
    272.5422,
  277.6225, 273.2487, 275.3552, 272.4922, 273.2926, 274.7328, 272.8897, 
    272.8784, 273.0069, 276.1583, 278.1846, 276.8491, 275.6223, 276.1849, 
    277.0156,
  273.8687, 273.6449, 273.9374, 272.7805, 275.0074, 274.9987, 273.0139, 
    272.9732, 272.8813, 273.4633, 276.8913, 274.2543, 273.6129, 273.1988, 
    273.6466,
  274.9979, 274.8626, 274.2088, 272.9085, 273.8365, 273.1766, 273.126, 
    273.0428, 272.9455, 272.8857, 273.2931, 273.0485, 273.0428, 273.2133, 
    273.0964,
  275.8553, 275.3617, 274.499, 273.9244, 272.3151, 273.1908, 272.8431, 
    272.9223, 272.5084, 272.637, 272.7693, 272.8947, 273.0255, 272.9823, 
    272.9578,
  276.0724, 274.8618, 274.5494, 273.2002, 272.5343, 272.4566, 272.8764, 
    272.2452, 270.5597, 272.6326, 272.5893, 272.8023, 272.7462, 272.4646, 
    272.383,
  276.23, 274.8969, 273.938, 272.5838, 272.4249, 272.5988, 272.4619, 
    272.3643, 272.7469, 272.4098, 272.3925, 272.4383, 272.2586, 272.1039, 
    271.8972,
  276.6676, 275.4913, 273.1216, 272.0234, 271.8857, 272.414, 272.5987, 
    272.5974, 272.0535, 271.8073, 272.0949, 272.0159, 271.7938, 270.874, 
    271.6342,
  277.2235, 275.7562, 272.6837, 271.8909, 271.8941, 272.5064, 272.5409, 
    272.3269, 271.9035, 271.9803, 271.6664, 271.6754, 271.5423, 271.6524, 
    271.696,
  277.3566, 274.7302, 272.2124, 272.5416, 272.4949, 272.6788, 272.5762, 
    272.2686, 272.2577, 272.005, 271.8077, 271.7408, 271.6421, 271.6953, 
    271.9101,
  276.3673, 274.6925, 272.8662, 272.9006, 272.9063, 272.8678, 272.418, 
    272.2749, 271.8727, 272.3254, 271.9345, 271.6787, 271.6968, 271.4205, 
    272.4687,
  280.7637, 273.4165, 275.6207, 272.54, 273.3736, 274.9236, 273.0414, 
    272.9306, 273.0971, 278.2652, 279.7242, 277.5707, 277.3481, 277.36, 
    277.0659,
  274.0148, 273.6371, 273.896, 272.9069, 275.7463, 275.1926, 273.0829, 
    273.031, 272.6332, 274.0144, 277.5831, 274.6515, 274.0124, 273.1117, 
    275.2844,
  275.0795, 274.8509, 274.2433, 273.0965, 275.0074, 273.1911, 273.3742, 
    273.081, 272.987, 272.8598, 273.9595, 272.863, 272.4184, 272.413, 272.808,
  275.9083, 275.4234, 274.5255, 274.0474, 272.4626, 273.3979, 273.101, 
    273.0981, 273.0374, 273.0129, 272.984, 272.8787, 272.3008, 272.3242, 
    272.6487,
  276.032, 274.9218, 274.5508, 273.2862, 272.454, 272.405, 273.1075, 
    272.3364, 271.7934, 273.0686, 272.9068, 272.5228, 272.3539, 272.0461, 
    272.4096,
  276.1551, 274.9294, 273.9627, 272.5667, 272.3421, 272.611, 272.5718, 
    272.6204, 272.887, 272.8424, 272.6635, 272.0137, 271.9534, 271.9763, 
    272.3952,
  276.5726, 275.5217, 273.1495, 272.1114, 271.98, 272.2558, 272.6806, 
    272.7221, 272.534, 272.1815, 272.0322, 271.5816, 271.6272, 271.8105, 
    272.3032,
  277.0966, 275.7927, 272.7841, 271.9696, 271.8982, 272.2888, 272.6042, 
    272.4533, 272.2378, 272.0264, 271.7528, 271.3823, 271.8668, 272.2121, 
    272.4376,
  277.2799, 274.7107, 272.3165, 272.2597, 272.3104, 272.5409, 272.4735, 
    272.3768, 272.2022, 271.6862, 271.1803, 271.7073, 272.0432, 272.4477, 
    272.263,
  276.4577, 274.6862, 272.7604, 272.8313, 272.8292, 272.6681, 272.1931, 
    271.9617, 271.6678, 271.5256, 271.6664, 271.7298, 272.2387, 272.5181, 
    272.947,
  277.2579, 273.5791, 275.6911, 272.5902, 273.2861, 274.866, 273.026, 
    272.9546, 273.1756, 279.3677, 280.3901, 277.7664, 277.4262, 277.1878, 
    277.244,
  274.1517, 273.8064, 273.9797, 273.0117, 275.3692, 275.2224, 272.7182, 
    272.9992, 272.9095, 274.2241, 278.43, 275.0877, 274.4089, 273.4264, 
    274.9189,
  275.2119, 275.0014, 274.3602, 273.2314, 274.64, 272.626, 273.2536, 
    272.9676, 272.9767, 272.8985, 274.4887, 273.4854, 273.0199, 273.1108, 
    273.1515,
  276.0671, 275.6948, 274.5885, 274.1452, 272.6302, 273.729, 272.6751, 
    272.9436, 272.5643, 272.99, 272.9874, 273.0251, 273.0041, 272.6747, 
    272.8498,
  276.2652, 275.0289, 274.5155, 273.3224, 272.2988, 272.341, 273.0606, 
    272.3601, 271.9756, 272.9119, 273.0015, 272.9062, 272.7691, 272.4696, 
    272.6606,
  276.2168, 274.9603, 273.8706, 272.5396, 272.1357, 272.5638, 272.5779, 
    272.6417, 272.9628, 272.8474, 272.8703, 272.707, 272.3365, 272.269, 
    272.6104,
  276.5042, 275.4936, 273.0984, 271.9978, 271.9551, 272.0184, 272.7244, 
    272.7377, 272.5179, 272.3599, 272.311, 272.1125, 271.7965, 272.2295, 
    272.473,
  276.886, 275.6464, 272.8051, 271.8991, 271.9523, 272.1191, 272.6383, 
    272.5094, 272.5222, 272.6055, 272.3598, 271.6498, 271.8857, 272.1853, 
    272.3587,
  276.8615, 274.6103, 272.424, 272.2945, 272.111, 272.2624, 272.5952, 
    272.719, 272.8725, 272.6011, 271.7117, 271.433, 271.999, 272.2047, 
    272.6362,
  275.9643, 274.5164, 272.8759, 272.6106, 272.6925, 272.6432, 272.4842, 
    272.516, 272.4908, 271.9386, 271.4854, 271.4188, 272.1585, 272.4953, 
    273.1761,
  280.1588, 274.176, 278.0297, 272.66, 273.0822, 274.1313, 273.0038, 
    272.9218, 273.1395, 277.5391, 280.1473, 278.3629, 279.101, 278.3588, 
    278.2272,
  274.2304, 273.8118, 274.0242, 273.0631, 274.1201, 273.6858, 273.0042, 
    272.9723, 272.8795, 273.926, 278.0524, 275.2498, 274.7857, 275.3572, 
    276.855,
  275.1786, 274.9709, 274.3713, 273.334, 274.729, 272.4655, 272.9485, 
    272.8742, 272.3843, 272.6693, 274.4673, 273.7037, 273.0596, 273.2854, 
    274.4349,
  276.0043, 275.6909, 274.6537, 274.2845, 273.0186, 274.5073, 272.2803, 
    272.6971, 271.9184, 272.7818, 272.8374, 272.9649, 273.0048, 272.9278, 
    272.9681,
  276.3297, 275.2707, 274.7897, 273.634, 272.4017, 272.4799, 273.2065, 
    271.8477, 271.9982, 273.3914, 272.8074, 272.7874, 272.9247, 272.8288, 
    272.8052,
  276.5244, 275.2671, 274.1126, 272.759, 272.0259, 272.3738, 272.5985, 
    272.6744, 273.0042, 272.8654, 272.7668, 272.7313, 272.8709, 272.7706, 
    272.7727,
  276.7728, 275.6684, 273.2332, 272.1085, 272.0391, 271.8868, 272.5393, 
    272.71, 272.5751, 272.3438, 272.4221, 272.694, 272.8102, 272.7458, 
    272.6889,
  277.0497, 275.6906, 272.9044, 272.0113, 272.0739, 271.9632, 272.4449, 
    272.5046, 272.496, 272.7203, 272.7556, 272.6693, 272.7707, 272.4893, 
    272.3226,
  276.938, 274.7628, 272.5117, 272.3428, 272.2399, 272.0495, 272.4564, 
    272.7675, 272.9336, 272.9336, 272.9155, 272.8222, 272.677, 272.1509, 
    272.3725,
  275.9918, 274.5935, 272.9892, 272.688, 272.6925, 272.6831, 272.5568, 
    272.8741, 273.0212, 273.0042, 272.8856, 272.6606, 272.4107, 272.0657, 
    273.0229,
  277.2008, 273.6194, 275.5648, 272.5146, 273.2099, 274.6242, 272.9715, 
    272.8744, 273.0703, 277.9944, 280.4358, 279.2127, 280.8711, 280.2487, 
    279.0269,
  274.2906, 273.8185, 273.9114, 272.9977, 275.0448, 274.8438, 272.986, 
    272.9479, 272.8454, 273.8584, 278.0948, 275.3691, 275.3576, 277.8404, 
    278.0978,
  275.0034, 274.8765, 274.2767, 273.2495, 274.5592, 272.7921, 273.2799, 
    272.9625, 272.9351, 272.8881, 274.5621, 273.8968, 273.0582, 273.4239, 
    275.1157,
  275.8433, 275.4332, 274.3457, 274.0514, 272.8384, 274.2225, 272.52, 
    272.8057, 272.6066, 272.8732, 272.9754, 273.0038, 272.9763, 272.8935, 
    272.9742,
  276.1061, 275.0228, 274.5451, 273.4215, 272.1509, 272.3193, 273.3135, 
    272.2834, 271.6009, 272.9759, 272.8522, 272.9238, 272.9212, 272.8288, 
    272.7289,
  276.4105, 275.1063, 274.0463, 272.7698, 272.0009, 272.1797, 272.4621, 
    272.7685, 273.2967, 272.6258, 272.6081, 272.7214, 272.8164, 272.8163, 
    272.735,
  276.7874, 275.6483, 273.2714, 272.2284, 272.1737, 272.0038, 272.3352, 
    272.5113, 272.3572, 272.1033, 272.2296, 272.3141, 272.4324, 272.658, 
    272.7393,
  277.1458, 275.7407, 273.032, 272.1569, 272.2008, 272.0883, 272.3379, 
    272.493, 272.464, 272.4005, 272.532, 272.7513, 272.7972, 272.7285, 
    272.6832,
  277.0294, 274.8671, 272.6943, 272.2971, 272.33, 272.134, 272.4897, 
    272.7726, 272.8688, 272.9026, 272.8937, 272.8665, 272.7997, 272.668, 
    272.58,
  276.0444, 274.64, 272.9167, 272.6556, 272.6721, 272.6385, 272.5249, 
    272.7017, 272.9188, 272.9828, 272.9156, 272.8096, 272.7026, 272.3766, 
    272.9654,
  275.5519, 273.5087, 274.8569, 272.5398, 273.0481, 274.2663, 272.2022, 
    271.9519, 272.1597, 274.7657, 276.8483, 275.9606, 275.9751, 277.4948, 
    278.8025,
  274.3099, 273.8723, 273.8364, 272.9428, 274.4138, 274.5631, 271.9526, 
    272.0846, 272.086, 272.9352, 275.6558, 275.0893, 274.0619, 274.7299, 
    276.6468,
  275.1906, 275.0038, 274.3994, 273.2411, 274.1623, 272.0884, 272.9337, 
    272.0728, 272.1328, 272.048, 272.9982, 273.5262, 273.0062, 273.2358, 
    274.3709,
  276.2, 275.6939, 274.4896, 274.0186, 272.8241, 274.0147, 271.9152, 
    272.0824, 272.3615, 272.1242, 272.8343, 272.8994, 272.8726, 272.8676, 
    273.1008,
  276.4092, 275.3236, 274.6637, 273.3875, 272.1766, 272.447, 273.3474, 
    271.0501, 270.5595, 273.0949, 272.9267, 272.9099, 272.8578, 272.779, 
    272.6591,
  276.6902, 275.3759, 274.2026, 272.8372, 272.0442, 272.1475, 272.5086, 
    272.826, 273.0505, 272.9058, 272.9455, 272.9361, 272.8938, 272.8056, 
    272.6978,
  276.9845, 275.888, 273.4469, 272.321, 272.2641, 272.1404, 272.1902, 
    272.6076, 272.5228, 272.4341, 272.6521, 272.9124, 272.8381, 272.7802, 
    272.7375,
  277.4921, 276.0341, 273.2512, 272.2963, 272.314, 272.2553, 272.2797, 
    272.5009, 272.6027, 272.8034, 272.914, 272.907, 272.7994, 272.7217, 
    272.7076,
  277.2783, 275.0465, 272.8667, 272.37, 272.3438, 272.0696, 272.5262, 
    272.7784, 272.8352, 272.9438, 272.9833, 272.9164, 272.8221, 272.6936, 
    272.7287,
  276.0869, 274.6623, 272.8804, 272.7026, 272.6719, 272.6699, 272.4599, 
    272.6686, 272.9073, 272.9883, 273.0289, 272.8914, 272.7362, 272.6908, 
    273.0596,
  279.2404, 274.0419, 278.0646, 272.6987, 273.5706, 276.0883, 272.9312, 
    272.874, 273.0444, 277.1561, 279.2295, 276.886, 276.1609, 276.8831, 
    276.5498,
  274.0646, 273.7154, 273.7238, 272.9438, 275.7325, 275.2671, 272.8848, 
    272.7101, 272.7545, 273.7474, 277.3479, 275.5177, 273.8887, 274.8721, 
    275.382,
  274.9185, 274.781, 274.2178, 273.1653, 274.2356, 272.548, 272.9383, 
    272.7499, 272.7897, 272.7618, 273.4618, 273.2718, 272.9733, 273.3051, 
    274.4591,
  275.9454, 275.4562, 274.309, 273.9332, 272.8382, 273.8748, 272.3533, 
    272.4243, 272.825, 272.7999, 272.9508, 272.8489, 272.7742, 272.8948, 
    273.715,
  276.3643, 275.2339, 274.6266, 273.4445, 272.2048, 272.4396, 273.4819, 
    271.9206, 271.487, 273.6219, 272.8186, 272.8787, 272.7879, 272.665, 
    272.5956,
  276.8567, 275.4499, 274.3016, 273.0205, 272.2043, 272.1923, 272.4937, 
    272.9746, 273.6288, 272.9687, 272.7876, 272.8961, 272.8404, 272.2642, 
    272.3685,
  277.2607, 276.0008, 273.5645, 272.5103, 272.4562, 272.3557, 272.1783, 
    272.6097, 272.5198, 272.4233, 272.6297, 272.2721, 271.8097, 271.9138, 
    272.684,
  277.7109, 276.1736, 273.5394, 272.5514, 272.5417, 272.5219, 272.1311, 
    272.4434, 272.6661, 272.7968, 272.4902, 272.3257, 271.6138, 272.6195, 
    272.7007,
  277.4166, 275.1023, 273.1573, 272.4358, 272.3214, 272.1212, 272.4252, 
    272.7014, 272.7926, 272.8782, 272.8218, 272.7372, 272.7314, 272.6955, 
    272.7379,
  276.1703, 274.6893, 272.9687, 272.5559, 272.6228, 272.5614, 272.3929, 
    272.5765, 272.4561, 272.9669, 272.9551, 272.8679, 272.723, 272.697, 
    273.0753,
  276.713, 274.2551, 276.8753, 273.3724, 273.7264, 277.6549, 272.9287, 
    272.903, 273.4205, 284.4755, 285.1221, 280.0549, 280.0976, 278.7163, 
    278.9743,
  274.0962, 273.7991, 273.9782, 273.3164, 277.9975, 279.6996, 272.9338, 
    272.9265, 272.8857, 275.4826, 282.4899, 276.4921, 274.5232, 276.9482, 
    277.8785,
  274.8137, 274.7716, 274.3521, 273.3762, 276.2747, 273.1876, 274.1651, 
    272.9625, 272.9232, 272.8518, 274.0307, 273.8061, 273.0268, 273.3972, 
    275.3516,
  275.8213, 275.3491, 274.2747, 274.0871, 273.0098, 276.102, 273.2011, 
    273.3167, 272.9712, 272.9666, 272.9488, 272.8777, 272.8269, 272.9822, 
    274.1599,
  276.1573, 275.0194, 274.5098, 273.491, 272.4723, 272.5841, 273.5896, 
    273.2717, 273.0194, 274.5382, 272.9557, 272.9127, 272.8313, 272.6992, 
    272.6822,
  276.5231, 275.1678, 274.113, 272.935, 272.2144, 272.3583, 272.5122, 
    272.9865, 274.4525, 273.0147, 273.0248, 272.8941, 272.8812, 272.7246, 
    272.6216,
  277.0439, 275.7812, 273.3415, 272.4027, 272.4099, 272.3149, 272.2412, 
    272.6774, 272.5215, 272.3784, 272.6829, 272.8352, 272.7612, 272.6753, 
    272.6559,
  277.5981, 276.0219, 273.3214, 272.4237, 272.4092, 272.3829, 272.0461, 
    272.4977, 272.5637, 272.7036, 272.7951, 272.7589, 272.5011, 272.5865, 
    272.6597,
  277.4576, 275.0083, 272.9706, 272.0711, 271.9678, 271.909, 272.3496, 
    272.7827, 272.7975, 272.849, 272.7616, 272.7053, 272.6742, 272.6002, 
    272.8133,
  276.2198, 274.5854, 272.6932, 272.1703, 272.244, 272.1089, 272.2468, 
    272.5148, 272.7076, 272.762, 272.7728, 272.7143, 272.5624, 272.5721, 
    273.1899,
  275.4336, 274.0086, 275.9201, 273.4407, 273.7078, 277.4742, 272.9205, 
    272.886, 273.485, 286.714, 288.477, 283.3762, 285.9019, 283.8677, 283.9285,
  274.1101, 273.7782, 273.9411, 273.4574, 277.122, 277.8047, 272.9232, 
    272.9029, 272.9046, 275.9063, 286.0387, 278.509, 276.0206, 283.7354, 
    282.7821,
  274.8278, 274.7649, 274.3235, 273.4651, 275.2802, 273.1886, 273.7702, 
    272.9283, 272.9143, 272.896, 274.7279, 274.8071, 273.0949, 273.8529, 
    277.8012,
  275.8635, 275.3487, 274.2906, 274.0842, 273.1297, 275.2067, 273.2307, 
    273.863, 272.9311, 272.9163, 272.9113, 272.8837, 272.8893, 273.3019, 
    275.2271,
  276.2364, 275.0278, 274.5235, 273.5851, 272.4673, 272.6155, 273.944, 
    273.3405, 273.0652, 275.8068, 273.0161, 272.8571, 272.8399, 272.767, 
    272.686,
  276.5691, 275.168, 274.1138, 273.0028, 272.3221, 272.299, 272.4404, 
    273.0557, 274.6088, 273.1491, 274.4776, 272.8594, 272.8739, 272.759, 
    272.6557,
  277.0863, 275.7628, 273.3215, 272.4481, 272.4893, 272.423, 272.2064, 
    272.5344, 272.4557, 272.3837, 272.6209, 272.8509, 272.8457, 272.7838, 
    272.7194,
  277.6838, 275.9642, 273.2478, 272.4821, 272.4613, 272.4755, 272.071, 
    272.4158, 272.5591, 272.7409, 272.8023, 272.857, 272.8217, 272.749, 
    272.7677,
  277.6046, 275.0263, 272.9072, 272.4016, 272.2497, 271.9834, 272.3502, 
    272.6757, 272.8276, 272.9626, 272.9636, 272.8976, 272.8353, 272.7233, 
    272.8134,
  276.3275, 274.6617, 272.9213, 272.6278, 272.634, 272.2666, 272.3486, 
    272.5835, 272.8025, 272.982, 273.0547, 272.8732, 272.7328, 272.6702, 
    273.1586,
  274.4872, 273.7008, 276.5768, 273.5479, 274.0886, 277.2379, 272.9171, 
    272.8792, 273.5482, 287.1035, 289.3036, 284.4927, 288.3771, 287.4292, 
    289.3368,
  273.9216, 273.5502, 273.7532, 273.4533, 279.35, 278.4798, 272.9619, 
    272.8958, 272.8965, 276.3719, 287.339, 279.4685, 277.2531, 288.0512, 
    288.3449,
  274.7598, 274.6783, 274.2009, 273.4413, 276.0672, 273.1891, 273.7706, 
    272.9713, 272.9027, 272.8897, 275.5143, 275.9037, 273.1689, 274.0156, 
    280.7956,
  275.8483, 275.3091, 274.2424, 273.9987, 273.0961, 275.8153, 273.2364, 
    273.9287, 272.9728, 272.887, 272.8834, 272.8724, 272.8864, 273.341, 
    276.5064,
  276.3148, 275.077, 274.5182, 273.5983, 272.4299, 272.5747, 274.3952, 
    273.3811, 273.0739, 274.2151, 272.9402, 272.8436, 272.8246, 272.7687, 
    272.7121,
  276.8001, 275.2876, 274.1645, 273.0504, 272.332, 272.1989, 272.3242, 
    273.1702, 274.1125, 273.738, 274.1162, 272.8431, 272.8441, 272.7446, 
    272.6759,
  277.4709, 276.1354, 273.5971, 272.5922, 272.5344, 272.4718, 272.1312, 
    272.4144, 272.4233, 272.4701, 272.6684, 272.8439, 272.7732, 272.7545, 
    272.6941,
  277.9716, 276.3522, 273.7386, 272.8255, 272.5804, 272.5979, 272.0271, 
    272.3206, 272.4377, 272.6518, 272.8136, 272.8629, 272.7189, 272.6264, 
    272.7491,
  277.7479, 275.3229, 273.2059, 272.4334, 272.2861, 272.2143, 272.0943, 
    272.437, 272.6074, 272.6844, 272.7503, 272.5656, 272.6796, 272.6611, 
    272.6984,
  276.4928, 274.7937, 273.0494, 272.7394, 272.7116, 272.1305, 272.2337, 
    272.3926, 272.5624, 272.682, 272.784, 272.6776, 272.574, 272.4937, 
    273.0894,
  274.9123, 273.8353, 276.6247, 273.9548, 274.7001, 276.8957, 272.8669, 
    272.8712, 273.5131, 286.9084, 289.1698, 284.4406, 288.1957, 287.6051, 
    290.554,
  273.5962, 273.4921, 273.8503, 273.8041, 281.0034, 279.2492, 272.9693, 
    272.9469, 272.9153, 276.3768, 287.6616, 280.4707, 279.068, 288.4808, 
    290.2241,
  274.4449, 274.5237, 274.3229, 273.8281, 278.7845, 273.2062, 273.9697, 
    273.0061, 272.9619, 272.9712, 276.6014, 277.6299, 273.625, 274.096, 
    281.9715,
  275.6748, 275.1413, 274.2346, 274.39, 273.6494, 277.5532, 273.2656, 
    274.7911, 272.9958, 272.9309, 272.8997, 272.9347, 272.9439, 273.4577, 
    277.1407,
  276.1445, 274.9131, 274.3941, 273.662, 272.8549, 272.8338, 275.2036, 
    273.4712, 273.0829, 275.8973, 273.1108, 272.8493, 272.8509, 272.8152, 
    272.7469,
  276.56, 275.1211, 274.0614, 272.8746, 272.4323, 272.4987, 272.4169, 
    273.5133, 276.3528, 275.2004, 275.3004, 272.8325, 272.8399, 272.7469, 
    272.6756,
  277.3025, 275.8415, 273.358, 272.4226, 272.4703, 272.5673, 272.3743, 
    272.6333, 272.5634, 272.5389, 272.6918, 272.8391, 272.8391, 272.7629, 
    272.6832,
  277.9917, 276.2326, 273.5077, 272.5996, 272.4897, 272.5493, 272.1166, 
    272.4925, 272.6417, 272.764, 272.845, 272.8794, 272.8367, 272.7551, 
    272.7593,
  277.8316, 275.4879, 273.3513, 272.1338, 271.8802, 272.1019, 272.1255, 
    272.5931, 272.7188, 272.7941, 272.8463, 272.8707, 272.815, 272.7453, 
    272.7913,
  276.8305, 275.2286, 273.1208, 272.5558, 272.309, 271.6907, 271.9033, 
    272.3005, 272.4935, 272.6437, 272.8499, 272.778, 272.7229, 272.6348, 
    273.1577,
  274.3991, 273.7768, 275.8335, 274.1709, 274.4199, 275.5328, 272.7982, 
    272.8318, 273.3348, 287.2235, 288.8983, 284.0172, 287.0425, 286.7821, 
    288.6121,
  273.5799, 273.5104, 274.0629, 273.9556, 277.3849, 276.917, 272.9313, 
    272.8776, 272.7687, 276.3467, 287.5812, 281.3407, 280.5276, 287.6961, 
    289.042,
  274.3416, 274.5337, 274.6311, 273.9371, 276.5168, 272.6873, 274.0765, 
    272.9547, 272.9081, 272.9893, 277.2021, 279.2519, 274.9246, 274.0301, 
    281.8031,
  275.6074, 275.1267, 274.4807, 274.5526, 273.9037, 277.2749, 273.2969, 
    274.8865, 272.9611, 272.947, 272.9581, 273.1028, 272.9915, 273.5235, 
    277.2545,
  275.938, 274.7928, 274.3931, 274.1989, 273.1308, 273.0826, 275.8336, 
    273.562, 273.07, 276.0146, 273.1772, 272.8651, 272.8633, 272.8662, 272.802,
  276.3593, 274.9771, 274.0098, 272.955, 272.8395, 272.6412, 272.3556, 
    273.679, 277.0745, 276.105, 275.9076, 272.8138, 272.8429, 272.7956, 
    272.7515,
  277.0752, 275.6185, 273.2352, 272.3586, 272.6649, 272.8029, 272.5037, 
    272.5993, 272.6222, 272.619, 272.6835, 272.8008, 272.8381, 272.7822, 
    272.7308,
  277.7996, 275.9915, 273.3013, 272.4975, 272.5095, 272.8096, 272.2019, 
    272.4072, 272.608, 272.7269, 272.8372, 272.867, 272.8382, 272.7746, 
    272.7998,
  277.741, 275.3373, 273.1165, 272.2536, 271.9516, 272.1458, 272.3232, 
    272.7287, 272.8538, 272.9349, 272.9268, 272.8896, 272.8533, 272.7888, 
    272.9945,
  277.0654, 275.3706, 272.8911, 272.5435, 272.3156, 271.8303, 272.43, 
    272.6624, 272.883, 272.9532, 273.0774, 272.8616, 272.8145, 272.6957, 
    273.2587,
  276.562, 273.8059, 275.2944, 274.1802, 274.0682, 274.4641, 272.7345, 
    272.5078, 272.6722, 281.1562, 287.4497, 283.3395, 284.8742, 285.1127, 
    286.2331,
  273.6652, 273.5172, 274.0293, 274.0123, 275.7304, 275.3548, 272.8163, 
    272.5058, 272.2378, 274.9931, 285.9301, 281.7635, 281.1473, 285.4304, 
    286.7089,
  274.3621, 274.579, 274.6064, 273.9422, 275.5488, 272.8352, 273.8551, 
    272.446, 272.4323, 272.9071, 278.0688, 281.0569, 276.6753, 274.0086, 
    281.0578,
  275.6834, 275.1562, 274.4814, 274.4941, 273.9296, 276.8839, 273.2584, 
    273.8144, 272.541, 272.9075, 272.9967, 273.5543, 273.1227, 273.5124, 
    277.5645,
  275.9427, 274.7999, 274.4421, 274.3439, 273.1577, 273.6251, 276.0678, 
    273.3111, 272.8832, 275.523, 273.1017, 272.7018, 272.8044, 272.8196, 
    272.8649,
  276.3964, 274.9258, 274.022, 273.1808, 273.0231, 273.0077, 272.6931, 
    273.8361, 276.5591, 276.1674, 275.7715, 272.7739, 272.7744, 272.7823, 
    272.7466,
  277.0909, 275.5655, 273.2268, 272.5002, 273.0553, 273.0962, 272.6544, 
    272.4533, 272.5923, 272.7084, 272.7503, 272.7918, 272.8404, 272.8014, 
    272.718,
  277.8438, 275.9167, 273.2798, 272.5245, 272.7034, 273.2038, 272.3452, 
    272.2225, 272.6071, 272.7433, 272.8144, 272.868, 272.8479, 272.7925, 
    272.7405,
  277.8217, 275.402, 273.0925, 272.3175, 272.0656, 272.3594, 272.122, 
    272.7169, 272.9001, 272.9893, 272.9188, 272.8921, 272.8693, 272.8172, 
    273.1926,
  277.3241, 275.6424, 273.108, 272.4545, 272.2977, 271.9115, 272.35, 
    272.6562, 272.9221, 272.9505, 273.1641, 272.8458, 272.8394, 272.6763, 
    273.3712,
  280.3509, 274.7863, 276.7858, 274.2893, 274.1751, 274.2298, 272.8154, 
    272.7716, 272.4754, 277.3114, 281.3319, 282.1646, 284.9293, 285.2046, 
    286.56,
  274.4344, 274.0073, 274.2206, 274.1497, 275.9526, 275.0471, 272.8193, 
    272.7537, 272.2081, 274.2938, 281.0982, 281.7822, 281.5359, 284.6557, 
    286.2341,
  274.9033, 274.8331, 274.6248, 274.06, 275.7155, 273.2813, 273.2283, 
    272.7093, 272.4532, 272.9913, 278.4995, 282.1751, 278.1616, 274.1779, 
    280.1685,
  276.0673, 275.3984, 274.4917, 274.4869, 273.9612, 275.882, 272.5621, 
    274.0278, 272.636, 272.8484, 273.0787, 274.1045, 273.2404, 273.4779, 
    276.8181,
  276.209, 275.06, 274.5861, 274.0182, 273.1576, 273.4848, 275.3623, 
    272.0544, 272.2197, 274.7399, 272.9285, 272.7253, 272.936, 273.045, 
    273.205,
  276.7558, 275.1859, 274.0948, 273.0568, 272.8207, 272.9069, 272.7737, 
    273.7493, 275.0993, 275.7279, 275.0151, 272.5721, 272.5044, 272.5775, 
    272.7536,
  277.3658, 275.6243, 273.2826, 272.5414, 272.8743, 273.026, 272.7472, 
    272.3562, 272.5527, 272.7516, 272.7672, 272.7571, 272.7541, 272.5817, 
    272.5999,
  277.9421, 275.9112, 273.3897, 272.5903, 272.7074, 273.0926, 272.4706, 
    272.209, 272.5201, 272.6702, 272.7561, 272.7911, 272.7448, 272.5406, 
    272.5404,
  277.8169, 275.3797, 273.1129, 272.449, 272.1786, 272.4112, 272.0942, 
    272.6148, 272.8292, 272.8824, 272.8437, 272.7129, 272.5513, 272.4868, 
    272.9633,
  277.203, 275.5735, 273.2179, 272.4599, 272.3949, 272.0152, 272.2073, 
    272.6062, 272.7424, 273.2038, 273.3915, 272.8418, 272.7375, 272.6261, 
    273.4028,
  280.1353, 275.5596, 276.705, 274.669, 274.5348, 273.888, 272.7908, 
    272.8291, 272.9425, 276.8592, 283.168, 283.7115, 286.0356, 286.7682, 
    288.5278,
  275.1132, 274.5292, 275.0169, 274.7505, 276.7535, 275.2752, 272.6274, 
    272.6729, 272.6813, 274.2413, 281.8799, 282.684, 282.2057, 286.7719, 
    288.3548,
  275.2123, 275.1449, 275.3382, 274.759, 276.4623, 273.4781, 273.3521, 
    272.7664, 272.6681, 273.1387, 278.9989, 282.9974, 279.8004, 274.6159, 
    281.0601,
  276.379, 275.6985, 275.0108, 275.1159, 274.5121, 276.5053, 272.7799, 
    273.1957, 272.4135, 272.695, 273.2486, 274.6281, 273.6019, 273.5182, 
    277.2579,
  277.0546, 275.794, 274.9972, 274.3296, 273.4782, 273.7502, 275.4073, 
    272.4896, 271.6346, 273.5755, 272.7585, 272.7357, 273.1579, 273.2191, 
    273.5775,
  277.32, 275.5976, 274.3015, 273.1942, 272.8633, 273.0026, 272.8978, 
    273.7005, 274.6403, 275.2319, 274.306, 272.4744, 272.5725, 272.7379, 
    273.1717,
  277.5314, 275.774, 273.3979, 272.6403, 272.8416, 272.9391, 272.7876, 
    272.2816, 272.5137, 272.7717, 272.7503, 272.4395, 272.4059, 272.5484, 
    272.8509,
  278.0081, 275.9812, 273.5492, 272.6905, 272.7233, 272.9761, 272.5092, 
    272.2305, 272.427, 272.7809, 272.7785, 272.6192, 272.3871, 272.4876, 
    272.7119,
  277.7564, 275.4305, 273.2191, 272.5547, 272.3039, 272.4094, 272.1254, 
    272.4276, 272.8303, 272.7944, 272.7854, 272.539, 272.2715, 272.4447, 
    272.9523,
  276.9515, 275.3599, 273.2441, 272.7621, 272.6375, 272.0728, 272.1749, 
    272.6872, 272.9205, 273.5417, 273.409, 272.6834, 272.1416, 272.4984, 
    273.3936 ;

 zg500 =
  5016.91, 5014.094, 5010.697, 5008.675, 5005.066, 5001.233, 4997.681, 
    4997.488, 4998.486, 4999.898, 5006.186, 5016.654, 5028.275, 5041.976, 
    5056.665,
  5016.206, 5011.117, 5006.529, 5002.919, 4996.127, 4988.95, 4984.727, 
    4978.8, 4975.673, 4977.88, 4981.002, 4991.537, 5003.511, 5020.288, 
    5035.089,
  5016.883, 5010.208, 5003.837, 4998.53, 4988.037, 4981.21, 4965.73, 
    4963.812, 4955.026, 4951.932, 4954.414, 4963.894, 4978.147, 4996.36, 
    5016.882,
  5019.993, 5010.633, 5002.139, 4992.454, 4982.087, 4964.761, 4957.208, 
    4939.52, 4934.744, 4930.263, 4931.304, 4938.6, 4954.128, 4975.777, 
    4999.714,
  5027.089, 5014.977, 5003.647, 4991.393, 4977.18, 4962.76, 4944.542, 
    4934.722, 4922.415, 4912.895, 4915.585, 4921.293, 4937.432, 4958.279, 
    4986.216,
  5036.703, 5023.073, 5008.766, 4994.757, 4977.094, 4960.743, 4944.885, 
    4928.109, 4915.823, 4911.226, 4908.43, 4915.216, 4929.794, 4952.054, 
    4979.129,
  5050.585, 5036.109, 5020.361, 5004.626, 4986.902, 4969.612, 4952.109, 
    4939.521, 4926.878, 4918.279, 4916.16, 4921.684, 4934.462, 4954.931, 
    4979.824,
  5068.113, 5052.827, 5036.68, 5020.674, 5001.375, 4984.267, 4967.755, 
    4953.129, 4942.083, 4936.523, 4934.627, 4938.709, 4950.445, 4968.409, 
    4990.536,
  5088.918, 5073, 5057.331, 5041.878, 5025.108, 5008.585, 4991.771, 4979.022, 
    4968.467, 4961.878, 4960.02, 4963.774, 4973.188, 4988.205, 5007.15,
  5113.09, 5094.551, 5078.841, 5064.938, 5048.704, 5034.159, 5020.718, 
    5007.645, 4997.554, 4991.007, 4990.138, 4993.506, 5001.812, 5014.681, 
    5031.246,
  4964.104, 4953.202, 4942.328, 4937.605, 4933.519, 4931.811, 4931.452, 
    4935.724, 4944.386, 4964.776, 4998.107, 5044.174, 5090.215, 5135.171, 
    5176.324,
  4966.034, 4951.333, 4938.549, 4930.847, 4927.159, 4929.619, 4933.533, 
    4937.159, 4945.868, 4968.191, 4998.967, 5042.122, 5085.641, 5128.601, 
    5164.531,
  4970.005, 4951.095, 4936.989, 4927.704, 4922.616, 4929.083, 4930.461, 
    4941.885, 4951.889, 4969.895, 4999.942, 5038.318, 5080.658, 5116.869, 
    5155.171,
  4978.435, 4955.083, 4938.616, 4924.114, 4920.709, 4917.529, 4931.375, 
    4933.136, 4948.755, 4968.777, 4997.368, 5032.902, 5072.035, 5109.239, 
    5144.242,
  4992.264, 4966.385, 4946.037, 4929.044, 4919.9, 4920.502, 4922.087, 
    4935.609, 4950.612, 4964.158, 4992.821, 5024.387, 5061.628, 5092.841, 
    5127.604,
  5011.583, 4985.819, 4960.647, 4941.922, 4925.928, 4919.717, 4923.883, 
    4927.897, 4938.792, 4961.302, 4983.667, 5014.085, 5048.043, 5081.281, 
    5112.135,
  5033.725, 5009.99, 4984.143, 4961.83, 4944.298, 4932.804, 4927.23, 
    4934.295, 4944.453, 4957.689, 4977.411, 5004.117, 5033.513, 5063.951, 
    5094.141,
  5056.603, 5035.175, 5011.28, 4988.604, 4966.053, 4950.838, 4941.718, 
    4938.495, 4942.396, 4956.289, 4973.072, 4994.976, 5022.196, 5051.031, 
    5079.662,
  5078.818, 5060.523, 5038.536, 5018.315, 4997.584, 4979.124, 4963.716, 
    4958.027, 4958.125, 4963.239, 4974.663, 4992.668, 5015.098, 5040.763, 
    5066.865,
  5101.377, 5084.47, 5065.735, 5046.689, 5025.541, 5007.605, 4991.872, 
    4978.499, 4972.05, 4973.283, 4982.025, 4995.739, 5015.118, 5037.717, 
    5061.255,
  4965.508, 4944.197, 4923.596, 4913.562, 4908.782, 4912.33, 4917.467, 
    4931.029, 4942.224, 4958.373, 4980.552, 5007.733, 5046.747, 5098.196, 
    5150.428,
  4968.215, 4941.938, 4923.159, 4914.503, 4911.2, 4913.987, 4919.35, 
    4928.817, 4938.674, 4961.417, 4987.802, 5021.46, 5068.485, 5125.148, 
    5172.837,
  4969.981, 4944.117, 4926.535, 4920.448, 4917.022, 4921.107, 4923.172, 
    4933.15, 4948.123, 4969.45, 4999.146, 5038.013, 5092.211, 5145.019, 
    5193.941,
  4976.406, 4948.28, 4932.371, 4924.872, 4926.513, 4922.168, 4930.667, 
    4933.588, 4949.201, 4977.421, 5013.403, 5057.654, 5114.255, 5169.787, 
    5215.858,
  4984.003, 4956.619, 4939.627, 4932.04, 4932.65, 4933.905, 4934.578, 
    4944.057, 4968.045, 4989.234, 5030.337, 5078.192, 5137.853, 5186.284, 
    5232.592,
  4995.375, 4966.984, 4948.457, 4940.18, 4938.078, 4939.297, 4945.333, 
    4953.818, 4970.108, 5007.158, 5046.791, 5099.585, 5157.061, 5208.498, 
    5249.951,
  5009.294, 4981.26, 4960.468, 4950.643, 4947.007, 4949.817, 4954.341, 
    4971.055, 4996.217, 5026.274, 5067.87, 5121.389, 5174.519, 5222.446, 
    5264.068,
  5026.051, 4998.171, 4975.44, 4963.4, 4956.414, 4958.649, 4967.528, 4982.09, 
    5004.496, 5041.886, 5086.996, 5139.354, 5192.006, 5238.196, 5278.934,
  5042.819, 5017.827, 4994.755, 4980.218, 4973.251, 4973.764, 4981.654, 
    5001.744, 5028.396, 5062.28, 5105.221, 5156.646, 5205.822, 5249.696, 
    5288.351,
  5060.666, 5037.698, 5016.102, 5000.58, 4990.569, 4989.736, 4998.146, 
    5014.641, 5039.758, 5075.888, 5121.016, 5170.665, 5217.324, 5259.624, 
    5295.835,
  5053.167, 5034.066, 5017.181, 5009.562, 5002.811, 4998.091, 5001.071, 
    5014.876, 5030.06, 5042.117, 5058.143, 5081.231, 5112.723, 5143.874, 
    5176.053,
  5046.434, 5026.462, 5013.63, 5007.519, 5001.949, 5002.713, 5010.118, 
    5021.775, 5033.044, 5050.947, 5070.96, 5100.558, 5134.02, 5168.096, 
    5195.719,
  5037.902, 5019.254, 5009.813, 5007.252, 5004.847, 5011.55, 5015.954, 
    5033.975, 5048.736, 5062.968, 5087.302, 5120.816, 5155.892, 5185.038, 
    5211.652,
  5029.856, 5012.571, 5007.586, 5006.389, 5010.77, 5010.862, 5030.393, 
    5034.533, 5049.026, 5074.232, 5106.404, 5142.636, 5176.698, 5205.834, 
    5229.465,
  5021.601, 5009.204, 5006.215, 5008.668, 5012.692, 5023.625, 5030.677, 
    5049.259, 5072.149, 5090.511, 5129.556, 5163.571, 5197.002, 5219.525, 
    5241.724,
  5016.2, 5005.823, 5005.415, 5009.868, 5015.449, 5027.671, 5044.927, 
    5056.488, 5074.915, 5116.541, 5152.265, 5185.941, 5214.141, 5236.432, 
    5254.701,
  5011.336, 5005.644, 5008.044, 5013.108, 5021.902, 5035.701, 5051.525, 
    5076.204, 5108.191, 5142.523, 5175.876, 5206.787, 5229.801, 5249.096, 
    5267.563,
  5009.104, 5006.202, 5009.635, 5016.567, 5026.64, 5043.299, 5064.335, 
    5088.217, 5123.378, 5164.26, 5197.128, 5224.087, 5246.213, 5265.849, 
    5286.25,
  5008.533, 5010.289, 5016.562, 5024.48, 5038.133, 5055.566, 5079.263, 
    5115.556, 5155.787, 5188.698, 5217.145, 5241.263, 5263.069, 5284.27, 
    5308.26,
  5013.157, 5015.617, 5023.226, 5034.171, 5049.35, 5071.506, 5101.128, 
    5136.22, 5173.045, 5207.396, 5235.589, 5260.025, 5284.029, 5309.16, 
    5336.947,
  5179.965, 5178.492, 5168.348, 5155.463, 5139.925, 5127.719, 5122.734, 
    5124.899, 5132.28, 5143.704, 5167.479, 5200.307, 5236.374, 5269.353, 
    5303.806,
  5170.919, 5168.969, 5160.629, 5150.466, 5135.013, 5128.077, 5126.967, 
    5128.158, 5136.224, 5157.32, 5186.104, 5224.292, 5258.864, 5296.95, 
    5325.595,
  5161.221, 5159.636, 5152.942, 5144.043, 5133.692, 5131.419, 5129.407, 
    5139.097, 5153.175, 5172.683, 5207.512, 5244.565, 5280.532, 5312.75, 
    5343.656,
  5150.37, 5148.356, 5143.239, 5136.951, 5133.415, 5130.764, 5138.978, 
    5140.056, 5155.931, 5189.007, 5226.767, 5263.86, 5300.461, 5333.773, 
    5363.617,
  5138.666, 5137.86, 5134.233, 5132.593, 5131.871, 5139.424, 5140.556, 
    5156.744, 5182.905, 5205.73, 5246.537, 5281.227, 5317.599, 5346.397, 
    5376.268,
  5125.947, 5125.923, 5123.713, 5126.611, 5131.405, 5140.32, 5153.741, 
    5163.222, 5184.769, 5227.385, 5263.923, 5299.275, 5332.004, 5361.696, 
    5388.354,
  5114.322, 5116.938, 5117.978, 5124.765, 5134.271, 5147.301, 5159.118, 
    5182.841, 5215.464, 5248.092, 5282.717, 5315.061, 5344.748, 5371.259, 
    5395.952,
  5104.532, 5108.853, 5112.482, 5123.481, 5136.456, 5152.312, 5169.974, 
    5191.905, 5223.057, 5262.836, 5296.661, 5327.369, 5355.673, 5381.037, 
    5404.72,
  5096.738, 5104.775, 5114.322, 5128.335, 5144.333, 5161.17, 5181.11, 
    5212.636, 5249.272, 5281.499, 5310.74, 5338.636, 5363.901, 5387.605, 
    5410.075,
  5091.924, 5102.128, 5115.279, 5132.816, 5151.35, 5172.238, 5196.762, 
    5226.804, 5260.731, 5293.474, 5322.507, 5347.812, 5371.587, 5394.847, 
    5417.328,
  5233.297, 5242.573, 5250.869, 5257.121, 5256.113, 5248.693, 5250.685, 
    5268.249, 5292.704, 5319.059, 5345.813, 5369.455, 5389.122, 5402.452, 
    5411.551,
  5225.122, 5234.228, 5244.375, 5252.137, 5251.38, 5246.3, 5250.322, 
    5267.345, 5293.993, 5328.791, 5358.56, 5385.494, 5404.92, 5420.778, 
    5428.75,
  5217.466, 5227.001, 5239.259, 5248.47, 5249.897, 5245.475, 5249.286, 
    5273.033, 5305.125, 5337.419, 5370.144, 5398.114, 5420.39, 5434.864, 
    5444.518,
  5210.694, 5220.647, 5233.517, 5243.054, 5247.887, 5241.056, 5251.527, 
    5265.611, 5300.106, 5342.21, 5379.124, 5408.378, 5432.768, 5448.653, 
    5459.307,
  5203.421, 5214.807, 5227.973, 5239.609, 5242.719, 5245.677, 5244.671, 
    5274.482, 5312.913, 5346.203, 5386.003, 5417.435, 5443.11, 5459.305, 
    5470.628,
  5195.087, 5208.192, 5220.829, 5232.602, 5236.883, 5238.519, 5248.397, 
    5265.25, 5300.565, 5352.047, 5390.25, 5425.393, 5450.791, 5469.892, 
    5480.67,
  5186.447, 5201.258, 5214.364, 5226.139, 5232.044, 5236.194, 5242.479, 
    5269.534, 5313.333, 5354.024, 5395.351, 5430.576, 5457.487, 5476.848, 
    5487.834,
  5178.374, 5194.044, 5205.89, 5217.756, 5223.616, 5230.45, 5239.363, 
    5258.304, 5300.479, 5353.015, 5396.491, 5433.473, 5461.814, 5481.93, 
    5493.266,
  5171.337, 5187.92, 5199.991, 5212.035, 5219.223, 5225.357, 5236.141, 
    5260.119, 5306.741, 5354.842, 5396.884, 5435.836, 5463.626, 5484.258, 
    5494.451,
  5165.549, 5181.38, 5192.499, 5204.688, 5212.793, 5220.438, 5232.735, 
    5251.987, 5297.253, 5350.659, 5396.982, 5436.067, 5464.341, 5484.622, 
    5494.305,
  5304.342, 5295.548, 5295.882, 5302.979, 5309.552, 5325.196, 5342.271, 
    5358.164, 5369.121, 5373.128, 5373.361, 5371.386, 5365.783, 5357.827, 
    5348.687,
  5302.169, 5294.971, 5295.469, 5302.486, 5307.183, 5324.304, 5345.019, 
    5361.892, 5373.83, 5384.091, 5386.797, 5387.224, 5382.823, 5378.602, 
    5371.389,
  5296.761, 5292.204, 5293.819, 5301.368, 5306.707, 5324.667, 5344.724, 
    5368.631, 5385.419, 5394, 5398.711, 5400.163, 5398.537, 5394.422, 5388.685,
  5286.5, 5286.844, 5289.351, 5296.836, 5305.753, 5317.615, 5348.11, 
    5365.288, 5386.204, 5400.51, 5409.357, 5410.796, 5411.138, 5407.304, 
    5403.961,
  5273.489, 5278.876, 5283.599, 5294.308, 5301.725, 5319.451, 5341.687, 
    5372.021, 5395.508, 5407.386, 5418.732, 5422.645, 5424.335, 5420.768, 
    5417.125,
  5254.693, 5265.227, 5273.691, 5286.361, 5295.998, 5309.705, 5342.491, 
    5365.466, 5390.757, 5413.823, 5426.14, 5434.199, 5437.083, 5435.911, 
    5431.647,
  5234.334, 5249.127, 5263.425, 5278.929, 5292.087, 5305.242, 5333.7, 
    5368.495, 5397.61, 5416.967, 5433.541, 5444.533, 5450.178, 5450.412, 
    5445.873,
  5216.446, 5233.226, 5249.754, 5268.624, 5283.405, 5297.624, 5326.244, 
    5357.964, 5388.279, 5416.993, 5437.504, 5451.803, 5460.655, 5463.021, 
    5460.061,
  5202.231, 5219.583, 5240.299, 5261.27, 5279.199, 5292.269, 5317.057, 
    5353.853, 5387.07, 5414.876, 5437.829, 5455.863, 5467.656, 5472.538, 
    5470.844,
  5192.268, 5208.158, 5228.499, 5250.641, 5270.745, 5286.146, 5308.207, 
    5340.504, 5373.452, 5406.508, 5434.354, 5455.415, 5470.299, 5477.965, 
    5478.793,
  5305.358, 5300.871, 5294.144, 5289.099, 5293.458, 5295.626, 5292.379, 
    5287.74, 5284.036, 5281.228, 5281.517, 5284.889, 5289.504, 5294.116, 
    5298.63,
  5286.63, 5287.205, 5287.807, 5285.776, 5291.618, 5298.938, 5302.233, 
    5300.458, 5296.928, 5297.403, 5298.584, 5302.704, 5306.599, 5312.124, 
    5317.446,
  5263.654, 5270.401, 5278.108, 5280.729, 5289.494, 5301.805, 5307.004, 
    5311.782, 5312.261, 5312.123, 5314.466, 5318.479, 5324.295, 5329.813, 
    5335.516,
  5242.844, 5254.558, 5267.319, 5273.342, 5284.738, 5298.534, 5312.775, 
    5315.891, 5319.169, 5322.978, 5327.643, 5332.045, 5338.673, 5344.876, 
    5352.235,
  5233.162, 5245.374, 5260.588, 5269.976, 5279.553, 5299.707, 5311.638, 
    5323.576, 5329.331, 5331.127, 5337.231, 5342.729, 5350.661, 5357.801, 
    5365.603,
  5226.101, 5239.761, 5254.969, 5265.957, 5274.018, 5293.788, 5313.596, 
    5324.348, 5330.586, 5338.459, 5344.56, 5352.694, 5361.12, 5370.716, 
    5378.206,
  5223.362, 5237.423, 5252.211, 5263.891, 5272.334, 5290.913, 5310.813, 
    5327.636, 5337.453, 5344.323, 5352.071, 5361.927, 5372.212, 5382.049, 
    5389.128,
  5227.12, 5233.905, 5246.946, 5259.743, 5267.698, 5285.156, 5308.469, 
    5325.439, 5337.292, 5348.973, 5358.99, 5370.699, 5382.082, 5392.369, 
    5399.688,
  5235.562, 5233.456, 5241.332, 5255.797, 5266.669, 5281.458, 5304.097, 
    5325.004, 5340.599, 5352.986, 5365.465, 5379.081, 5391.451, 5401.956, 
    5409.507,
  5236.447, 5235.798, 5235.167, 5246.569, 5260.008, 5274.4, 5297.864, 
    5320.193, 5337.777, 5354.221, 5370.062, 5385.445, 5399.146, 5411.028, 
    5419.344,
  5189.159, 5203.968, 5215.478, 5223.44, 5229.025, 5236.602, 5246.618, 
    5260.452, 5272.687, 5280.221, 5285.386, 5288.685, 5289.299, 5289.144, 
    5288.142,
  5178.89, 5194.617, 5210.849, 5222.227, 5228.845, 5236.762, 5248.552, 
    5261.236, 5274.012, 5286.897, 5294.02, 5298.26, 5299.556, 5300.271, 
    5301.036,
  5172.854, 5187.007, 5206.907, 5220.326, 5230.471, 5238.87, 5247.091, 
    5263.788, 5278.894, 5290.09, 5299.066, 5304.24, 5308.128, 5311.642, 
    5313.863,
  5170.753, 5182.937, 5203.995, 5218.175, 5232.72, 5237.202, 5249.517, 
    5257.836, 5274.701, 5289.965, 5301.91, 5308.493, 5315.835, 5322.102, 
    5325.923,
  5172.601, 5183.566, 5203.731, 5219.771, 5232.457, 5243.738, 5247.486, 
    5262.686, 5278.038, 5289.948, 5303.888, 5313.342, 5324.413, 5332.469, 
    5337.424,
  5178.046, 5187.582, 5205.437, 5220.679, 5233.58, 5242.775, 5252.994, 
    5260.569, 5273.249, 5292.228, 5305.4, 5319.125, 5331.617, 5342.624, 
    5348.202,
  5187.005, 5195.575, 5210.832, 5223.472, 5236.031, 5247.348, 5254.516, 
    5266.46, 5279.765, 5293.312, 5308.444, 5324.034, 5338.991, 5351.27, 
    5358.839,
  5199.008, 5205.745, 5215.714, 5226.112, 5235.663, 5248.203, 5258.082, 
    5266.497, 5277.391, 5294.585, 5310.23, 5327.639, 5344.357, 5358.208, 
    5368.391,
  5208.95, 5213.72, 5220.992, 5228.733, 5236.859, 5249.751, 5260.122, 
    5271.437, 5282.702, 5295.508, 5311.163, 5330.1, 5347.673, 5363.331, 
    5375.363,
  5217.959, 5216.681, 5220.942, 5227.639, 5233.813, 5246.147, 5260.129, 
    5269.937, 5280.294, 5294.26, 5311.1, 5330.016, 5348.852, 5365.774, 
    5380.043,
  5192.384, 5205.438, 5215.158, 5224.75, 5233.345, 5240.052, 5243.388, 
    5244.624, 5242.972, 5235.956, 5226.518, 5214.022, 5199.841, 5183.782, 
    5168.864,
  5199.021, 5212.179, 5223.279, 5235.164, 5244.153, 5251.625, 5257.303, 
    5257.88, 5253.743, 5248.113, 5237.729, 5225.554, 5209.609, 5194.519, 
    5178.134,
  5205.566, 5219.032, 5231.092, 5244.436, 5254.935, 5265.354, 5269.203, 
    5272.688, 5269.524, 5261.404, 5250.039, 5237.431, 5222.654, 5206.666, 
    5190.938,
  5213.3, 5226.396, 5239.056, 5251.309, 5264.364, 5271.541, 5279.899, 
    5280.945, 5279.647, 5273.201, 5263.478, 5250.427, 5237.452, 5222.321, 
    5207.994,
  5221.381, 5233.851, 5245.186, 5257.06, 5267.042, 5277.339, 5282.323, 
    5288.116, 5290.839, 5284.379, 5276.771, 5264.917, 5254.244, 5239.292, 
    5226.601,
  5229.981, 5240.3, 5248.925, 5259.097, 5266.519, 5272.774, 5279.607, 
    5284.469, 5289.961, 5293.032, 5288.383, 5280.828, 5272.388, 5261.104, 
    5249.101,
  5236.389, 5245.388, 5251.334, 5258.739, 5264.065, 5268.586, 5270.746, 
    5278.42, 5288.415, 5296.308, 5297.727, 5296.008, 5291.599, 5284.2, 5274.32,
  5245.249, 5248.621, 5251.905, 5257.456, 5260.324, 5262.636, 5263.725, 
    5266.707, 5278.134, 5294.647, 5303.193, 5309.187, 5311.121, 5309.617, 
    5303.824,
  5252.888, 5248.955, 5250.459, 5253.612, 5257.513, 5259.897, 5259.658, 
    5262.485, 5272.241, 5290.655, 5305.022, 5318.432, 5327.104, 5331.493, 
    5330.609,
  5256.843, 5248.46, 5245.545, 5247.674, 5250.773, 5254.899, 5256.134, 
    5257.296, 5265.06, 5284.442, 5303.331, 5321.813, 5336.14, 5345.407, 
    5349.899,
  5245.714, 5251.382, 5256.781, 5257.951, 5254.151, 5244.2, 5226.433, 
    5208.703, 5190.147, 5170.822, 5155.607, 5142.221, 5131.884, 5121.303, 
    5112.952,
  5254.055, 5259.832, 5265.454, 5267.5, 5264.291, 5252.561, 5240.485, 
    5219.061, 5199.003, 5183.482, 5169.865, 5158.667, 5147.72, 5139.366, 
    5130.569,
  5261.853, 5267.823, 5272.977, 5276.75, 5272.032, 5266.896, 5247.613, 
    5234.315, 5215.811, 5198.223, 5184.817, 5175.122, 5166.261, 5157.767, 
    5149.686,
  5271.296, 5275.298, 5280.504, 5281.731, 5281.186, 5270.293, 5261.3, 
    5242.014, 5225.578, 5211.481, 5200.654, 5191.027, 5184.255, 5176.478, 
    5169.761,
  5282.146, 5283.975, 5286.732, 5287.049, 5285.61, 5278.843, 5266.948, 
    5253.226, 5243.82, 5225.342, 5216.87, 5207.673, 5203.202, 5195.937, 
    5191.14,
  5295.458, 5293.977, 5291.349, 5290.221, 5285.975, 5279.778, 5273.031, 
    5260.479, 5249.489, 5241.138, 5232.531, 5226.289, 5221.931, 5217.487, 
    5212.709,
  5307.862, 5303.92, 5296.983, 5292.693, 5286.697, 5281.212, 5274.415, 
    5268.302, 5263.282, 5255.952, 5249.601, 5246.141, 5242.819, 5240.065, 
    5235.638,
  5318.601, 5309.989, 5300.093, 5293.664, 5285.965, 5279.844, 5275.907, 
    5270.552, 5268.465, 5268.531, 5266.382, 5265.468, 5264.399, 5262.895, 
    5259.472,
  5322.581, 5311.316, 5300.638, 5292.498, 5286.596, 5280.233, 5276.083, 
    5274.514, 5276.444, 5279.735, 5281.706, 5284.617, 5286.021, 5285.755, 
    5282.938,
  5326.018, 5306.965, 5292.997, 5285.806, 5280.672, 5275.892, 5273.604, 
    5272.65, 5276.351, 5285.532, 5292.944, 5299.606, 5303.709, 5305.986, 
    5304.857,
  5286.047, 5286.089, 5279.389, 5267.708, 5254.691, 5241.557, 5228.175, 
    5218.905, 5211.26, 5202.066, 5192.552, 5182.223, 5170.966, 5156.526, 
    5141.234,
  5289.386, 5288.774, 5282.357, 5272.01, 5260.885, 5247.267, 5240.012, 
    5231.692, 5224.035, 5217.88, 5209.976, 5201.14, 5188.545, 5174.721, 
    5157.427,
  5292.017, 5291.443, 5285.95, 5278.349, 5266.672, 5259.236, 5248.211, 
    5243.581, 5239.481, 5234.688, 5227.872, 5220.077, 5208.922, 5193.379, 
    5174.53,
  5297.159, 5295.493, 5290.867, 5282.344, 5274.546, 5263.611, 5259.703, 
    5255.35, 5251.355, 5249.138, 5245.415, 5237.917, 5227.746, 5213.396, 
    5193.997,
  5305.445, 5302.949, 5298.111, 5290.668, 5282.288, 5275.327, 5268.454, 
    5264.347, 5266.351, 5262.802, 5261.165, 5254.744, 5246.928, 5231.966, 
    5214.314,
  5313.308, 5309.233, 5304.083, 5298.103, 5288.793, 5280.884, 5278.292, 
    5275.923, 5274.303, 5275.287, 5274.153, 5269.817, 5263.15, 5251.22, 
    5234.606,
  5316.578, 5309.727, 5305.792, 5303.944, 5297.745, 5290.274, 5284.526, 
    5283.837, 5284.733, 5285.509, 5285.023, 5282.914, 5277.591, 5268.526, 
    5254.337,
  5325.146, 5310.465, 5302.66, 5302.361, 5299.668, 5294.714, 5290.134, 
    5290.118, 5289.909, 5292.245, 5293.321, 5292.599, 5289.583, 5283.279, 
    5272.602,
  5345.56, 5325.15, 5308.95, 5302.488, 5302.091, 5300.154, 5293.805, 
    5294.016, 5294.909, 5296.844, 5299.027, 5299.902, 5298.848, 5295.197, 
    5287.623,
  5368.561, 5349.22, 5329.172, 5313.71, 5305.136, 5302.057, 5297.365, 
    5295.704, 5296.79, 5298.334, 5301.667, 5303.881, 5304.86, 5304.163, 
    5300.296,
  5275.86, 5275.384, 5275.735, 5279.208, 5284.864, 5290.639, 5292.921, 
    5291.918, 5286.478, 5274.062, 5255.934, 5230.146, 5200.646, 5167.651, 
    5137.034,
  5275.185, 5275.539, 5277.714, 5283.134, 5289.435, 5295.869, 5300.306, 
    5300.674, 5294.598, 5285.352, 5268.713, 5246.341, 5215.927, 5183.788, 
    5151.195,
  5275.197, 5278.432, 5282.064, 5288.543, 5294.352, 5301.81, 5305.694, 
    5306.476, 5303.426, 5294.993, 5281.369, 5261.471, 5234.688, 5201.327, 
    5167.821,
  5278.212, 5281.469, 5286.967, 5291.425, 5300.312, 5304.396, 5311.317, 
    5312.213, 5309.131, 5302.297, 5292.229, 5275.17, 5251.996, 5222.582, 
    5189.093,
  5282.329, 5287.58, 5292.696, 5297.118, 5303.139, 5310.545, 5314.079, 
    5315.154, 5314.446, 5307.554, 5300.287, 5287.195, 5269.496, 5242.292, 
    5212.761,
  5287.925, 5292.833, 5296.567, 5301.736, 5306.422, 5311.949, 5317.114, 
    5318.34, 5316.495, 5311.881, 5305.566, 5295.944, 5283.022, 5262.489, 
    5236.214,
  5291.48, 5297.318, 5300.743, 5305.014, 5308.475, 5313.753, 5316.246, 
    5318.531, 5317.502, 5314.127, 5308.642, 5302.108, 5292.584, 5277.812, 
    5256.675,
  5304.238, 5301.531, 5302.307, 5307.157, 5310.125, 5314.201, 5316.881, 
    5318.322, 5317.405, 5315.392, 5310.933, 5305.636, 5299.094, 5289.758, 
    5274.126,
  5326.863, 5320.697, 5315.542, 5313.171, 5313.803, 5315.406, 5316.562, 
    5317.676, 5316.918, 5315.642, 5312.528, 5308.328, 5302.812, 5296.289, 
    5285.798,
  5343.165, 5339.347, 5334.811, 5330.228, 5326.192, 5324.682, 5323.792, 
    5323.016, 5321.83, 5319.787, 5316.542, 5312.122, 5306.634, 5301.155, 
    5293.827,
  5251.763, 5260.902, 5269.228, 5277.066, 5288.11, 5299.447, 5308.009, 
    5312.054, 5311.063, 5302.132, 5287.738, 5266.623, 5241.256, 5209.567, 
    5177.359,
  5245.167, 5253.845, 5262.583, 5272.606, 5283.858, 5297.001, 5307.873, 
    5312.179, 5310.284, 5304.662, 5291.986, 5274.888, 5250.978, 5222.822, 
    5189.547,
  5237.389, 5246.647, 5256.537, 5269.037, 5282.602, 5297.208, 5305.062, 
    5311.613, 5309.498, 5304.488, 5294.5, 5280.439, 5260.698, 5233.213, 
    5201.235,
  5231.418, 5240.75, 5252.066, 5265.605, 5281.539, 5294.546, 5306.271, 
    5309.15, 5308.941, 5303.489, 5295.796, 5284.629, 5268.727, 5246.38, 
    5215.193,
  5227.111, 5237.185, 5249.392, 5264.746, 5280.836, 5296.641, 5303.847, 
    5308.825, 5306.753, 5301.902, 5295.577, 5286.929, 5275.517, 5255.209, 
    5229.076,
  5226.634, 5237.727, 5249.69, 5265.203, 5280.812, 5294.471, 5304.35, 
    5306.834, 5305.433, 5300.988, 5295.566, 5289.091, 5281.166, 5266.29, 
    5243.177,
  5230.159, 5241.324, 5253.09, 5267.462, 5282.26, 5294.477, 5301.26, 
    5304.509, 5302.849, 5299.071, 5295.505, 5291.7, 5285.552, 5273.674, 
    5254.646,
  5238.441, 5248.674, 5258.529, 5270.674, 5281.673, 5291.904, 5298.268, 
    5300.674, 5299.402, 5297.773, 5296, 5295.317, 5291.324, 5282.569, 5267.492,
  5249.758, 5256.78, 5264.111, 5273.378, 5282.33, 5289.633, 5293.133, 
    5294.754, 5294.988, 5296.147, 5298.121, 5299.564, 5296.59, 5288.95, 
    5276.877,
  5267.415, 5270.023, 5273.588, 5278.202, 5282.481, 5287.09, 5290.784, 
    5293.849, 5296.225, 5299.109, 5302.018, 5303.542, 5301.007, 5295.648, 
    5286.039,
  5240.426, 5254.739, 5268.713, 5281.27, 5291.639, 5297.704, 5299.336, 
    5299.871, 5295.539, 5285.706, 5273.326, 5257.298, 5235.28, 5202.33, 
    5168.703,
  5240.312, 5254.481, 5267.333, 5279.488, 5287.854, 5294.535, 5299.804, 
    5296.642, 5293.093, 5287.196, 5275.797, 5263.014, 5240.735, 5211.92, 
    5177.46,
  5237.771, 5251.519, 5264.259, 5276.653, 5286.353, 5292.788, 5292.742, 
    5299.026, 5293.899, 5287.663, 5278.953, 5268.806, 5249.321, 5221.267, 
    5189.549,
  5234.522, 5246.917, 5259.569, 5270.955, 5279.865, 5288.01, 5292.064, 
    5289.479, 5291.29, 5288.074, 5282.417, 5274.755, 5259.305, 5236.167, 
    5207.143,
  5229.445, 5241.11, 5252.788, 5265.016, 5273.91, 5281.082, 5286.609, 
    5291.935, 5291.174, 5287.456, 5285.181, 5280.534, 5268.969, 5248.25, 
    5224.75,
  5223.088, 5234.341, 5244.505, 5255.168, 5264.914, 5273.135, 5280.833, 
    5284.704, 5287.8, 5287.855, 5286.32, 5285.467, 5277.979, 5262.88, 5242.982,
  5215.365, 5226.282, 5236.184, 5246.496, 5256.751, 5267.151, 5274.681, 
    5282.98, 5286.344, 5285.33, 5285.919, 5288.358, 5284.211, 5272.805, 
    5257.274,
  5208.197, 5218.368, 5227.299, 5237.239, 5246.843, 5258.285, 5268.209, 
    5275.191, 5280.447, 5282.688, 5283.761, 5288.683, 5288.849, 5282.636, 
    5270.78,
  5203.366, 5212.855, 5221.81, 5231.834, 5242.805, 5253.646, 5263.269, 
    5271.636, 5275.877, 5276.535, 5278.865, 5286.035, 5289.636, 5286.758, 
    5279.196,
  5203.491, 5211.044, 5218.999, 5228.037, 5238.06, 5248.763, 5258.043, 
    5264.233, 5268.178, 5270.687, 5274.191, 5282.211, 5287.81, 5288.456, 
    5284.163,
  5249.843, 5262.465, 5273.87, 5280.917, 5286.406, 5287.833, 5285.498, 
    5281.08, 5274.612, 5265.375, 5254.438, 5240.072, 5223.165, 5203.435, 
    5182.851,
  5257.386, 5268.612, 5278.341, 5284.423, 5288.618, 5290.567, 5291.464, 
    5285.134, 5278.958, 5273.957, 5265.377, 5254.501, 5238.778, 5223.438, 
    5203.328,
  5261.681, 5271.672, 5280.183, 5286.549, 5290.86, 5293.722, 5292.104, 
    5292.554, 5286.956, 5280.917, 5273.979, 5265.333, 5253.327, 5238.332, 
    5220.104,
  5265.013, 5272.916, 5280.274, 5285.881, 5289.485, 5293.253, 5293.625, 
    5289.188, 5284.924, 5285.052, 5280.288, 5273.648, 5264.075, 5252.712, 
    5236.466,
  5266.04, 5272.431, 5277.875, 5283.208, 5288.002, 5290.345, 5291.59, 
    5292.044, 5291.055, 5284.935, 5284.34, 5278.725, 5272.265, 5261.616, 
    5249.028,
  5265.087, 5269.762, 5273.923, 5277.268, 5281.295, 5284.855, 5286.717, 
    5285.57, 5284.653, 5283.909, 5284.239, 5282.19, 5277.583, 5270.851, 
    5260.545,
  5260.104, 5263.78, 5266.766, 5269.806, 5273.014, 5276.939, 5279.845, 
    5282.21, 5282.279, 5281.468, 5280.666, 5281.438, 5279.41, 5275.035, 
    5267.687,
  5251.095, 5254.042, 5256.635, 5259.331, 5261.796, 5265.104, 5269.352, 
    5271.485, 5273.175, 5275.083, 5275.451, 5277.851, 5279.462, 5278.201, 
    5274.269,
  5237.33, 5240.332, 5243.367, 5246.604, 5249.706, 5253.264, 5256.766, 
    5261.171, 5264.501, 5266.571, 5267.986, 5270.778, 5274.527, 5276.711, 
    5275.671,
  5223.299, 5225.555, 5228.62, 5231.765, 5234.328, 5237.743, 5241.48, 
    5245.518, 5250.028, 5255.177, 5258.867, 5261.993, 5267.755, 5273.376, 
    5275.691,
  5230.404, 5243.575, 5255.063, 5262.056, 5266.922, 5267.575, 5264.476, 
    5260.01, 5252.032, 5238.927, 5223.808, 5203.75, 5178.957, 5144.257, 
    5105.12,
  5243.954, 5255.89, 5265.736, 5271.428, 5274.795, 5273.187, 5271.795, 
    5263.397, 5253.788, 5243.789, 5228.844, 5211.086, 5186.249, 5156.041, 
    5117.616,
  5254.946, 5266.055, 5273.957, 5279.56, 5280.323, 5281.69, 5274.765, 
    5271.599, 5261.528, 5249.104, 5234.337, 5218.042, 5195.751, 5167.114, 
    5131.293,
  5264.501, 5272.295, 5278.662, 5282.755, 5284.705, 5282.484, 5279.51, 
    5270.829, 5260.393, 5251.915, 5239.11, 5224.241, 5205.673, 5181.847, 
    5149.819,
  5269.225, 5276.06, 5281.249, 5285.154, 5286.554, 5285.393, 5279.236, 
    5273.664, 5266.013, 5253.385, 5243.172, 5229.994, 5215.249, 5194.334, 
    5168.819,
  5272.328, 5277.868, 5281.47, 5284.384, 5283.585, 5281.51, 5276.477, 
    5268.299, 5259.315, 5252.089, 5243.99, 5234.518, 5223.216, 5209.158, 
    5189.492,
  5271.87, 5276.634, 5279.029, 5280.222, 5278.688, 5274.725, 5268.555, 
    5262.886, 5256.095, 5249.037, 5242.571, 5236.311, 5228.175, 5219.346, 
    5206.267,
  5270.124, 5272.065, 5272.264, 5271.16, 5267.238, 5262.519, 5256.353, 
    5249.937, 5243.675, 5239.693, 5236.817, 5234.186, 5230.928, 5226.879, 
    5220.396,
  5262.498, 5262.459, 5260.834, 5257.464, 5252.567, 5246.77, 5239.814, 
    5234.562, 5230.734, 5228.041, 5227.717, 5228.291, 5228.413, 5228.586, 
    5227.87,
  5250.296, 5246.404, 5241.75, 5237.071, 5230.811, 5225.419, 5220.595, 
    5216.823, 5214.113, 5213.78, 5214.985, 5218.611, 5222.401, 5226.681, 
    5231.1,
  5222.274, 5234.953, 5245.081, 5250.515, 5252.183, 5247.919, 5237.128, 
    5223.309, 5204.506, 5180.521, 5156.657, 5131.463, 5110.468, 5093.508, 
    5081.869,
  5235.162, 5246.94, 5256.185, 5260.949, 5261.344, 5255.113, 5246.755, 
    5228.175, 5208.709, 5190.274, 5169.125, 5147.171, 5126.549, 5112.619, 
    5102.437,
  5245.717, 5257.933, 5265.455, 5270.227, 5267.675, 5265.193, 5250.652, 
    5240.905, 5221.751, 5200.412, 5181.572, 5162.358, 5144.318, 5131.272, 
    5122.172,
  5255.834, 5266.132, 5272.458, 5275.31, 5274.72, 5266.23, 5258.266, 5238.84, 
    5221.31, 5206.992, 5192.018, 5176.338, 5161.025, 5149.257, 5142.932,
  5263.529, 5271.776, 5276.902, 5278.54, 5276.057, 5270.814, 5257.029, 
    5247.026, 5230.775, 5210.683, 5200.105, 5187.93, 5176.647, 5166.194, 
    5161.545,
  5268.829, 5275.124, 5277.886, 5278.572, 5274.548, 5267.062, 5256.038, 
    5238.822, 5222.29, 5211.791, 5204.07, 5197.014, 5188.88, 5181.646, 
    5178.469,
  5270.641, 5275.639, 5276.544, 5275.045, 5269.839, 5261.163, 5248.534, 
    5236.328, 5222.651, 5209.274, 5204.781, 5202.668, 5198.036, 5193.662, 
    5191.778,
  5269.952, 5272.006, 5270.795, 5267.774, 5260.67, 5251.322, 5238.916, 
    5224.552, 5210.896, 5203.725, 5202.7, 5204.753, 5204.977, 5203.439, 
    5204.232,
  5264.199, 5265.038, 5262.499, 5257.749, 5250.084, 5240.093, 5228.963, 
    5218.546, 5208.621, 5201.071, 5199.656, 5203.994, 5208.402, 5210.1, 
    5212.85,
  5255.861, 5254.3, 5250.144, 5245.59, 5238.142, 5230.783, 5222.93, 5213.558, 
    5204.57, 5199.004, 5197.291, 5202.19, 5208.414, 5213.464, 5218.468,
  5277.063, 5281.623, 5281.402, 5273.778, 5261.999, 5245.187, 5224.044, 
    5206.8, 5191.819, 5178.229, 5167.671, 5157.44, 5145.125, 5129.858, 
    5110.511,
  5283.711, 5288.588, 5287.582, 5281.045, 5269.045, 5249.729, 5235.595, 
    5211.227, 5193.445, 5183.919, 5174.413, 5165.69, 5154.127, 5140.584, 
    5122.132,
  5287.635, 5293.384, 5291.784, 5287.407, 5273.435, 5262.165, 5235.423, 
    5224.444, 5202.303, 5188.406, 5179.872, 5172.238, 5162.742, 5149.415, 
    5131.572,
  5290.22, 5295.183, 5294.816, 5289.693, 5279.297, 5260.547, 5247.322, 
    5222.165, 5204.003, 5190.932, 5183.684, 5176.924, 5169.633, 5159.382, 
    5143.321,
  5289.838, 5294.816, 5295.489, 5290.607, 5281.036, 5266.566, 5246.492, 
    5231.908, 5212.235, 5193.41, 5187.139, 5180.228, 5175.864, 5166.357, 
    5154.135,
  5287.228, 5292.712, 5293.447, 5289.764, 5279.272, 5265.126, 5249.59, 
    5230.333, 5211.146, 5197.455, 5189.414, 5182.762, 5180.04, 5174.433, 
    5165.018,
  5282.541, 5288.575, 5290.087, 5285.757, 5276.98, 5263.5, 5248.732, 5235.03, 
    5218.262, 5201.374, 5191.637, 5185.256, 5182.015, 5179.761, 5173.471,
  5277.21, 5282.81, 5284.044, 5279.927, 5270.523, 5258.872, 5247.412, 
    5233.127, 5217.542, 5203.209, 5193.06, 5186.591, 5183.612, 5183.452, 
    5181.321,
  5270.13, 5275.657, 5276.276, 5271.519, 5264.11, 5254.306, 5244.609, 
    5233.516, 5219.706, 5203.979, 5192.104, 5186.55, 5183.397, 5183.71, 
    5185.259,
  5263.209, 5266.496, 5265.813, 5261.985, 5254.349, 5247.114, 5238.283, 
    5225.708, 5212.393, 5200.115, 5189.35, 5184.226, 5182.164, 5182.617, 
    5186.999,
  5297.39, 5299.072, 5298.632, 5292.287, 5283.429, 5269.472, 5251.694, 
    5233.711, 5211.77, 5183.736, 5160.298, 5135.355, 5109.747, 5078.981, 
    5044.902,
  5292.872, 5295.721, 5295.68, 5291.195, 5283.158, 5267.958, 5256.326, 
    5230.514, 5208.009, 5186.792, 5162.396, 5136.788, 5109.464, 5080.505, 
    5044.776,
  5286.226, 5290.632, 5291.215, 5289.374, 5280.313, 5272.289, 5250.681, 
    5241.168, 5216.673, 5190.192, 5163.976, 5139.023, 5109.967, 5080.557, 
    5045.886,
  5279, 5283.245, 5284.94, 5283.233, 5277.321, 5264.646, 5254.709, 5230.601, 
    5211.128, 5193.036, 5165.814, 5140.262, 5112.07, 5084.418, 5051.19,
  5269.542, 5274.105, 5277.063, 5275.768, 5271.462, 5262.255, 5246.728, 
    5236.124, 5217.154, 5190.188, 5168.38, 5140.831, 5114.774, 5086.499, 
    5058.025,
  5259.606, 5263.637, 5265.977, 5265.659, 5260.8, 5252.811, 5241.84, 
    5223.377, 5206.114, 5189.341, 5167.309, 5142.13, 5117.213, 5092.311, 
    5066.38,
  5248.89, 5252.48, 5254.4, 5253.74, 5250.252, 5242.373, 5231.247, 5220.579, 
    5205.156, 5185.086, 5164.707, 5142.494, 5118.422, 5096.526, 5074.36,
  5239.938, 5241.177, 5241.049, 5240.421, 5235.396, 5228.815, 5219.092, 
    5205.978, 5191.792, 5177.982, 5160.158, 5140.05, 5119.759, 5101.509, 
    5084.487,
  5233.479, 5233.583, 5232.134, 5228.731, 5223.66, 5216.211, 5206.226, 
    5197.088, 5185.127, 5169.857, 5153.391, 5135.851, 5118.723, 5104.191, 
    5092.696,
  5232.644, 5228.138, 5223.251, 5218.662, 5210.997, 5201.925, 5192.3, 
    5180.915, 5169.313, 5158.424, 5144.38, 5128.977, 5115.912, 5106.584, 
    5101.105,
  5281.218, 5276.957, 5274.274, 5270.771, 5266.627, 5259.299, 5248.202, 
    5238.133, 5223.783, 5202.497, 5181.308, 5158.146, 5131.968, 5102.703, 
    5069.742,
  5272.461, 5268.619, 5265.436, 5260.644, 5254.925, 5245.54, 5239.006, 
    5220.961, 5206.686, 5193.804, 5172.432, 5150.396, 5124.207, 5099.736, 
    5063.798,
  5267.511, 5262.524, 5257.912, 5253.106, 5243.796, 5239.299, 5222.366, 
    5220.728, 5200.69, 5181.929, 5161.979, 5143.215, 5117.719, 5092.61, 
    5058.345,
  5263.383, 5256.81, 5250.697, 5243.867, 5236.521, 5224.765, 5219.056, 
    5197.066, 5186.51, 5173.692, 5152.502, 5134.622, 5112.194, 5088.606, 
    5055.298,
  5262.564, 5255.016, 5246.985, 5238.883, 5229.905, 5220.016, 5204.919, 
    5197.09, 5179.415, 5159.204, 5144.983, 5125.576, 5106.584, 5081.614, 
    5052.418,
  5264.369, 5254.986, 5244.132, 5234.44, 5221.906, 5210.218, 5196.701, 
    5177.756, 5162.499, 5149.641, 5132.457, 5116.648, 5098.705, 5077.008, 
    5049.225,
  5268.796, 5257.954, 5244.544, 5231.674, 5217.217, 5202.194, 5185.033, 
    5170.617, 5152.3, 5133.606, 5119.204, 5105.373, 5088.984, 5069.81, 5044.12,
  5272.726, 5258.862, 5242.577, 5227.142, 5208.681, 5191.682, 5171.856, 
    5151.656, 5132.134, 5117.073, 5102.187, 5090.486, 5077.882, 5062.541, 
    5040.222,
  5274.462, 5259.167, 5241.364, 5222.172, 5202.023, 5180.682, 5157.664, 
    5137.049, 5116.004, 5096.752, 5083.736, 5075.108, 5065.598, 5053.549, 
    5035.061,
  5272.007, 5252.312, 5232.415, 5211.758, 5187.965, 5164.478, 5139.969, 
    5114.888, 5093.181, 5077.172, 5066.243, 5059.666, 5053.277, 5044.931, 
    5030.801,
  5247.519, 5243.82, 5241.659, 5239.821, 5239.079, 5237.379, 5234.385, 
    5231.862, 5225.039, 5212.034, 5198.766, 5183.333, 5166.209, 5144.132, 
    5123.599,
  5251.107, 5246.157, 5243.507, 5240.976, 5239.461, 5235.875, 5234.764, 
    5224.654, 5216.943, 5209.376, 5193.226, 5175.771, 5154.658, 5134.603, 
    5110.349,
  5259.21, 5252.996, 5248.687, 5245.955, 5240.372, 5239.743, 5230.691, 
    5230.104, 5216.322, 5199.78, 5182.489, 5163.92, 5139.253, 5117.428, 
    5096.805,
  5266.31, 5259.05, 5253.973, 5248.732, 5245.336, 5236.464, 5233.163, 
    5216.752, 5206.383, 5195.471, 5170.09, 5146.867, 5121.932, 5099.578, 
    5083.744,
  5269.522, 5262.181, 5256.215, 5250.339, 5243.911, 5237.795, 5226.575, 
    5218.441, 5201.068, 5176.838, 5156.534, 5127.25, 5101.733, 5080.917, 
    5072.199,
  5265.218, 5258.143, 5252.126, 5246.533, 5239.203, 5230.821, 5219.742, 
    5204.613, 5186.06, 5165.899, 5137.382, 5108.891, 5081.611, 5067.738, 
    5063.258,
  5252.57, 5246.414, 5240.538, 5236.088, 5229.361, 5221.482, 5209.789, 
    5196.205, 5174.534, 5148.68, 5120.003, 5091.396, 5064.733, 5057.265, 
    5056.452,
  5234.598, 5228.083, 5222.224, 5219.892, 5213.878, 5207.544, 5194.776, 
    5179.185, 5158.178, 5136.101, 5105.225, 5076.898, 5054.043, 5051.324, 
    5053.683,
  5212.994, 5206.74, 5202.032, 5199.809, 5195.553, 5190.158, 5179.574, 
    5166.917, 5145.985, 5121.709, 5092.551, 5067.386, 5048.121, 5048.847, 
    5052.994,
  5191.191, 5183.183, 5178.706, 5177.079, 5174.043, 5169.965, 5161.11, 
    5148.43, 5130.38, 5109.844, 5083.407, 5061.424, 5047.13, 5049.788, 
    5053.629,
  5228.762, 5219.91, 5213.69, 5211.3, 5213.462, 5218.079, 5224.466, 5231.421, 
    5235.199, 5235.623, 5232.128, 5223.748, 5206.036, 5181.104, 5152.628,
  5229.608, 5221.052, 5215.69, 5212.356, 5211.71, 5215.639, 5221.391, 
    5225.83, 5229.629, 5232.643, 5226.058, 5217.139, 5196.6, 5172.952, 
    5137.749,
  5227.065, 5218.874, 5214.09, 5212.243, 5211.686, 5214.812, 5217.337, 
    5225.177, 5226.033, 5226.406, 5220.982, 5210.574, 5189.185, 5162.202, 
    5127.738,
  5216.752, 5208.862, 5204.678, 5203.743, 5205.179, 5206.741, 5212.173, 
    5211.077, 5218.542, 5218.343, 5213.337, 5202.43, 5182.8, 5156.345, 
    5123.846,
  5203.173, 5194.98, 5190.111, 5189.403, 5190.688, 5195.117, 5197.625, 
    5208.263, 5206.115, 5209.026, 5205.805, 5195.01, 5176.832, 5151.26, 
    5124.383,
  5188.243, 5177.935, 5170.313, 5168.432, 5168.362, 5172.822, 5179.837, 
    5183.616, 5192.658, 5196.154, 5193.617, 5186.845, 5171.25, 5149.233, 
    5126.139,
  5171.63, 5159.516, 5149.083, 5143.214, 5141.838, 5145.695, 5153.285, 
    5166.147, 5173.439, 5178.054, 5182.85, 5177.446, 5164.878, 5145.789, 
    5127.722,
  5153.96, 5137.848, 5122.715, 5114.1, 5109.513, 5113.082, 5121.546, 
    5132.843, 5147.247, 5160.629, 5166.372, 5165.381, 5158.175, 5142.865, 
    5128.719,
  5135.67, 5116.436, 5097.573, 5083.996, 5078.051, 5080.161, 5089.489, 
    5105.419, 5122.504, 5136.574, 5148.712, 5152.862, 5149.349, 5138.014, 
    5128.041,
  5121.864, 5096.868, 5073.785, 5060.333, 5054.359, 5055.15, 5063.233, 
    5076.412, 5096.176, 5116.088, 5131.388, 5138.76, 5140.424, 5132.794, 
    5126.378,
  5180.27, 5180.952, 5177.129, 5172.559, 5172.58, 5183.149, 5197.637, 
    5215.868, 5234.411, 5249.079, 5256.522, 5258.363, 5248.831, 5232.56, 
    5209.271,
  5172.116, 5177.03, 5176.242, 5174.681, 5172.105, 5181.821, 5195.746, 
    5213.041, 5229.958, 5247.419, 5254.252, 5257.508, 5247.605, 5236.352, 
    5212.226,
  5163.067, 5170.188, 5174.845, 5175.475, 5176.394, 5183.038, 5194.028, 
    5212.845, 5228.185, 5242.538, 5250.741, 5254.949, 5247.507, 5237.188, 
    5215.702,
  5151.46, 5158.931, 5166.773, 5171.909, 5177.58, 5180.779, 5192.875, 
    5200.865, 5219.801, 5234.077, 5244.963, 5249.585, 5246.373, 5238.924, 
    5220.384,
  5141.406, 5148.624, 5157.063, 5166.109, 5172.664, 5182.106, 5185.215, 
    5201.23, 5211.072, 5224.196, 5235.685, 5242.732, 5243.077, 5238.763, 
    5223.982,
  5130.844, 5137.687, 5145.703, 5155.798, 5164.518, 5172.625, 5182.724, 
    5189.285, 5200.297, 5214.075, 5222.927, 5233.956, 5237.591, 5238.259, 
    5227.188,
  5122.014, 5125.957, 5134.124, 5143.4, 5152.982, 5163.23, 5171.183, 
    5183.637, 5193.224, 5201.085, 5213.605, 5223.829, 5231.504, 5235.808, 
    5228.955,
  5117.701, 5115.094, 5119.305, 5129.424, 5136.968, 5146.696, 5155.675, 
    5164.331, 5175.485, 5189.914, 5201.139, 5212.643, 5224.438, 5232.405, 
    5230.726,
  5123.647, 5114.233, 5110.288, 5113.506, 5119.581, 5126.924, 5135.297, 
    5147.269, 5159.206, 5171.83, 5186.891, 5202.541, 5216.249, 5227.68, 
    5230.945,
  5136.955, 5121.29, 5111.661, 5107.243, 5105.218, 5107.121, 5111.968, 
    5118.871, 5131.402, 5150.116, 5170.308, 5189.357, 5207.038, 5222.521, 
    5230.135,
  5166.443, 5176.715, 5178.353, 5176.41, 5182.771, 5194.721, 5212.447, 
    5231.94, 5248.074, 5257.18, 5259.762, 5260.392, 5259.748, 5260.354, 
    5263.69,
  5163.791, 5175.647, 5177.819, 5176.208, 5179.634, 5194.903, 5214.743, 
    5233.191, 5249.041, 5262.979, 5267.715, 5269.73, 5269.513, 5271.801, 
    5275.119,
  5161.693, 5174.913, 5179.393, 5177.432, 5181.781, 5198.221, 5216.36, 5240, 
    5258.969, 5269.481, 5275.254, 5278.048, 5279.882, 5281.311, 5284.94,
  5159.071, 5172.783, 5180.298, 5179.492, 5187.15, 5196.544, 5224.451, 
    5237.845, 5258.786, 5271.999, 5281.903, 5284.327, 5287.055, 5289.771, 
    5293.886,
  5156.231, 5171.868, 5180.165, 5185.262, 5188.144, 5209.114, 5220.508, 
    5249.346, 5264.931, 5276.845, 5284.965, 5289.966, 5292.989, 5295.799, 
    5299.789,
  5154.062, 5170.16, 5179.967, 5187.712, 5193.326, 5205.876, 5229.537, 
    5243.235, 5259.282, 5278.263, 5285.14, 5292.569, 5294.583, 5300.783, 
    5303.697,
  5152.873, 5168.857, 5180.624, 5189.705, 5197.927, 5211.417, 5225.943, 
    5248.038, 5265, 5275.157, 5285.994, 5292.283, 5296.893, 5303.112, 5306.25,
  5152.22, 5166.289, 5177.784, 5189.44, 5197.204, 5210.453, 5225.708, 
    5238.613, 5252.886, 5270.271, 5281.322, 5289.789, 5296.69, 5304.356, 
    5308.57,
  5153.568, 5164.005, 5174.582, 5186.144, 5196.617, 5207.729, 5220.825, 
    5237.843, 5251.744, 5263.511, 5274.599, 5287.031, 5295.427, 5305.14, 
    5310.016,
  5158.061, 5160.572, 5166.67, 5176.67, 5187.219, 5199.875, 5212.606, 
    5225.595, 5238.556, 5255.227, 5269.112, 5282.754, 5293.333, 5305.479, 
    5311.778,
  5179.295, 5188.037, 5196.963, 5208.076, 5218.706, 5228.229, 5237.067, 
    5247.824, 5260.752, 5272.379, 5284.86, 5297.944, 5307.689, 5316.051, 
    5320.374,
  5185.59, 5194.024, 5203.247, 5214.847, 5224.227, 5234.959, 5246.198, 
    5256.984, 5268.495, 5284.483, 5298.092, 5311.296, 5320.621, 5328.816, 
    5333.195,
  5193.289, 5202.824, 5213.074, 5224.759, 5233.691, 5247.035, 5254.564, 
    5269.806, 5284.804, 5296.701, 5310.554, 5322.482, 5332.851, 5339.699, 
    5344.627,
  5203.27, 5212.369, 5222.948, 5231.547, 5246.359, 5250.931, 5269.289, 
    5276.313, 5291.164, 5306.269, 5320.969, 5331.632, 5342.029, 5348.989, 
    5354.71,
  5212.955, 5222.152, 5230.84, 5241.187, 5250.793, 5269.097, 5276.354, 
    5293.407, 5308.586, 5316.949, 5330.298, 5339.981, 5350.303, 5356.374, 
    5362.861,
  5222.059, 5230.933, 5236.054, 5246.409, 5259.292, 5274.052, 5293.525, 
    5302.729, 5312.585, 5327.398, 5337.792, 5347.687, 5356.513, 5363.904, 
    5370.292,
  5229.751, 5238.742, 5244.224, 5252.589, 5268.949, 5288.342, 5300.837, 
    5317.776, 5330.879, 5338.196, 5346.577, 5354.77, 5363.08, 5370.14, 
    5376.742,
  5237.109, 5245.096, 5250.399, 5259.516, 5275.738, 5296.598, 5313.774, 
    5325.61, 5334.976, 5345.603, 5353.358, 5360.771, 5368.437, 5375.666, 
    5382.921,
  5241.519, 5251.522, 5260.001, 5270.45, 5287.793, 5306.995, 5323.088, 
    5338.366, 5348.753, 5354.489, 5360.06, 5366.498, 5372.841, 5380.207, 
    5387.645,
  5245.331, 5256.347, 5265.812, 5278.788, 5296.194, 5316.149, 5332.591, 
    5343.944, 5351.257, 5358.526, 5364.104, 5370.071, 5376.392, 5384.041, 
    5392.186,
  5240.112, 5251.866, 5264.082, 5275.493, 5283.355, 5290.862, 5301.363, 
    5313.294, 5322.33, 5326.989, 5330.083, 5333.201, 5335, 5336.209, 5336.493,
  5236.513, 5250.23, 5264.1, 5277.718, 5284.743, 5296.09, 5311.351, 5324.758, 
    5333.318, 5343.018, 5348.009, 5352.631, 5354.023, 5356.1, 5356.787,
  5234.443, 5250.496, 5266.021, 5280.355, 5288.604, 5305.362, 5319.176, 
    5337.038, 5350.112, 5357.908, 5364.211, 5368.78, 5372.472, 5374.412, 
    5375.841,
  5235.08, 5251.203, 5269.1, 5280.727, 5297.417, 5307.25, 5332.784, 5343.915, 
    5359.016, 5369.288, 5378.347, 5382.692, 5387.702, 5390.472, 5394.226,
  5237.257, 5254.351, 5272.229, 5286.388, 5300.442, 5324.022, 5338.823, 
    5358.505, 5374.094, 5380.539, 5389.783, 5394.105, 5400.648, 5403.901, 
    5409.159,
  5242.277, 5259.454, 5274.413, 5290.629, 5307.614, 5327.57, 5353.244, 
    5365.849, 5378.468, 5390.997, 5397.628, 5403.643, 5409.771, 5415.724, 
    5422.324,
  5249.745, 5266.83, 5281.612, 5296.715, 5316.872, 5340.938, 5358.766, 
    5378.417, 5392.387, 5398.752, 5404.36, 5410.429, 5417.031, 5424.607, 
    5432.078,
  5258.803, 5274.22, 5288.839, 5306.271, 5325.439, 5348.852, 5369.22, 
    5383.07, 5393.34, 5402.842, 5409.252, 5415.251, 5422.207, 5430.904, 
    5440.074,
  5268.702, 5284.815, 5301.382, 5319.617, 5340.57, 5360.002, 5376.014, 
    5391.396, 5401.668, 5407.854, 5413.308, 5419.499, 5426.138, 5434.861, 
    5444.638,
  5280.459, 5296.537, 5314.03, 5333.296, 5352.585, 5370.551, 5384.717, 
    5394.314, 5401.911, 5409.703, 5416.377, 5422.738, 5429.174, 5437.596, 
    5447.791,
  5330.029, 5328.655, 5329.221, 5330.101, 5331.757, 5333.585, 5333.157, 
    5333.634, 5335.52, 5335.011, 5334.288, 5334.414, 5335.211, 5336.735, 
    5340.983,
  5336.923, 5337.289, 5339.112, 5342.858, 5346.072, 5347.898, 5351.479, 
    5353.715, 5352.224, 5353.489, 5351.961, 5351.56, 5349.957, 5351.81, 
    5356.164,
  5342.023, 5344.667, 5348.456, 5354.995, 5357.811, 5365.524, 5365.351, 
    5369.693, 5371.817, 5372.119, 5369.882, 5368, 5366.219, 5366.896, 5371.729,
  5345.73, 5348.854, 5356.612, 5362.163, 5372.425, 5374.582, 5382.62, 
    5385.477, 5387.398, 5388.186, 5388.392, 5384.527, 5383.495, 5384.616, 
    5392.208,
  5347.36, 5352.423, 5362.476, 5370.391, 5380.179, 5389.116, 5395.848, 
    5397.672, 5406.145, 5404.476, 5406.557, 5402.805, 5403.725, 5403.664, 
    5413.415,
  5346.623, 5354.695, 5364.813, 5375.607, 5387.092, 5396.442, 5406.806, 
    5413.74, 5416.429, 5420.37, 5422.393, 5422.06, 5422.988, 5425.92, 5434.16,
  5345.283, 5357.011, 5368.963, 5379.761, 5391.521, 5405.554, 5414.025, 
    5422.73, 5429.842, 5433.597, 5436.202, 5439.635, 5441.58, 5445.903, 
    5452.587,
  5343.806, 5357.442, 5370.459, 5382.831, 5394.913, 5408.944, 5421.311, 
    5431.363, 5436.557, 5442.243, 5447.418, 5452.591, 5457.292, 5462.771, 
    5469.189,
  5342.451, 5358.555, 5374.188, 5385.908, 5399.655, 5414.915, 5426.225, 
    5436.55, 5443.604, 5448.923, 5454.276, 5461.466, 5468.219, 5474.778, 
    5480.816,
  5340.567, 5357.616, 5373.945, 5387.463, 5402.642, 5418.813, 5432.26, 
    5441.774, 5446.193, 5451.213, 5457.654, 5465.47, 5473.582, 5482.157, 
    5489.213,
  5308.567, 5307.993, 5307.438, 5307.585, 5309.482, 5313.463, 5317.985, 
    5327.013, 5338.665, 5351.071, 5365.227, 5381.955, 5399.473, 5417.17, 
    5435.825,
  5321.622, 5322.442, 5322.452, 5323.44, 5324.514, 5326.498, 5332.784, 
    5339.43, 5348.021, 5362.765, 5377.605, 5396.707, 5414.904, 5436.91, 
    5455.023,
  5334.289, 5336.895, 5338.073, 5340.308, 5339.268, 5344.305, 5343.555, 
    5352.897, 5362.213, 5373.564, 5388.402, 5407.927, 5429.651, 5450.845, 
    5471.807,
  5346.87, 5350.065, 5353.643, 5353.938, 5357.297, 5353.641, 5359.184, 
    5359.632, 5366.71, 5379.569, 5396.732, 5416.889, 5441.496, 5465.637, 
    5487.698,
  5357.767, 5362.441, 5366.782, 5368.811, 5369.064, 5369.877, 5367.244, 
    5369.167, 5379.556, 5386.07, 5404.372, 5425.492, 5451.871, 5475.622, 
    5499.106,
  5367.805, 5374.092, 5378.4, 5381.888, 5381.823, 5379.473, 5379.174, 
    5378.653, 5380.857, 5395.732, 5412.343, 5435.769, 5461.423, 5487.547, 
    5509.473,
  5377.488, 5384.912, 5390.311, 5394.323, 5394.386, 5393.051, 5388.564, 
    5390.494, 5397.036, 5407.072, 5424.179, 5447.502, 5472.343, 5496.925, 
    5517.183,
  5386.709, 5394.104, 5400.108, 5405.257, 5406.381, 5405.174, 5403.431, 
    5403.086, 5406.742, 5419.931, 5438.236, 5460.414, 5484.071, 5506.762, 
    5524.926,
  5395.051, 5402.467, 5409.819, 5414.958, 5418.354, 5418.758, 5417.303, 
    5419.547, 5426.205, 5437.423, 5453.627, 5474.75, 5495.691, 5514.86, 
    5530.265,
  5401.742, 5408.901, 5416.579, 5422.427, 5427.395, 5430.342, 5432.068, 
    5434.104, 5439.867, 5452.176, 5468.638, 5487.137, 5505.513, 5522.314, 
    5534.759,
  5279.298, 5286.591, 5295.213, 5304.855, 5315.617, 5326.273, 5337.517, 
    5352.788, 5369.523, 5386.384, 5406.951, 5429.469, 5450.629, 5468.962, 
    5483.907,
  5290.241, 5297.826, 5306.131, 5316.768, 5326.522, 5337.798, 5353.895, 
    5368.445, 5385.037, 5409.106, 5431.485, 5455.73, 5474.913, 5492.955, 
    5505.776,
  5300.778, 5308.389, 5316.995, 5327.911, 5338.501, 5354.867, 5366.698, 
    5389.9, 5411.064, 5431.578, 5454.819, 5476.716, 5497.129, 5513.335, 
    5526.355,
  5311.77, 5318.31, 5328.252, 5336.947, 5352.915, 5361.221, 5386.413, 
    5398.915, 5422.468, 5448.724, 5473.572, 5495.023, 5515.861, 5531.625, 
    5542.831,
  5321.357, 5328.214, 5336.522, 5347.285, 5359.413, 5379.025, 5392.147, 
    5419.135, 5446.651, 5463.857, 5490.148, 5510.621, 5531.746, 5544.808, 
    5554.775,
  5330.958, 5337.195, 5343.128, 5353.465, 5365.763, 5381.445, 5405.524, 
    5424.273, 5447.057, 5478.646, 5501.419, 5524.323, 5543.007, 5556.592, 
    5563.439,
  5339.724, 5345.233, 5349.833, 5357.494, 5369.478, 5387.817, 5407.645, 
    5437.146, 5465.805, 5488.639, 5512.11, 5535.009, 5552.277, 5563.932, 
    5568.299,
  5349.897, 5353.183, 5355.746, 5361.493, 5369.593, 5386.55, 5411.099, 
    5435.627, 5462.479, 5493.392, 5519.265, 5541.524, 5558.438, 5568.862, 
    5571.742,
  5358.354, 5360.707, 5362.258, 5364.297, 5371.978, 5386.664, 5409.852, 
    5441.017, 5472.232, 5499.225, 5523.901, 5546.3, 5562.116, 5571.437, 
    5572.851,
  5365.575, 5366.852, 5367.214, 5367.032, 5371.168, 5385.274, 5409.361, 
    5437.675, 5468.193, 5499.396, 5526.64, 5548.671, 5564.164, 5572.535, 
    5573.733,
  5267.594, 5276.451, 5291.233, 5307.388, 5324.418, 5340.968, 5359.341, 
    5381.324, 5401.738, 5416.643, 5428.011, 5434.999, 5438.333, 5437.896, 
    5435.721,
  5275.511, 5283.5, 5296.978, 5313.73, 5328.585, 5346.414, 5369.282, 5390.49, 
    5411.058, 5432.181, 5443.959, 5452.105, 5453.753, 5453.732, 5450.938,
  5283.536, 5290.836, 5304.417, 5319.723, 5335.135, 5357.65, 5376.131, 
    5406.996, 5431.454, 5447.36, 5460.412, 5467.635, 5471.774, 5472.293, 
    5469.496,
  5291.305, 5298.598, 5311.652, 5324.512, 5344.465, 5357.863, 5392.897, 
    5411.026, 5438.492, 5460.639, 5475.711, 5483.43, 5488.941, 5489.429, 
    5490.085,
  5297.763, 5306.581, 5318.375, 5333.336, 5350.507, 5375.771, 5395.269, 
    5432.418, 5459.878, 5473.514, 5490.138, 5498.337, 5506.028, 5506.096, 
    5507.668,
  5303.944, 5313.674, 5324.489, 5339.671, 5357.611, 5378.525, 5411.629, 
    5434.645, 5460.386, 5487.373, 5501.825, 5513.129, 5519.083, 5522.421, 
    5523.543,
  5309.023, 5319.813, 5331.614, 5346.353, 5365.771, 5389.62, 5415.309, 
    5450.115, 5478.714, 5497.099, 5513.14, 5525.206, 5531.614, 5535.015, 
    5536.508,
  5313.595, 5324.687, 5336.052, 5351.188, 5368.278, 5392.532, 5422.557, 
    5449.264, 5475.316, 5502.05, 5520.532, 5533.356, 5541.278, 5545.411, 
    5547.707,
  5316.633, 5328.192, 5341.01, 5356.257, 5374.795, 5396.298, 5423.092, 
    5455.85, 5484.15, 5506.315, 5524.985, 5539.633, 5548.052, 5552.74, 
    5555.098,
  5319.625, 5329.859, 5341.792, 5355.881, 5372.961, 5395.261, 5421.981, 
    5449.811, 5476.74, 5504.114, 5526.209, 5542.617, 5552.357, 5557.637, 
    5560.056,
  5266.047, 5278.92, 5288.533, 5298.713, 5306.675, 5313.591, 5316.041, 
    5318.034, 5319.972, 5323.182, 5330.02, 5341.613, 5355.23, 5369.658, 5384.3,
  5267.557, 5280.482, 5291.515, 5303.717, 5313.095, 5320.568, 5324.916, 
    5326.18, 5325.99, 5330.513, 5337.711, 5350.259, 5363.874, 5379.547, 
    5394.832,
  5267.414, 5279.264, 5293.084, 5306.955, 5318.073, 5328.539, 5330.912, 
    5332.137, 5333.003, 5336.849, 5345.302, 5357.495, 5373.334, 5389.187, 
    5406.329,
  5266.899, 5275.6, 5292.317, 5306.052, 5322.02, 5329.694, 5338.16, 5335.969, 
    5337.445, 5342.065, 5352.495, 5365.758, 5382.997, 5402.043, 5423.591,
  5265.997, 5271.859, 5288.975, 5305.292, 5322.662, 5336.672, 5341.896, 
    5342.662, 5344.891, 5348.913, 5360.91, 5374.864, 5394.573, 5413.375, 
    5439.604,
  5264.137, 5267.497, 5282.471, 5301.211, 5319.118, 5335.525, 5346.438, 
    5349.484, 5350.878, 5358.023, 5369.466, 5385.167, 5404.517, 5428.06, 
    5454.667,
  5260.84, 5264.266, 5276.868, 5296.403, 5316.358, 5335.993, 5348.606, 
    5354.566, 5359.708, 5365.931, 5378.211, 5395.128, 5415.048, 5438.091, 
    5465.533,
  5257.59, 5261.637, 5270.86, 5289.046, 5308.896, 5330.922, 5348.506, 
    5358.054, 5363.58, 5372.667, 5385.458, 5402.247, 5423.977, 5447.534, 
    5474.274,
  5254.709, 5260.125, 5268.471, 5284.555, 5303.938, 5326.502, 5345.818, 
    5358.887, 5368.574, 5377.904, 5390.924, 5408.042, 5428.95, 5452.46, 
    5477.618,
  5252.738, 5258.986, 5265.464, 5277.861, 5295.649, 5317.532, 5340.149, 
    5356.701, 5368.471, 5381.058, 5394.704, 5410.959, 5431.066, 5453.944, 
    5477.543,
  5315.11, 5305.102, 5296.673, 5290.034, 5282.746, 5276.529, 5273.621, 
    5278.057, 5288.293, 5301.558, 5317.27, 5335.545, 5353.518, 5370.298, 
    5387.093,
  5316.386, 5306.143, 5299.322, 5294.845, 5290.203, 5284.372, 5281.185, 
    5282.692, 5289.389, 5303.734, 5320.164, 5339.523, 5358.249, 5377.173, 
    5395.257,
  5314.812, 5305.37, 5299.357, 5296.13, 5293.706, 5291.028, 5286.496, 
    5287.333, 5294.051, 5304.95, 5321.521, 5341.313, 5361.592, 5379.846, 
    5400.049,
  5308.545, 5301.551, 5296.49, 5294.078, 5294.228, 5293.303, 5290.221, 
    5288.039, 5291.621, 5303.33, 5320.805, 5340.483, 5362.455, 5382.625, 
    5405.301,
  5297.498, 5293.989, 5290.899, 5289.62, 5291.249, 5293.444, 5292.755, 
    5289.767, 5293.519, 5301.607, 5318.707, 5337.851, 5360.853, 5380.226, 
    5404.683,
  5282.547, 5282.472, 5281.582, 5281.96, 5284.411, 5288.837, 5291.632, 
    5290.412, 5290.817, 5300.03, 5313.125, 5333.914, 5356.017, 5378.055, 
    5401.386,
  5265.353, 5268.775, 5269.842, 5271.857, 5275.326, 5281.321, 5286.404, 
    5289.06, 5289.715, 5295.269, 5307.595, 5327.072, 5348.475, 5371.033, 
    5393.526,
  5248.078, 5252.782, 5255.043, 5258.312, 5262.711, 5270.284, 5277.544, 
    5282.936, 5283.566, 5288.948, 5299.355, 5317.112, 5338.908, 5361.957, 
    5384.577,
  5230.706, 5236.289, 5240.538, 5243.718, 5248.211, 5256.474, 5265.475, 
    5273.77, 5278.261, 5281.491, 5290.077, 5306.157, 5326.317, 5349.349, 
    5371.682,
  5213.73, 5219.636, 5223.929, 5227.738, 5232.574, 5240.2, 5250.979, 
    5261.003, 5268.646, 5274.078, 5280.892, 5293.557, 5312.488, 5334.751, 
    5358.052,
  5292.804, 5293.843, 5291.066, 5281.473, 5269.601, 5261.586, 5267.482, 
    5283.483, 5300.159, 5311.08, 5319.597, 5326.917, 5337.375, 5349.74, 
    5363.941,
  5271.646, 5278.762, 5283.24, 5280.612, 5273.066, 5263.755, 5269.541, 
    5281.583, 5297.887, 5313.455, 5322.417, 5331.132, 5342.246, 5356.457, 
    5370.444,
  5248.181, 5261.614, 5272.478, 5277.269, 5273.951, 5270.307, 5267.346, 
    5282.214, 5296.663, 5310.869, 5322.502, 5331.778, 5344.171, 5357.964, 
    5374.042,
  5223.605, 5241.424, 5258.222, 5270.542, 5273.271, 5270.008, 5270.186, 
    5273.689, 5288.684, 5305.06, 5318.441, 5329.314, 5342.365, 5357.271, 
    5374.928,
  5199.188, 5220.884, 5242.029, 5261.943, 5271.124, 5272.38, 5270.337, 
    5273.564, 5283.64, 5295.431, 5311.097, 5323.337, 5337.171, 5351.141, 
    5369.95,
  5175.072, 5199.45, 5224.675, 5248.686, 5264.563, 5270.211, 5270.833, 
    5272.281, 5277.423, 5289.019, 5300.345, 5314.676, 5328.862, 5343.638, 
    5361.15,
  5153.899, 5181.171, 5209.324, 5236.54, 5256.955, 5268.207, 5270.815, 
    5273.671, 5278.222, 5282.678, 5291.566, 5303.025, 5316.86, 5332.238, 
    5347.796,
  5136.969, 5164.893, 5194.574, 5223.575, 5246.134, 5261.51, 5268.953, 
    5271.977, 5274.874, 5280.003, 5285.372, 5291.993, 5303.569, 5318.021, 
    5333.613,
  5125.116, 5153.555, 5184.333, 5213.907, 5237.42, 5253.978, 5263.562, 
    5269.84, 5273.451, 5276.237, 5279.509, 5284.533, 5290.289, 5302.093, 
    5315.891,
  5119.539, 5145.96, 5174.749, 5202.398, 5225.472, 5242.883, 5254.088, 
    5261.268, 5265.834, 5270.296, 5273.403, 5276.43, 5280.198, 5287.531, 
    5299.018,
  5167.016, 5161.914, 5160.405, 5163.83, 5169.875, 5173.607, 5183.064, 
    5197.787, 5209.045, 5212.517, 5219.128, 5226.534, 5234.539, 5240.672, 
    5249.209,
  5156.191, 5150.679, 5149.7, 5154.202, 5162.06, 5167.629, 5179.987, 
    5193.339, 5205.378, 5214.872, 5223.599, 5233.404, 5242.848, 5252.047, 
    5262.035,
  5146.132, 5140.618, 5141.152, 5146.53, 5158.076, 5166.164, 5174.533, 
    5194.889, 5208.222, 5217.061, 5228.009, 5239.207, 5251.073, 5261.287, 
    5272.44,
  5136.317, 5131.203, 5131.891, 5138.403, 5152.992, 5160.058, 5174.341, 
    5184.523, 5203.375, 5217.664, 5231.396, 5243.433, 5257.495, 5269.512, 
    5283.454,
  5126.777, 5122.985, 5123.496, 5133.373, 5147.937, 5162.785, 5166.44, 
    5185.328, 5203.505, 5217.7, 5233.02, 5246.786, 5261.36, 5274.41, 5288.933,
  5116.944, 5113.329, 5114.212, 5123.693, 5141.38, 5155.195, 5166.963, 
    5174.706, 5193.658, 5216.923, 5232.721, 5248.967, 5262.709, 5277.712, 
    5291.783,
  5105.68, 5103.664, 5106.798, 5116.973, 5136.133, 5153.822, 5162.127, 
    5175.845, 5193.98, 5212.195, 5231.905, 5247.91, 5262.782, 5276.328, 
    5290.26,
  5093.209, 5091.921, 5097.228, 5108.931, 5127.932, 5147.847, 5160.92, 
    5168.394, 5182.814, 5206.421, 5226.388, 5243.693, 5259.565, 5273.043, 
    5286.386,
  5080.514, 5080.129, 5090.712, 5104.916, 5126.029, 5145.149, 5158.11, 
    5169.256, 5181.671, 5199.471, 5219.408, 5238.38, 5253.468, 5266.625, 
    5278.697,
  5071.25, 5069.561, 5081.988, 5098.258, 5120.943, 5142.161, 5157.231, 
    5165.92, 5176.339, 5194.555, 5215.471, 5232.681, 5247.519, 5259.852, 
    5270.255,
  5120.631, 5111.266, 5102.017, 5094.027, 5086.611, 5081.461, 5079.477, 
    5082.503, 5090.765, 5097.025, 5102.496, 5106.153, 5108.553, 5111.517, 
    5118.575,
  5114.728, 5103.945, 5095.146, 5087.284, 5080.731, 5076.784, 5075.572, 
    5077.145, 5085.056, 5094.032, 5099.682, 5103.618, 5105.949, 5108.998, 
    5116.424,
  5107.222, 5095.72, 5088.024, 5081.292, 5076.341, 5073.878, 5071.477, 
    5076.88, 5085.618, 5091.938, 5098.212, 5102.254, 5104.611, 5108.761, 
    5116.308,
  5096.622, 5086.12, 5079.254, 5074.095, 5071.953, 5069.818, 5071.128, 
    5071.368, 5081.736, 5089.793, 5097.773, 5101.417, 5105.374, 5110.352, 
    5120.288,
  5083.747, 5074.168, 5069.658, 5067.655, 5067.794, 5070.122, 5069.066, 
    5073.753, 5082.917, 5090.096, 5098.177, 5103.007, 5108.51, 5114.704, 
    5126.04,
  5068.66, 5060.645, 5057.737, 5058.301, 5060.118, 5064.673, 5067.797, 
    5070.899, 5079.699, 5091.904, 5100.144, 5106.575, 5113.21, 5122.689, 
    5134.433,
  5053.681, 5047.378, 5047.056, 5050.304, 5053.95, 5060.879, 5063.573, 
    5072.299, 5083.586, 5093.933, 5103.77, 5111.584, 5120.532, 5131.469, 
    5144.001,
  5041.194, 5035.311, 5035.488, 5041.99, 5046.655, 5055.939, 5061.714, 
    5068.885, 5081.357, 5095.521, 5106.795, 5117.399, 5128.736, 5141.142, 
    5155.088,
  5031.869, 5025.542, 5027.749, 5037.106, 5043.467, 5053.294, 5060.348, 
    5071.195, 5084.748, 5097.437, 5110.759, 5123.693, 5136.625, 5150.298, 
    5164.578,
  5026.285, 5017.734, 5023.104, 5032.618, 5039.347, 5051.131, 5060.253, 
    5069.147, 5083.426, 5099.283, 5114.627, 5128.856, 5143.628, 5158.505, 
    5173.359,
  5088.929, 5084.696, 5079.434, 5072.782, 5068.599, 5063.489, 5057.007, 
    5051.805, 5048.183, 5045.645, 5050.028, 5056.357, 5061.39, 5066.655, 
    5075.825,
  5071.022, 5066.466, 5063.085, 5056.914, 5054.698, 5049.742, 5048.78, 
    5042.288, 5039.011, 5040.17, 5044.633, 5052.438, 5058.555, 5064.313, 
    5072.37,
  5054.66, 5049.335, 5045.866, 5042.383, 5040.996, 5042.072, 5034.31, 
    5036.557, 5031.837, 5033.01, 5038.819, 5047.26, 5054.133, 5060.855, 
    5067.91,
  5037.585, 5031.555, 5028.173, 5026.96, 5027.565, 5027.722, 5031.257, 
    5022.536, 5025.347, 5026.27, 5032.969, 5040.438, 5048.801, 5055.418, 
    5063.881,
  5018.294, 5011.857, 5010.724, 5013.219, 5017.323, 5022.11, 5020.229, 
    5022.348, 5018.123, 5021.413, 5027.474, 5034.693, 5042.753, 5048.938, 
    5058.175,
  4996.848, 4989.711, 4992.167, 4999.695, 5006.082, 5011.399, 5015.91, 
    5014.562, 5015.573, 5019.312, 5022.89, 5029.972, 5036.118, 5043.089, 
    5051.72,
  4973.886, 4967.954, 4972.411, 4986.688, 4997.121, 5004.528, 5007.082, 
    5010.73, 5012.638, 5014.98, 5020.374, 5024.813, 5030.553, 5036.848, 
    5045.53,
  4959.478, 4957.303, 4964.509, 4979.318, 4989.455, 4997.699, 5001.839, 
    5004.041, 5007.186, 5012.198, 5015.885, 5019.977, 5025.624, 5031.96, 
    5041.436,
  4956.414, 4958.098, 4966.094, 4980.459, 4987.599, 4994.316, 4997.796, 
    5001.667, 5005.864, 5010.266, 5013.403, 5017.482, 5022.647, 5029.486, 
    5039.58,
  4960.883, 4963.455, 4972.548, 4982.541, 4987.175, 4993.793, 4996.528, 
    5000.243, 5006.171, 5011.543, 5013.239, 5017.073, 5023.116, 5030.83, 
    5041.985,
  5076.95, 5075.854, 5075.317, 5074.65, 5074.686, 5073.528, 5072.964, 
    5073.444, 5073.117, 5068.408, 5063.33, 5057.373, 5052.721, 5046.865, 
    5044.544,
  5061.723, 5058.688, 5057.326, 5055.68, 5055.002, 5054.448, 5056.201, 
    5054.765, 5055.2, 5056.177, 5052.046, 5048.536, 5044.815, 5042.31, 
    5040.804,
  5042.623, 5039.188, 5036.783, 5036.802, 5036.431, 5038.977, 5035.554, 
    5043.005, 5042.261, 5041.912, 5040.402, 5038.898, 5037.579, 5036.419, 
    5037.445,
  5021.683, 5018.449, 5017.747, 5018.354, 5020.036, 5021.806, 5027.029, 
    5021.835, 5029.529, 5030.361, 5030.577, 5028.762, 5031.114, 5031.426, 
    5035.808,
  4994.168, 4991.959, 4993.614, 4998.267, 5003.174, 5008.281, 5011.067, 
    5017.286, 5015.236, 5016.542, 5019.634, 5019.246, 5024.348, 5026.596, 
    5033.696,
  4971.346, 4969.044, 4971.399, 4978.526, 4987.51, 4995.513, 5001.981, 
    5003.187, 5007.285, 5010.493, 5010.802, 5013.129, 5018.329, 5024.125, 
    5031.51,
  4956.561, 4952.651, 4958.044, 4963.328, 4976.984, 4989.753, 4994.515, 
    4999.254, 4999.904, 5001.419, 5004.625, 5007.766, 5013.816, 5021.719, 
    5030.123,
  4954.983, 4950.01, 4955.121, 4959.153, 4973.29, 4987.836, 4992.892, 
    4992.528, 4992.476, 4996.172, 4998.17, 5002.935, 5010.438, 5019.963, 
    5029.61,
  4969.387, 4963.819, 4963.69, 4966.997, 4978.727, 4988.772, 4989.843, 
    4990.537, 4988.652, 4989.771, 4992.939, 4999.366, 5007.158, 5018.076, 
    5028.57,
  4978.798, 4974.665, 4974.474, 4977.106, 4982.198, 4986.666, 4986.056, 
    4983.813, 4982.514, 4985.991, 4989.743, 4995.733, 5004.363, 5015.863, 
    5027.585,
  5100.354, 5099.584, 5100.279, 5101.729, 5106.011, 5109.836, 5114.629, 
    5120.433, 5124.212, 5124.861, 5125.893, 5126.113, 5124.057, 5120.688, 
    5115.611,
  5079.938, 5079.788, 5082.914, 5086.222, 5089.196, 5093.654, 5099.239, 
    5100.411, 5103.824, 5108.664, 5108.201, 5109.14, 5107.129, 5105.252, 
    5099.139,
  5054.524, 5053.325, 5055.926, 5062.882, 5069.504, 5078.682, 5077.514, 
    5088.479, 5085.807, 5088.417, 5090.087, 5091.663, 5090.823, 5088.792, 
    5085.437,
  5034.188, 5028.625, 5030.017, 5034.338, 5044.358, 5050.962, 5065.508, 
    5060.344, 5071.298, 5072.877, 5075.022, 5075.347, 5076.336, 5075.094, 
    5072.191,
  5020.375, 5009.763, 5008.364, 5012.939, 5019.805, 5030.023, 5033.629, 
    5046.994, 5046.989, 5050.357, 5056.109, 5057.525, 5060.148, 5059.83, 
    5060.764,
  5013.727, 4999.768, 4994.874, 4997.584, 5002.323, 5008.082, 5016.706, 
    5019.394, 5028.232, 5035.652, 5038.344, 5042.092, 5045.794, 5048.192, 
    5050.202,
  5013.844, 4998.553, 4994.144, 4996.473, 4996.85, 4997.438, 5000.942, 
    5007.707, 5012.616, 5016.086, 5022.711, 5027.291, 5033.003, 5036.893, 
    5041.006,
  5019.212, 5002.743, 4991.275, 4986.277, 4985.427, 4990.072, 4993.552, 
    4996.073, 4999.423, 5005.483, 5010.664, 5016.958, 5023.245, 5028.406, 
    5033.722,
  5025.912, 5009.738, 4998.929, 4993.755, 4993.998, 4996.341, 4996.883, 
    4998.176, 4996.717, 4998.745, 5003.242, 5009.572, 5014.857, 5021.824, 
    5028.451,
  5034.897, 5018.513, 5005.983, 5001.292, 4999.439, 5000.465, 4998.735, 
    4995.57, 4992.862, 4994.843, 4998.02, 5003.552, 5009.305, 5017.834, 
    5025.604,
  5125.722, 5117.797, 5111.668, 5108.459, 5108.258, 5110.023, 5113.647, 
    5121.172, 5128.792, 5135.788, 5144.067, 5152.825, 5159.833, 5166.532, 
    5171.156,
  5115.079, 5103.31, 5091.895, 5085.634, 5083.325, 5086.282, 5092.509, 
    5097.057, 5104.675, 5115.406, 5122.464, 5131.939, 5139.174, 5148.129, 
    5152.182,
  5108.447, 5092.419, 5077.167, 5068.074, 5062.945, 5068.891, 5068.133, 
    5082.475, 5087.203, 5096.47, 5105.375, 5115.015, 5123.184, 5130.967, 
    5138.404,
  5101.512, 5082.447, 5066.301, 5054.508, 5050.048, 5047.042, 5059.477, 
    5058.403, 5073.999, 5083.973, 5094.208, 5102.317, 5111.807, 5120.041, 
    5126.852,
  5097.292, 5077.272, 5059.019, 5049.283, 5042.269, 5042.016, 5040.53, 
    5052.271, 5060.676, 5071.162, 5084.431, 5092.95, 5102.426, 5109.622, 
    5117.902,
  5094.398, 5074.299, 5056.145, 5044.597, 5036.792, 5034.112, 5035.575, 
    5036.29, 5045.668, 5061.583, 5072.423, 5084.619, 5093.771, 5102.865, 
    5110.141,
  5093.811, 5075.589, 5056.569, 5043.159, 5033.666, 5029.244, 5027.303, 
    5031.781, 5037.367, 5047.022, 5061.012, 5073.312, 5083.617, 5093.835, 
    5101.823,
  5094.181, 5076.896, 5057.554, 5041.75, 5028.997, 5022.525, 5020.317, 
    5019.783, 5023.972, 5034.795, 5047.14, 5059.668, 5072.918, 5084.799, 
    5093.683,
  5096.555, 5081.59, 5063.417, 5045.786, 5032.06, 5022.55, 5018.029, 
    5017.177, 5016.853, 5022.09, 5033.908, 5048.107, 5062.098, 5075.523, 
    5085.718,
  5098.792, 5084.155, 5066.617, 5048.86, 5031.66, 5020.556, 5017.009, 
    5014.624, 5013.461, 5016.57, 5025.661, 5038.73, 5053.618, 5068.055, 
    5079.489,
  5184.299, 5168.317, 5151.971, 5136.222, 5123.608, 5114.601, 5108.626, 
    5108.255, 5110.004, 5114.175, 5122.533, 5132.308, 5142.793, 5153.675, 
    5165.382,
  5181.928, 5163.775, 5145.43, 5127.885, 5113.475, 5101.583, 5096.912, 
    5090.444, 5090.77, 5095.424, 5101.337, 5112.323, 5122.027, 5134.328, 
    5142.701,
  5179.973, 5161.916, 5142.594, 5124.912, 5107.504, 5098.082, 5083.954, 
    5083.068, 5076.444, 5076.629, 5080.67, 5089.768, 5101.04, 5112.342, 
    5123.221,
  5178.342, 5160.767, 5142.888, 5124.007, 5106.617, 5091.058, 5084.074, 
    5070.202, 5067.719, 5065.351, 5066.12, 5072.048, 5081.545, 5094.025, 
    5104.955,
  5176.562, 5161.771, 5145.758, 5127.116, 5109.04, 5092.65, 5077.563, 
    5070.269, 5060.991, 5056.201, 5057.158, 5060.228, 5068.206, 5077.034, 
    5089.693,
  5175.259, 5163.27, 5148.498, 5130.927, 5110.94, 5093.117, 5077.667, 
    5063.186, 5054.19, 5050.602, 5050.909, 5055.131, 5061.625, 5069.585, 
    5080.477,
  5174.513, 5166.882, 5153.071, 5135.44, 5115.248, 5094.461, 5076.285, 
    5062.667, 5051.224, 5044.606, 5046.959, 5052.709, 5059.591, 5067.116, 
    5077.6,
  5176.395, 5168.82, 5154.59, 5137.531, 5115.329, 5094.142, 5074.979, 
    5058.087, 5045.588, 5040.01, 5043.06, 5051.731, 5059.934, 5068.552, 
    5079.693,
  5178.653, 5170.867, 5156.572, 5136.746, 5113.899, 5092.012, 5071.792, 5056, 
    5043.097, 5035.613, 5039.577, 5050.754, 5060.8, 5071.876, 5083.353,
  5181.353, 5168.173, 5150.66, 5129.621, 5105.924, 5085.091, 5066.343, 
    5048.903, 5037.091, 5031.061, 5035.994, 5049.161, 5062.251, 5075.827, 
    5086.946,
  5259.777, 5250.472, 5245.604, 5236.17, 5224.272, 5208.981, 5189.2, 
    5174.134, 5157.215, 5135.962, 5120.919, 5108.889, 5100.728, 5095.964, 
    5095.747,
  5258.22, 5252.359, 5247.334, 5237.155, 5223.109, 5203.147, 5190.41, 
    5161.955, 5141.872, 5127.601, 5110.115, 5097.576, 5088.78, 5086.248, 
    5085.244,
  5259.867, 5256.716, 5250.007, 5239.727, 5219.418, 5205.418, 5171.182, 
    5165.728, 5135.802, 5114.921, 5098.204, 5086.205, 5076.996, 5074.816, 
    5077.324,
  5263.501, 5259.422, 5251.534, 5236.451, 5216.924, 5190.941, 5172.312, 
    5132.8, 5119.832, 5101.838, 5086.108, 5073.602, 5066.183, 5063.843, 
    5068.669,
  5268.409, 5262.888, 5253.053, 5234.454, 5211.51, 5183.039, 5151.568, 
    5132.901, 5108.729, 5085.6, 5073.791, 5061.218, 5055.721, 5051.863, 
    5059.299,
  5273.339, 5265.887, 5251.297, 5229.256, 5199.239, 5167.065, 5135.039, 
    5106.021, 5086.3, 5073.733, 5060.5, 5051.551, 5046.202, 5043.572, 5048.718,
  5279.43, 5270.221, 5251.207, 5224.757, 5191.445, 5152.514, 5117.732, 
    5094.702, 5076.438, 5061.122, 5051.364, 5044.01, 5039.992, 5038.554, 
    5041.459,
  5286.12, 5271.718, 5248.826, 5219.323, 5179.461, 5139.834, 5102.747, 
    5076.208, 5060.58, 5052.51, 5044.037, 5038.167, 5036.541, 5036.291, 
    5038.639,
  5290.996, 5274.985, 5251.77, 5217.932, 5176.906, 5133.229, 5094.314, 
    5069.537, 5054.909, 5046, 5038.517, 5034.436, 5034.136, 5034.352, 5037.571,
  5295.632, 5275.861, 5249.011, 5213.736, 5170.94, 5127.734, 5089.229, 
    5059.978, 5045.739, 5041.083, 5034.44, 5032.105, 5033.217, 5035.202, 
    5039.409,
  5338.474, 5333.484, 5326.592, 5307.413, 5280.249, 5245.187, 5203.405, 
    5173.65, 5151.187, 5129.483, 5116.438, 5108.652, 5103.664, 5101.027, 
    5100.669,
  5340.541, 5339.309, 5327.779, 5304.542, 5273.26, 5227.386, 5192.047, 
    5146.794, 5120.932, 5107.901, 5097.75, 5092.893, 5089.188, 5089.177, 
    5087.601,
  5348.604, 5345.146, 5330.134, 5307.675, 5268.887, 5230.776, 5168.706, 
    5143.478, 5114.583, 5097.396, 5087.084, 5084.665, 5080.932, 5080.37, 
    5078.485,
  5356.327, 5350.316, 5335.491, 5308.692, 5273.867, 5222.467, 5179.667, 
    5130.218, 5104.767, 5092.942, 5083.38, 5077.042, 5073.149, 5070.731, 
    5069.425,
  5364.415, 5356.718, 5341.432, 5315.884, 5281.168, 5234.87, 5180.116, 
    5143.725, 5118.657, 5093.044, 5082.492, 5072.16, 5068.177, 5063.745, 
    5062.793,
  5371.086, 5363.438, 5346.66, 5323.238, 5288.533, 5245.495, 5198.775, 
    5151.789, 5120.765, 5101.515, 5085.087, 5073.69, 5066.68, 5061.421, 
    5058.762,
  5377.924, 5370.534, 5353.836, 5331.977, 5301.306, 5261.918, 5215.373, 
    5174.084, 5142.187, 5114.6, 5093.7, 5078.689, 5067.891, 5061.546, 5057.933,
  5384.884, 5376.434, 5360.667, 5339.562, 5309.894, 5275.012, 5235.744, 
    5191.017, 5154.884, 5128.057, 5104.864, 5085.795, 5072.444, 5064.729, 
    5061.66,
  5391.721, 5383.375, 5368.462, 5348.504, 5323.258, 5289.914, 5252.138, 
    5213.69, 5175.915, 5144.063, 5116.438, 5095.144, 5078.415, 5068.895, 
    5066.51,
  5396.308, 5387.213, 5374.254, 5355.427, 5329.307, 5299.145, 5265.853, 
    5227.463, 5189.579, 5157.286, 5129.304, 5105.208, 5086.042, 5073.516, 
    5071.403,
  5375.866, 5381.691, 5380.299, 5369.069, 5349.762, 5320.814, 5280.719, 
    5243.806, 5205.633, 5159.906, 5123.705, 5097.753, 5084.477, 5071.914, 
    5064.718,
  5383.135, 5388.782, 5386.651, 5377.186, 5360.035, 5330.22, 5302.663, 
    5256.349, 5215.071, 5178.188, 5139.08, 5108.422, 5090.63, 5081.557, 
    5073.642,
  5391.178, 5396.996, 5393.572, 5387.04, 5367.166, 5351.537, 5309.614, 
    5286.105, 5247.537, 5201.977, 5159.918, 5124.614, 5099.965, 5090.988, 
    5085.314,
  5399.917, 5403.598, 5402.37, 5393.313, 5381.644, 5354.971, 5336.443, 
    5297.405, 5259.074, 5223.985, 5182.899, 5144.888, 5114.438, 5098.059, 
    5093.998,
  5408.195, 5410.905, 5410.667, 5402.245, 5390.72, 5371.806, 5345.81, 
    5317.637, 5290.887, 5245.912, 5207.391, 5166.782, 5134.309, 5109.846, 
    5100.778,
  5415.235, 5419.21, 5417.497, 5411.308, 5397.886, 5379.287, 5359.232, 
    5330.109, 5297.093, 5266.78, 5230.646, 5190.406, 5155.017, 5126.176, 
    5110.791,
  5421.641, 5425.464, 5423.565, 5417.065, 5405.484, 5389.501, 5367.07, 
    5344.954, 5318.975, 5284.664, 5248.726, 5212.934, 5175.918, 5145.55, 
    5124.135,
  5426.075, 5429.092, 5427.489, 5421.471, 5408.69, 5393.215, 5374.68, 
    5350.491, 5322.615, 5295.624, 5264.256, 5229.903, 5195.407, 5162.696, 
    5139.615,
  5427.322, 5430.026, 5427.9, 5421.071, 5411.3, 5396.745, 5377.176, 5356.671, 
    5332.987, 5304.008, 5274.058, 5242.021, 5210.634, 5178.119, 5153.277,
  5424.265, 5425.65, 5424.45, 5418.813, 5406.823, 5391.959, 5374.296, 
    5351.877, 5327.973, 5304.337, 5278.03, 5248.951, 5219.309, 5189.664, 
    5163.714,
  5423.144, 5437.361, 5446.691, 5447.655, 5441.532, 5428.567, 5406.219, 
    5380.248, 5345.682, 5300.563, 5255.206, 5210.509, 5178.315, 5159.667, 
    5152.984,
  5423.698, 5439.086, 5448.154, 5449.993, 5445.507, 5432.71, 5418.354, 
    5388.472, 5355.995, 5322.413, 5282.808, 5242.71, 5205.289, 5185.17, 
    5174.906,
  5426.854, 5443.121, 5450.569, 5454.535, 5448.015, 5443.076, 5420.385, 
    5405.696, 5378.288, 5343.645, 5307.353, 5271.83, 5236.756, 5209.215, 
    5196.295,
  5432.209, 5446.289, 5454.32, 5455.835, 5452.82, 5441.915, 5431.729, 
    5408.938, 5382.231, 5359.114, 5327.165, 5295.507, 5264.209, 5235.198, 
    5216.841,
  5438.228, 5449.522, 5457.026, 5457.944, 5455.186, 5447.226, 5433.293, 
    5417.863, 5399.292, 5367.836, 5342.213, 5312.665, 5285.125, 5258.504, 
    5235.137,
  5442.683, 5451.844, 5456.931, 5457.934, 5453.4, 5445.005, 5433.633, 
    5414.613, 5393.361, 5372.792, 5348.981, 5323.05, 5298.187, 5273.837, 
    5252.517,
  5445.994, 5453.217, 5455.313, 5454.357, 5449.686, 5441.21, 5427.523, 
    5412.823, 5393.933, 5370.812, 5348.383, 5325.896, 5303.003, 5280.973, 
    5261.542,
  5447.698, 5451.003, 5450.417, 5447.982, 5440.213, 5430.162, 5416.767, 
    5399.395, 5380.355, 5361.993, 5341.677, 5320.599, 5300.024, 5280.385, 
    5263.358,
  5446.881, 5447.22, 5443.341, 5436.461, 5428, 5415.951, 5401.102, 5385.865, 
    5368.165, 5347.996, 5327.889, 5308.479, 5289.538, 5272.026, 5257.2,
  5442.322, 5437.282, 5430.582, 5422.033, 5409.269, 5394.877, 5380.18, 
    5362.539, 5344.964, 5327.931, 5309.364, 5290.54, 5273.059, 5257.657, 
    5245.05,
  5465.753, 5482.748, 5494.926, 5498.979, 5498.833, 5492.716, 5479.396, 
    5465.587, 5446.812, 5423.677, 5403.208, 5384.017, 5365.799, 5352.416, 
    5344.86,
  5473.21, 5489.752, 5500.086, 5504.989, 5504.279, 5497.042, 5488.245, 
    5469.708, 5452.171, 5435.875, 5415.348, 5396.19, 5376.832, 5360.41, 
    5347.087,
  5483.512, 5498.724, 5506.122, 5511.105, 5507.774, 5505.433, 5490.557, 
    5481.102, 5462.094, 5441.441, 5422.617, 5403.791, 5383.811, 5365.723, 
    5348.693,
  5493.903, 5505.37, 5513.012, 5514.817, 5513.795, 5502.818, 5496.143, 
    5477.219, 5461.046, 5444.836, 5423.561, 5405.504, 5385.307, 5367.117, 
    5348.126,
  5503.324, 5513.108, 5518.616, 5519.112, 5515.081, 5508.771, 5493.55, 
    5480.451, 5463.301, 5441.426, 5422.664, 5401.105, 5382.615, 5361.537, 
    5342.916,
  5510.885, 5518.87, 5521.29, 5521.111, 5514.528, 5504.074, 5491.918, 
    5473.853, 5454.558, 5435.648, 5415.283, 5393.228, 5373.023, 5351.742, 
    5331.787,
  5519.458, 5525.018, 5524.206, 5519.912, 5511.601, 5500.248, 5484.111, 
    5467.135, 5446.756, 5424.9, 5402.803, 5380.375, 5357.62, 5335.388, 
    5313.935,
  5526.258, 5526.866, 5523.117, 5516.534, 5504.188, 5489.787, 5472.782, 
    5453.354, 5431.429, 5409.535, 5385.813, 5361.686, 5337.435, 5313.794, 
    5291.088,
  5531.906, 5529.312, 5521.224, 5509.215, 5494.957, 5477.35, 5457.158, 
    5437.109, 5413.773, 5388.689, 5363.377, 5337.62, 5311.348, 5286.137, 
    5261.898,
  5531.69, 5522.692, 5511.431, 5498.745, 5480.064, 5459.172, 5437.06, 
    5411.828, 5387.042, 5361.963, 5335.368, 5307.507, 5279.5, 5253.507, 
    5228.207,
  5522.199, 5537.662, 5552.486, 5562.635, 5570.654, 5575.654, 5578.098, 
    5577.662, 5572.53, 5560.517, 5547.333, 5531.355, 5511.355, 5487.393, 
    5463.615,
  5514.332, 5533.665, 5552.437, 5566.089, 5575.141, 5579.453, 5580.354, 
    5576.144, 5570.471, 5562.486, 5546.156, 5526.125, 5503.285, 5477.667, 
    5449.536,
  5505.579, 5528.972, 5549.92, 5566.373, 5574.853, 5581.566, 5580.667, 
    5579.478, 5567.194, 5551.148, 5534.725, 5515.885, 5489.382, 5461.252, 
    5428.979,
  5497.282, 5522.042, 5546.068, 5562.919, 5575.382, 5575.866, 5576.859, 
    5567.555, 5561.686, 5548.628, 5522.563, 5499.749, 5471.675, 5439.912, 
    5402.37,
  5489.678, 5515.375, 5540.625, 5558.495, 5569.576, 5574.12, 5570.359, 
    5562.995, 5548.457, 5526.167, 5507.829, 5476.433, 5446.524, 5408.527, 
    5369.317,
  5484.307, 5509.756, 5533.785, 5552.797, 5562.677, 5563.494, 5557.622, 
    5544.128, 5528.934, 5508.729, 5481.069, 5447.091, 5411.016, 5368.424, 
    5325.768,
  5482.907, 5507.765, 5529.03, 5545.131, 5552.885, 5552.012, 5543.394, 
    5528.825, 5506.558, 5478.526, 5447.171, 5409.169, 5365.367, 5318.984, 
    5269.486,
  5485.332, 5506.317, 5524.27, 5537.3, 5540.107, 5535.521, 5522.25, 5503.393, 
    5478.952, 5448.089, 5408.895, 5362.846, 5314.011, 5261.356, 5208.376,
  5489.636, 5507.461, 5520.748, 5526.463, 5526.099, 5516.853, 5499.771, 
    5476.442, 5444.016, 5404.393, 5358.324, 5308.208, 5254.021, 5197.185, 
    5147.023,
  5493.355, 5505.06, 5512.525, 5515.638, 5507.521, 5492.2, 5469.26, 5436.997, 
    5399.04, 5353.358, 5302.866, 5246.935, 5187.887, 5135.156, 5089.808,
  5516.728, 5514.63, 5510.786, 5506.859, 5506.73, 5509.365, 5516.027, 
    5524.736, 5531.662, 5535.065, 5536.718, 5532.82, 5521.363, 5503.814, 
    5479.319,
  5501.769, 5502.256, 5501.561, 5500.29, 5500.875, 5503.044, 5508.832, 
    5512.346, 5518.674, 5523.497, 5519.812, 5513.448, 5500.408, 5482.305, 
    5454.708,
  5483.593, 5486.835, 5488.325, 5490.552, 5491.703, 5496.37, 5496.937, 
    5506.444, 5502.923, 5503.297, 5500.915, 5492.782, 5476.585, 5455.282, 
    5426.937,
  5462.044, 5467.64, 5471.482, 5474.141, 5478.435, 5479.511, 5486.888, 
    5482.126, 5489.636, 5485.6, 5477.608, 5468.266, 5450.809, 5427.594, 
    5395.218,
  5438.367, 5444.344, 5449.102, 5454.378, 5458.316, 5464.43, 5463.312, 
    5473.666, 5463.507, 5461.547, 5454.745, 5440.904, 5423.342, 5396.255, 
    5363.815,
  5413.074, 5418.073, 5422.199, 5427.502, 5431.699, 5437.168, 5441.677, 
    5438.483, 5441.091, 5435.591, 5423.875, 5409.889, 5390.029, 5362.601, 
    5330.555,
  5386.708, 5390.161, 5392.817, 5397.335, 5403.192, 5407.834, 5411.029, 
    5414.43, 5409.079, 5400.636, 5392.042, 5375.373, 5353.218, 5324.981, 
    5292.547,
  5360.461, 5361.455, 5361.995, 5365.579, 5369.326, 5375.732, 5378.87, 
    5377.812, 5375.227, 5369.46, 5356.398, 5339.209, 5316.607, 5288.298, 
    5255.189,
  5337.388, 5336.707, 5336.347, 5338.783, 5341.878, 5344.771, 5347.106, 
    5348.467, 5344.61, 5336.999, 5325.958, 5308.689, 5284.16, 5254.453, 
    5219.261,
  5318.851, 5316.443, 5317.246, 5319.876, 5322.253, 5326.595, 5330.427, 
    5330.652, 5327.734, 5319.509, 5303.74, 5280.884, 5252.492, 5219.538, 
    5181.205,
  5506.228, 5481.876, 5460.354, 5442.147, 5427.611, 5415.068, 5404.516, 
    5398.608, 5392.194, 5385.144, 5381.569, 5378.271, 5373.736, 5366.864, 
    5357.947,
  5475.431, 5451.258, 5432.811, 5416.272, 5403.247, 5392.603, 5388.96, 
    5380.286, 5378.044, 5376.358, 5370.875, 5366.601, 5359.642, 5351.515, 
    5338.71,
  5446.493, 5425.731, 5408.986, 5395.947, 5383.922, 5379.255, 5369.292, 
    5373.348, 5365.29, 5362.684, 5357.903, 5352.322, 5342.659, 5331.691, 
    5317.998,
  5422.314, 5404.605, 5389.826, 5377.773, 5368.886, 5360.562, 5360.909, 
    5351.41, 5353.64, 5349.092, 5342.967, 5335.487, 5324.626, 5312.018, 
    5294.959,
  5404.769, 5388.725, 5374.605, 5364.104, 5356.038, 5350.851, 5343.254, 
    5345.025, 5336.977, 5331.95, 5326.501, 5316.243, 5305.192, 5289.052, 
    5270.489,
  5390.192, 5374.978, 5360.948, 5350.852, 5341.298, 5335.592, 5331.326, 
    5324.313, 5321.311, 5316.853, 5307.896, 5297.466, 5284.909, 5265.835, 
    5241.847,
  5378.214, 5363.87, 5349.416, 5338.288, 5329.464, 5322.495, 5316.809, 
    5313.766, 5307.139, 5299.295, 5291.708, 5280.772, 5263.751, 5239.178, 
    5208.554,
  5367.392, 5352.76, 5337.939, 5326.818, 5316.208, 5310.316, 5304.879, 
    5298.847, 5293.4, 5288.009, 5278.556, 5262.833, 5239.534, 5208.394, 
    5171.18,
  5357.26, 5343.309, 5329.007, 5317.792, 5309.307, 5302.753, 5295.923, 
    5291.053, 5285.675, 5276.326, 5261.953, 5239.457, 5208.548, 5170.565, 
    5127.758,
  5347.652, 5332.768, 5318.987, 5309.836, 5300.195, 5293.378, 5289.223, 
    5283.241, 5275.062, 5260.494, 5238.719, 5208.314, 5170.683, 5127.874, 
    5080.961,
  5571.661, 5544.717, 5517.583, 5492.14, 5468.352, 5443.679, 5415.108, 
    5393.268, 5371.391, 5345.272, 5327.481, 5313.37, 5302.556, 5292.617, 
    5285.143,
  5556.394, 5530.631, 5506.82, 5483.531, 5461.44, 5433.423, 5415.058, 
    5379.79, 5357.544, 5341.391, 5322.853, 5307.661, 5294.952, 5284.118, 
    5272.812,
  5542.342, 5520.661, 5499.309, 5479.766, 5454.965, 5436.905, 5400.946, 
    5390.13, 5359.434, 5335.439, 5316.225, 5300.654, 5284.562, 5271.41, 
    5258.003,
  5529.6, 5510.826, 5492.448, 5472.65, 5451.222, 5424.236, 5405.238, 5368.73, 
    5349.182, 5330.88, 5308.166, 5290.722, 5273.369, 5257.558, 5240.117,
  5519.269, 5503.621, 5488.11, 5469.027, 5448.113, 5423.497, 5395.107, 
    5374.371, 5348.268, 5318.819, 5300.394, 5277.757, 5260.479, 5239.125, 
    5220.886,
  5509.387, 5495.906, 5481.119, 5463.831, 5441.063, 5416.723, 5391.229, 
    5360.486, 5334.23, 5311.634, 5287.942, 5264.395, 5243.89, 5219.357, 
    5195.599,
  5500.562, 5490.216, 5476.462, 5458.498, 5436.512, 5411.178, 5382.959, 
    5356.761, 5328.56, 5299.756, 5274.374, 5249.148, 5223.283, 5195.491, 
    5165.466,
  5492.714, 5482.332, 5467.51, 5449.779, 5425.139, 5399.823, 5371.376, 
    5340.734, 5311.898, 5285.948, 5258.161, 5229.617, 5200.086, 5166.912, 
    5130.91,
  5485.719, 5476.076, 5460.363, 5439.781, 5415.314, 5387.168, 5355.697, 
    5327.328, 5298.347, 5267.871, 5237.908, 5206.413, 5171.407, 5133.151, 
    5091.284,
  5477.358, 5463.275, 5445.063, 5424.228, 5396.244, 5366.437, 5335.67, 
    5304.551, 5274.726, 5246.251, 5213.946, 5178.003, 5139.126, 5095.32, 
    5052.383,
  5590.833, 5583.125, 5574.046, 5567.603, 5563.003, 5553.458, 5541.217, 
    5528.753, 5509.945, 5480.666, 5453.624, 5424.586, 5395.03, 5361.152, 
    5329.357,
  5580.264, 5573.269, 5565.105, 5559.544, 5553.311, 5544.248, 5535.724, 
    5512.144, 5493.062, 5473.849, 5446.658, 5416.686, 5384.272, 5350.776, 
    5313.164,
  5567.623, 5561.004, 5553.596, 5548.956, 5540.798, 5534.45, 5517.54, 
    5517.747, 5489.265, 5460.119, 5433.589, 5406.187, 5371.027, 5334.004, 
    5293.229,
  5551.177, 5544.938, 5538.757, 5533.375, 5526.433, 5516.491, 5508.332, 
    5483.337, 5472.125, 5452.59, 5420.61, 5390.686, 5355.361, 5315.535, 
    5270.487,
  5532.454, 5526.457, 5520.987, 5515.914, 5509.36, 5500.564, 5487.715, 
    5477.506, 5455.293, 5427.001, 5403.96, 5369.942, 5334.878, 5291.297, 
    5245.173,
  5510.779, 5505.904, 5500.141, 5496.571, 5489.853, 5482.145, 5469.83, 
    5449.898, 5431.646, 5410.436, 5381.755, 5347.851, 5309.854, 5264.993, 
    5216.166,
  5489.335, 5485.786, 5480.441, 5476.459, 5470.899, 5462.21, 5449.309, 
    5433.882, 5411.349, 5385.363, 5357.781, 5323.322, 5281.897, 5234.995, 
    5183.79,
  5468.341, 5464.374, 5459.426, 5456.389, 5449.935, 5441.552, 5427.25, 
    5408.247, 5387.51, 5364.652, 5333.775, 5296.231, 5253.478, 5205.23, 
    5151.854,
  5447.01, 5444.536, 5439.959, 5434.853, 5427.977, 5417.865, 5402.96, 
    5386.878, 5365.229, 5338.321, 5305.886, 5267.65, 5223.297, 5172.355, 
    5120.011,
  5423.532, 5418.789, 5414.273, 5410.575, 5403.257, 5392.247, 5377.078, 
    5358.001, 5336.499, 5310.925, 5277.375, 5237.419, 5191.823, 5141.02, 
    5090.627,
  5517.455, 5512.293, 5507.888, 5499.82, 5493.542, 5484.724, 5474.166, 
    5465.418, 5453.586, 5435.125, 5418.304, 5400.216, 5379.392, 5355.873, 
    5331.572,
  5490.237, 5484.247, 5480.406, 5472.72, 5465.461, 5457.898, 5453.34, 
    5434.425, 5422.632, 5413.38, 5395.191, 5377.716, 5357.318, 5337.345, 
    5311.766,
  5460.555, 5454.334, 5449.334, 5442.982, 5435.785, 5431.896, 5416.41, 
    5421.586, 5397.627, 5384.499, 5370.058, 5355.805, 5335.327, 5314.975, 
    5291.454,
  5427.981, 5423.041, 5417.741, 5411.942, 5406.055, 5398.043, 5397.687, 
    5376.663, 5377.098, 5363.735, 5347.475, 5333.115, 5315.482, 5296.023, 
    5271.762,
  5393.287, 5389.322, 5383.944, 5380.018, 5375.552, 5370.381, 5361.571, 
    5364.594, 5348.244, 5337.09, 5326.803, 5310.854, 5295.526, 5274.919, 
    5252.673,
  5358.154, 5355.711, 5350.534, 5349.464, 5344.899, 5342.616, 5338.054, 
    5328.216, 5324.474, 5317.309, 5303.496, 5290.498, 5275.187, 5255.448, 
    5232.088,
  5323.497, 5323.06, 5319.668, 5318.929, 5316.608, 5314.169, 5310.254, 
    5308.905, 5300.608, 5290.718, 5281.871, 5268.704, 5252.843, 5233.222, 
    5210.179,
  5293.46, 5292.925, 5290.154, 5291.16, 5289.049, 5288.721, 5284.669, 
    5278.965, 5274.074, 5268.748, 5258.109, 5245.323, 5230.585, 5211.39, 
    5188.33,
  5265.366, 5265.181, 5263.412, 5262.471, 5260.606, 5259.009, 5255.963, 
    5253.802, 5248.316, 5240.645, 5232.544, 5221.369, 5206.294, 5187.736, 
    5165.579,
  5237.98, 5235.561, 5233.453, 5233.529, 5232.262, 5229.929, 5226.298, 
    5221.001, 5217.037, 5212.893, 5205.708, 5195.29, 5181.966, 5164.838, 
    5143.142,
  5408.126, 5408.875, 5410.273, 5408.608, 5406.838, 5400.918, 5392.885, 
    5386.962, 5374.955, 5356.693, 5340.987, 5324.803, 5306.666, 5288.769, 
    5273.188,
  5370.484, 5372.963, 5375.022, 5372.682, 5367.946, 5363.025, 5361.42, 
    5344.729, 5332.937, 5326.778, 5309.178, 5294.542, 5277.442, 5263.974, 
    5247.425,
  5330.997, 5333.812, 5335.135, 5333.648, 5328.909, 5326.226, 5311, 5323.906, 
    5296.122, 5286.759, 5275.225, 5264.283, 5248.763, 5236.066, 5224.129,
  5282.564, 5286.091, 5287.609, 5286.187, 5282.765, 5276.971, 5281.146, 
    5259.137, 5266.034, 5253.287, 5241.798, 5232.979, 5223.521, 5212.758, 
    5202.156,
  5236.986, 5238.161, 5238.276, 5239.025, 5239.3, 5237.31, 5230.081, 
    5238.702, 5222.747, 5219.332, 5214.219, 5205.715, 5199.586, 5189.664, 
    5182.522,
  5192.671, 5193.929, 5193.497, 5196.416, 5196.08, 5197.837, 5196.736, 
    5188.783, 5191.24, 5191.689, 5184.019, 5181.464, 5176.301, 5170.18, 
    5163.747,
  5152.96, 5154.154, 5153.398, 5155.458, 5157.707, 5159.175, 5160.202, 
    5165.233, 5162.378, 5159.566, 5160.612, 5158.53, 5154.268, 5150.296, 
    5145.138,
  5113.528, 5113.463, 5112.968, 5117.572, 5120.297, 5125.844, 5128.629, 
    5129.738, 5133.095, 5137.643, 5137.176, 5136.542, 5135.463, 5132.673, 
    5128.39,
  5075.795, 5075.178, 5075.048, 5078.628, 5083.506, 5090.59, 5097.45, 
    5105.767, 5109.574, 5111.565, 5114.872, 5117.034, 5116.038, 5114.486, 
    5110.648,
  5044.486, 5039.186, 5036.812, 5040.14, 5045.235, 5053.418, 5062.209, 
    5070.539, 5079.453, 5088.085, 5093.308, 5096.604, 5097.422, 5096.285, 
    5091.741,
  5224.399, 5238.136, 5251.224, 5261.798, 5272.659, 5281.124, 5291.166, 
    5304.122, 5311.897, 5315.335, 5319.88, 5321.423, 5317.078, 5309.807, 
    5299.475,
  5195.491, 5209.279, 5224.256, 5236.329, 5245.211, 5256.112, 5267.915, 
    5273.175, 5280.495, 5291.19, 5290.184, 5290.27, 5285.165, 5279.554, 
    5265.775,
  5165.917, 5179.578, 5193.711, 5205.36, 5215.849, 5228.144, 5229.991, 
    5253.185, 5248.242, 5253.254, 5256.479, 5256.322, 5250.775, 5243.199, 
    5233.243,
  5133.329, 5144.476, 5157.349, 5167.43, 5179.565, 5183.91, 5206.138, 
    5197.581, 5219.556, 5220.914, 5218.33, 5217.166, 5215.977, 5208.027, 
    5197.831,
  5100.796, 5106.548, 5115.079, 5126.008, 5137.381, 5149.094, 5151.604, 
    5174.444, 5169.658, 5176.833, 5179.561, 5177.804, 5178.826, 5170.477, 
    5165.485,
  5074.271, 5075.224, 5078.057, 5083.935, 5089.462, 5097.659, 5107.61, 
    5108.199, 5126.564, 5135.164, 5133.407, 5138.501, 5138.689, 5135.513, 
    5131.774,
  5046.169, 5041.042, 5039.358, 5042.039, 5048.772, 5055.349, 5063.235, 
    5077.637, 5084.048, 5088.05, 5096.759, 5100.545, 5101.893, 5102.42, 
    5100.969,
  5030.703, 5017.257, 5007.18, 5003.684, 5002.348, 5008.357, 5015.567, 
    5022.493, 5035.208, 5049.216, 5056.217, 5062.895, 5068.624, 5071.272, 
    5071.726,
  5029.379, 5010.183, 4993.032, 4981.579, 4975.263, 4973.563, 4976.848, 
    4987.562, 4997.231, 5006.659, 5018.511, 5029.355, 5036.333, 5041.784, 
    5045.333,
  5043.798, 5018.139, 4996.816, 4980.689, 4966.506, 4960.277, 4959.285, 
    4962.875, 4973.139, 4986.667, 4997.746, 5006.9, 5014.442, 5020.351, 
    5023.787,
  5119.12, 5126.327, 5134.681, 5143.821, 5153.664, 5161.391, 5169.375, 
    5178.623, 5185.541, 5191.001, 5198.596, 5206.385, 5211.924, 5217.967, 
    5223.692,
  5098.463, 5103.446, 5109.565, 5117.56, 5124.863, 5134.707, 5144.686, 
    5149.104, 5156.092, 5166.463, 5170, 5177.023, 5181.898, 5189.018, 5191.477,
  5076.995, 5079.866, 5083.424, 5091.358, 5096.728, 5110.297, 5110.951, 
    5128.878, 5128.404, 5135.929, 5142.054, 5149.215, 5153.757, 5159.022, 
    5165.183,
  5061.95, 5059.639, 5060.785, 5063.229, 5070.327, 5072.378, 5090.42, 
    5085.813, 5103.171, 5108.155, 5113.741, 5119.12, 5125.925, 5131.089, 
    5135.903,
  5055.49, 5047.494, 5043.609, 5042.66, 5045.342, 5051.238, 5051.301, 
    5067.65, 5068.474, 5073.754, 5084.831, 5088.563, 5097.112, 5101.213, 
    5109.058,
  5059.386, 5045.682, 5035.269, 5030.439, 5026.743, 5026.868, 5032.051, 
    5029.033, 5037.91, 5044.683, 5046.934, 5053.568, 5059.604, 5064.936, 
    5071.678,
  5069.571, 5052.456, 5037.264, 5025.959, 5019.002, 5013.855, 5010.863, 
    5012.998, 5011.502, 5009.609, 5014.739, 5017.525, 5020.837, 5025.533, 
    5030.926,
  5084.678, 5065.847, 5047.205, 5032.25, 5017.768, 5008.112, 4999.755, 
    4991.602, 4987.38, 4985.345, 4981.489, 4979.731, 4980.571, 4982.047, 
    4985.548,
  5096.709, 5078.778, 5059.582, 5042.191, 5026.225, 5011.544, 4998.356, 
    4988.594, 4977.62, 4967.314, 4960.647, 4954.088, 4948.486, 4945.655, 
    4945.131,
  5108.284, 5088.592, 5068.551, 5050.395, 5030.653, 5013.758, 4997.893, 
    4982.684, 4971.068, 4960.952, 4951.256, 4942.322, 4935.669, 4930.895, 
    4927.916,
  5065.998, 5066.786, 5068.811, 5073.296, 5078.947, 5086.042, 5095.158, 
    5106.7, 5117.778, 5129.006, 5142.254, 5156.019, 5166.945, 5178.183, 
    5188.891,
  5061.762, 5058.326, 5056.12, 5056.619, 5057.647, 5062.751, 5069.673, 
    5075.002, 5084.533, 5097.09, 5105.771, 5118.095, 5128.285, 5141.72, 
    5149.204,
  5060.593, 5052.851, 5046.859, 5044.335, 5041.678, 5046.714, 5044.34, 
    5056.254, 5056.164, 5064.667, 5073.358, 5084.283, 5093.251, 5102.459, 
    5113.931,
  5059.878, 5049.403, 5041.178, 5033.486, 5029.562, 5024.063, 5031.119, 
    5025.041, 5035.443, 5039.096, 5044.823, 5052.24, 5061.401, 5070.213, 
    5077.91,
  5055.407, 5043.559, 5034.201, 5025.438, 5019.504, 5014.031, 5007.596, 
    5011.331, 5006.51, 5009.33, 5016.982, 5020.568, 5029.544, 5035.004, 
    5045.235,
  5047.962, 5033.875, 5022.502, 5013.96, 5005.423, 4999.714, 4996.212, 
    4989.081, 4989.437, 4989.292, 4987.806, 4991.069, 4996.771, 5002.384, 
    5010.31,
  5040.831, 5024.857, 5010.37, 4998.977, 4990.438, 4983.068, 4977.43, 
    4975.716, 4971.414, 4968.249, 4969.976, 4970.454, 4971.639, 4974.563, 
    4979.825,
  5037.598, 5017.046, 4998.132, 4984.273, 4971.016, 4962.545, 4955.604, 
    4950.363, 4948.333, 4949.086, 4948.359, 4950.041, 4952.81, 4955.621, 
    4958.796,
  5038.517, 5015.174, 4991.908, 4972.841, 4957.182, 4944.716, 4934.341, 
    4928.611, 4923.218, 4921.199, 4923.516, 4927.194, 4931.24, 4935.966, 
    4940.206,
  5044.979, 5015.372, 4988.504, 4966.032, 4944.923, 4929.413, 4917.037, 
    4906.894, 4901.08, 4898.219, 4897.354, 4899.66, 4905.066, 4912.647, 
    4919.666,
  5024.129, 5016.272, 5010.939, 5009.276, 5010.748, 5016.003, 5028.472, 
    5046.977, 5066.55, 5087.953, 5108.851, 5130.638, 5150.609, 5169.159, 
    5186.035,
  5018.775, 5010.791, 5004.744, 5001.459, 4999.067, 5002.021, 5007.302, 
    5015.518, 5031.119, 5052.199, 5069.813, 5090.177, 5106.735, 5127.98, 
    5140.41,
  5012.231, 5003.189, 4996.797, 4993.518, 4991.31, 4994.037, 4991.654, 
    5002.131, 5005.003, 5016.827, 5032.25, 5049.732, 5066.16, 5081.085, 
    5097.489,
  5004.913, 4993.789, 4986.847, 4981.917, 4980.738, 4977.927, 4986.418, 
    4979.167, 4990.802, 4996.235, 5005.651, 5016.962, 5031.301, 5045.975, 
    5058.376,
  4998.011, 4984.703, 4974.602, 4967.743, 4963.674, 4964.564, 4961.488, 
    4972.743, 4971.445, 4975.778, 4984.65, 4991.71, 5003.117, 5012.131, 
    5025.964,
  4994.341, 4978.031, 4964.154, 4953.603, 4945.077, 4940.485, 4942.009, 
    4938.984, 4947.835, 4958.073, 4962.931, 4972.479, 4981.31, 4989.879, 
    4999.971,
  4990.78, 4973.829, 4956.684, 4941.937, 4929.519, 4919.906, 4914.003, 
    4916.267, 4918.684, 4923.97, 4935.617, 4947.292, 4956.772, 4967.188, 
    4977.11,
  4987.298, 4969.198, 4948.807, 4931.083, 4913.069, 4899.688, 4890.208, 
    4884.482, 4885.561, 4894.296, 4904.436, 4916.087, 4928.951, 4941.362, 
    4953.759,
  4982.15, 4964.264, 4941.351, 4920.687, 4899.715, 4882.027, 4869.143, 
    4864.008, 4862.064, 4864.732, 4873.34, 4885.603, 4898.408, 4912.062, 
    4926.512,
  4977.893, 4957.876, 4932.165, 4909.862, 4886.161, 4866.236, 4851.729, 
    4842.457, 4841.646, 4846.226, 4853.199, 4861.521, 4871.943, 4884.434, 
    4899.026,
  4980.397, 4982.752, 4983.446, 4982.842, 4982.374, 4980.878, 4979.621, 
    4980.392, 4982.1, 4988.305, 5002.136, 5021.707, 5045.371, 5072.52, 
    5103.509,
  4966.796, 4969.836, 4970.506, 4969.137, 4966.979, 4966.118, 4966.107, 
    4962.639, 4963.207, 4969.713, 4977.696, 4994.643, 5013.891, 5042.021, 
    5068.792,
  4954.397, 4958.774, 4958.869, 4956.835, 4952.777, 4952.643, 4947.471, 
    4953.216, 4948.928, 4950.909, 4956.926, 4969.734, 4986.723, 5007.343, 
    5035.388,
  4946.007, 4948.678, 4946.421, 4941.619, 4937.186, 4931.836, 4936.101, 
    4928.362, 4936.05, 4937.264, 4941.418, 4948.803, 4963.186, 4983.049, 
    5006.151,
  4941.487, 4939.589, 4933.488, 4924.706, 4917.607, 4913.716, 4909.561, 
    4917.449, 4915.641, 4919.769, 4926.883, 4931.694, 4943.365, 4956.87, 
    4980.917,
  4941.238, 4932.983, 4923.359, 4909.889, 4898.526, 4892.338, 4890.718, 
    4887.748, 4894.195, 4902.922, 4908.404, 4916.671, 4926.021, 4938.312, 
    4956.897,
  4932.187, 4925.015, 4912.72, 4896.705, 4883.283, 4873.201, 4868.553, 
    4870.063, 4871.361, 4875.867, 4887.915, 4899.54, 4909.662, 4920.714, 
    4935.954,
  4930.773, 4917.581, 4901.332, 4883.653, 4865.196, 4853.559, 4844.992, 
    4841.11, 4844.03, 4852.917, 4863.785, 4878.634, 4893.975, 4907.396, 
    4920.868,
  4921.962, 4910.083, 4890.765, 4868.91, 4850.68, 4836.531, 4826.635, 
    4822.043, 4820.888, 4826.156, 4838.263, 4855.859, 4875.101, 4892.618, 
    4907.306,
  4911.017, 4896.647, 4874.71, 4854.864, 4834.837, 4818.61, 4806.333, 
    4799.104, 4799.588, 4806.217, 4817.456, 4833.976, 4856.431, 4878.381, 
    4896.333,
  4904.511, 4910.949, 4921.29, 4932.018, 4943.628, 4954.419, 4967.398, 
    4981.441, 4994.711, 5006.061, 5020.342, 5036.419, 5052.448, 5068.809, 
    5087.949,
  4883.843, 4892.065, 4903.016, 4915.092, 4926.615, 4939.526, 4953.254, 
    4964.682, 4977.867, 4993.109, 5004.854, 5019.066, 5032.609, 5050.233, 
    5064.156,
  4867.868, 4878.125, 4890.363, 4902.887, 4914.215, 4929.449, 4937.627, 
    4955.53, 4964.419, 4975.845, 4988.524, 5002.033, 5014.706, 5026.988, 
    5041.448,
  4863.202, 4874.433, 4887.021, 4898.099, 4910.616, 4916.373, 4933.011, 
    4933.328, 4949.613, 4959.87, 4971.336, 4982.407, 4995.694, 5008.487, 
    5020.583,
  4866.657, 4877.997, 4890.284, 4900.081, 4906.194, 4913.063, 4913.136, 
    4925.587, 4930.434, 4937.159, 4951.951, 4961.518, 4975.651, 4985.353, 
    4998.816,
  4880.504, 4892.444, 4900.126, 4905.713, 4904.756, 4901.388, 4902.225, 
    4898.824, 4905.143, 4916.284, 4924.382, 4937.066, 4950.653, 4963.241, 
    4976.166,
  4896.979, 4905.703, 4907.025, 4905.42, 4900.314, 4892.071, 4884.698, 
    4885.458, 4886.412, 4888.28, 4898.052, 4908.915, 4921.612, 4935.622, 
    4948.899,
  4906.92, 4906.905, 4900.812, 4894.42, 4882.476, 4870.154, 4861.287, 
    4856.424, 4857.297, 4865.143, 4871.135, 4879.997, 4892.807, 4907.222, 
    4922.131,
  4904.735, 4903.367, 4892.259, 4878.948, 4858.62, 4841.563, 4831.452, 
    4833.079, 4835.054, 4839.013, 4844.973, 4853.96, 4864.293, 4878.481, 
    4893.956,
  4897.462, 4888.017, 4873.159, 4853.865, 4832.206, 4817.455, 4808.111, 
    4805.358, 4808.203, 4815.508, 4821.676, 4829.702, 4840.31, 4854.694, 
    4870.648,
  4874.289, 4895.923, 4919.682, 4942.997, 4966.357, 4984.958, 5000.778, 
    5014.079, 5024.401, 5030.637, 5036.781, 5043.54, 5048.107, 5051.335, 
    5054.664,
  4854.52, 4873.731, 4895.395, 4918.846, 4940.454, 4961.029, 4979.506, 
    4990.689, 5001.056, 5013.269, 5020.009, 5028.953, 5034.799, 5041.618, 
    5044.562,
  4850.296, 4865.073, 4881.107, 4901.511, 4920.109, 4943.065, 4951.989, 
    4974.158, 4982.195, 4993.115, 5002.888, 5013.009, 5021.517, 5028.922, 
    5035.483,
  4863.864, 4870.108, 4879.534, 4890.971, 4906.029, 4917.292, 4939.862, 
    4942.469, 4961.719, 4974.253, 4986.419, 4996.063, 5007.404, 5017.034, 
    5026.382,
  4884.568, 4884.091, 4886.003, 4890.783, 4897.331, 4909.863, 4915.548, 
    4935.052, 4943.892, 4953.042, 4968.639, 4978.449, 4991.764, 5002.202, 
    5015.64,
  4900.384, 4898.246, 4895.984, 4896.741, 4896.868, 4900.273, 4909.668, 
    4913.578, 4924.917, 4940.98, 4950.319, 4963.908, 4976.3, 4989.571, 5003.83,
  4909.497, 4905.47, 4901.655, 4898.531, 4897.511, 4897.169, 4898.292, 
    4906.393, 4914.71, 4922.193, 4935.302, 4948.701, 4961.625, 4976.407, 
    4991.751,
  4897.491, 4891.467, 4886.399, 4883.066, 4878.514, 4877.608, 4879.754, 
    4883.574, 4892.352, 4907.406, 4920.812, 4934.213, 4948.952, 4964.435, 
    4980.241,
  4883.344, 4877.138, 4868.092, 4859.899, 4852.488, 4848.592, 4848.771, 
    4856.902, 4869.05, 4883.791, 4901.189, 4919.21, 4935.341, 4951.846, 
    4968.281,
  4871.889, 4862.064, 4851.967, 4842.752, 4833.058, 4826.252, 4823.57, 
    4825.134, 4835.813, 4856.416, 4880.12, 4901.978, 4921.417, 4938.983, 
    4955.301,
  4880.137, 4885.191, 4898.547, 4921.685, 4953.523, 4986.65, 5019.658, 
    5053.098, 5082.953, 5107.693, 5131.026, 5153.288, 5170.657, 5185.031, 
    5194.908,
  4883.574, 4882.078, 4887.257, 4903.662, 4927.61, 4960.776, 4996.169, 
    5026.35, 5056.328, 5088.221, 5112.25, 5134.625, 5152.387, 5168.627, 
    5176.943,
  4892.368, 4887.552, 4886.56, 4894.633, 4909.615, 4941.823, 4967.749, 
    5009.217, 5036.984, 5064.447, 5090.99, 5114.375, 5133.569, 5148.226, 
    5160.836,
  4899.952, 4891.761, 4890.89, 4891.681, 4902, 4913.858, 4953.004, 4971.647, 
    5011.617, 5043.073, 5071.425, 5093.773, 5115.377, 5131.291, 5143.072,
  4899.112, 4892.182, 4889.05, 4889.468, 4896.011, 4910.839, 4923.072, 
    4962.575, 4992.295, 5018.073, 5050.646, 5073.208, 5096.421, 5111.479, 
    5126.14,
  4887.312, 4880.222, 4880.715, 4885.966, 4890.812, 4899.589, 4918.224, 
    4932.436, 4964.6, 5001.922, 5027.973, 5055.077, 5076.821, 5094.774, 
    5108.142,
  4877.951, 4866.574, 4866.845, 4873.35, 4884.117, 4893.714, 4905.279, 
    4926.98, 4952.974, 4976.383, 5008.312, 5035.493, 5057.204, 5076.228, 
    5089.989,
  4874.233, 4860.826, 4854.77, 4860.145, 4870.652, 4884.194, 4896.738, 
    4908.69, 4929.109, 4960.745, 4990.332, 5016.363, 5040.136, 5059.252, 
    5073.834,
  4877.256, 4862.632, 4853.063, 4850.198, 4856.123, 4869.731, 4883.986, 
    4903.531, 4923.606, 4944.937, 4971.929, 4999.774, 5023.369, 5042.887, 
    5058.696,
  4880.977, 4862.992, 4850.587, 4845.422, 4843.975, 4852.795, 4866.663, 
    4883.549, 4903.554, 4929.959, 4957.912, 4985.126, 5009.313, 5029.626, 
    5046.263,
  4888.061, 4883.078, 4894.118, 4906.678, 4920.168, 4932.75, 4945.669, 
    4963.853, 4987.19, 5014.395, 5046.465, 5082.549, 5118.226, 5154.585, 
    5188.473,
  4895.812, 4890.301, 4894.559, 4908.191, 4921.203, 4935.53, 4952.296, 
    4968.957, 4991.32, 5022.529, 5054.27, 5089.408, 5123.854, 5160.155, 
    5191.614,
  4902.174, 4896.803, 4897.08, 4908.808, 4922.18, 4941.375, 4955.072, 
    4979.015, 5003.82, 5029.614, 5061.327, 5094.018, 5129.738, 5161.868, 
    5194.208,
  4903.588, 4901.442, 4900.761, 4907.694, 4923.731, 4936.335, 4963.188, 
    4977.158, 5004.275, 5033.672, 5065.771, 5097.665, 5132.235, 5165.823, 
    5195.653,
  4898.86, 4894.347, 4901.297, 4907.437, 4920.832, 4940.719, 4957.083, 
    4984.937, 5012.656, 5035.758, 5067.879, 5099.696, 5134.504, 5163.98, 
    5193.603,
  4896.977, 4886.451, 4892.247, 4903.918, 4917.963, 4934.862, 4959.326, 
    4979.585, 5003.497, 5038.17, 5066.817, 5101.13, 5133.978, 5166.257, 
    5192.564,
  4892.847, 4883.62, 4883.253, 4896.375, 4913.643, 4932.913, 4951.918, 
    4979.825, 5009.144, 5034.97, 5066.692, 5099.876, 5131.887, 5162.681, 
    5189.142,
  4893.554, 4880.292, 4877.584, 4888.564, 4905.356, 4925.575, 4947.867, 
    4967.951, 4994.353, 5028.856, 5062.365, 5095.341, 5128.723, 5159.399, 
    5185.863,
  4894.21, 4881.104, 4875.655, 4881.432, 4897.839, 4918.652, 4940.369, 
    4964.613, 4992.306, 5020.834, 5053.933, 5088.957, 5122.211, 5152.859, 
    5179.49,
  4901.508, 4884.496, 4875.251, 4877.931, 4890.705, 4910.428, 4933.655, 
    4953.537, 4977.442, 5009.034, 5044.677, 5081.063, 5115.163, 5146.729, 
    5173.714,
  4923.603, 4917.463, 4909.653, 4900.937, 4891.984, 4883.74, 4877.111, 
    4877.938, 4886.26, 4895.984, 4910.355, 4931.065, 4956.036, 4983.99, 
    5015.356,
  4926.397, 4921.628, 4912.511, 4901.866, 4890.254, 4879.087, 4872.461, 
    4872.333, 4879.182, 4896.875, 4916.635, 4941.479, 4968.61, 5000.859, 
    5032.114,
  4931.536, 4926.45, 4919.622, 4908.82, 4895.249, 4886.729, 4875.382, 
    4880.913, 4894.558, 4909.787, 4931.727, 4958.528, 4988.353, 5018.542, 
    5052.77,
  4935.269, 4933.688, 4929.85, 4918.799, 4911.735, 4896.303, 4899.244, 
    4896.443, 4908.633, 4929.314, 4955.541, 4981.945, 5013.558, 5046.23, 
    5080.625,
  4940.602, 4940.935, 4941.438, 4936.84, 4932.092, 4927.589, 4924.259, 
    4927.884, 4949.074, 4959.658, 4986.876, 5012.226, 5045.185, 5073.641, 
    5107.488,
  4946.198, 4950.02, 4952.884, 4953.641, 4953.253, 4952.36, 4958.327, 
    4964.252, 4972.95, 4997.552, 5020.057, 5047.166, 5075.833, 5106.02, 
    5133.055,
  4954.391, 4958.776, 4965.305, 4970.986, 4975.466, 4982.122, 4986.444, 
    4999.195, 5016.796, 5032.622, 5053.079, 5078.597, 5104.341, 5131.433, 
    5155.499,
  4962.824, 4968.481, 4976.162, 4985.431, 4991.83, 5001.691, 5013.608, 
    5025.247, 5037.891, 5059.003, 5080.898, 5104.687, 5129.906, 5154.062, 
    5175.239,
  4973.542, 4978.132, 4987.302, 4998.35, 5008.415, 5019.708, 5031.202, 
    5048.232, 5066.117, 5084.084, 5103.614, 5127.526, 5150.458, 5172.064, 
    5190.21,
  4985.647, 4987.097, 4994.513, 5007.088, 5017.94, 5032.385, 5046.864, 
    5062.182, 5078.84, 5099.912, 5122.4, 5145.658, 5167.72, 5188.297, 5204.586,
  4922.211, 4903.181, 4884.238, 4871.526, 4867.901, 4874.566, 4885.814, 
    4894.698, 4905.692, 4919.621, 4938.085, 4958.261, 4977.532, 4996.636, 
    5014.867,
  4919.37, 4893.636, 4868.749, 4851.191, 4846.628, 4856.365, 4876.026, 
    4888.543, 4899.998, 4918.277, 4937.095, 4955.53, 4972.152, 4989.997, 
    5005.716,
  4924.99, 4894.036, 4866.147, 4845.595, 4839.003, 4852.26, 4868.346, 
    4886.546, 4904.933, 4920.767, 4938.826, 4954.487, 4970.228, 4983.835, 
    5000.255,
  4939.134, 4907.154, 4878.93, 4855.833, 4850.451, 4852.279, 4874.414, 
    4887.219, 4905.036, 4923.884, 4942.634, 4956.073, 4970.576, 4984.233, 
    5001.086,
  4961.394, 4930.369, 4902.317, 4882.191, 4869.844, 4876.483, 4880.581, 
    4898.626, 4919.968, 4932.221, 4949.437, 4960.73, 4975.421, 4989.023, 
    5009.42,
  4991.92, 4962.422, 4934.49, 4914.834, 4901.94, 4897.902, 4909.338, 
    4917.669, 4927.542, 4946.273, 4959.549, 4974.277, 4990.276, 5008.591, 
    5026.711,
  5025.896, 5002.097, 4976.816, 4956.301, 4943.251, 4938.085, 4935.7, 
    4947.056, 4961.383, 4972.865, 4987.055, 5002.747, 5018.301, 5034.319, 
    5051.33,
  5058.432, 5042.542, 5023.613, 5008.024, 4993.87, 4988.596, 4989.495, 
    4992.181, 4998.746, 5012.639, 5025.01, 5037.973, 5051.1, 5064.731, 
    5077.508,
  5085.945, 5075.192, 5061.739, 5050.477, 5041.354, 5036.15, 5034.132, 
    5039.186, 5045.65, 5052.387, 5060.545, 5070.484, 5079.543, 5088.312, 
    5096.844,
  5109.011, 5101.945, 5094.163, 5086.016, 5078.923, 5075.566, 5074.421, 
    5074.515, 5077.127, 5083.124, 5088.965, 5094.573, 5099.691, 5104.584, 
    5108.665,
  4896.062, 4888.802, 4898.074, 4913.99, 4930.31, 4942.751, 4951.557, 
    4957.786, 4963.261, 4968.803, 4978.539, 4994.399, 5023.328, 5063.2, 
    5103.405,
  4916.868, 4903.36, 4903.459, 4914.43, 4929.399, 4941.377, 4950.833, 
    4955.738, 4957.034, 4962.104, 4970.137, 4982.615, 5006.031, 5046.769, 
    5086.364,
  4946.878, 4930.339, 4924.928, 4929.59, 4937.478, 4948.49, 4950.48, 
    4951.955, 4954.632, 4959.063, 4966.081, 4974.953, 4994.309, 5027.802, 
    5070.559,
  4978.835, 4960.106, 4950.799, 4946.607, 4950.53, 4947.674, 4951.29, 
    4950.42, 4954.051, 4960.319, 4967.106, 4972.402, 4987.723, 5018.53, 
    5058.889,
  5013.327, 4992, 4976.547, 4967.175, 4960.404, 4960.434, 4957.063, 4956.97, 
    4963.971, 4966.339, 4972.01, 4974.591, 4987.354, 5009.381, 5048.003,
  5050.185, 5027.917, 5007.641, 4994.547, 4982.295, 4972.914, 4971.021, 
    4971.179, 4971.211, 4976.318, 4979.276, 4982.087, 4991.928, 5011.813, 
    5042.125,
  5085.873, 5064.467, 5043.324, 5026.092, 5011.532, 5000.508, 4987.706, 
    4982.892, 4984.088, 4986.739, 4989.232, 4993.689, 5001.036, 5016.633, 
    5041.104,
  5117.467, 5098.617, 5078.031, 5061.883, 5045.684, 5032.285, 5020.166, 
    5009.901, 5001.616, 5000.73, 5002.918, 5007.671, 5015.501, 5028.472, 
    5047.365,
  5144.005, 5127.118, 5108.753, 5091.266, 5075.73, 5062.292, 5050.188, 
    5041.178, 5033.099, 5027.664, 5025.403, 5028.361, 5034.111, 5044.014, 
    5057.677,
  5166.811, 5150.376, 5135.017, 5119.276, 5102.335, 5088.536, 5076.758, 
    5067.367, 5059.401, 5054.358, 5051.221, 5051.508, 5054.887, 5062.078, 
    5071.973,
  4999.549, 4996.577, 4995.256, 4994.186, 4996.722, 5002.297, 5011.153, 
    5021.668, 5032.737, 5041.798, 5052.2, 5063.813, 5077.564, 5095.591, 
    5122.378,
  5014.455, 5007.77, 5006.241, 5004.413, 5006.122, 5009.509, 5018.381, 
    5027.069, 5036.678, 5048.784, 5060.535, 5074.784, 5089.984, 5112.499, 
    5139.061,
  5030.347, 5020.396, 5015.834, 5014.484, 5014.44, 5019.034, 5022.677, 
    5032.213, 5042.178, 5052.906, 5066.414, 5082.626, 5101.387, 5123.594, 
    5151.397,
  5055.673, 5038.375, 5026.24, 5020.188, 5019.267, 5019.403, 5026.509, 
    5031.034, 5040.028, 5052.881, 5067.287, 5084.926, 5106.702, 5132.218, 
    5160.714,
  5086.513, 5066.958, 5048.549, 5036.64, 5029.002, 5028.15, 5028.413, 
    5034.593, 5043.936, 5050.653, 5064.497, 5080.902, 5104.021, 5129.762, 
    5159.209,
  5115.772, 5095.848, 5074.79, 5059.426, 5046.39, 5040.304, 5038.536, 
    5039.913, 5041.416, 5051.274, 5058.158, 5072.192, 5093.819, 5123.356, 
    5154.12,
  5146.051, 5127.345, 5106.029, 5087.873, 5070.465, 5059.078, 5050.847, 
    5050.089, 5050.771, 5051.28, 5052.708, 5060.855, 5079.171, 5108.307, 
    5141.514,
  5172.796, 5154.453, 5134.199, 5116.771, 5097.424, 5080.835, 5067.167, 
    5057.943, 5052.643, 5051.787, 5050.008, 5051.458, 5066.152, 5093.69, 
    5128.191,
  5199.969, 5182.115, 5162.065, 5143.817, 5126.065, 5109.069, 5090.334, 
    5076.315, 5064.768, 5056.726, 5051.403, 5048.979, 5057.305, 5081.045, 
    5114.379,
  5225.374, 5204.339, 5183.971, 5165.216, 5145.801, 5129.869, 5113.841, 
    5096.729, 5080.194, 5067.453, 5057.742, 5052.896, 5056.222, 5074.798, 
    5105.613,
  5056.982, 5054.894, 5054.738, 5053.935, 5053.139, 5047.966, 5038.137, 
    5028.377, 5015.195, 4997.222, 4989.709, 4995.328, 5009.975, 5033.348, 
    5063.376,
  5069.632, 5064.238, 5063.719, 5061.454, 5061.051, 5053.077, 5048.083, 
    5028.768, 5009.311, 4992.959, 4982.855, 4988.734, 5005.139, 5031.507, 
    5062.513,
  5085.488, 5074.236, 5069.856, 5069.119, 5064.972, 5064.384, 5049.626, 
    5039.582, 5021.252, 4998.954, 4987.55, 4992.747, 5010.581, 5034.699, 
    5068.992,
  5109.509, 5091.43, 5079.542, 5072.045, 5071.888, 5063.823, 5062.079, 
    5044.386, 5025.04, 5012.361, 5003.882, 5009.152, 5026.232, 5052.677, 
    5087.774,
  5138.555, 5116.604, 5098.462, 5084.473, 5076.631, 5073.976, 5066.323, 
    5056.009, 5048.864, 5031.942, 5028.33, 5032.595, 5051.419, 5074.394, 
    5111.339,
  5164.241, 5142.763, 5121.489, 5103.804, 5089.351, 5078.965, 5076.666, 
    5068.227, 5057.356, 5053.982, 5053.095, 5060.326, 5078.71, 5106.538, 
    5138.9,
  5190.129, 5167.786, 5145.876, 5127.129, 5109.993, 5096.143, 5085.349, 
    5082.421, 5080.05, 5076.149, 5078.158, 5088.928, 5107.48, 5135.112, 
    5166.003,
  5210.85, 5191.609, 5169.226, 5148.632, 5129.129, 5114.153, 5102.77, 
    5094.544, 5090.954, 5095.27, 5102.154, 5115.772, 5136.47, 5162.562, 
    5189.994,
  5226.874, 5211.314, 5191.691, 5170.945, 5151.071, 5134.299, 5120.981, 
    5113.619, 5110.18, 5112.528, 5121.33, 5137.482, 5157.328, 5181.408, 
    5206.136,
  5236.729, 5225.25, 5208.844, 5189.157, 5167.882, 5150.527, 5137.893, 
    5128.533, 5123.637, 5124.953, 5133.471, 5149.138, 5169.375, 5191.818, 
    5215.317,
  5049.583, 5039.839, 5031.986, 5022.063, 5012.87, 5001.711, 4989.397, 
    4982.276, 4978.281, 4977.634, 4984.078, 4997.27, 5017.593, 5043.602, 
    5072.545,
  5047.871, 5036.729, 5028.675, 5018.814, 5008.952, 4992.546, 4986.921, 
    4970.6, 4965.548, 4967.926, 4978.176, 4994.569, 5016.677, 5046.19, 5073.53,
  5052.403, 5039.022, 5028.971, 5018.396, 5004.974, 4994.888, 4973.514, 
    4966.948, 4956.718, 4960.493, 4972.35, 4993.073, 5017.994, 5046.125, 
    5075.662,
  5060.045, 5045.542, 5032.798, 5019.412, 5005.371, 4985.77, 4973.862, 
    4958.939, 4952.298, 4956.217, 4972.552, 4994.409, 5022.08, 5052.967, 
    5082.738,
  5069.351, 5052.86, 5039.042, 5022.374, 5005.281, 4986.983, 4970.269, 
    4959.191, 4957.106, 4960.51, 4978.334, 5001.178, 5030.418, 5059.53, 
    5091.383,
  5080.956, 5063.904, 5045.799, 5028.718, 5009.169, 4991.446, 4977.797, 
    4968.504, 4964.434, 4973.553, 4990.515, 5014.071, 5042.562, 5074.117, 
    5102.63,
  5094.984, 5076.951, 5058.147, 5040.366, 5021.496, 5004.906, 4990.1, 
    4982.624, 4983.93, 4992.344, 5008.856, 5032.091, 5059.583, 5089.299, 
    5116.567,
  5111.271, 5093.664, 5075.762, 5057.1, 5038.703, 5023.385, 5012.065, 
    5004.824, 5004.854, 5015.652, 5032.875, 5055.733, 5082.602, 5109.31, 
    5133.731,
  5128.816, 5113.67, 5096.942, 5079.885, 5064.813, 5051.222, 5040.053, 
    5035.751, 5038.474, 5047.436, 5062.784, 5083.988, 5107.602, 5131.027, 
    5153.792,
  5148.208, 5134.423, 5120.151, 5105.674, 5091.862, 5082.073, 5075.51, 
    5071.981, 5074.193, 5083.321, 5097.691, 5116.199, 5135.955, 5156.016, 
    5176.792,
  5020.44, 5015.797, 5015.517, 5017.051, 5019.692, 5021.459, 5022.641, 
    5023.945, 5025.403, 5024.188, 5021.329, 5016.608, 5010.672, 5006.822, 
    5009.406,
  4997.392, 4992.236, 4992.062, 4995.917, 5001.352, 5005.501, 5011.68, 
    5013.122, 5014.563, 5017.035, 5014.553, 5010.617, 5005.613, 5006.157, 
    5011.151,
  4985.415, 4978.076, 4977.548, 4980.299, 4987.033, 4995.845, 4997.48, 
    5007.337, 5009.279, 5011.212, 5009.305, 5007.684, 5008.042, 5011.724, 
    5019.909,
  4979.259, 4971.548, 4970.419, 4972.293, 4978.978, 4984.201, 4994.228, 
    4997.154, 5002.082, 5006.191, 5009.573, 5012.688, 5019.702, 5026.627, 
    5037.805,
  4980.991, 4972.349, 4968.576, 4970.889, 4974.596, 4982.323, 4987.371, 
    4996.283, 5005.483, 5008.851, 5018.459, 5025.697, 5036.171, 5043.459, 
    5056.104,
  4987.994, 4978.557, 4972.806, 4974.21, 4976.74, 4983.045, 4992.062, 
    5000.588, 5008.732, 5022.549, 5033.464, 5044.303, 5054.319, 5063.757, 
    5073.782,
  5002.58, 4993.044, 4986.218, 4985.825, 4988.941, 4995.646, 5002.356, 
    5015.511, 5029.879, 5042.286, 5054.12, 5065.031, 5074.132, 5082.714, 
    5090.935,
  5025.882, 5015.406, 5007.798, 5006.685, 5008.552, 5016.812, 5027.422, 
    5038.737, 5050.786, 5065.006, 5076.359, 5085.871, 5094.006, 5101.073, 
    5108.118,
  5060.846, 5050.641, 5043.028, 5040.97, 5043.286, 5049.212, 5057.141, 
    5069.512, 5080.93, 5090.634, 5099.243, 5107.663, 5114.375, 5120.875, 
    5127.24,
  5100.164, 5089.464, 5082.19, 5078.452, 5078.474, 5083.437, 5090.801, 
    5098.505, 5106.952, 5115.834, 5123.638, 5130.527, 5136.498, 5142.307, 
    5147.607,
  4992.59, 5005.084, 5021.617, 5039.306, 5057.44, 5071.424, 5080.973, 
    5087.993, 5090.59, 5087.291, 5081.114, 5073.832, 5067.278, 5063.187, 
    5060.302,
  4971.395, 4982.998, 5000.405, 5021.354, 5040.846, 5058.668, 5072.468, 
    5078.511, 5079.946, 5078.689, 5070.841, 5063.54, 5056.085, 5051.228, 
    5044.502,
  4957.079, 4964.841, 4982.079, 5003.872, 5027.108, 5049.549, 5058.519, 
    5070.789, 5071.403, 5069.079, 5062.194, 5054.784, 5048.551, 5042.291, 
    5035.647,
  4952.689, 4957.973, 4973.242, 4992.608, 5016.605, 5033.85, 5053.942, 
    5055.372, 5062.135, 5058.892, 5055.634, 5051.837, 5048.698, 5042.401, 
    5036.209,
  4959.579, 4962.642, 4974.169, 4992.443, 5011.607, 5032.964, 5042.414, 
    5053.21, 5055.366, 5056.659, 5059.439, 5057.338, 5055.424, 5050.76, 
    5048.54,
  4977.043, 4979.247, 4986.169, 5001.25, 5016.201, 5029.923, 5043.769, 
    5049.757, 5056.918, 5063.57, 5066.136, 5066.714, 5065.168, 5063.303, 
    5061.045,
  4999.885, 5001.519, 5005.66, 5016.437, 5029.587, 5042.758, 5051.262, 
    5062.685, 5070.281, 5074.8, 5077.024, 5077.411, 5076.048, 5074.972, 
    5073.867,
  5031.78, 5032.29, 5034.383, 5042.435, 5050.172, 5061.452, 5070.522, 
    5077.066, 5081.759, 5086.557, 5087.884, 5088.232, 5087.211, 5085.828, 
    5084.562,
  5066.081, 5066.104, 5066.655, 5071.204, 5077.023, 5083.737, 5088.996, 
    5095.894, 5100.077, 5102.501, 5103.105, 5102.513, 5100.605, 5098.748, 
    5096.932,
  5100.73, 5098.539, 5098.268, 5100.058, 5102.837, 5107.942, 5112.515, 
    5115.574, 5117.644, 5119.064, 5118.546, 5117.071, 5114.66, 5111.984, 
    5109.354,
  4955.167, 4960.253, 4970.896, 4985.971, 5006.194, 5027.478, 5046.991, 
    5062.315, 5074.889, 5080.797, 5080.739, 5071.562, 5057.969, 5042.428, 
    5029.245,
  4949.076, 4954.425, 4966.125, 4982.89, 5003.609, 5025.229, 5044.648, 
    5059.185, 5070, 5076.426, 5074.282, 5064.938, 5052.196, 5039.263, 5025.288,
  4951.061, 4957.166, 4969.797, 4987.246, 5008.59, 5032.089, 5045.663, 
    5059.809, 5069.414, 5072.494, 5068.968, 5060.326, 5051.239, 5037.967, 
    5025.028,
  4960.643, 4966.526, 4981.466, 4997.839, 5020.856, 5034.204, 5052.437, 
    5058.16, 5066.798, 5066.582, 5064.214, 5059.839, 5053.166, 5044.123, 
    5033.432,
  4975.797, 4983.541, 4996.782, 5013.986, 5029.206, 5046.538, 5052.015, 
    5060.631, 5062.362, 5064.21, 5063.875, 5061.873, 5059.29, 5053.038, 
    5047.327,
  4996.845, 5003.387, 5012.926, 5027.948, 5039.575, 5047.143, 5053.686, 
    5056.814, 5059.09, 5063.838, 5065.562, 5065.538, 5064.129, 5062.484, 
    5059.453,
  5019.069, 5023.997, 5030.144, 5038.908, 5047.089, 5053.361, 5054.943, 
    5060.305, 5064.562, 5068.579, 5069.304, 5070.301, 5070.022, 5070.351, 
    5069.633,
  5042.219, 5043.089, 5044.726, 5050.208, 5053.043, 5057.271, 5061.564, 
    5065.395, 5068.356, 5071.855, 5073.334, 5074.55, 5074.554, 5075.549, 
    5076.525,
  5068.275, 5066.297, 5064.722, 5064.767, 5066.296, 5068.531, 5070.25, 
    5074.356, 5077.508, 5079.734, 5080.58, 5080.979, 5081.183, 5081.599, 
    5082.424,
  5094.41, 5088.48, 5084.038, 5081.845, 5079.743, 5079.751, 5081.316, 
    5082.806, 5084.32, 5086.285, 5087.798, 5088.555, 5088.421, 5088.632, 
    5089.146,
  5002.965, 4990.354, 4981.157, 4976.066, 4975.069, 4979.156, 4987.27, 
    5001.142, 5012.854, 5022.452, 5032.27, 5043.293, 5050.738, 5055.113, 
    5053.924,
  5004.357, 4990.907, 4980.304, 4975.286, 4975.941, 4982.004, 4997.098, 
    5008.7, 5017.165, 5028.413, 5038.344, 5046.646, 5051.406, 5053.225, 
    5050.022,
  5013.713, 5000.393, 4989.577, 4985.5, 4986.517, 4998.474, 5005.331, 
    5017.565, 5028.58, 5037.639, 5045.337, 5051.44, 5055.849, 5056.296, 
    5053.549,
  5027.64, 5015.298, 5007.521, 5001.761, 5006.846, 5009.119, 5022.679, 
    5028.283, 5037.548, 5045.729, 5053.807, 5059.043, 5063.708, 5063.062, 
    5059.22,
  5041.913, 5032.334, 5026.688, 5022.693, 5022.708, 5029.638, 5033.29, 
    5040.948, 5051.675, 5055.454, 5063.349, 5067.875, 5071.978, 5070.103, 
    5066.448,
  5051.778, 5044.827, 5039.332, 5037.125, 5037.68, 5039.013, 5047.396, 
    5052.849, 5057.459, 5065.748, 5072.17, 5077.392, 5079.882, 5078.54, 
    5073.369,
  5057.691, 5054.066, 5050.526, 5048.137, 5048.938, 5052.887, 5055.133, 
    5061.844, 5069.32, 5075.788, 5081.046, 5085.765, 5087.192, 5085.603, 
    5081.122,
  5061.25, 5058.107, 5054.991, 5055.301, 5056.19, 5060.014, 5065.842, 
    5071.103, 5076.378, 5083.532, 5089.155, 5093.065, 5094.636, 5093.584, 
    5090.206,
  5063.923, 5062.46, 5061.795, 5062.396, 5064.911, 5068.932, 5073.31, 
    5080.07, 5087.046, 5092.298, 5096.539, 5099.961, 5101.469, 5101.347, 
    5099.653,
  5062.651, 5060.265, 5062.045, 5065.734, 5069.932, 5075.867, 5082.885, 
    5089.08, 5094.706, 5100.373, 5105.097, 5108.678, 5110.978, 5112.088, 
    5111.638,
  5121.573, 5106.523, 5091.364, 5078.039, 5067.324, 5054.617, 5039.704, 
    5028.876, 5020.189, 5016.082, 5019.673, 5025.721, 5029.735, 5031.958, 
    5032.376,
  5113.419, 5100.753, 5089.072, 5080.852, 5074.169, 5062.471, 5055.392, 
    5043.863, 5034.344, 5030.792, 5029.373, 5030.394, 5030.771, 5030.68, 
    5029.617,
  5109.947, 5100.905, 5092.987, 5089.05, 5081.521, 5078.802, 5066.119, 
    5061.013, 5054.458, 5048.739, 5044.586, 5042.404, 5038.404, 5033.948, 
    5028.428,
  5109.875, 5102.833, 5098.969, 5094.375, 5092.947, 5085.603, 5083.701, 
    5075.27, 5066.911, 5062.587, 5057.459, 5050.981, 5043.868, 5034.732, 
    5025.579,
  5111.338, 5106.348, 5105.467, 5103.394, 5101.975, 5099.069, 5095.086, 
    5087.583, 5086.749, 5075.947, 5071.403, 5061.223, 5052.34, 5038.464, 
    5026.312,
  5114.22, 5111.536, 5110.86, 5111.149, 5110.893, 5108.435, 5106.818, 
    5102.432, 5095.29, 5090.368, 5082.976, 5073.513, 5063.141, 5050.481, 
    5037.604,
  5117.345, 5117.938, 5118.43, 5119.498, 5120.286, 5120.704, 5117.347, 
    5114.407, 5111.488, 5105.239, 5097.515, 5089.257, 5079.275, 5068.895, 
    5057.909,
  5122.359, 5123.77, 5124.931, 5127.749, 5128.747, 5129.434, 5128.905, 
    5126.443, 5122.029, 5118.22, 5112.69, 5105.873, 5097.97, 5089.7, 5081.27,
  5127.206, 5130.159, 5133.395, 5136.181, 5138.759, 5140.188, 5139.308, 
    5138.829, 5137.633, 5134.302, 5129.774, 5125.069, 5119.227, 5112.84, 
    5106.245,
  5132.674, 5135.803, 5140.133, 5143.983, 5146.796, 5149.065, 5151.209, 
    5151.56, 5150.712, 5149.506, 5147.579, 5144.621, 5140.867, 5136.466, 
    5131.823,
  5161.758, 5163.032, 5164.397, 5163.073, 5160.948, 5156.094, 5149.22, 
    5140.353, 5129.874, 5115.979, 5102.975, 5090.866, 5080.844, 5074.526, 
    5073.911,
  5149.686, 5150.412, 5152.024, 5151.489, 5150.048, 5146.122, 5141.991, 
    5131.201, 5119.084, 5107.246, 5092.338, 5078.155, 5064.994, 5059.106, 
    5059.27,
  5143.765, 5145.071, 5146.583, 5147.826, 5146.667, 5145.51, 5134.158, 
    5128.459, 5115.449, 5100.483, 5083.322, 5066.008, 5050.002, 5043.834, 
    5049.582,
  5144.526, 5146.294, 5148.15, 5148.593, 5146.903, 5141.354, 5136.108, 
    5123.052, 5111.125, 5096.625, 5078.145, 5057.877, 5040.996, 5035.047, 
    5043.34,
  5148.939, 5150.591, 5152.502, 5152.096, 5149.585, 5143.343, 5135.172, 
    5126.712, 5115.344, 5096.865, 5080.278, 5059.43, 5044.95, 5039.012, 
    5048.126,
  5154.922, 5156.55, 5156.886, 5156.092, 5151.856, 5146.691, 5139.891, 
    5129.677, 5117.148, 5104.048, 5087.912, 5072.031, 5060.563, 5056.663, 
    5062.304,
  5161.205, 5163.154, 5162.514, 5161.605, 5158.434, 5153.74, 5146.205, 
    5138.888, 5128.549, 5115.836, 5102.484, 5090.795, 5082.592, 5080.29, 
    5084.475,
  5168.011, 5169.332, 5168.691, 5168.154, 5164.879, 5161.372, 5155.994, 
    5148.255, 5139.034, 5130.084, 5120.789, 5112.593, 5107.774, 5107.326, 
    5111.446,
  5175.058, 5177.076, 5177.38, 5176.724, 5175.034, 5172.001, 5166.749, 
    5161.614, 5155.088, 5147.837, 5140.939, 5135.734, 5132.981, 5133.604, 
    5137.472,
  5182.898, 5183.713, 5185.109, 5185.699, 5184.776, 5183.021, 5179.595, 
    5174.451, 5169.232, 5164.962, 5161.308, 5158.868, 5158.082, 5160.115, 
    5165.031,
  5121.28, 5128.687, 5140.771, 5153.421, 5166.603, 5176.375, 5182.747, 
    5187.881, 5189.047, 5185.931, 5180.553, 5173.698, 5164.929, 5155.878, 
    5148.325,
  5123.11, 5128.114, 5135.242, 5144.225, 5151.555, 5157.734, 5164.546, 
    5164.877, 5163.562, 5161.378, 5153.304, 5145.576, 5135.055, 5129.417, 
    5122.15,
  5123.935, 5127.161, 5131.559, 5138.073, 5141.392, 5149.051, 5143.336, 
    5150.032, 5142.759, 5137.941, 5129.195, 5120.562, 5110.496, 5103.292, 
    5102.471,
  5126.884, 5127.981, 5130.905, 5132.637, 5135.337, 5134.174, 5139.373, 
    5130.048, 5129.671, 5121.746, 5112.422, 5101.561, 5095.066, 5093.847, 
    5098.446,
  5134.163, 5132.836, 5133.662, 5133.561, 5133.749, 5133.06, 5128.196, 
    5128.283, 5119.255, 5109.287, 5103.18, 5096.521, 5097.525, 5099.64, 
    5105.548,
  5140.957, 5138.716, 5137.017, 5136.101, 5133.794, 5131.906, 5128.563, 
    5120.873, 5115.457, 5111.313, 5107.677, 5107, 5109.042, 5112.345, 5116.579,
  5147.761, 5145.638, 5143.153, 5141.378, 5139.235, 5135.548, 5129.865, 
    5125.833, 5121.094, 5118.429, 5119.005, 5121.696, 5125.411, 5130.348, 
    5136.462,
  5154.894, 5152.441, 5149.098, 5146.39, 5142.872, 5140.199, 5136.217, 
    5132.181, 5131.251, 5133.863, 5138.013, 5143.739, 5150.593, 5157.601, 
    5165.191,
  5161.674, 5158.97, 5155.854, 5152.372, 5149.924, 5147.106, 5145.335, 
    5146.209, 5149.542, 5155.122, 5162.599, 5170.64, 5178.512, 5186.061, 
    5193.217,
  5168.857, 5164.362, 5160.404, 5156.89, 5154.646, 5155.137, 5157.817, 
    5163.086, 5170.944, 5180.214, 5189.521, 5198.191, 5205.703, 5211.443, 
    5214.864,
  5098.555, 5105.259, 5119.336, 5133.985, 5152.921, 5167.702, 5182.573, 
    5199.529, 5212.476, 5223.112, 5233.701, 5243.813, 5250.306, 5255.726, 
    5257.58,
  5106.96, 5110.175, 5120.171, 5133.119, 5145.974, 5160.708, 5178.495, 
    5188.565, 5202.008, 5214.984, 5221.599, 5228.82, 5231.562, 5234.692, 
    5231.377,
  5113.787, 5116.162, 5122.877, 5133.28, 5144.092, 5158.282, 5164.007, 
    5184.205, 5189.892, 5198.157, 5204.603, 5208.913, 5208.748, 5205.832, 
    5200.737,
  5118.217, 5118.246, 5124.33, 5129.444, 5139.972, 5146.537, 5162.265, 
    5163.265, 5178.148, 5184.25, 5186.082, 5185.073, 5181.812, 5177.011, 
    5168.769,
  5122.119, 5120.298, 5124.051, 5128.454, 5134.974, 5143.186, 5148.007, 
    5159.549, 5162.031, 5160.201, 5165.673, 5161.026, 5157.514, 5149.583, 
    5143.567,
  5128.963, 5124.001, 5122.129, 5124.131, 5127.59, 5132.62, 5140.21, 
    5141.477, 5146.273, 5150.796, 5147.981, 5144.712, 5141.281, 5136.028, 
    5131.422,
  5135.808, 5133.25, 5128.872, 5127.749, 5128.999, 5131.692, 5133.863, 
    5137.989, 5139.426, 5139.699, 5142.643, 5143.74, 5141.897, 5137.238, 
    5130.776,
  5145.709, 5138.263, 5133.587, 5131.292, 5131.457, 5134.806, 5139.671, 
    5143.83, 5148.592, 5153.607, 5153.931, 5151.961, 5148.832, 5143.828, 
    5136.952,
  5151.497, 5148.541, 5146.763, 5146.286, 5148.941, 5154.068, 5160.802, 
    5166.769, 5167.861, 5164.348, 5160.146, 5155.379, 5150.677, 5147.344, 
    5143.194,
  5151.39, 5152.242, 5155.017, 5160.131, 5167.292, 5175.171, 5181.21, 
    5182.143, 5178.732, 5171.893, 5161.334, 5150.322, 5142.947, 5141.101, 
    5142.624,
  5163.227, 5163.681, 5167.154, 5173.262, 5180.809, 5186.954, 5192.622, 
    5198.818, 5205.626, 5215.742, 5228.882, 5243.335, 5258.786, 5274.993, 
    5292.476,
  5164.986, 5166.438, 5169.963, 5177.634, 5187.004, 5193.779, 5201.75, 
    5205.893, 5212.937, 5223.358, 5232.878, 5245.351, 5258.236, 5272.721, 
    5285.882,
  5164.946, 5167.485, 5172.138, 5180.142, 5187.588, 5197.769, 5202.633, 
    5213.163, 5217.151, 5223.039, 5231.576, 5241.426, 5252.739, 5263.504, 
    5275.63,
  5162.313, 5166.256, 5172.71, 5178.923, 5188.46, 5195.346, 5205.209, 
    5208.288, 5216.97, 5223.944, 5229.568, 5236.735, 5245.167, 5254.381, 
    5261.846,
  5158.536, 5160.812, 5170.306, 5178.277, 5186.619, 5194.117, 5199.918, 
    5207.819, 5211.654, 5212.967, 5218.625, 5221.891, 5228.671, 5233.885, 
    5242.17,
  5158.057, 5157.441, 5165.757, 5175.032, 5184.221, 5191.12, 5196.292, 
    5197.544, 5200.441, 5203.604, 5204.919, 5206.436, 5210.464, 5214.007, 
    5219.136,
  5162.809, 5157.838, 5164.128, 5174.273, 5182.487, 5188.234, 5190.174, 
    5190.53, 5187.737, 5182.15, 5179.67, 5178.886, 5181.14, 5185.227, 5191.382,
  5168.272, 5162.25, 5169.355, 5176.277, 5184.662, 5188.961, 5190.051, 
    5184.79, 5177.558, 5169.929, 5162.564, 5157.735, 5158.608, 5162.306, 
    5167.961,
  5174.474, 5178.04, 5183.854, 5192.533, 5199.237, 5201.88, 5197.746, 
    5189.201, 5175.936, 5160.528, 5147.644, 5141.273, 5139.771, 5144.171, 
    5150.369,
  5190.683, 5196.871, 5204.034, 5210.367, 5212.825, 5211.44, 5203.855, 
    5190.152, 5171.299, 5150.648, 5131.533, 5119.916, 5118.203, 5123.701, 
    5132.322,
  5280.925, 5268.982, 5259.799, 5253.287, 5248.632, 5243.238, 5237.778, 
    5234.409, 5231.646, 5231.621, 5235.208, 5241.167, 5250.329, 5261.221, 
    5276.143,
  5271.608, 5260.789, 5253.829, 5249.393, 5247.806, 5245.321, 5244.613, 
    5242.062, 5240.88, 5240.013, 5239.34, 5241.652, 5245.752, 5255.075, 
    5266.279,
  5260.241, 5251.288, 5244.333, 5242.75, 5243.91, 5246.794, 5246.462, 
    5247.465, 5246.885, 5246.199, 5245.855, 5245.577, 5247.205, 5250.767, 
    5260.484,
  5246.836, 5239.375, 5233.165, 5231.811, 5236.07, 5241.318, 5246.963, 
    5246.895, 5247.885, 5248.408, 5248.647, 5249.143, 5250.985, 5253.462, 
    5259.227,
  5233.062, 5226.293, 5221.283, 5222.186, 5227.786, 5237.706, 5241.217, 
    5247.973, 5247.533, 5247.749, 5247.008, 5246.588, 5248.282, 5251.233, 
    5257.272,
  5218.768, 5213.044, 5209.008, 5212.272, 5219.219, 5230.753, 5238.175, 
    5240.167, 5242.439, 5242.861, 5240.814, 5239.862, 5240.117, 5243.292, 
    5248.675,
  5205.698, 5201.354, 5200.544, 5208.503, 5217.851, 5228.599, 5234.514, 
    5238.812, 5237.681, 5234.041, 5229.582, 5225.748, 5223.633, 5225.524, 
    5231.789,
  5195.578, 5193.968, 5198.33, 5207.663, 5216.598, 5226.543, 5231.909, 
    5233.105, 5230.606, 5226.983, 5220.451, 5213.839, 5207.676, 5205.286, 
    5208.993,
  5190.369, 5193.062, 5202.078, 5212.464, 5222.098, 5230.167, 5232.546, 
    5231.705, 5228.278, 5223.114, 5216.11, 5206.053, 5194.956, 5186.41, 
    5185.779,
  5190.554, 5199.219, 5209.647, 5218.729, 5226.019, 5229.077, 5229.273, 
    5226.783, 5225.048, 5221.531, 5212.714, 5199.047, 5183.156, 5170.339, 
    5165.331,
  5284.223, 5292.753, 5300.054, 5303.064, 5303.104, 5302.048, 5301.346, 
    5301.06, 5296.824, 5293.356, 5293.651, 5298.333, 5304.034, 5309.219, 
    5313.639,
  5261.095, 5272.433, 5282.558, 5288.803, 5290.755, 5290.648, 5293.145, 
    5293.363, 5292.953, 5291.775, 5287.514, 5288.23, 5290.042, 5295.711, 
    5297.871,
  5237.865, 5252.467, 5264.717, 5274.755, 5278.841, 5282.836, 5281.76, 
    5288.643, 5288.876, 5289.151, 5288.013, 5285.702, 5283.598, 5281.879, 
    5282.423,
  5215.643, 5232.836, 5246.892, 5258.258, 5265.118, 5268.3, 5275.72, 
    5275.028, 5282.009, 5284.745, 5285.428, 5284.035, 5282.144, 5278.838, 
    5274.104,
  5195.825, 5213.978, 5230.551, 5243.521, 5252.38, 5258.463, 5262.128, 
    5271.781, 5275.314, 5278.531, 5281.747, 5279.083, 5274.425, 5268.629, 
    5264.305,
  5180.408, 5198.949, 5215.478, 5229.116, 5237.943, 5245.049, 5252.667, 
    5257.864, 5267.044, 5274.025, 5275.093, 5271.896, 5266.517, 5259.272, 
    5251.99,
  5168.172, 5187.63, 5204.623, 5217.853, 5227.877, 5235.694, 5243.176, 
    5252.825, 5261.653, 5267.437, 5269.54, 5266.594, 5260.763, 5251.101, 
    5239.498,
  5160.568, 5179.689, 5195.022, 5207.675, 5217.434, 5226.907, 5235.875, 
    5244.491, 5255.07, 5262.845, 5265.136, 5265.038, 5258.501, 5245.395, 
    5228.009,
  5155.269, 5174.049, 5189.504, 5202.298, 5212.533, 5221.875, 5231.618, 
    5242.625, 5252.79, 5260.051, 5265.62, 5264.907, 5255.876, 5239.815, 
    5217.98,
  5154.264, 5170.814, 5184.468, 5196.968, 5207.076, 5217.374, 5228.004, 
    5238.647, 5249.475, 5259.628, 5265.595, 5264.119, 5254.375, 5236.646, 
    5211.36,
  5224.07, 5231.092, 5242.814, 5256.864, 5271.896, 5283.762, 5292.431, 
    5300.063, 5304.688, 5306.195, 5306.774, 5304.82, 5301.457, 5299.094, 
    5299.934,
  5210.066, 5216.489, 5226.953, 5241.089, 5255.167, 5268.026, 5280.374, 
    5286.644, 5292.809, 5297.914, 5299.792, 5299.589, 5297.238, 5294.498, 
    5292.139,
  5195.246, 5202.621, 5213.088, 5227.097, 5241.858, 5256.613, 5264.759, 
    5278.927, 5283.701, 5288.276, 5292.035, 5294.312, 5293.24, 5290.286, 
    5286.298,
  5178.535, 5185.963, 5198.222, 5211.612, 5227.281, 5240.134, 5257.332, 
    5262.017, 5274.195, 5280.195, 5284.772, 5286.987, 5287.46, 5284.223, 
    5278.517,
  5163.324, 5170.114, 5182.332, 5197.751, 5213.047, 5229.935, 5240.609, 
    5258.587, 5264.683, 5270.285, 5276.654, 5279.676, 5279.91, 5275.178, 
    5268.277,
  5149.918, 5156.099, 5166.429, 5181.608, 5197.768, 5214.102, 5231.358, 
    5242.002, 5254.321, 5264.165, 5268.975, 5272.699, 5272.382, 5266.889, 
    5257.405,
  5139.286, 5146.372, 5155.593, 5168.993, 5186.031, 5202.706, 5218.104, 
    5234.927, 5246.393, 5254.716, 5262.524, 5266.621, 5265.843, 5258.944, 
    5245.394,
  5130.531, 5139.909, 5148.155, 5158.916, 5173.311, 5191.454, 5208.126, 
    5222.181, 5234.788, 5247.282, 5255.969, 5261.24, 5260.859, 5251.779, 
    5233.146,
  5124.778, 5134.888, 5144.596, 5154.921, 5167.907, 5183.689, 5199.897, 
    5215.754, 5228.479, 5240.383, 5250.845, 5258.265, 5257.64, 5245.722, 
    5222.207,
  5124.791, 5132.935, 5141.433, 5150.682, 5163.209, 5178.55, 5194.164, 
    5207.315, 5220.977, 5235.763, 5248.266, 5256.954, 5256.334, 5241.926, 
    5217.946,
  5261.351, 5232.215, 5206.916, 5188.038, 5179.811, 5181.411, 5191.453, 
    5205.039, 5221.08, 5238.297, 5255.713, 5269.536, 5278.342, 5281.751, 
    5282.405,
  5246.909, 5217.633, 5194.149, 5178.246, 5171.256, 5175.606, 5187.634, 
    5200.309, 5216.023, 5234.176, 5249.654, 5262.03, 5270.742, 5275.071, 
    5275.467,
  5231.266, 5203.673, 5183.116, 5170.54, 5166.811, 5173.343, 5181.823, 
    5199.99, 5213.651, 5229.091, 5243.532, 5255.345, 5262.695, 5266.479, 
    5267.267,
  5214.208, 5189.209, 5171.363, 5161.718, 5162.35, 5167.701, 5182.848, 
    5192.551, 5210.036, 5225.624, 5238.208, 5248.125, 5254.829, 5257.788, 
    5256.412,
  5198.398, 5176.996, 5162.311, 5155.836, 5158.6, 5167.818, 5177.844, 
    5195.77, 5209.936, 5220.577, 5233.669, 5241.584, 5247.028, 5247.771, 
    5245.375,
  5183.382, 5166.25, 5153.801, 5150.014, 5154.738, 5164.55, 5178.224, 
    5190.478, 5203.733, 5219.113, 5228.345, 5235.743, 5239.67, 5238.7, 
    5233.538,
  5171.595, 5160.349, 5150.062, 5148.397, 5153.695, 5164.464, 5175.388, 
    5191.625, 5205.233, 5215.676, 5224.496, 5231.185, 5232.822, 5230.356, 
    5220.952,
  5163.983, 5156.633, 5149.121, 5148.251, 5152.036, 5163.105, 5174.136, 
    5186.791, 5198.877, 5212.193, 5220.821, 5227.183, 5227.472, 5223.297, 
    5209.093,
  5160.325, 5155.65, 5153.222, 5149.618, 5153.049, 5161.478, 5172.292, 
    5185.883, 5198.643, 5209.926, 5218.291, 5224.083, 5224.151, 5216.205, 
    5200.155,
  5158.605, 5155.879, 5154.904, 5151.257, 5151.28, 5158.663, 5170.002, 
    5181.402, 5193.562, 5206.273, 5216.674, 5221.39, 5221.484, 5211.698, 5200,
  5329.404, 5314.024, 5296.086, 5273.505, 5248.91, 5223.325, 5200.719, 
    5185.137, 5176.155, 5176.073, 5186.512, 5208.991, 5235.299, 5255.67, 
    5271.803,
  5300.101, 5286.966, 5270.922, 5250.234, 5227.81, 5203.36, 5189.404, 
    5176.119, 5169.811, 5174.31, 5185.816, 5207.967, 5232.438, 5252.435, 
    5265.949,
  5269.369, 5259.351, 5245.31, 5229.196, 5207.465, 5194.706, 5173.106, 
    5172.772, 5167.493, 5174.267, 5186.167, 5206.829, 5229.043, 5246.141, 
    5259.214,
  5238.444, 5231.156, 5220.052, 5205.776, 5189.077, 5172.52, 5169.064, 
    5158.683, 5164.131, 5172.739, 5187, 5205.816, 5225.403, 5241.23, 5250.453,
  5214.453, 5208.575, 5200.008, 5186.958, 5173.537, 5163.874, 5155.411, 
    5160.784, 5164.599, 5172.897, 5188.01, 5204.807, 5221.643, 5233.562, 
    5241.341,
  5196.021, 5190.72, 5181.91, 5170.334, 5158.451, 5151.626, 5151.195, 
    5154.569, 5162.088, 5175.348, 5188.358, 5204.094, 5217.531, 5227.202, 
    5232.084,
  5184.492, 5177.397, 5168.784, 5157.341, 5149.664, 5146.615, 5148.63, 
    5156.866, 5167.105, 5177.347, 5190.294, 5203.322, 5214.541, 5221.106, 
    5221.707,
  5174.906, 5167.372, 5157.059, 5146.966, 5141.881, 5144.031, 5149.049, 
    5156.86, 5167.121, 5179.807, 5192.005, 5203.094, 5211.741, 5216.185, 
    5213.028,
  5166.773, 5159.101, 5150.527, 5143.182, 5141.696, 5145.615, 5151.235, 
    5161.724, 5172.839, 5183.521, 5193.762, 5203.676, 5210.312, 5211.314, 
    5206.531,
  5162.898, 5156.768, 5149.689, 5142.787, 5141.639, 5145.812, 5153.62, 
    5163.317, 5174.053, 5185.223, 5195.166, 5203.628, 5208.695, 5208.328, 
    5208.727,
  5299.877, 5282.601, 5268.4, 5254.344, 5242.774, 5231.41, 5221.241, 
    5214.553, 5209.832, 5205.539, 5205.786, 5209.023, 5218.341, 5233.542, 
    5250.92,
  5264.499, 5245.264, 5229.787, 5215.469, 5204.59, 5194.181, 5191.034, 
    5184.559, 5182.557, 5182.969, 5184.471, 5189.601, 5200.416, 5218.928, 
    5237.736,
  5229.304, 5211.25, 5195.804, 5184.011, 5175.467, 5174.316, 5164.348, 
    5168.713, 5164.54, 5165.502, 5168.014, 5174.371, 5186.153, 5204.763, 
    5226.524,
  5207.233, 5189.781, 5175.617, 5166.413, 5160.687, 5155.489, 5158.016, 
    5150.884, 5152.856, 5153.242, 5156.317, 5162.911, 5175.727, 5195.744, 
    5218.286,
  5194.023, 5178.649, 5166.063, 5156.387, 5150.901, 5148.385, 5144.308, 
    5146.864, 5143.811, 5143.204, 5148.94, 5155.831, 5170.297, 5188.708, 
    5212.271,
  5189.025, 5173.279, 5158.73, 5149.152, 5141.367, 5138.575, 5137.467, 
    5135.186, 5137.337, 5141.081, 5145.595, 5154.875, 5168.848, 5188.616, 
    5211.387,
  5188.367, 5172.499, 5157.221, 5145.969, 5138.028, 5131.881, 5128.335, 
    5129.56, 5133.187, 5138.303, 5147.238, 5158.806, 5173.668, 5192.401, 
    5213.748,
  5191.822, 5174.665, 5157.434, 5144.448, 5134.22, 5128.11, 5125.341, 
    5127.055, 5133.513, 5143.695, 5155.254, 5167.99, 5182.867, 5200.271, 
    5218.439,
  5199.071, 5182.357, 5164.514, 5150.212, 5141.174, 5134.738, 5131.53, 
    5135.375, 5142.979, 5153.261, 5165.726, 5178.491, 5192.592, 5207.811, 
    5222.838,
  5209.89, 5192.328, 5174.096, 5158.61, 5147.256, 5142.109, 5141.481, 
    5144.967, 5152.865, 5164.373, 5175.881, 5188.737, 5201.44, 5214.707, 
    5227.057,
  5290.714, 5265.595, 5242.954, 5219.83, 5199.88, 5182.759, 5168.401, 
    5160.407, 5155.033, 5149.311, 5146.408, 5145.779, 5149.804, 5159.324, 
    5174.772,
  5275.08, 5249.563, 5225.666, 5201.51, 5181.108, 5161.359, 5153.55, 
    5143.517, 5140.459, 5137.169, 5133.726, 5132.515, 5134.923, 5144.339, 
    5159.456,
  5267.179, 5242.339, 5216.998, 5193.536, 5170.531, 5156.806, 5142.132, 
    5140.553, 5136.224, 5132.599, 5127.861, 5126.593, 5128.106, 5135.194, 
    5150.536,
  5266.771, 5240.742, 5214.497, 5189.839, 5168.593, 5148.989, 5143.413, 
    5136.184, 5133.135, 5129.421, 5124.834, 5123.604, 5126.951, 5136.151, 
    5151.787,
  5271.043, 5245.254, 5219.82, 5194.994, 5173.577, 5156.274, 5142.77, 
    5138.367, 5134.571, 5129.502, 5125.338, 5125.439, 5130.619, 5140.484, 
    5157.799,
  5279.924, 5252.936, 5225.91, 5202.821, 5179.653, 5160.863, 5149.317, 
    5140.147, 5134.415, 5130.995, 5128.94, 5131.034, 5138.141, 5150.696, 
    5166.672,
  5291.735, 5266.067, 5238.228, 5215.41, 5194.715, 5175.312, 5157.396, 
    5147.48, 5139.859, 5135.017, 5134.297, 5139.071, 5147.437, 5160.696, 
    5177.071,
  5307.157, 5280.443, 5251.384, 5227.854, 5206.26, 5188.791, 5172.019, 
    5158.105, 5147.775, 5143.738, 5143.795, 5149.416, 5159.507, 5174.068, 
    5192.177,
  5324.995, 5299.105, 5270.285, 5245.259, 5224.179, 5206.66, 5189.6, 
    5176.853, 5165.697, 5159.062, 5158.409, 5164.431, 5175.52, 5191.149, 
    5210.254,
  5345.164, 5316, 5286.816, 5260.562, 5236.012, 5219.5, 5206.709, 5194.662, 
    5183.879, 5178.068, 5177.891, 5183.971, 5195.471, 5211.193, 5229.139,
  5301.953, 5271.786, 5242.655, 5212.382, 5183.648, 5157.846, 5132.897, 5117, 
    5103.785, 5090.821, 5082.248, 5076.817, 5075.032, 5079.283, 5090.469,
  5316.898, 5284.203, 5252.131, 5220.143, 5190.825, 5159.662, 5141.202, 
    5117.434, 5102.518, 5093.87, 5086.806, 5082.393, 5079.798, 5084.012, 
    5093.497,
  5335.024, 5301.002, 5266.694, 5234.693, 5200.332, 5176.776, 5143.415, 
    5129.763, 5112.869, 5099.873, 5091.737, 5088.473, 5087.063, 5090.515, 
    5100.78,
  5354.527, 5318.663, 5283.107, 5246.886, 5216.404, 5181.57, 5161.892, 
    5134.555, 5116.485, 5107.182, 5099.996, 5095.536, 5096.374, 5101.11, 
    5114.659,
  5375.239, 5339.075, 5303.296, 5265.738, 5232.904, 5201.932, 5173.193, 
    5152.478, 5138.874, 5119.824, 5114.56, 5108.676, 5112.21, 5117.062, 
    5132.385,
  5394.145, 5358.34, 5321.09, 5284.784, 5249.38, 5217.709, 5193.84, 5169.551, 
    5150.662, 5140.382, 5133.372, 5130.032, 5133.05, 5140.638, 5154.11,
  5410.727, 5378.216, 5341.966, 5305.912, 5271.626, 5239.608, 5211.939, 
    5194.126, 5178.551, 5165.798, 5157.668, 5156.271, 5158.832, 5166.965, 
    5179.1,
  5423.658, 5392.641, 5358.22, 5324.109, 5290.111, 5258.76, 5232.817, 5214.1, 
    5199.362, 5190.485, 5185.535, 5184.147, 5187.535, 5195.03, 5205.98,
  5434.565, 5405.707, 5374.673, 5342.495, 5310.74, 5280.013, 5252.26, 
    5235.581, 5224.846, 5216.115, 5211.488, 5211.582, 5214.98, 5221.677, 
    5230.385,
  5441.305, 5411.133, 5381.808, 5353.583, 5323.104, 5296.387, 5271.246, 
    5251.798, 5241.72, 5237.285, 5235.295, 5236.599, 5239.604, 5245.241, 
    5251.759,
  5277.076, 5247.836, 5216.808, 5180.212, 5144.789, 5112.677, 5080.955, 
    5059.109, 5043.912, 5030.458, 5022.54, 5017.792, 5015.929, 5017.196, 
    5024.673,
  5276.079, 5247.922, 5218.382, 5183.034, 5149.541, 5114.352, 5091.035, 
    5063.965, 5044.635, 5032.934, 5023.572, 5018.229, 5016.433, 5020.639, 
    5028.449,
  5275.671, 5249.473, 5222.779, 5190.652, 5156.547, 5133.54, 5097.035, 
    5079.865, 5060.758, 5045.458, 5034, 5028.615, 5027.687, 5032.177, 5041.015,
  5275.52, 5250.786, 5228.766, 5196.826, 5170.781, 5139.266, 5122.386, 
    5095.796, 5077.693, 5065.484, 5057.501, 5051.143, 5052.786, 5057.307, 
    5069.265,
  5275.383, 5253.47, 5236.048, 5207.536, 5184.474, 5159.991, 5139.938, 
    5119.529, 5112.008, 5093.537, 5089.276, 5082.492, 5086.608, 5088.921, 
    5100.715,
  5275.772, 5256.287, 5241.163, 5218.69, 5197.282, 5176.486, 5162.243, 
    5146.601, 5132.092, 5125.363, 5120.328, 5117.081, 5119.25, 5123.602, 
    5132.049,
  5276.582, 5260.585, 5248.171, 5231.368, 5213.914, 5198.298, 5182.669, 
    5172.565, 5164.861, 5157.797, 5152.53, 5151.91, 5153.02, 5157.118, 
    5163.034,
  5279.379, 5265.903, 5255.19, 5243.278, 5227.477, 5215.698, 5205.5, 
    5197.657, 5188.978, 5186.045, 5183.965, 5183.314, 5184.528, 5188.075, 
    5192.452,
  5284.127, 5272.947, 5263.821, 5256.408, 5244.726, 5235.72, 5225.835, 
    5221.931, 5217.916, 5214.922, 5212.625, 5213.238, 5213.977, 5216.398, 
    5218.822,
  5290.878, 5280.296, 5272.539, 5267.445, 5257.151, 5251.967, 5247.009, 
    5243.732, 5240.024, 5239.374, 5239.049, 5239.804, 5240.725, 5243.089, 
    5245.011,
  5181.213, 5165.707, 5147.877, 5124.596, 5098.744, 5070.687, 5040.175, 
    5020.875, 5006.39, 4997.396, 4996.369, 5001.143, 5008.67, 5019.099, 
    5032.034,
  5185.78, 5172.559, 5155.232, 5135.476, 5112.388, 5083.059, 5062.489, 
    5036.297, 5016.018, 5005.978, 5000.773, 5002.261, 5006.658, 5016.105, 
    5026.66,
  5194.965, 5182.864, 5167.637, 5152.509, 5127.826, 5113.97, 5078.095, 
    5063.412, 5044.352, 5026.621, 5013.227, 5008.041, 5008.537, 5014.177, 
    5023.266,
  5207.421, 5196.143, 5184.649, 5167.127, 5153.189, 5125.216, 5113.686, 
    5086.418, 5066.127, 5051.029, 5037.935, 5023.922, 5019.124, 5018.937, 
    5026.245,
  5221.472, 5211.93, 5203.301, 5188.83, 5174.386, 5156.493, 5133.798, 
    5111.339, 5099.83, 5073.503, 5061.846, 5045.642, 5037.104, 5030.146, 
    5033.904,
  5236.907, 5229.935, 5221.106, 5210.859, 5196.684, 5179.15, 5163.37, 
    5141.115, 5117.638, 5101.219, 5083.645, 5067.942, 5056.393, 5047.772, 
    5046.276,
  5253.056, 5248.203, 5240.855, 5232.852, 5222.241, 5208.303, 5188.37, 
    5170.11, 5150.764, 5128.842, 5108.544, 5091.911, 5077.341, 5067.111, 
    5062.055,
  5270.267, 5266.625, 5260.157, 5254.4, 5244.261, 5233.113, 5218.73, 
    5199.972, 5177.371, 5156.708, 5135.798, 5116.93, 5100.632, 5088.787, 
    5081.41,
  5287.468, 5284.554, 5279.844, 5275.311, 5268.991, 5258.991, 5244.539, 
    5229.816, 5211.833, 5190.079, 5166.862, 5146.459, 5128.106, 5114.115, 
    5104.545,
  5304.691, 5301.423, 5298.469, 5294.277, 5287.302, 5280.476, 5270.786, 
    5256.317, 5238.766, 5220.237, 5199.234, 5178.144, 5158.897, 5143.478, 
    5132.234,
  5205.749, 5193.532, 5179.445, 5161.033, 5140.401, 5117.3, 5088.255, 
    5063.886, 5040.306, 5018.733, 5007.248, 5004.081, 5009.648, 5025.249, 
    5057.521,
  5217.974, 5206.022, 5190.184, 5170.512, 5149.305, 5120.64, 5097.61, 
    5063.713, 5037.722, 5017.867, 5004.323, 5000.265, 5001.923, 5015.911, 
    5040.54,
  5231.077, 5220.166, 5204.024, 5186.277, 5158.966, 5139.417, 5101.046, 
    5078.111, 5049.405, 5023.958, 5005.856, 4999.877, 5000.361, 5008.289, 
    5028.614,
  5244.874, 5233.803, 5219.079, 5197.899, 5176.897, 5143.587, 5121.902, 
    5084.442, 5055.05, 5032.221, 5013.006, 5002.527, 5002.755, 5008.612, 
    5024.378,
  5256.275, 5246.324, 5233.193, 5213.017, 5190.679, 5163.384, 5130.922, 
    5102.028, 5078.166, 5043.819, 5024.608, 5008.356, 5007.37, 5008.464, 
    5022.1,
  5265.747, 5256.458, 5242.658, 5225.095, 5201.525, 5174.479, 5146.704, 
    5114.284, 5085.792, 5062.79, 5037.904, 5019.478, 5013.745, 5014.045, 
    5022.994,
  5272.661, 5264.86, 5252.042, 5235.416, 5213.76, 5187.149, 5156.807, 
    5130.768, 5107.076, 5081.318, 5056.713, 5034.785, 5022.412, 5020.045, 
    5024.157,
  5278.31, 5270.23, 5257.871, 5242.07, 5219.439, 5193.73, 5166.081, 5139.041, 
    5115.379, 5095.945, 5075.074, 5053.231, 5035.928, 5028.536, 5029.606,
  5282.304, 5274.96, 5262.767, 5247.205, 5225.574, 5199.399, 5171.586, 
    5148.961, 5128.98, 5110.901, 5090.987, 5071.273, 5053.454, 5039.604, 
    5034.933,
  5285.681, 5276.804, 5265.063, 5248.35, 5224.809, 5200.521, 5175.444, 
    5152.102, 5132.92, 5118.441, 5104.35, 5087.191, 5070.495, 5056.384, 
    5045.317,
  5207.026, 5206.018, 5201.89, 5192.436, 5179.86, 5162.428, 5140.527, 
    5120.168, 5099.689, 5079.863, 5064.806, 5053.165, 5047.684, 5046.605, 
    5054.798,
  5208.872, 5204.125, 5194.618, 5181.52, 5164.428, 5141.893, 5124.52, 
    5098.109, 5079.306, 5064.755, 5048.892, 5038.46, 5029.694, 5028.39, 
    5032.027,
  5206.172, 5197.858, 5183.958, 5168.969, 5147.061, 5131.199, 5098.546, 
    5084.953, 5064.311, 5052.116, 5037.788, 5025.804, 5015.592, 5010.864, 
    5012.654,
  5200.735, 5188.344, 5171.638, 5152.023, 5130.794, 5104.49, 5089.841, 
    5061.719, 5053.663, 5043.66, 5030.373, 5014.593, 5003.843, 4996.5, 
    4997.617,
  5193.568, 5177.947, 5159.711, 5137.519, 5115.517, 5094.081, 5069.093, 
    5060.223, 5048.595, 5038.655, 5024.634, 5006.002, 4994.068, 4984.552, 
    4985.484,
  5186.042, 5168.397, 5147.694, 5125.624, 5102.113, 5081.444, 5066.041, 
    5051.365, 5044.79, 5037.286, 5020.575, 5001.609, 4987.69, 4978.187, 
    4976.536,
  5180.286, 5162.122, 5141.185, 5119.433, 5098.429, 5078.398, 5061.954, 
    5054.792, 5048.038, 5036.928, 5020.875, 5001.164, 4985.146, 4975.674, 
    4972.411,
  5178.208, 5159.989, 5138.831, 5117.124, 5095.263, 5076.89, 5064.441, 
    5054.505, 5047.639, 5039.653, 5024.39, 5004.942, 4987.75, 4978.075, 
    4974.875,
  5180.236, 5163.01, 5142.448, 5121.256, 5100.419, 5081.877, 5067.286, 
    5060.582, 5053.672, 5044.274, 5030.518, 5012.561, 4994.616, 4984.027, 
    4981.346,
  5186.395, 5169.28, 5150.088, 5128.602, 5105.966, 5087.63, 5073.727, 
    5063.249, 5056.46, 5048.839, 5037.792, 5022.589, 5005.34, 4993.229, 
    4989.929,
  5169.21, 5166.477, 5162.876, 5158.297, 5154.098, 5149.624, 5145.339, 
    5143.601, 5140.547, 5136.88, 5134.933, 5133.12, 5131.82, 5130.841, 
    5130.922,
  5163.226, 5155.919, 5146.833, 5137.865, 5128.483, 5120.356, 5116.166, 
    5109.62, 5106.374, 5104.894, 5100.696, 5100.267, 5098.006, 5099.718, 
    5098.1,
  5153.208, 5141.942, 5127.473, 5114.59, 5099.705, 5092.96, 5077.326, 
    5078.304, 5069.716, 5068.727, 5066.91, 5067.997, 5067.292, 5067.971, 
    5068.485,
  5146.741, 5132.203, 5114.682, 5097.497, 5081.697, 5067.042, 5064.434, 
    5050.907, 5050.829, 5048.049, 5047.398, 5047.189, 5046.393, 5046, 5044.082,
  5146.613, 5130.707, 5112.276, 5092.198, 5075.696, 5063.109, 5049.763, 
    5048.396, 5040.877, 5037.964, 5037.576, 5034.446, 5031.319, 5026.28, 
    5024.013,
  5150.572, 5134.167, 5113.948, 5093.773, 5073.646, 5059.208, 5049.481, 
    5038.672, 5034.621, 5033.084, 5028.68, 5023.716, 5017.179, 5009.608, 
    5003.917,
  5157.772, 5142.156, 5121.975, 5100.334, 5080.409, 5061.788, 5047.174, 
    5039.623, 5032.055, 5025.216, 5020.398, 5013.389, 5003.746, 4993.718, 
    4985.015,
  5165.862, 5149.727, 5129.851, 5108.352, 5085.082, 5064.942, 5048.493, 
    5034.93, 5025.204, 5018.637, 5011.107, 5002.361, 4991.068, 4979.066, 
    4968.548,
  5173.159, 5157.971, 5138.818, 5117.293, 5094.298, 5071.332, 5050.824, 
    5035.55, 5022.291, 5011.073, 5001.394, 4991.141, 4978.632, 4966.145, 
    4955.288,
  5178.775, 5162.21, 5144.094, 5124.111, 5100.062, 5076.431, 5054.097, 
    5033.377, 5016.879, 5004.214, 4992.855, 4981.422, 4968.57, 4955.883, 
    4945.305,
  5176.677, 5174.774, 5172.436, 5168.506, 5163.885, 5157.759, 5151.833, 
    5149.626, 5145.755, 5141.632, 5142.724, 5146.204, 5152.428, 5159.802, 
    5170.776,
  5172.997, 5167.647, 5161.17, 5152.725, 5143.58, 5133.863, 5126.527, 
    5114.926, 5110.811, 5110.276, 5106.891, 5109.692, 5113.004, 5123.432, 
    5130.566,
  5173.832, 5167.334, 5158.632, 5149.172, 5136.616, 5126.722, 5109.558, 
    5105.577, 5089.813, 5081.65, 5077.82, 5077.139, 5078.627, 5083.71, 
    5093.238,
  5178.16, 5169.941, 5159.597, 5147.321, 5133.318, 5116.855, 5105.07, 
    5081.735, 5075.144, 5063.921, 5053.031, 5048.282, 5047.798, 5051.338, 
    5057.488,
  5181.764, 5172.605, 5161.153, 5145.903, 5128.918, 5110.528, 5088.382, 
    5074.864, 5051.791, 5038.19, 5030.298, 5021.884, 5021.786, 5020.954, 
    5028.113,
  5184.753, 5173.664, 5158.27, 5140.905, 5118.679, 5096.391, 5072.636, 
    5045.334, 5026.529, 5012.053, 4998.292, 4993.469, 4994.555, 4997.297, 
    5003.654,
  5187.003, 5173.863, 5155.532, 5133.572, 5108.75, 5079.145, 5048.737, 
    5020.182, 4992.216, 4970.474, 4960.436, 4957.865, 4961.041, 4969.314, 
    4978.635,
  5188.986, 5171.362, 5149.054, 5123.221, 5091.254, 5056.298, 5017.594, 
    4978.71, 4948.213, 4927.114, 4915.074, 4914.167, 4923.495, 4937.762, 
    4953.167,
  5189.586, 5170.719, 5145.904, 5115.021, 5078.036, 5033.466, 4983.671, 
    4941.27, 4903.599, 4877.963, 4867.857, 4872.523, 4886.357, 4906.236, 
    4926.127,
  5191.289, 5168.387, 5139.475, 5103.917, 5058.377, 5007.437, 4951.351, 
    4900.434, 4858.631, 4833.828, 4824.925, 4834.258, 4854.272, 4879.576, 
    4903.47,
  5221.204, 5219.215, 5217.509, 5217.266, 5217.519, 5217.478, 5215.975, 
    5219.054, 5217.405, 5213.406, 5212.906, 5213.454, 5213.498, 5214.994, 
    5217.69,
  5223.806, 5222.071, 5218.052, 5215.012, 5208.769, 5204.589, 5200.268, 
    5188.722, 5184.46, 5182.908, 5175.195, 5172.708, 5170.335, 5172.727, 
    5171.844,
  5230.106, 5227.7, 5221.917, 5215.686, 5205.215, 5197.289, 5179.865, 
    5179.954, 5161.855, 5151.88, 5145.066, 5140.34, 5136.092, 5135.061, 
    5137.581,
  5234.863, 5228.495, 5218.709, 5205.906, 5192.304, 5174.228, 5164.267, 
    5135.045, 5128.021, 5113.705, 5100.204, 5092.999, 5089.581, 5089.603, 
    5092.484,
  5236.061, 5226.157, 5212.754, 5195.688, 5174.237, 5154.283, 5127.425, 
    5114.936, 5084.837, 5063.354, 5050.224, 5036.559, 5033.847, 5031.51, 
    5039.73,
  5233.63, 5219.366, 5200.083, 5176.783, 5151.245, 5124.156, 5095.506, 
    5060.471, 5034.526, 5012.609, 4989.654, 4975.961, 4969.625, 4969.086, 
    4978.125,
  5229.216, 5211.201, 5186.622, 5159.78, 5128.576, 5094.137, 5057.283, 
    5023.195, 4989.057, 4959.435, 4939.426, 4922.613, 4911.79, 4909.905, 
    4917.704,
  5222.595, 5198.779, 5170.962, 5137.908, 5101.475, 5061.122, 5018.405, 
    4979.638, 4949.655, 4924.425, 4897.914, 4875.183, 4860.157, 4854.859, 
    4862.441,
  5214.409, 5189.567, 5157.275, 5119.53, 5077.868, 5031.424, 4989.052, 
    4957.514, 4924.639, 4890.745, 4859.467, 4831.384, 4810.374, 4802.063, 
    4809.179,
  5208.348, 5176.404, 5140.372, 5099.14, 5052.715, 5007.918, 4968.866, 
    4935.001, 4900.52, 4866.274, 4831.014, 4797.889, 4772.998, 4762.443, 
    4770.412,
  5300.206, 5294.299, 5288.229, 5280.356, 5271.519, 5260.518, 5245.934, 
    5236.986, 5225.402, 5210.868, 5202.72, 5197.891, 5195.594, 5196.188, 
    5200.839,
  5292.26, 5287.211, 5280.448, 5271.963, 5260.386, 5245.601, 5235.147, 
    5211.934, 5198.604, 5188.946, 5175.079, 5167.486, 5162.359, 5163.585, 
    5164.939,
  5285.209, 5280.58, 5271.962, 5262.538, 5246.159, 5234.303, 5205.354, 
    5199.122, 5172.942, 5154.94, 5141.805, 5132.183, 5124.663, 5122.552, 
    5125.196,
  5277.69, 5271.563, 5261.306, 5245.971, 5228.766, 5203.207, 5189.173, 
    5150.684, 5135.679, 5116.489, 5100.04, 5088.367, 5081.325, 5078.136, 
    5079.178,
  5270.542, 5261.544, 5248.336, 5229.809, 5205.402, 5180.545, 5146.451, 
    5130.54, 5099.598, 5072.513, 5059.277, 5042.592, 5035.976, 5028.647, 
    5031.553,
  5261.182, 5248.733, 5230.625, 5206.179, 5178.078, 5146.467, 5115.667, 
    5078.941, 5054.813, 5035.268, 5014.575, 4999.439, 4990.37, 4983.073, 
    4982.512,
  5251.204, 5234.787, 5210.601, 5183.749, 5151.183, 5114.701, 5081.548, 
    5055.279, 5026.915, 4998.669, 4979.045, 4963.158, 4951.694, 4943.787, 
    4939.634,
  5238.157, 5215.891, 5189.542, 5156.525, 5120.022, 5086.511, 5055.26, 
    5021.786, 4992.23, 4968.372, 4948.381, 4933.242, 4921.959, 4911.344, 
    4903.004,
  5222.806, 5199.342, 5168.076, 5132.888, 5097.841, 5065.295, 5032.617, 
    5000.404, 4968.372, 4943.505, 4926.929, 4913.806, 4899.879, 4884.695, 
    4870.182,
  5207.846, 5178.85, 5146.496, 5110.908, 5078.821, 5046.993, 5011.089, 
    4973.111, 4945.22, 4928.851, 4915.74, 4900.852, 4882.352, 4860.514, 
    4837.609,
  5350.989, 5355.964, 5357.429, 5353.867, 5347.85, 5338.058, 5324.455, 
    5313.105, 5295.044, 5270.035, 5246.187, 5220.782, 5195.291, 5169.375, 
    5148.402,
  5334.287, 5339.408, 5339.382, 5335.522, 5327.742, 5316.244, 5305.569, 
    5281.059, 5260.561, 5241.791, 5212.076, 5184.712, 5155.312, 5133.287, 
    5107.344,
  5316.577, 5321.747, 5319.862, 5317.191, 5306.828, 5299.45, 5273.882, 
    5267.074, 5235.318, 5206.426, 5176.985, 5147.761, 5116.62, 5090.592, 
    5066.726,
  5298.355, 5302.204, 5300.965, 5295.464, 5286.603, 5268.831, 5258.263, 
    5219.608, 5198.537, 5169.454, 5138.578, 5108.759, 5078.373, 5053.095, 
    5030.447,
  5280.176, 5283.023, 5281.553, 5275.542, 5263.8, 5249.214, 5220.683, 
    5207.621, 5172.549, 5133.554, 5105.671, 5070.289, 5043.084, 5017.12, 
    5000.405,
  5262.756, 5264.642, 5261.814, 5254.25, 5239.96, 5220.655, 5197.654, 
    5160.604, 5130.32, 5100.634, 5066.45, 5036.21, 5012.394, 4991.463, 
    4976.073,
  5248.354, 5248.671, 5243.954, 5233.366, 5217.999, 5194.455, 5166.295, 
    5139.073, 5105.604, 5067.841, 5036.305, 5009.9, 4988.003, 4969.885, 
    4954.361,
  5237.078, 5233.788, 5225.835, 5212.915, 5192.651, 5167.91, 5138.543, 
    5103.14, 5068.263, 5036.491, 5009.358, 4987.465, 4969.305, 4951.737, 
    4934.76,
  5224.616, 5219.382, 5208.619, 5191.777, 5169.761, 5141.818, 5110.889, 
    5078.124, 5043.233, 5013.233, 4990.746, 4971.641, 4952.592, 4933.157, 
    4913.713,
  5211.508, 5202.288, 5189.028, 5170.757, 5145.329, 5116.066, 5082.984, 
    5046.002, 5016.06, 4994.72, 4975.93, 4957.159, 4937.322, 4916.093, 4893.84,
  5246.489, 5260, 5274.195, 5286.835, 5299.531, 5308.977, 5318.171, 5326.925, 
    5331.749, 5331.82, 5330.799, 5325.519, 5315.507, 5300.158, 5282.018,
  5231.547, 5246.124, 5259.509, 5272.93, 5282.873, 5293.929, 5302.421, 
    5306.375, 5309.792, 5312.928, 5306.354, 5299.314, 5285.434, 5270.875, 
    5247.541,
  5212.735, 5228.574, 5242.795, 5256.345, 5267.218, 5278.337, 5280.346, 
    5292.039, 5288.39, 5286.073, 5280.765, 5270.875, 5254.031, 5234.291, 
    5210.665,
  5192.14, 5208.606, 5224.226, 5236.993, 5248.851, 5255.284, 5267.704, 
    5259.097, 5267.073, 5261.091, 5251.78, 5238.096, 5220.872, 5198.043, 
    5171.31,
  5170.477, 5186.929, 5203.246, 5216.917, 5227.987, 5237.115, 5238.081, 
    5248.321, 5239.366, 5230.64, 5223.709, 5204.454, 5185.652, 5157.104, 
    5133.61,
  5151.44, 5165.694, 5181.694, 5195.85, 5206.259, 5213.582, 5218.937, 
    5212.975, 5212.957, 5205.405, 5188.738, 5169.148, 5146.139, 5118.743, 
    5093.23,
  5136.136, 5147.065, 5161.234, 5174.055, 5184.785, 5190.858, 5193.308, 
    5195.117, 5186.629, 5172.106, 5157.187, 5133.536, 5107.394, 5079.903, 
    5053.763,
  5127.656, 5134.857, 5144.783, 5156.273, 5164.895, 5170.608, 5171.483, 
    5165.853, 5157.663, 5144.672, 5121.335, 5095.949, 5069.665, 5042.563, 
    5015.924,
  5121.689, 5128.118, 5135.603, 5143.091, 5148.604, 5151.583, 5150.466, 
    5145.591, 5131.563, 5110.492, 5087.42, 5062.138, 5033.942, 5006.214, 
    4979.304,
  5121.573, 5126.467, 5130.935, 5135.298, 5138.192, 5137.553, 5131.309, 
    5119.018, 5102.116, 5081.108, 5054.777, 5028.071, 5001.28, 4975.146, 
    4947.213,
  5070.486, 5073.565, 5080.797, 5090.636, 5104.85, 5120.699, 5140.559, 
    5165.574, 5190.327, 5210.774, 5228.364, 5244.318, 5256.688, 5268.252, 
    5278.448,
  5058.879, 5062.389, 5069.442, 5079.27, 5089.709, 5104.338, 5121.936, 
    5140.128, 5162.59, 5186.892, 5204.241, 5220.552, 5233.281, 5245.477, 
    5252.1,
  5051.671, 5055.039, 5062.383, 5072.784, 5082.998, 5097.635, 5108.03, 
    5128.365, 5142.734, 5161.459, 5179.976, 5195.785, 5208.504, 5216.599, 
    5226.062,
  5045.761, 5048.508, 5058.209, 5068.327, 5080.363, 5089.626, 5106.532, 
    5113.026, 5131.224, 5144.93, 5159.578, 5172.092, 5183.183, 5191.58, 
    5195.32,
  5041.613, 5043.901, 5054.335, 5066.537, 5078.508, 5091.508, 5099.708, 
    5112.888, 5121.675, 5130.17, 5142.517, 5149.736, 5158.386, 5161.24, 
    5166.016,
  5041.955, 5040.413, 5051.783, 5064.968, 5078.435, 5088.821, 5100.739, 
    5105.482, 5114.028, 5122.208, 5127.371, 5131.333, 5135.049, 5134.618, 
    5134.488,
  5044.365, 5041.981, 5049.704, 5063.271, 5076.849, 5087.438, 5094.679, 
    5102.232, 5106.306, 5106.908, 5109.805, 5108.988, 5107.589, 5102.983, 
    5098.198,
  5050.209, 5046.398, 5050.72, 5061.187, 5072.051, 5080.263, 5086.388, 
    5088.522, 5090.031, 5091.205, 5088.154, 5083.77, 5077.779, 5069.724, 
    5059.73,
  5059.25, 5055.692, 5055.112, 5060.345, 5066.641, 5072.294, 5074.803, 
    5076.042, 5072.992, 5067.064, 5060.603, 5052.889, 5042.475, 5030.333, 
    5016.101,
  5070.359, 5065.338, 5062.986, 5063.005, 5063.142, 5063.623, 5061.916, 
    5057.397, 5051.546, 5044.131, 5034.063, 5021.854, 5007.96, 4991.885, 
    4973.485,
  5033.944, 5017.806, 5003.918, 4992.293, 4982.29, 4974.183, 4968.271, 
    4969.061, 4976.799, 4989.065, 5006.152, 5026.237, 5045.485, 5065.402, 
    5087.038,
  5024.259, 5008.662, 4995.59, 4983.206, 4972.511, 4961.97, 4957.198, 
    4950.917, 4954.191, 4967.054, 4983.552, 5005.396, 5026.664, 5050.236, 
    5069.506,
  5019.288, 5004.672, 4992.141, 4980.878, 4968.3, 4958.402, 4945.97, 
    4944.196, 4940.91, 4947.91, 4963.314, 4985.849, 5008.832, 5031.613, 
    5054.442,
  5017.223, 5003.494, 4991.809, 4978.809, 4967.391, 4955.332, 4947.098, 
    4936.276, 4932.558, 4935.461, 4946.8, 4967.365, 4991.693, 5015.999, 
    5037.529,
  5017.44, 5004.528, 4994.105, 4981.482, 4970.748, 4959.606, 4949.243, 
    4940.472, 4935.936, 4931.302, 4939.326, 4952.923, 4976.065, 4997.716, 
    5020.508,
  5019.136, 5005.625, 4994.458, 4983.072, 4972.749, 4964.198, 4956.873, 
    4947.348, 4940.661, 4938.021, 4939.122, 4946.349, 4961.941, 4980.761, 
    4999.847,
  5022.317, 5008.912, 4996.119, 4984.402, 4974.186, 4965.849, 4959.507, 
    4955.965, 4951.886, 4947.147, 4945.596, 4948.063, 4955.53, 4967.102, 
    4980.73,
  5028.324, 5012.341, 4996.805, 4983.253, 4970.625, 4961.466, 4956.495, 
    4952.8, 4950.504, 4950.325, 4949.74, 4950.171, 4951.547, 4955.576, 
    4961.351,
  5035.765, 5019.423, 5001.088, 4984.431, 4968.211, 4956.52, 4948.789, 
    4945.82, 4944.181, 4942.624, 4941.637, 4941.616, 4941.626, 4942.152, 
    4942.655,
  5044.276, 5025.252, 5005.7, 4986.743, 4967.852, 4953.366, 4943.768, 
    4937.36, 4933.734, 4931.682, 4929.492, 4926.797, 4923.136, 4919.119, 
    4914.616,
  5075.027, 5068.882, 5062.326, 5053.927, 5044.554, 5031.743, 5014.509, 
    5000.851, 4985.784, 4969.611, 4959.016, 4951.369, 4945.744, 4942.164, 
    4941.431,
  5062.641, 5056.536, 5049.079, 5039.353, 5027.36, 5009.977, 4997.31, 
    4974.658, 4959.877, 4948.246, 4935.321, 4927.317, 4919.914, 4917.646, 
    4913.404,
  5053.876, 5046.534, 5037.188, 5027.559, 5011.063, 4998.722, 4971.464, 
    4964.446, 4943.455, 4929.479, 4915.593, 4907.286, 4898.439, 4893.311, 
    4890.701,
  5045.617, 5037.841, 5028.183, 5014.498, 4997.562, 4975.525, 4964.341, 
    4938.906, 4928.728, 4917.004, 4902.817, 4891.38, 4881.697, 4875.509, 
    4870.874,
  5037.938, 5030.011, 5020.686, 5005.111, 4986.577, 4966.91, 4944.408, 
    4936.06, 4920.797, 4904.449, 4893.368, 4879.067, 4869.684, 4861.02, 
    4858.698,
  5029.316, 5022.878, 5012.805, 4997.693, 4977.343, 4955.191, 4937.924, 
    4918.303, 4906.849, 4898.262, 4883.683, 4870.32, 4859.738, 4852.511, 
    4849.948,
  5020.304, 5015.663, 5006.887, 4994.852, 4974.443, 4949.83, 4928.349, 
    4915.586, 4901.959, 4886.708, 4874.192, 4861.641, 4850.992, 4845.201, 
    4843.831,
  5012.272, 5009.162, 5003.2, 4990.672, 4967.947, 4944.434, 4923.143, 
    4904.009, 4888.2, 4876.204, 4862.273, 4850.253, 4841.06, 4835.163, 4834.95,
  5004.723, 5002.777, 4997.598, 4985.499, 4967.295, 4942.983, 4919.515, 
    4900.333, 4881.603, 4863.218, 4847.268, 4834.556, 4825.357, 4821.519, 
    4822.884,
  5003.381, 4999.12, 4994.162, 4983.373, 4963.901, 4942.129, 4918.021, 
    4893.616, 4871.179, 4850.89, 4831.959, 4816.227, 4805.233, 4800.321, 
    4802.162,
  5078.076, 5088.17, 5098.341, 5106.371, 5113.229, 5117.208, 5119.141, 
    5119.875, 5114.986, 5105.646, 5095.616, 5084.51, 5072.472, 5061.064, 
    5051.945,
  5058.603, 5066.913, 5074.988, 5082.759, 5087.475, 5091.922, 5094.613, 
    5090.214, 5084.989, 5079.707, 5066.433, 5055.145, 5041.863, 5033.732, 
    5022.043,
  5047.484, 5053.487, 5058.773, 5064.987, 5067.855, 5074.227, 5065.905, 
    5070.747, 5057.78, 5048.113, 5036.51, 5025.069, 5011.575, 5000.425, 
    4991.459,
  5040.892, 5045.021, 5048.432, 5051.197, 5052.796, 5049.796, 5053.727, 
    5036.703, 5033.745, 5021.921, 5006.118, 4991.342, 4977.32, 4965.04, 
    4953.34,
  5037.441, 5040.042, 5041.827, 5042.375, 5041.942, 5038.813, 5028.338, 
    5024.853, 5005.619, 4986.982, 4973.22, 4952.204, 4936.676, 4919.599, 
    4910.032,
  5037.642, 5036.922, 5035.381, 5033.308, 5027.395, 5021.144, 5011.345, 
    4991.472, 4973.907, 4954.183, 4929.738, 4907.71, 4889.083, 4872.378, 
    4862.059,
  5041.148, 5038.402, 5033.144, 5028.02, 5020.202, 5008.255, 4990.795, 
    4971.958, 4946.36, 4918.154, 4894.025, 4869.769, 4848.348, 4831.869, 
    4821.594,
  5049.535, 5043.188, 5035.259, 5026.338, 5012.307, 4995.973, 4975.28, 
    4949.693, 4923.504, 4897.301, 4868.286, 4840.542, 4816.343, 4798.064, 
    4788.062,
  5061.209, 5052.869, 5041.754, 5029.4, 5013.41, 4994.213, 4971.441, 4946.53, 
    4916.546, 4882.969, 4850.478, 4818.382, 4790.266, 4770.148, 4759.896,
  5075.93, 5064.222, 5051.691, 5037.286, 5018.63, 4998.426, 4973.644, 
    4943.603, 4911.607, 4876.9, 4840.899, 4805.164, 4774.208, 4751.412, 
    4739.828,
  5051.277, 5057.664, 5072.805, 5092.708, 5116.441, 5137.491, 5158.846, 
    5179.927, 5198.32, 5213.203, 5225.749, 5235.376, 5240.582, 5242.003, 
    5240.519,
  5052.652, 5058.632, 5067.631, 5085.196, 5104, 5124.311, 5144.148, 5160.524, 
    5176.511, 5193.561, 5202.585, 5210.558, 5212.122, 5213.859, 5206.857,
  5053.278, 5058.651, 5065.979, 5078.542, 5092.965, 5113.979, 5123.055, 
    5147.269, 5156.384, 5166.896, 5174.659, 5179.793, 5179.627, 5176.29, 
    5171.166,
  5052.842, 5056.048, 5062.509, 5069.528, 5082.419, 5090.925, 5111.885, 
    5111.826, 5131.306, 5141.206, 5145.966, 5148.205, 5147.359, 5143.761, 
    5134.639,
  5053.485, 5053.091, 5057.744, 5063.368, 5071.638, 5082.919, 5088.894, 
    5103.596, 5109.774, 5109.048, 5118.453, 5116.464, 5116.409, 5108.838, 
    5103.348,
  5056.188, 5051.971, 5050.701, 5053.877, 5058.564, 5064.701, 5074.101, 
    5075.453, 5082.251, 5091.481, 5091.598, 5090.96, 5088.904, 5081.874, 
    5073.396,
  5061.827, 5055.771, 5051.078, 5048.688, 5051.678, 5055.906, 5060.229, 
    5067.632, 5070.948, 5069.264, 5070.183, 5068.305, 5062.965, 5054.808, 
    5043.839,
  5066.896, 5060.329, 5054.549, 5052.292, 5049.52, 5049.688, 5051.016, 
    5050.642, 5051.289, 5053.364, 5050.801, 5045.575, 5038.308, 5028.071, 
    5015.418,
  5065.928, 5058.871, 5052.36, 5047.71, 5044.843, 5043.465, 5041.646, 
    5041.314, 5038.166, 5032.479, 5027.105, 5020.213, 5010.197, 4998.611, 
    4984.798,
  5061.404, 5051.074, 5042.262, 5036.619, 5031.259, 5027.274, 5023.356, 
    5017.818, 5012.812, 5007.985, 5000.621, 4990.888, 4979.342, 4966.988, 
    4953.005,
  5061.824, 5049.009, 5039.227, 5034.908, 5031.499, 5029.071, 5029.516, 
    5038.226, 5051.409, 5068.461, 5091.699, 5122.748, 5157.716, 5189.366, 
    5217.708,
  5061.49, 5050.657, 5042.122, 5040.246, 5040.291, 5039.406, 5043.341, 
    5050.098, 5063.867, 5086.187, 5112.036, 5145.046, 5175.969, 5206.084, 
    5231.269,
  5061.16, 5051.625, 5045.234, 5045.228, 5047.994, 5052.059, 5055.033, 
    5068.76, 5085.511, 5104.863, 5132.993, 5162.825, 5190.971, 5214.861, 
    5238.443,
  5059.913, 5050.759, 5048.36, 5047.028, 5054.971, 5057.713, 5070.633, 
    5077.617, 5097.132, 5119.778, 5148.419, 5174.762, 5199.656, 5222.926, 
    5241.426,
  5058.949, 5048.824, 5047.481, 5048.312, 5055.369, 5066.84, 5075.633, 
    5091.418, 5114.362, 5131.054, 5157.053, 5179.421, 5202.453, 5219.954, 
    5236.099,
  5058.879, 5048.755, 5043.351, 5045.862, 5052.892, 5063.225, 5079.824, 
    5094.368, 5108.862, 5134.636, 5154.852, 5177.182, 5196.79, 5213.531, 
    5226.51,
  5055.736, 5048.459, 5042.379, 5040.848, 5046.116, 5057.312, 5070.758, 
    5089.563, 5110.585, 5127.437, 5147.918, 5167.18, 5183.797, 5197.626, 
    5207.971,
  5051.571, 5045.696, 5039.841, 5037.758, 5038.652, 5045.298, 5058.754, 
    5072.897, 5089.864, 5111.707, 5131.654, 5148.923, 5165.527, 5178.257, 
    5187.82,
  5039.703, 5034.625, 5030.537, 5028.564, 5027.679, 5032.603, 5041.35, 
    5057.084, 5074.262, 5091.034, 5107.984, 5126.141, 5141.598, 5154.242, 
    5163.354,
  5025.468, 5019.47, 5014.313, 5013.107, 5013.568, 5016.1, 5022.251, 
    5033.424, 5047.9, 5066.029, 5084.123, 5101.133, 5116.369, 5129.458, 
    5138.821,
  5106.018, 5095.672, 5084.41, 5072.747, 5060.401, 5046.901, 5029.889, 
    5018.1, 5009.977, 5006.869, 5011.451, 5023.024, 5040.246, 5058.782, 
    5077.641,
  5094.265, 5083.924, 5072.589, 5061.95, 5050.234, 5034.628, 5020.307, 
    5005.615, 4999.447, 5002.936, 5012.787, 5030.624, 5050.342, 5071.931, 
    5092.319,
  5084.5, 5075.249, 5065.26, 5056.539, 5043.77, 5031.953, 5009.729, 5004.521, 
    5001.924, 5008.464, 5023.344, 5044.408, 5066.196, 5087.894, 5115.283,
  5075.817, 5067.337, 5058.888, 5049.907, 5041.177, 5024.665, 5013.808, 
    4999.987, 5004.157, 5018.755, 5041.078, 5063.256, 5087.746, 5116.567, 
    5146.366,
  5066.528, 5060.062, 5054.047, 5047.026, 5041.024, 5027.688, 5014.838, 
    5007.591, 5024.565, 5035.412, 5062.129, 5085.105, 5115.524, 5143.895, 
    5171.815,
  5055.465, 5051.112, 5047.387, 5042.813, 5038.074, 5030.572, 5020.811, 
    5021.43, 5029.161, 5057.717, 5082.709, 5110.551, 5141.758, 5170.594, 
    5193.587,
  5042.685, 5041.193, 5040.008, 5039.227, 5037.796, 5035.022, 5027.665, 
    5033.283, 5054.363, 5078.184, 5104.535, 5134.413, 5164.029, 5189.298, 
    5209.659,
  5027.379, 5026.616, 5028.573, 5032.006, 5032.515, 5034.402, 5036.042, 
    5042.549, 5063.796, 5092.934, 5122.393, 5151.916, 5181.074, 5204.067, 
    5221.939,
  5009.606, 5007.442, 5012.382, 5022.038, 5029.307, 5033.991, 5038.155, 
    5051.977, 5079.538, 5106.833, 5135.067, 5165.291, 5191.669, 5212.625, 
    5228.149,
  4987.762, 4981.145, 4987.166, 5000.068, 5013.198, 5025.295, 5036.531, 
    5051.763, 5079.116, 5110.347, 5141.061, 5171.36, 5196.999, 5217.342, 
    5230.257,
  5097.769, 5083.916, 5074.954, 5072.387, 5071.059, 5069.216, 5067.02, 
    5066.809, 5065.781, 5064.901, 5066.174, 5071.089, 5078.797, 5088.789, 
    5099.886,
  5089.184, 5071.64, 5061.695, 5059.188, 5058.962, 5059.113, 5057.879, 
    5054.269, 5050.983, 5049.481, 5050.635, 5057.207, 5067.763, 5081.398, 
    5093.263,
  5081.439, 5058.674, 5048.444, 5046.751, 5048.818, 5051.438, 5046.383, 
    5044.379, 5038.723, 5036.369, 5039.823, 5050.033, 5064.066, 5078.515, 
    5094.625,
  5071.823, 5045.927, 5033.678, 5031.387, 5037.704, 5038.915, 5042.295, 
    5032.773, 5031.359, 5029.964, 5039.237, 5051.421, 5069.04, 5089.259, 
    5106.641,
  5062.818, 5031.624, 5017.888, 5018.208, 5027.834, 5034.365, 5032.182, 
    5032.333, 5029.683, 5033.585, 5045.957, 5063.116, 5086.786, 5105.887, 
    5119.461,
  5054.935, 5018.525, 5001.881, 5005.126, 5017.262, 5027.512, 5029.334, 
    5029.936, 5032.27, 5044.041, 5060.484, 5084.754, 5107.316, 5122.87, 
    5129.806,
  5047.731, 5008.4, 4990.483, 4997.387, 5013.272, 5024.616, 5026.784, 
    5032.664, 5042.173, 5058.733, 5081.834, 5106.826, 5125.958, 5136.651, 
    5138.499,
  5043.014, 5001.252, 4982.637, 4992.699, 5009.257, 5022.148, 5027.354, 
    5036.629, 5052.632, 5076.816, 5103.69, 5128.198, 5143.7, 5150.511, 
    5147.788,
  5041.034, 4997.054, 4980.158, 4993.588, 5011.798, 5023.633, 5030.462, 
    5046.501, 5068.872, 5096.796, 5124.961, 5147.503, 5159.931, 5164.473, 
    5159.152,
  5041.976, 4995.66, 4979.42, 4993.293, 5011.966, 5025.446, 5036.307, 
    5056.855, 5083.553, 5115.083, 5143.716, 5164.923, 5176.766, 5179.122, 
    5173.519,
  5104.166, 5062.714, 5033.79, 5022.152, 5024.423, 5032.058, 5034.106, 
    5037.114, 5038.078, 5038.003, 5038.354, 5039.276, 5041.406, 5045.388, 
    5053.957,
  5109.419, 5068.773, 5040.826, 5029.643, 5032.335, 5035.19, 5038.019, 
    5036.225, 5036.002, 5036.912, 5037.609, 5039.234, 5041.973, 5046.323, 
    5052.001,
  5118.586, 5079.173, 5052.56, 5041.579, 5040.266, 5045.76, 5040.312, 
    5039.075, 5036.684, 5035.623, 5036.87, 5039.711, 5043.039, 5047.284, 
    5053.164,
  5129.186, 5092.563, 5068.099, 5053.617, 5053.654, 5048.892, 5048.637, 
    5039.897, 5034.791, 5033.569, 5035.344, 5037.807, 5042.683, 5047.341, 
    5053.811,
  5143.292, 5108.242, 5086.519, 5071.13, 5067.224, 5062.686, 5053.997, 
    5045.417, 5039.005, 5034.567, 5037.125, 5040.311, 5047.06, 5051.217, 
    5057.704,
  5160.547, 5123.891, 5104.237, 5090.337, 5082.762, 5074.498, 5066.369, 
    5056.02, 5049.658, 5048.342, 5049.837, 5052.6, 5056.171, 5059.375, 
    5062.046,
  5179.126, 5140.481, 5122.878, 5109.522, 5100.321, 5091.321, 5079.866, 
    5072.054, 5067.015, 5063.725, 5062.342, 5063.046, 5063.729, 5066.519, 
    5069.551,
  5200.032, 5158.16, 5137.854, 5126.781, 5115.528, 5106.773, 5097.093, 
    5088.323, 5079.674, 5074.987, 5072.031, 5071.526, 5072.499, 5075.976, 
    5081.536,
  5220.092, 5178.618, 5153.997, 5141.757, 5131.946, 5124.434, 5115.271, 
    5107.626, 5098.543, 5090.917, 5085.106, 5084.293, 5087.097, 5093.424, 
    5101.302,
  5238.085, 5196.833, 5167.914, 5153.802, 5144.08, 5138.917, 5133.722, 
    5126.513, 5116.116, 5109.011, 5104.494, 5104.872, 5108.47, 5115.217, 
    5122.271,
  5272.583, 5238.435, 5203.131, 5166.612, 5134.628, 5111.873, 5094.193, 
    5085.696, 5079.112, 5070.026, 5062.96, 5055.397, 5049.953, 5044.99, 
    5044.802,
  5288.412, 5255.5, 5220.438, 5183.454, 5149.308, 5117.156, 5104.603, 
    5089.401, 5080.996, 5075.129, 5067.371, 5060.609, 5054.062, 5047.809, 
    5044.109,
  5304.924, 5273.691, 5239.087, 5204.547, 5164.261, 5139.943, 5107.375, 
    5101.013, 5089.455, 5082.234, 5073.51, 5066.702, 5059.117, 5054.32, 
    5049.294,
  5319.131, 5288.749, 5257.388, 5221.117, 5186.357, 5147.051, 5127.31, 
    5106.385, 5095.624, 5089.023, 5081.572, 5073.711, 5066.836, 5060.673, 
    5055.733,
  5333.388, 5303.133, 5274.186, 5239.036, 5205.525, 5169.429, 5138.181, 
    5120.129, 5110.528, 5098.379, 5092.481, 5083.545, 5077.726, 5068.999, 
    5063.788,
  5345.072, 5315.392, 5286.234, 5254.353, 5220.84, 5186.26, 5154.684, 
    5130.847, 5116.608, 5109.56, 5102.938, 5095.606, 5089.244, 5081.473, 
    5074.358,
  5354.065, 5327.549, 5298.786, 5267.711, 5236.133, 5203.797, 5171.704, 
    5145.438, 5131.278, 5121.017, 5114.088, 5108.417, 5101.539, 5093.842, 
    5085.22,
  5359.806, 5335.983, 5307.314, 5277.503, 5245.515, 5214.59, 5185.375, 
    5158.532, 5139.6, 5130.388, 5124.072, 5118.506, 5112.317, 5104.272, 
    5093.704,
  5362.716, 5342.052, 5315.307, 5284.619, 5253.594, 5223.235, 5194.856, 
    5170.104, 5151.496, 5139.961, 5132.434, 5126.903, 5120.165, 5111.245, 
    5099.395,
  5364.069, 5341.626, 5314.793, 5285.719, 5253.037, 5222.488, 5197.158, 
    5174.158, 5155.256, 5144.089, 5137.145, 5131.206, 5124.228, 5114.642, 
    5101.046,
  5409.601, 5384.834, 5354.381, 5322.114, 5290.472, 5259.274, 5225.589, 
    5201.287, 5175.863, 5147.022, 5125.797, 5107.054, 5092.953, 5080.219, 
    5073.162,
  5410.117, 5384.368, 5354.493, 5322.779, 5290.304, 5253.674, 5227.46, 
    5186.274, 5161.4, 5141.836, 5119.873, 5103.19, 5089.423, 5078.615, 
    5069.913,
  5409.302, 5383.102, 5352.979, 5321.835, 5284.712, 5256.106, 5209.561, 
    5190.404, 5152.117, 5127.068, 5110.168, 5097.046, 5085.034, 5075.635, 
    5067.123,
  5406.614, 5378.407, 5348.561, 5313.021, 5275.65, 5231.878, 5200.657, 
    5151.52, 5129.131, 5106.47, 5093.186, 5085.045, 5080.109, 5073.034, 
    5066.05,
  5403.285, 5374.588, 5342.802, 5304.007, 5262.136, 5216.207, 5167.702, 
    5137.46, 5103.021, 5080.323, 5073.448, 5069.24, 5071.269, 5068.474, 
    5065.042,
  5398.494, 5367.713, 5331.005, 5288.913, 5240.099, 5187.809, 5140.154, 
    5094.252, 5064.681, 5051.121, 5044.037, 5049.579, 5057.298, 5061.866, 
    5062.343,
  5393.086, 5361.363, 5320.88, 5273.434, 5217.911, 5160.677, 5107.212, 
    5066.058, 5036.109, 5019.187, 5019.267, 5029.064, 5040.833, 5051.191, 
    5054.879,
  5387.631, 5351.443, 5305.632, 5252.219, 5188.816, 5126.894, 5071.511, 
    5025.487, 4998.223, 4989.812, 4994.52, 5008.644, 5025.87, 5039.241, 
    5045.665,
  5382.403, 5345.412, 5296.921, 5236.681, 5168.875, 5100.475, 5040.916, 
    4999.472, 4974.357, 4965.645, 4975.62, 4994.295, 5012.895, 5026.991, 
    5033.912,
  5377.979, 5334.979, 5279.88, 5214.803, 5139.501, 5070.24, 5015.231, 
    4973.682, 4951.655, 4950.904, 4965.1, 4985.045, 5003.19, 5016.219, 
    5021.487,
  5346.058, 5295.255, 5243.748, 5192.291, 5145.1, 5098.292, 5046.657, 
    5011.37, 4983.521, 4957.521, 4948.878, 4951.78, 4963.781, 4981.077, 
    5003.088,
  5348.996, 5296.648, 5240.183, 5185.396, 5134.771, 5076.273, 5035.226, 
    4975.2, 4942.365, 4926.328, 4916.952, 4920.889, 4932.8, 4956.763, 4979.138,
  5355.167, 5302.137, 5241.625, 5185.601, 5125.519, 5081.961, 5009.867, 
    4979.775, 4933.995, 4907.019, 4894.612, 4898.893, 4912.118, 4935.409, 
    4963.32,
  5362.916, 5307.974, 5246.944, 5184.256, 5129.608, 5066.78, 5026.263, 
    4961.57, 4922.312, 4900.114, 4887.33, 4888.407, 4903.951, 4928.875, 
    4956.749,
  5371.941, 5317.738, 5256.543, 5192.727, 5137.668, 5082.916, 5026.682, 
    4978.184, 4941.226, 4904.081, 4893.697, 4891.532, 4908.819, 4931.2, 
    4959.849,
  5380.666, 5327.923, 5266.265, 5204.911, 5148.315, 5097.819, 5047.339, 
    4992.838, 4948.334, 4922.756, 4908.716, 4908.676, 4924.783, 4947.438, 
    4969.517,
  5390.568, 5341.65, 5283.052, 5222.195, 5169.169, 5120.999, 5068.993, 
    5023.208, 4982.418, 4949.543, 4933.88, 4934.561, 4946.861, 4965.487, 
    4980.503,
  5400.542, 5353.853, 5298.46, 5240.278, 5186.218, 5141.639, 5096.072, 
    5049.276, 5008.773, 4980.917, 4965.384, 4963.398, 4972.117, 4983.93, 
    4991.948,
  5409.808, 5367.601, 5317.428, 5261.288, 5210.1, 5166.16, 5122.299, 
    5082.387, 5046.95, 5016.253, 4998.181, 4992.763, 4994.47, 4998.339, 
    5000.099,
  5417.346, 5376.428, 5329.922, 5278.584, 5225.724, 5183.916, 5145.449, 
    5106.036, 5072.292, 5045.5, 5026.466, 5016.207, 5010.872, 5006.836, 
    5001.066,
  5417.716, 5384.351, 5350.047, 5311.114, 5272.017, 5231.913, 5187.29, 
    5150.679, 5111.872, 5070.562, 5039.029, 5014, 4998.613, 4990.369, 4991.618,
  5418.924, 5387.547, 5355.4, 5320.27, 5284.99, 5242.818, 5211.121, 5163.681, 
    5125.612, 5092.36, 5059.732, 5032.624, 5010.532, 4998.622, 4992.176,
  5417.679, 5388.421, 5357.437, 5327.329, 5290.253, 5263.296, 5212.939, 
    5188.47, 5151.223, 5114.639, 5080.157, 5051.982, 5027.126, 5010.23, 
    4998.976,
  5410.849, 5382.968, 5355.231, 5324.975, 5295.816, 5259.349, 5235.005, 
    5193.292, 5160.112, 5130.322, 5098.536, 5069.63, 5043.794, 5023.87, 
    5009.873,
  5401.409, 5375.23, 5349.93, 5321.81, 5295.254, 5266.202, 5233.028, 
    5207.503, 5177.385, 5139.716, 5112.055, 5082.168, 5058.172, 5035.515, 
    5020.353,
  5387.423, 5362.811, 5337.823, 5313.543, 5287.423, 5261.235, 5235.97, 
    5202.977, 5172.181, 5146.558, 5118.46, 5090.856, 5065.684, 5043.657, 
    5026.565,
  5370.809, 5348.491, 5324.534, 5302.014, 5279.122, 5255.615, 5229.43, 
    5205.767, 5178.517, 5148.224, 5119.9, 5093.531, 5067.287, 5045.348, 
    5026.709,
  5351.991, 5329.387, 5306.145, 5286.097, 5263.605, 5243.265, 5220.91, 
    5195.368, 5168.858, 5144.948, 5117.984, 5090.619, 5064.149, 5041.536, 
    5022.294,
  5332.151, 5310.146, 5288.787, 5268.769, 5249.292, 5230.03, 5209.214, 
    5188.986, 5165.28, 5138.889, 5110.978, 5083.545, 5056.396, 5033.705, 
    5013.423,
  5312.89, 5288.197, 5267.493, 5249.511, 5230.867, 5213.622, 5195.863, 
    5174.612, 5152.378, 5129.412, 5102.422, 5073.313, 5046.21, 5023.033, 
    5002.068,
  5323.524, 5290.958, 5262.263, 5237.886, 5220.254, 5205.839, 5192.206, 
    5184.491, 5177.089, 5166.431, 5158.817, 5150.649, 5141.177, 5129.247, 
    5118.006,
  5320.211, 5285.875, 5255.628, 5229.254, 5208.902, 5190.29, 5182.103, 
    5166.773, 5159.652, 5155.484, 5147.96, 5141.051, 5132.36, 5123.278, 
    5110.887,
  5320.779, 5285.319, 5253.834, 5227.085, 5202.11, 5188.459, 5164.42, 
    5162.082, 5148.158, 5140.829, 5134.613, 5129.569, 5121.382, 5111.963, 
    5101.361,
  5323.241, 5287.051, 5254.747, 5224.79, 5200.636, 5174.911, 5163.566, 
    5140.381, 5135.184, 5128.972, 5121.347, 5116.094, 5109.626, 5101.901, 
    5089.591,
  5327.715, 5291.607, 5259.094, 5228.422, 5201.632, 5177.197, 5152.816, 
    5139.944, 5124.414, 5113.166, 5108.71, 5101.681, 5096.996, 5087.743, 
    5078.429,
  5332.116, 5295.949, 5262.545, 5232.282, 5202.486, 5175.854, 5152.646, 
    5129.269, 5113.223, 5103.817, 5095.027, 5089.109, 5083.782, 5075.454, 
    5064.353,
  5336.12, 5302.283, 5269.025, 5238.84, 5209.229, 5180.625, 5152.965, 
    5131.336, 5110.158, 5093.277, 5083.477, 5076.775, 5069.561, 5060.77, 
    5048.426,
  5340.212, 5306.781, 5273.436, 5243.896, 5212.502, 5184.396, 5156.388, 
    5129.479, 5105.41, 5088.012, 5073.47, 5063.989, 5056.108, 5045.61, 
    5032.147,
  5344.177, 5312.643, 5280.691, 5251.112, 5221.412, 5191.991, 5161.823, 
    5134.929, 5107.84, 5084.935, 5065.987, 5052.603, 5039.665, 5028.218, 
    5015.916,
  5346.515, 5314.386, 5283.706, 5255.117, 5224.403, 5195.775, 5166.814, 
    5136.718, 5108.684, 5083.951, 5061.383, 5042.277, 5028.285, 5016.791, 
    5008.154,
  5347.691, 5319.251, 5293.052, 5268.705, 5247.098, 5226.345, 5203.96, 
    5186.632, 5167.684, 5148.247, 5135.462, 5128.772, 5129.159, 5132.512, 
    5137.528,
  5347.757, 5317.707, 5291.268, 5266.395, 5246.115, 5222.797, 5207.618, 
    5181.719, 5161.685, 5144.878, 5128.748, 5118.591, 5116.179, 5120.143, 
    5124.623,
  5347.149, 5316.474, 5289.211, 5265.785, 5242.888, 5228.163, 5201.922, 
    5188.51, 5165.642, 5142.965, 5123.988, 5110.862, 5104.343, 5106.541, 
    5112.451,
  5345.059, 5312.917, 5285.214, 5260.359, 5239.669, 5218.342, 5206.495, 
    5182.271, 5161.38, 5143.113, 5121.7, 5105.98, 5097.107, 5096.127, 5099.531,
  5342.505, 5309.36, 5281.497, 5256.672, 5236.187, 5217.653, 5199.757, 
    5186.216, 5168.112, 5141.448, 5121.961, 5102.49, 5092.422, 5086.775, 
    5090.106,
  5338.309, 5303.484, 5274.166, 5250.539, 5229.118, 5210.939, 5197.295, 
    5179.756, 5162.081, 5143.777, 5122.153, 5102.678, 5089.834, 5082.331, 
    5081.446,
  5332.133, 5298.009, 5268.027, 5244.643, 5224.073, 5207.145, 5191.44, 
    5180.327, 5164.927, 5144.604, 5123.043, 5103.382, 5087.35, 5077.932, 
    5072.857,
  5324.346, 5289.042, 5258.165, 5235.767, 5215.167, 5199.554, 5185.697, 
    5172.012, 5157.26, 5142.729, 5123.712, 5104.037, 5086.703, 5073.96, 
    5065.193,
  5315.161, 5281.084, 5251.404, 5228.305, 5208.801, 5193.483, 5179.366, 
    5168.424, 5154.245, 5137.954, 5120.722, 5102.763, 5085.326, 5070.638, 
    5058.09,
  5305.031, 5269.49, 5240.029, 5219.088, 5199.779, 5184.379, 5170.988, 
    5156.867, 5142.585, 5129.042, 5113.889, 5098.339, 5081.702, 5067.141, 
    5054.572,
  5307.778, 5269.66, 5240.018, 5219.187, 5204.417, 5189.23, 5174.527, 
    5168.746, 5166.813, 5160.299, 5151.858, 5137.5, 5123.04, 5110.836, 
    5107.983,
  5313.324, 5271.022, 5240.906, 5217.633, 5203.723, 5185.231, 5175.259, 
    5163.299, 5161.655, 5156.939, 5149.02, 5136.623, 5122.533, 5110.136, 
    5103.592,
  5318.486, 5272.891, 5242.452, 5218.625, 5203.159, 5189.93, 5171.738, 
    5166.004, 5160.65, 5154.506, 5146.347, 5135.381, 5122.598, 5109.464, 
    5101.237,
  5322.819, 5273.691, 5242.178, 5216.773, 5202.822, 5185.301, 5175.372, 
    5161.456, 5156.117, 5150.204, 5142.57, 5132.734, 5122.003, 5110.302, 
    5100.479,
  5325.919, 5274.518, 5242.87, 5216.622, 5202.07, 5187.586, 5173.579, 
    5163.223, 5155.176, 5146.554, 5138.584, 5128.052, 5119.031, 5108.599, 
    5100.443,
  5326.182, 5273.042, 5240.022, 5214.229, 5198.313, 5183.608, 5172.879, 
    5159.478, 5150.22, 5140.973, 5132.11, 5121.874, 5113.138, 5104.158, 
    5097.115,
  5323.425, 5273.082, 5239.083, 5213.418, 5196.314, 5181.696, 5169.162, 
    5157.52, 5146.278, 5134.434, 5123.781, 5113.189, 5103.649, 5095.691, 
    5089.545,
  5319.577, 5269.941, 5234.702, 5209.64, 5190.709, 5175.696, 5163.26, 
    5150.024, 5137.006, 5124.736, 5112.294, 5101.264, 5091.546, 5084.189, 
    5078.63,
  5315.706, 5267.988, 5234.304, 5207.982, 5188.124, 5171.646, 5156.951, 
    5142.761, 5127.884, 5112.747, 5098.724, 5086.419, 5076.007, 5069.213, 
    5064.471,
  5310.582, 5262.147, 5228.536, 5203.438, 5181.867, 5163.378, 5147.936, 
    5131.049, 5114.593, 5097.962, 5082.4, 5068.733, 5057.936, 5051.244, 
    5047.574,
  5336.96, 5293.757, 5256.798, 5226.369, 5202, 5182.56, 5164.37, 5153.049, 
    5144.915, 5136.152, 5131.636, 5125.979, 5120.909, 5113.726, 5106.691,
  5337.541, 5292.789, 5255.078, 5223.566, 5199.4, 5175.517, 5163.983, 
    5144.909, 5136.878, 5130.493, 5124.041, 5118.714, 5113.915, 5110.231, 
    5104.955,
  5335.867, 5290.922, 5252.775, 5221.983, 5196.178, 5178.462, 5153.085, 
    5145.358, 5130.56, 5120.876, 5114.761, 5109.921, 5105.522, 5102.44, 
    5100.016,
  5330.586, 5286.118, 5248.472, 5216.288, 5190.824, 5164.44, 5151.473, 
    5126.193, 5117.354, 5109.372, 5101.946, 5097.441, 5094.626, 5092.89, 
    5092.376,
  5324.37, 5281.053, 5244.833, 5212.242, 5186.263, 5160.877, 5134.82, 
    5122.173, 5104.559, 5090.063, 5085.984, 5080.631, 5080.188, 5079.029, 
    5081.246,
  5315.897, 5273.896, 5237.734, 5205.826, 5176.129, 5147.668, 5124.218, 
    5096.732, 5080.326, 5071.224, 5062.685, 5059.885, 5060.369, 5062.597, 
    5065.991,
  5305.962, 5268.181, 5231.918, 5200.172, 5169.042, 5138.007, 5106.83, 
    5084.539, 5062.867, 5045.475, 5037.058, 5035.072, 5036.708, 5041.773, 
    5047.82,
  5296.243, 5260.55, 5223.987, 5191.671, 5156.285, 5122.608, 5089.923, 
    5058.49, 5032.781, 5017.063, 5006.793, 5005.146, 5008.857, 5017.75, 
    5026.95,
  5287.379, 5254.188, 5219.252, 5185.028, 5148.354, 5110.421, 5071.477, 
    5038.64, 5008.849, 4984.983, 4972.615, 4971.309, 4977.291, 4989.509, 
    5003.872,
  5280.087, 5246.576, 5211.701, 5175.89, 5134.608, 5093.316, 5052.301, 
    5012.033, 4977.144, 4949.859, 4935.338, 4933.289, 4942.138, 4957.705, 
    4977.603,
  5202.927, 5172.902, 5148.093, 5125.718, 5106.002, 5086.863, 5067.766, 
    5055.583, 5045.229, 5036.445, 5035.917, 5039.318, 5044.461, 5050.906, 
    5058.783,
  5199.43, 5167.589, 5141.252, 5115.884, 5093.721, 5069.117, 5055.844, 
    5033.97, 5023.114, 5018.856, 5015.918, 5019.65, 5026.76, 5037.024, 5045.65,
  5197.337, 5164.175, 5135.647, 5108.369, 5081.445, 5063.833, 5033.725, 
    5025.827, 5007.774, 4996.934, 4993.685, 4997.042, 5005.759, 5017.705, 
    5030.826,
  5193.908, 5158.239, 5127.659, 5096.083, 5069.175, 5040.213, 5026.844, 
    4996.127, 4985.3, 4976.105, 4969.247, 4970.949, 4981.278, 4998.142, 
    5014.779,
  5190.73, 5152.954, 5120.029, 5086.179, 5057.736, 5032.326, 5003.947, 
    4989.667, 4968.361, 4948.329, 4943, 4941.4, 4953.856, 4973.039, 4997.186,
  5186.472, 5144.941, 5108.46, 5074.484, 5043.72, 5016.14, 4993.014, 
    4963.271, 4941.514, 4926.708, 4913.266, 4911.727, 4923.114, 4947.816, 
    4977.402,
  5181.467, 5138.36, 5099.837, 5064.92, 5034.607, 5005.943, 4976.865, 
    4952.982, 4927.162, 4901.743, 4885.778, 4882.82, 4893.027, 4921.828, 
    4957.126,
  5176.062, 5129.571, 5088.729, 5052.987, 5021.127, 4992.244, 4963.111, 
    4931.183, 4901.75, 4878.359, 4858.022, 4852.584, 4864.289, 4896.674, 
    4939.853,
  5170.865, 5123.688, 5082.616, 5045.849, 5014.852, 4983.271, 4949.374, 
    4918.569, 4886.52, 4856.056, 4833.019, 4826.607, 4839.456, 4875.42, 
    4926.011,
  5166.289, 5114.786, 5072.674, 5036.839, 5004.239, 4971.406, 4937.068, 
    4900.193, 4866.146, 4836.368, 4813.378, 4805.776, 4819.846, 4861.353, 
    4915.841,
  5129.912, 5081.58, 5046.263, 5017.958, 4999.131, 4984.742, 4974.133, 
    4970.429, 4969.601, 4974.578, 4986.448, 5002.956, 5022.52, 5039.679, 
    5056.934,
  5110.282, 5061.994, 5029.177, 5001.833, 4983.5, 4967.636, 4962.08, 4953.15, 
    4954.979, 4960.926, 4971.53, 4987.814, 5007.175, 5030.132, 5048.314,
  5092.129, 5045.856, 5014.509, 4987.619, 4968.841, 4958.701, 4944.557, 
    4945.875, 4942.053, 4947.614, 4958.953, 4973.431, 4993.651, 5014.766, 
    5037.553,
  5073.209, 5029.597, 4997.818, 4970.533, 4953.336, 4938.37, 4937.766, 
    4926.616, 4932.506, 4935.452, 4946.51, 4960.923, 4979.824, 5003.964, 
    5028.368,
  5056.658, 5013.899, 4981.034, 4953.635, 4936.184, 4926.586, 4918.268, 
    4919.729, 4918.176, 4923.805, 4934.386, 4948.302, 4967.494, 4989.475, 
    5017.201,
  5040.956, 4996.917, 4960.125, 4932.739, 4913.864, 4904.856, 4903.183, 
    4900.316, 4904.219, 4911.896, 4920.644, 4936.156, 4954.668, 4978.533, 
    5006.235,
  5027.541, 4983.868, 4943.199, 4913.804, 4893.084, 4884.235, 4880.632, 
    4884.961, 4888.866, 4896.192, 4908.06, 4923.653, 4942.77, 4966.669, 
    4995.342,
  5019.359, 4972.502, 4927.243, 4894.616, 4869.401, 4858.693, 4857.272, 
    4861.332, 4869.268, 4881.471, 4894.25, 4911.294, 4932.097, 4957.25, 
    4988.12,
  5017.054, 4968.937, 4920.173, 4882.457, 4853.884, 4838.897, 4835.284, 
    4843.292, 4853.415, 4866.009, 4881.769, 4900.77, 4922.996, 4949.713, 
    4982.377,
  5021.017, 4968.335, 4916.034, 4876.138, 4842.033, 4824.097, 4819.845, 
    4826.508, 4839.59, 4855.567, 4873.048, 4893.366, 4917.388, 4946.759, 
    4982.876,
  5032.557, 4993.119, 4960.844, 4937.852, 4925.505, 4923.08, 4928.734, 
    4940.915, 4952.162, 4960.052, 4970.882, 4990.277, 5017.595, 5049.138, 
    5078.564,
  5006.956, 4962.175, 4928.576, 4903.645, 4895.022, 4897.754, 4911.79, 
    4923.292, 4936.193, 4948.713, 4961.648, 4983.733, 5013.061, 5048.712, 
    5076.984,
  4986.545, 4937.644, 4902.021, 4876.931, 4874.672, 4884.337, 4895.805, 
    4917.97, 4931.116, 4941.726, 4955.375, 4978.978, 5012.095, 5045.42, 
    5075.178,
  4968.704, 4917.179, 4879.131, 4853.846, 4853.856, 4863.371, 4891.594, 
    4905.548, 4923.703, 4936.208, 4951.92, 4977.703, 5013.774, 5049.056, 
    5077.544,
  4958.499, 4905.621, 4865.169, 4838.864, 4837.518, 4855.117, 4879.485, 
    4910.126, 4925.081, 4934.735, 4951.125, 4980.276, 5017.679, 5050.094, 
    5079.612,
  4957.289, 4903.104, 4861.69, 4834.849, 4831.314, 4846.805, 4884.112, 
    4905.67, 4921.381, 4936.261, 4954.336, 4986.543, 5023.235, 5056.105, 
    5084.138,
  4964.77, 4913.489, 4873.495, 4847.576, 4841.441, 4858.72, 4887.079, 
    4914.935, 4928.512, 4940.847, 4961.622, 4994.707, 5029.835, 5060.774, 
    5088.789,
  4981.802, 4931.583, 4893.498, 4870.69, 4863.322, 4878.312, 4901.406, 
    4916.295, 4929.793, 4948.062, 4971.498, 5004.281, 5037.623, 5068.531, 
    5095.921,
  5003.653, 4955.216, 4919.349, 4896.896, 4890.837, 4898.58, 4913.103, 
    4929.057, 4943.163, 4959.348, 4983.307, 5014.81, 5045.428, 5075.634, 
    5102.461,
  5032.119, 4981.296, 4944.955, 4924.303, 4914.127, 4917.997, 4928.17, 
    4938.098, 4951.797, 4971.124, 4996.173, 5025.626, 5054.931, 5084.299, 
    5110.851,
  5039.333, 4992.756, 4951.955, 4919.501, 4892.571, 4869.741, 4855.527, 
    4867.909, 4907.269, 4947.762, 4980.851, 5010.924, 5034.936, 5057.592, 
    5082.934,
  5032.187, 4987.288, 4949.385, 4920.095, 4896.537, 4870.911, 4861.036, 
    4871.649, 4910.608, 4951.53, 4982.82, 5009.11, 5029.899, 5053.544, 
    5078.488,
  5031.163, 4989.551, 4955.218, 4931.156, 4908.859, 4896.232, 4881.2, 
    4893.02, 4930.052, 4960.751, 4986.383, 5007.271, 5027.347, 5047.739, 
    5075.448,
  5033.281, 4994.456, 4964.431, 4941.436, 4928.507, 4910.196, 4912.937, 
    4918.703, 4944.434, 4969.019, 4990.903, 5006.427, 5026.32, 5049.201, 
    5078.46,
  5038.856, 5003.524, 4976.579, 4956.384, 4945.322, 4938.574, 4936.069, 
    4942.8, 4965.297, 4975.89, 4993.928, 5007.197, 5028.811, 5051.982, 
    5083.729,
  5046.033, 5013.057, 4988.063, 4970.455, 4959.613, 4952.801, 4954.47, 
    4960.437, 4966.897, 4983.839, 4996.048, 5012.848, 5035.414, 5062.99, 
    5093.405,
  5054.112, 5024.065, 5001.227, 4984.109, 4973.001, 4968.247, 4965.178, 
    4970.694, 4980.614, 4990.288, 5002.9, 5023.607, 5047.483, 5075.887, 
    5106.616,
  5063.396, 5033.52, 5010.836, 4995.279, 4982.274, 4975.296, 4974.391, 
    4977.073, 4983.744, 4998.71, 5016.912, 5040.023, 5065.296, 5093.841, 
    5124.308,
  5073.927, 5044.733, 5021.91, 5006.011, 4995.237, 4989.144, 4986.396, 
    4992.315, 5003.772, 5018.375, 5038.003, 5061.27, 5085.089, 5113.271, 
    5141.548,
  5087.569, 5055.76, 5032.059, 5017.645, 5007.005, 5002.94, 5004.639, 
    5010.846, 5022.666, 5041.056, 5061.808, 5083.584, 5106.86, 5132.647, 
    5159.285,
  5106.44, 5080.213, 5057.04, 5037.677, 5019.111, 5000.201, 4977.594, 
    4963.324, 4952.836, 4955.694, 4965.642, 4976.135, 4991.439, 5004.748, 
    5022.677,
  5097.475, 5073.111, 5053.274, 5039.106, 5027.562, 5012.54, 5004.883, 
    4994.104, 4988.175, 4994.422, 5002.874, 5015.41, 5024.82, 5038.811, 
    5053.903,
  5093.806, 5070.77, 5054.699, 5046.132, 5036.524, 5038.007, 5025.872, 
    5026.414, 5029.082, 5031.677, 5037.612, 5046.035, 5057.296, 5067.501, 
    5079.277,
  5093.34, 5070.455, 5057.888, 5048.834, 5050.074, 5042.417, 5052.695, 
    5050.274, 5051.321, 5057.945, 5066.061, 5071.827, 5079.986, 5088.75, 
    5100.056,
  5096.427, 5075.035, 5062.807, 5056.52, 5058.78, 5062.982, 5065.932, 
    5068.82, 5078.408, 5077.996, 5085.024, 5088.664, 5097.227, 5101.399, 
    5111.218,
  5104.219, 5083.402, 5067.931, 5062.283, 5063.402, 5066.468, 5074.822, 
    5078.92, 5081.151, 5089.202, 5092.917, 5097.374, 5103.081, 5109.664, 
    5117.534,
  5116.222, 5096.927, 5080.305, 5071.054, 5069.212, 5074.021, 5076.996, 
    5084.409, 5089.206, 5089.978, 5092.377, 5098.139, 5104.212, 5111.233, 
    5120.185,
  5131.876, 5112.773, 5095.38, 5083.684, 5075.068, 5073.479, 5076.077, 
    5078.164, 5078.157, 5081.011, 5085.217, 5092.594, 5102.297, 5113.048, 
    5125.362,
  5150.343, 5131.388, 5114.893, 5102.211, 5092.196, 5084.712, 5078.378, 
    5076.858, 5075.258, 5075.034, 5079.225, 5090.56, 5103.522, 5117.806, 
    5135.303,
  5170.923, 5148.567, 5133.421, 5121.802, 5109.64, 5100.389, 5092.881, 
    5084.875, 5079.759, 5080.259, 5086.822, 5098.815, 5114.509, 5134, 5155.432,
  5220.375, 5205.972, 5196.5, 5185.473, 5173.897, 5160.727, 5142.17, 5125.2, 
    5101.208, 5067.478, 5029.519, 4984.564, 4941.575, 4913.162, 4911.73,
  5228.468, 5210.33, 5198.65, 5185.315, 5173.568, 5157.153, 5147.191, 
    5124.822, 5106.449, 5083.542, 5050.164, 5012.755, 4971.25, 4941.52, 
    4929.261,
  5237.888, 5216.486, 5201.08, 5187.2, 5171.006, 5160.654, 5140.217, 
    5133.556, 5117.06, 5097.951, 5073.385, 5042.05, 5007.96, 4975.935, 
    4957.738,
  5247.719, 5223.098, 5203.192, 5185.772, 5169.777, 5152.413, 5143.492, 
    5125.408, 5118.286, 5108.778, 5091.973, 5068.897, 5043.998, 5018.46, 
    4999.535,
  5258.359, 5231.98, 5208.232, 5187.487, 5169.46, 5152.507, 5135.341, 
    5125.202, 5117.622, 5114.081, 5106.702, 5090.527, 5074.483, 5056.52, 
    5043.956,
  5268.209, 5240.977, 5214.131, 5189.853, 5167.645, 5148.169, 5131.678, 
    5114.222, 5108.732, 5113.891, 5113.695, 5107.258, 5097.383, 5087.491, 
    5079.459,
  5277.232, 5250.534, 5222.589, 5196.306, 5171.031, 5148.32, 5127.22, 
    5110.958, 5103.547, 5108.596, 5115.161, 5117.057, 5114.584, 5111.64, 
    5108.574,
  5285.84, 5257.492, 5229.872, 5202.675, 5174.738, 5150.146, 5127.878, 
    5106.171, 5094.525, 5100.687, 5111.705, 5120.322, 5124.726, 5127.808, 
    5130.292,
  5292.484, 5265.488, 5238.696, 5210.099, 5182.685, 5157.741, 5134.408, 
    5113.352, 5099.218, 5098.143, 5108.673, 5121.562, 5130.785, 5137.735, 
    5144.303,
  5299.965, 5271.871, 5243.742, 5216.113, 5188.566, 5164.863, 5144.587, 
    5124.182, 5109.857, 5107.241, 5115.1, 5126.406, 5135.78, 5144.765, 5153.93,
  5355.981, 5326.38, 5297.473, 5263.915, 5232.907, 5200.637, 5169.739, 
    5141.989, 5124.05, 5100.173, 5067.523, 5021.561, 4976.563, 4944.202, 
    4928.658,
  5351.06, 5321.69, 5292.868, 5259.036, 5228.493, 5191.595, 5172.68, 
    5137.495, 5124.239, 5107.69, 5077.199, 5038.033, 4994.041, 4965.452, 
    4948.879,
  5347.191, 5318.854, 5289.676, 5257.885, 5223.585, 5197.738, 5160.024, 
    5144.338, 5128.746, 5116.83, 5090.916, 5058.259, 5019.946, 4987.533, 
    4968.266,
  5342.936, 5314.542, 5285.886, 5253.06, 5220.972, 5186.705, 5166.863, 
    5139.151, 5133.017, 5124.634, 5106.779, 5080.872, 5049.688, 5020.094, 
    4995.177,
  5339.449, 5311.549, 5283.96, 5250.799, 5219.117, 5186.771, 5160.135, 
    5141.645, 5138.381, 5132.694, 5121.024, 5100.812, 5077.285, 5050.764, 
    5028.369,
  5335.788, 5308.359, 5279.568, 5248.461, 5214.736, 5182.046, 5161.892, 
    5140.82, 5138.752, 5139.254, 5132.06, 5118.944, 5099.515, 5078.279, 
    5056.693,
  5332.925, 5306.339, 5278.255, 5247.893, 5213.245, 5181.882, 5160.951, 
    5143.83, 5141.7, 5144.32, 5140.547, 5132.626, 5117.74, 5100.635, 5080.706,
  5330.973, 5303.351, 5276.035, 5245.604, 5209.553, 5180.213, 5162.81, 
    5144.197, 5141.072, 5147.075, 5146.356, 5141.555, 5130.492, 5117.83, 
    5101.494,
  5328.84, 5302.345, 5276.231, 5245.389, 5211.373, 5181.749, 5164.894, 
    5148.553, 5142.658, 5148.126, 5148.575, 5145.812, 5138.058, 5128.428, 
    5116.231,
  5327.512, 5299.734, 5274.324, 5244.892, 5210.313, 5181.941, 5168.139, 
    5152.041, 5143.677, 5147.205, 5149.052, 5146.71, 5141.245, 5134.668, 
    5125.716,
  5363.641, 5339.406, 5317.307, 5293.528, 5271.25, 5242.751, 5212.103, 
    5189.458, 5172.267, 5161.963, 5153.77, 5139.383, 5118.431, 5091.135, 
    5067.996,
  5356.197, 5330.413, 5307.174, 5282.782, 5259.038, 5223.611, 5199.417, 
    5174.083, 5160.559, 5157.359, 5150.334, 5139.425, 5119.973, 5099.142, 
    5073.688,
  5351.137, 5325.09, 5300.742, 5276.394, 5248.268, 5220.945, 5182.394, 
    5172.104, 5155.412, 5151.914, 5146.519, 5137.93, 5120.707, 5100.441, 
    5079.272,
  5347.38, 5320.208, 5295.381, 5267.909, 5240.723, 5200.834, 5183.671, 
    5157.288, 5149.217, 5146.429, 5143.004, 5135.332, 5119.805, 5102.641, 
    5083.263,
  5345.27, 5318.164, 5292.833, 5263.992, 5235.181, 5199.702, 5173.156, 
    5159.643, 5144.718, 5141.454, 5138.934, 5131.396, 5116.456, 5099.837, 
    5083.715,
  5343.809, 5316.353, 5289.373, 5260.158, 5229.612, 5193.378, 5173.421, 
    5152.759, 5139.773, 5138.712, 5134.661, 5127.045, 5111.92, 5097.597, 
    5082.847,
  5343.054, 5316.787, 5289.683, 5258.854, 5229.535, 5193.789, 5172.671, 
    5155.662, 5141.375, 5136.265, 5131.005, 5121.772, 5106.627, 5093.005, 
    5077.709,
  5343.332, 5316.447, 5288.616, 5257.005, 5227.205, 5193.193, 5174.304, 
    5155.065, 5140.31, 5135.878, 5128.638, 5117.875, 5102.787, 5088.603, 
    5071.946,
  5343.697, 5318.057, 5290.663, 5257.772, 5229.804, 5196.5, 5177.265, 
    5160.671, 5145.506, 5137.643, 5127.701, 5115.898, 5099.641, 5082.197, 
    5061.629,
  5344.814, 5317.875, 5290.17, 5257.424, 5229.798, 5198.261, 5180.821, 
    5164.518, 5148.809, 5140.771, 5129.409, 5116.726, 5098.496, 5077.496, 
    5053.343,
  5373.774, 5347.798, 5319.373, 5286.067, 5256.653, 5227.247, 5198.209, 
    5178.599, 5159.162, 5140.243, 5127.388, 5120.497, 5117.604, 5116.428, 
    5115.388,
  5374.928, 5347.784, 5317.612, 5282.135, 5250.947, 5216.196, 5194.536, 
    5167.038, 5147.209, 5133.685, 5120.252, 5113.44, 5108.698, 5106.944, 
    5102.167,
  5375.737, 5348.472, 5317.043, 5281.729, 5246.582, 5220.038, 5183.438, 
    5170.616, 5146.559, 5128.886, 5114.224, 5107.233, 5099.391, 5094.106, 
    5086.706,
  5375.724, 5347.312, 5316.019, 5278.25, 5244.349, 5208.186, 5188.14, 
    5158.401, 5138.584, 5125.053, 5108.918, 5098.274, 5087.177, 5078.224, 
    5068.836,
  5375.142, 5346.871, 5316.385, 5278.007, 5243.201, 5210.59, 5180.275, 
    5163.466, 5141.007, 5118.296, 5102.374, 5085.583, 5071.463, 5058.58, 
    5049.583,
  5373.578, 5345.242, 5314.3, 5276.672, 5240.181, 5207.933, 5181.826, 
    5155.483, 5131.501, 5114.066, 5092.643, 5072.959, 5054.947, 5040.93, 
    5030.864,
  5371.219, 5344.098, 5314.065, 5276.778, 5241.474, 5209.941, 5181.309, 
    5160.199, 5134.989, 5110.107, 5085.802, 5064.124, 5043.215, 5029.715, 
    5019.203,
  5368.357, 5341.585, 5311.465, 5275.253, 5239.859, 5210.145, 5182.907, 
    5158.085, 5131.49, 5109.697, 5084.36, 5060.333, 5039.044, 5025.993, 
    5018.252,
  5364.515, 5339.929, 5311.114, 5275.964, 5242.768, 5213.641, 5185.98, 
    5163.625, 5138.004, 5113.66, 5087.306, 5063.268, 5041.963, 5029.82, 
    5022.542,
  5360.647, 5336.086, 5307.406, 5274.316, 5242.432, 5215.363, 5189.559, 
    5165.789, 5140.989, 5119.714, 5095.717, 5072.855, 5052.992, 5042.352, 
    5036.199,
  5404.487, 5382.597, 5357.474, 5327.497, 5293.623, 5259.089, 5225.065, 
    5200.962, 5179.593, 5155.401, 5136.762, 5121.581, 5110.751, 5102.846, 
    5101.42,
  5396.3, 5374.178, 5348.963, 5317.473, 5283.208, 5245.351, 5221.877, 
    5191.798, 5168.791, 5150.2, 5129.988, 5112.227, 5097.538, 5089.253, 
    5084.752,
  5388.841, 5367.954, 5341.716, 5311.237, 5274.404, 5249.124, 5209.548, 
    5196.627, 5172.724, 5147.845, 5124.246, 5104.447, 5085.345, 5073.434, 
    5068.063,
  5382.249, 5361.107, 5335.596, 5302.391, 5268.731, 5233.801, 5216.061, 
    5188.604, 5167.262, 5148.714, 5122.749, 5099.007, 5076.844, 5060.003, 
    5051.571,
  5377.543, 5356.475, 5331.942, 5298.346, 5266.381, 5236.491, 5210.101, 
    5194.284, 5177.341, 5149.238, 5126.043, 5097.212, 5072.861, 5049.664, 
    5038.506,
  5373.902, 5353.319, 5328.111, 5296.289, 5263.11, 5233.416, 5212.835, 
    5193.09, 5174.975, 5155.348, 5130.302, 5100.822, 5072.609, 5046.173, 
    5029.754,
  5371.232, 5352.409, 5327.779, 5297.729, 5267.131, 5238.29, 5213.77, 
    5200.189, 5184.716, 5162.491, 5136.357, 5106.65, 5074.503, 5044.758, 
    5023.597,
  5369.253, 5351.676, 5327.761, 5299.971, 5269.535, 5241.55, 5218.397, 
    5200.848, 5185.237, 5168.247, 5143.863, 5113.791, 5080.045, 5046.208, 
    5020.267,
  5367.597, 5351.61, 5329.907, 5304.834, 5277.907, 5250.179, 5224.505, 
    5207.81, 5193.474, 5174.235, 5150.279, 5121.626, 5087.385, 5050.532, 
    5020.109,
  5365.765, 5350.112, 5331.085, 5308.881, 5282.602, 5256.345, 5231.657, 
    5210.409, 5194.649, 5177.869, 5156.391, 5130.035, 5096.881, 5058.643, 
    5023.718,
  5445.806, 5422.126, 5396.785, 5368.527, 5342.764, 5322.634, 5307.936, 
    5297.342, 5281.997, 5258.688, 5236.381, 5212.519, 5193.63, 5177.657, 
    5166.429,
  5448.025, 5424.377, 5398.851, 5371.346, 5345.724, 5322.916, 5312.894, 
    5294.888, 5278.69, 5260.435, 5237.131, 5212.401, 5191.189, 5175.07, 
    5159.895,
  5449.66, 5426.621, 5401.414, 5375.802, 5348.592, 5331.743, 5309.744, 
    5302.104, 5283.02, 5259.24, 5235.951, 5211.654, 5188.338, 5170.162, 
    5151.695,
  5449.199, 5426.385, 5401.989, 5376.291, 5351.566, 5327.711, 5315.232, 
    5293.324, 5276.27, 5257.808, 5232.538, 5208.224, 5184.971, 5165.207, 
    5143.096,
  5446.818, 5424.795, 5401.688, 5376.822, 5353.412, 5331.739, 5310.874, 
    5297.705, 5278.978, 5251.956, 5229.903, 5202.194, 5180.199, 5156.828, 
    5133.613,
  5441.596, 5419.664, 5396.597, 5373.828, 5350.773, 5329.286, 5311.026, 
    5288.648, 5268.562, 5246.929, 5223.091, 5195.914, 5173.376, 5148.771, 
    5122.965,
  5433.661, 5413.506, 5390.501, 5368.54, 5347.74, 5327.892, 5307.917, 
    5290.139, 5268.727, 5242.343, 5216.373, 5189.174, 5164.661, 5139.194, 
    5110.096,
  5424.613, 5403.864, 5380.314, 5360.18, 5339.982, 5322.056, 5303.795, 
    5282.618, 5260.204, 5236.052, 5209.438, 5181.192, 5156.219, 5129.187, 
    5098.646,
  5414.797, 5394.138, 5371.183, 5350.829, 5332.786, 5315.598, 5297.3, 
    5278.443, 5256.159, 5229.698, 5202.026, 5172.73, 5146.716, 5118.497, 
    5086.958,
  5405.125, 5381.934, 5358.899, 5340.669, 5322.542, 5305.29, 5287.549, 
    5266.014, 5243.952, 5219.754, 5193.139, 5163.577, 5137.5, 5108.717, 
    5076.762,
  5533.108, 5509.543, 5486.41, 5460.799, 5437.783, 5414.406, 5391.234, 
    5373.114, 5355.959, 5336.781, 5322.623, 5308.337, 5295.289, 5282.988, 
    5274.46,
  5522.261, 5499.324, 5477.164, 5452.445, 5429.372, 5403.064, 5387.121, 
    5361.613, 5346.23, 5334.903, 5320.477, 5307.251, 5294.648, 5283.951, 
    5274.146,
  5509.405, 5488.252, 5466.049, 5444.119, 5418.833, 5401.515, 5371.242, 
    5363.454, 5342.932, 5327.524, 5314.505, 5302.768, 5289.45, 5278.585, 
    5268.074,
  5493.628, 5473.836, 5453.085, 5430.974, 5408.884, 5383.174, 5369.599, 
    5341.723, 5330.43, 5319.109, 5304.158, 5292.087, 5279.74, 5268.559, 
    5257.519,
  5477.814, 5459.622, 5440.133, 5419.351, 5397.669, 5376.041, 5351.896, 
    5340.722, 5321.051, 5302.432, 5290.235, 5274.426, 5263.209, 5250.227, 
    5241.17,
  5461.466, 5445.003, 5425.562, 5405.895, 5382.151, 5359.866, 5339.812, 
    5316.731, 5298.946, 5283.477, 5265.422, 5249.542, 5236.771, 5224.911, 
    5216.151,
  5446.859, 5432.112, 5412.886, 5392.383, 5369.539, 5345.843, 5322.195, 
    5301.774, 5277.974, 5253.22, 5233.22, 5215.023, 5200.284, 5189.81, 
    5182.293,
  5434.366, 5418.637, 5398.574, 5377.44, 5351.504, 5326.723, 5300.021, 
    5270.578, 5241.793, 5216.505, 5191.919, 5171.762, 5157.211, 5148.158, 
    5143.29,
  5422.805, 5408.07, 5387.586, 5363.648, 5336.306, 5306.343, 5272.362, 
    5240.127, 5207.214, 5175.172, 5149.828, 5130.041, 5116.715, 5109.203, 
    5106.344,
  5414.371, 5397.32, 5374.095, 5347.649, 5314.347, 5278.137, 5239.797, 
    5200.8, 5166.568, 5136.615, 5113.193, 5096.193, 5085.745, 5080.071, 
    5077.89,
  5454.753, 5435.97, 5421.438, 5406.688, 5394.879, 5380.817, 5363.196, 
    5348.423, 5331.439, 5313.116, 5301.019, 5291.369, 5284.423, 5277.903, 
    5274.465,
  5439.324, 5424.114, 5411.787, 5398.317, 5386.243, 5367.133, 5353.85, 
    5327.283, 5309.495, 5296.864, 5283.466, 5275.727, 5269.936, 5268.251, 
    5265.534,
  5429.352, 5418.119, 5405.938, 5394.274, 5376.937, 5362.631, 5330.27, 
    5317.107, 5290.174, 5272.216, 5259.765, 5252.95, 5247.636, 5247.113, 
    5247.831,
  5424.149, 5413.033, 5401.609, 5386.071, 5367.006, 5340.221, 5320.819, 
    5279.657, 5260.921, 5244.884, 5231.288, 5222.767, 5219.125, 5218.381, 
    5221.434,
  5421.729, 5411.588, 5399.034, 5380.25, 5357.089, 5328.389, 5289.833, 
    5266.771, 5238.788, 5214.255, 5202.98, 5189.937, 5185.145, 5180.778, 
    5185.278,
  5421.825, 5409.795, 5393.889, 5371.527, 5342.842, 5307.901, 5269.423, 
    5230.479, 5205.506, 5190.171, 5172.588, 5160.03, 5151.563, 5145.821, 
    5146.098,
  5422.593, 5408.792, 5390.35, 5363.614, 5332.379, 5290.419, 5244.953, 
    5215.989, 5189.415, 5166.886, 5149.91, 5136.773, 5125.076, 5117.622, 
    5113.519,
  5423.165, 5406.104, 5384.516, 5353.501, 5317.297, 5271.315, 5225.841, 
    5194.729, 5169.066, 5151.928, 5133.266, 5118.586, 5105.568, 5095.798, 
    5088.451,
  5423.218, 5404.848, 5380.368, 5345.808, 5307.839, 5257.748, 5213.751, 
    5189.208, 5162.941, 5140.727, 5119.825, 5103.762, 5088.529, 5077.128, 
    5067.26,
  5423.43, 5400.74, 5373.079, 5337.148, 5295.213, 5245.057, 5206.809, 
    5179.602, 5152.195, 5129.847, 5107.229, 5089.192, 5073.385, 5061.73, 
    5051.344,
  5441.712, 5415.572, 5388.348, 5358.289, 5327.541, 5293.655, 5258.684, 
    5232.291, 5205.948, 5180.793, 5166.658, 5160.173, 5160.018, 5165.544, 
    5175.458,
  5448.057, 5420.855, 5391.331, 5358.988, 5326.385, 5284.986, 5256.168, 
    5217.609, 5189.177, 5169.947, 5154.354, 5146.551, 5145.057, 5150.836, 
    5159.911,
  5454.002, 5426.624, 5395.181, 5363.186, 5325.505, 5293.948, 5244.462, 
    5223.845, 5191.525, 5164.482, 5145.601, 5136.642, 5132.177, 5136.122, 
    5144.572,
  5458.045, 5429.734, 5398.099, 5362.974, 5327.537, 5283.724, 5253.05, 
    5211.156, 5181.674, 5161.05, 5140.622, 5129.066, 5123.619, 5124.969, 
    5131.398,
  5461.407, 5433.079, 5401.673, 5365.692, 5330.126, 5290.1, 5247.433, 
    5220.577, 5190.588, 5157.005, 5137.746, 5121.708, 5115.736, 5114.162, 
    5119.652,
  5463.206, 5434.68, 5402.027, 5367.653, 5330.095, 5290.265, 5252.574, 
    5215.194, 5181.631, 5157.625, 5134.191, 5116.824, 5107.732, 5105.021, 
    5109.518,
  5463.597, 5436.685, 5404.099, 5369.852, 5333.774, 5294.595, 5254.058, 
    5223.08, 5189.955, 5158.496, 5132.525, 5113.175, 5099.749, 5095.336, 
    5097.712,
  5463.034, 5435.891, 5402.924, 5370.038, 5333.066, 5295.621, 5257.078, 
    5221.725, 5187.062, 5159.203, 5132.769, 5110.879, 5094.424, 5086.689, 
    5085.88,
  5461.241, 5435.769, 5403.813, 5370.674, 5335.479, 5297.903, 5258.89, 
    5226.609, 5193.512, 5161.897, 5133.486, 5109.627, 5090.336, 5079.222, 
    5075.079,
  5458.592, 5431.468, 5400.115, 5368.886, 5333.016, 5296.278, 5259.033, 
    5224.341, 5191.627, 5162.297, 5134.508, 5109.107, 5087.686, 5073.785, 
    5066.352,
  5497.081, 5467.053, 5437.551, 5406.764, 5376.479, 5345.138, 5309.008, 
    5279.282, 5247.766, 5213.065, 5186.432, 5166.417, 5154.583, 5151.333, 
    5157.686,
  5497.796, 5467.668, 5438.365, 5407.887, 5378.425, 5343.099, 5316.968, 
    5274.439, 5243.067, 5215.883, 5188.024, 5166.062, 5151.423, 5145.405, 
    5148.134,
  5496.625, 5466.989, 5437.459, 5408.748, 5376.423, 5351.776, 5307.612, 
    5288.136, 5249.881, 5216.308, 5187.472, 5164.955, 5147.426, 5138.934, 
    5138.203,
  5492.412, 5462.574, 5433.603, 5403.677, 5374.612, 5339.49, 5314.502, 
    5268.302, 5239.113, 5212.274, 5184.365, 5161.322, 5143.495, 5132.361, 
    5129.661,
  5486.446, 5457.139, 5428.576, 5399.283, 5369.669, 5338.358, 5301.606, 
    5275.235, 5239.801, 5202.627, 5179.661, 5155.456, 5138.695, 5124.404, 
    5120.806,
  5477.549, 5448.318, 5419.421, 5390.999, 5359.686, 5327.916, 5294.747, 
    5254.676, 5219.397, 5193.71, 5169.655, 5149.693, 5132.147, 5118.04, 
    5111.576,
  5466.372, 5438.9, 5410.296, 5381.027, 5350.098, 5315.905, 5279.101, 
    5245.918, 5211.144, 5182.029, 5159.543, 5142.209, 5124.506, 5111.094, 
    5101.865,
  5453.654, 5426.95, 5397.414, 5368.276, 5334.353, 5299.119, 5261.549, 
    5222.437, 5190.34, 5168.578, 5149.486, 5133.522, 5117, 5103.02, 5092.468,
  5440.26, 5415.417, 5386.564, 5355.3, 5320.022, 5282.264, 5242.415, 
    5208.138, 5180.655, 5158.126, 5140.063, 5124.75, 5108.235, 5094.136, 
    5083.774,
  5427.41, 5401.351, 5370.745, 5339.012, 5300.46, 5262.434, 5223.68, 
    5189.326, 5165.016, 5147.321, 5131.502, 5115.864, 5099.556, 5085.789, 
    5076.408,
  5429.18, 5409.384, 5386.724, 5360.991, 5336.649, 5313.485, 5288.626, 
    5270.586, 5250.89, 5228.266, 5209.423, 5194.103, 5182.182, 5174.137, 
    5171.302,
  5414.376, 5392.031, 5367.962, 5342.023, 5316.785, 5290.467, 5271.303, 
    5242.339, 5220.357, 5204.37, 5184.36, 5170.957, 5161.72, 5159.973, 
    5158.116,
  5398.296, 5375.448, 5350.233, 5324.812, 5296.026, 5277.897, 5241.865, 
    5230.353, 5199.107, 5174.218, 5155.268, 5144.125, 5139.108, 5141.178, 
    5144.816,
  5382.224, 5358.917, 5333.448, 5305.119, 5278.043, 5246.715, 5229.227, 
    5187.526, 5163.744, 5142.488, 5123.99, 5116.889, 5117.894, 5124.219, 
    5131.76,
  5368.556, 5345.34, 5318.618, 5288.239, 5257.901, 5231.074, 5194.698, 
    5176.616, 5145.127, 5112.849, 5101.649, 5096.211, 5101.804, 5109.838, 
    5120.156,
  5357.649, 5331.93, 5302.359, 5270.754, 5239.509, 5207.636, 5177.713, 
    5140.877, 5114.354, 5099.275, 5087.619, 5086.269, 5091.957, 5100.281, 
    5109.839,
  5347.23, 5320.978, 5289.095, 5256.35, 5223.228, 5191.924, 5158.717, 
    5135.796, 5113.65, 5093.644, 5083.598, 5082.327, 5085.32, 5092.304, 
    5099.961,
  5338.495, 5309.921, 5275.826, 5241.69, 5208.782, 5177.803, 5149.188, 
    5122.393, 5102.396, 5091.382, 5083.542, 5080.465, 5081.009, 5084.821, 
    5090.191,
  5331.311, 5301.623, 5265.716, 5231.137, 5198.627, 5169.849, 5144.04, 
    5125.702, 5108.879, 5093.456, 5082.988, 5077.439, 5074.797, 5075.643, 
    5078.88,
  5325.729, 5291.963, 5254.729, 5220.615, 5190.469, 5164.463, 5143.231, 
    5122.375, 5106.187, 5093.107, 5082.414, 5073.637, 5068.167, 5066.293, 
    5067.562,
  5285.19, 5257.106, 5231.075, 5203.16, 5175.385, 5149.103, 5123.287, 
    5106.149, 5093.216, 5083.774, 5084.299, 5095.126, 5112.88, 5132.834, 
    5153.121,
  5276.226, 5246.082, 5218.157, 5187.328, 5158.242, 5126.354, 5107.915, 
    5083.051, 5068.018, 5061.388, 5060.538, 5070.104, 5089.032, 5113.19, 
    5135.896,
  5269.115, 5238.431, 5208.714, 5178.071, 5145.521, 5124.953, 5090.18, 
    5079.12, 5059.517, 5045.502, 5040.386, 5050.426, 5070.26, 5094.406, 
    5121.421,
  5262.188, 5231.241, 5201.78, 5170.04, 5140.964, 5111.569, 5095.356, 
    5066.393, 5049.583, 5038.552, 5030.438, 5038.028, 5056.596, 5081.925, 
    5108.914,
  5258.568, 5228.459, 5199.4, 5168.75, 5142.622, 5117.591, 5091.791, 
    5073.979, 5057.373, 5038.477, 5031.554, 5033.423, 5050.554, 5070.841, 
    5098.974,
  5256.864, 5227.304, 5198.422, 5171.169, 5144.148, 5121.22, 5099.584, 
    5076.031, 5057.04, 5046.969, 5038.248, 5038.246, 5049.806, 5067.969, 
    5091.755,
  5257.911, 5230.199, 5202.14, 5177.035, 5153.523, 5130.957, 5106.758, 
    5088.221, 5070.434, 5054.855, 5046.661, 5046.408, 5052.5, 5067.928, 
    5087.449,
  5260.658, 5234.05, 5207.174, 5184.181, 5159.829, 5138.768, 5116.231, 
    5094.173, 5074.599, 5062.953, 5054.634, 5053.81, 5057.692, 5070.011, 
    5085.365,
  5266.98, 5242.157, 5216.423, 5194.705, 5172.893, 5150.323, 5125.956, 
    5105.603, 5086.042, 5070.01, 5059.761, 5057.646, 5060.581, 5070.09, 
    5083.353,
  5275.584, 5250.19, 5226.585, 5206.307, 5182.141, 5159.562, 5135.694, 
    5111.994, 5090.733, 5074.762, 5063.49, 5059.474, 5060.923, 5069.206, 
    5080.953,
  5274.243, 5238.24, 5205.558, 5172.02, 5142.307, 5115.976, 5090.421, 
    5073.784, 5061.435, 5049.23, 5045.489, 5050.368, 5066.802, 5092.999, 
    5124.096,
  5281.656, 5243.937, 5208.722, 5172.553, 5140.966, 5107.736, 5090.052, 
    5063.647, 5048.918, 5039.694, 5032.141, 5030.311, 5035.286, 5059.608, 
    5089.963,
  5291.651, 5252.483, 5214.24, 5177.255, 5139.992, 5115.043, 5080.561, 
    5067.85, 5050.112, 5037.048, 5026.259, 5019.066, 5018.877, 5031.695, 
    5060.394,
  5301.099, 5260.443, 5220.504, 5179.565, 5142.851, 5106.719, 5088.187, 
    5061.111, 5047.399, 5037.991, 5026.445, 5016.069, 5013.427, 5022.886, 
    5045.493,
  5312.454, 5271.113, 5229.789, 5186.933, 5148.411, 5114.158, 5085.236, 
    5068.378, 5056.401, 5042.619, 5032.213, 5019.373, 5018.076, 5022.763, 
    5044.078,
  5323.406, 5281.722, 5237.806, 5194.754, 5152.663, 5116.601, 5091.537, 
    5070.591, 5058.185, 5052.583, 5043.816, 5035.169, 5031.823, 5038.237, 
    5053.915,
  5335.114, 5294.998, 5250.204, 5206.406, 5163.884, 5125.967, 5095.764, 
    5079.325, 5069.954, 5063.209, 5058.86, 5056.053, 5056.365, 5061.862, 
    5074.41,
  5346.599, 5307.866, 5262.132, 5217.687, 5173.262, 5134.636, 5103.949, 
    5083.187, 5073.375, 5071.98, 5072.572, 5073.953, 5078.286, 5086.201, 
    5097.143,
  5358.921, 5323.307, 5278.529, 5234.207, 5191.064, 5150.004, 5114.61, 
    5092.776, 5082.651, 5079.845, 5081.82, 5086.993, 5093.188, 5102.412, 
    5113.159,
  5370.902, 5337.445, 5295.263, 5251.389, 5206.161, 5165.631, 5130.158, 
    5101.634, 5087.852, 5085.453, 5089.018, 5095.767, 5104.129, 5113.878, 
    5124.828,
  5348.679, 5306.256, 5258.361, 5208.819, 5164.389, 5138.485, 5114.596, 
    5098.539, 5086.397, 5076.581, 5082.741, 5099.737, 5123.761, 5151.623, 
    5178.894,
  5345.92, 5305.146, 5258.047, 5209.241, 5167.885, 5140.078, 5126.151, 
    5102.157, 5086.452, 5078.524, 5078.709, 5091.911, 5113.072, 5142.844, 
    5166.959,
  5344.124, 5306.096, 5259.766, 5213.852, 5172.673, 5155.646, 5130.326, 
    5117.236, 5100.508, 5084.27, 5077.942, 5084.572, 5101.171, 5124.827, 
    5153.159,
  5341.628, 5306.154, 5262.091, 5215.687, 5180.559, 5157.211, 5148.994, 
    5128.893, 5108.337, 5092.746, 5079.885, 5078.374, 5088.961, 5110.506, 
    5135.746,
  5340.482, 5308.291, 5266.012, 5221.425, 5188.813, 5170.539, 5159.088, 
    5142.861, 5132.043, 5107.445, 5090.819, 5076.854, 5078.504, 5090.915, 
    5115.366,
  5339.717, 5310.434, 5268.808, 5227.318, 5193.631, 5176.353, 5173.101, 
    5160.354, 5143.625, 5127.089, 5110.064, 5089.629, 5076.598, 5077.559, 
    5095.051,
  5340.214, 5314.378, 5274.437, 5234.773, 5202.37, 5184.239, 5179.505, 
    5175.22, 5165.787, 5149.186, 5130.293, 5112.703, 5092.916, 5076.983, 
    5078.505,
  5341.532, 5318.469, 5280.505, 5242.262, 5208.263, 5188.142, 5186.434, 
    5185.137, 5177.547, 5167.441, 5152.516, 5134.562, 5116.373, 5098.501, 
    5084.612,
  5344.433, 5324.562, 5289.881, 5252.474, 5220.441, 5196.741, 5189.469, 
    5193.149, 5192.428, 5184.934, 5172.811, 5157.881, 5140.709, 5123.828, 
    5108.133,
  5348.314, 5330.727, 5299.835, 5263.708, 5229.632, 5205.011, 5194.328, 
    5195.787, 5198.203, 5196.341, 5189.396, 5177.529, 5163.822, 5149.352, 
    5135.635,
  5315.725, 5298.936, 5281.152, 5260.623, 5240.042, 5227.013, 5204.231, 
    5179.663, 5153.112, 5138.117, 5147.826, 5160.447, 5172.204, 5179.445, 
    5184.97,
  5302.558, 5286.023, 5270.01, 5250.305, 5235.198, 5227.084, 5212.787, 
    5182.84, 5156.334, 5141.485, 5148.202, 5161.316, 5174.026, 5184.562, 
    5190.752,
  5291.82, 5275.942, 5259.95, 5242.997, 5234.283, 5235.067, 5215.465, 
    5197.638, 5173.843, 5151.412, 5149.268, 5159.698, 5173.789, 5184.935, 
    5193.006,
  5283.586, 5265.094, 5248.23, 5236.128, 5236.966, 5234.198, 5228.092, 
    5207.915, 5184.083, 5165.449, 5150.756, 5157.438, 5170.166, 5185.368, 
    5195.592,
  5278.424, 5257.474, 5243.811, 5236.893, 5242.068, 5242.887, 5234.855, 
    5218.631, 5204.797, 5179.101, 5163.082, 5152.518, 5163.778, 5179.129, 
    5193.389,
  5278.708, 5256.743, 5242.549, 5239.384, 5244.596, 5248.094, 5244.546, 
    5231.093, 5212.101, 5194.696, 5175.874, 5157.01, 5154.6, 5171.34, 5188.324,
  5286.055, 5262.244, 5248.586, 5245.345, 5251.071, 5256.497, 5251.396, 
    5243.395, 5229.662, 5210.248, 5189.576, 5170.724, 5154.222, 5159.586, 
    5178.478,
  5300.766, 5273.486, 5255.66, 5251.909, 5255.065, 5261.641, 5260.849, 
    5252.441, 5237.964, 5222.568, 5204.3, 5185.364, 5167.836, 5156.462, 
    5166.951,
  5316.565, 5291.431, 5268.436, 5260.947, 5262.849, 5267.688, 5266.915, 
    5262.118, 5252.341, 5236.76, 5218.458, 5200.224, 5182.921, 5168.161, 
    5160.527,
  5331.409, 5310.228, 5284.712, 5268.99, 5267.037, 5270.329, 5272.144, 
    5267.415, 5258.735, 5246.475, 5231.126, 5214.292, 5197.223, 5182.7, 
    5170.245,
  5270.064, 5267.675, 5265.128, 5258.854, 5253.381, 5251.713, 5240.846, 
    5226.942, 5209.08, 5188.538, 5185.479, 5190.6, 5194.576, 5191.699, 
    5183.364,
  5256.793, 5256.167, 5256.442, 5254.365, 5255.193, 5251.025, 5243.029, 
    5224.011, 5205.502, 5190.277, 5185.805, 5190.138, 5192.281, 5188.785, 
    5178.927,
  5253.254, 5252.663, 5256.102, 5259.953, 5259.417, 5257.362, 5243.073, 
    5230.886, 5214.068, 5194.431, 5185.619, 5188.917, 5190.418, 5186.681, 
    5175.859,
  5260.184, 5259.55, 5264.568, 5267.074, 5267.267, 5258.08, 5251.332, 
    5233.727, 5215.384, 5199.902, 5185.869, 5185.763, 5189.41, 5185.963, 
    5176.72,
  5275.149, 5273.838, 5277.217, 5277.04, 5274.751, 5266.784, 5254.9, 
    5240.795, 5227.626, 5205.012, 5190.744, 5182.334, 5187.264, 5186.169, 
    5180.923,
  5289.078, 5287.169, 5286.555, 5284.845, 5280.09, 5271.676, 5262.099, 
    5246.758, 5230.195, 5213.764, 5196.082, 5182.148, 5185.699, 5188.254, 
    5185.645,
  5298.731, 5295.382, 5293.241, 5289.958, 5285.042, 5277.303, 5265.67, 
    5254.568, 5241.63, 5224.005, 5205.574, 5189.774, 5185.188, 5191.09, 
    5191.197,
  5305.384, 5297.905, 5293.75, 5289.516, 5284.477, 5278.258, 5269.026, 
    5257.838, 5245.674, 5232.729, 5216.889, 5200.639, 5190.549, 5192.436, 
    5196.6,
  5309.219, 5301.314, 5292.814, 5287.034, 5283.118, 5278.107, 5269.622, 
    5261.358, 5252.832, 5241.869, 5227.599, 5212.5, 5200.105, 5194.939, 
    5199.026,
  5309.423, 5303.17, 5295.175, 5285.39, 5279.958, 5276.499, 5270.491, 
    5262.646, 5253.885, 5246.086, 5236.304, 5223.812, 5210.983, 5202.108, 
    5200.666,
  5292.786, 5289.949, 5286.886, 5282.022, 5276.565, 5268.86, 5257.485, 
    5246.473, 5233.481, 5216.563, 5201.722, 5195.371, 5194.889, 5196.052, 
    5197.511,
  5300.417, 5295.289, 5290.951, 5284.609, 5277.604, 5266.998, 5258.464, 
    5242.595, 5228.651, 5214.152, 5199.282, 5194.016, 5195.172, 5196.744, 
    5196.291,
  5307.668, 5301.455, 5294.59, 5287.654, 5278.081, 5270.266, 5254.213, 
    5244.459, 5229.984, 5213.458, 5197.32, 5191.435, 5191.852, 5192.355, 
    5189.3,
  5309.027, 5302.145, 5294.956, 5285.942, 5275.964, 5264.338, 5255.741, 
    5239.605, 5227.246, 5214.071, 5197.379, 5188.354, 5186.611, 5185.743, 
    5180.787,
  5308.558, 5301.504, 5293.857, 5283.24, 5273.884, 5264.318, 5250.834, 
    5241.357, 5230.293, 5214.254, 5199.056, 5186.444, 5182.754, 5178.45, 
    5172.826,
  5305.943, 5298.516, 5290.137, 5279.504, 5270.205, 5261.787, 5251.7, 
    5238.557, 5227.437, 5216.034, 5201.079, 5187.119, 5179.921, 5172.722, 
    5164.136,
  5303.886, 5297.479, 5289.104, 5278.658, 5271.508, 5263.628, 5252.39, 
    5242.646, 5231.547, 5218.126, 5203.261, 5188.917, 5176.952, 5167.724, 
    5154.82,
  5302.237, 5296.907, 5289.825, 5281.124, 5274.191, 5267.417, 5256.964, 
    5244.303, 5231.409, 5220.023, 5206.194, 5191.593, 5176.451, 5164.102, 
    5148.578,
  5300.664, 5298.1, 5293.997, 5288.116, 5282.829, 5275.597, 5264.037, 
    5251.755, 5237.548, 5223.431, 5209.295, 5195.166, 5178.845, 5162.327, 
    5145.273,
  5299.888, 5297.9, 5297.629, 5294.847, 5290.104, 5283.349, 5272.108, 
    5257.19, 5241.406, 5226.143, 5212.401, 5199.39, 5183.288, 5164.459, 
    5146.054,
  5336.579, 5324.366, 5313.89, 5302.496, 5290.613, 5278.035, 5264.065, 
    5252.198, 5240.142, 5227.128, 5215.689, 5204.242, 5197.083, 5193.694, 
    5191.296,
  5334.757, 5321.566, 5310.424, 5298.353, 5286.537, 5271.751, 5261.343, 
    5244.561, 5232.336, 5222.88, 5212.047, 5200.989, 5194.294, 5191.417, 
    5191.07,
  5334.234, 5321.61, 5310.323, 5299.539, 5285.504, 5275.289, 5255.679, 
    5246.019, 5231.431, 5218.73, 5208.026, 5198.174, 5190.108, 5185.906, 
    5184.508,
  5335.187, 5322.669, 5312.094, 5300.111, 5287.978, 5271.824, 5260.086, 
    5239.246, 5226.306, 5215.281, 5204.068, 5194.416, 5185.43, 5179.682, 
    5175.955,
  5336.336, 5325.223, 5316.275, 5304.973, 5292.91, 5277.624, 5258.091, 
    5243.619, 5227.876, 5210.533, 5200.244, 5188.561, 5180.375, 5172.062, 
    5167.739,
  5337.64, 5327.82, 5319.547, 5309.351, 5295.71, 5279.622, 5261.857, 
    5240.469, 5222.987, 5208.395, 5194.782, 5182.205, 5173.4, 5164.388, 
    5159.522,
  5338.556, 5331.29, 5324.156, 5314.135, 5300.988, 5284.246, 5263.949, 
    5245.158, 5226.527, 5206.42, 5190.208, 5176.399, 5165.396, 5155.485, 
    5150.001,
  5340.562, 5334.075, 5326.455, 5316.729, 5302.24, 5285.766, 5266.312, 
    5244.749, 5224.378, 5205.409, 5186.879, 5169.851, 5156.272, 5145.106, 
    5139.018,
  5343.27, 5337.612, 5329.916, 5319.299, 5305.594, 5288.678, 5268.464, 
    5248.761, 5228.373, 5206.412, 5184.469, 5163.729, 5146, 5132.194, 5126.265,
  5348.697, 5340.637, 5331.583, 5320.688, 5305.061, 5287.743, 5269.023, 
    5248.486, 5228.318, 5206.753, 5183.243, 5158.891, 5137.473, 5121.797, 
    5117.767,
  5339.441, 5327.639, 5318.339, 5305.983, 5292.312, 5276.251, 5258.632, 
    5244.766, 5231.084, 5216.526, 5206.402, 5198.561, 5193.404, 5191.076, 
    5191.738,
  5337.585, 5326.02, 5315.432, 5301.428, 5286.368, 5267.413, 5254.93, 
    5234.998, 5222.218, 5211.752, 5200.791, 5192.459, 5186.502, 5184.458, 
    5184.682,
  5337.227, 5325.6, 5313.036, 5298.128, 5279.88, 5266.337, 5243.137, 
    5235.318, 5218.076, 5205.317, 5194.542, 5185.785, 5178.318, 5175.216, 
    5175.458,
  5336.949, 5322.871, 5308.265, 5290.291, 5272.124, 5251.295, 5240.221, 
    5217.741, 5208.597, 5198.021, 5186.868, 5176.982, 5169.078, 5165.311, 
    5165.525,
  5336.389, 5320.76, 5303.374, 5282.549, 5262.247, 5243.066, 5223.13, 
    5214.357, 5199.519, 5186.834, 5177.408, 5165.456, 5157.49, 5152.505, 
    5154.083,
  5335.432, 5316.266, 5293.666, 5270.203, 5245.998, 5225.152, 5208.989, 
    5193.06, 5183.223, 5175.302, 5163.881, 5152.61, 5143.12, 5139.406, 
    5141.607,
  5333.326, 5310.815, 5282.757, 5254.576, 5228.051, 5205.627, 5189.803, 
    5181.063, 5172.401, 5161.395, 5150.617, 5137.267, 5126.159, 5124.427, 
    5129.555,
  5330.636, 5301.429, 5267.018, 5235.195, 5205.295, 5185.044, 5172.309, 
    5163.339, 5157.009, 5149.588, 5136.952, 5120.993, 5109.977, 5112.015, 
    5121.312,
  5327.836, 5294.282, 5255.954, 5219.972, 5190.347, 5170.787, 5160.279, 
    5155.943, 5150.088, 5139.354, 5124.387, 5106.537, 5099.521, 5107.368, 
    5120.009,
  5328.132, 5288.136, 5246.796, 5209.573, 5178.818, 5160.738, 5153.25, 
    5148.404, 5142.862, 5133.227, 5117.411, 5104.531, 5105.314, 5115.325, 
    5128.44,
  5300.11, 5288.958, 5280.089, 5271.908, 5265.716, 5259.091, 5252.855, 
    5249.483, 5244.771, 5238.82, 5235.761, 5230.974, 5225.025, 5218.289, 
    5214.984,
  5282.122, 5269.368, 5258.116, 5248.252, 5240.283, 5233.639, 5232.143, 
    5224.508, 5224.038, 5224.657, 5222.499, 5222.292, 5220.279, 5217.389, 
    5216.264,
  5265.633, 5250.712, 5236.826, 5225.809, 5213.983, 5209.94, 5197.404, 
    5204.143, 5197.439, 5201.415, 5205.875, 5210.155, 5212.464, 5213.417, 
    5214.522,
  5253.701, 5235.521, 5219.018, 5202.163, 5188.639, 5174.086, 5173.407, 
    5159.52, 5169.495, 5173.953, 5184.117, 5192.809, 5202.002, 5207.371, 
    5212.694,
  5245.535, 5224.637, 5204.425, 5184.776, 5166.747, 5150.698, 5135.106, 
    5135.038, 5130.333, 5139.482, 5158.318, 5173, 5188.28, 5197.902, 5208.053,
  5242.107, 5218.424, 5194.256, 5171.896, 5148.704, 5130.686, 5116.31, 
    5103.205, 5103.18, 5113.054, 5128.765, 5152.476, 5172.507, 5188.88, 
    5201.668,
  5242.738, 5218.859, 5193.604, 5170.122, 5147.302, 5126.12, 5109.1, 5100.41, 
    5093.195, 5095.066, 5111.982, 5136.089, 5157.991, 5178.377, 5194.288,
  5249.054, 5225.205, 5199.436, 5175.792, 5150.156, 5129.089, 5112.128, 
    5100.6, 5094.506, 5095.814, 5105.13, 5125.471, 5147.841, 5169.226, 5187.99,
  5259.887, 5236.876, 5211.849, 5187.938, 5162.417, 5137.124, 5117.964, 
    5108.82, 5101.354, 5097.923, 5104.066, 5120.566, 5139.587, 5161.292, 
    5182.302,
  5275.113, 5250.408, 5226.277, 5200.328, 5169.975, 5142.843, 5122.835, 
    5111.121, 5107.453, 5104.344, 5108.429, 5120.447, 5136.622, 5157.937, 
    5180.747,
  5275.029, 5262.151, 5250.612, 5239.976, 5231.156, 5223.279, 5217.033, 
    5215.503, 5215.283, 5217.292, 5224.909, 5234.424, 5244.205, 5250.41, 
    5251.077,
  5271.85, 5256.431, 5242.21, 5228.72, 5217.149, 5206.265, 5201.593, 
    5194.795, 5196.1, 5201.173, 5208.753, 5221.943, 5233.914, 5244.593, 
    5246.437,
  5270, 5252.206, 5235.832, 5220.979, 5206.134, 5197.495, 5183.72, 5183.801, 
    5178.795, 5184.122, 5195.205, 5210.788, 5226.522, 5239.014, 5243.787,
  5263.608, 5243.159, 5224.115, 5205.436, 5190.842, 5176.163, 5173.021, 
    5161.126, 5164.323, 5167.118, 5180.706, 5199.467, 5220.223, 5235.371, 
    5242.957,
  5256.303, 5233.58, 5210.993, 5190.243, 5172.388, 5159.778, 5148.768, 
    5151.468, 5148.305, 5152.404, 5167.424, 5189.584, 5214.994, 5232.446, 
    5243.522,
  5247.747, 5221.231, 5194.365, 5170.6, 5149.87, 5135.923, 5129.278, 
    5126.814, 5133.641, 5141.512, 5154.261, 5182.346, 5210.685, 5232.355, 
    5245.451,
  5239.517, 5210.895, 5180.397, 5153.459, 5130.851, 5115.242, 5107.884, 
    5113.172, 5120.819, 5129.738, 5146.018, 5176.952, 5208.963, 5233.021, 
    5250.121,
  5233.101, 5201.188, 5166.983, 5138.645, 5113.185, 5098.039, 5092.789, 
    5097.172, 5109.604, 5123.26, 5140.583, 5175.293, 5210.367, 5236.512, 
    5257.461,
  5228.859, 5195.715, 5160.672, 5130.939, 5106.15, 5090.942, 5086.288, 
    5095.247, 5107.999, 5119.76, 5140.681, 5178.631, 5214.098, 5242.373, 
    5266.523,
  5228.664, 5192.932, 5158.326, 5129.496, 5105.616, 5091.974, 5089.897, 
    5096.475, 5108.505, 5121.511, 5147.522, 5186.444, 5221.878, 5251.399, 
    5277.694,
  5276.955, 5254.873, 5237.14, 5223.667, 5215.466, 5210.353, 5208.551, 
    5210.5, 5212.99, 5214.692, 5218.232, 5222.7, 5231.211, 5243.055, 5259.118,
  5254.396, 5231.365, 5213.945, 5201.319, 5194.437, 5190.979, 5192.788, 
    5193.454, 5199.039, 5206.227, 5210.262, 5215.374, 5221.488, 5235.073, 
    5250.102,
  5231.849, 5208.621, 5191.687, 5180.691, 5174.095, 5175.317, 5172.923, 
    5182.894, 5186.613, 5194.678, 5201.57, 5207.968, 5214.691, 5225.961, 
    5241.887,
  5209.736, 5186.732, 5170.661, 5158.663, 5153.375, 5150.823, 5159.545, 
    5159.338, 5172.717, 5183.251, 5193.67, 5201.31, 5210.312, 5222.273, 
    5237.581,
  5189.047, 5166.959, 5150.313, 5139.151, 5133.023, 5132.198, 5135.335, 
    5149.923, 5159.583, 5172.228, 5185.868, 5196.082, 5207.686, 5219.961, 
    5235.046,
  5171.162, 5148.982, 5132.425, 5121.261, 5113.801, 5112.474, 5119.006, 
    5129.209, 5146.494, 5165.57, 5178.735, 5193.764, 5207.085, 5222.417, 
    5235.937,
  5154.929, 5134.455, 5118.322, 5108.142, 5101.486, 5099.076, 5104.09, 
    5121.984, 5141.314, 5159.208, 5177.362, 5193.65, 5210.54, 5226.248, 
    5239.161,
  5142.598, 5123.275, 5107.917, 5099.043, 5092.26, 5090.082, 5096.957, 
    5112.189, 5134.776, 5159.228, 5177.665, 5197.679, 5217.291, 5232.719, 
    5245.57,
  5134.191, 5116.488, 5102.655, 5094.751, 5089.499, 5088.377, 5096.137, 
    5117.465, 5141.123, 5162.803, 5183.714, 5206.846, 5225.352, 5240.569, 
    5254.452,
  5130.744, 5113.361, 5101.208, 5094.772, 5090.198, 5092.09, 5103.776, 
    5123.147, 5146.77, 5171.24, 5195.023, 5217.893, 5236.097, 5252.878, 
    5269.723,
  5287.585, 5266.829, 5248.687, 5230.771, 5216.297, 5204.552, 5196.761, 
    5193.228, 5192.77, 5193.437, 5197.703, 5203.401, 5209.928, 5217.183, 
    5228.666,
  5252.384, 5229.483, 5210.3, 5192.422, 5180.141, 5171.99, 5172.007, 
    5171.353, 5175.834, 5183.365, 5191.476, 5200.604, 5209.959, 5221.446, 
    5234.967,
  5215.838, 5192.309, 5173.029, 5158.5, 5150.204, 5151.279, 5148.457, 
    5160.692, 5167.522, 5177.444, 5187.982, 5199.33, 5211.187, 5223.694, 
    5240.842,
  5178.622, 5157.074, 5139.885, 5129.512, 5125.273, 5127.136, 5140.198, 
    5144.607, 5159.021, 5172.564, 5186.871, 5199.385, 5213.384, 5228.508, 
    5246.966,
  5148.264, 5129.918, 5117.253, 5110.398, 5109.526, 5115.888, 5124.687, 
    5143.886, 5157.554, 5170.399, 5186.408, 5200.537, 5215.602, 5230.702, 
    5250.546,
  5126.176, 5111.094, 5099.716, 5096.011, 5096.995, 5104.848, 5120.93, 
    5134.794, 5152.09, 5170.639, 5186.598, 5202.927, 5218.009, 5234.679, 
    5253.57,
  5111.087, 5099.042, 5090.271, 5088.493, 5092.778, 5101.707, 5115.15, 
    5136.638, 5155.225, 5171.062, 5188.873, 5205.126, 5220.414, 5236.318, 
    5255.452,
  5103.031, 5093.073, 5085.504, 5086.122, 5090.073, 5100.525, 5116.13, 
    5133.325, 5152.293, 5173.093, 5191.362, 5208.094, 5223.698, 5240.17, 
    5259.843,
  5100.715, 5092.488, 5087.339, 5088.65, 5094.392, 5104.269, 5118.643, 
    5139.802, 5159.743, 5177.533, 5195.377, 5212.328, 5227.994, 5245.292, 
    5264.9,
  5104.21, 5094.902, 5090.997, 5092.984, 5098.388, 5109.633, 5126.18, 
    5144.527, 5163.55, 5183.566, 5201.722, 5218.393, 5234.759, 5252.943, 
    5273.105,
  5309.006, 5289.173, 5270.894, 5253.311, 5239.026, 5227.052, 5217.771, 
    5212.668, 5209.453, 5207.238, 5208.696, 5214.011, 5223.412, 5235.891, 
    5251.498,
  5272.919, 5250.58, 5230.335, 5211.53, 5197.751, 5186.285, 5182.162, 
    5176.312, 5175.231, 5179.427, 5185.154, 5197.582, 5213.425, 5235.262, 
    5255.602,
  5237.296, 5214.599, 5194.46, 5180.026, 5167.15, 5165.054, 5154.007, 
    5159.743, 5158.715, 5165.433, 5174.961, 5192.354, 5214.169, 5239.083, 
    5263.406,
  5203.46, 5183.266, 5166.997, 5154.261, 5146.231, 5139.738, 5144.372, 
    5140.039, 5147.046, 5158.499, 5174.505, 5195.756, 5222.337, 5250.767, 
    5274.866,
  5178.228, 5160.986, 5146.534, 5136.394, 5131.288, 5129.449, 5130.158, 
    5139.756, 5152.217, 5161.748, 5182.643, 5206.722, 5236.109, 5262.538, 
    5288.084,
  5159.038, 5142.917, 5130.364, 5123.239, 5118.984, 5120.345, 5128.208, 
    5137.292, 5151.68, 5172.806, 5195.245, 5222.688, 5251.097, 5278.217, 
    5302.847,
  5144.494, 5131.855, 5121.995, 5116.931, 5115.949, 5120.125, 5130.072, 
    5148.781, 5167.413, 5187.624, 5211.974, 5239.478, 5266.484, 5293.74, 
    5318.078,
  5136.312, 5126.766, 5118.408, 5115.747, 5116.506, 5126.168, 5141.601, 
    5159.3, 5178.934, 5203.938, 5229.096, 5256.273, 5283.378, 5309.206, 
    5331.913,
  5134.539, 5127.827, 5121.777, 5122.035, 5127.485, 5139.944, 5156.823, 
    5177.023, 5198.699, 5221.249, 5246.299, 5272.776, 5298.465, 5322.784, 
    5342.68,
  5138.573, 5132.167, 5128.967, 5131.841, 5139.648, 5155.515, 5172.895, 
    5191.844, 5213.183, 5237.309, 5262.339, 5287.557, 5312.346, 5334.423, 
    5351.664,
  5384.3, 5360.994, 5338.706, 5313.687, 5291.472, 5270.933, 5253.62, 
    5242.823, 5234.172, 5227.582, 5226.032, 5227.863, 5234.183, 5245.438, 
    5260.401,
  5346.771, 5320.348, 5294.967, 5269.34, 5249.328, 5230.249, 5220.52, 
    5208.048, 5202.094, 5200, 5198.232, 5203.136, 5210.115, 5226.387, 5243.643,
  5305.859, 5279.559, 5254.201, 5234.654, 5214.278, 5205.932, 5186.41, 
    5186.698, 5177.803, 5178.378, 5179.456, 5185.99, 5196.395, 5213.486, 
    5236.349,
  5266.967, 5243.74, 5223.486, 5203.275, 5187.553, 5171.845, 5169.789, 
    5157.484, 5160.313, 5159.654, 5165.48, 5173.985, 5190.094, 5211.78, 
    5239.268,
  5238.415, 5218.819, 5198.215, 5180.302, 5165.344, 5154.945, 5146.251, 
    5148.425, 5147.109, 5151.247, 5159.773, 5172.552, 5194.481, 5220.011, 
    5251.254,
  5217.112, 5197.543, 5177.176, 5161.112, 5146.328, 5139.113, 5135.71, 
    5135.505, 5140.251, 5149.529, 5161.845, 5183.384, 5210.319, 5240.165, 
    5268.443,
  5199.503, 5182.104, 5162.872, 5149.279, 5138.54, 5133.293, 5131.569, 
    5137.914, 5145.379, 5159.151, 5180.437, 5207.423, 5235.863, 5263.587, 
    5289.132,
  5186.954, 5170.731, 5154.234, 5144.138, 5136.283, 5136.074, 5138.773, 
    5147.966, 5162.347, 5185.7, 5210.086, 5237.592, 5263.348, 5288.489, 
    5309.757,
  5179.715, 5167.229, 5156.332, 5151.461, 5149.444, 5151.986, 5159.449, 
    5174.899, 5195.667, 5218.002, 5242.678, 5267.469, 5291.129, 5311.742, 
    5328.487,
  5178.822, 5170.027, 5165.144, 5165.019, 5167.029, 5175.238, 5188.188, 
    5206.441, 5227.558, 5251.727, 5274.444, 5297.2, 5316.075, 5332.08, 
    5343.347,
  5474.637, 5461.804, 5445.409, 5421.892, 5394.461, 5361.68, 5326.402, 
    5298.247, 5271.093, 5248.6, 5235.162, 5229.26, 5228.868, 5231.91, 5237.285,
  5447.49, 5432.745, 5414.06, 5388.1, 5358.372, 5323.553, 5295.965, 5261.84, 
    5238.832, 5225.032, 5211.908, 5210.215, 5210.98, 5218.537, 5224.405,
  5421.681, 5406.626, 5383.939, 5358.043, 5323.728, 5299.894, 5255.244, 
    5240.078, 5210.805, 5199.013, 5190.922, 5192.706, 5195.635, 5203.811, 
    5213.439,
  5392.728, 5376.393, 5352.461, 5323.458, 5292.068, 5255.01, 5236.239, 
    5197.82, 5185.891, 5177.112, 5174.25, 5176.457, 5183.825, 5193.475, 
    5205.602,
  5361.596, 5345.132, 5320.314, 5292.755, 5260.305, 5231.168, 5197.442, 
    5187.198, 5168.871, 5159.746, 5161.974, 5165.372, 5175.424, 5185.902, 
    5201.771,
  5330.67, 5314.461, 5289.952, 5261.835, 5230.603, 5201.899, 5179.517, 
    5158.998, 5152.047, 5152.855, 5153.831, 5161.33, 5171.637, 5185.633, 
    5202.983,
  5303.781, 5288.127, 5262.71, 5236.976, 5208.732, 5184.032, 5164.412, 
    5155.877, 5150.39, 5148.992, 5154.154, 5163.423, 5175.304, 5191.886, 
    5212.307,
  5278.41, 5262.562, 5239.957, 5217.649, 5192.964, 5174.578, 5159.425, 
    5150.852, 5150.531, 5157.187, 5164.932, 5176.586, 5190.471, 5208.425, 
    5229.717,
  5256.57, 5244.238, 5227.986, 5211.17, 5193.869, 5179.997, 5172.261, 
    5172.371, 5175.797, 5181.613, 5190.878, 5202.268, 5215.356, 5231.937, 
    5252.188,
  5240.728, 5233.187, 5223.7, 5214.41, 5207.121, 5202.487, 5201.43, 5203.064, 
    5207.833, 5215.3, 5223.356, 5232.685, 5243.982, 5258.119, 5275.221,
  5385.678, 5394.238, 5405, 5413.973, 5422.636, 5426.488, 5426.658, 5425.574, 
    5418.598, 5403.975, 5387.628, 5367.057, 5345.285, 5325.028, 5309.861,
  5358.406, 5367.269, 5377.566, 5386.174, 5393.436, 5397.981, 5400.55, 
    5392.767, 5381.521, 5370.26, 5350.784, 5332.507, 5312.03, 5299.34, 
    5286.489,
  5335.752, 5345.492, 5355.052, 5365.656, 5371.385, 5378.241, 5366.771, 
    5368.037, 5348.271, 5331.793, 5312.778, 5295.468, 5278.328, 5267.194, 
    5262.961,
  5316.938, 5326.016, 5337.064, 5345.121, 5352.477, 5348.372, 5351.124, 
    5326.131, 5313.073, 5293.539, 5274.469, 5256.492, 5245.835, 5240.185, 
    5241.874,
  5301.464, 5311.081, 5322.125, 5329.995, 5333.278, 5331.806, 5315.25, 
    5306.434, 5281.101, 5250.77, 5238.413, 5221.553, 5217.737, 5216.622, 
    5226.146,
  5292.865, 5301.84, 5309.643, 5314.988, 5314.745, 5307.958, 5294.016, 
    5267.582, 5242.515, 5224.121, 5205.547, 5196.226, 5196.917, 5203.914, 
    5217.709,
  5288.194, 5296.08, 5301.859, 5304.368, 5301.853, 5290.89, 5270.261, 
    5248.936, 5223.606, 5197.774, 5184.484, 5182.534, 5187.766, 5199.766, 
    5218.294,
  5285.994, 5293.075, 5297.56, 5297.865, 5289.947, 5276.151, 5259.71, 
    5236.261, 5209.716, 5189.986, 5180.1, 5181.106, 5190.65, 5205.403, 
    5227.021,
  5287.085, 5294.159, 5296.054, 5291.977, 5283.35, 5276.071, 5262.407, 
    5244.109, 5218.292, 5194.629, 5185.674, 5188.096, 5198.148, 5215.323, 
    5239.834,
  5288.182, 5292.955, 5292.615, 5288.597, 5285.974, 5281.259, 5269.033, 
    5250.568, 5227.952, 5209.249, 5200.296, 5201.662, 5213.502, 5233.014, 
    5259.108,
  5386.936, 5361.53, 5341.679, 5327.037, 5318.035, 5312.896, 5310.941, 
    5313.696, 5317.432, 5321.788, 5328.091, 5336.528, 5345.527, 5356.077, 
    5367.639,
  5355.475, 5332.268, 5317.177, 5305.916, 5298.853, 5295.411, 5296.261, 
    5295.309, 5298.365, 5303.352, 5307.099, 5314.022, 5321.803, 5334.305, 
    5343.652,
  5331.721, 5314.661, 5303.702, 5295.858, 5290.12, 5289.607, 5285.508, 
    5288.785, 5286.969, 5288.105, 5291.642, 5297.098, 5303.642, 5312.667, 
    5324.982,
  5316.669, 5303.933, 5294.948, 5288.153, 5284.657, 5281.311, 5282.597, 
    5274.1, 5276.303, 5276.124, 5277.284, 5281.299, 5288.88, 5297.355, 
    5307.501,
  5307.157, 5297.756, 5291.316, 5286.663, 5281.322, 5277.916, 5270.633, 
    5267.02, 5258.518, 5255.02, 5258.159, 5261.637, 5269.87, 5278.012, 5290.27,
  5300.503, 5294.873, 5289.938, 5285.405, 5279.134, 5271.589, 5260.573, 
    5245.903, 5236.205, 5231.252, 5229.466, 5235.085, 5245.858, 5258.394, 
    5272.229,
  5297.806, 5295.771, 5291.819, 5285.497, 5275.853, 5262.287, 5245.13, 
    5227.379, 5209.206, 5197.67, 5197.397, 5205.446, 5218.663, 5236.327, 
    5254.938,
  5297.712, 5298.327, 5293.738, 5285.961, 5273.578, 5258.014, 5236.56, 
    5210.075, 5185.972, 5173.47, 5170.255, 5179.928, 5198.338, 5219.772, 
    5245.149,
  5302.017, 5303.169, 5297.337, 5287.583, 5274.206, 5255.549, 5230.953, 
    5203.528, 5179.966, 5168.086, 5166.589, 5174.345, 5191.645, 5217.007, 
    5245.904,
  5307.763, 5306.588, 5299.544, 5289.598, 5275.622, 5257.905, 5234.204, 
    5206.369, 5184.479, 5174.369, 5172.756, 5180.516, 5198.868, 5225.965, 
    5258.299,
  5479.059, 5471.021, 5463.071, 5448.407, 5432.143, 5413.135, 5393.068, 
    5375.271, 5355.886, 5334.06, 5316.902, 5303.662, 5294.542, 5289.6, 
    5290.786,
  5438.657, 5434.628, 5430.666, 5419.282, 5406.249, 5387.868, 5374.254, 
    5351.906, 5334.343, 5320.093, 5303.889, 5291.351, 5282.044, 5278.786, 
    5278.129,
  5398.179, 5399.556, 5397.786, 5391.953, 5379.821, 5370.537, 5347.214, 
    5339.759, 5318.329, 5300.69, 5287.047, 5278.915, 5272.829, 5270.516, 
    5270.292,
  5360.004, 5365.698, 5367.339, 5364.881, 5356.655, 5342.344, 5333.558, 
    5305.944, 5292.67, 5279.831, 5267.428, 5262.152, 5263.559, 5265.785, 
    5267.206,
  5340.5, 5345.826, 5347.297, 5344.76, 5336.521, 5325.409, 5304.856, 
    5296.101, 5272.492, 5250.786, 5245.178, 5245.826, 5258.634, 5263.687, 
    5268.719,
  5330.975, 5332.912, 5331.466, 5327.606, 5317.665, 5304.154, 5287.195, 
    5260.735, 5239.241, 5224.668, 5220.725, 5235.089, 5256.338, 5266.046, 
    5273.482,
  5323.754, 5323.821, 5320.544, 5313.549, 5302.989, 5286.319, 5266.58, 
    5245.438, 5222.072, 5200.782, 5205.165, 5231.915, 5256.688, 5271.319, 
    5281.58,
  5318.296, 5315.147, 5308.835, 5299.98, 5286.814, 5269.735, 5248.365, 
    5220.793, 5197.425, 5188.267, 5200.637, 5231.731, 5259.026, 5277.684, 
    5290.097,
  5308.401, 5305.621, 5299.917, 5290.413, 5276.253, 5256.297, 5232.729, 
    5209.198, 5191.869, 5185.639, 5204.176, 5236.571, 5264.884, 5284.749, 
    5299.509,
  5305.76, 5302.371, 5294.757, 5283.202, 5266.32, 5244.307, 5220.856, 
    5197.837, 5184.764, 5191.089, 5214.104, 5244.023, 5272.47, 5293.199, 
    5310.743,
  5362.576, 5337.509, 5318.756, 5305.106, 5300.518, 5302.663, 5313.227, 
    5331.871, 5352.422, 5368.3, 5378.917, 5379.694, 5372.52, 5359.038, 
    5343.454,
  5335.582, 5307.773, 5287.007, 5273.693, 5270.773, 5276.306, 5292.504, 
    5309.852, 5331.65, 5350.976, 5359.058, 5358.371, 5350.042, 5338.204, 
    5320.26,
  5320.191, 5289.967, 5270.112, 5258.859, 5257.144, 5267.487, 5277.131, 
    5302.458, 5320.612, 5334.373, 5340.029, 5337.926, 5328.057, 5313.625, 
    5299.011,
  5313.836, 5286.402, 5267.781, 5257.249, 5259.709, 5261.942, 5283.021, 
    5289.691, 5308.498, 5317.304, 5321.114, 5316.2, 5307.063, 5294.072, 
    5284.466,
  5314.515, 5292.521, 5276.912, 5269.37, 5267.266, 5274.849, 5277.805, 
    5290.587, 5299.013, 5299.026, 5303.798, 5295.686, 5288.41, 5280.583, 
    5277.522,
  5315.346, 5297.097, 5282.381, 5275.561, 5272.785, 5272.875, 5277.622, 
    5279.253, 5282.62, 5286.682, 5283.218, 5278.792, 5276.896, 5276.497, 
    5277.821,
  5313.384, 5298.85, 5286.37, 5277.839, 5272.919, 5272.375, 5271.199, 
    5272.743, 5273.283, 5269.801, 5267.831, 5269.711, 5272.857, 5278.48, 
    5286.002,
  5307.975, 5295.15, 5282.01, 5274.273, 5266.771, 5262.31, 5258.798, 
    5256.754, 5254.477, 5253.957, 5256.546, 5266.651, 5276.247, 5287.333, 
    5297.496,
  5302.019, 5290.731, 5278.442, 5268.885, 5260.093, 5253.836, 5247.884, 
    5246.326, 5242.884, 5243.715, 5255.675, 5272.182, 5285.714, 5299.102, 
    5310.236,
  5297.168, 5284.801, 5271.886, 5261.42, 5249.907, 5240.963, 5234.564, 
    5232.366, 5231.241, 5245.171, 5266.146, 5283.825, 5299.575, 5313.359, 
    5324.346,
  5514.575, 5473.435, 5435.478, 5396.912, 5363.134, 5329.664, 5295.004, 
    5267.668, 5248.63, 5237.238, 5240.592, 5254.625, 5272.016, 5285.569, 
    5298.152,
  5490.775, 5452.045, 5417.809, 5383.102, 5355.478, 5322.469, 5303.61, 
    5276.927, 5264.217, 5262.616, 5269.662, 5282.522, 5292.799, 5302.153, 
    5307.373,
  5467.877, 5433.286, 5401.578, 5373.948, 5347.674, 5329.402, 5305.121, 
    5295.233, 5289.869, 5290.892, 5296.945, 5304.79, 5310.388, 5311.755, 
    5310.01,
  5443.837, 5413.262, 5384.799, 5361.732, 5341.461, 5324.936, 5314.43, 
    5307.056, 5304.649, 5310.619, 5316.539, 5321.343, 5320.42, 5315.941, 
    5306.513,
  5421.105, 5392.693, 5369.666, 5350.363, 5336.487, 5326.688, 5317.075, 
    5315.323, 5321.021, 5324.158, 5329.185, 5331.187, 5326.684, 5315.439, 
    5302.851,
  5396.5, 5371.878, 5351.826, 5337.391, 5326.929, 5319.914, 5318.719, 
    5315.287, 5320.776, 5329.43, 5335.079, 5335.465, 5329.252, 5316.138, 
    5308.003,
  5373.479, 5352.707, 5333.198, 5323.012, 5316.844, 5314.469, 5314.375, 
    5319.038, 5323.619, 5331.387, 5336.248, 5338.481, 5329.688, 5320.302, 
    5318.297,
  5352.28, 5330.549, 5311.905, 5305.042, 5301.39, 5303.626, 5305.077, 
    5312.069, 5317.646, 5328.906, 5335.037, 5338.18, 5330.983, 5328.993, 
    5330.728,
  5332.022, 5308.016, 5289.998, 5283.803, 5284.795, 5291.028, 5295.999, 
    5305.155, 5314.359, 5324.635, 5332.663, 5334.752, 5335.329, 5339.655, 
    5342.173,
  5313.515, 5285.076, 5266.706, 5261.968, 5265.987, 5275.851, 5284.148, 
    5293.964, 5304.979, 5317.568, 5328.646, 5335.419, 5343.452, 5350.717, 
    5355.49,
  5613.039, 5586.1, 5555.892, 5519.273, 5484.822, 5449.135, 5417.746, 
    5395.184, 5381.773, 5369.491, 5356.932, 5331.802, 5307.542, 5288.726, 
    5276.276,
  5593.559, 5564.301, 5531.639, 5494.073, 5459.584, 5422.675, 5401.895, 
    5380.373, 5372.422, 5369.546, 5358.147, 5335.836, 5310.472, 5294.638, 
    5281.413,
  5572.927, 5540.702, 5505.724, 5469.623, 5432.939, 5412.351, 5377.433, 
    5373.022, 5367.359, 5370.544, 5359.209, 5339.812, 5315.451, 5298.926, 
    5285.479,
  5548.67, 5513.758, 5477.166, 5439.461, 5409.188, 5376.788, 5368.013, 
    5354.904, 5362.942, 5368.739, 5362.274, 5344.881, 5324.308, 5307.693, 
    5293.843,
  5522.342, 5485.946, 5448.071, 5413.866, 5382.429, 5360.783, 5346.438, 
    5351.762, 5364.812, 5368.619, 5364.969, 5351.655, 5334.96, 5319.934, 
    5306.434,
  5495.332, 5457.163, 5420.1, 5384.532, 5353.706, 5336.188, 5335.648, 
    5342.371, 5355.365, 5369.924, 5367.662, 5359.281, 5346.535, 5335.024, 
    5322.404,
  5468.865, 5433.178, 5393.964, 5359.35, 5331.47, 5323.044, 5327.333, 
    5344.094, 5360.3, 5370.855, 5372.185, 5366.994, 5358.172, 5349.083, 
    5338.519,
  5448.207, 5411.886, 5370.942, 5335.104, 5312.426, 5311.994, 5326.522, 
    5344.152, 5360.017, 5374.229, 5377.812, 5375.319, 5369.669, 5362.873, 
    5353.788,
  5431.905, 5396.607, 5354.936, 5322.458, 5306.971, 5313.149, 5332.038, 
    5351.484, 5368.048, 5380.505, 5384.781, 5384.636, 5381.169, 5375.781, 
    5367.563,
  5422.004, 5385.24, 5346.433, 5319.204, 5309.92, 5320.954, 5340.196, 
    5357.784, 5373.848, 5387.007, 5393.027, 5394.52, 5393.227, 5388.938, 
    5381.21,
  5616.679, 5587.196, 5557.678, 5520.15, 5480.566, 5437.066, 5397.127, 
    5367.821, 5353.668, 5344.96, 5334.973, 5321.39, 5308.903, 5302.354, 
    5298.731,
  5596.858, 5568.814, 5535.945, 5495.916, 5453.646, 5407.02, 5380.564, 
    5361.039, 5353.778, 5351.628, 5341.415, 5328.787, 5314.727, 5306.918, 
    5301.549,
  5578.498, 5549.083, 5514.515, 5473.597, 5428.292, 5399.504, 5363.83, 
    5364.561, 5361.564, 5360.945, 5350.242, 5339.446, 5324.773, 5313.418, 
    5304.245,
  5560.571, 5530.211, 5493.236, 5449.818, 5409.855, 5376.08, 5369.39, 
    5365.842, 5369.251, 5368.021, 5360.703, 5349.441, 5335.404, 5321.434, 
    5308.706,
  5543.623, 5511.546, 5473.753, 5433.213, 5397.692, 5378.192, 5371.794, 
    5377.469, 5382.284, 5376.528, 5370.516, 5357.995, 5344.701, 5328.246, 
    5313.348,
  5526.556, 5495.164, 5457.87, 5420.718, 5392.08, 5379.756, 5382.646, 
    5387.215, 5387.716, 5386.049, 5378.423, 5366.411, 5351.491, 5334.123, 
    5316.555,
  5511.99, 5481.775, 5446.788, 5417.399, 5398.289, 5394.416, 5395.716, 
    5400.663, 5400.764, 5395.8, 5386.583, 5373.975, 5357.312, 5338.996, 
    5318.626,
  5499.008, 5471.792, 5440.926, 5418.865, 5407.773, 5407.875, 5410.892, 
    5412.395, 5409.951, 5405.255, 5395.263, 5381.177, 5363.128, 5343.072, 
    5321.079,
  5489.453, 5466.182, 5439.704, 5426.326, 5423.171, 5424.098, 5424.725, 
    5424.957, 5422.304, 5415.311, 5403.964, 5388.309, 5368.766, 5347.245, 
    5323.813,
  5483.378, 5462.246, 5441.338, 5434.341, 5434.529, 5435.649, 5436.893, 
    5435.635, 5431.622, 5424.346, 5412.472, 5395.596, 5374.991, 5352.866, 
    5328.963,
  5589.954, 5562.534, 5535.387, 5503.277, 5470.018, 5444.811, 5431.008, 
    5421.411, 5409.024, 5390.622, 5371.287, 5350.359, 5330.02, 5309.993, 
    5294.739,
  5572.844, 5547.697, 5521.528, 5488.636, 5461.495, 5439.537, 5434.237, 
    5418.576, 5405.161, 5389.91, 5369.309, 5346.606, 5323.607, 5304.962, 
    5286.377,
  5558.862, 5533.607, 5509.257, 5479.892, 5454.984, 5445.904, 5429.774, 
    5424.104, 5407.877, 5388.543, 5365.509, 5341.701, 5316.879, 5295.55, 
    5276.694,
  5545.115, 5521.048, 5496.593, 5469.746, 5451.547, 5441.362, 5433.093, 
    5418.374, 5401.903, 5385.532, 5360.678, 5335.972, 5310.536, 5289.302, 
    5268.051,
  5531.379, 5509.062, 5485.407, 5462.406, 5451.979, 5442.297, 5430.753, 
    5421.007, 5405.67, 5380.274, 5357.34, 5330.372, 5306.211, 5281.904, 
    5260.846,
  5518.617, 5497.83, 5474.238, 5457.764, 5448.82, 5440.69, 5431.493, 
    5415.512, 5397.299, 5377.246, 5353.621, 5327.982, 5304.209, 5280.438, 
    5258.169,
  5506.193, 5487.507, 5466.248, 5454.631, 5449.745, 5441.711, 5430.804, 
    5417.791, 5399.43, 5375.627, 5352.455, 5329.276, 5305.95, 5283.386, 
    5260.877,
  5496.355, 5478.761, 5460.01, 5453.299, 5448.773, 5441.724, 5431.144, 
    5414.55, 5394.845, 5374.987, 5354.626, 5333.938, 5313.5, 5292.831, 
    5271.572,
  5489.084, 5472.99, 5457.398, 5453.772, 5450.76, 5443.352, 5431.83, 
    5416.654, 5397.756, 5377.492, 5358.945, 5341.828, 5324.673, 5306.525, 
    5287.753,
  5484.512, 5469.238, 5456.678, 5456.154, 5451.962, 5444.635, 5432.732, 
    5415.848, 5397.521, 5380.271, 5365.017, 5351.271, 5338.127, 5324.15, 5309,
  5566.935, 5534.088, 5501.464, 5470.969, 5446.318, 5425.045, 5408.752, 
    5397.098, 5384.746, 5367.338, 5351.1, 5334.15, 5318.195, 5300.707, 5286.8,
  5551.78, 5517.146, 5483.941, 5455.402, 5433.359, 5413.324, 5404.116, 
    5386.661, 5373.021, 5358.335, 5342.062, 5326.648, 5309.765, 5293.336, 
    5275.566,
  5537.731, 5501.604, 5469.695, 5445.307, 5424.248, 5413.166, 5394.086, 
    5386.449, 5367.823, 5351.049, 5336.302, 5322.708, 5305.504, 5286.792, 
    5267.379,
  5522.445, 5486.606, 5458.556, 5435.859, 5419.136, 5403.75, 5394.693, 
    5373.216, 5358.483, 5346.783, 5334.561, 5321.724, 5304.618, 5285.779, 
    5265.312,
  5508.695, 5475.45, 5451.062, 5431.745, 5418.01, 5404.208, 5385.854, 
    5374.489, 5357.473, 5343.904, 5335.035, 5321.979, 5306.259, 5286.861, 
    5268.087,
  5496.43, 5466.777, 5445.36, 5429.711, 5415.023, 5400.212, 5384.836, 
    5365.19, 5351.771, 5344.939, 5335.643, 5323.78, 5308.298, 5290.992, 
    5272.552,
  5487.138, 5461.989, 5442.95, 5429.63, 5415.91, 5400.044, 5381.989, 
    5367.857, 5354.972, 5344.847, 5335.782, 5324.005, 5308.945, 5293.121, 
    5276.329,
  5480.539, 5458.43, 5441.783, 5429.926, 5413.999, 5398.701, 5381.67, 
    5364.973, 5352.318, 5344.413, 5334.643, 5322.443, 5308.333, 5293.641, 
    5279.444,
  5476.89, 5458.104, 5443.169, 5431.218, 5416.296, 5400.265, 5382.726, 
    5368.563, 5355.029, 5343.08, 5331.689, 5318.905, 5304.974, 5291.422, 
    5279.872,
  5475.894, 5458.243, 5445.698, 5434.133, 5417.895, 5401.991, 5384.782, 
    5367.444, 5352.458, 5339.723, 5327.102, 5314.095, 5301.191, 5289.036, 
    5279.4,
  5569.098, 5531.782, 5494.471, 5462.472, 5441.341, 5421.383, 5400.716, 
    5384.721, 5368.502, 5351.862, 5345.648, 5344.216, 5341.725, 5335.788, 
    5327.692,
  5556.294, 5517.998, 5482.311, 5455.271, 5435.149, 5412.085, 5397.282, 
    5372.42, 5357.811, 5348.636, 5343.025, 5341.519, 5339.131, 5334.434, 
    5326.279,
  5545.083, 5507.402, 5473.926, 5452.106, 5429.163, 5412.386, 5383.464, 
    5374.123, 5353.201, 5341.999, 5337.609, 5336.081, 5333.672, 5330.256, 
    5323.121,
  5533.149, 5496.789, 5467.731, 5445.897, 5423.903, 5399.131, 5382.853, 
    5354.867, 5342.486, 5333.668, 5327.942, 5326.816, 5325.206, 5323.271, 
    5318.209,
  5523.092, 5488.958, 5464.705, 5442.521, 5420.097, 5396.122, 5370.287, 
    5354.833, 5334.663, 5320.202, 5316.169, 5313.302, 5313.496, 5311.874, 
    5310.008,
  5514.015, 5482.58, 5460.928, 5438.289, 5413.617, 5388.616, 5364.654, 
    5338.132, 5319.162, 5307.824, 5299.613, 5298.099, 5298.427, 5298.783, 
    5298.643,
  5507.223, 5479.926, 5459.391, 5436.201, 5411.757, 5384.253, 5356.245, 
    5332.537, 5310.514, 5293.335, 5284.96, 5282.128, 5282.208, 5283.866, 
    5285.089,
  5502.095, 5477.839, 5457.358, 5434.018, 5406.971, 5378.777, 5349.249, 
    5319.902, 5296.345, 5281.315, 5271.62, 5267.542, 5267.502, 5269.749, 
    5272.379,
  5499.949, 5479.095, 5458.456, 5434.757, 5408.078, 5377.019, 5344.99, 
    5316.301, 5291.151, 5272.539, 5262.416, 5257.217, 5254.961, 5256.248, 
    5259.687,
  5500.547, 5480.434, 5460.66, 5437.358, 5408.007, 5377.252, 5345.794, 
    5314.091, 5288.107, 5269.776, 5257.771, 5250.516, 5247.037, 5246.835, 
    5249.836,
  5543.875, 5510.218, 5479.23, 5451.689, 5427.705, 5403.568, 5378.557, 
    5360.312, 5344.108, 5328.703, 5322.453, 5321.354, 5325.769, 5331.902, 
    5334.466,
  5529.141, 5496.139, 5467.322, 5440.252, 5414.755, 5385.305, 5367.532, 
    5340.551, 5325.25, 5315.511, 5309.594, 5310.907, 5317.256, 5327.809, 
    5333.181,
  5517.105, 5486.245, 5459.437, 5433.03, 5403.141, 5381.354, 5345.759, 
    5334.666, 5312.501, 5299.741, 5294.448, 5298.208, 5306.213, 5320.713, 
    5330.299,
  5507.599, 5478.82, 5452.802, 5423.438, 5393.323, 5359.553, 5340.932, 
    5308.103, 5295.257, 5285.329, 5280.728, 5284.943, 5295.468, 5312.937, 
    5327.064,
  5501.166, 5475.378, 5449.755, 5418.761, 5386.269, 5354.071, 5319.608, 
    5303.815, 5284.367, 5269.311, 5266.804, 5271.246, 5284.382, 5303.308, 
    5322.979,
  5497.545, 5473.678, 5446.952, 5414.712, 5378.128, 5342.214, 5310.681, 
    5282.099, 5265.924, 5259.12, 5255.888, 5262.05, 5275.012, 5296.488, 
    5318.125,
  5496.735, 5475.127, 5448.339, 5415.443, 5378.255, 5337.745, 5299.923, 
    5276.308, 5260.981, 5250.21, 5249.165, 5255.75, 5267.804, 5290.396, 
    5314.145,
  5498.084, 5478.28, 5451.298, 5417.752, 5377.036, 5335.003, 5295.647, 
    5265.754, 5250.913, 5246.398, 5245.743, 5253.335, 5265.067, 5287.679, 
    5311.702,
  5501.57, 5483.902, 5458.106, 5426.708, 5387.624, 5342.314, 5298.13, 
    5268.531, 5252.018, 5245.715, 5244.142, 5252.299, 5264.643, 5287.032, 
    5311.613,
  5506.872, 5490.484, 5468.717, 5438.228, 5397.816, 5354.323, 5309.188, 
    5272.83, 5253.589, 5248.045, 5247.619, 5254.287, 5268.391, 5289.766, 
    5313.011,
  5462.864, 5446.002, 5429.719, 5407.245, 5379.789, 5350.747, 5321.835, 
    5302.299, 5292.426, 5290.683, 5296.401, 5307.507, 5320.896, 5337.447, 
    5353.432,
  5455.841, 5439.582, 5419.543, 5391.028, 5357.647, 5320.584, 5296.778, 
    5274.263, 5269.115, 5273.834, 5284.415, 5300.073, 5317.153, 5338.743, 
    5358.036,
  5451.818, 5434.231, 5409.217, 5375.63, 5334.752, 5305.42, 5265.491, 
    5257.553, 5251.96, 5261.542, 5274.986, 5294.522, 5315.296, 5338.702, 
    5360.584,
  5448.095, 5428.365, 5398.725, 5358.681, 5316.726, 5276.234, 5255.343, 
    5234.726, 5240.524, 5252.559, 5271.027, 5290.682, 5314.907, 5341.117, 
    5365.891,
  5445.759, 5423.615, 5390.148, 5346.739, 5304.192, 5266.782, 5237.457, 
    5230.122, 5237.947, 5249.859, 5269.185, 5290.231, 5316.689, 5342.674, 
    5370.325,
  5443.533, 5420.027, 5383.12, 5339.253, 5295.574, 5259.844, 5235.618, 
    5228.306, 5235.204, 5253.533, 5270.187, 5293.059, 5319.226, 5348.14, 
    5374.44,
  5442.681, 5419.03, 5380.662, 5338.072, 5297.517, 5264.669, 5242.412, 
    5238.251, 5247.7, 5259.187, 5275.459, 5298.797, 5324.828, 5353.347, 
    5379.148,
  5443.128, 5419.375, 5381.679, 5341.208, 5302.69, 5273.228, 5255.933, 
    5250.928, 5255.495, 5268.088, 5284.141, 5306.702, 5332.758, 5360.512, 
    5385.054,
  5445.396, 5422.968, 5387.361, 5350.238, 5316.257, 5288.988, 5271.681, 
    5268.093, 5271.641, 5280.989, 5295.722, 5319.079, 5342.988, 5368.745, 
    5390.485,
  5448.779, 5427.535, 5395.819, 5362.99, 5330.507, 5306.112, 5290.969, 
    5284.37, 5286.35, 5296.261, 5311.805, 5332.865, 5354.774, 5377.583, 
    5396.216,
  5452.634, 5426.56, 5400.36, 5371.704, 5342.372, 5314.523, 5292.417, 
    5280.141, 5278.935, 5287.796, 5304.759, 5328.945, 5350.547, 5375.26, 
    5401.013,
  5436.967, 5409.988, 5381.588, 5349.48, 5317.14, 5286.533, 5270.658, 
    5257.717, 5257.46, 5271.62, 5293.427, 5322.344, 5349.25, 5381.481, 5407.55,
  5422.065, 5394.865, 5363.928, 5330.173, 5295.805, 5275.447, 5248.16, 
    5244.768, 5247.372, 5264.573, 5290.052, 5321.814, 5354.564, 5386.842, 
    5415.243,
  5408.03, 5379.545, 5346.617, 5311.264, 5280.702, 5254.026, 5244.352, 
    5232.631, 5241.438, 5264.121, 5294.314, 5327.207, 5363.687, 5398.761, 
    5426.075,
  5394.652, 5365.938, 5332.286, 5298.492, 5271.932, 5250.887, 5237.729, 
    5236.084, 5255.165, 5270.898, 5304.958, 5338.556, 5376.668, 5408.561, 
    5436.705,
  5382.98, 5353.888, 5320.089, 5290.627, 5266.489, 5250.088, 5242.844, 
    5246.053, 5257.738, 5287.232, 5318.782, 5354.88, 5390.883, 5423.246, 
    5448.279,
  5373.317, 5345.102, 5313.621, 5288.756, 5269.357, 5258.274, 5252.759, 
    5260.692, 5281.391, 5305.765, 5337.153, 5372.398, 5405.396, 5435.849, 
    5460.396,
  5366.753, 5339.706, 5311.444, 5290.708, 5274.772, 5267.979, 5268.747, 
    5278.224, 5296.77, 5324.484, 5356.816, 5388.656, 5420.334, 5448.572, 
    5473.768,
  5363.697, 5339.17, 5315.688, 5297.988, 5286.855, 5283.514, 5286.47, 
    5300.473, 5321.414, 5346.015, 5374.425, 5404.183, 5433.536, 5460.974, 
    5486.356,
  5364.663, 5342.596, 5323.053, 5308.528, 5299.791, 5299.248, 5305.901, 
    5318.669, 5337.672, 5362.91, 5390.504, 5418.224, 5446.186, 5473.045, 
    5498.513,
  5467.982, 5458.217, 5446.27, 5429.66, 5412.243, 5392.479, 5369.712, 
    5351.455, 5336.636, 5328.864, 5329.928, 5344.714, 5369.011, 5393.77, 
    5413.461,
  5450.536, 5438.287, 5422.533, 5404.595, 5384.221, 5359.787, 5340.349, 
    5321.404, 5306.559, 5306.299, 5313.825, 5337.179, 5366.596, 5397.502, 
    5417.8,
  5432.166, 5417.253, 5398.42, 5379.806, 5352.643, 5338.311, 5305.169, 
    5297.754, 5286.357, 5291.249, 5305.438, 5336.286, 5371.056, 5400.516, 
    5423.482,
  5412.419, 5393.195, 5373.234, 5348.305, 5326.33, 5298.564, 5290.722, 
    5270.732, 5271.884, 5282.432, 5307.261, 5342.584, 5380.104, 5409.64, 
    5433.459,
  5388.092, 5368.463, 5345.876, 5322.24, 5298.398, 5280.286, 5265.442, 
    5265.487, 5273.406, 5285.489, 5317.813, 5355.512, 5392.335, 5420.509, 
    5445.206,
  5364.258, 5343.751, 5320.465, 5297.185, 5276.437, 5262.768, 5257.731, 
    5260.602, 5271.533, 5298.972, 5334.759, 5372.899, 5407.189, 5435.82, 
    5458.134,
  5342.065, 5323.836, 5300.023, 5280.757, 5264.965, 5257.589, 5256.686, 
    5269.468, 5289.742, 5320.294, 5357.45, 5392.609, 5425.086, 5450.456, 
    5471.601,
  5326.958, 5307.55, 5286.7, 5272.575, 5262.255, 5262.139, 5269.474, 
    5285.714, 5310.786, 5346.818, 5381.799, 5414.549, 5443.154, 5466.078, 
    5486.237,
  5315.792, 5299.74, 5285.566, 5277.222, 5274.454, 5279.148, 5291.121, 
    5314.803, 5344.341, 5376.928, 5407.352, 5436.311, 5460.021, 5481.049, 
    5499.516,
  5313.879, 5300.967, 5293.058, 5290.149, 5292.983, 5304.044, 5323.155, 
    5347.14, 5375.208, 5405.026, 5431.868, 5455.851, 5476.896, 5496.87, 
    5514.28,
  5448.405, 5463.053, 5476.646, 5484.226, 5488.5, 5488.583, 5484.237, 
    5478.823, 5467.724, 5452.21, 5434.208, 5416.461, 5401.555, 5399.384, 
    5409.712,
  5444.398, 5456.942, 5465.997, 5471.131, 5472.476, 5469.891, 5466.438, 
    5454.387, 5442.743, 5429.269, 5411.141, 5394.283, 5387.606, 5398.192, 
    5411.836,
  5438.787, 5447.921, 5452.864, 5456.371, 5453.234, 5452.924, 5437.973, 
    5436.06, 5419.254, 5405.379, 5389.017, 5380.536, 5387.304, 5402.712, 
    5417.416,
  5429.539, 5433.55, 5435.526, 5433.506, 5431.206, 5421.472, 5420.64, 
    5400.576, 5393.021, 5382.847, 5374.791, 5378.263, 5395.937, 5412.302, 
    5427.601,
  5415.954, 5415.698, 5413.373, 5409.595, 5403.024, 5396.85, 5384.293, 
    5384.602, 5374.105, 5365.889, 5370.67, 5386.781, 5408.359, 5422.487, 
    5436.302,
  5393.22, 5389.254, 5382.875, 5376.799, 5368.35, 5362.407, 5357.314, 
    5351.313, 5351.939, 5360.062, 5376.498, 5400.822, 5419.92, 5436.918, 
    5449.748,
  5366.495, 5360.835, 5352.025, 5344.662, 5337.412, 5333.297, 5330.944, 
    5337.931, 5345.31, 5363.061, 5390.601, 5415.578, 5436.859, 5453.693, 
    5467.223,
  5338.708, 5330.479, 5319.347, 5312.1, 5306.72, 5307.657, 5313.269, 
    5322.872, 5344.019, 5377.292, 5408.208, 5434.605, 5456.359, 5472.644, 
    5487.145,
  5312.332, 5302.71, 5293.9, 5289.334, 5288.986, 5294.065, 5306.113, 
    5329.141, 5362.744, 5398.563, 5429.042, 5456.602, 5476.363, 5494.849, 
    5508.987,
  5293.047, 5284.34, 5278.674, 5276.888, 5280.872, 5292.967, 5314.293, 
    5347.364, 5386.815, 5422.751, 5453.19, 5478.375, 5499.184, 5516.495, 
    5530.795,
  5426.039, 5444.271, 5465.355, 5487.668, 5508.745, 5527.082, 5542.301, 
    5555.428, 5561.288, 5558.271, 5543.837, 5522.126, 5494.911, 5466.087, 
    5458.174,
  5417.563, 5438.173, 5460.161, 5483.686, 5504.047, 5522.32, 5538.472, 
    5548.037, 5551.418, 5546.594, 5530.68, 5504.863, 5472.801, 5453.852, 
    5447.3,
  5412.338, 5434.78, 5457.713, 5480.502, 5501.228, 5522.348, 5532.951, 
    5542.91, 5545.255, 5533.398, 5516.665, 5488.378, 5461.317, 5450.912, 
    5447.005,
  5410.537, 5432.18, 5455.644, 5476.368, 5499.414, 5514.665, 5531.41, 
    5532.757, 5531.857, 5521.915, 5502.659, 5476.923, 5464.714, 5458.271, 
    5458.533,
  5411.238, 5431.782, 5454.342, 5474.802, 5494.493, 5515.264, 5522.919, 
    5530.369, 5524.745, 5508.594, 5490.749, 5471.404, 5472.107, 5467.519, 
    5472.194,
  5413.628, 5431.333, 5450.78, 5469.796, 5488.421, 5505.125, 5516.342, 
    5517.707, 5510.334, 5498.258, 5479.837, 5473.161, 5478.385, 5478.804, 
    5483.636,
  5415.488, 5431.167, 5448.604, 5463.831, 5481.9, 5498.556, 5505.715, 
    5508.34, 5501.26, 5485.726, 5474.523, 5477.934, 5482.488, 5486.306, 
    5491.314,
  5414.194, 5428.349, 5441.529, 5455.505, 5470.954, 5486.321, 5494.721, 
    5495.44, 5487.4, 5477.286, 5474.996, 5482.298, 5486.966, 5492.462, 
    5497.805,
  5406.945, 5419.844, 5432.717, 5446.73, 5462.473, 5475.858, 5483.424, 
    5486.031, 5479.296, 5475.92, 5480.731, 5487.184, 5491.672, 5497.616, 
    5504.868,
  5392.877, 5405.096, 5417.356, 5432.644, 5448.59, 5463.668, 5472.472, 
    5475.958, 5475.745, 5481.614, 5489.227, 5494.706, 5500.825, 5507.911, 
    5515.81,
  5406.937, 5414.755, 5430.234, 5453.36, 5477.201, 5500.03, 5523.39, 
    5545.124, 5563.402, 5577.545, 5587.421, 5593.408, 5592.476, 5588.115, 
    5582.315,
  5407.522, 5416.307, 5433.146, 5456.132, 5476.417, 5499.469, 5521.476, 
    5541.873, 5556.807, 5571.01, 5577.521, 5580.235, 5575.106, 5569.204, 
    5558.396,
  5411.984, 5425.224, 5442.443, 5463.228, 5481.565, 5506.56, 5521.435, 
    5539.869, 5553.295, 5562.246, 5567.277, 5565.776, 5557.449, 5546.456, 
    5534.723,
  5421.51, 5434.938, 5452.297, 5468.918, 5490.574, 5503.373, 5526.262, 
    5534.413, 5547.847, 5554.619, 5555.625, 5549.54, 5539.799, 5527.684, 
    5514.284,
  5430.26, 5444.966, 5461.868, 5479.308, 5494.075, 5512.994, 5521.897, 
    5536.763, 5543.647, 5545.458, 5543.564, 5533.87, 5523.672, 5510.185, 
    5497.047,
  5437.338, 5453.265, 5468.518, 5484.374, 5497.305, 5509.458, 5525.514, 
    5533.489, 5538.698, 5537.493, 5529.508, 5518.094, 5509.775, 5498.426, 
    5485.908,
  5444.113, 5460.118, 5474.897, 5487.776, 5500.345, 5514.108, 5524.366, 
    5533.064, 5533.416, 5525.47, 5515.288, 5506.157, 5499.656, 5491.306, 
    5481.346,
  5450.305, 5465.893, 5479.207, 5490.668, 5502.305, 5515.465, 5528.034, 
    5530.2, 5524.591, 5512.957, 5502.979, 5498.655, 5495.773, 5490.653, 
    5484.289,
  5456.899, 5471.999, 5483.923, 5495.346, 5508.687, 5521.45, 5529.043, 
    5527.441, 5516.12, 5505.009, 5499.459, 5498.402, 5495.781, 5493.832, 
    5492.526,
  5464.248, 5476.688, 5487.612, 5499.297, 5513.114, 5526.767, 5532.445, 
    5526.155, 5513.951, 5506.66, 5502.715, 5500.561, 5500.028, 5499.914, 
    5500.975,
  5361.019, 5380.636, 5397.504, 5422.181, 5444.334, 5461.445, 5482.102, 
    5506.573, 5534.5, 5559.386, 5580.388, 5600.555, 5615.636, 5628.015, 
    5637.084,
  5361.899, 5378.096, 5394.929, 5418.898, 5439.244, 5459.111, 5478.438, 
    5499.843, 5524.028, 5550.961, 5570.714, 5588.715, 5602.304, 5614.591, 
    5620.863,
  5362.049, 5377.855, 5395.852, 5418.975, 5439.074, 5460.927, 5474.962, 
    5498.088, 5520.22, 5543.193, 5561.98, 5577.345, 5589.575, 5597.814, 
    5604.367,
  5369.667, 5382.869, 5401.273, 5420.927, 5442.233, 5456.986, 5480.825, 
    5492.414, 5514.264, 5534.634, 5553.298, 5566.314, 5576.529, 5583.267, 
    5586.738,
  5385.372, 5396.239, 5412.023, 5430.419, 5446.973, 5466.287, 5476.57, 
    5496.991, 5513.567, 5525.656, 5542.702, 5553.498, 5561.604, 5564.601, 
    5567.368,
  5409.9, 5417.638, 5427.923, 5442.412, 5455.202, 5468.043, 5484.326, 
    5494.769, 5506.602, 5522.364, 5531.232, 5540.575, 5546.306, 5547.453, 
    5546.902,
  5436.089, 5440.993, 5447.406, 5456.773, 5467.637, 5478.028, 5486.992, 
    5500.36, 5509.726, 5514.094, 5519.958, 5524.359, 5526.591, 5525.616, 
    5523.106,
  5457.675, 5460.219, 5464.004, 5470.164, 5476.723, 5485.334, 5493.271, 
    5496.785, 5499.881, 5503.989, 5505.539, 5506.715, 5506.958, 5506.497, 
    5503.699,
  5473.621, 5475.062, 5477.754, 5482.192, 5487.808, 5491.717, 5493.39, 
    5494.915, 5494.417, 5492.69, 5492.421, 5493.207, 5492.792, 5492.34, 
    5491.064,
  5485.208, 5486.519, 5489.419, 5493.212, 5496.323, 5498.69, 5497.949, 
    5494.694, 5490.99, 5490.277, 5490.172, 5489.08, 5487.706, 5487.112, 
    5486.777,
  5361.836, 5362.96, 5366.846, 5368.917, 5377.577, 5391.655, 5424.848, 
    5471.535, 5510.427, 5546.751, 5578.216, 5609.381, 5633.59, 5654.314, 
    5668.46,
  5371.448, 5372.174, 5369.06, 5373.499, 5377.172, 5387.747, 5419.227, 
    5465.429, 5504.069, 5544.107, 5576.463, 5606.23, 5629.959, 5649.714, 
    5662.099,
  5383.583, 5381.027, 5379.615, 5381.646, 5382.286, 5395.158, 5420.1, 
    5468.838, 5506.965, 5541.442, 5572.886, 5601.182, 5623.907, 5641.063, 
    5654.015,
  5402.757, 5399.226, 5396.456, 5394.857, 5398.175, 5398.695, 5433.525, 
    5465.219, 5503.318, 5539.159, 5567.983, 5593.786, 5615.83, 5632.638, 
    5643.375,
  5421.129, 5419.57, 5416.997, 5416.635, 5415.098, 5423.804, 5436.781, 
    5482.153, 5511.8, 5536.358, 5562.772, 5586.08, 5606.183, 5620.687, 
    5630.872,
  5437.405, 5437.588, 5435.81, 5434.973, 5435.447, 5437.663, 5457.307, 
    5480.312, 5503.351, 5535.11, 5555.523, 5578.274, 5594.77, 5608.288, 
    5615.958,
  5448.107, 5447.899, 5447.663, 5446.982, 5449.766, 5455, 5465.208, 5490.287, 
    5511.846, 5529.86, 5549.479, 5568.142, 5582.272, 5593.646, 5598.979,
  5456.977, 5456.002, 5455.486, 5456.673, 5458.646, 5465.314, 5476.094, 
    5488.084, 5502.713, 5523.695, 5541.171, 5556.033, 5569.295, 5578.255, 
    5582.762,
  5467.206, 5465.667, 5464.936, 5465.4, 5469.105, 5473.703, 5481.726, 
    5494.764, 5508.9, 5520.347, 5532.509, 5544.486, 5554.297, 5561.051, 
    5564.711,
  5478.273, 5474.992, 5473.703, 5473.382, 5474.646, 5478.656, 5484.949, 
    5490.954, 5499.979, 5511.528, 5522.104, 5530.709, 5538.701, 5543.931, 
    5546.688,
  5412.146, 5403.84, 5396.208, 5393.956, 5396.852, 5408.846, 5427.097, 
    5451.517, 5476.692, 5501.026, 5529.867, 5559.441, 5589.355, 5617.569, 
    5643.765,
  5410.001, 5399.517, 5389.437, 5385.593, 5384.546, 5395.87, 5414.981, 
    5437.572, 5463.785, 5495.922, 5528.971, 5560.798, 5592.051, 5622.405, 
    5647.263,
  5406.566, 5393.266, 5381.484, 5375.012, 5374.31, 5385.538, 5400.782, 
    5433.563, 5463.712, 5493.247, 5529.104, 5562.413, 5596.394, 5623.305, 
    5649.188,
  5399.403, 5384.528, 5370.56, 5360.728, 5358.308, 5366.289, 5395.825, 
    5416.807, 5453.149, 5490.244, 5530.741, 5564.482, 5600.159, 5627.825, 
    5651.361,
  5392.874, 5376.389, 5358.106, 5345.046, 5338.695, 5355.953, 5374.368, 
    5422.259, 5459.748, 5490.8, 5532.561, 5567.611, 5602.748, 5627.922, 
    5650.001,
  5388.642, 5369.047, 5345.142, 5324.691, 5318.634, 5336.52, 5374.274, 
    5409.354, 5449.338, 5495.811, 5534.732, 5572.231, 5603.802, 5629.387, 
    5648.449,
  5387.554, 5365.484, 5336.482, 5312.609, 5310.618, 5334.553, 5369.424, 
    5422.621, 5465.873, 5499.167, 5540.781, 5574.603, 5604.473, 5626.705, 
    5643.685,
  5392.349, 5369.982, 5341.478, 5321.411, 5319.843, 5346.5, 5384.313, 
    5423.703, 5462.23, 5506.031, 5544.531, 5575.938, 5603.839, 5623.532, 
    5638.035,
  5402.519, 5383.988, 5361.854, 5347.399, 5350.079, 5371.344, 5404.827, 
    5446.755, 5482.254, 5514.897, 5547.699, 5576.866, 5600.322, 5617.13, 
    5628.753,
  5417.17, 5403.766, 5389.383, 5380.603, 5382.771, 5402.051, 5428.114, 
    5456.324, 5485.736, 5519.447, 5550.626, 5575.474, 5595.682, 5609.678, 
    5618.475,
  5452.635, 5446.671, 5441.157, 5435.812, 5431.708, 5427.032, 5424.797, 
    5428.084, 5433.674, 5438.922, 5448.679, 5463.88, 5482.802, 5509.118, 
    5541.27,
  5434.813, 5427.14, 5420.651, 5415.624, 5413.446, 5412.555, 5413.357, 
    5414.546, 5421.801, 5432.445, 5443.509, 5461.111, 5481.518, 5509.593, 
    5540.54,
  5416.41, 5406.679, 5399.704, 5396.129, 5396.068, 5399.601, 5399.786, 
    5408.212, 5417.622, 5428.177, 5441.57, 5462.215, 5486.464, 5512.646, 
    5545.29,
  5397.676, 5385.52, 5377.192, 5373.303, 5377.287, 5382.579, 5393.827, 
    5394.607, 5408.534, 5424.815, 5442.77, 5466.454, 5492.489, 5522.408, 
    5554.297,
  5380.34, 5364.089, 5352.789, 5350.279, 5356.728, 5368.905, 5379.203, 
    5394.36, 5409.04, 5424.896, 5446.469, 5473.128, 5501.538, 5530.487, 
    5562.752,
  5362.155, 5339.356, 5319.648, 5316.632, 5331.21, 5351.679, 5372.124, 
    5384.479, 5402.14, 5428.185, 5451.812, 5481.657, 5510.186, 5542.589, 
    5572.542,
  5346.576, 5316.23, 5290.591, 5286.402, 5306.577, 5338.107, 5362.252, 
    5386.007, 5409.036, 5432.257, 5460.513, 5490.459, 5520.021, 5552.283, 
    5581.746,
  5340.014, 5306.636, 5279.729, 5275.145, 5297.396, 5333.125, 5361.697, 
    5382.445, 5408.003, 5440.102, 5469.612, 5500.195, 5531.054, 5563.757, 
    5591.463,
  5344.358, 5315.37, 5293.156, 5289.907, 5312.425, 5341.143, 5366.576, 
    5392.772, 5420.913, 5449.808, 5479.16, 5511.004, 5542.174, 5573.532, 
    5599.164,
  5359.032, 5336.87, 5321.943, 5320.689, 5335.076, 5355.729, 5377.85, 
    5399.563, 5427.497, 5458.517, 5489.846, 5521.851, 5553.228, 5582.393, 
    5606.17,
  5492.014, 5486.07, 5481.481, 5475.573, 5471.494, 5466.345, 5461.291, 
    5458.947, 5455.503, 5451.255, 5449.902, 5449.803, 5451.177, 5454.226, 
    5468.586,
  5468.798, 5462.3, 5456.706, 5450.757, 5445.871, 5442.185, 5441.823, 
    5437.242, 5436.445, 5437.05, 5435.686, 5438.497, 5441.986, 5448.349, 
    5462.79,
  5445.734, 5438.489, 5430.8, 5425.213, 5420.219, 5420.604, 5414.96, 
    5422.909, 5418.992, 5421.204, 5423.257, 5427.663, 5433.767, 5441.671, 
    5460.065,
  5423.504, 5413.83, 5404.55, 5396.788, 5393.001, 5391.761, 5400.256, 
    5396.392, 5405.384, 5407.467, 5413.102, 5419.262, 5428.314, 5440.243, 
    5463.138,
  5401.711, 5388.404, 5375.173, 5365.734, 5362.171, 5366.162, 5370.361, 
    5386.617, 5388.779, 5396.795, 5405.643, 5414.502, 5426.699, 5442.93, 
    5471.03,
  5380.753, 5363.344, 5345.722, 5332.588, 5328.523, 5337.69, 5353.074, 
    5364.518, 5378.609, 5391.281, 5401.823, 5415.548, 5430.328, 5453.854, 
    5483.422,
  5363.528, 5342.759, 5319.074, 5302.151, 5299.964, 5312.61, 5334.167, 
    5357.848, 5373.748, 5388.695, 5404.568, 5421.157, 5439.874, 5468.767, 
    5501.84,
  5352.317, 5329.472, 5302.008, 5283.924, 5283.695, 5302.951, 5329.85, 
    5352.272, 5373.76, 5393.848, 5412.934, 5430.892, 5456.479, 5488.96, 
    5521.901,
  5349.738, 5330.056, 5304.96, 5291.606, 5296.03, 5314.833, 5338.458, 
    5362.326, 5384.327, 5404.347, 5424.722, 5447.359, 5478.646, 5511.894, 
    5540.952,
  5355.122, 5341.597, 5325.729, 5317.181, 5321.208, 5335.26, 5354.5, 
    5374.928, 5398.105, 5420.735, 5442.036, 5469.926, 5502.75, 5533.768, 
    5561.142,
  5495.188, 5508.374, 5521.623, 5531.501, 5540.712, 5545.746, 5548.486, 
    5550.325, 5547.07, 5539.999, 5532.076, 5520.872, 5508.052, 5492.939, 
    5477.792,
  5483.209, 5492.945, 5502.664, 5511.696, 5517.979, 5523.907, 5527.602, 
    5526.561, 5526.091, 5525.08, 5517.184, 5509.955, 5499.499, 5489.692, 
    5474.432,
  5473.873, 5479.521, 5485.576, 5492.95, 5496.763, 5503.813, 5500.521, 
    5509.393, 5505.051, 5505.167, 5502.887, 5499.771, 5494.442, 5489.256, 
    5478.58,
  5460.929, 5464.018, 5466.448, 5468.872, 5472.27, 5472.822, 5482.261, 
    5475.273, 5486.287, 5486.859, 5489.447, 5490.474, 5492.022, 5490.813, 
    5487.254,
  5440.45, 5443.042, 5443.297, 5443.729, 5444.4, 5446.567, 5445.553, 
    5459.583, 5459.387, 5467.548, 5476.03, 5483.438, 5490.729, 5493.925, 
    5497.29,
  5420.557, 5419.532, 5417.017, 5414.825, 5411.055, 5411.992, 5416.811, 
    5421.477, 5437.323, 5452.604, 5463.913, 5478.811, 5490.835, 5499.956, 
    5506.917,
  5400.792, 5397.99, 5392.637, 5386.662, 5381.173, 5378.602, 5382.539, 
    5398.544, 5415.224, 5434.865, 5455.835, 5475.978, 5493.468, 5507.049, 
    5518.202,
  5385.817, 5381.149, 5373.277, 5364.375, 5354.423, 5350.833, 5354.395, 
    5368.67, 5394.004, 5424.755, 5449.791, 5475.423, 5498.514, 5516.267, 
    5529.236,
  5375.952, 5371.971, 5362.349, 5351.746, 5341.884, 5335.584, 5337.733, 
    5355.98, 5383.706, 5416.404, 5447.791, 5479.146, 5505.311, 5526.955, 
    5539.274,
  5374.031, 5368.532, 5359.068, 5349.349, 5338.916, 5332.304, 5332.82, 
    5348.638, 5379.098, 5416.776, 5452.47, 5486.277, 5516.598, 5538.865, 
    5549.656,
  5446.109, 5445.508, 5452.254, 5460.607, 5467.627, 5485.546, 5506.056, 
    5522.703, 5538.79, 5552.389, 5563.392, 5568.724, 5565.35, 5551.586, 
    5537.022,
  5449.068, 5447.619, 5455.409, 5465.531, 5472.492, 5488.425, 5504.127, 
    5518.568, 5533.942, 5549.296, 5559.642, 5563.379, 5557.123, 5544.998, 
    5530.363,
  5453.736, 5451.877, 5460.308, 5470.827, 5478.489, 5494.12, 5503.646, 
    5519.705, 5533.257, 5546.231, 5556.146, 5557.104, 5548.754, 5535.28, 
    5524.922,
  5457.645, 5457.201, 5465.375, 5472.814, 5485.377, 5491.574, 5509.578, 
    5517.119, 5533.453, 5544.446, 5551.5, 5548.484, 5540.146, 5529.465, 
    5520.918,
  5457.993, 5462.552, 5469.646, 5477.692, 5485.343, 5499.435, 5505.185, 
    5521.438, 5531.165, 5538.6, 5544.091, 5538.928, 5531.911, 5522.396, 
    5517.036,
  5451.312, 5462.084, 5470.415, 5477.924, 5485.941, 5493.935, 5508.793, 
    5515.587, 5525.393, 5533.729, 5534.296, 5529.813, 5524.195, 5518.69, 
    5514.457,
  5444.203, 5455.52, 5468.015, 5475.399, 5483.385, 5493.616, 5501.473, 
    5513.874, 5520.54, 5523.324, 5523.311, 5520.897, 5517.788, 5515.198, 
    5511.337,
  5431.915, 5442.558, 5457.662, 5469.002, 5475.039, 5486.028, 5495.098, 
    5502.007, 5507.255, 5512.354, 5512, 5512.165, 5513.017, 5514.112, 5509.816,
  5419.229, 5429.28, 5444.317, 5457.226, 5464.915, 5475.253, 5483.393, 
    5492.262, 5496.658, 5499.433, 5502.014, 5506.749, 5511.484, 5513.714, 
    5508.663,
  5408.248, 5415.851, 5427.995, 5442.07, 5451.922, 5462.231, 5471.194, 
    5477.959, 5483.86, 5490.713, 5497.506, 5505.674, 5512.685, 5514.975, 
    5509.331,
  5568.248, 5538.429, 5513.756, 5491.227, 5476.259, 5475.69, 5477.102, 
    5483.97, 5489.793, 5501.746, 5511.904, 5523.655, 5534.474, 5542.906, 
    5543.799,
  5566.415, 5542.133, 5520.6, 5503.062, 5492.374, 5489.096, 5488.631, 
    5492.294, 5497.891, 5509.049, 5519.029, 5532.104, 5541.75, 5545.379, 
    5539.066,
  5561.635, 5543.514, 5526.705, 5512.389, 5502.993, 5505.033, 5498.316, 
    5500.489, 5507.129, 5517.27, 5529.028, 5541.665, 5545.85, 5542.145, 
    5531.093,
  5552.032, 5539.029, 5528.463, 5515.549, 5510.527, 5504.608, 5508.632, 
    5508.164, 5515.912, 5527.078, 5539.828, 5546.87, 5545.705, 5536.663, 
    5520.71,
  5538.727, 5530.363, 5525.089, 5517.949, 5510.529, 5511.882, 5512.165, 
    5514.927, 5527.129, 5537.393, 5546.006, 5547.928, 5540.882, 5525.754, 
    5509.402,
  5520.726, 5516.688, 5515.503, 5513.74, 5511.477, 5511.237, 5516.349, 
    5524.283, 5532.737, 5544.133, 5548.631, 5544.481, 5532.521, 5515.777, 
    5499.964,
  5502.381, 5502.178, 5505.398, 5506.802, 5508.539, 5513.435, 5518.116, 
    5528.288, 5540.019, 5547.17, 5547.856, 5538.787, 5522.635, 5506.292, 
    5493.646,
  5482.623, 5484.735, 5491.869, 5497.94, 5502.494, 5509.798, 5520.601, 
    5531.084, 5541.7, 5548.546, 5544.07, 5530.088, 5513.877, 5502.407, 5491.96,
  5463.722, 5467.296, 5479.078, 5490.619, 5498.906, 5508.846, 5520.243, 
    5534.459, 5545.493, 5546.079, 5537.358, 5522.115, 5510.272, 5502.713, 
    5493.577,
  5443.897, 5449.028, 5463.233, 5480.205, 5493.014, 5507.477, 5521.261, 
    5534.733, 5542.395, 5541.946, 5530.674, 5519.29, 5512.735, 5506.556, 
    5501.323,
  5661.018, 5652.478, 5642.845, 5627.917, 5612.383, 5597.251, 5582.411, 
    5573.143, 5565.336, 5556.574, 5551.308, 5549.704, 5551.439, 5554.346, 
    5555.788,
  5643.371, 5637.388, 5631.542, 5619.564, 5607.515, 5593.781, 5584.814, 
    5573.624, 5566.501, 5562.425, 5559.742, 5560.22, 5560.605, 5559.101, 
    5554.509,
  5620.963, 5617.119, 5613.439, 5607.022, 5597.578, 5592.245, 5577.028, 
    5574.743, 5566.792, 5562.535, 5562.526, 5563.779, 5561.357, 5555.834, 
    5545.306,
  5590.722, 5590.206, 5589.167, 5587.219, 5583.44, 5577.07, 5575.086, 
    5563.39, 5561.659, 5561.172, 5562.013, 5562.113, 5557.562, 5546.979, 
    5531.561,
  5554.913, 5557.687, 5560.176, 5563.438, 5565.504, 5566.034, 5561.146, 
    5561.14, 5556.556, 5556.389, 5559.617, 5556.391, 5548.335, 5533.042, 
    5515.671,
  5513.226, 5518.16, 5524.327, 5534.501, 5541.951, 5548.731, 5550.442, 
    5549.704, 5550.774, 5553.269, 5553.57, 5548.893, 5537.163, 5520.023, 
    5503.21,
  5469.917, 5477.187, 5487.227, 5503.198, 5518.652, 5530.815, 5537.317, 
    5541.98, 5544.033, 5547.416, 5547.521, 5540.549, 5525.144, 5509.026, 
    5495.171,
  5439.719, 5448.063, 5458.749, 5476.841, 5496.045, 5514.027, 5524.585, 
    5530.932, 5536.569, 5543.034, 5541.214, 5530.834, 5515.516, 5502.408, 
    5489.514,
  5421.265, 5431.255, 5445.422, 5463.756, 5483.453, 5500.801, 5513.293, 
    5523.884, 5532.308, 5538.053, 5535.068, 5523.613, 5509.824, 5497.471, 
    5484.027,
  5404.596, 5414.667, 5431.811, 5452.109, 5472.466, 5489.835, 5504.442, 
    5516.887, 5528.31, 5535.348, 5529.816, 5518.841, 5507.875, 5494.702, 
    5482.426,
  5656.5, 5653.018, 5651.109, 5646.511, 5641.773, 5634.523, 5625.911, 
    5618.838, 5609.273, 5598.986, 5591.771, 5584.76, 5580.06, 5575.5, 5572.59,
  5636.984, 5633.116, 5630.188, 5625.049, 5619.132, 5612.368, 5607.753, 
    5598.126, 5593.007, 5587.935, 5580.43, 5575.617, 5571.29, 5568.435, 
    5563.413,
  5610.271, 5605.128, 5599.51, 5593.896, 5587.915, 5585.535, 5576.546, 
    5580.582, 5571.28, 5568.186, 5564.231, 5561.499, 5557.68, 5554.499, 
    5548.985,
  5580.783, 5573.085, 5565.011, 5557.726, 5551.872, 5547.396, 5551.609, 
    5541.893, 5548.667, 5547.503, 5545.943, 5544.503, 5542.576, 5540.232, 
    5533.506,
  5550.031, 5539.078, 5526.822, 5517.241, 5510.089, 5507.323, 5505.342, 
    5519.085, 5515.631, 5520.231, 5524.546, 5525.421, 5525.868, 5523.033, 
    5518.024,
  5512.523, 5495.996, 5478.27, 5466.077, 5457.513, 5458.795, 5465.024, 
    5470.355, 5484.481, 5496.894, 5500.934, 5507.493, 5508.435, 5507.523, 
    5502.203,
  5470.387, 5449.933, 5429.945, 5415.34, 5406.578, 5408.219, 5419.319, 
    5439.538, 5454.727, 5468.356, 5481.703, 5489.775, 5492.85, 5492.803, 
    5487.468,
  5428.436, 5404.575, 5378.326, 5362.051, 5354.197, 5363.508, 5382.45, 
    5404.407, 5428.134, 5450.715, 5465.077, 5475.358, 5479.777, 5478.493, 
    5475.087,
  5389.245, 5363.873, 5343.401, 5329.433, 5325.184, 5337.024, 5361.371, 
    5391.211, 5416.69, 5437.354, 5453.524, 5464.526, 5467.745, 5467.649, 
    5464.843,
  5359.455, 5342.927, 5332.187, 5320.009, 5312.565, 5327.594, 5354.391, 
    5383.197, 5410.711, 5434.267, 5448.941, 5457.293, 5459.004, 5459.439, 
    5464.192,
  5605.525, 5608.707, 5611.403, 5611.518, 5612.655, 5611.546, 5610.555, 
    5610.334, 5605.985, 5599.038, 5593.559, 5587.322, 5579.935, 5571.795, 
    5564.409,
  5582.136, 5585.456, 5587.214, 5586.618, 5584.847, 5582.833, 5581.122, 
    5573.474, 5570.404, 5568.755, 5562.646, 5558.51, 5553.427, 5549.014, 
    5542.616,
  5556.902, 5560.739, 5562.287, 5561.657, 5558.252, 5556.152, 5546.039, 
    5549.676, 5539.402, 5536.307, 5533.266, 5531.274, 5527.439, 5524.646, 
    5521.254,
  5531.831, 5534.147, 5533.872, 5531.435, 5526.411, 5521.657, 5521.035, 
    5506.888, 5507.633, 5504.583, 5501.154, 5499.845, 5499.923, 5499.235, 
    5497.605,
  5508.759, 5510.287, 5509.449, 5506.991, 5502.465, 5494.723, 5483.658, 
    5483.389, 5469.812, 5462.545, 5464.596, 5462.928, 5467.054, 5468.318, 
    5472.047,
  5492.751, 5491.072, 5485.671, 5477.915, 5465.743, 5454.161, 5441.334, 
    5425.002, 5418.831, 5416.069, 5414.232, 5419.376, 5426.955, 5435.33, 
    5443.317,
  5471.043, 5466.077, 5456.156, 5444.482, 5429.476, 5410.399, 5391.689, 
    5379.865, 5368.144, 5362.755, 5368.753, 5378.002, 5390.971, 5405.578, 
    5418.932,
  5450.317, 5440.869, 5426.836, 5409.129, 5387.293, 5365.933, 5345.025, 
    5328.329, 5322.884, 5327.018, 5334.833, 5348.931, 5367.189, 5386.541, 
    5404.072,
  5422.393, 5411.158, 5395.508, 5376.181, 5355.736, 5333.94, 5314.352, 
    5302.14, 5296.199, 5301.542, 5315.656, 5334.405, 5355.291, 5377.153, 
    5396.771,
  5400.318, 5388.382, 5373.575, 5358.151, 5339.932, 5318.831, 5296.733, 
    5281.059, 5280.803, 5292.971, 5311.029, 5331.991, 5355.401, 5377.725, 
    5397.352,
  5522.362, 5525.948, 5532.148, 5537.558, 5544.329, 5550.561, 5556.087, 
    5563.685, 5570.106, 5574.431, 5578.95, 5580.989, 5580.188, 5577.816, 
    5575.258,
  5489.116, 5490.65, 5493.911, 5498.773, 5502.764, 5510.58, 5519.47, 
    5524.283, 5532.744, 5542.84, 5547.864, 5552.55, 5553.422, 5554.362, 
    5549.582,
  5466.389, 5462.383, 5459.779, 5462.372, 5466.901, 5477.071, 5477.979, 
    5493.833, 5495.777, 5506.521, 5514.507, 5521.33, 5523.282, 5523.714, 
    5522.5,
  5452.137, 5449.02, 5446.683, 5444.68, 5446.21, 5447.436, 5458.419, 
    5454.344, 5466.993, 5474.009, 5481.031, 5486.825, 5491.506, 5492.211, 
    5489.874,
  5437.756, 5434.335, 5432.107, 5431.8, 5432.451, 5434.216, 5433.792, 
    5441.234, 5443.055, 5443.513, 5451.622, 5453.153, 5457.375, 5457.222, 
    5458.472,
  5424.225, 5422.032, 5419.927, 5419.229, 5418.716, 5419.631, 5422.25, 
    5419.209, 5420.602, 5422.971, 5421.314, 5422.052, 5424.043, 5424.422, 
    5425.005,
  5413.688, 5412.339, 5410.996, 5409.081, 5408.119, 5406.117, 5403.221, 
    5402.281, 5397.674, 5391.573, 5389.758, 5388.403, 5388.798, 5390.854, 
    5393.7,
  5404.23, 5403.99, 5402.606, 5400.824, 5397.461, 5393.808, 5388.19, 
    5379.161, 5370.582, 5363.692, 5357.863, 5355.71, 5358.209, 5362.432, 
    5369.203,
  5391.953, 5390.498, 5387.814, 5384.761, 5380.116, 5374.062, 5365.824, 
    5356.32, 5343.176, 5331.351, 5325.01, 5326.121, 5331.094, 5341.608, 
    5353.836,
  5381.535, 5378.357, 5374.622, 5370.564, 5364.542, 5357.848, 5348.613, 
    5334.16, 5317.629, 5306.425, 5302.291, 5306.002, 5317.541, 5332.683, 
    5351.854,
  5572.342, 5576.714, 5582.497, 5585.302, 5587.961, 5585.773, 5579.62, 
    5573.836, 5562.922, 5546.793, 5533.692, 5521.067, 5509.807, 5501.652, 
    5498.804,
  5545.964, 5551.485, 5555.909, 5557.082, 5555.794, 5552.059, 5547.985, 
    5532.769, 5521.979, 5510.34, 5494.33, 5481.907, 5471.193, 5466.719, 
    5460.753,
  5518.629, 5524.211, 5526.853, 5527.609, 5525.124, 5524.542, 5509.206, 
    5509.588, 5489.334, 5474.697, 5460.217, 5448.558, 5437.545, 5432.675, 
    5431.297,
  5490.993, 5494.487, 5496.5, 5496.47, 5494.001, 5486.876, 5486.742, 
    5466.065, 5460.943, 5448.104, 5434.286, 5423.547, 5416.651, 5413.329, 
    5412.42,
  5462.943, 5465.151, 5465.887, 5464.382, 5461.584, 5456.643, 5446.687, 
    5447.768, 5434.744, 5424.177, 5418.778, 5410.097, 5406.018, 5402.208, 
    5404.134,
  5435.491, 5435.121, 5434.202, 5432.761, 5429.422, 5426.254, 5422.308, 
    5413.446, 5411.658, 5411.032, 5406.631, 5404.245, 5402.791, 5402.388, 
    5404.124,
  5415.122, 5413.772, 5411.608, 5409.905, 5407.765, 5404.754, 5401.738, 
    5401.721, 5398.349, 5395.904, 5397.118, 5399.21, 5400.577, 5402.589, 
    5405.838,
  5399.136, 5396.449, 5393.905, 5392.296, 5389.432, 5387.38, 5384.115, 
    5380.59, 5381.032, 5384.655, 5388.631, 5392.22, 5397.647, 5401.716, 
    5405.266,
  5386.372, 5384.426, 5381.47, 5379.114, 5375.802, 5371.553, 5367.439, 
    5365.297, 5363.889, 5365.559, 5372.187, 5381.824, 5389.631, 5398.109, 
    5404.91,
  5376.821, 5373.534, 5370.443, 5367.324, 5362.021, 5356.101, 5349.257, 
    5343.043, 5341.004, 5345.299, 5354.217, 5367.491, 5381.288, 5393.539, 
    5403.577,
  5537.889, 5562.251, 5586.783, 5608.752, 5629.493, 5644.991, 5656.654, 
    5665.619, 5669.41, 5666.881, 5661.52, 5650.232, 5632.618, 5608.641, 
    5580.224,
  5519.409, 5542.928, 5566.01, 5587.895, 5605.727, 5622.166, 5635.156, 
    5640.416, 5644.254, 5646.331, 5638.183, 5626.166, 5606.908, 5585.479, 
    5555.832,
  5501.444, 5524.376, 5546.336, 5567.702, 5584.255, 5602.482, 5605.387, 
    5621.459, 5618.279, 5617.859, 5611.731, 5600.04, 5580.755, 5557.797, 
    5534.724,
  5482.505, 5501.556, 5521.534, 5539.731, 5558.22, 5568.178, 5587.995, 
    5582.09, 5593.098, 5590.561, 5583.873, 5571.163, 5555.407, 5536.93, 
    5518.732,
  5464.037, 5480.039, 5496.196, 5513.182, 5528.317, 5544.999, 5547.909, 
    5565.041, 5561.267, 5557.104, 5554.934, 5543.287, 5532.121, 5517.887, 
    5506.266,
  5448.034, 5458.889, 5471.199, 5486.098, 5498.685, 5510.439, 5522.217, 
    5521.818, 5527.405, 5530.215, 5524.67, 5518.865, 5511.965, 5503.841, 
    5497.089,
  5433.242, 5440.411, 5449.348, 5459.43, 5471.406, 5481.465, 5489.224, 
    5498.996, 5500.961, 5499.633, 5500.523, 5498.638, 5495.19, 5492.029, 
    5489.159,
  5416.73, 5421.277, 5427.31, 5435.22, 5443.214, 5452.368, 5460.388, 
    5465.668, 5472.149, 5478.528, 5480.103, 5481.091, 5481.966, 5482.605, 
    5484.518,
  5401.541, 5404.771, 5408.545, 5413.575, 5419.528, 5426.46, 5433.84, 
    5442.938, 5450.008, 5455.594, 5461.991, 5467.514, 5471.881, 5475.601, 
    5482.149,
  5389.282, 5390.084, 5391.823, 5395.414, 5399.274, 5404.575, 5410.768, 
    5417.829, 5427.073, 5438.26, 5447.945, 5456.827, 5465.672, 5473.183, 
    5483.969,
  5527.392, 5550.096, 5574.014, 5598.701, 5622.871, 5646.336, 5669.091, 
    5690.646, 5707.166, 5717.697, 5724.575, 5726.814, 5722.753, 5712.345, 
    5696.849,
  5510.066, 5533.08, 5556.267, 5580.498, 5603.711, 5627.641, 5651.551, 
    5670.118, 5687.008, 5702.733, 5709.37, 5712.413, 5708.062, 5700.399, 
    5683.761,
  5492.04, 5513.464, 5536.81, 5561.712, 5584.876, 5612.011, 5628.207, 
    5657.179, 5670.106, 5682.999, 5691.754, 5695.88, 5692.307, 5683.553, 
    5668.735,
  5474.625, 5492.076, 5514.979, 5538.622, 5564.362, 5584.244, 5616.086, 
    5624.02, 5649.461, 5663.672, 5673.063, 5676.699, 5675.828, 5667.29, 
    5652.696,
  5456.89, 5471.892, 5491.35, 5516.008, 5540.408, 5567.873, 5583.924, 
    5616.371, 5627.824, 5640.519, 5653.016, 5656.719, 5656.958, 5648.434, 
    5637.564,
  5440.808, 5452.138, 5468.13, 5490.195, 5514.267, 5539.455, 5567.602, 
    5582.11, 5603.168, 5624.054, 5630.663, 5637.971, 5638.661, 5633.361, 
    5621.518,
  5425.775, 5435.035, 5447.914, 5466.537, 5490.157, 5515.274, 5538.858, 
    5567.913, 5587.937, 5598.473, 5611.548, 5618.9, 5619.398, 5614.274, 
    5602.047,
  5411.417, 5419.083, 5429.473, 5444.479, 5464.208, 5489.527, 5515.048, 
    5535.213, 5556.976, 5577.721, 5589.46, 5596.025, 5599.055, 5594.744, 
    5585.717,
  5396.502, 5404.404, 5414.696, 5427.413, 5444.687, 5465.487, 5490.417, 
    5517.137, 5538.27, 5553.12, 5565.546, 5574.471, 5577.853, 5575.751, 
    5569.439,
  5383.057, 5389.123, 5398.747, 5411.802, 5426.792, 5446.968, 5468.769, 
    5490.066, 5510.794, 5529.835, 5544.158, 5553.583, 5558.411, 5558.188, 
    5555.864,
  5541.181, 5558.196, 5584.181, 5608.087, 5631.09, 5651.756, 5671.36, 
    5691.652, 5709.109, 5722.837, 5733.923, 5741.023, 5743.425, 5741.109, 
    5733.476,
  5529.958, 5544.889, 5564.712, 5590.523, 5613.532, 5634.869, 5655.896, 
    5672.926, 5690.394, 5708.2, 5719.337, 5727.184, 5730.492, 5729.97, 
    5723.448,
  5516.544, 5531.435, 5548, 5569.179, 5594.772, 5619.919, 5634.521, 5660.312, 
    5674.459, 5689.23, 5702.331, 5711.758, 5716.392, 5715.974, 5712.005,
  5501.123, 5515.326, 5530.17, 5547.18, 5569.687, 5590.881, 5620.911, 
    5630.126, 5654.799, 5671.159, 5684.922, 5694.622, 5701.403, 5702.43, 
    5698.918,
  5481.007, 5496.381, 5511.071, 5527.15, 5545.333, 5569.69, 5586.777, 
    5618.754, 5633.646, 5648.74, 5666.38, 5676.364, 5684.855, 5686.471, 
    5685.38,
  5457.808, 5472.163, 5487.232, 5504.177, 5519.728, 5539.755, 5564.437, 
    5582.201, 5605.936, 5629.595, 5643.654, 5657.696, 5666.374, 5670.724, 
    5670.457,
  5432.396, 5445.95, 5461.537, 5478.748, 5497.081, 5515.142, 5534.068, 
    5561.443, 5583.031, 5600.109, 5621.234, 5636.346, 5646.783, 5653.119, 
    5654.748,
  5405.854, 5418.119, 5432.024, 5449.437, 5467.014, 5487.382, 5507.39, 
    5526.255, 5548.999, 5575.257, 5595.712, 5612.209, 5626.037, 5634.548, 
    5639.146,
  5381.199, 5392.423, 5405.705, 5421.891, 5439.747, 5458.699, 5478.868, 
    5502.846, 5525.698, 5545.949, 5567.429, 5588.166, 5603.661, 5615.294, 
    5621.574,
  5358.048, 5368.957, 5381.127, 5395.143, 5410.828, 5429.622, 5449.747, 
    5470.439, 5494.052, 5519.32, 5542.419, 5562.86, 5580.797, 5595.359, 
    5603.769,
  5509.694, 5520.297, 5537.893, 5558.469, 5582.671, 5607.169, 5633.249, 
    5661.984, 5687.927, 5711.893, 5731.241, 5747.594, 5756.333, 5761.317, 
    5759.467,
  5512.596, 5525.945, 5542.604, 5561.885, 5581.826, 5605.808, 5630.747, 
    5656.003, 5679.848, 5706.207, 5724.787, 5739.925, 5749.014, 5754.388, 
    5753.614,
  5508.929, 5528.155, 5543.389, 5563.565, 5582.074, 5606.237, 5625.989, 
    5654.276, 5676.911, 5697.362, 5715.737, 5730.16, 5739.567, 5744.789, 
    5745.797,
  5501.242, 5521.682, 5539.205, 5557.081, 5578.912, 5594.53, 5624.56, 
    5639.009, 5664.837, 5686.787, 5704.277, 5717.617, 5727.978, 5733.636, 
    5735.425,
  5490.308, 5509.513, 5528.073, 5549.131, 5567.716, 5592.811, 5605.958, 
    5635.186, 5655.605, 5671.451, 5690.065, 5702.61, 5713.631, 5719.625, 
    5723.84,
  5476.699, 5492.876, 5511.367, 5531.396, 5552.695, 5571.933, 5597.376, 
    5611.437, 5633.432, 5655.995, 5670.965, 5685.963, 5696.63, 5704.291, 
    5708.992,
  5455.648, 5471.745, 5490.386, 5510.757, 5532.761, 5554.917, 5573.676, 
    5598.157, 5617.098, 5632.121, 5650.276, 5664.675, 5676.469, 5685.743, 
    5691.875,
  5429.038, 5444.765, 5462.686, 5483.785, 5504.547, 5527.481, 5549.777, 
    5567.293, 5585.914, 5607.588, 5624.893, 5639.553, 5652.927, 5663.329, 
    5671.168,
  5397.377, 5412.625, 5431.261, 5452.886, 5475.451, 5497.52, 5518.747, 
    5542.122, 5562.327, 5578.203, 5594.021, 5609.581, 5623.306, 5635.366, 
    5645.554,
  5363.188, 5377.875, 5396.352, 5417.268, 5439.202, 5462.576, 5484.222, 
    5504.086, 5523.956, 5544.335, 5561.943, 5576.873, 5590.675, 5603.486, 
    5614.688,
  5408.028, 5419.442, 5446.003, 5477.659, 5514.65, 5552.683, 5597.686, 
    5638.625, 5675.561, 5703.415, 5725.379, 5746.485, 5761.916, 5772.467, 
    5776.045,
  5411.137, 5420.767, 5445.417, 5477.868, 5511.896, 5551.624, 5593.919, 
    5631.834, 5665.537, 5698.242, 5722.015, 5742.607, 5759.643, 5772.018, 
    5777.113,
  5421.917, 5427.236, 5450.024, 5480.077, 5514.241, 5553.752, 5589.912, 
    5630.569, 5662.995, 5690.575, 5716.021, 5736.927, 5755.062, 5767.35, 
    5775.548,
  5433.847, 5437.218, 5456.779, 5481.948, 5516.816, 5544.103, 5591.43, 
    5615.563, 5651.09, 5682.58, 5709.109, 5729.818, 5748.682, 5762.132, 
    5771.006,
  5439.868, 5448.761, 5463.998, 5488.978, 5515.747, 5551.524, 5574.601, 
    5619.096, 5645.806, 5672.152, 5699.401, 5720.399, 5739.496, 5752.688, 
    5762.951,
  5440.914, 5453.403, 5469.386, 5491.637, 5517.186, 5541.967, 5577.207, 
    5599.94, 5628.933, 5663.683, 5685.991, 5709.888, 5727.255, 5742.289, 
    5752.356,
  5437.691, 5451.588, 5469.012, 5491.993, 5517.234, 5541.6, 5564.616, 
    5600.216, 5626.759, 5646.34, 5672.606, 5694.476, 5712.186, 5727.104, 
    5737.579,
  5429.852, 5443.745, 5460.39, 5483.959, 5507.943, 5533.263, 5557.566, 
    5577.703, 5602.523, 5632.395, 5656.204, 5676.137, 5694.626, 5709.125, 
    5720.563,
  5415.236, 5430.332, 5448.017, 5470.228, 5496.291, 5521.221, 5545.981, 
    5572.968, 5596.373, 5615.952, 5636.307, 5656.538, 5673.407, 5687.785, 
    5699.013,
  5397.384, 5410.092, 5428.725, 5450.337, 5474.186, 5502.118, 5527.446, 
    5549.447, 5571.657, 5595.394, 5616.254, 5634.802, 5650.968, 5665.247, 
    5676.419,
  5404.65, 5403.135, 5419.979, 5450.5, 5489.672, 5533.583, 5576.719, 
    5625.407, 5659.897, 5688.709, 5709.652, 5725.387, 5734.022, 5738.012, 
    5737.481,
  5406.057, 5407.406, 5422.15, 5452.005, 5488.996, 5532.574, 5576.658, 
    5623.18, 5655.694, 5690.769, 5714.301, 5732.509, 5743.137, 5751.069, 
    5753.121,
  5412.553, 5414.897, 5430.263, 5456.935, 5492.436, 5537.222, 5575.712, 
    5627.452, 5662.13, 5692.034, 5717.365, 5737.093, 5751.757, 5760.404, 
    5765.929,
  5419.683, 5423.277, 5439.359, 5461.266, 5496.098, 5527.093, 5582.402, 
    5616.008, 5656.245, 5691.343, 5719.606, 5739.688, 5757.065, 5767.821, 
    5776.326,
  5424.325, 5432.067, 5447.258, 5469.455, 5495.626, 5535.97, 5568.122, 
    5624.852, 5660.607, 5690.212, 5718.829, 5740.646, 5759.832, 5771.952, 
    5781.827,
  5428.276, 5436.341, 5452.966, 5472.618, 5497.04, 5527.063, 5572.395, 
    5608.159, 5646.229, 5688.525, 5714.897, 5739.683, 5758.176, 5773.825, 
    5783.824,
  5430.993, 5439.127, 5457.127, 5475.078, 5501.107, 5529.501, 5561.773, 
    5610.656, 5650.911, 5679.822, 5710.258, 5734.68, 5754.391, 5770.634, 
    5781.626,
  5429.673, 5439.189, 5455.014, 5474.701, 5497.096, 5525.79, 5555.95, 
    5590.56, 5627.926, 5669.342, 5701.035, 5725.693, 5747.07, 5763.964, 
    5776.479,
  5425.033, 5435.014, 5451.103, 5470.939, 5494.188, 5519.694, 5546.684, 
    5585.947, 5624.792, 5657.452, 5686.898, 5714.002, 5735.478, 5753.079, 
    5765.774,
  5417.957, 5426.553, 5442.476, 5461.519, 5482.801, 5509.432, 5535.228, 
    5564.243, 5599.817, 5637.387, 5670.22, 5697.847, 5720.287, 5738.356, 
    5751.433,
  5479.718, 5481.107, 5488.431, 5504.18, 5529.154, 5555.154, 5584.204, 
    5609.91, 5633.073, 5647.614, 5656.79, 5657.728, 5657.523, 5663.001, 
    5667.58,
  5465.314, 5462.721, 5463.733, 5478.108, 5501.983, 5533.909, 5570.214, 
    5599.594, 5624.052, 5646.159, 5657.919, 5662.224, 5665.564, 5673.874, 
    5679.915,
  5453.689, 5446.487, 5444.036, 5455.768, 5479.546, 5516.961, 5552.235, 
    5595.968, 5625.075, 5645.041, 5659.697, 5667.946, 5677.248, 5687.367, 
    5696.752,
  5444.784, 5434.116, 5429.521, 5436.65, 5462.075, 5493.674, 5546.424, 
    5578.739, 5616.211, 5643.372, 5662.942, 5674.95, 5689.932, 5703.103, 
    5713.485,
  5438.935, 5427.644, 5421.082, 5427.835, 5449.27, 5488.757, 5527.917, 
    5582.706, 5618.131, 5643.149, 5665.611, 5683.075, 5702.464, 5715.777, 
    5728.181,
  5436.272, 5426.208, 5418.317, 5424.889, 5444.428, 5478.907, 5530.178, 
    5569.25, 5608.033, 5645.468, 5668.402, 5691.584, 5711.317, 5727.913, 
    5739.963,
  5435.583, 5428.937, 5423.148, 5429.476, 5449.617, 5482.372, 5526.282, 
    5577.025, 5616.714, 5645.009, 5672.665, 5697.864, 5718.828, 5736.195, 
    5749.721,
  5436.776, 5434.271, 5429.913, 5437.867, 5455.665, 5487.989, 5530.926, 
    5569.875, 5607.125, 5645.813, 5674.979, 5701.549, 5723.835, 5742.274, 
    5757.529,
  5438.482, 5440.57, 5441.062, 5450.152, 5468.556, 5496.96, 5535.219, 
    5578.668, 5615.239, 5647.17, 5675.274, 5703.439, 5725.616, 5745.341, 
    5761.595,
  5441.221, 5444.859, 5448.723, 5459.921, 5476.8, 5504.863, 5538.565, 
    5573.746, 5607.497, 5643.789, 5673.902, 5701.696, 5724.543, 5745.139, 
    5762.324,
  5545.29, 5546.539, 5556.211, 5567.605, 5582.409, 5594.658, 5605.561, 
    5614.878, 5622.538, 5627.171, 5628.45, 5621.37, 5613.774, 5603.717, 
    5599.71,
  5530.135, 5528.733, 5531.978, 5545.73, 5560.468, 5579.433, 5595.292, 
    5605.585, 5615.816, 5625.171, 5628.579, 5625.264, 5619.879, 5613.956, 
    5612.302,
  5511.664, 5509.488, 5509.79, 5518.745, 5535.044, 5560.454, 5577.426, 
    5601.581, 5611.379, 5621.229, 5627.396, 5628.226, 5626.618, 5623.203, 
    5624.141,
  5493.101, 5488.391, 5488.142, 5491.744, 5506.279, 5525.759, 5561.383, 
    5579.466, 5603.035, 5616.663, 5626.403, 5630.091, 5633.612, 5633.148, 
    5638.432,
  5475.103, 5468.584, 5465.946, 5469.107, 5477.75, 5500.819, 5527.197, 
    5568.9, 5593.481, 5609.093, 5623.235, 5631.776, 5639.497, 5641.969, 
    5650.723,
  5458.706, 5452.196, 5448.202, 5449.185, 5454.858, 5470.183, 5503.19, 
    5537.273, 5573.283, 5602.904, 5618.149, 5633.047, 5643.578, 5651.88, 
    5662.021,
  5448.741, 5443.75, 5438.291, 5435.115, 5438.536, 5450.225, 5475.217, 
    5520.301, 5562.059, 5591.337, 5613.433, 5632.555, 5647.435, 5658.252, 
    5672.167,
  5444.053, 5438.005, 5428.434, 5422.489, 5419.775, 5431.422, 5454.365, 
    5493.233, 5540.838, 5581.603, 5607.995, 5631.153, 5650.772, 5664.667, 
    5681.969,
  5441.152, 5433.953, 5422.723, 5412.405, 5406.382, 5415.146, 5438.101, 
    5481.094, 5531.908, 5572.422, 5601.913, 5630.293, 5652.305, 5670.091, 
    5689.145,
  5440.277, 5430.946, 5419.586, 5406.917, 5396.005, 5403.396, 5427.391, 
    5465.472, 5516.88, 5564.132, 5597.576, 5628.915, 5653.962, 5675.017, 
    5696.373,
  5588.331, 5595.296, 5603.701, 5609.851, 5618.247, 5625.691, 5631.091, 
    5637.016, 5640.856, 5642.736, 5645.695, 5649.95, 5657.368, 5667.718, 
    5677.605,
  5573.541, 5580.96, 5589.277, 5597.749, 5606.213, 5614.849, 5624.781, 
    5631.167, 5637.325, 5644.799, 5649.392, 5655.947, 5664.484, 5678.406, 
    5690.374,
  5551.892, 5561.047, 5569.316, 5580.312, 5588.186, 5603.262, 5608.857, 
    5625.625, 5633.891, 5641.909, 5649.509, 5657.607, 5669.111, 5683.747, 
    5699.406,
  5532.219, 5535.888, 5543.946, 5552.398, 5566.219, 5574.464, 5596.56, 
    5602.916, 5621.265, 5634.426, 5646.473, 5655.185, 5668.792, 5686.111, 
    5704.951,
  5519.109, 5519.318, 5520.137, 5525.837, 5534.826, 5551.794, 5564.005, 
    5591.088, 5608.62, 5621.929, 5638.081, 5650.755, 5665.065, 5684.159, 
    5705.475,
  5504.312, 5502.191, 5500.796, 5503.777, 5507.587, 5518.257, 5536.57, 
    5555.218, 5579.542, 5607.327, 5626.543, 5643.267, 5658.073, 5679.944, 
    5703.349,
  5491.157, 5487.263, 5484.389, 5484.213, 5487.855, 5494.489, 5505.218, 
    5528.583, 5559.094, 5585.386, 5611.666, 5633.123, 5650.229, 5671.449, 
    5697.395,
  5478.543, 5472.021, 5467.444, 5467.493, 5468.701, 5473.976, 5483.063, 
    5496.056, 5522.776, 5561.188, 5592.836, 5620.362, 5640.892, 5662.103, 
    5689.627,
  5467.597, 5458.656, 5451.012, 5447.518, 5448.034, 5453.254, 5461.732, 
    5477.27, 5500.902, 5535.929, 5571.86, 5605.297, 5629.871, 5651.916, 
    5679.335,
  5459.104, 5445.741, 5436.412, 5432.373, 5429.586, 5431.49, 5439.973, 
    5452.312, 5474.295, 5511.124, 5550.888, 5589.096, 5617.957, 5641.862, 
    5669.23 ;
}
