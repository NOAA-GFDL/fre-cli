netcdf \20030101.grid_spec.tile4 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 
    125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125,
  125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 
    125.7828, 125.7828, 125.7828, 125.7828, 125.7828, 125.7828,
  126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 
    126.5727, 126.5727, 126.5727, 126.5727, 126.5727, 126.5727,
  127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 
    127.3698, 127.3698, 127.3698, 127.3698, 127.3698, 127.3698,
  128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 
    128.1741, 128.1741, 128.1741, 128.1741, 128.1741, 128.1741,
  128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 
    128.9857, 128.9857, 128.9857, 128.9857, 128.9857, 128.9857,
  129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 
    129.8047, 129.8047, 129.8047, 129.8047, 129.8047, 129.8047,
  130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 
    130.6309, 130.6309, 130.6309, 130.6309, 130.6309, 130.6309,
  131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 
    131.4646, 131.4646, 131.4646, 131.4646, 131.4646, 131.4646,
  132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 
    132.3056, 132.3056, 132.3056, 132.3056, 132.3056, 132.3056,
  133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 
    133.1541, 133.1541, 133.1541, 133.1541, 133.1541, 133.1541,
  134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 
    134.01, 134.01, 134.01, 134.01, 134.01, 134.01, 134.01,
  134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 
    134.8733, 134.8733, 134.8733, 134.8733, 134.8733, 134.8733,
  135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 135.744, 
    135.744,
  136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 
    136.6221, 136.6221, 136.6221, 136.6221, 136.6221, 136.6221,
  137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 
    137.5075, 137.5075, 137.5075, 137.5075, 137.5075, 137.5075,
  138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 
    138.4002, 138.4002, 138.4002, 138.4002, 138.4002, 138.4002,
  139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 
    139.3002, 139.3002, 139.3002, 139.3002, 139.3002, 139.3002,
  140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 
    140.2074, 140.2074, 140.2074, 140.2074, 140.2074, 140.2074,
  141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 
    141.1216, 141.1216, 141.1216, 141.1216, 141.1216, 141.1216,
  142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 142.043, 
    142.043,
  142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 
    142.9712, 142.9712, 142.9712, 142.9712, 142.9712, 142.9712,
  143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 
    143.9063, 143.9063, 143.9063, 143.9063, 143.9063, 143.9063,
  144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 
    144.8482, 144.8482, 144.8482, 144.8482, 144.8482, 144.8482,
  145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 
    145.7966, 145.7966, 145.7966, 145.7966, 145.7966, 145.7966,
  146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 
    146.7514, 146.7514, 146.7514, 146.7514, 146.7514, 146.7514,
  147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 
    147.7126, 147.7126, 147.7126, 147.7126, 147.7126, 147.7126,
  148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 
    148.6799, 148.6799, 148.6799, 148.6799, 148.6799, 148.6799,
  149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 
    149.6532, 149.6532, 149.6532, 149.6532, 149.6532, 149.6532,
  150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 
    150.6322, 150.6322, 150.6322, 150.6322, 150.6322, 150.6322,
  151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 
    151.6168, 151.6168, 151.6168, 151.6168, 151.6168, 151.6168,
  152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 
    152.6068, 152.6068, 152.6068, 152.6068, 152.6068, 152.6068,
  153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 
    153.6019, 153.6019, 153.6019, 153.6019, 153.6019, 153.6019,
  154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 
    154.6019, 154.6019, 154.6019, 154.6019, 154.6019, 154.6019,
  155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 
    155.6065, 155.6065, 155.6065, 155.6065, 155.6065, 155.6065,
  156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 
    156.6156, 156.6156, 156.6156, 156.6156, 156.6156, 156.6156,
  157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 
    157.6287, 157.6287, 157.6287, 157.6287, 157.6287, 157.6287,
  158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 
    158.6458, 158.6458, 158.6458, 158.6458, 158.6458, 158.6458,
  159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 
    159.6663, 159.6663, 159.6663, 159.6663, 159.6663, 159.6663,
  160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 
    160.6902, 160.6902, 160.6902, 160.6902, 160.6902, 160.6902,
  161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 161.717, 
    161.717,
  162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 
    162.7465, 162.7465, 162.7465, 162.7465, 162.7465, 162.7465,
  163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 
    163.7783, 163.7783, 163.7783, 163.7783, 163.7783, 163.7783,
  164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 
    164.8122, 164.8122, 164.8122, 164.8122, 164.8122, 164.8122,
  165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 
    165.8477, 165.8477, 165.8477, 165.8477, 165.8477, 165.8477,
  166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 
    166.8846, 166.8846, 166.8846, 166.8846, 166.8846, 166.8846,
  167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 
    167.9225, 167.9225, 167.9225, 167.9225, 167.9225, 167.9225,
  168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 
    168.9611, 168.9611, 168.9611, 168.9611, 168.9611, 168.9611,
  170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 
    170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170,
  171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 
    171.0389, 171.0389, 171.0389, 171.0389, 171.0389, 171.0389,
  172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 
    172.0775, 172.0775, 172.0775, 172.0775, 172.0775, 172.0775,
  173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 
    173.1154, 173.1154, 173.1154, 173.1154, 173.1154, 173.1154,
  174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 
    174.1523, 174.1523, 174.1523, 174.1523, 174.1523, 174.1523,
  175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 
    175.1878, 175.1878, 175.1878, 175.1878, 175.1878, 175.1878,
  176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 
    176.2217, 176.2217, 176.2217, 176.2217, 176.2217, 176.2217,
  177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 
    177.2535, 177.2535, 177.2535, 177.2535, 177.2535, 177.2535,
  178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 178.283, 
    178.283,
  179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 
    179.3098, 179.3098, 179.3098, 179.3098, 179.3098, 179.3098,
  180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 
    180.3337, 180.3337, 180.3337, 180.3337, 180.3337, 180.3337,
  181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 
    181.3542, 181.3542, 181.3542, 181.3542, 181.3542, 181.3542,
  182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 
    182.3713, 182.3713, 182.3713, 182.3713, 182.3713, 182.3713,
  183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 
    183.3844, 183.3844, 183.3844, 183.3844, 183.3844, 183.3844,
  184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 
    184.3935, 184.3935, 184.3935, 184.3935, 184.3935, 184.3935,
  185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 
    185.3981, 185.3981, 185.3981, 185.3981, 185.3981, 185.3981,
  186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 
    186.3981, 186.3981, 186.3981, 186.3981, 186.3981, 186.3981,
  187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 
    187.3932, 187.3932, 187.3932, 187.3932, 187.3932, 187.3932,
  188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 
    188.3832, 188.3832, 188.3832, 188.3832, 188.3832, 188.3832,
  189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 
    189.3678, 189.3678, 189.3678, 189.3678, 189.3678, 189.3678,
  190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 
    190.3468, 190.3468, 190.3468, 190.3468, 190.3468, 190.3468,
  191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 
    191.3201, 191.3201, 191.3201, 191.3201, 191.3201, 191.3201,
  192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 
    192.2874, 192.2874, 192.2874, 192.2874, 192.2874, 192.2874,
  193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 
    193.2486, 193.2486, 193.2486, 193.2486, 193.2486, 193.2486,
  194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 
    194.2034, 194.2034, 194.2034, 194.2034, 194.2034, 194.2034,
  195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 
    195.1518, 195.1518, 195.1518, 195.1518, 195.1518, 195.1518,
  196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 
    196.0937, 196.0937, 196.0937, 196.0937, 196.0937, 196.0937,
  197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 
    197.0288, 197.0288, 197.0288, 197.0288, 197.0288, 197.0288,
  197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 197.957, 
    197.957,
  198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 
    198.8784, 198.8784, 198.8784, 198.8784, 198.8784, 198.8784,
  199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 
    199.7926, 199.7926, 199.7926, 199.7926, 199.7926, 199.7926,
  200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 
    200.6998, 200.6998, 200.6998, 200.6998, 200.6998, 200.6998,
  201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 
    201.5998, 201.5998, 201.5998, 201.5998, 201.5998, 201.5998,
  202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 
    202.4925, 202.4925, 202.4925, 202.4925, 202.4925, 202.4925,
  203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 
    203.3779, 203.3779, 203.3779, 203.3779, 203.3779, 203.3779,
  204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 204.256, 
    204.256,
  205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 
    205.1267, 205.1267, 205.1267, 205.1267, 205.1267, 205.1267,
  205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 
    205.99, 205.99, 205.99, 205.99, 205.99, 205.99, 205.99,
  206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 
    206.8459, 206.8459, 206.8459, 206.8459, 206.8459, 206.8459,
  207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 
    207.6944, 207.6944, 207.6944, 207.6944, 207.6944, 207.6944,
  208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 
    208.5354, 208.5354, 208.5354, 208.5354, 208.5354, 208.5354,
  209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 
    209.3691, 209.3691, 209.3691, 209.3691, 209.3691, 209.3691,
  210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 
    210.1953, 210.1953, 210.1953, 210.1953, 210.1953, 210.1953,
  211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 
    211.0143, 211.0143, 211.0143, 211.0143, 211.0143, 211.0143,
  211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 
    211.8259, 211.8259, 211.8259, 211.8259, 211.8259, 211.8259,
  212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 
    212.6302, 212.6302, 212.6302, 212.6302, 212.6302, 212.6302,
  213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 
    213.4273, 213.4273, 213.4273, 213.4273, 213.4273, 213.4273,
  214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 
    214.2172, 214.2172, 214.2172, 214.2172, 214.2172, 214.2172,
  215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 
    215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215 ;

 grid_lat =
  35.26439, 34.52972, 33.79504, 33.06036, 32.32569, 31.59101, 30.85634, 
    30.12167, 29.38699, 28.65232, 27.91764, 27.18297, 26.44829, 25.71362, 
    24.97894, 24.24427, 23.50959, 22.77492, 22.04024, 21.30557, 20.57089, 
    19.83622, 19.10155, 18.36687, 17.63219, 16.89752, 16.16285, 15.42817, 
    14.6935, 13.95882, 13.22415, 12.48947, 11.7548, 11.02012, 10.28545, 
    9.550773, 8.816097, 8.081423, 7.346748, 6.612073, 5.877398, 5.142724, 
    4.408049, 3.673374, 2.938699, 2.204024, 1.46935, 0.7346748, 0, 
    -0.7346748, -1.46935, -2.204024, -2.938699, -3.673374, -4.408049, 
    -5.142724, -5.877398, -6.612073, -7.346748, -8.081423, -8.816097, 
    -9.550773, -10.28545, -11.02012, -11.7548, -12.48947, -13.22415, 
    -13.95882, -14.6935, -15.42817, -16.16285, -16.89752, -17.63219, 
    -18.36687, -19.10155, -19.83622, -20.57089, -21.30557, -22.04024, 
    -22.77492, -23.50959, -24.24427, -24.97894, -25.71362, -26.44829, 
    -27.18297, -27.91764, -28.65232, -29.38699, -30.12167, -30.85634, 
    -31.59101, -32.32569, -33.06036, -33.79504, -34.52972, -35.26439,
  35.62921, 34.89117, 34.15289, 33.41436, 32.67561, 31.93662, 31.19741, 
    30.45796, 29.7183, 28.97841, 28.23831, 27.49799, 26.75747, 26.01674, 
    25.2758, 24.53467, 23.79335, 23.05183, 22.31014, 21.56826, 20.8262, 
    20.08398, 19.34159, 18.59904, 17.85633, 17.11348, 16.37048, 15.62734, 
    14.88407, 14.14067, 13.39715, 12.65351, 11.90976, 11.16591, 10.42197, 
    9.677926, 8.933801, 8.189597, 7.445321, 6.700978, 5.956575, 5.21212, 
    4.467618, 3.723077, 2.978501, 2.233899, 1.489277, 0.744642, 0, -0.744642, 
    -1.489277, -2.233899, -2.978501, -3.723077, -4.467618, -5.21212, 
    -5.956575, -6.700978, -7.445321, -8.189597, -8.933801, -9.677926, 
    -10.42197, -11.16591, -11.90976, -12.65351, -13.39715, -14.14067, 
    -14.88407, -15.62734, -16.37048, -17.11348, -17.85633, -18.59904, 
    -19.34159, -20.08398, -20.8262, -21.56826, -22.31014, -23.05183, 
    -23.79335, -24.53467, -25.2758, -26.01674, -26.75747, -27.49799, 
    -28.23831, -28.97841, -29.7183, -30.45796, -31.19741, -31.93662, 
    -32.67561, -33.41436, -34.15289, -34.89117, -35.62921,
  35.98892, 35.24767, 34.50594, 33.76374, 33.02107, 32.27793, 31.53433, 
    30.79028, 30.04578, 29.30084, 28.55546, 27.80966, 27.06343, 26.31679, 
    25.56974, 24.82229, 24.07445, 23.32623, 22.57764, 21.82868, 21.07937, 
    20.32972, 19.57973, 18.82941, 18.07879, 17.32786, 16.57663, 15.82513, 
    15.07335, 14.32132, 13.56903, 12.81652, 12.06378, 11.31083, 10.55768, 
    9.804344, 9.050837, 8.297169, 7.543353, 6.789403, 6.035332, 5.281153, 
    4.526879, 3.772523, 3.0181, 2.263623, 1.509105, 0.7545591, 0, -0.7545591, 
    -1.509105, -2.263623, -3.0181, -3.772523, -4.526879, -5.281153, 
    -6.035332, -6.789403, -7.543353, -8.297169, -9.050837, -9.804344, 
    -10.55768, -11.31083, -12.06378, -12.81652, -13.56903, -14.32132, 
    -15.07335, -15.82513, -16.57663, -17.32786, -18.07879, -18.82941, 
    -19.57973, -20.32972, -21.07937, -21.82868, -22.57764, -23.32623, 
    -24.07445, -24.82229, -25.56974, -26.31679, -27.06343, -27.80966, 
    -28.55546, -29.30084, -30.04578, -30.79028, -31.53433, -32.27793, 
    -33.02107, -33.76374, -34.50594, -35.24767, -35.98892,
  36.34341, 35.59911, 34.8541, 34.10837, 33.36194, 32.61481, 31.86699, 
    31.11849, 30.36931, 29.61947, 28.86897, 28.11782, 27.36604, 26.61363, 
    25.86061, 25.10699, 24.35277, 23.59798, 22.84263, 22.08672, 21.33028, 
    20.57332, 19.81585, 19.05788, 18.29944, 17.54054, 16.7812, 16.02143, 
    15.26124, 14.50067, 13.73972, 12.97841, 12.21676, 11.45479, 10.69252, 
    9.929964, 9.167146, 8.404083, 7.640796, 6.877304, 6.113627, 5.349786, 
    4.5858, 3.82169, 3.057476, 2.29318, 1.528821, 0.7644209, 0, -0.7644209, 
    -1.528821, -2.29318, -3.057476, -3.82169, -4.5858, -5.349786, -6.113627, 
    -6.877304, -7.640796, -8.404083, -9.167146, -9.929964, -10.69252, 
    -11.45479, -12.21676, -12.97841, -13.73972, -14.50067, -15.26124, 
    -16.02143, -16.7812, -17.54054, -18.29944, -19.05788, -19.81585, 
    -20.57332, -21.33028, -22.08672, -22.84263, -23.59798, -24.35277, 
    -25.10699, -25.86061, -26.61363, -27.36604, -28.11782, -28.86897, 
    -29.61947, -30.36931, -31.11849, -31.86699, -32.61481, -33.36194, 
    -34.10837, -34.8541, -35.59911, -36.34341,
  36.69255, 35.94537, 35.19722, 34.44813, 33.6981, 32.94714, 32.19525, 
    31.44245, 30.68875, 29.93416, 29.17869, 28.42235, 27.66517, 26.90714, 
    26.14829, 25.38863, 24.62818, 23.86696, 23.10497, 22.34225, 21.5788, 
    20.81466, 20.04982, 19.28433, 18.51819, 17.75143, 16.98408, 16.21614, 
    15.44765, 14.67863, 13.90911, 13.1391, 12.36863, 11.59772, 10.82641, 
    10.05472, 9.282667, 8.510284, 7.737598, 6.964634, 6.19142, 5.417983, 
    4.64435, 3.870549, 3.096608, 2.322554, 1.548416, 0.7742223, 1.272222e-14, 
    -0.7742223, -1.548416, -2.322554, -3.096608, -3.870549, -4.64435, 
    -5.417983, -6.19142, -6.964634, -7.737598, -8.510284, -9.282667, 
    -10.05472, -10.82641, -11.59772, -12.36863, -13.1391, -13.90911, 
    -14.67863, -15.44765, -16.21614, -16.98408, -17.75143, -18.51819, 
    -19.28433, -20.04982, -20.81466, -21.5788, -22.34225, -23.10497, 
    -23.86696, -24.62818, -25.38863, -26.14829, -26.90714, -27.66517, 
    -28.42235, -29.17869, -29.93416, -30.68875, -31.44245, -32.19525, 
    -32.94714, -33.6981, -34.44813, -35.19722, -35.94537, -36.69255,
  37.03624, 36.28631, 35.53519, 34.78289, 34.02942, 33.27477, 32.51897, 
    31.76203, 31.00396, 30.24478, 29.48449, 28.72311, 27.96067, 27.19717, 
    26.43264, 25.66709, 24.90054, 24.13302, 23.36455, 22.59513, 21.82482, 
    21.05361, 20.28154, 19.50863, 18.73492, 17.96042, 17.18516, 16.40917, 
    15.63248, 14.85512, 14.07711, 13.2985, 12.5193, 11.73955, 10.95929, 
    10.17854, 9.397336, 8.615713, 7.833705, 7.051345, 6.268667, 5.485706, 
    4.702497, 3.919074, 3.135473, 2.35173, 1.56788, 0.7839577, 1.272222e-14, 
    -0.7839577, -1.56788, -2.35173, -3.135473, -3.919074, -4.702497, 
    -5.485706, -6.268667, -7.051345, -7.833705, -8.615713, -9.397336, 
    -10.17854, -10.95929, -11.73955, -12.5193, -13.2985, -14.07711, 
    -14.85512, -15.63248, -16.40917, -17.18516, -17.96042, -18.73492, 
    -19.50863, -20.28154, -21.05361, -21.82482, -22.59513, -23.36455, 
    -24.13302, -24.90054, -25.66709, -26.43264, -27.19717, -27.96067, 
    -28.72311, -29.48449, -30.24478, -31.00396, -31.76203, -32.51897, 
    -33.27477, -34.02942, -34.78289, -35.53519, -36.28631, -37.03624,
  37.37434, 36.62183, 35.86789, 35.11252, 34.35575, 33.59758, 32.83802, 
    32.0771, 31.31481, 30.55118, 29.78622, 29.01996, 28.25241, 27.48358, 
    26.71351, 25.94222, 25.16972, 24.39604, 23.6212, 22.84524, 22.06818, 
    21.29005, 20.51087, 19.73068, 18.9495, 18.16737, 17.38433, 16.6004, 
    15.81561, 15.03002, 14.24364, 13.45652, 12.66869, 11.88019, 11.09107, 
    10.30135, 9.511086, 8.720308, 7.929061, 7.137385, 6.345323, 5.552916, 
    4.760206, 3.967237, 3.17405, 2.38069, 1.587199, 0.7936214, 1.272222e-14, 
    -0.7936214, -1.587199, -2.38069, -3.17405, -3.967237, -4.760206, 
    -5.552916, -6.345323, -7.137385, -7.929061, -8.720308, -9.511086, 
    -10.30135, -11.09107, -11.88019, -12.66869, -13.45652, -14.24364, 
    -15.03002, -15.81561, -16.6004, -17.38433, -18.16737, -18.9495, 
    -19.73068, -20.51087, -21.29005, -22.06818, -22.84524, -23.6212, 
    -24.39604, -25.16972, -25.94222, -26.71351, -27.48358, -28.25241, 
    -29.01996, -29.78622, -30.55118, -31.31481, -32.0771, -32.83802, 
    -33.59758, -34.35575, -35.11252, -35.86789, -36.62183, -37.37434,
  37.70675, 36.95179, 36.19517, 35.4369, 34.67698, 33.91543, 33.15226, 
    32.3875, 31.62114, 30.85322, 30.08375, 29.31275, 28.54023, 27.76624, 
    26.99077, 26.21387, 25.43556, 24.65587, 23.87482, 23.09244, 22.30877, 
    21.52384, 20.73768, 19.95033, 19.16182, 18.37219, 17.58147, 16.78971, 
    15.99695, 15.20323, 14.40859, 13.61306, 12.81671, 12.01956, 11.22167, 
    10.42309, 9.623848, 8.824006, 8.023608, 7.222704, 6.421341, 5.619571, 
    4.817443, 4.015007, 3.212315, 2.409416, 1.606363, 0.8032075, 
    1.272222e-14, -0.8032075, -1.606363, -2.409416, -3.212315, -4.015007, 
    -4.817443, -5.619571, -6.421341, -7.222704, -8.023608, -8.824006, 
    -9.623848, -10.42309, -11.22167, -12.01956, -12.81671, -13.61306, 
    -14.40859, -15.20323, -15.99695, -16.78971, -17.58147, -18.37219, 
    -19.16182, -19.95033, -20.73768, -21.52384, -22.30877, -23.09244, 
    -23.87482, -24.65587, -25.43556, -26.21387, -26.99077, -27.76624, 
    -28.54023, -29.31275, -30.08375, -30.85322, -31.62114, -32.3875, 
    -33.15226, -33.91543, -34.67698, -35.4369, -36.19517, -36.95179, -37.70675,
  38.03334, 37.27608, 36.51693, 35.75588, 34.99296, 34.22818, 33.46156, 
    32.6931, 31.92283, 31.15076, 30.37692, 29.60133, 28.82401, 28.04498, 
    27.26427, 26.48191, 25.69794, 24.91236, 24.12524, 23.33659, 22.54645, 
    21.75485, 20.96184, 20.16746, 19.37174, 18.57473, 17.77647, 16.97701, 
    16.17639, 15.37465, 14.57185, 13.76804, 12.96326, 12.15757, 11.35102, 
    10.54366, 9.735553, 8.926742, 8.117288, 7.307246, 6.496675, 5.68563, 
    4.874171, 4.062356, 3.250242, 2.437891, 1.62536, 0.8127099, 1.272222e-14, 
    -0.8127099, -1.62536, -2.437891, -3.250242, -4.062356, -4.874171, 
    -5.68563, -6.496675, -7.307246, -8.117288, -8.926742, -9.735553, 
    -10.54366, -11.35102, -12.15757, -12.96326, -13.76804, -14.57185, 
    -15.37465, -16.17639, -16.97701, -17.77647, -18.57473, -19.37174, 
    -20.16746, -20.96184, -21.75485, -22.54645, -23.33659, -24.12524, 
    -24.91236, -25.69794, -26.48191, -27.26427, -28.04498, -28.82401, 
    -29.60133, -30.37692, -31.15076, -31.92283, -32.6931, -33.46156, 
    -34.22818, -34.99296, -35.75588, -36.51693, -37.27608, -38.03334,
  38.354, 37.59457, 36.83301, 36.06934, 35.30357, 34.5357, 33.76576, 
    32.99376, 32.21972, 31.44366, 30.6656, 29.88556, 29.10357, 28.31966, 
    27.53386, 26.74619, 25.95669, 25.16539, 24.37232, 23.57754, 22.78106, 
    21.98295, 21.18322, 20.38194, 19.57915, 18.77489, 17.96921, 17.16216, 
    16.3538, 15.54417, 14.73334, 13.92135, 13.10826, 12.29414, 11.47903, 
    10.66301, 9.846126, 9.028447, 8.210036, 7.390956, 6.571271, 5.751048, 
    4.930352, 4.10925, 3.287808, 2.466094, 1.644176, 0.8221223, 1.272222e-14, 
    -0.8221223, -1.644176, -2.466094, -3.287808, -4.10925, -4.930352, 
    -5.751048, -6.571271, -7.390956, -8.210036, -9.028447, -9.846126, 
    -10.66301, -11.47903, -12.29414, -13.10826, -13.92135, -14.73334, 
    -15.54417, -16.3538, -17.16216, -17.96921, -18.77489, -19.57915, 
    -20.38194, -21.18322, -21.98295, -22.78106, -23.57754, -24.37232, 
    -25.16539, -25.95669, -26.74619, -27.53386, -28.31966, -29.10357, 
    -29.88556, -30.6656, -31.44366, -32.21972, -32.99376, -33.76576, 
    -34.5357, -35.30357, -36.06934, -36.83301, -37.59457, -38.354,
  38.66859, 37.90713, 37.14331, 36.37715, 35.60866, 34.83784, 34.06473, 
    33.28933, 32.51167, 31.73176, 30.94962, 30.16529, 29.37879, 28.59014, 
    27.79938, 27.00655, 26.21167, 25.41478, 24.61593, 23.81515, 23.01249, 
    22.20798, 21.40168, 20.59364, 19.7839, 18.97252, 18.15956, 17.34505, 
    16.52908, 15.71168, 14.89293, 14.07288, 13.2516, 12.42916, 11.60561, 
    10.78103, 9.955491, 9.129053, 8.30179, 7.473776, 6.645081, 5.815781, 
    4.985948, 4.155657, 3.324986, 2.494007, 1.662799, 0.8314381, 
    1.272222e-14, -0.8314381, -1.662799, -2.494007, -3.324986, -4.155657, 
    -4.985948, -5.815781, -6.645081, -7.473776, -8.30179, -9.129053, 
    -9.955491, -10.78103, -11.60561, -12.42916, -13.2516, -14.07288, 
    -14.89293, -15.71168, -16.52908, -17.34505, -18.15956, -18.97252, 
    -19.7839, -20.59364, -21.40168, -22.20798, -23.01249, -23.81515, 
    -24.61593, -25.41478, -26.21167, -27.00655, -27.79938, -28.59014, 
    -29.37879, -30.16529, -30.94962, -31.73176, -32.51167, -33.28933, 
    -34.06473, -34.83784, -35.60866, -36.37715, -37.14331, -37.90713, 
    -38.66859,
  38.977, 38.21363, 37.44768, 36.67916, 35.90809, 35.13448, 34.35833, 
    33.57967, 32.79853, 32.01491, 31.22885, 30.44036, 29.64949, 28.85626, 
    28.0607, 27.26284, 26.46273, 25.6604, 24.85591, 24.04927, 23.24056, 
    22.42981, 21.61708, 20.80241, 19.98587, 19.16751, 18.34738, 17.52556, 
    16.7021, 15.87706, 15.05052, 14.22254, 13.39319, 12.56255, 11.73068, 
    10.89766, 10.06357, 9.228487, 8.392486, 7.555646, 6.718051, 5.87978, 
    5.040917, 4.201545, 3.361748, 2.52161, 1.681216, 0.8406506, 1.272222e-14, 
    -0.8406506, -1.681216, -2.52161, -3.361748, -4.201545, -5.040917, 
    -5.87978, -6.718051, -7.555646, -8.392486, -9.228487, -10.06357, 
    -10.89766, -11.73068, -12.56255, -13.39319, -14.22254, -15.05052, 
    -15.87706, -16.7021, -17.52556, -18.34738, -19.16751, -19.98587, 
    -20.80241, -21.61708, -22.42981, -23.24056, -24.04927, -24.85591, 
    -25.6604, -26.46273, -27.26284, -28.0607, -28.85626, -29.64949, 
    -30.44036, -31.22885, -32.01491, -32.79853, -33.57967, -34.35833, 
    -35.13448, -35.90809, -36.67916, -37.44768, -38.21363, -38.977,
  39.27911, 38.51395, 37.746, 36.97525, 36.20173, 35.42545, 34.64641, 
    33.86464, 33.08015, 32.29297, 31.50312, 30.71063, 29.91554, 29.11786, 
    28.31764, 27.51491, 26.70972, 25.9021, 25.0921, 24.27976, 23.46515, 
    22.6483, 21.82927, 21.00812, 20.18491, 19.35971, 18.53256, 17.70355, 
    16.87274, 16.0402, 15.20599, 14.37021, 13.53292, 12.6942, 11.85414, 
    11.0128, 10.17029, 9.326677, 8.482054, 7.636507, 6.790126, 5.943, 
    5.095221, 4.246879, 3.398068, 2.548881, 1.699411, 0.8497528, 
    1.272222e-14, -0.8497528, -1.699411, -2.548881, -3.398068, -4.246879, 
    -5.095221, -5.943, -6.790126, -7.636507, -8.482054, -9.326677, -10.17029, 
    -11.0128, -11.85414, -12.6942, -13.53292, -14.37021, -15.20599, -16.0402, 
    -16.87274, -17.70355, -18.53256, -19.35971, -20.18491, -21.00812, 
    -21.82927, -22.6483, -23.46515, -24.27976, -25.0921, -25.9021, -26.70972, 
    -27.51491, -28.31764, -29.11786, -29.91554, -30.71063, -31.50312, 
    -32.29297, -33.08015, -33.86464, -34.64641, -35.42545, -36.20173, 
    -36.97525, -37.746, -38.51395, -39.27911,
  39.57478, 38.80796, 38.03813, 37.26529, 36.48944, 35.71062, 34.92882, 
    34.14407, 33.35638, 32.56578, 31.77229, 30.97594, 30.17676, 29.37479, 
    28.57006, 27.76261, 26.95247, 26.13971, 25.32435, 24.50646, 23.68609, 
    22.86328, 22.03811, 21.21062, 20.38089, 19.54898, 18.71496, 17.8789, 
    17.04088, 16.20097, 15.35924, 14.51579, 13.67069, 12.82403, 11.97589, 
    11.12637, 10.27556, 9.423547, 8.570426, 7.716295, 6.86125, 6.00539, 
    5.148814, 4.291623, 3.433917, 2.575799, 1.717372, 0.8587376, 
    1.272222e-14, -0.8587376, -1.717372, -2.575799, -3.433917, -4.291623, 
    -5.148814, -6.00539, -6.86125, -7.716295, -8.570426, -9.423547, 
    -10.27556, -11.12637, -11.97589, -12.82403, -13.67069, -14.51579, 
    -15.35924, -16.20097, -17.04088, -17.8789, -18.71496, -19.54898, 
    -20.38089, -21.21062, -22.03811, -22.86328, -23.68609, -24.50646, 
    -25.32435, -26.13971, -26.95247, -27.76261, -28.57006, -29.37479, 
    -30.17676, -30.97594, -31.77229, -32.56578, -33.35638, -34.14407, 
    -34.92882, -35.71062, -36.48944, -37.26529, -38.03813, -38.80796, 
    -39.57478,
  39.8639, 39.09554, 38.32394, 37.54912, 36.77109, 35.98985, 35.20542, 
    34.41782, 33.62707, 32.83318, 32.03619, 31.23613, 30.43301, 29.62689, 
    28.81779, 28.00576, 27.19084, 26.37307, 25.55252, 24.72922, 23.90323, 
    23.07462, 22.24345, 21.40977, 20.57367, 19.7352, 18.89445, 18.05148, 
    17.20639, 16.35925, 15.51014, 14.65916, 13.80638, 12.95192, 12.09585, 
    11.23828, 10.3793, 9.519018, 8.657532, 7.794946, 6.931367, 6.066901, 
    5.201655, 4.335741, 3.469266, 2.602343, 1.735083, 0.8675976, 
    1.272222e-14, -0.8675976, -1.735083, -2.602343, -3.469266, -4.335741, 
    -5.201655, -6.066901, -6.931367, -7.794946, -8.657532, -9.519018, 
    -10.3793, -11.23828, -12.09585, -12.95192, -13.80638, -14.65916, 
    -15.51014, -16.35925, -17.20639, -18.05148, -18.89445, -19.7352, 
    -20.57367, -21.40977, -22.24345, -23.07462, -23.90323, -24.72922, 
    -25.55252, -26.37307, -27.19084, -28.00576, -28.81779, -29.62689, 
    -30.43301, -31.23613, -32.03619, -32.83318, -33.62707, -34.41782, 
    -35.20542, -35.98985, -36.77109, -37.54912, -38.32394, -39.09554, -39.8639,
  40.14635, 39.37654, 38.6033, 37.82662, 37.04652, 36.26299, 35.47607, 
    34.68575, 33.89207, 33.09504, 32.29469, 31.49104, 30.68413, 29.874, 
    29.06068, 28.24422, 27.42466, 26.60204, 25.77643, 24.94787, 24.11643, 
    23.28216, 22.44514, 21.60542, 20.76309, 19.91821, 19.07088, 18.22116, 
    17.36914, 16.51492, 15.65857, 14.8002, 13.9399, 13.07777, 12.21391, 
    11.34843, 10.48143, 9.613013, 8.743299, 7.872395, 7.000417, 6.12748, 
    5.253699, 4.379195, 3.504085, 2.628489, 1.752529, 0.8763254, 
    1.272222e-14, -0.8763254, -1.752529, -2.628489, -3.504085, -4.379195, 
    -5.253699, -6.12748, -7.000417, -7.872395, -8.743299, -9.613013, 
    -10.48143, -11.34843, -12.21391, -13.07777, -13.9399, -14.8002, 
    -15.65857, -16.51492, -17.36914, -18.22116, -19.07088, -19.91821, 
    -20.76309, -21.60542, -22.44514, -23.28216, -24.11643, -24.94787, 
    -25.77643, -26.60204, -27.42466, -28.24422, -29.06068, -29.874, 
    -30.68413, -31.49104, -32.29469, -33.09504, -33.89207, -34.68575, 
    -35.47607, -36.26299, -37.04652, -37.82662, -38.6033, -39.37654, -40.14635,
  40.42199, 39.65086, 38.87608, 38.09766, 37.3156, 36.52991, 35.74061, 
    34.94771, 34.15122, 33.35118, 32.5476, 31.74052, 30.92996, 30.11596, 
    29.29857, 28.47782, 27.65377, 26.82645, 25.99593, 25.16227, 24.32551, 
    23.48574, 22.64302, 21.79742, 20.94901, 20.09789, 19.24412, 18.38779, 
    17.52901, 16.66785, 15.80442, 14.93881, 14.07113, 13.20149, 12.32998, 
    11.45673, 10.58185, 9.705451, 8.827652, 7.948575, 7.068341, 6.187074, 
    5.304901, 4.421948, 3.538343, 2.654216, 1.769696, 0.8849133, 
    1.272222e-14, -0.8849133, -1.769696, -2.654216, -3.538343, -4.421948, 
    -5.304901, -6.187074, -7.068341, -7.948575, -8.827652, -9.705451, 
    -10.58185, -11.45673, -12.32998, -13.20149, -14.07113, -14.93881, 
    -15.80442, -16.66785, -17.52901, -18.38779, -19.24412, -20.09789, 
    -20.94901, -21.79742, -22.64302, -23.48574, -24.32551, -25.16227, 
    -25.99593, -26.82645, -27.65377, -28.47782, -29.29857, -30.11596, 
    -30.92996, -31.74052, -32.5476, -33.35118, -34.15122, -34.94771, 
    -35.74061, -36.52991, -37.3156, -38.09766, -38.87608, -39.65086, -40.42199,
  40.69072, 39.91835, 39.14214, 38.36209, 37.57819, 36.79046, 35.9989, 
    35.20354, 34.40438, 33.60146, 32.79479, 31.98441, 31.17034, 30.35262, 
    29.5313, 28.70641, 27.87801, 27.04614, 26.21087, 25.37224, 24.53034, 
    23.68522, 22.83695, 21.98561, 21.13129, 20.27407, 19.41402, 18.55125, 
    17.68585, 16.81791, 15.94755, 15.07486, 14.19996, 13.32295, 12.44396, 
    11.5631, 10.68048, 9.79625, 8.910519, 8.023417, 7.135077, 6.245632, 
    5.355214, 4.463961, 3.57201, 2.679499, 1.786567, 0.8933536, 1.272222e-14, 
    -0.8933536, -1.786567, -2.679499, -3.57201, -4.463961, -5.355214, 
    -6.245632, -7.135077, -8.023417, -8.910519, -9.79625, -10.68048, 
    -11.5631, -12.44396, -13.32295, -14.19996, -15.07486, -15.94755, 
    -16.81791, -17.68585, -18.55125, -19.41402, -20.27407, -21.13129, 
    -21.98561, -22.83695, -23.68522, -24.53034, -25.37224, -26.21087, 
    -27.04614, -27.87801, -28.70641, -29.5313, -30.35262, -31.17034, 
    -31.98441, -32.79479, -33.60146, -34.40438, -35.20354, -35.9989, 
    -36.79046, -37.57819, -38.36209, -39.14214, -39.91835, -40.69072,
  40.9524, 40.1789, 39.40136, 38.61978, 37.83415, 37.04449, 36.2508, 
    35.45309, 34.6514, 33.84572, 33.03609, 32.22254, 31.4051, 30.5838, 
    29.75869, 28.92981, 28.09721, 27.26094, 26.42107, 25.57764, 24.73074, 
    23.88042, 23.02677, 22.16986, 21.30978, 20.44661, 19.58045, 18.71139, 
    17.83953, 16.96498, 16.08784, 15.20823, 14.32627, 13.44206, 12.55573, 
    11.66742, 10.77724, 9.885328, 8.99182, 8.096853, 7.200565, 6.303097, 
    5.404592, 4.505196, 3.605054, 2.704315, 1.803126, 0.9016382, 
    1.272222e-14, -0.9016382, -1.803126, -2.704315, -3.605054, -4.505196, 
    -5.404592, -6.303097, -7.200565, -8.096853, -8.99182, -9.885328, 
    -10.77724, -11.66742, -12.55573, -13.44206, -14.32627, -15.20823, 
    -16.08784, -16.96498, -17.83953, -18.71139, -19.58045, -20.44661, 
    -21.30978, -22.16986, -23.02677, -23.88042, -24.73074, -25.57764, 
    -26.42107, -27.26094, -28.09721, -28.92981, -29.75869, -30.5838, 
    -31.4051, -32.22254, -33.03609, -33.84572, -34.6514, -35.45309, -36.2508, 
    -37.04449, -37.83415, -38.61978, -39.40136, -40.1789, -40.9524,
  41.20691, 40.43238, 39.6536, 38.87059, 38.08334, 37.29186, 36.49615, 
    35.69623, 34.89211, 34.08381, 33.27135, 32.45477, 31.63409, 30.80936, 
    29.9806, 29.14787, 28.31122, 27.47071, 26.62638, 25.77831, 24.92656, 
    24.0712, 23.21232, 22.35, 21.48432, 20.61537, 19.74325, 18.86807, 
    17.98992, 17.10892, 16.22518, 15.33881, 14.44994, 13.5587, 12.66521, 
    11.7696, 10.87202, 9.972599, 9.071482, 8.168813, 7.26474, 6.359414, 
    5.452987, 4.545611, 3.637443, 2.72864, 1.819359, 0.9097592, 1.272222e-14, 
    -0.9097592, -1.819359, -2.72864, -3.637443, -4.545611, -5.452987, 
    -6.359414, -7.26474, -8.168813, -9.071482, -9.972599, -10.87202, 
    -11.7696, -12.66521, -13.5587, -14.44994, -15.33881, -16.22518, 
    -17.10892, -17.98992, -18.86807, -19.74325, -20.61537, -21.48432, -22.35, 
    -23.21232, -24.0712, -24.92656, -25.77831, -26.62638, -27.47071, 
    -28.31122, -29.14787, -29.9806, -30.80936, -31.63409, -32.45477, 
    -33.27135, -34.08381, -34.89211, -35.69623, -36.49615, -37.29186, 
    -38.08334, -38.87059, -39.6536, -40.43238, -41.20691,
  41.45414, 40.67865, 39.89874, 39.1144, 38.32563, 37.53244, 36.73482, 
    35.9328, 35.12637, 34.31557, 33.50042, 32.68093, 31.85715, 31.02912, 
    30.19686, 29.36043, 28.51988, 27.67526, 26.82663, 25.97407, 25.11763, 
    24.2574, 23.39345, 22.52588, 21.65476, 20.7802, 19.9023, 19.02115, 
    18.13688, 17.2496, 16.35942, 15.46647, 14.57087, 13.67276, 12.77227, 
    11.86955, 10.96474, 10.05798, 9.149424, 8.239225, 7.327541, 6.414529, 
    5.50035, 4.585167, 3.669145, 2.752449, 1.835248, 0.9177083, 1.272222e-14, 
    -0.9177083, -1.835248, -2.752449, -3.669145, -4.585167, -5.50035, 
    -6.414529, -7.327541, -8.239225, -9.149424, -10.05798, -10.96474, 
    -11.86955, -12.77227, -13.67276, -14.57087, -15.46647, -16.35942, 
    -17.2496, -18.13688, -19.02115, -19.9023, -20.7802, -21.65476, -22.52588, 
    -23.39345, -24.2574, -25.11763, -25.97407, -26.82663, -27.67526, 
    -28.51988, -29.36043, -30.19686, -31.02912, -31.85715, -32.68093, 
    -33.50042, -34.31557, -35.12637, -35.9328, -36.73482, -37.53244, 
    -38.32563, -39.1144, -39.89874, -40.67865, -41.45414,
  41.69396, 40.9176, 40.13664, 39.35107, 38.56088, 37.76608, 36.96666, 
    36.16264, 35.35404, 34.54086, 33.72313, 32.90088, 32.07413, 31.24292, 
    30.4073, 29.56732, 28.72301, 27.87444, 27.02167, 26.16477, 25.3038, 
    24.43885, 23.57, 22.69734, 21.82095, 20.94095, 20.05743, 19.1705, 
    18.28028, 17.38689, 16.49044, 15.59108, 14.68893, 13.78413, 12.87683, 
    11.96717, 11.0553, 10.14138, 9.225567, 8.308019, 7.388902, 6.468383, 
    5.546633, 4.623823, 3.700126, 2.775718, 1.850776, 0.9254774, 
    1.272222e-14, -0.9254774, -1.850776, -2.775718, -3.700126, -4.623823, 
    -5.546633, -6.468383, -7.388902, -8.308019, -9.225567, -10.14138, 
    -11.0553, -11.96717, -12.87683, -13.78413, -14.68893, -15.59108, 
    -16.49044, -17.38689, -18.28028, -19.1705, -20.05743, -20.94095, 
    -21.82095, -22.69734, -23.57, -24.43885, -25.3038, -26.16477, -27.02167, 
    -27.87444, -28.72301, -29.56732, -30.4073, -31.24292, -32.07413, 
    -32.90088, -33.72313, -34.54086, -35.35404, -36.16264, -36.96666, 
    -37.76608, -38.56088, -39.35107, -40.13664, -40.9176, -41.69396,
  41.92625, 41.14911, 40.36718, 39.58046, 38.78895, 37.99264, 37.19153, 
    36.38563, 35.57495, 34.75951, 33.93933, 33.11443, 32.28485, 31.45062, 
    30.61178, 29.76838, 28.92046, 28.06809, 27.21133, 26.35024, 25.48491, 
    24.6154, 23.74181, 22.86423, 21.98275, 21.09747, 20.20851, 19.31597, 
    18.41997, 17.52065, 16.61812, 15.71253, 14.804, 13.8927, 12.97877, 
    12.06235, 11.14361, 10.22272, 9.299832, 8.375121, 7.448759, 6.520922, 
    5.591787, 4.661538, 3.730354, 2.798423, 1.865928, 0.9330581, 
    1.272222e-14, -0.9330581, -1.865928, -2.798423, -3.730354, -4.661538, 
    -5.591787, -6.520922, -7.448759, -8.375121, -9.299832, -10.22272, 
    -11.14361, -12.06235, -12.97877, -13.8927, -14.804, -15.71253, -16.61812, 
    -17.52065, -18.41997, -19.31597, -20.20851, -21.09747, -21.98275, 
    -22.86423, -23.74181, -24.6154, -25.48491, -26.35024, -27.21133, 
    -28.06809, -28.92046, -29.76838, -30.61178, -31.45062, -32.28485, 
    -33.11443, -33.93933, -34.75951, -35.57495, -36.38563, -37.19153, 
    -37.99264, -38.78895, -39.58046, -40.36718, -41.14911, -41.92625,
  42.15091, 41.37305, 40.59023, 39.80246, 39.00971, 38.21198, 37.40928, 
    36.6016, 35.78897, 34.97139, 34.14888, 33.32146, 32.48917, 31.65205, 
    30.81012, 29.96344, 29.11207, 28.25605, 27.39545, 26.53034, 25.6608, 
    24.7869, 23.90874, 23.0264, 22.13999, 21.24961, 20.35538, 19.45741, 
    18.55582, 17.65075, 16.74232, 15.83068, 14.91598, 13.99836, 13.07798, 
    12.155, 11.22959, 10.30191, 9.372141, 8.44046, 7.507047, 6.572086, 
    5.635764, 4.69827, 3.759796, 2.820537, 1.880687, 0.9404421, 1.272222e-14, 
    -0.9404421, -1.880687, -2.820537, -3.759796, -4.69827, -5.635764, 
    -6.572086, -7.507047, -8.44046, -9.372141, -10.30191, -11.22959, -12.155, 
    -13.07798, -13.99836, -14.91598, -15.83068, -16.74232, -17.65075, 
    -18.55582, -19.45741, -20.35538, -21.24961, -22.13999, -23.0264, 
    -23.90874, -24.7869, -25.6608, -26.53034, -27.39545, -28.25605, 
    -29.11207, -29.96344, -30.81012, -31.65205, -32.48917, -33.32146, 
    -34.14888, -34.97139, -35.78897, -36.6016, -37.40928, -38.21198, 
    -39.00971, -39.80246, -40.59023, -41.37305, -42.15091,
  42.36781, 41.5893, 40.80568, 40.01692, 39.22302, 38.42397, 37.61977, 
    36.81043, 35.99594, 35.17633, 34.35161, 33.5218, 32.68693, 31.84704, 
    31.00217, 30.15236, 29.29767, 28.43815, 27.57387, 26.70489, 25.8313, 
    24.95318, 24.07061, 23.18369, 22.29253, 21.39723, 20.49791, 19.59469, 
    18.68769, 17.77705, 16.86292, 15.94542, 15.02473, 14.10098, 13.17436, 
    12.24501, 11.31312, 10.37886, 9.442413, 8.503963, 7.563702, 6.621819, 
    5.678512, 4.733978, 3.788419, 2.842036, 1.895035, 0.947621, 1.272222e-14, 
    -0.947621, -1.895035, -2.842036, -3.788419, -4.733978, -5.678512, 
    -6.621819, -7.563702, -8.503963, -9.442413, -10.37886, -11.31312, 
    -12.24501, -13.17436, -14.10098, -15.02473, -15.94542, -16.86292, 
    -17.77705, -18.68769, -19.59469, -20.49791, -21.39723, -22.29253, 
    -23.18369, -24.07061, -24.95318, -25.8313, -26.70489, -27.57387, 
    -28.43815, -29.29767, -30.15236, -31.00217, -31.84704, -32.68693, 
    -33.5218, -34.35161, -35.17633, -35.99594, -36.81043, -37.61977, 
    -38.42397, -39.22302, -40.01692, -40.80568, -41.5893, -42.36781,
  42.57683, 41.79774, 41.01338, 40.22372, 39.42876, 38.62848, 37.82288, 
    37.01196, 36.19573, 35.3742, 34.54738, 33.7153, 32.87798, 32.03546, 
    31.18778, 30.33498, 29.47712, 28.61425, 27.74643, 26.87375, 25.99627, 
    25.11408, 24.22728, 23.33596, 22.44022, 21.54018, 20.63595, 19.72766, 
    18.81544, 17.89944, 16.97978, 16.05663, 15.13014, 14.20047, 13.2678, 
    12.33229, 11.39412, 10.45349, 9.510569, 8.565559, 7.618658, 6.670065, 
    5.719984, 4.768622, 3.816189, 2.862896, 1.908957, 0.9545865, 
    1.272222e-14, -0.9545865, -1.908957, -2.862896, -3.816189, -4.768622, 
    -5.719984, -6.670065, -7.618658, -8.565559, -9.510569, -10.45349, 
    -11.39412, -12.33229, -13.2678, -14.20047, -15.13014, -16.05663, 
    -16.97978, -17.89944, -18.81544, -19.72766, -20.63595, -21.54018, 
    -22.44022, -23.33596, -24.22728, -25.11408, -25.99627, -26.87375, 
    -27.74643, -28.61425, -29.47712, -30.33498, -31.18778, -32.03546, 
    -32.87798, -33.7153, -34.54738, -35.3742, -36.19573, -37.01196, 
    -37.82288, -38.62848, -39.42876, -40.22372, -41.01338, -41.79774, 
    -42.57683,
  42.77788, 41.99827, 41.21324, 40.42275, 39.6268, 38.82537, 38.01846, 
    37.20607, 36.38819, 35.56485, 34.73605, 33.90181, 33.06216, 32.21714, 
    31.36679, 30.51114, 29.65025, 28.78417, 27.91298, 27.03675, 26.15555, 
    25.26947, 24.3786, 23.48304, 22.5829, 21.6783, 20.76936, 19.85619, 
    18.93895, 18.01776, 17.09279, 16.16418, 15.2321, 14.29671, 13.3582, 
    12.41673, 11.47251, 10.52571, 9.576528, 8.625175, 7.671851, 6.716765, 
    5.760129, 4.802159, 3.843073, 2.883091, 1.922435, 0.9613302, 
    1.272222e-14, -0.9613302, -1.922435, -2.883091, -3.843073, -4.802159, 
    -5.760129, -6.716765, -7.671851, -8.625175, -9.576528, -10.52571, 
    -11.47251, -12.41673, -13.3582, -14.29671, -15.2321, -16.16418, 
    -17.09279, -18.01776, -18.93895, -19.85619, -20.76936, -21.6783, 
    -22.5829, -23.48304, -24.3786, -25.26947, -26.15555, -27.03675, 
    -27.91298, -28.78417, -29.65025, -30.51114, -31.36679, -32.21714, 
    -33.06216, -33.90181, -34.73605, -35.56485, -36.38819, -37.20607, 
    -38.01846, -38.82537, -39.6268, -40.42275, -41.21324, -41.99827, -42.77788,
  42.97084, 42.19077, 41.40512, 40.61388, 39.81702, 39.01452, 38.20639, 
    37.39261, 36.57319, 35.74813, 34.91746, 34.08119, 33.23934, 32.39194, 
    31.53904, 30.68068, 29.8169, 28.94778, 28.07337, 27.19374, 26.30898, 
    25.41917, 24.52441, 23.6248, 22.72045, 21.81147, 20.89799, 19.98014, 
    19.05806, 18.1319, 17.20181, 16.26795, 15.33048, 14.38959, 13.44545, 
    12.49824, 11.54817, 10.59543, 9.640213, 8.682739, 7.723217, 6.761864, 
    5.7989, 4.834549, 3.869038, 2.902596, 1.935454, 0.9678438, 1.272222e-14, 
    -0.9678438, -1.935454, -2.902596, -3.869038, -4.834549, -5.7989, 
    -6.761864, -7.723217, -8.682739, -9.640213, -10.59543, -11.54817, 
    -12.49824, -13.44545, -14.38959, -15.33048, -16.26795, -17.20181, 
    -18.1319, -19.05806, -19.98014, -20.89799, -21.81147, -22.72045, 
    -23.6248, -24.52441, -25.41917, -26.30898, -27.19374, -28.07337, 
    -28.94778, -29.8169, -30.68068, -31.53904, -32.39194, -33.23934, 
    -34.08119, -34.91746, -35.74813, -36.57319, -37.39261, -38.20639, 
    -39.01452, -39.81702, -40.61388, -41.40512, -42.19077, -42.97084,
  43.1556, 42.37512, 41.58892, 40.79699, 39.99928, 39.1958, 38.38652, 
    37.57145, 36.75058, 35.92393, 35.09149, 34.25329, 33.40936, 32.55971, 
    31.7044, 30.84346, 29.97694, 29.10491, 28.22743, 27.34457, 26.45642, 
    25.56305, 24.66457, 23.76108, 22.85269, 21.93953, 21.02171, 20.09937, 
    19.17266, 18.24172, 17.30672, 16.36782, 15.42518, 14.479, 13.52945, 
    12.57673, 11.62103, 10.66257, 9.701547, 8.738181, 7.772693, 6.805305, 
    5.836247, 4.865752, 3.894052, 2.921387, 1.947996, 0.9741191, 
    1.272222e-14, -0.9741191, -1.947996, -2.921387, -3.894052, -4.865752, 
    -5.836247, -6.805305, -7.772693, -8.738181, -9.701547, -10.66257, 
    -11.62103, -12.57673, -13.52945, -14.479, -15.42518, -16.36782, 
    -17.30672, -18.24172, -19.17266, -20.09937, -21.02171, -21.93953, 
    -22.85269, -23.76108, -24.66457, -25.56305, -26.45642, -27.34457, 
    -28.22743, -29.10491, -29.97694, -30.84346, -31.7044, -32.55971, 
    -33.40936, -34.25329, -35.09149, -35.92393, -36.75058, -37.57145, 
    -38.38652, -39.1958, -39.99928, -40.79699, -41.58892, -42.37512, -43.1556,
  43.33206, 42.55122, 41.76453, 40.97196, 40.17348, 39.36908, 38.55875, 
    37.74247, 36.92025, 36.09208, 35.25799, 34.41798, 33.57207, 32.7203, 
    31.86271, 30.99933, 30.13022, 29.25543, 28.37503, 27.4891, 26.59771, 
    25.70096, 24.79893, 23.89175, 22.97951, 22.06234, 21.14038, 20.21375, 
    19.28261, 18.34711, 17.4074, 16.46367, 15.51608, 14.56483, 13.61009, 
    12.65208, 11.691, 10.72705, 9.760451, 8.791431, 7.820215, 6.847034, 
    5.872125, 4.895727, 3.918083, 2.93944, 1.960045, 0.9801481, 1.272222e-14, 
    -0.9801481, -1.960045, -2.93944, -3.918083, -4.895727, -5.872125, 
    -6.847034, -7.820215, -8.791431, -9.760451, -10.72705, -11.691, 
    -12.65208, -13.61009, -14.56483, -15.51608, -16.46367, -17.4074, 
    -18.34711, -19.28261, -20.21375, -21.14038, -22.06234, -22.97951, 
    -23.89175, -24.79893, -25.70096, -26.59771, -27.4891, -28.37503, 
    -29.25543, -30.13022, -30.99933, -31.86271, -32.7203, -33.57207, 
    -34.41798, -35.25799, -36.09208, -36.92025, -37.74247, -38.55875, 
    -39.36908, -40.17348, -40.97196, -41.76453, -42.55122, -43.33206,
  43.50012, 42.71897, 41.93184, 41.13869, 40.3395, 39.53426, 38.72294, 
    37.90554, 37.08205, 36.25248, 35.41682, 34.57511, 33.72735, 32.87358, 
    32.01384, 31.14815, 30.27658, 29.39919, 28.51603, 27.62718, 26.73272, 
    25.83275, 24.92736, 24.01665, 23.10075, 22.17978, 21.25386, 20.32315, 
    19.38778, 18.44792, 17.50373, 16.55539, 15.60307, 14.64697, 13.68729, 
    12.72422, 11.75798, 10.78878, 9.816853, 8.842422, 7.865723, 6.886996, 
    5.906484, 4.924435, 3.941099, 2.956731, 1.971586, 0.9859229, 
    1.272222e-14, -0.9859229, -1.971586, -2.956731, -3.941099, -4.924435, 
    -5.906484, -6.886996, -7.865723, -8.842422, -9.816853, -10.78878, 
    -11.75798, -12.72422, -13.68729, -14.64697, -15.60307, -16.55539, 
    -17.50373, -18.44792, -19.38778, -20.32315, -21.25386, -22.17978, 
    -23.10075, -24.01665, -24.92736, -25.83275, -26.73272, -27.62718, 
    -28.51603, -29.39919, -30.27658, -31.14815, -32.01384, -32.87358, 
    -33.72735, -34.57511, -35.41682, -36.25248, -37.08205, -37.90554, 
    -38.72294, -39.53426, -40.3395, -41.13869, -41.93184, -42.71897, -43.50012,
  43.65969, 42.87827, 42.09073, 41.29707, 40.49723, 39.69121, 38.87898, 
    38.06054, 37.23587, 36.40498, 35.56787, 34.72456, 33.87507, 33.01942, 
    32.15764, 31.28979, 30.4159, 29.53604, 28.65027, 27.75867, 26.86131, 
    25.95829, 25.0497, 24.13567, 23.21629, 22.2917, 21.36204, 20.42744, 
    19.48806, 18.54405, 17.5956, 16.64287, 15.68605, 14.72534, 13.76093, 
    12.79304, 11.82189, 10.84769, 9.870676, 8.891085, 7.909157, 6.925138, 
    5.939281, 4.951838, 3.963069, 2.973237, 1.982603, 0.9914355, 
    1.272222e-14, -0.9914355, -1.982603, -2.973237, -3.963069, -4.951838, 
    -5.939281, -6.925138, -7.909157, -8.891085, -9.870676, -10.84769, 
    -11.82189, -12.79304, -13.76093, -14.72534, -15.68605, -16.64287, 
    -17.5956, -18.54405, -19.48806, -20.42744, -21.36204, -22.2917, 
    -23.21629, -24.13567, -25.0497, -25.95829, -26.86131, -27.75867, 
    -28.65027, -29.53604, -30.4159, -31.28979, -32.15764, -33.01942, 
    -33.87507, -34.72456, -35.56787, -36.40498, -37.23587, -38.06054, 
    -38.87898, -39.69121, -40.49723, -41.29707, -42.09073, -42.87827, 
    -43.65969,
  43.81068, 43.02901, 42.24112, 41.44698, 40.64656, 39.83982, 39.02676, 
    38.20735, 37.38158, 36.54947, 35.71101, 34.8662, 34.01508, 33.15767, 
    32.29399, 31.4241, 30.54803, 29.66586, 28.77763, 27.88343, 26.98333, 
    26.07744, 25.16584, 24.24865, 23.32599, 22.39799, 21.46477, 20.5265, 
    19.58331, 18.63538, 17.68288, 16.72599, 15.7649, 14.79981, 13.83093, 
    12.85847, 11.88264, 10.90369, 9.92185, 8.937356, 7.950458, 6.96141, 
    5.970469, 4.977899, 3.983964, 2.988935, 1.993082, 0.9966785, 
    1.272222e-14, -0.9966785, -1.993082, -2.988935, -3.983964, -4.977899, 
    -5.970469, -6.96141, -7.950458, -8.937356, -9.92185, -10.90369, 
    -11.88264, -12.85847, -13.83093, -14.79981, -15.7649, -16.72599, 
    -17.68288, -18.63538, -19.58331, -20.5265, -21.46477, -22.39799, 
    -23.32599, -24.24865, -25.16584, -26.07744, -26.98333, -27.88343, 
    -28.77763, -29.66586, -30.54803, -31.4241, -32.29399, -33.15767, 
    -34.01508, -34.8662, -35.71101, -36.54947, -37.38158, -38.20735, 
    -39.02676, -39.83982, -40.64656, -41.44698, -42.24112, -43.02901, 
    -43.81068,
  43.95298, 43.17111, 42.38291, 41.58834, 40.78738, 39.97999, 39.16616, 
    38.34586, 37.51908, 36.68583, 35.8461, 34.99992, 34.14728, 33.28822, 
    32.42276, 31.55096, 30.67286, 29.78851, 28.89797, 28.00133, 27.09867, 
    26.19007, 25.27564, 24.35549, 23.42973, 22.49851, 21.56195, 20.6202, 
    19.67343, 18.7218, 17.76548, 16.80466, 15.83954, 14.87031, 13.89719, 
    12.9204, 11.94017, 10.95672, 9.970306, 8.981172, 7.989569, 6.995759, 
    6.000007, 5.002581, 4.003754, 3.003803, 2.003006, 1.001644, 1.272222e-14, 
    -1.001644, -2.003006, -3.003803, -4.003754, -5.002581, -6.000007, 
    -6.995759, -7.989569, -8.981172, -9.970306, -10.95672, -11.94017, 
    -12.9204, -13.89719, -14.87031, -15.83954, -16.80466, -17.76548, 
    -18.7218, -19.67343, -20.6202, -21.56195, -22.49851, -23.42973, 
    -24.35549, -25.27564, -26.19007, -27.09867, -28.00133, -28.89797, 
    -29.78851, -30.67286, -31.55096, -32.42276, -33.28822, -34.14728, 
    -34.99992, -35.8461, -36.68583, -37.51908, -38.34586, -39.16616, 
    -39.97999, -40.78738, -41.58834, -42.38291, -43.17111, -43.95298,
  44.08652, 43.30448, 42.516, 41.72106, 40.91961, 40.11162, 39.29708, 
    38.47596, 37.64825, 36.81395, 35.97306, 35.12558, 34.27153, 33.41094, 
    32.54383, 31.67025, 30.79025, 29.90387, 29.01118, 28.11226, 27.20719, 
    26.29606, 25.37897, 24.45604, 23.52739, 22.59314, 21.65344, 20.70844, 
    19.7583, 18.80319, 17.84328, 16.87877, 15.90985, 14.93673, 13.95963, 
    12.97877, 11.99438, 11.0067, 10.01598, 9.02247, 8.026436, 7.02814, 
    6.027852, 5.025849, 4.022411, 3.017821, 2.012363, 1.006326, 1.272222e-14, 
    -1.006326, -2.012363, -3.017821, -4.022411, -5.025849, -6.027852, 
    -7.02814, -8.026436, -9.02247, -10.01598, -11.0067, -11.99438, -12.97877, 
    -13.95963, -14.93673, -15.90985, -16.87877, -17.84328, -18.80319, 
    -19.7583, -20.70844, -21.65344, -22.59314, -23.52739, -24.45604, 
    -25.37897, -26.29606, -27.20719, -28.11226, -29.01118, -29.90387, 
    -30.79025, -31.67025, -32.54383, -33.41094, -34.27153, -35.12558, 
    -35.97306, -36.81395, -37.64825, -38.47596, -39.29708, -40.11162, 
    -40.91961, -41.72106, -42.516, -43.30448, -44.08652,
  44.21122, 43.42903, 42.64032, 41.84503, 41.04314, 40.23461, 39.41943, 
    38.59755, 37.76899, 36.93372, 36.09175, 35.24308, 34.38773, 33.52573, 
    32.65709, 31.78186, 30.90008, 30.01182, 29.11712, 28.21608, 27.30877, 
    26.39529, 25.47573, 24.55021, 23.61885, 22.68178, 21.73915, 20.79111, 
    19.83782, 18.87945, 17.91618, 16.94822, 15.97575, 14.99899, 14.01815, 
    13.03348, 12.0452, 11.05355, 10.0588, 9.061195, 8.061007, 7.058504, 
    6.053965, 5.047671, 4.039908, 3.030967, 2.021138, 1.010717, 1.272222e-14, 
    -1.010717, -2.021138, -3.030967, -4.039908, -5.047671, -6.053965, 
    -7.058504, -8.061007, -9.061195, -10.0588, -11.05355, -12.0452, 
    -13.03348, -14.01815, -14.99899, -15.97575, -16.94822, -17.91618, 
    -18.87945, -19.83782, -20.79111, -21.73915, -22.68178, -23.61885, 
    -24.55021, -25.47573, -26.39529, -27.30877, -28.21608, -29.11712, 
    -30.01182, -30.90008, -31.78186, -32.65709, -33.52573, -34.38773, 
    -35.24308, -36.09175, -36.93372, -37.76899, -38.59755, -39.41943, 
    -40.23461, -41.04314, -41.84503, -42.64032, -43.42903, -44.21122,
  44.32701, 43.54469, 42.75576, 41.96017, 41.15789, 40.34887, 39.5331, 
    38.71054, 37.8812, 37.04504, 36.20208, 35.35233, 34.49578, 33.63246, 
    32.76241, 31.88566, 31.00225, 30.11224, 29.2157, 28.3127, 27.40331, 
    26.48764, 25.56579, 24.63787, 23.704, 22.76431, 21.81896, 20.8681, 
    19.91188, 18.95048, 17.9841, 17.01292, 16.03714, 15.05699, 14.07269, 
    13.08447, 12.09256, 11.09722, 10.09871, 9.097291, 8.09323, 7.086808, 
    6.078306, 5.068013, 4.05622, 3.043222, 2.029319, 1.014811, 1.272222e-14, 
    -1.014811, -2.029319, -3.043222, -4.05622, -5.068013, -6.078306, 
    -7.086808, -8.09323, -9.097291, -10.09871, -11.09722, -12.09256, 
    -13.08447, -14.07269, -15.05699, -16.03714, -17.01292, -17.9841, 
    -18.95048, -19.91188, -20.8681, -21.81896, -22.76431, -23.704, -24.63787, 
    -25.56579, -26.48764, -27.40331, -28.3127, -29.2157, -30.11224, 
    -31.00225, -31.88566, -32.76241, -33.63246, -34.49578, -35.35233, 
    -36.20208, -37.04504, -37.8812, -38.71054, -39.5331, -40.34887, 
    -41.15789, -41.96017, -42.75576, -43.54469, -44.32701,
  44.4338, 43.65138, 42.86227, 42.06641, 41.26377, 40.45432, 39.63801, 
    38.81484, 37.98478, 37.14782, 36.30396, 35.45321, 34.59556, 33.73105, 
    32.85971, 31.98156, 31.09665, 30.20505, 29.3068, 28.40199, 27.4907, 
    26.57302, 25.64905, 24.71892, 23.78273, 22.84064, 21.89278, 20.9393, 
    19.98038, 19.0162, 18.04693, 17.07278, 16.09396, 15.11067, 14.12316, 
    13.13165, 12.1364, 11.13764, 10.13566, 9.130703, 8.123061, 7.113011, 
    6.100842, 5.086846, 4.071321, 3.054569, 2.036894, 1.018601, 1.272222e-14, 
    -1.018601, -2.036894, -3.054569, -4.071321, -5.086846, -6.100842, 
    -7.113011, -8.123061, -9.130703, -10.13566, -11.13764, -12.1364, 
    -13.13165, -14.12316, -15.11067, -16.09396, -17.07278, -18.04693, 
    -19.0162, -19.98038, -20.9393, -21.89278, -22.84064, -23.78273, 
    -24.71892, -25.64905, -26.57302, -27.4907, -28.40199, -29.3068, 
    -30.20505, -31.09665, -31.98156, -32.85971, -33.73105, -34.59556, 
    -35.45321, -36.30396, -37.14782, -37.98478, -38.81484, -39.63801, 
    -40.45432, -41.26377, -42.06641, -42.86227, -43.65138, -44.4338,
  44.53154, 43.74903, 42.95976, 42.16367, 41.36071, 40.55087, 39.73409, 
    38.91036, 38.07965, 37.24197, 36.39729, 35.54563, 34.68699, 33.8214, 
    32.94887, 32.06945, 31.18319, 30.29012, 29.39032, 28.48387, 27.57083, 
    26.65132, 25.72542, 24.79326, 23.85496, 22.91066, 21.9605, 21.00464, 
    20.04325, 19.0765, 18.1046, 17.12773, 16.1461, 15.15995, 14.16949, 
    13.17497, 12.17664, 11.17476, 10.16958, 9.161384, 8.150454, 7.137073, 
    6.121536, 5.104141, 4.08519, 3.06499, 2.04385, 1.022082, 1.272222e-14, 
    -1.022082, -2.04385, -3.06499, -4.08519, -5.104141, -6.121536, -7.137073, 
    -8.150454, -9.161384, -10.16958, -11.17476, -12.17664, -13.17497, 
    -14.16949, -15.15995, -16.1461, -17.12773, -18.1046, -19.0765, -20.04325, 
    -21.00464, -21.9605, -22.91066, -23.85496, -24.79326, -25.72542, 
    -26.65132, -27.57083, -28.48387, -29.39032, -30.29012, -31.18319, 
    -32.06945, -32.94887, -33.8214, -34.68699, -35.54563, -36.39729, 
    -37.24197, -38.07965, -38.91036, -39.73409, -40.55087, -41.36071, 
    -42.16367, -42.95976, -43.74903, -44.53154,
  44.62016, 43.83758, 43.04817, 42.25187, 41.44865, 40.63845, 39.82125, 
    38.99702, 38.16574, 37.3274, 36.48199, 35.62952, 34.76999, 33.90341, 
    33.02983, 32.14926, 31.26176, 30.36738, 29.46618, 28.55823, 27.64362, 
    26.72244, 25.7948, 24.86081, 23.92059, 22.97429, 22.02205, 21.06402, 
    20.10039, 19.13132, 18.15702, 17.17768, 16.19351, 15.20475, 14.21162, 
    13.21437, 12.21324, 11.2085, 10.20043, 9.189286, 8.175366, 7.158958, 
    6.140359, 5.119872, 4.097805, 3.074468, 2.050177, 1.025248, 1.272222e-14, 
    -1.025248, -2.050177, -3.074468, -4.097805, -5.119872, -6.140359, 
    -7.158958, -8.175366, -9.189286, -10.20043, -11.2085, -12.21324, 
    -13.21437, -14.21162, -15.20475, -16.19351, -17.17768, -18.15702, 
    -19.13132, -20.10039, -21.06402, -22.02205, -22.97429, -23.92059, 
    -24.86081, -25.7948, -26.72244, -27.64362, -28.55823, -29.46618, 
    -30.36738, -31.26176, -32.14926, -33.02983, -33.90341, -34.76999, 
    -35.62952, -36.48199, -37.3274, -38.16574, -38.99702, -39.82125, 
    -40.63845, -41.44865, -42.25187, -43.04817, -43.83758, -44.62016,
  44.6996, 43.91697, 43.12745, 42.33097, 41.5275, 40.717, 39.89942, 39.07475, 
    38.24297, 37.40405, 36.55799, 35.70479, 34.84446, 33.97701, 33.10248, 
    32.22089, 31.33229, 30.43673, 29.53428, 28.625, 27.70898, 26.78632, 
    25.85711, 24.92148, 23.97954, 23.03145, 22.07734, 21.11737, 20.15172, 
    19.18058, 18.20412, 17.22256, 16.23612, 15.24501, 14.24948, 13.24977, 
    12.24614, 11.23884, 10.22816, 9.21437, 8.197762, 7.178632, 6.157281, 
    5.134015, 4.109146, 3.08299, 2.055866, 1.028095, 1.272222e-14, -1.028095, 
    -2.055866, -3.08299, -4.109146, -5.134015, -6.157281, -7.178632, 
    -8.197762, -9.21437, -10.22816, -11.23884, -12.24614, -13.24977, 
    -14.24948, -15.24501, -16.23612, -17.22256, -18.20412, -19.18058, 
    -20.15172, -21.11737, -22.07734, -23.03145, -23.97954, -24.92148, 
    -25.85711, -26.78632, -27.70898, -28.625, -29.53428, -30.43673, 
    -31.33229, -32.22089, -33.10248, -33.97701, -34.84446, -35.70479, 
    -36.55799, -37.40405, -38.24297, -39.07475, -39.89942, -40.717, -41.5275, 
    -42.33097, -43.12745, -43.91697, -44.6996,
  44.76982, 43.98714, 43.19752, 42.40089, 41.59722, 40.78645, 39.96855, 
    39.1435, 38.31126, 37.47184, 36.62521, 35.77137, 34.91034, 34.04213, 
    33.16676, 32.28428, 31.39471, 30.49811, 29.59455, 28.6841, 27.76684, 
    26.84286, 25.91227, 24.97519, 24.03174, 23.08206, 22.1263, 21.16462, 
    20.19719, 19.2242, 18.24584, 17.26232, 16.27386, 15.28068, 14.28303, 
    13.28114, 12.27528, 11.26572, 10.25273, 9.236594, 8.217607, 7.196066, 
    6.172276, 5.146547, 4.119196, 3.090542, 2.060907, 1.030618, 1.272222e-14, 
    -1.030618, -2.060907, -3.090542, -4.119196, -5.146547, -6.172276, 
    -7.196066, -8.217607, -9.236594, -10.25273, -11.26572, -12.27528, 
    -13.28114, -14.28303, -15.28068, -16.27386, -17.26232, -18.24584, 
    -19.2242, -20.19719, -21.16462, -22.1263, -23.08206, -24.03174, 
    -24.97519, -25.91227, -26.84286, -27.76684, -28.6841, -29.59455, 
    -30.49811, -31.39471, -32.28428, -33.16676, -34.04213, -34.91034, 
    -35.77137, -36.62521, -37.47184, -38.31126, -39.1435, -39.96855, 
    -40.78645, -41.59722, -42.40089, -43.19752, -43.98714, -44.76982,
  44.83077, 44.04806, 43.25835, 42.4616, 41.65775, 40.84675, 40.02857, 
    39.20319, 38.37057, 37.53071, 36.68359, 35.8292, 34.96757, 34.0987, 
    33.22261, 32.33934, 31.44894, 30.55145, 29.64693, 28.73546, 27.81712, 
    26.892, 25.96022, 25.02188, 24.07711, 23.12605, 22.16886, 21.20569, 
    20.23672, 19.26213, 18.28212, 17.2969, 16.30668, 15.3117, 14.3122, 
    13.30842, 12.30063, 11.2891, 10.2741, 9.255927, 8.23487, 7.211231, 
    6.18532, 5.15745, 4.127939, 3.097111, 2.065293, 1.032812, 1.272222e-14, 
    -1.032812, -2.065293, -3.097111, -4.127939, -5.15745, -6.18532, 
    -7.211231, -8.23487, -9.255927, -10.2741, -11.2891, -12.30063, -13.30842, 
    -14.3122, -15.3117, -16.30668, -17.2969, -18.28212, -19.26213, -20.23672, 
    -21.20569, -22.16886, -23.12605, -24.07711, -25.02188, -25.96022, 
    -26.892, -27.81712, -28.73546, -29.64693, -30.55145, -31.44894, 
    -32.33934, -33.22261, -34.0987, -34.96757, -35.8292, -36.68359, 
    -37.53071, -38.37057, -39.20319, -40.02857, -40.84675, -41.65775, 
    -42.4616, -43.25835, -44.04806, -44.83077,
  44.88241, 44.09967, 43.3099, 42.51304, 41.70904, 40.89785, 40.07944, 
    39.25378, 38.42085, 37.58062, 36.73308, 35.87823, 35.01609, 34.14666, 
    33.26997, 32.38604, 31.49493, 30.59668, 29.69135, 28.77902, 27.85977, 
    26.93369, 26.00089, 25.06149, 24.1156, 23.16338, 22.20498, 21.24054, 
    20.27026, 19.29432, 18.31291, 17.32624, 16.33454, 15.33803, 14.33696, 
    13.33158, 12.32215, 11.30894, 10.29224, 9.272337, 8.249522, 7.224104, 
    6.196393, 5.166705, 4.135361, 3.102689, 2.069016, 1.034675, 1.272222e-14, 
    -1.034675, -2.069016, -3.102689, -4.135361, -5.166705, -6.196393, 
    -7.224104, -8.249522, -9.272337, -10.29224, -11.30894, -12.32215, 
    -13.33158, -14.33696, -15.33803, -16.33454, -17.32624, -18.31291, 
    -19.29432, -20.27026, -21.24054, -22.20498, -23.16338, -24.1156, 
    -25.06149, -26.00089, -26.93369, -27.85977, -28.77902, -29.69135, 
    -30.59668, -31.49493, -32.38604, -33.26997, -34.14666, -35.01609, 
    -35.87823, -36.73308, -37.58062, -38.42085, -39.25378, -40.07944, 
    -40.89785, -41.70904, -42.51304, -43.3099, -44.09967, -44.88241,
  44.9247, 44.14195, 43.35213, 42.55518, 41.75106, 40.93972, 40.12112, 
    39.29524, 38.46204, 37.62151, 36.77364, 35.91842, 35.05586, 34.18597, 
    33.30878, 32.42432, 31.53263, 30.63375, 29.72776, 28.81473, 27.89473, 
    26.96786, 26.03424, 25.09396, 24.14717, 23.19399, 22.23459, 21.26912, 
    20.29777, 19.32071, 18.33815, 17.3503, 16.35738, 15.35962, 14.35726, 
    13.35057, 12.3398, 11.32522, 10.30712, 9.285798, 8.261543, 7.234665, 
    6.205477, 5.174297, 4.14145, 3.107264, 2.07207, 1.036204, 1.272222e-14, 
    -1.036204, -2.07207, -3.107264, -4.14145, -5.174297, -6.205477, 
    -7.234665, -8.261543, -9.285798, -10.30712, -11.32522, -12.3398, 
    -13.35057, -14.35726, -15.35962, -16.35738, -17.3503, -18.33815, 
    -19.32071, -20.29777, -21.26912, -22.23459, -23.19399, -24.14717, 
    -25.09396, -26.03424, -26.96786, -27.89473, -28.81473, -29.72776, 
    -30.63375, -31.53263, -32.42432, -33.30878, -34.18597, -35.05586, 
    -35.91842, -36.77364, -37.62151, -38.46204, -39.29524, -40.12112, 
    -40.93972, -41.75106, -42.55518, -43.35213, -44.14195, -44.9247,
  44.95763, 44.17486, 43.385, 42.58799, 41.78378, 40.97232, 40.15358, 
    39.32752, 38.49412, 37.65335, 36.80522, 35.94971, 35.08683, 34.21658, 
    33.33901, 32.45413, 31.56199, 30.66263, 29.75613, 28.84255, 27.92197, 
    26.99449, 26.06021, 25.11926, 24.17175, 23.21784, 22.25766, 21.29139, 
    20.3192, 19.34128, 18.35783, 17.36906, 16.37519, 15.37645, 14.37309, 
    13.36537, 12.35355, 11.33791, 10.31872, 9.29629, 8.270913, 7.242897, 
    6.212557, 5.180215, 4.146196, 3.11083, 2.074451, 1.037395, 1.272222e-14, 
    -1.037395, -2.074451, -3.11083, -4.146196, -5.180215, -6.212557, 
    -7.242897, -8.270913, -9.29629, -10.31872, -11.33791, -12.35355, 
    -13.36537, -14.37309, -15.37645, -16.37519, -17.36906, -18.35783, 
    -19.34128, -20.3192, -21.29139, -22.25766, -23.21784, -24.17175, 
    -25.11926, -26.06021, -26.99449, -27.92197, -28.84255, -29.75613, 
    -30.66263, -31.56199, -32.45413, -33.33901, -34.21658, -35.08683, 
    -35.94971, -36.80522, -37.65335, -38.49412, -39.32752, -40.15358, 
    -40.97232, -41.78378, -42.58799, -43.385, -44.17486, -44.95763,
  44.98116, 44.19839, 43.4085, 42.61144, 41.80717, 40.99562, 40.17678, 
    39.3506, 38.51705, 37.67612, 36.8278, 35.97208, 35.10897, 34.23848, 
    33.36062, 32.47544, 31.58298, 30.68328, 29.77641, 28.86244, 27.94145, 
    27.01353, 26.0788, 25.13736, 24.18934, 23.2349, 22.27417, 21.30732, 
    20.33454, 19.356, 18.3719, 17.38247, 16.38792, 15.38849, 14.38441, 
    13.37596, 12.36339, 11.34698, 10.32702, 9.303797, 8.277617, 7.248786, 
    6.217623, 5.184449, 4.149592, 3.113382, 2.076154, 1.038247, 1.272222e-14, 
    -1.038247, -2.076154, -3.113382, -4.149592, -5.184449, -6.217623, 
    -7.248786, -8.277617, -9.303797, -10.32702, -11.34698, -12.36339, 
    -13.37596, -14.38441, -15.38849, -16.38792, -17.38247, -18.3719, -19.356, 
    -20.33454, -21.30732, -22.27417, -23.2349, -24.18934, -25.13736, 
    -26.0788, -27.01353, -27.94145, -28.86244, -29.77641, -30.68328, 
    -31.58298, -32.47544, -33.36062, -34.23848, -35.10897, -35.97208, 
    -36.8278, -37.67612, -38.51705, -39.3506, -40.17678, -40.99562, 
    -41.80717, -42.61144, -43.4085, -44.19839, -44.98116,
  44.99529, 44.21251, 43.4226, 42.62552, 41.82121, 41.00961, 40.1907, 
    39.36445, 38.53082, 37.68979, 36.84136, 35.98551, 35.12226, 34.25162, 
    33.3736, 32.48825, 31.59559, 30.69568, 29.78859, 28.87439, 27.95315, 
    27.02497, 26.08995, 25.14822, 24.19991, 23.24514, 22.28408, 21.31689, 
    20.34374, 19.36483, 18.38036, 17.39053, 16.39557, 15.39572, 14.39121, 
    13.38232, 12.3693, 11.35243, 10.332, 9.308306, 8.281642, 7.252323, 
    6.220666, 5.186993, 4.151631, 3.114914, 2.077178, 1.038759, 1.272222e-14, 
    -1.038759, -2.077178, -3.114914, -4.151631, -5.186993, -6.220666, 
    -7.252323, -8.281642, -9.308306, -10.332, -11.35243, -12.3693, -13.38232, 
    -14.39121, -15.39572, -16.39557, -17.39053, -18.38036, -19.36483, 
    -20.34374, -21.31689, -22.28408, -23.24514, -24.19991, -25.14822, 
    -26.08995, -27.02497, -27.95315, -28.87439, -29.78859, -30.69568, 
    -31.59559, -32.48825, -33.3736, -34.25162, -35.12226, -35.98551, 
    -36.84136, -37.68979, -38.53082, -39.36445, -40.1907, -41.00961, 
    -41.82121, -42.62552, -43.4226, -44.21251, -44.99529,
  45, 44.21722, 43.42731, 42.63021, 41.82589, 41.01428, 40.19535, 39.36907, 
    38.53541, 37.69435, 36.84588, 35.98999, 35.12669, 34.256, 33.37793, 
    32.49251, 31.59979, 30.69982, 29.79265, 28.87837, 27.95705, 27.02878, 
    26.09367, 25.15185, 24.20343, 23.24856, 22.28739, 21.32008, 20.34682, 
    19.36778, 18.38318, 17.39322, 16.39812, 15.39813, 14.39348, 13.38444, 
    12.37127, 11.35425, 10.33367, 9.30981, 8.282985, 7.253503, 6.221681, 
    5.187841, 4.152311, 3.115426, 2.077519, 1.03893, 1.272222e-14, -1.03893, 
    -2.077519, -3.115426, -4.152311, -5.187841, -6.221681, -7.253503, 
    -8.282985, -9.30981, -10.33367, -11.35425, -12.37127, -13.38444, 
    -14.39348, -15.39813, -16.39812, -17.39322, -18.38318, -19.36778, 
    -20.34682, -21.32008, -22.28739, -23.24856, -24.20343, -25.15185, 
    -26.09367, -27.02878, -27.95705, -28.87837, -29.79265, -30.69982, 
    -31.59979, -32.49251, -33.37793, -34.256, -35.12669, -35.98999, 
    -36.84588, -37.69435, -38.53541, -39.36907, -40.19535, -41.01428, 
    -41.82589, -42.63021, -43.42731, -44.21722, -45,
  44.99529, 44.21251, 43.4226, 42.62552, 41.82121, 41.00961, 40.1907, 
    39.36445, 38.53082, 37.68979, 36.84136, 35.98551, 35.12226, 34.25162, 
    33.3736, 32.48825, 31.59559, 30.69568, 29.78859, 28.87439, 27.95315, 
    27.02497, 26.08995, 25.14822, 24.19991, 23.24514, 22.28408, 21.31689, 
    20.34374, 19.36483, 18.38036, 17.39053, 16.39557, 15.39572, 14.39121, 
    13.38232, 12.3693, 11.35243, 10.332, 9.308306, 8.281642, 7.252323, 
    6.220666, 5.186993, 4.151631, 3.114914, 2.077178, 1.038759, 1.272222e-14, 
    -1.038759, -2.077178, -3.114914, -4.151631, -5.186993, -6.220666, 
    -7.252323, -8.281642, -9.308306, -10.332, -11.35243, -12.3693, -13.38232, 
    -14.39121, -15.39572, -16.39557, -17.39053, -18.38036, -19.36483, 
    -20.34374, -21.31689, -22.28408, -23.24514, -24.19991, -25.14822, 
    -26.08995, -27.02497, -27.95315, -28.87439, -29.78859, -30.69568, 
    -31.59559, -32.48825, -33.3736, -34.25162, -35.12226, -35.98551, 
    -36.84136, -37.68979, -38.53082, -39.36445, -40.1907, -41.00961, 
    -41.82121, -42.62552, -43.4226, -44.21251, -44.99529,
  44.98116, 44.19839, 43.4085, 42.61144, 41.80717, 40.99562, 40.17678, 
    39.3506, 38.51705, 37.67612, 36.8278, 35.97208, 35.10897, 34.23848, 
    33.36062, 32.47544, 31.58298, 30.68328, 29.77641, 28.86244, 27.94145, 
    27.01353, 26.0788, 25.13736, 24.18934, 23.2349, 22.27417, 21.30732, 
    20.33454, 19.356, 18.3719, 17.38247, 16.38792, 15.38849, 14.38441, 
    13.37596, 12.36339, 11.34698, 10.32702, 9.303797, 8.277617, 7.248786, 
    6.217623, 5.184449, 4.149592, 3.113382, 2.076154, 1.038247, 1.272222e-14, 
    -1.038247, -2.076154, -3.113382, -4.149592, -5.184449, -6.217623, 
    -7.248786, -8.277617, -9.303797, -10.32702, -11.34698, -12.36339, 
    -13.37596, -14.38441, -15.38849, -16.38792, -17.38247, -18.3719, -19.356, 
    -20.33454, -21.30732, -22.27417, -23.2349, -24.18934, -25.13736, 
    -26.0788, -27.01353, -27.94145, -28.86244, -29.77641, -30.68328, 
    -31.58298, -32.47544, -33.36062, -34.23848, -35.10897, -35.97208, 
    -36.8278, -37.67612, -38.51705, -39.3506, -40.17678, -40.99562, 
    -41.80717, -42.61144, -43.4085, -44.19839, -44.98116,
  44.95763, 44.17486, 43.385, 42.58799, 41.78378, 40.97232, 40.15358, 
    39.32752, 38.49412, 37.65335, 36.80522, 35.94971, 35.08683, 34.21658, 
    33.33901, 32.45413, 31.56199, 30.66263, 29.75613, 28.84255, 27.92197, 
    26.99449, 26.06021, 25.11926, 24.17175, 23.21784, 22.25766, 21.29139, 
    20.3192, 19.34128, 18.35783, 17.36906, 16.37519, 15.37645, 14.37309, 
    13.36537, 12.35355, 11.33791, 10.31872, 9.29629, 8.270913, 7.242897, 
    6.212557, 5.180215, 4.146196, 3.11083, 2.074451, 1.037395, 1.272222e-14, 
    -1.037395, -2.074451, -3.11083, -4.146196, -5.180215, -6.212557, 
    -7.242897, -8.270913, -9.29629, -10.31872, -11.33791, -12.35355, 
    -13.36537, -14.37309, -15.37645, -16.37519, -17.36906, -18.35783, 
    -19.34128, -20.3192, -21.29139, -22.25766, -23.21784, -24.17175, 
    -25.11926, -26.06021, -26.99449, -27.92197, -28.84255, -29.75613, 
    -30.66263, -31.56199, -32.45413, -33.33901, -34.21658, -35.08683, 
    -35.94971, -36.80522, -37.65335, -38.49412, -39.32752, -40.15358, 
    -40.97232, -41.78378, -42.58799, -43.385, -44.17486, -44.95763,
  44.9247, 44.14195, 43.35213, 42.55518, 41.75106, 40.93972, 40.12112, 
    39.29524, 38.46204, 37.62151, 36.77364, 35.91842, 35.05586, 34.18597, 
    33.30878, 32.42432, 31.53263, 30.63375, 29.72776, 28.81473, 27.89473, 
    26.96786, 26.03424, 25.09396, 24.14717, 23.19399, 22.23459, 21.26912, 
    20.29777, 19.32071, 18.33815, 17.3503, 16.35738, 15.35962, 14.35726, 
    13.35057, 12.3398, 11.32522, 10.30712, 9.285798, 8.261543, 7.234665, 
    6.205477, 5.174297, 4.14145, 3.107264, 2.07207, 1.036204, 1.272222e-14, 
    -1.036204, -2.07207, -3.107264, -4.14145, -5.174297, -6.205477, 
    -7.234665, -8.261543, -9.285798, -10.30712, -11.32522, -12.3398, 
    -13.35057, -14.35726, -15.35962, -16.35738, -17.3503, -18.33815, 
    -19.32071, -20.29777, -21.26912, -22.23459, -23.19399, -24.14717, 
    -25.09396, -26.03424, -26.96786, -27.89473, -28.81473, -29.72776, 
    -30.63375, -31.53263, -32.42432, -33.30878, -34.18597, -35.05586, 
    -35.91842, -36.77364, -37.62151, -38.46204, -39.29524, -40.12112, 
    -40.93972, -41.75106, -42.55518, -43.35213, -44.14195, -44.9247,
  44.88241, 44.09967, 43.3099, 42.51304, 41.70904, 40.89785, 40.07944, 
    39.25378, 38.42085, 37.58062, 36.73308, 35.87823, 35.01609, 34.14666, 
    33.26997, 32.38604, 31.49493, 30.59668, 29.69135, 28.77902, 27.85977, 
    26.93369, 26.00089, 25.06149, 24.1156, 23.16338, 22.20498, 21.24054, 
    20.27026, 19.29432, 18.31291, 17.32624, 16.33454, 15.33803, 14.33696, 
    13.33158, 12.32215, 11.30894, 10.29224, 9.272337, 8.249522, 7.224104, 
    6.196393, 5.166705, 4.135361, 3.102689, 2.069016, 1.034675, 1.272222e-14, 
    -1.034675, -2.069016, -3.102689, -4.135361, -5.166705, -6.196393, 
    -7.224104, -8.249522, -9.272337, -10.29224, -11.30894, -12.32215, 
    -13.33158, -14.33696, -15.33803, -16.33454, -17.32624, -18.31291, 
    -19.29432, -20.27026, -21.24054, -22.20498, -23.16338, -24.1156, 
    -25.06149, -26.00089, -26.93369, -27.85977, -28.77902, -29.69135, 
    -30.59668, -31.49493, -32.38604, -33.26997, -34.14666, -35.01609, 
    -35.87823, -36.73308, -37.58062, -38.42085, -39.25378, -40.07944, 
    -40.89785, -41.70904, -42.51304, -43.3099, -44.09967, -44.88241,
  44.83077, 44.04806, 43.25835, 42.4616, 41.65775, 40.84675, 40.02857, 
    39.20319, 38.37057, 37.53071, 36.68359, 35.8292, 34.96757, 34.0987, 
    33.22261, 32.33934, 31.44894, 30.55145, 29.64693, 28.73546, 27.81712, 
    26.892, 25.96022, 25.02188, 24.07711, 23.12605, 22.16886, 21.20569, 
    20.23672, 19.26213, 18.28212, 17.2969, 16.30668, 15.3117, 14.3122, 
    13.30842, 12.30063, 11.2891, 10.2741, 9.255927, 8.23487, 7.211231, 
    6.18532, 5.15745, 4.127939, 3.097111, 2.065293, 1.032812, 1.272222e-14, 
    -1.032812, -2.065293, -3.097111, -4.127939, -5.15745, -6.18532, 
    -7.211231, -8.23487, -9.255927, -10.2741, -11.2891, -12.30063, -13.30842, 
    -14.3122, -15.3117, -16.30668, -17.2969, -18.28212, -19.26213, -20.23672, 
    -21.20569, -22.16886, -23.12605, -24.07711, -25.02188, -25.96022, 
    -26.892, -27.81712, -28.73546, -29.64693, -30.55145, -31.44894, 
    -32.33934, -33.22261, -34.0987, -34.96757, -35.8292, -36.68359, 
    -37.53071, -38.37057, -39.20319, -40.02857, -40.84675, -41.65775, 
    -42.4616, -43.25835, -44.04806, -44.83077,
  44.76982, 43.98714, 43.19752, 42.40089, 41.59722, 40.78645, 39.96855, 
    39.1435, 38.31126, 37.47184, 36.62521, 35.77137, 34.91034, 34.04213, 
    33.16676, 32.28428, 31.39471, 30.49811, 29.59455, 28.6841, 27.76684, 
    26.84286, 25.91227, 24.97519, 24.03174, 23.08206, 22.1263, 21.16462, 
    20.19719, 19.2242, 18.24584, 17.26232, 16.27386, 15.28068, 14.28303, 
    13.28114, 12.27528, 11.26572, 10.25273, 9.236594, 8.217607, 7.196066, 
    6.172276, 5.146547, 4.119196, 3.090542, 2.060907, 1.030618, 1.272222e-14, 
    -1.030618, -2.060907, -3.090542, -4.119196, -5.146547, -6.172276, 
    -7.196066, -8.217607, -9.236594, -10.25273, -11.26572, -12.27528, 
    -13.28114, -14.28303, -15.28068, -16.27386, -17.26232, -18.24584, 
    -19.2242, -20.19719, -21.16462, -22.1263, -23.08206, -24.03174, 
    -24.97519, -25.91227, -26.84286, -27.76684, -28.6841, -29.59455, 
    -30.49811, -31.39471, -32.28428, -33.16676, -34.04213, -34.91034, 
    -35.77137, -36.62521, -37.47184, -38.31126, -39.1435, -39.96855, 
    -40.78645, -41.59722, -42.40089, -43.19752, -43.98714, -44.76982,
  44.6996, 43.91697, 43.12745, 42.33097, 41.5275, 40.717, 39.89942, 39.07475, 
    38.24297, 37.40405, 36.55799, 35.70479, 34.84446, 33.97701, 33.10248, 
    32.22089, 31.33229, 30.43673, 29.53428, 28.625, 27.70898, 26.78632, 
    25.85711, 24.92148, 23.97954, 23.03145, 22.07734, 21.11737, 20.15172, 
    19.18058, 18.20412, 17.22256, 16.23612, 15.24501, 14.24948, 13.24977, 
    12.24614, 11.23884, 10.22816, 9.21437, 8.197762, 7.178632, 6.157281, 
    5.134015, 4.109146, 3.08299, 2.055866, 1.028095, 1.272222e-14, -1.028095, 
    -2.055866, -3.08299, -4.109146, -5.134015, -6.157281, -7.178632, 
    -8.197762, -9.21437, -10.22816, -11.23884, -12.24614, -13.24977, 
    -14.24948, -15.24501, -16.23612, -17.22256, -18.20412, -19.18058, 
    -20.15172, -21.11737, -22.07734, -23.03145, -23.97954, -24.92148, 
    -25.85711, -26.78632, -27.70898, -28.625, -29.53428, -30.43673, 
    -31.33229, -32.22089, -33.10248, -33.97701, -34.84446, -35.70479, 
    -36.55799, -37.40405, -38.24297, -39.07475, -39.89942, -40.717, -41.5275, 
    -42.33097, -43.12745, -43.91697, -44.6996,
  44.62016, 43.83758, 43.04817, 42.25187, 41.44865, 40.63845, 39.82125, 
    38.99702, 38.16574, 37.3274, 36.48199, 35.62952, 34.76999, 33.90341, 
    33.02983, 32.14926, 31.26176, 30.36738, 29.46618, 28.55823, 27.64362, 
    26.72244, 25.7948, 24.86081, 23.92059, 22.97429, 22.02205, 21.06402, 
    20.10039, 19.13132, 18.15702, 17.17768, 16.19351, 15.20475, 14.21162, 
    13.21437, 12.21324, 11.2085, 10.20043, 9.189286, 8.175366, 7.158958, 
    6.140359, 5.119872, 4.097805, 3.074468, 2.050177, 1.025248, 1.272222e-14, 
    -1.025248, -2.050177, -3.074468, -4.097805, -5.119872, -6.140359, 
    -7.158958, -8.175366, -9.189286, -10.20043, -11.2085, -12.21324, 
    -13.21437, -14.21162, -15.20475, -16.19351, -17.17768, -18.15702, 
    -19.13132, -20.10039, -21.06402, -22.02205, -22.97429, -23.92059, 
    -24.86081, -25.7948, -26.72244, -27.64362, -28.55823, -29.46618, 
    -30.36738, -31.26176, -32.14926, -33.02983, -33.90341, -34.76999, 
    -35.62952, -36.48199, -37.3274, -38.16574, -38.99702, -39.82125, 
    -40.63845, -41.44865, -42.25187, -43.04817, -43.83758, -44.62016,
  44.53154, 43.74903, 42.95976, 42.16367, 41.36071, 40.55087, 39.73409, 
    38.91036, 38.07965, 37.24197, 36.39729, 35.54563, 34.68699, 33.8214, 
    32.94887, 32.06945, 31.18319, 30.29012, 29.39032, 28.48387, 27.57083, 
    26.65132, 25.72542, 24.79326, 23.85496, 22.91066, 21.9605, 21.00464, 
    20.04325, 19.0765, 18.1046, 17.12773, 16.1461, 15.15995, 14.16949, 
    13.17497, 12.17664, 11.17476, 10.16958, 9.161384, 8.150454, 7.137073, 
    6.121536, 5.104141, 4.08519, 3.06499, 2.04385, 1.022082, 1.272222e-14, 
    -1.022082, -2.04385, -3.06499, -4.08519, -5.104141, -6.121536, -7.137073, 
    -8.150454, -9.161384, -10.16958, -11.17476, -12.17664, -13.17497, 
    -14.16949, -15.15995, -16.1461, -17.12773, -18.1046, -19.0765, -20.04325, 
    -21.00464, -21.9605, -22.91066, -23.85496, -24.79326, -25.72542, 
    -26.65132, -27.57083, -28.48387, -29.39032, -30.29012, -31.18319, 
    -32.06945, -32.94887, -33.8214, -34.68699, -35.54563, -36.39729, 
    -37.24197, -38.07965, -38.91036, -39.73409, -40.55087, -41.36071, 
    -42.16367, -42.95976, -43.74903, -44.53154,
  44.4338, 43.65138, 42.86227, 42.06641, 41.26377, 40.45432, 39.63801, 
    38.81484, 37.98478, 37.14782, 36.30396, 35.45321, 34.59556, 33.73105, 
    32.85971, 31.98156, 31.09665, 30.20505, 29.3068, 28.40199, 27.4907, 
    26.57302, 25.64905, 24.71892, 23.78273, 22.84064, 21.89278, 20.9393, 
    19.98038, 19.0162, 18.04693, 17.07278, 16.09396, 15.11067, 14.12316, 
    13.13165, 12.1364, 11.13764, 10.13566, 9.130703, 8.123061, 7.113011, 
    6.100842, 5.086846, 4.071321, 3.054569, 2.036894, 1.018601, 1.272222e-14, 
    -1.018601, -2.036894, -3.054569, -4.071321, -5.086846, -6.100842, 
    -7.113011, -8.123061, -9.130703, -10.13566, -11.13764, -12.1364, 
    -13.13165, -14.12316, -15.11067, -16.09396, -17.07278, -18.04693, 
    -19.0162, -19.98038, -20.9393, -21.89278, -22.84064, -23.78273, 
    -24.71892, -25.64905, -26.57302, -27.4907, -28.40199, -29.3068, 
    -30.20505, -31.09665, -31.98156, -32.85971, -33.73105, -34.59556, 
    -35.45321, -36.30396, -37.14782, -37.98478, -38.81484, -39.63801, 
    -40.45432, -41.26377, -42.06641, -42.86227, -43.65138, -44.4338,
  44.32701, 43.54469, 42.75576, 41.96017, 41.15789, 40.34887, 39.5331, 
    38.71054, 37.8812, 37.04504, 36.20208, 35.35233, 34.49578, 33.63246, 
    32.76241, 31.88566, 31.00225, 30.11224, 29.2157, 28.3127, 27.40331, 
    26.48764, 25.56579, 24.63787, 23.704, 22.76431, 21.81896, 20.8681, 
    19.91188, 18.95048, 17.9841, 17.01292, 16.03714, 15.05699, 14.07269, 
    13.08447, 12.09256, 11.09722, 10.09871, 9.097291, 8.09323, 7.086808, 
    6.078306, 5.068013, 4.05622, 3.043222, 2.029319, 1.014811, 1.272222e-14, 
    -1.014811, -2.029319, -3.043222, -4.05622, -5.068013, -6.078306, 
    -7.086808, -8.09323, -9.097291, -10.09871, -11.09722, -12.09256, 
    -13.08447, -14.07269, -15.05699, -16.03714, -17.01292, -17.9841, 
    -18.95048, -19.91188, -20.8681, -21.81896, -22.76431, -23.704, -24.63787, 
    -25.56579, -26.48764, -27.40331, -28.3127, -29.2157, -30.11224, 
    -31.00225, -31.88566, -32.76241, -33.63246, -34.49578, -35.35233, 
    -36.20208, -37.04504, -37.8812, -38.71054, -39.5331, -40.34887, 
    -41.15789, -41.96017, -42.75576, -43.54469, -44.32701,
  44.21122, 43.42903, 42.64032, 41.84503, 41.04314, 40.23461, 39.41943, 
    38.59755, 37.76899, 36.93372, 36.09175, 35.24308, 34.38773, 33.52573, 
    32.65709, 31.78186, 30.90008, 30.01182, 29.11712, 28.21608, 27.30877, 
    26.39529, 25.47573, 24.55021, 23.61885, 22.68178, 21.73915, 20.79111, 
    19.83782, 18.87945, 17.91618, 16.94822, 15.97575, 14.99899, 14.01815, 
    13.03348, 12.0452, 11.05355, 10.0588, 9.061195, 8.061007, 7.058504, 
    6.053965, 5.047671, 4.039908, 3.030967, 2.021138, 1.010717, 1.272222e-14, 
    -1.010717, -2.021138, -3.030967, -4.039908, -5.047671, -6.053965, 
    -7.058504, -8.061007, -9.061195, -10.0588, -11.05355, -12.0452, 
    -13.03348, -14.01815, -14.99899, -15.97575, -16.94822, -17.91618, 
    -18.87945, -19.83782, -20.79111, -21.73915, -22.68178, -23.61885, 
    -24.55021, -25.47573, -26.39529, -27.30877, -28.21608, -29.11712, 
    -30.01182, -30.90008, -31.78186, -32.65709, -33.52573, -34.38773, 
    -35.24308, -36.09175, -36.93372, -37.76899, -38.59755, -39.41943, 
    -40.23461, -41.04314, -41.84503, -42.64032, -43.42903, -44.21122,
  44.08652, 43.30448, 42.516, 41.72106, 40.91961, 40.11162, 39.29708, 
    38.47596, 37.64825, 36.81395, 35.97306, 35.12558, 34.27153, 33.41094, 
    32.54383, 31.67025, 30.79025, 29.90387, 29.01118, 28.11226, 27.20719, 
    26.29606, 25.37897, 24.45604, 23.52739, 22.59314, 21.65344, 20.70844, 
    19.7583, 18.80319, 17.84328, 16.87877, 15.90985, 14.93673, 13.95963, 
    12.97877, 11.99438, 11.0067, 10.01598, 9.02247, 8.026436, 7.02814, 
    6.027852, 5.025849, 4.022411, 3.017821, 2.012363, 1.006326, 1.272222e-14, 
    -1.006326, -2.012363, -3.017821, -4.022411, -5.025849, -6.027852, 
    -7.02814, -8.026436, -9.02247, -10.01598, -11.0067, -11.99438, -12.97877, 
    -13.95963, -14.93673, -15.90985, -16.87877, -17.84328, -18.80319, 
    -19.7583, -20.70844, -21.65344, -22.59314, -23.52739, -24.45604, 
    -25.37897, -26.29606, -27.20719, -28.11226, -29.01118, -29.90387, 
    -30.79025, -31.67025, -32.54383, -33.41094, -34.27153, -35.12558, 
    -35.97306, -36.81395, -37.64825, -38.47596, -39.29708, -40.11162, 
    -40.91961, -41.72106, -42.516, -43.30448, -44.08652,
  43.95298, 43.17111, 42.38291, 41.58834, 40.78738, 39.97999, 39.16616, 
    38.34586, 37.51908, 36.68583, 35.8461, 34.99992, 34.14728, 33.28822, 
    32.42276, 31.55096, 30.67286, 29.78851, 28.89797, 28.00133, 27.09867, 
    26.19007, 25.27564, 24.35549, 23.42973, 22.49851, 21.56195, 20.6202, 
    19.67343, 18.7218, 17.76548, 16.80466, 15.83954, 14.87031, 13.89719, 
    12.9204, 11.94017, 10.95672, 9.970306, 8.981172, 7.989569, 6.995759, 
    6.000007, 5.002581, 4.003754, 3.003803, 2.003006, 1.001644, 1.272222e-14, 
    -1.001644, -2.003006, -3.003803, -4.003754, -5.002581, -6.000007, 
    -6.995759, -7.989569, -8.981172, -9.970306, -10.95672, -11.94017, 
    -12.9204, -13.89719, -14.87031, -15.83954, -16.80466, -17.76548, 
    -18.7218, -19.67343, -20.6202, -21.56195, -22.49851, -23.42973, 
    -24.35549, -25.27564, -26.19007, -27.09867, -28.00133, -28.89797, 
    -29.78851, -30.67286, -31.55096, -32.42276, -33.28822, -34.14728, 
    -34.99992, -35.8461, -36.68583, -37.51908, -38.34586, -39.16616, 
    -39.97999, -40.78738, -41.58834, -42.38291, -43.17111, -43.95298,
  43.81068, 43.02901, 42.24112, 41.44698, 40.64656, 39.83982, 39.02676, 
    38.20735, 37.38158, 36.54947, 35.71101, 34.8662, 34.01508, 33.15767, 
    32.29399, 31.4241, 30.54803, 29.66586, 28.77763, 27.88343, 26.98333, 
    26.07744, 25.16584, 24.24865, 23.32599, 22.39799, 21.46477, 20.5265, 
    19.58331, 18.63538, 17.68288, 16.72599, 15.7649, 14.79981, 13.83093, 
    12.85847, 11.88264, 10.90369, 9.92185, 8.937356, 7.950458, 6.96141, 
    5.970469, 4.977899, 3.983964, 2.988935, 1.993082, 0.9966785, 
    1.272222e-14, -0.9966785, -1.993082, -2.988935, -3.983964, -4.977899, 
    -5.970469, -6.96141, -7.950458, -8.937356, -9.92185, -10.90369, 
    -11.88264, -12.85847, -13.83093, -14.79981, -15.7649, -16.72599, 
    -17.68288, -18.63538, -19.58331, -20.5265, -21.46477, -22.39799, 
    -23.32599, -24.24865, -25.16584, -26.07744, -26.98333, -27.88343, 
    -28.77763, -29.66586, -30.54803, -31.4241, -32.29399, -33.15767, 
    -34.01508, -34.8662, -35.71101, -36.54947, -37.38158, -38.20735, 
    -39.02676, -39.83982, -40.64656, -41.44698, -42.24112, -43.02901, 
    -43.81068,
  43.65969, 42.87827, 42.09073, 41.29707, 40.49723, 39.69121, 38.87898, 
    38.06054, 37.23587, 36.40498, 35.56787, 34.72456, 33.87507, 33.01942, 
    32.15764, 31.28979, 30.4159, 29.53604, 28.65027, 27.75867, 26.86131, 
    25.95829, 25.0497, 24.13567, 23.21629, 22.2917, 21.36204, 20.42744, 
    19.48806, 18.54405, 17.5956, 16.64287, 15.68605, 14.72534, 13.76093, 
    12.79304, 11.82189, 10.84769, 9.870676, 8.891085, 7.909157, 6.925138, 
    5.939281, 4.951838, 3.963069, 2.973237, 1.982603, 0.9914355, 
    1.272222e-14, -0.9914355, -1.982603, -2.973237, -3.963069, -4.951838, 
    -5.939281, -6.925138, -7.909157, -8.891085, -9.870676, -10.84769, 
    -11.82189, -12.79304, -13.76093, -14.72534, -15.68605, -16.64287, 
    -17.5956, -18.54405, -19.48806, -20.42744, -21.36204, -22.2917, 
    -23.21629, -24.13567, -25.0497, -25.95829, -26.86131, -27.75867, 
    -28.65027, -29.53604, -30.4159, -31.28979, -32.15764, -33.01942, 
    -33.87507, -34.72456, -35.56787, -36.40498, -37.23587, -38.06054, 
    -38.87898, -39.69121, -40.49723, -41.29707, -42.09073, -42.87827, 
    -43.65969,
  43.50012, 42.71897, 41.93184, 41.13869, 40.3395, 39.53426, 38.72294, 
    37.90554, 37.08205, 36.25248, 35.41682, 34.57511, 33.72735, 32.87358, 
    32.01384, 31.14815, 30.27658, 29.39919, 28.51603, 27.62718, 26.73272, 
    25.83275, 24.92736, 24.01665, 23.10075, 22.17978, 21.25386, 20.32315, 
    19.38778, 18.44792, 17.50373, 16.55539, 15.60307, 14.64697, 13.68729, 
    12.72422, 11.75798, 10.78878, 9.816853, 8.842422, 7.865723, 6.886996, 
    5.906484, 4.924435, 3.941099, 2.956731, 1.971586, 0.9859229, 
    1.272222e-14, -0.9859229, -1.971586, -2.956731, -3.941099, -4.924435, 
    -5.906484, -6.886996, -7.865723, -8.842422, -9.816853, -10.78878, 
    -11.75798, -12.72422, -13.68729, -14.64697, -15.60307, -16.55539, 
    -17.50373, -18.44792, -19.38778, -20.32315, -21.25386, -22.17978, 
    -23.10075, -24.01665, -24.92736, -25.83275, -26.73272, -27.62718, 
    -28.51603, -29.39919, -30.27658, -31.14815, -32.01384, -32.87358, 
    -33.72735, -34.57511, -35.41682, -36.25248, -37.08205, -37.90554, 
    -38.72294, -39.53426, -40.3395, -41.13869, -41.93184, -42.71897, -43.50012,
  43.33206, 42.55122, 41.76453, 40.97196, 40.17348, 39.36908, 38.55875, 
    37.74247, 36.92025, 36.09208, 35.25799, 34.41798, 33.57207, 32.7203, 
    31.86271, 30.99933, 30.13022, 29.25543, 28.37503, 27.4891, 26.59771, 
    25.70096, 24.79893, 23.89175, 22.97951, 22.06234, 21.14038, 20.21375, 
    19.28261, 18.34711, 17.4074, 16.46367, 15.51608, 14.56483, 13.61009, 
    12.65208, 11.691, 10.72705, 9.760451, 8.791431, 7.820215, 6.847034, 
    5.872125, 4.895727, 3.918083, 2.93944, 1.960045, 0.9801481, 1.272222e-14, 
    -0.9801481, -1.960045, -2.93944, -3.918083, -4.895727, -5.872125, 
    -6.847034, -7.820215, -8.791431, -9.760451, -10.72705, -11.691, 
    -12.65208, -13.61009, -14.56483, -15.51608, -16.46367, -17.4074, 
    -18.34711, -19.28261, -20.21375, -21.14038, -22.06234, -22.97951, 
    -23.89175, -24.79893, -25.70096, -26.59771, -27.4891, -28.37503, 
    -29.25543, -30.13022, -30.99933, -31.86271, -32.7203, -33.57207, 
    -34.41798, -35.25799, -36.09208, -36.92025, -37.74247, -38.55875, 
    -39.36908, -40.17348, -40.97196, -41.76453, -42.55122, -43.33206,
  43.1556, 42.37512, 41.58892, 40.79699, 39.99928, 39.1958, 38.38652, 
    37.57145, 36.75058, 35.92393, 35.09149, 34.25329, 33.40936, 32.55971, 
    31.7044, 30.84346, 29.97694, 29.10491, 28.22743, 27.34457, 26.45642, 
    25.56305, 24.66457, 23.76108, 22.85269, 21.93953, 21.02171, 20.09937, 
    19.17266, 18.24172, 17.30672, 16.36782, 15.42518, 14.479, 13.52945, 
    12.57673, 11.62103, 10.66257, 9.701547, 8.738181, 7.772693, 6.805305, 
    5.836247, 4.865752, 3.894052, 2.921387, 1.947996, 0.9741191, 
    1.272222e-14, -0.9741191, -1.947996, -2.921387, -3.894052, -4.865752, 
    -5.836247, -6.805305, -7.772693, -8.738181, -9.701547, -10.66257, 
    -11.62103, -12.57673, -13.52945, -14.479, -15.42518, -16.36782, 
    -17.30672, -18.24172, -19.17266, -20.09937, -21.02171, -21.93953, 
    -22.85269, -23.76108, -24.66457, -25.56305, -26.45642, -27.34457, 
    -28.22743, -29.10491, -29.97694, -30.84346, -31.7044, -32.55971, 
    -33.40936, -34.25329, -35.09149, -35.92393, -36.75058, -37.57145, 
    -38.38652, -39.1958, -39.99928, -40.79699, -41.58892, -42.37512, -43.1556,
  42.97084, 42.19077, 41.40512, 40.61388, 39.81702, 39.01452, 38.20639, 
    37.39261, 36.57319, 35.74813, 34.91746, 34.08119, 33.23934, 32.39194, 
    31.53904, 30.68068, 29.8169, 28.94778, 28.07337, 27.19374, 26.30898, 
    25.41917, 24.52441, 23.6248, 22.72045, 21.81147, 20.89799, 19.98014, 
    19.05806, 18.1319, 17.20181, 16.26795, 15.33048, 14.38959, 13.44545, 
    12.49824, 11.54817, 10.59543, 9.640213, 8.682739, 7.723217, 6.761864, 
    5.7989, 4.834549, 3.869038, 2.902596, 1.935454, 0.9678438, 1.272222e-14, 
    -0.9678438, -1.935454, -2.902596, -3.869038, -4.834549, -5.7989, 
    -6.761864, -7.723217, -8.682739, -9.640213, -10.59543, -11.54817, 
    -12.49824, -13.44545, -14.38959, -15.33048, -16.26795, -17.20181, 
    -18.1319, -19.05806, -19.98014, -20.89799, -21.81147, -22.72045, 
    -23.6248, -24.52441, -25.41917, -26.30898, -27.19374, -28.07337, 
    -28.94778, -29.8169, -30.68068, -31.53904, -32.39194, -33.23934, 
    -34.08119, -34.91746, -35.74813, -36.57319, -37.39261, -38.20639, 
    -39.01452, -39.81702, -40.61388, -41.40512, -42.19077, -42.97084,
  42.77788, 41.99827, 41.21324, 40.42275, 39.6268, 38.82537, 38.01846, 
    37.20607, 36.38819, 35.56485, 34.73605, 33.90181, 33.06216, 32.21714, 
    31.36679, 30.51114, 29.65025, 28.78417, 27.91298, 27.03675, 26.15555, 
    25.26947, 24.3786, 23.48304, 22.5829, 21.6783, 20.76936, 19.85619, 
    18.93895, 18.01776, 17.09279, 16.16418, 15.2321, 14.29671, 13.3582, 
    12.41673, 11.47251, 10.52571, 9.576528, 8.625175, 7.671851, 6.716765, 
    5.760129, 4.802159, 3.843073, 2.883091, 1.922435, 0.9613302, 
    1.272222e-14, -0.9613302, -1.922435, -2.883091, -3.843073, -4.802159, 
    -5.760129, -6.716765, -7.671851, -8.625175, -9.576528, -10.52571, 
    -11.47251, -12.41673, -13.3582, -14.29671, -15.2321, -16.16418, 
    -17.09279, -18.01776, -18.93895, -19.85619, -20.76936, -21.6783, 
    -22.5829, -23.48304, -24.3786, -25.26947, -26.15555, -27.03675, 
    -27.91298, -28.78417, -29.65025, -30.51114, -31.36679, -32.21714, 
    -33.06216, -33.90181, -34.73605, -35.56485, -36.38819, -37.20607, 
    -38.01846, -38.82537, -39.6268, -40.42275, -41.21324, -41.99827, -42.77788,
  42.57683, 41.79774, 41.01338, 40.22372, 39.42876, 38.62848, 37.82288, 
    37.01196, 36.19573, 35.3742, 34.54738, 33.7153, 32.87798, 32.03546, 
    31.18778, 30.33498, 29.47712, 28.61425, 27.74643, 26.87375, 25.99627, 
    25.11408, 24.22728, 23.33596, 22.44022, 21.54018, 20.63595, 19.72766, 
    18.81544, 17.89944, 16.97978, 16.05663, 15.13014, 14.20047, 13.2678, 
    12.33229, 11.39412, 10.45349, 9.510569, 8.565559, 7.618658, 6.670065, 
    5.719984, 4.768622, 3.816189, 2.862896, 1.908957, 0.9545865, 
    1.272222e-14, -0.9545865, -1.908957, -2.862896, -3.816189, -4.768622, 
    -5.719984, -6.670065, -7.618658, -8.565559, -9.510569, -10.45349, 
    -11.39412, -12.33229, -13.2678, -14.20047, -15.13014, -16.05663, 
    -16.97978, -17.89944, -18.81544, -19.72766, -20.63595, -21.54018, 
    -22.44022, -23.33596, -24.22728, -25.11408, -25.99627, -26.87375, 
    -27.74643, -28.61425, -29.47712, -30.33498, -31.18778, -32.03546, 
    -32.87798, -33.7153, -34.54738, -35.3742, -36.19573, -37.01196, 
    -37.82288, -38.62848, -39.42876, -40.22372, -41.01338, -41.79774, 
    -42.57683,
  42.36781, 41.5893, 40.80568, 40.01692, 39.22302, 38.42397, 37.61977, 
    36.81043, 35.99594, 35.17633, 34.35161, 33.5218, 32.68693, 31.84704, 
    31.00217, 30.15236, 29.29767, 28.43815, 27.57387, 26.70489, 25.8313, 
    24.95318, 24.07061, 23.18369, 22.29253, 21.39723, 20.49791, 19.59469, 
    18.68769, 17.77705, 16.86292, 15.94542, 15.02473, 14.10098, 13.17436, 
    12.24501, 11.31312, 10.37886, 9.442413, 8.503963, 7.563702, 6.621819, 
    5.678512, 4.733978, 3.788419, 2.842036, 1.895035, 0.947621, 1.272222e-14, 
    -0.947621, -1.895035, -2.842036, -3.788419, -4.733978, -5.678512, 
    -6.621819, -7.563702, -8.503963, -9.442413, -10.37886, -11.31312, 
    -12.24501, -13.17436, -14.10098, -15.02473, -15.94542, -16.86292, 
    -17.77705, -18.68769, -19.59469, -20.49791, -21.39723, -22.29253, 
    -23.18369, -24.07061, -24.95318, -25.8313, -26.70489, -27.57387, 
    -28.43815, -29.29767, -30.15236, -31.00217, -31.84704, -32.68693, 
    -33.5218, -34.35161, -35.17633, -35.99594, -36.81043, -37.61977, 
    -38.42397, -39.22302, -40.01692, -40.80568, -41.5893, -42.36781,
  42.15091, 41.37305, 40.59023, 39.80246, 39.00971, 38.21198, 37.40928, 
    36.6016, 35.78897, 34.97139, 34.14888, 33.32146, 32.48917, 31.65205, 
    30.81012, 29.96344, 29.11207, 28.25605, 27.39545, 26.53034, 25.6608, 
    24.7869, 23.90874, 23.0264, 22.13999, 21.24961, 20.35538, 19.45741, 
    18.55582, 17.65075, 16.74232, 15.83068, 14.91598, 13.99836, 13.07798, 
    12.155, 11.22959, 10.30191, 9.372141, 8.44046, 7.507047, 6.572086, 
    5.635764, 4.69827, 3.759796, 2.820537, 1.880687, 0.9404421, 1.272222e-14, 
    -0.9404421, -1.880687, -2.820537, -3.759796, -4.69827, -5.635764, 
    -6.572086, -7.507047, -8.44046, -9.372141, -10.30191, -11.22959, -12.155, 
    -13.07798, -13.99836, -14.91598, -15.83068, -16.74232, -17.65075, 
    -18.55582, -19.45741, -20.35538, -21.24961, -22.13999, -23.0264, 
    -23.90874, -24.7869, -25.6608, -26.53034, -27.39545, -28.25605, 
    -29.11207, -29.96344, -30.81012, -31.65205, -32.48917, -33.32146, 
    -34.14888, -34.97139, -35.78897, -36.6016, -37.40928, -38.21198, 
    -39.00971, -39.80246, -40.59023, -41.37305, -42.15091,
  41.92625, 41.14911, 40.36718, 39.58046, 38.78895, 37.99264, 37.19153, 
    36.38563, 35.57495, 34.75951, 33.93933, 33.11443, 32.28485, 31.45062, 
    30.61178, 29.76838, 28.92046, 28.06809, 27.21133, 26.35024, 25.48491, 
    24.6154, 23.74181, 22.86423, 21.98275, 21.09747, 20.20851, 19.31597, 
    18.41997, 17.52065, 16.61812, 15.71253, 14.804, 13.8927, 12.97877, 
    12.06235, 11.14361, 10.22272, 9.299832, 8.375121, 7.448759, 6.520922, 
    5.591787, 4.661538, 3.730354, 2.798423, 1.865928, 0.9330581, 
    1.272222e-14, -0.9330581, -1.865928, -2.798423, -3.730354, -4.661538, 
    -5.591787, -6.520922, -7.448759, -8.375121, -9.299832, -10.22272, 
    -11.14361, -12.06235, -12.97877, -13.8927, -14.804, -15.71253, -16.61812, 
    -17.52065, -18.41997, -19.31597, -20.20851, -21.09747, -21.98275, 
    -22.86423, -23.74181, -24.6154, -25.48491, -26.35024, -27.21133, 
    -28.06809, -28.92046, -29.76838, -30.61178, -31.45062, -32.28485, 
    -33.11443, -33.93933, -34.75951, -35.57495, -36.38563, -37.19153, 
    -37.99264, -38.78895, -39.58046, -40.36718, -41.14911, -41.92625,
  41.69396, 40.9176, 40.13664, 39.35107, 38.56088, 37.76608, 36.96666, 
    36.16264, 35.35404, 34.54086, 33.72313, 32.90088, 32.07413, 31.24292, 
    30.4073, 29.56732, 28.72301, 27.87444, 27.02167, 26.16477, 25.3038, 
    24.43885, 23.57, 22.69734, 21.82095, 20.94095, 20.05743, 19.1705, 
    18.28028, 17.38689, 16.49044, 15.59108, 14.68893, 13.78413, 12.87683, 
    11.96717, 11.0553, 10.14138, 9.225567, 8.308019, 7.388902, 6.468383, 
    5.546633, 4.623823, 3.700126, 2.775718, 1.850776, 0.9254774, 
    1.272222e-14, -0.9254774, -1.850776, -2.775718, -3.700126, -4.623823, 
    -5.546633, -6.468383, -7.388902, -8.308019, -9.225567, -10.14138, 
    -11.0553, -11.96717, -12.87683, -13.78413, -14.68893, -15.59108, 
    -16.49044, -17.38689, -18.28028, -19.1705, -20.05743, -20.94095, 
    -21.82095, -22.69734, -23.57, -24.43885, -25.3038, -26.16477, -27.02167, 
    -27.87444, -28.72301, -29.56732, -30.4073, -31.24292, -32.07413, 
    -32.90088, -33.72313, -34.54086, -35.35404, -36.16264, -36.96666, 
    -37.76608, -38.56088, -39.35107, -40.13664, -40.9176, -41.69396,
  41.45414, 40.67865, 39.89874, 39.1144, 38.32563, 37.53244, 36.73482, 
    35.9328, 35.12637, 34.31557, 33.50042, 32.68093, 31.85715, 31.02912, 
    30.19686, 29.36043, 28.51988, 27.67526, 26.82663, 25.97407, 25.11763, 
    24.2574, 23.39345, 22.52588, 21.65476, 20.7802, 19.9023, 19.02115, 
    18.13688, 17.2496, 16.35942, 15.46647, 14.57087, 13.67276, 12.77227, 
    11.86955, 10.96474, 10.05798, 9.149424, 8.239225, 7.327541, 6.414529, 
    5.50035, 4.585167, 3.669145, 2.752449, 1.835248, 0.9177083, 1.272222e-14, 
    -0.9177083, -1.835248, -2.752449, -3.669145, -4.585167, -5.50035, 
    -6.414529, -7.327541, -8.239225, -9.149424, -10.05798, -10.96474, 
    -11.86955, -12.77227, -13.67276, -14.57087, -15.46647, -16.35942, 
    -17.2496, -18.13688, -19.02115, -19.9023, -20.7802, -21.65476, -22.52588, 
    -23.39345, -24.2574, -25.11763, -25.97407, -26.82663, -27.67526, 
    -28.51988, -29.36043, -30.19686, -31.02912, -31.85715, -32.68093, 
    -33.50042, -34.31557, -35.12637, -35.9328, -36.73482, -37.53244, 
    -38.32563, -39.1144, -39.89874, -40.67865, -41.45414,
  41.20691, 40.43238, 39.6536, 38.87059, 38.08334, 37.29186, 36.49615, 
    35.69623, 34.89211, 34.08381, 33.27135, 32.45477, 31.63409, 30.80936, 
    29.9806, 29.14787, 28.31122, 27.47071, 26.62638, 25.77831, 24.92656, 
    24.0712, 23.21232, 22.35, 21.48432, 20.61537, 19.74325, 18.86807, 
    17.98992, 17.10892, 16.22518, 15.33881, 14.44994, 13.5587, 12.66521, 
    11.7696, 10.87202, 9.972599, 9.071482, 8.168813, 7.26474, 6.359414, 
    5.452987, 4.545611, 3.637443, 2.72864, 1.819359, 0.9097592, 1.272222e-14, 
    -0.9097592, -1.819359, -2.72864, -3.637443, -4.545611, -5.452987, 
    -6.359414, -7.26474, -8.168813, -9.071482, -9.972599, -10.87202, 
    -11.7696, -12.66521, -13.5587, -14.44994, -15.33881, -16.22518, 
    -17.10892, -17.98992, -18.86807, -19.74325, -20.61537, -21.48432, -22.35, 
    -23.21232, -24.0712, -24.92656, -25.77831, -26.62638, -27.47071, 
    -28.31122, -29.14787, -29.9806, -30.80936, -31.63409, -32.45477, 
    -33.27135, -34.08381, -34.89211, -35.69623, -36.49615, -37.29186, 
    -38.08334, -38.87059, -39.6536, -40.43238, -41.20691,
  40.9524, 40.1789, 39.40136, 38.61978, 37.83415, 37.04449, 36.2508, 
    35.45309, 34.6514, 33.84572, 33.03609, 32.22254, 31.4051, 30.5838, 
    29.75869, 28.92981, 28.09721, 27.26094, 26.42107, 25.57764, 24.73074, 
    23.88042, 23.02677, 22.16986, 21.30978, 20.44661, 19.58045, 18.71139, 
    17.83953, 16.96498, 16.08784, 15.20823, 14.32627, 13.44206, 12.55573, 
    11.66742, 10.77724, 9.885328, 8.99182, 8.096853, 7.200565, 6.303097, 
    5.404592, 4.505196, 3.605054, 2.704315, 1.803126, 0.9016382, 
    1.272222e-14, -0.9016382, -1.803126, -2.704315, -3.605054, -4.505196, 
    -5.404592, -6.303097, -7.200565, -8.096853, -8.99182, -9.885328, 
    -10.77724, -11.66742, -12.55573, -13.44206, -14.32627, -15.20823, 
    -16.08784, -16.96498, -17.83953, -18.71139, -19.58045, -20.44661, 
    -21.30978, -22.16986, -23.02677, -23.88042, -24.73074, -25.57764, 
    -26.42107, -27.26094, -28.09721, -28.92981, -29.75869, -30.5838, 
    -31.4051, -32.22254, -33.03609, -33.84572, -34.6514, -35.45309, -36.2508, 
    -37.04449, -37.83415, -38.61978, -39.40136, -40.1789, -40.9524,
  40.69072, 39.91835, 39.14214, 38.36209, 37.57819, 36.79046, 35.9989, 
    35.20354, 34.40438, 33.60146, 32.79479, 31.98441, 31.17034, 30.35262, 
    29.5313, 28.70641, 27.87801, 27.04614, 26.21087, 25.37224, 24.53034, 
    23.68522, 22.83695, 21.98561, 21.13129, 20.27407, 19.41402, 18.55125, 
    17.68585, 16.81791, 15.94755, 15.07486, 14.19996, 13.32295, 12.44396, 
    11.5631, 10.68048, 9.79625, 8.910519, 8.023417, 7.135077, 6.245632, 
    5.355214, 4.463961, 3.57201, 2.679499, 1.786567, 0.8933536, 1.272222e-14, 
    -0.8933536, -1.786567, -2.679499, -3.57201, -4.463961, -5.355214, 
    -6.245632, -7.135077, -8.023417, -8.910519, -9.79625, -10.68048, 
    -11.5631, -12.44396, -13.32295, -14.19996, -15.07486, -15.94755, 
    -16.81791, -17.68585, -18.55125, -19.41402, -20.27407, -21.13129, 
    -21.98561, -22.83695, -23.68522, -24.53034, -25.37224, -26.21087, 
    -27.04614, -27.87801, -28.70641, -29.5313, -30.35262, -31.17034, 
    -31.98441, -32.79479, -33.60146, -34.40438, -35.20354, -35.9989, 
    -36.79046, -37.57819, -38.36209, -39.14214, -39.91835, -40.69072,
  40.42199, 39.65086, 38.87608, 38.09766, 37.3156, 36.52991, 35.74061, 
    34.94771, 34.15122, 33.35118, 32.5476, 31.74052, 30.92996, 30.11596, 
    29.29857, 28.47782, 27.65377, 26.82645, 25.99593, 25.16227, 24.32551, 
    23.48574, 22.64302, 21.79742, 20.94901, 20.09789, 19.24412, 18.38779, 
    17.52901, 16.66785, 15.80442, 14.93881, 14.07113, 13.20149, 12.32998, 
    11.45673, 10.58185, 9.705451, 8.827652, 7.948575, 7.068341, 6.187074, 
    5.304901, 4.421948, 3.538343, 2.654216, 1.769696, 0.8849133, 
    1.272222e-14, -0.8849133, -1.769696, -2.654216, -3.538343, -4.421948, 
    -5.304901, -6.187074, -7.068341, -7.948575, -8.827652, -9.705451, 
    -10.58185, -11.45673, -12.32998, -13.20149, -14.07113, -14.93881, 
    -15.80442, -16.66785, -17.52901, -18.38779, -19.24412, -20.09789, 
    -20.94901, -21.79742, -22.64302, -23.48574, -24.32551, -25.16227, 
    -25.99593, -26.82645, -27.65377, -28.47782, -29.29857, -30.11596, 
    -30.92996, -31.74052, -32.5476, -33.35118, -34.15122, -34.94771, 
    -35.74061, -36.52991, -37.3156, -38.09766, -38.87608, -39.65086, -40.42199,
  40.14635, 39.37654, 38.6033, 37.82662, 37.04652, 36.26299, 35.47607, 
    34.68575, 33.89207, 33.09504, 32.29469, 31.49104, 30.68413, 29.874, 
    29.06068, 28.24422, 27.42466, 26.60204, 25.77643, 24.94787, 24.11643, 
    23.28216, 22.44514, 21.60542, 20.76309, 19.91821, 19.07088, 18.22116, 
    17.36914, 16.51492, 15.65857, 14.8002, 13.9399, 13.07777, 12.21391, 
    11.34843, 10.48143, 9.613013, 8.743299, 7.872395, 7.000417, 6.12748, 
    5.253699, 4.379195, 3.504085, 2.628489, 1.752529, 0.8763254, 
    1.272222e-14, -0.8763254, -1.752529, -2.628489, -3.504085, -4.379195, 
    -5.253699, -6.12748, -7.000417, -7.872395, -8.743299, -9.613013, 
    -10.48143, -11.34843, -12.21391, -13.07777, -13.9399, -14.8002, 
    -15.65857, -16.51492, -17.36914, -18.22116, -19.07088, -19.91821, 
    -20.76309, -21.60542, -22.44514, -23.28216, -24.11643, -24.94787, 
    -25.77643, -26.60204, -27.42466, -28.24422, -29.06068, -29.874, 
    -30.68413, -31.49104, -32.29469, -33.09504, -33.89207, -34.68575, 
    -35.47607, -36.26299, -37.04652, -37.82662, -38.6033, -39.37654, -40.14635,
  39.8639, 39.09554, 38.32394, 37.54912, 36.77109, 35.98985, 35.20542, 
    34.41782, 33.62707, 32.83318, 32.03619, 31.23613, 30.43301, 29.62689, 
    28.81779, 28.00576, 27.19084, 26.37307, 25.55252, 24.72922, 23.90323, 
    23.07462, 22.24345, 21.40977, 20.57367, 19.7352, 18.89445, 18.05148, 
    17.20639, 16.35925, 15.51014, 14.65916, 13.80638, 12.95192, 12.09585, 
    11.23828, 10.3793, 9.519018, 8.657532, 7.794946, 6.931367, 6.066901, 
    5.201655, 4.335741, 3.469266, 2.602343, 1.735083, 0.8675976, 
    1.272222e-14, -0.8675976, -1.735083, -2.602343, -3.469266, -4.335741, 
    -5.201655, -6.066901, -6.931367, -7.794946, -8.657532, -9.519018, 
    -10.3793, -11.23828, -12.09585, -12.95192, -13.80638, -14.65916, 
    -15.51014, -16.35925, -17.20639, -18.05148, -18.89445, -19.7352, 
    -20.57367, -21.40977, -22.24345, -23.07462, -23.90323, -24.72922, 
    -25.55252, -26.37307, -27.19084, -28.00576, -28.81779, -29.62689, 
    -30.43301, -31.23613, -32.03619, -32.83318, -33.62707, -34.41782, 
    -35.20542, -35.98985, -36.77109, -37.54912, -38.32394, -39.09554, -39.8639,
  39.57478, 38.80796, 38.03813, 37.26529, 36.48944, 35.71062, 34.92882, 
    34.14407, 33.35638, 32.56578, 31.77229, 30.97594, 30.17676, 29.37479, 
    28.57006, 27.76261, 26.95247, 26.13971, 25.32435, 24.50646, 23.68609, 
    22.86328, 22.03811, 21.21062, 20.38089, 19.54898, 18.71496, 17.8789, 
    17.04088, 16.20097, 15.35924, 14.51579, 13.67069, 12.82403, 11.97589, 
    11.12637, 10.27556, 9.423547, 8.570426, 7.716295, 6.86125, 6.00539, 
    5.148814, 4.291623, 3.433917, 2.575799, 1.717372, 0.8587376, 
    1.272222e-14, -0.8587376, -1.717372, -2.575799, -3.433917, -4.291623, 
    -5.148814, -6.00539, -6.86125, -7.716295, -8.570426, -9.423547, 
    -10.27556, -11.12637, -11.97589, -12.82403, -13.67069, -14.51579, 
    -15.35924, -16.20097, -17.04088, -17.8789, -18.71496, -19.54898, 
    -20.38089, -21.21062, -22.03811, -22.86328, -23.68609, -24.50646, 
    -25.32435, -26.13971, -26.95247, -27.76261, -28.57006, -29.37479, 
    -30.17676, -30.97594, -31.77229, -32.56578, -33.35638, -34.14407, 
    -34.92882, -35.71062, -36.48944, -37.26529, -38.03813, -38.80796, 
    -39.57478,
  39.27911, 38.51395, 37.746, 36.97525, 36.20173, 35.42545, 34.64641, 
    33.86464, 33.08015, 32.29297, 31.50312, 30.71063, 29.91554, 29.11786, 
    28.31764, 27.51491, 26.70972, 25.9021, 25.0921, 24.27976, 23.46515, 
    22.6483, 21.82927, 21.00812, 20.18491, 19.35971, 18.53256, 17.70355, 
    16.87274, 16.0402, 15.20599, 14.37021, 13.53292, 12.6942, 11.85414, 
    11.0128, 10.17029, 9.326677, 8.482054, 7.636507, 6.790126, 5.943, 
    5.095221, 4.246879, 3.398068, 2.548881, 1.699411, 0.8497528, 
    1.272222e-14, -0.8497528, -1.699411, -2.548881, -3.398068, -4.246879, 
    -5.095221, -5.943, -6.790126, -7.636507, -8.482054, -9.326677, -10.17029, 
    -11.0128, -11.85414, -12.6942, -13.53292, -14.37021, -15.20599, -16.0402, 
    -16.87274, -17.70355, -18.53256, -19.35971, -20.18491, -21.00812, 
    -21.82927, -22.6483, -23.46515, -24.27976, -25.0921, -25.9021, -26.70972, 
    -27.51491, -28.31764, -29.11786, -29.91554, -30.71063, -31.50312, 
    -32.29297, -33.08015, -33.86464, -34.64641, -35.42545, -36.20173, 
    -36.97525, -37.746, -38.51395, -39.27911,
  38.977, 38.21363, 37.44768, 36.67916, 35.90809, 35.13448, 34.35833, 
    33.57967, 32.79853, 32.01491, 31.22885, 30.44036, 29.64949, 28.85626, 
    28.0607, 27.26284, 26.46273, 25.6604, 24.85591, 24.04927, 23.24056, 
    22.42981, 21.61708, 20.80241, 19.98587, 19.16751, 18.34738, 17.52556, 
    16.7021, 15.87706, 15.05052, 14.22254, 13.39319, 12.56255, 11.73068, 
    10.89766, 10.06357, 9.228487, 8.392486, 7.555646, 6.718051, 5.87978, 
    5.040917, 4.201545, 3.361748, 2.52161, 1.681216, 0.8406506, 1.272222e-14, 
    -0.8406506, -1.681216, -2.52161, -3.361748, -4.201545, -5.040917, 
    -5.87978, -6.718051, -7.555646, -8.392486, -9.228487, -10.06357, 
    -10.89766, -11.73068, -12.56255, -13.39319, -14.22254, -15.05052, 
    -15.87706, -16.7021, -17.52556, -18.34738, -19.16751, -19.98587, 
    -20.80241, -21.61708, -22.42981, -23.24056, -24.04927, -24.85591, 
    -25.6604, -26.46273, -27.26284, -28.0607, -28.85626, -29.64949, 
    -30.44036, -31.22885, -32.01491, -32.79853, -33.57967, -34.35833, 
    -35.13448, -35.90809, -36.67916, -37.44768, -38.21363, -38.977,
  38.66859, 37.90713, 37.14331, 36.37715, 35.60866, 34.83784, 34.06473, 
    33.28933, 32.51167, 31.73176, 30.94962, 30.16529, 29.37879, 28.59014, 
    27.79938, 27.00655, 26.21167, 25.41478, 24.61593, 23.81515, 23.01249, 
    22.20798, 21.40168, 20.59364, 19.7839, 18.97252, 18.15956, 17.34505, 
    16.52908, 15.71168, 14.89293, 14.07288, 13.2516, 12.42916, 11.60561, 
    10.78103, 9.955491, 9.129053, 8.30179, 7.473776, 6.645081, 5.815781, 
    4.985948, 4.155657, 3.324986, 2.494007, 1.662799, 0.8314381, 
    1.272222e-14, -0.8314381, -1.662799, -2.494007, -3.324986, -4.155657, 
    -4.985948, -5.815781, -6.645081, -7.473776, -8.30179, -9.129053, 
    -9.955491, -10.78103, -11.60561, -12.42916, -13.2516, -14.07288, 
    -14.89293, -15.71168, -16.52908, -17.34505, -18.15956, -18.97252, 
    -19.7839, -20.59364, -21.40168, -22.20798, -23.01249, -23.81515, 
    -24.61593, -25.41478, -26.21167, -27.00655, -27.79938, -28.59014, 
    -29.37879, -30.16529, -30.94962, -31.73176, -32.51167, -33.28933, 
    -34.06473, -34.83784, -35.60866, -36.37715, -37.14331, -37.90713, 
    -38.66859,
  38.354, 37.59457, 36.83301, 36.06934, 35.30357, 34.5357, 33.76576, 
    32.99376, 32.21972, 31.44366, 30.6656, 29.88556, 29.10357, 28.31966, 
    27.53386, 26.74619, 25.95669, 25.16539, 24.37232, 23.57754, 22.78106, 
    21.98295, 21.18322, 20.38194, 19.57915, 18.77489, 17.96921, 17.16216, 
    16.3538, 15.54417, 14.73334, 13.92135, 13.10826, 12.29414, 11.47903, 
    10.66301, 9.846126, 9.028447, 8.210036, 7.390956, 6.571271, 5.751048, 
    4.930352, 4.10925, 3.287808, 2.466094, 1.644176, 0.8221223, 1.272222e-14, 
    -0.8221223, -1.644176, -2.466094, -3.287808, -4.10925, -4.930352, 
    -5.751048, -6.571271, -7.390956, -8.210036, -9.028447, -9.846126, 
    -10.66301, -11.47903, -12.29414, -13.10826, -13.92135, -14.73334, 
    -15.54417, -16.3538, -17.16216, -17.96921, -18.77489, -19.57915, 
    -20.38194, -21.18322, -21.98295, -22.78106, -23.57754, -24.37232, 
    -25.16539, -25.95669, -26.74619, -27.53386, -28.31966, -29.10357, 
    -29.88556, -30.6656, -31.44366, -32.21972, -32.99376, -33.76576, 
    -34.5357, -35.30357, -36.06934, -36.83301, -37.59457, -38.354,
  38.03334, 37.27608, 36.51693, 35.75588, 34.99296, 34.22818, 33.46156, 
    32.6931, 31.92283, 31.15076, 30.37692, 29.60133, 28.82401, 28.04498, 
    27.26427, 26.48191, 25.69794, 24.91236, 24.12524, 23.33659, 22.54645, 
    21.75485, 20.96184, 20.16746, 19.37174, 18.57473, 17.77647, 16.97701, 
    16.17639, 15.37465, 14.57185, 13.76804, 12.96326, 12.15757, 11.35102, 
    10.54366, 9.735553, 8.926742, 8.117288, 7.307246, 6.496675, 5.68563, 
    4.874171, 4.062356, 3.250242, 2.437891, 1.62536, 0.8127099, 1.272222e-14, 
    -0.8127099, -1.62536, -2.437891, -3.250242, -4.062356, -4.874171, 
    -5.68563, -6.496675, -7.307246, -8.117288, -8.926742, -9.735553, 
    -10.54366, -11.35102, -12.15757, -12.96326, -13.76804, -14.57185, 
    -15.37465, -16.17639, -16.97701, -17.77647, -18.57473, -19.37174, 
    -20.16746, -20.96184, -21.75485, -22.54645, -23.33659, -24.12524, 
    -24.91236, -25.69794, -26.48191, -27.26427, -28.04498, -28.82401, 
    -29.60133, -30.37692, -31.15076, -31.92283, -32.6931, -33.46156, 
    -34.22818, -34.99296, -35.75588, -36.51693, -37.27608, -38.03334,
  37.70675, 36.95179, 36.19517, 35.4369, 34.67698, 33.91543, 33.15226, 
    32.3875, 31.62114, 30.85322, 30.08375, 29.31275, 28.54023, 27.76624, 
    26.99077, 26.21387, 25.43556, 24.65587, 23.87482, 23.09244, 22.30877, 
    21.52384, 20.73768, 19.95033, 19.16182, 18.37219, 17.58147, 16.78971, 
    15.99695, 15.20323, 14.40859, 13.61306, 12.81671, 12.01956, 11.22167, 
    10.42309, 9.623848, 8.824006, 8.023608, 7.222704, 6.421341, 5.619571, 
    4.817443, 4.015007, 3.212315, 2.409416, 1.606363, 0.8032075, 
    1.272222e-14, -0.8032075, -1.606363, -2.409416, -3.212315, -4.015007, 
    -4.817443, -5.619571, -6.421341, -7.222704, -8.023608, -8.824006, 
    -9.623848, -10.42309, -11.22167, -12.01956, -12.81671, -13.61306, 
    -14.40859, -15.20323, -15.99695, -16.78971, -17.58147, -18.37219, 
    -19.16182, -19.95033, -20.73768, -21.52384, -22.30877, -23.09244, 
    -23.87482, -24.65587, -25.43556, -26.21387, -26.99077, -27.76624, 
    -28.54023, -29.31275, -30.08375, -30.85322, -31.62114, -32.3875, 
    -33.15226, -33.91543, -34.67698, -35.4369, -36.19517, -36.95179, -37.70675,
  37.37434, 36.62183, 35.86789, 35.11252, 34.35575, 33.59758, 32.83802, 
    32.0771, 31.31481, 30.55118, 29.78622, 29.01996, 28.25241, 27.48358, 
    26.71351, 25.94222, 25.16972, 24.39604, 23.6212, 22.84524, 22.06818, 
    21.29005, 20.51087, 19.73068, 18.9495, 18.16737, 17.38433, 16.6004, 
    15.81561, 15.03002, 14.24364, 13.45652, 12.66869, 11.88019, 11.09107, 
    10.30135, 9.511086, 8.720308, 7.929061, 7.137385, 6.345323, 5.552916, 
    4.760206, 3.967237, 3.17405, 2.38069, 1.587199, 0.7936214, 1.272222e-14, 
    -0.7936214, -1.587199, -2.38069, -3.17405, -3.967237, -4.760206, 
    -5.552916, -6.345323, -7.137385, -7.929061, -8.720308, -9.511086, 
    -10.30135, -11.09107, -11.88019, -12.66869, -13.45652, -14.24364, 
    -15.03002, -15.81561, -16.6004, -17.38433, -18.16737, -18.9495, 
    -19.73068, -20.51087, -21.29005, -22.06818, -22.84524, -23.6212, 
    -24.39604, -25.16972, -25.94222, -26.71351, -27.48358, -28.25241, 
    -29.01996, -29.78622, -30.55118, -31.31481, -32.0771, -32.83802, 
    -33.59758, -34.35575, -35.11252, -35.86789, -36.62183, -37.37434,
  37.03624, 36.28631, 35.53519, 34.78289, 34.02942, 33.27477, 32.51897, 
    31.76203, 31.00396, 30.24478, 29.48449, 28.72311, 27.96067, 27.19717, 
    26.43264, 25.66709, 24.90054, 24.13302, 23.36455, 22.59513, 21.82482, 
    21.05361, 20.28154, 19.50863, 18.73492, 17.96042, 17.18516, 16.40917, 
    15.63248, 14.85512, 14.07711, 13.2985, 12.5193, 11.73955, 10.95929, 
    10.17854, 9.397336, 8.615713, 7.833705, 7.051345, 6.268667, 5.485706, 
    4.702497, 3.919074, 3.135473, 2.35173, 1.56788, 0.7839577, 1.272222e-14, 
    -0.7839577, -1.56788, -2.35173, -3.135473, -3.919074, -4.702497, 
    -5.485706, -6.268667, -7.051345, -7.833705, -8.615713, -9.397336, 
    -10.17854, -10.95929, -11.73955, -12.5193, -13.2985, -14.07711, 
    -14.85512, -15.63248, -16.40917, -17.18516, -17.96042, -18.73492, 
    -19.50863, -20.28154, -21.05361, -21.82482, -22.59513, -23.36455, 
    -24.13302, -24.90054, -25.66709, -26.43264, -27.19717, -27.96067, 
    -28.72311, -29.48449, -30.24478, -31.00396, -31.76203, -32.51897, 
    -33.27477, -34.02942, -34.78289, -35.53519, -36.28631, -37.03624,
  36.69255, 35.94537, 35.19722, 34.44813, 33.6981, 32.94714, 32.19525, 
    31.44245, 30.68875, 29.93416, 29.17869, 28.42235, 27.66517, 26.90714, 
    26.14829, 25.38863, 24.62818, 23.86696, 23.10497, 22.34225, 21.5788, 
    20.81466, 20.04982, 19.28433, 18.51819, 17.75143, 16.98408, 16.21614, 
    15.44765, 14.67863, 13.90911, 13.1391, 12.36863, 11.59772, 10.82641, 
    10.05472, 9.282667, 8.510284, 7.737598, 6.964634, 6.19142, 5.417983, 
    4.64435, 3.870549, 3.096608, 2.322554, 1.548416, 0.7742223, 1.272222e-14, 
    -0.7742223, -1.548416, -2.322554, -3.096608, -3.870549, -4.64435, 
    -5.417983, -6.19142, -6.964634, -7.737598, -8.510284, -9.282667, 
    -10.05472, -10.82641, -11.59772, -12.36863, -13.1391, -13.90911, 
    -14.67863, -15.44765, -16.21614, -16.98408, -17.75143, -18.51819, 
    -19.28433, -20.04982, -20.81466, -21.5788, -22.34225, -23.10497, 
    -23.86696, -24.62818, -25.38863, -26.14829, -26.90714, -27.66517, 
    -28.42235, -29.17869, -29.93416, -30.68875, -31.44245, -32.19525, 
    -32.94714, -33.6981, -34.44813, -35.19722, -35.94537, -36.69255,
  36.34341, 35.59911, 34.8541, 34.10837, 33.36194, 32.61481, 31.86699, 
    31.11849, 30.36931, 29.61947, 28.86897, 28.11782, 27.36604, 26.61363, 
    25.86061, 25.10699, 24.35277, 23.59798, 22.84263, 22.08672, 21.33028, 
    20.57332, 19.81585, 19.05788, 18.29944, 17.54054, 16.7812, 16.02143, 
    15.26124, 14.50067, 13.73972, 12.97841, 12.21676, 11.45479, 10.69252, 
    9.929964, 9.167146, 8.404083, 7.640796, 6.877304, 6.113627, 5.349786, 
    4.5858, 3.82169, 3.057476, 2.29318, 1.528821, 0.7644209, 1.272222e-14, 
    -0.7644209, -1.528821, -2.29318, -3.057476, -3.82169, -4.5858, -5.349786, 
    -6.113627, -6.877304, -7.640796, -8.404083, -9.167146, -9.929964, 
    -10.69252, -11.45479, -12.21676, -12.97841, -13.73972, -14.50067, 
    -15.26124, -16.02143, -16.7812, -17.54054, -18.29944, -19.05788, 
    -19.81585, -20.57332, -21.33028, -22.08672, -22.84263, -23.59798, 
    -24.35277, -25.10699, -25.86061, -26.61363, -27.36604, -28.11782, 
    -28.86897, -29.61947, -30.36931, -31.11849, -31.86699, -32.61481, 
    -33.36194, -34.10837, -34.8541, -35.59911, -36.34341,
  35.98892, 35.24767, 34.50594, 33.76374, 33.02107, 32.27793, 31.53433, 
    30.79028, 30.04578, 29.30084, 28.55546, 27.80966, 27.06343, 26.31679, 
    25.56974, 24.82229, 24.07445, 23.32623, 22.57764, 21.82868, 21.07937, 
    20.32972, 19.57973, 18.82941, 18.07879, 17.32786, 16.57663, 15.82513, 
    15.07335, 14.32132, 13.56903, 12.81652, 12.06378, 11.31083, 10.55768, 
    9.804344, 9.050837, 8.297169, 7.543353, 6.789403, 6.035332, 5.281153, 
    4.526879, 3.772523, 3.0181, 2.263623, 1.509105, 0.7545591, 1.272222e-14, 
    -0.7545591, -1.509105, -2.263623, -3.0181, -3.772523, -4.526879, 
    -5.281153, -6.035332, -6.789403, -7.543353, -8.297169, -9.050837, 
    -9.804344, -10.55768, -11.31083, -12.06378, -12.81652, -13.56903, 
    -14.32132, -15.07335, -15.82513, -16.57663, -17.32786, -18.07879, 
    -18.82941, -19.57973, -20.32972, -21.07937, -21.82868, -22.57764, 
    -23.32623, -24.07445, -24.82229, -25.56974, -26.31679, -27.06343, 
    -27.80966, -28.55546, -29.30084, -30.04578, -30.79028, -31.53433, 
    -32.27793, -33.02107, -33.76374, -34.50594, -35.24767, -35.98892,
  35.62921, 34.89117, 34.15289, 33.41436, 32.67561, 31.93662, 31.19741, 
    30.45796, 29.7183, 28.97841, 28.23831, 27.49799, 26.75747, 26.01674, 
    25.2758, 24.53467, 23.79335, 23.05183, 22.31014, 21.56826, 20.8262, 
    20.08398, 19.34159, 18.59904, 17.85633, 17.11348, 16.37048, 15.62734, 
    14.88407, 14.14067, 13.39715, 12.65351, 11.90976, 11.16591, 10.42197, 
    9.677926, 8.933801, 8.189597, 7.445321, 6.700978, 5.956575, 5.21212, 
    4.467618, 3.723077, 2.978501, 2.233899, 1.489277, 0.744642, 1.272222e-14, 
    -0.744642, -1.489277, -2.233899, -2.978501, -3.723077, -4.467618, 
    -5.21212, -5.956575, -6.700978, -7.445321, -8.189597, -8.933801, 
    -9.677926, -10.42197, -11.16591, -11.90976, -12.65351, -13.39715, 
    -14.14067, -14.88407, -15.62734, -16.37048, -17.11348, -17.85633, 
    -18.59904, -19.34159, -20.08398, -20.8262, -21.56826, -22.31014, 
    -23.05183, -23.79335, -24.53467, -25.2758, -26.01674, -26.75747, 
    -27.49799, -28.23831, -28.97841, -29.7183, -30.45796, -31.19741, 
    -31.93662, -32.67561, -33.41436, -34.15289, -34.89117, -35.62921,
  35.26439, 34.52972, 33.79504, 33.06036, 32.32569, 31.59101, 30.85634, 
    30.12167, 29.38699, 28.65232, 27.91764, 27.18297, 26.44829, 25.71362, 
    24.97894, 24.24427, 23.50959, 22.77492, 22.04024, 21.30557, 20.57089, 
    19.83622, 19.10155, 18.36687, 17.63219, 16.89752, 16.16285, 15.42817, 
    14.6935, 13.95882, 13.22415, 12.48947, 11.7548, 11.02012, 10.28545, 
    9.550773, 8.816097, 8.081423, 7.346748, 6.612073, 5.877398, 5.142724, 
    4.408049, 3.673374, 2.938699, 2.204024, 1.46935, 0.7346748, 1.272222e-14, 
    -0.7346748, -1.46935, -2.204024, -2.938699, -3.673374, -4.408049, 
    -5.142724, -5.877398, -6.612073, -7.346748, -8.081423, -8.816097, 
    -9.550773, -10.28545, -11.02012, -11.7548, -12.48947, -13.22415, 
    -13.95882, -14.6935, -15.42817, -16.16285, -16.89752, -17.63219, 
    -18.36687, -19.10155, -19.83622, -20.57089, -21.30557, -22.04024, 
    -22.77492, -23.50959, -24.24427, -24.97894, -25.71362, -26.44829, 
    -27.18297, -27.91764, -28.65232, -29.38699, -30.12167, -30.85634, 
    -31.59101, -32.32569, -33.06036, -33.79504, -34.52972, -35.26439 ;

 grid_lont =
  125.3905, 125.3905, 125.3906, 125.3906, 125.3906, 125.3907, 125.3907, 
    125.3907, 125.3908, 125.3908, 125.3908, 125.3908, 125.3909, 125.3909, 
    125.3909, 125.391, 125.391, 125.391, 125.391, 125.3911, 125.3911, 
    125.3911, 125.3911, 125.3911, 125.3912, 125.3912, 125.3912, 125.3912, 
    125.3912, 125.3912, 125.3913, 125.3913, 125.3913, 125.3913, 125.3913, 
    125.3913, 125.3913, 125.3913, 125.3913, 125.3914, 125.3914, 125.3914, 
    125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 
    125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 125.3914, 
    125.3914, 125.3913, 125.3913, 125.3913, 125.3913, 125.3913, 125.3913, 
    125.3913, 125.3913, 125.3913, 125.3912, 125.3912, 125.3912, 125.3912, 
    125.3912, 125.3912, 125.3911, 125.3911, 125.3911, 125.3911, 125.3911, 
    125.391, 125.391, 125.391, 125.391, 125.3909, 125.3909, 125.3909, 
    125.3908, 125.3908, 125.3908, 125.3908, 125.3907, 125.3907, 125.3907, 
    125.3906, 125.3906, 125.3906, 125.3905, 125.3905,
  126.1769, 126.1769, 126.1769, 126.177, 126.177, 126.177, 126.177, 126.1771, 
    126.1771, 126.1771, 126.1772, 126.1772, 126.1772, 126.1772, 126.1773, 
    126.1773, 126.1773, 126.1773, 126.1774, 126.1774, 126.1774, 126.1774, 
    126.1775, 126.1775, 126.1775, 126.1775, 126.1775, 126.1776, 126.1776, 
    126.1776, 126.1776, 126.1776, 126.1776, 126.1776, 126.1777, 126.1777, 
    126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 
    126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 
    126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 
    126.1777, 126.1777, 126.1777, 126.1777, 126.1777, 126.1776, 126.1776, 
    126.1776, 126.1776, 126.1776, 126.1776, 126.1776, 126.1775, 126.1775, 
    126.1775, 126.1775, 126.1775, 126.1774, 126.1774, 126.1774, 126.1774, 
    126.1773, 126.1773, 126.1773, 126.1773, 126.1772, 126.1772, 126.1772, 
    126.1772, 126.1771, 126.1771, 126.1771, 126.177, 126.177, 126.177, 
    126.177, 126.1769, 126.1769, 126.1769,
  126.9704, 126.9704, 126.9704, 126.9705, 126.9705, 126.9705, 126.9705, 
    126.9706, 126.9706, 126.9706, 126.9707, 126.9707, 126.9707, 126.9707, 
    126.9708, 126.9708, 126.9708, 126.9708, 126.9709, 126.9709, 126.9709, 
    126.9709, 126.971, 126.971, 126.971, 126.971, 126.971, 126.9711, 
    126.9711, 126.9711, 126.9711, 126.9711, 126.9711, 126.9711, 126.9712, 
    126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 
    126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 
    126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 
    126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9712, 126.9711, 
    126.9711, 126.9711, 126.9711, 126.9711, 126.9711, 126.9711, 126.971, 
    126.971, 126.971, 126.971, 126.971, 126.9709, 126.9709, 126.9709, 
    126.9709, 126.9708, 126.9708, 126.9708, 126.9708, 126.9707, 126.9707, 
    126.9707, 126.9707, 126.9706, 126.9706, 126.9706, 126.9705, 126.9705, 
    126.9705, 126.9705, 126.9704, 126.9704, 126.9704,
  127.7711, 127.7711, 127.7711, 127.7712, 127.7712, 127.7712, 127.7712, 
    127.7713, 127.7713, 127.7713, 127.7714, 127.7714, 127.7714, 127.7714, 
    127.7715, 127.7715, 127.7715, 127.7715, 127.7716, 127.7716, 127.7716, 
    127.7716, 127.7717, 127.7717, 127.7717, 127.7717, 127.7717, 127.7718, 
    127.7718, 127.7718, 127.7718, 127.7718, 127.7718, 127.7719, 127.7719, 
    127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 
    127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 
    127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 
    127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 127.7719, 
    127.7718, 127.7718, 127.7718, 127.7718, 127.7718, 127.7718, 127.7717, 
    127.7717, 127.7717, 127.7717, 127.7717, 127.7716, 127.7716, 127.7716, 
    127.7716, 127.7715, 127.7715, 127.7715, 127.7715, 127.7714, 127.7714, 
    127.7714, 127.7714, 127.7713, 127.7713, 127.7713, 127.7712, 127.7712, 
    127.7712, 127.7712, 127.7711, 127.7711, 127.7711,
  128.579, 128.5791, 128.5791, 128.5791, 128.5791, 128.5792, 128.5792, 
    128.5792, 128.5793, 128.5793, 128.5793, 128.5793, 128.5794, 128.5794, 
    128.5794, 128.5795, 128.5795, 128.5795, 128.5795, 128.5796, 128.5796, 
    128.5796, 128.5796, 128.5797, 128.5797, 128.5797, 128.5797, 128.5797, 
    128.5797, 128.5798, 128.5798, 128.5798, 128.5798, 128.5798, 128.5798, 
    128.5798, 128.5798, 128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 
    128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 
    128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 128.5799, 
    128.5799, 128.5799, 128.5799, 128.5798, 128.5798, 128.5798, 128.5798, 
    128.5798, 128.5798, 128.5798, 128.5798, 128.5797, 128.5797, 128.5797, 
    128.5797, 128.5797, 128.5797, 128.5796, 128.5796, 128.5796, 128.5796, 
    128.5795, 128.5795, 128.5795, 128.5795, 128.5794, 128.5794, 128.5794, 
    128.5793, 128.5793, 128.5793, 128.5793, 128.5792, 128.5792, 128.5792, 
    128.5791, 128.5791, 128.5791, 128.5791, 128.579,
  129.3943, 129.3943, 129.3943, 129.3944, 129.3944, 129.3944, 129.3945, 
    129.3945, 129.3945, 129.3946, 129.3946, 129.3946, 129.3946, 129.3947, 
    129.3947, 129.3947, 129.3947, 129.3948, 129.3948, 129.3948, 129.3949, 
    129.3949, 129.3949, 129.3949, 129.3949, 129.395, 129.395, 129.395, 
    129.395, 129.395, 129.3951, 129.3951, 129.3951, 129.3951, 129.3951, 
    129.3951, 129.3951, 129.3951, 129.3951, 129.3952, 129.3952, 129.3952, 
    129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 
    129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 129.3952, 
    129.3952, 129.3951, 129.3951, 129.3951, 129.3951, 129.3951, 129.3951, 
    129.3951, 129.3951, 129.3951, 129.395, 129.395, 129.395, 129.395, 
    129.395, 129.3949, 129.3949, 129.3949, 129.3949, 129.3949, 129.3948, 
    129.3948, 129.3948, 129.3947, 129.3947, 129.3947, 129.3947, 129.3946, 
    129.3946, 129.3946, 129.3946, 129.3945, 129.3945, 129.3945, 129.3944, 
    129.3944, 129.3944, 129.3943, 129.3943, 129.3943,
  130.2169, 130.2169, 130.2169, 130.217, 130.217, 130.217, 130.2171, 
    130.2171, 130.2171, 130.2172, 130.2172, 130.2172, 130.2172, 130.2173, 
    130.2173, 130.2173, 130.2173, 130.2174, 130.2174, 130.2174, 130.2175, 
    130.2175, 130.2175, 130.2175, 130.2175, 130.2176, 130.2176, 130.2176, 
    130.2176, 130.2176, 130.2177, 130.2177, 130.2177, 130.2177, 130.2177, 
    130.2177, 130.2177, 130.2177, 130.2177, 130.2178, 130.2178, 130.2178, 
    130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 
    130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 130.2178, 
    130.2178, 130.2177, 130.2177, 130.2177, 130.2177, 130.2177, 130.2177, 
    130.2177, 130.2177, 130.2177, 130.2176, 130.2176, 130.2176, 130.2176, 
    130.2176, 130.2175, 130.2175, 130.2175, 130.2175, 130.2175, 130.2174, 
    130.2174, 130.2174, 130.2173, 130.2173, 130.2173, 130.2173, 130.2172, 
    130.2172, 130.2172, 130.2172, 130.2171, 130.2171, 130.2171, 130.217, 
    130.217, 130.217, 130.2169, 130.2169, 130.2169,
  131.0469, 131.0469, 131.0469, 131.047, 131.047, 131.047, 131.047, 131.0471, 
    131.0471, 131.0471, 131.0471, 131.0472, 131.0472, 131.0472, 131.0473, 
    131.0473, 131.0473, 131.0473, 131.0474, 131.0474, 131.0474, 131.0474, 
    131.0475, 131.0475, 131.0475, 131.0475, 131.0475, 131.0476, 131.0476, 
    131.0476, 131.0476, 131.0476, 131.0477, 131.0477, 131.0477, 131.0477, 
    131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 
    131.0477, 131.0478, 131.0478, 131.0478, 131.0478, 131.0478, 131.0478, 
    131.0478, 131.0478, 131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 
    131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 131.0477, 
    131.0476, 131.0476, 131.0476, 131.0476, 131.0476, 131.0475, 131.0475, 
    131.0475, 131.0475, 131.0475, 131.0474, 131.0474, 131.0474, 131.0474, 
    131.0473, 131.0473, 131.0473, 131.0473, 131.0472, 131.0472, 131.0472, 
    131.0471, 131.0471, 131.0471, 131.0471, 131.047, 131.047, 131.047, 
    131.047, 131.0469, 131.0469, 131.0469,
  131.8842, 131.8842, 131.8843, 131.8843, 131.8843, 131.8844, 131.8844, 
    131.8844, 131.8845, 131.8845, 131.8845, 131.8845, 131.8846, 131.8846, 
    131.8846, 131.8846, 131.8847, 131.8847, 131.8847, 131.8848, 131.8848, 
    131.8848, 131.8848, 131.8848, 131.8849, 131.8849, 131.8849, 131.8849, 
    131.8849, 131.885, 131.885, 131.885, 131.885, 131.885, 131.885, 131.885, 
    131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 
    131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 
    131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 131.8851, 
    131.8851, 131.8851, 131.8851, 131.885, 131.885, 131.885, 131.885, 
    131.885, 131.885, 131.885, 131.8849, 131.8849, 131.8849, 131.8849, 
    131.8849, 131.8848, 131.8848, 131.8848, 131.8848, 131.8848, 131.8847, 
    131.8847, 131.8847, 131.8846, 131.8846, 131.8846, 131.8846, 131.8845, 
    131.8845, 131.8845, 131.8845, 131.8844, 131.8844, 131.8844, 131.8843, 
    131.8843, 131.8843, 131.8842, 131.8842,
  132.729, 132.729, 132.729, 132.7291, 132.7291, 132.7291, 132.7292, 
    132.7292, 132.7292, 132.7292, 132.7293, 132.7293, 132.7293, 132.7294, 
    132.7294, 132.7294, 132.7294, 132.7295, 132.7295, 132.7295, 132.7295, 
    132.7296, 132.7296, 132.7296, 132.7296, 132.7296, 132.7297, 132.7297, 
    132.7297, 132.7297, 132.7297, 132.7298, 132.7298, 132.7298, 132.7298, 
    132.7298, 132.7298, 132.7298, 132.7298, 132.7299, 132.7299, 132.7299, 
    132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 
    132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 132.7299, 
    132.7299, 132.7298, 132.7298, 132.7298, 132.7298, 132.7298, 132.7298, 
    132.7298, 132.7298, 132.7297, 132.7297, 132.7297, 132.7297, 132.7297, 
    132.7296, 132.7296, 132.7296, 132.7296, 132.7296, 132.7295, 132.7295, 
    132.7295, 132.7295, 132.7294, 132.7294, 132.7294, 132.7294, 132.7293, 
    132.7293, 132.7293, 132.7292, 132.7292, 132.7292, 132.7292, 132.7291, 
    132.7291, 132.7291, 132.729, 132.729, 132.729,
  133.5812, 133.5812, 133.5812, 133.5813, 133.5813, 133.5813, 133.5813, 
    133.5814, 133.5814, 133.5814, 133.5815, 133.5815, 133.5815, 133.5815, 
    133.5816, 133.5816, 133.5816, 133.5816, 133.5817, 133.5817, 133.5817, 
    133.5817, 133.5818, 133.5818, 133.5818, 133.5818, 133.5818, 133.5819, 
    133.5819, 133.5819, 133.5819, 133.5819, 133.582, 133.582, 133.582, 
    133.582, 133.582, 133.582, 133.582, 133.582, 133.582, 133.582, 133.582, 
    133.5821, 133.5821, 133.5821, 133.5821, 133.5821, 133.5821, 133.5821, 
    133.5821, 133.5821, 133.5821, 133.582, 133.582, 133.582, 133.582, 
    133.582, 133.582, 133.582, 133.582, 133.582, 133.582, 133.582, 133.5819, 
    133.5819, 133.5819, 133.5819, 133.5819, 133.5818, 133.5818, 133.5818, 
    133.5818, 133.5818, 133.5817, 133.5817, 133.5817, 133.5817, 133.5816, 
    133.5816, 133.5816, 133.5816, 133.5815, 133.5815, 133.5815, 133.5815, 
    133.5814, 133.5814, 133.5814, 133.5813, 133.5813, 133.5813, 133.5813, 
    133.5812, 133.5812, 133.5812,
  134.4408, 134.4408, 134.4408, 134.4408, 134.4409, 134.4409, 134.4409, 
    134.4409, 134.441, 134.441, 134.441, 134.4411, 134.4411, 134.4411, 
    134.4411, 134.4412, 134.4412, 134.4412, 134.4413, 134.4413, 134.4413, 
    134.4413, 134.4413, 134.4414, 134.4414, 134.4414, 134.4414, 134.4415, 
    134.4415, 134.4415, 134.4415, 134.4415, 134.4415, 134.4416, 134.4416, 
    134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 
    134.4416, 134.4417, 134.4417, 134.4417, 134.4417, 134.4417, 134.4417, 
    134.4417, 134.4417, 134.4417, 134.4417, 134.4416, 134.4416, 134.4416, 
    134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 134.4416, 
    134.4415, 134.4415, 134.4415, 134.4415, 134.4415, 134.4415, 134.4414, 
    134.4414, 134.4414, 134.4414, 134.4413, 134.4413, 134.4413, 134.4413, 
    134.4413, 134.4412, 134.4412, 134.4412, 134.4411, 134.4411, 134.4411, 
    134.4411, 134.441, 134.441, 134.441, 134.4409, 134.4409, 134.4409, 
    134.4409, 134.4408, 134.4408, 134.4408, 134.4408,
  135.3077, 135.3078, 135.3078, 135.3078, 135.3079, 135.3079, 135.3079, 
    135.308, 135.308, 135.308, 135.308, 135.3081, 135.3081, 135.3081, 
    135.3082, 135.3082, 135.3082, 135.3082, 135.3082, 135.3083, 135.3083, 
    135.3083, 135.3083, 135.3084, 135.3084, 135.3084, 135.3084, 135.3084, 
    135.3085, 135.3085, 135.3085, 135.3085, 135.3085, 135.3085, 135.3086, 
    135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 
    135.3086, 135.3086, 135.3086, 135.3087, 135.3087, 135.3087, 135.3087, 
    135.3087, 135.3087, 135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 
    135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 135.3086, 135.3085, 
    135.3085, 135.3085, 135.3085, 135.3085, 135.3085, 135.3084, 135.3084, 
    135.3084, 135.3084, 135.3084, 135.3083, 135.3083, 135.3083, 135.3083, 
    135.3082, 135.3082, 135.3082, 135.3082, 135.3082, 135.3081, 135.3081, 
    135.3081, 135.308, 135.308, 135.308, 135.308, 135.3079, 135.3079, 
    135.3079, 135.3078, 135.3078, 135.3078, 135.3077,
  136.1821, 136.1822, 136.1822, 136.1822, 136.1823, 136.1823, 136.1823, 
    136.1823, 136.1824, 136.1824, 136.1824, 136.1824, 136.1825, 136.1825, 
    136.1825, 136.1826, 136.1826, 136.1826, 136.1826, 136.1827, 136.1827, 
    136.1827, 136.1827, 136.1828, 136.1828, 136.1828, 136.1828, 136.1828, 
    136.1828, 136.1829, 136.1829, 136.1829, 136.1829, 136.1829, 136.1829, 
    136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 
    136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 
    136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 136.183, 
    136.183, 136.183, 136.1829, 136.1829, 136.1829, 136.1829, 136.1829, 
    136.1829, 136.1828, 136.1828, 136.1828, 136.1828, 136.1828, 136.1828, 
    136.1827, 136.1827, 136.1827, 136.1827, 136.1826, 136.1826, 136.1826, 
    136.1826, 136.1825, 136.1825, 136.1825, 136.1824, 136.1824, 136.1824, 
    136.1824, 136.1823, 136.1823, 136.1823, 136.1823, 136.1822, 136.1822, 
    136.1822, 136.1821,
  137.0639, 137.0639, 137.0639, 137.064, 137.064, 137.064, 137.0641, 
    137.0641, 137.0641, 137.0641, 137.0642, 137.0642, 137.0642, 137.0642, 
    137.0643, 137.0643, 137.0643, 137.0643, 137.0644, 137.0644, 137.0644, 
    137.0645, 137.0645, 137.0645, 137.0645, 137.0645, 137.0646, 137.0646, 
    137.0646, 137.0646, 137.0646, 137.0646, 137.0647, 137.0647, 137.0647, 
    137.0647, 137.0647, 137.0647, 137.0647, 137.0647, 137.0647, 137.0648, 
    137.0648, 137.0648, 137.0648, 137.0648, 137.0648, 137.0648, 137.0648, 
    137.0648, 137.0648, 137.0648, 137.0648, 137.0648, 137.0648, 137.0647, 
    137.0647, 137.0647, 137.0647, 137.0647, 137.0647, 137.0647, 137.0647, 
    137.0647, 137.0646, 137.0646, 137.0646, 137.0646, 137.0646, 137.0646, 
    137.0645, 137.0645, 137.0645, 137.0645, 137.0645, 137.0644, 137.0644, 
    137.0644, 137.0643, 137.0643, 137.0643, 137.0643, 137.0642, 137.0642, 
    137.0642, 137.0642, 137.0641, 137.0641, 137.0641, 137.0641, 137.064, 
    137.064, 137.064, 137.0639, 137.0639, 137.0639,
  137.953, 137.953, 137.953, 137.953, 137.9531, 137.9531, 137.9531, 137.9532, 
    137.9532, 137.9532, 137.9532, 137.9533, 137.9533, 137.9533, 137.9533, 
    137.9534, 137.9534, 137.9534, 137.9534, 137.9535, 137.9535, 137.9535, 
    137.9535, 137.9536, 137.9536, 137.9536, 137.9536, 137.9536, 137.9537, 
    137.9537, 137.9537, 137.9537, 137.9537, 137.9537, 137.9538, 137.9538, 
    137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 
    137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 
    137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 
    137.9538, 137.9538, 137.9538, 137.9538, 137.9538, 137.9537, 137.9537, 
    137.9537, 137.9537, 137.9537, 137.9537, 137.9536, 137.9536, 137.9536, 
    137.9536, 137.9536, 137.9535, 137.9535, 137.9535, 137.9535, 137.9534, 
    137.9534, 137.9534, 137.9534, 137.9533, 137.9533, 137.9533, 137.9533, 
    137.9532, 137.9532, 137.9532, 137.9532, 137.9531, 137.9531, 137.9531, 
    137.953, 137.953, 137.953, 137.953,
  138.8493, 138.8493, 138.8494, 138.8494, 138.8494, 138.8494, 138.8495, 
    138.8495, 138.8495, 138.8496, 138.8496, 138.8496, 138.8496, 138.8497, 
    138.8497, 138.8497, 138.8497, 138.8498, 138.8498, 138.8498, 138.8498, 
    138.8499, 138.8499, 138.8499, 138.8499, 138.8499, 138.85, 138.85, 138.85, 
    138.85, 138.85, 138.8501, 138.8501, 138.8501, 138.8501, 138.8501, 
    138.8501, 138.8501, 138.8501, 138.8502, 138.8502, 138.8502, 138.8502, 
    138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 
    138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 138.8502, 
    138.8501, 138.8501, 138.8501, 138.8501, 138.8501, 138.8501, 138.8501, 
    138.8501, 138.85, 138.85, 138.85, 138.85, 138.85, 138.8499, 138.8499, 
    138.8499, 138.8499, 138.8499, 138.8498, 138.8498, 138.8498, 138.8498, 
    138.8497, 138.8497, 138.8497, 138.8497, 138.8496, 138.8496, 138.8496, 
    138.8496, 138.8495, 138.8495, 138.8495, 138.8494, 138.8494, 138.8494, 
    138.8494, 138.8493, 138.8493,
  139.7529, 139.7529, 139.7529, 139.753, 139.753, 139.753, 139.7531, 
    139.7531, 139.7531, 139.7531, 139.7532, 139.7532, 139.7532, 139.7532, 
    139.7533, 139.7533, 139.7533, 139.7533, 139.7534, 139.7534, 139.7534, 
    139.7534, 139.7534, 139.7535, 139.7535, 139.7535, 139.7535, 139.7536, 
    139.7536, 139.7536, 139.7536, 139.7536, 139.7536, 139.7537, 139.7537, 
    139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 
    139.7538, 139.7538, 139.7538, 139.7538, 139.7538, 139.7538, 139.7538, 
    139.7538, 139.7538, 139.7538, 139.7538, 139.7538, 139.7537, 139.7537, 
    139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 139.7537, 
    139.7536, 139.7536, 139.7536, 139.7536, 139.7536, 139.7536, 139.7535, 
    139.7535, 139.7535, 139.7535, 139.7534, 139.7534, 139.7534, 139.7534, 
    139.7534, 139.7533, 139.7533, 139.7533, 139.7533, 139.7532, 139.7532, 
    139.7532, 139.7532, 139.7531, 139.7531, 139.7531, 139.7531, 139.753, 
    139.753, 139.753, 139.7529, 139.7529, 139.7529,
  140.6636, 140.6637, 140.6637, 140.6637, 140.6637, 140.6638, 140.6638, 
    140.6638, 140.6638, 140.6639, 140.6639, 140.6639, 140.6639, 140.664, 
    140.664, 140.664, 140.664, 140.6641, 140.6641, 140.6641, 140.6641, 
    140.6642, 140.6642, 140.6642, 140.6642, 140.6642, 140.6643, 140.6643, 
    140.6643, 140.6643, 140.6643, 140.6644, 140.6644, 140.6644, 140.6644, 
    140.6644, 140.6644, 140.6644, 140.6644, 140.6644, 140.6645, 140.6645, 
    140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 
    140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 140.6645, 
    140.6644, 140.6644, 140.6644, 140.6644, 140.6644, 140.6644, 140.6644, 
    140.6644, 140.6644, 140.6643, 140.6643, 140.6643, 140.6643, 140.6643, 
    140.6642, 140.6642, 140.6642, 140.6642, 140.6642, 140.6641, 140.6641, 
    140.6641, 140.6641, 140.664, 140.664, 140.664, 140.664, 140.6639, 
    140.6639, 140.6639, 140.6639, 140.6638, 140.6638, 140.6638, 140.6638, 
    140.6637, 140.6637, 140.6637, 140.6637, 140.6636,
  141.5814, 141.5815, 141.5815, 141.5815, 141.5815, 141.5816, 141.5816, 
    141.5816, 141.5816, 141.5817, 141.5817, 141.5817, 141.5818, 141.5818, 
    141.5818, 141.5818, 141.5818, 141.5819, 141.5819, 141.5819, 141.5819, 
    141.582, 141.582, 141.582, 141.582, 141.582, 141.5821, 141.5821, 
    141.5821, 141.5821, 141.5821, 141.5822, 141.5822, 141.5822, 141.5822, 
    141.5822, 141.5822, 141.5822, 141.5822, 141.5823, 141.5823, 141.5823, 
    141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 
    141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 141.5823, 
    141.5823, 141.5822, 141.5822, 141.5822, 141.5822, 141.5822, 141.5822, 
    141.5822, 141.5822, 141.5821, 141.5821, 141.5821, 141.5821, 141.5821, 
    141.582, 141.582, 141.582, 141.582, 141.582, 141.5819, 141.5819, 
    141.5819, 141.5819, 141.5818, 141.5818, 141.5818, 141.5818, 141.5818, 
    141.5817, 141.5817, 141.5817, 141.5816, 141.5816, 141.5816, 141.5816, 
    141.5815, 141.5815, 141.5815, 141.5815, 141.5814,
  142.5062, 142.5063, 142.5063, 142.5063, 142.5063, 142.5064, 142.5064, 
    142.5064, 142.5065, 142.5065, 142.5065, 142.5065, 142.5065, 142.5066, 
    142.5066, 142.5066, 142.5067, 142.5067, 142.5067, 142.5067, 142.5067, 
    142.5068, 142.5068, 142.5068, 142.5068, 142.5069, 142.5069, 142.5069, 
    142.5069, 142.5069, 142.5069, 142.507, 142.507, 142.507, 142.507, 
    142.507, 142.507, 142.507, 142.507, 142.507, 142.5071, 142.5071, 
    142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 
    142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 142.5071, 
    142.507, 142.507, 142.507, 142.507, 142.507, 142.507, 142.507, 142.507, 
    142.507, 142.5069, 142.5069, 142.5069, 142.5069, 142.5069, 142.5069, 
    142.5068, 142.5068, 142.5068, 142.5068, 142.5067, 142.5067, 142.5067, 
    142.5067, 142.5067, 142.5066, 142.5066, 142.5066, 142.5065, 142.5065, 
    142.5065, 142.5065, 142.5065, 142.5064, 142.5064, 142.5064, 142.5063, 
    142.5063, 142.5063, 142.5063, 142.5062,
  143.4379, 143.438, 143.438, 143.438, 143.438, 143.4381, 143.4381, 143.4381, 
    143.4381, 143.4382, 143.4382, 143.4382, 143.4382, 143.4383, 143.4383, 
    143.4383, 143.4383, 143.4384, 143.4384, 143.4384, 143.4384, 143.4385, 
    143.4385, 143.4385, 143.4385, 143.4385, 143.4386, 143.4386, 143.4386, 
    143.4386, 143.4386, 143.4386, 143.4387, 143.4387, 143.4387, 143.4387, 
    143.4387, 143.4387, 143.4387, 143.4387, 143.4388, 143.4388, 143.4388, 
    143.4388, 143.4388, 143.4388, 143.4388, 143.4388, 143.4388, 143.4388, 
    143.4388, 143.4388, 143.4388, 143.4388, 143.4388, 143.4388, 143.4387, 
    143.4387, 143.4387, 143.4387, 143.4387, 143.4387, 143.4387, 143.4387, 
    143.4386, 143.4386, 143.4386, 143.4386, 143.4386, 143.4386, 143.4385, 
    143.4385, 143.4385, 143.4385, 143.4385, 143.4384, 143.4384, 143.4384, 
    143.4384, 143.4383, 143.4383, 143.4383, 143.4383, 143.4382, 143.4382, 
    143.4382, 143.4382, 143.4381, 143.4381, 143.4381, 143.4381, 143.438, 
    143.438, 143.438, 143.438, 143.4379,
  144.3764, 144.3764, 144.3765, 144.3765, 144.3765, 144.3765, 144.3766, 
    144.3766, 144.3766, 144.3766, 144.3767, 144.3767, 144.3767, 144.3767, 
    144.3768, 144.3768, 144.3768, 144.3768, 144.3769, 144.3769, 144.3769, 
    144.3769, 144.377, 144.377, 144.377, 144.377, 144.377, 144.377, 144.3771, 
    144.3771, 144.3771, 144.3771, 144.3771, 144.3771, 144.3772, 144.3772, 
    144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 
    144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 
    144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 
    144.3772, 144.3772, 144.3772, 144.3772, 144.3772, 144.3771, 144.3771, 
    144.3771, 144.3771, 144.3771, 144.3771, 144.377, 144.377, 144.377, 
    144.377, 144.377, 144.377, 144.3769, 144.3769, 144.3769, 144.3769, 
    144.3768, 144.3768, 144.3768, 144.3768, 144.3767, 144.3767, 144.3767, 
    144.3767, 144.3766, 144.3766, 144.3766, 144.3766, 144.3765, 144.3765, 
    144.3765, 144.3765, 144.3764, 144.3764,
  145.3216, 145.3216, 145.3216, 145.3216, 145.3217, 145.3217, 145.3217, 
    145.3217, 145.3217, 145.3218, 145.3218, 145.3218, 145.3219, 145.3219, 
    145.3219, 145.3219, 145.3219, 145.322, 145.322, 145.322, 145.322, 
    145.3221, 145.3221, 145.3221, 145.3221, 145.3221, 145.3222, 145.3222, 
    145.3222, 145.3222, 145.3222, 145.3222, 145.3223, 145.3223, 145.3223, 
    145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 
    145.3223, 145.3224, 145.3224, 145.3224, 145.3224, 145.3224, 145.3224, 
    145.3224, 145.3224, 145.3224, 145.3224, 145.3223, 145.3223, 145.3223, 
    145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 145.3223, 
    145.3223, 145.3222, 145.3222, 145.3222, 145.3222, 145.3222, 145.3222, 
    145.3221, 145.3221, 145.3221, 145.3221, 145.3221, 145.322, 145.322, 
    145.322, 145.322, 145.3219, 145.3219, 145.3219, 145.3219, 145.3219, 
    145.3218, 145.3218, 145.3218, 145.3217, 145.3217, 145.3217, 145.3217, 
    145.3217, 145.3216, 145.3216, 145.3216, 145.3216,
  146.2732, 146.2732, 146.2733, 146.2733, 146.2733, 146.2733, 146.2734, 
    146.2734, 146.2734, 146.2734, 146.2735, 146.2735, 146.2735, 146.2735, 
    146.2736, 146.2736, 146.2736, 146.2736, 146.2736, 146.2737, 146.2737, 
    146.2737, 146.2737, 146.2737, 146.2738, 146.2738, 146.2738, 146.2738, 
    146.2738, 146.2738, 146.2739, 146.2739, 146.2739, 146.2739, 146.2739, 
    146.2739, 146.2739, 146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 
    146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 
    146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 146.274, 
    146.2739, 146.2739, 146.2739, 146.2739, 146.2739, 146.2739, 146.2739, 
    146.2738, 146.2738, 146.2738, 146.2738, 146.2738, 146.2738, 146.2737, 
    146.2737, 146.2737, 146.2737, 146.2737, 146.2736, 146.2736, 146.2736, 
    146.2736, 146.2736, 146.2735, 146.2735, 146.2735, 146.2735, 146.2734, 
    146.2734, 146.2734, 146.2734, 146.2733, 146.2733, 146.2733, 146.2733, 
    146.2732, 146.2732,
  147.2313, 147.2313, 147.2313, 147.2313, 147.2314, 147.2314, 147.2314, 
    147.2314, 147.2314, 147.2315, 147.2315, 147.2315, 147.2315, 147.2316, 
    147.2316, 147.2316, 147.2316, 147.2316, 147.2317, 147.2317, 147.2317, 
    147.2317, 147.2318, 147.2318, 147.2318, 147.2318, 147.2318, 147.2318, 
    147.2319, 147.2319, 147.2319, 147.2319, 147.2319, 147.2319, 147.2319, 
    147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 
    147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 
    147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 147.232, 
    147.232, 147.232, 147.2319, 147.2319, 147.2319, 147.2319, 147.2319, 
    147.2319, 147.2319, 147.2318, 147.2318, 147.2318, 147.2318, 147.2318, 
    147.2318, 147.2317, 147.2317, 147.2317, 147.2317, 147.2316, 147.2316, 
    147.2316, 147.2316, 147.2316, 147.2315, 147.2315, 147.2315, 147.2315, 
    147.2314, 147.2314, 147.2314, 147.2314, 147.2314, 147.2313, 147.2313, 
    147.2313, 147.2313,
  148.1955, 148.1955, 148.1956, 148.1956, 148.1956, 148.1956, 148.1957, 
    148.1957, 148.1957, 148.1957, 148.1957, 148.1958, 148.1958, 148.1958, 
    148.1958, 148.1959, 148.1959, 148.1959, 148.1959, 148.1959, 148.196, 
    148.196, 148.196, 148.196, 148.196, 148.196, 148.1961, 148.1961, 
    148.1961, 148.1961, 148.1961, 148.1962, 148.1962, 148.1962, 148.1962, 
    148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 
    148.1963, 148.1963, 148.1963, 148.1963, 148.1963, 148.1963, 148.1963, 
    148.1963, 148.1963, 148.1963, 148.1963, 148.1963, 148.1962, 148.1962, 
    148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 148.1962, 
    148.1962, 148.1962, 148.1961, 148.1961, 148.1961, 148.1961, 148.1961, 
    148.196, 148.196, 148.196, 148.196, 148.196, 148.196, 148.1959, 148.1959, 
    148.1959, 148.1959, 148.1959, 148.1958, 148.1958, 148.1958, 148.1958, 
    148.1957, 148.1957, 148.1957, 148.1957, 148.1957, 148.1956, 148.1956, 
    148.1956, 148.1956, 148.1955, 148.1955,
  149.1658, 149.1658, 149.1659, 149.1659, 149.1659, 149.1659, 149.166, 
    149.166, 149.166, 149.166, 149.166, 149.1661, 149.1661, 149.1661, 
    149.1661, 149.1662, 149.1662, 149.1662, 149.1662, 149.1662, 149.1662, 
    149.1663, 149.1663, 149.1663, 149.1663, 149.1663, 149.1664, 149.1664, 
    149.1664, 149.1664, 149.1664, 149.1664, 149.1664, 149.1665, 149.1665, 
    149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 
    149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 
    149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 
    149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 149.1665, 
    149.1664, 149.1664, 149.1664, 149.1664, 149.1664, 149.1664, 149.1664, 
    149.1663, 149.1663, 149.1663, 149.1663, 149.1663, 149.1662, 149.1662, 
    149.1662, 149.1662, 149.1662, 149.1662, 149.1661, 149.1661, 149.1661, 
    149.1661, 149.166, 149.166, 149.166, 149.166, 149.166, 149.1659, 
    149.1659, 149.1659, 149.1659, 149.1658, 149.1658,
  150.142, 150.142, 150.142, 150.1421, 150.1421, 150.1421, 150.1421, 
    150.1422, 150.1422, 150.1422, 150.1422, 150.1422, 150.1423, 150.1423, 
    150.1423, 150.1423, 150.1423, 150.1423, 150.1424, 150.1424, 150.1424, 
    150.1424, 150.1424, 150.1425, 150.1425, 150.1425, 150.1425, 150.1425, 
    150.1425, 150.1426, 150.1426, 150.1426, 150.1426, 150.1426, 150.1426, 
    150.1426, 150.1426, 150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 
    150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 
    150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 150.1427, 
    150.1427, 150.1427, 150.1427, 150.1426, 150.1426, 150.1426, 150.1426, 
    150.1426, 150.1426, 150.1426, 150.1426, 150.1425, 150.1425, 150.1425, 
    150.1425, 150.1425, 150.1425, 150.1424, 150.1424, 150.1424, 150.1424, 
    150.1424, 150.1423, 150.1423, 150.1423, 150.1423, 150.1423, 150.1423, 
    150.1422, 150.1422, 150.1422, 150.1422, 150.1422, 150.1421, 150.1421, 
    150.1421, 150.1421, 150.142, 150.142, 150.142,
  151.1239, 151.1239, 151.1239, 151.1239, 151.1239, 151.1239, 151.124, 
    151.124, 151.124, 151.124, 151.1241, 151.1241, 151.1241, 151.1241, 
    151.1241, 151.1241, 151.1242, 151.1242, 151.1242, 151.1242, 151.1242, 
    151.1243, 151.1243, 151.1243, 151.1243, 151.1243, 151.1243, 151.1244, 
    151.1244, 151.1244, 151.1244, 151.1244, 151.1244, 151.1244, 151.1245, 
    151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 
    151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 
    151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 
    151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1245, 151.1244, 
    151.1244, 151.1244, 151.1244, 151.1244, 151.1244, 151.1244, 151.1243, 
    151.1243, 151.1243, 151.1243, 151.1243, 151.1243, 151.1242, 151.1242, 
    151.1242, 151.1242, 151.1242, 151.1241, 151.1241, 151.1241, 151.1241, 
    151.1241, 151.1241, 151.124, 151.124, 151.124, 151.124, 151.1239, 
    151.1239, 151.1239, 151.1239, 151.1239, 151.1239,
  152.1112, 152.1112, 152.1112, 152.1112, 152.1112, 152.1113, 152.1113, 
    152.1113, 152.1113, 152.1113, 152.1113, 152.1114, 152.1114, 152.1114, 
    152.1114, 152.1115, 152.1115, 152.1115, 152.1115, 152.1115, 152.1115, 
    152.1116, 152.1116, 152.1116, 152.1116, 152.1116, 152.1116, 152.1116, 
    152.1117, 152.1117, 152.1117, 152.1117, 152.1117, 152.1117, 152.1117, 
    152.1117, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 
    152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 
    152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 152.1118, 
    152.1118, 152.1118, 152.1118, 152.1118, 152.1117, 152.1117, 152.1117, 
    152.1117, 152.1117, 152.1117, 152.1117, 152.1117, 152.1116, 152.1116, 
    152.1116, 152.1116, 152.1116, 152.1116, 152.1116, 152.1115, 152.1115, 
    152.1115, 152.1115, 152.1115, 152.1115, 152.1114, 152.1114, 152.1114, 
    152.1114, 152.1113, 152.1113, 152.1113, 152.1113, 152.1113, 152.1113, 
    152.1112, 152.1112, 152.1112, 152.1112, 152.1112,
  153.1037, 153.1037, 153.1037, 153.1038, 153.1038, 153.1038, 153.1038, 
    153.1038, 153.1039, 153.1039, 153.1039, 153.1039, 153.1039, 153.1039, 
    153.104, 153.104, 153.104, 153.104, 153.104, 153.104, 153.1041, 153.1041, 
    153.1041, 153.1041, 153.1041, 153.1042, 153.1042, 153.1042, 153.1042, 
    153.1042, 153.1042, 153.1042, 153.1042, 153.1042, 153.1043, 153.1043, 
    153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 
    153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 
    153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 
    153.1043, 153.1043, 153.1043, 153.1043, 153.1043, 153.1042, 153.1042, 
    153.1042, 153.1042, 153.1042, 153.1042, 153.1042, 153.1042, 153.1042, 
    153.1041, 153.1041, 153.1041, 153.1041, 153.1041, 153.104, 153.104, 
    153.104, 153.104, 153.104, 153.104, 153.1039, 153.1039, 153.1039, 
    153.1039, 153.1039, 153.1039, 153.1038, 153.1038, 153.1038, 153.1038, 
    153.1038, 153.1037, 153.1037, 153.1037,
  154.1013, 154.1013, 154.1013, 154.1013, 154.1013, 154.1014, 154.1014, 
    154.1014, 154.1014, 154.1014, 154.1015, 154.1015, 154.1015, 154.1015, 
    154.1015, 154.1015, 154.1016, 154.1016, 154.1016, 154.1016, 154.1016, 
    154.1016, 154.1017, 154.1017, 154.1017, 154.1017, 154.1017, 154.1017, 
    154.1017, 154.1018, 154.1018, 154.1018, 154.1018, 154.1018, 154.1018, 
    154.1018, 154.1018, 154.1018, 154.1018, 154.1019, 154.1019, 154.1019, 
    154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 
    154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 154.1019, 
    154.1019, 154.1018, 154.1018, 154.1018, 154.1018, 154.1018, 154.1018, 
    154.1018, 154.1018, 154.1018, 154.1018, 154.1017, 154.1017, 154.1017, 
    154.1017, 154.1017, 154.1017, 154.1017, 154.1016, 154.1016, 154.1016, 
    154.1016, 154.1016, 154.1016, 154.1015, 154.1015, 154.1015, 154.1015, 
    154.1015, 154.1015, 154.1014, 154.1014, 154.1014, 154.1014, 154.1014, 
    154.1013, 154.1013, 154.1013, 154.1013, 154.1013,
  155.1036, 155.1037, 155.1037, 155.1037, 155.1037, 155.1037, 155.1037, 
    155.1037, 155.1038, 155.1038, 155.1038, 155.1038, 155.1038, 155.1039, 
    155.1039, 155.1039, 155.1039, 155.1039, 155.1039, 155.1039, 155.104, 
    155.104, 155.104, 155.104, 155.104, 155.104, 155.104, 155.104, 155.1041, 
    155.1041, 155.1041, 155.1041, 155.1041, 155.1041, 155.1041, 155.1041, 
    155.1041, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 
    155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 
    155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 155.1042, 
    155.1042, 155.1042, 155.1041, 155.1041, 155.1041, 155.1041, 155.1041, 
    155.1041, 155.1041, 155.1041, 155.1041, 155.104, 155.104, 155.104, 
    155.104, 155.104, 155.104, 155.104, 155.104, 155.1039, 155.1039, 
    155.1039, 155.1039, 155.1039, 155.1039, 155.1039, 155.1038, 155.1038, 
    155.1038, 155.1038, 155.1038, 155.1037, 155.1037, 155.1037, 155.1037, 
    155.1037, 155.1037, 155.1037, 155.1036,
  156.1105, 156.1105, 156.1105, 156.1106, 156.1106, 156.1106, 156.1106, 
    156.1106, 156.1106, 156.1107, 156.1107, 156.1107, 156.1107, 156.1107, 
    156.1107, 156.1107, 156.1108, 156.1108, 156.1108, 156.1108, 156.1108, 
    156.1108, 156.1108, 156.1109, 156.1109, 156.1109, 156.1109, 156.1109, 
    156.1109, 156.1109, 156.1109, 156.1109, 156.111, 156.111, 156.111, 
    156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 
    156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 
    156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 156.111, 
    156.111, 156.111, 156.111, 156.111, 156.111, 156.1109, 156.1109, 
    156.1109, 156.1109, 156.1109, 156.1109, 156.1109, 156.1109, 156.1109, 
    156.1108, 156.1108, 156.1108, 156.1108, 156.1108, 156.1108, 156.1108, 
    156.1107, 156.1107, 156.1107, 156.1107, 156.1107, 156.1107, 156.1107, 
    156.1106, 156.1106, 156.1106, 156.1106, 156.1106, 156.1106, 156.1105, 
    156.1105, 156.1105,
  157.1217, 157.1217, 157.1217, 157.1217, 157.1217, 157.1217, 157.1217, 
    157.1217, 157.1218, 157.1218, 157.1218, 157.1218, 157.1218, 157.1218, 
    157.1219, 157.1219, 157.1219, 157.1219, 157.1219, 157.1219, 157.1219, 
    157.1219, 157.122, 157.122, 157.122, 157.122, 157.122, 157.122, 157.122, 
    157.122, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 
    157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 
    157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 
    157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 
    157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 157.1221, 
    157.1221, 157.1221, 157.122, 157.122, 157.122, 157.122, 157.122, 157.122, 
    157.122, 157.122, 157.1219, 157.1219, 157.1219, 157.1219, 157.1219, 
    157.1219, 157.1219, 157.1219, 157.1218, 157.1218, 157.1218, 157.1218, 
    157.1218, 157.1218, 157.1217, 157.1217, 157.1217, 157.1217, 157.1217, 
    157.1217, 157.1217, 157.1217,
  158.1368, 158.1368, 158.1368, 158.1368, 158.1368, 158.1368, 158.1369, 
    158.1369, 158.1369, 158.1369, 158.1369, 158.1369, 158.1369, 158.1369, 
    158.137, 158.137, 158.137, 158.137, 158.137, 158.137, 158.137, 158.1371, 
    158.1371, 158.1371, 158.1371, 158.1371, 158.1371, 158.1371, 158.1371, 
    158.1371, 158.1371, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 
    158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 
    158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 
    158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 
    158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 158.1372, 
    158.1372, 158.1371, 158.1371, 158.1371, 158.1371, 158.1371, 158.1371, 
    158.1371, 158.1371, 158.1371, 158.1371, 158.137, 158.137, 158.137, 
    158.137, 158.137, 158.137, 158.137, 158.1369, 158.1369, 158.1369, 
    158.1369, 158.1369, 158.1369, 158.1369, 158.1369, 158.1368, 158.1368, 
    158.1368, 158.1368, 158.1368, 158.1368,
  159.1556, 159.1556, 159.1556, 159.1557, 159.1557, 159.1557, 159.1557, 
    159.1557, 159.1557, 159.1557, 159.1557, 159.1557, 159.1558, 159.1558, 
    159.1558, 159.1558, 159.1558, 159.1558, 159.1558, 159.1559, 159.1559, 
    159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 
    159.1559, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 
    159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 
    159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 
    159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 
    159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.156, 159.1559, 
    159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 159.1559, 
    159.1559, 159.1559, 159.1558, 159.1558, 159.1558, 159.1558, 159.1558, 
    159.1558, 159.1558, 159.1557, 159.1557, 159.1557, 159.1557, 159.1557, 
    159.1557, 159.1557, 159.1557, 159.1557, 159.1556, 159.1556, 159.1556,
  160.1779, 160.1779, 160.1779, 160.1779, 160.1779, 160.1779, 160.1779, 
    160.1779, 160.178, 160.178, 160.178, 160.178, 160.178, 160.178, 160.178, 
    160.178, 160.1781, 160.1781, 160.1781, 160.1781, 160.1781, 160.1781, 
    160.1781, 160.1781, 160.1781, 160.1781, 160.1782, 160.1782, 160.1782, 
    160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 
    160.1782, 160.1782, 160.1782, 160.1782, 160.1783, 160.1783, 160.1783, 
    160.1783, 160.1783, 160.1783, 160.1783, 160.1783, 160.1783, 160.1783, 
    160.1783, 160.1783, 160.1783, 160.1783, 160.1783, 160.1783, 160.1782, 
    160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 
    160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1782, 160.1781, 
    160.1781, 160.1781, 160.1781, 160.1781, 160.1781, 160.1781, 160.1781, 
    160.1781, 160.1781, 160.178, 160.178, 160.178, 160.178, 160.178, 160.178, 
    160.178, 160.178, 160.1779, 160.1779, 160.1779, 160.1779, 160.1779, 
    160.1779, 160.1779, 160.1779,
  161.2033, 161.2033, 161.2033, 161.2033, 161.2033, 161.2033, 161.2033, 
    161.2033, 161.2033, 161.2033, 161.2034, 161.2034, 161.2034, 161.2034, 
    161.2034, 161.2034, 161.2034, 161.2034, 161.2034, 161.2034, 161.2035, 
    161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 
    161.2035, 161.2035, 161.2035, 161.2035, 161.2036, 161.2036, 161.2036, 
    161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 
    161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 
    161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 
    161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 161.2036, 
    161.2036, 161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 
    161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 161.2035, 161.2034, 
    161.2034, 161.2034, 161.2034, 161.2034, 161.2034, 161.2034, 161.2034, 
    161.2034, 161.2034, 161.2033, 161.2033, 161.2033, 161.2033, 161.2033, 
    161.2033, 161.2033, 161.2033, 161.2033, 161.2033,
  162.2314, 162.2315, 162.2315, 162.2315, 162.2315, 162.2315, 162.2315, 
    162.2315, 162.2315, 162.2315, 162.2315, 162.2316, 162.2316, 162.2316, 
    162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 
    162.2316, 162.2316, 162.2316, 162.2317, 162.2317, 162.2317, 162.2317, 
    162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 
    162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2318, 162.2318, 
    162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 
    162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 162.2318, 
    162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 
    162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 162.2317, 
    162.2317, 162.2317, 162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 
    162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 162.2316, 
    162.2316, 162.2315, 162.2315, 162.2315, 162.2315, 162.2315, 162.2315, 
    162.2315, 162.2315, 162.2315, 162.2315, 162.2314,
  163.2621, 163.2621, 163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 
    163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 
    163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 
    163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 
    163.2623, 163.2623, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 
    163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 
    163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 
    163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 
    163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 163.2624, 
    163.2624, 163.2624, 163.2624, 163.2623, 163.2623, 163.2623, 163.2623, 
    163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 
    163.2623, 163.2623, 163.2623, 163.2623, 163.2623, 163.2622, 163.2622, 
    163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 163.2622, 
    163.2622, 163.2622, 163.2622, 163.2621, 163.2621,
  164.295, 164.295, 164.295, 164.295, 164.295, 164.295, 164.295, 164.2951, 
    164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 
    164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 164.2952, 
    164.2952, 164.2952, 164.2952, 164.2952, 164.2951, 164.2951, 164.2951, 
    164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 164.2951, 
    164.2951, 164.2951, 164.2951, 164.2951, 164.295, 164.295, 164.295, 
    164.295, 164.295, 164.295, 164.295,
  165.3297, 165.3297, 165.3297, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 165.3299, 
    165.3299, 165.3299, 165.3299, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 165.3298, 
    165.3298, 165.3298, 165.3297, 165.3297, 165.3297,
  166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 
    166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 166.3661, 
    166.3661, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 
    166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 166.366, 
    166.366,
  167.4034, 167.4034, 167.4034, 167.4034, 167.4034, 167.4034, 167.4034, 
    167.4034, 167.4034, 167.4034, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 167.4035, 
    167.4035, 167.4035, 167.4034, 167.4034, 167.4034, 167.4034, 167.4034, 
    167.4034, 167.4034, 167.4034, 167.4034, 167.4034,
  168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 
    168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 
    168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 
    168.4418, 168.4418, 168.4418, 168.4418, 168.4418, 168.4417, 168.4417, 
    168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 
    168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 168.4417, 
    168.4417, 168.4417, 168.4417, 168.4417, 168.4417,
  169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 169.4805, 
    169.4805, 169.4805, 169.4805, 169.4805, 169.4805,
  170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 170.5195, 
    170.5195, 170.5195, 170.5195, 170.5195, 170.5195,
  171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 
    171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 
    171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 
    171.5582, 171.5582, 171.5582, 171.5582, 171.5582, 171.5583, 171.5583, 
    171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 
    171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 171.5583, 
    171.5583, 171.5583, 171.5583, 171.5583, 171.5583,
  172.5966, 172.5966, 172.5966, 172.5966, 172.5966, 172.5966, 172.5966, 
    172.5966, 172.5966, 172.5966, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 172.5965, 
    172.5965, 172.5965, 172.5966, 172.5966, 172.5966, 172.5966, 172.5966, 
    172.5966, 172.5966, 172.5966, 172.5966, 172.5966,
  173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 
    173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 173.6339, 
    173.6339, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 
    173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 173.634, 
    173.634,
  174.6703, 174.6703, 174.6703, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 174.6701, 
    174.6701, 174.6701, 174.6701, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 174.6702, 
    174.6702, 174.6702, 174.6703, 174.6703, 174.6703,
  175.705, 175.705, 175.705, 175.705, 175.705, 175.705, 175.705, 175.7049, 
    175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 
    175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 175.7048, 
    175.7048, 175.7048, 175.7048, 175.7048, 175.7049, 175.7049, 175.7049, 
    175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 175.7049, 
    175.7049, 175.7049, 175.7049, 175.7049, 175.705, 175.705, 175.705, 
    175.705, 175.705, 175.705, 175.705,
  176.7379, 176.7379, 176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 
    176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 
    176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 
    176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 
    176.7377, 176.7377, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 
    176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 
    176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 
    176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 
    176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 176.7376, 
    176.7376, 176.7376, 176.7376, 176.7377, 176.7377, 176.7377, 176.7377, 
    176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 
    176.7377, 176.7377, 176.7377, 176.7377, 176.7377, 176.7378, 176.7378, 
    176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 176.7378, 
    176.7378, 176.7378, 176.7378, 176.7379, 176.7379,
  177.7686, 177.7685, 177.7685, 177.7685, 177.7685, 177.7685, 177.7685, 
    177.7685, 177.7685, 177.7685, 177.7685, 177.7684, 177.7684, 177.7684, 
    177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 
    177.7684, 177.7684, 177.7684, 177.7683, 177.7683, 177.7683, 177.7683, 
    177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 
    177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7682, 177.7682, 
    177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 
    177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 177.7682, 
    177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 
    177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 177.7683, 
    177.7683, 177.7683, 177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 
    177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 177.7684, 
    177.7684, 177.7685, 177.7685, 177.7685, 177.7685, 177.7685, 177.7685, 
    177.7685, 177.7685, 177.7685, 177.7685, 177.7686,
  178.7967, 178.7967, 178.7967, 178.7967, 178.7967, 178.7967, 178.7967, 
    178.7967, 178.7967, 178.7967, 178.7966, 178.7966, 178.7966, 178.7966, 
    178.7966, 178.7966, 178.7966, 178.7966, 178.7966, 178.7966, 178.7965, 
    178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 
    178.7965, 178.7965, 178.7965, 178.7965, 178.7964, 178.7964, 178.7964, 
    178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 
    178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 
    178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 
    178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 178.7964, 
    178.7964, 178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 
    178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 178.7965, 178.7966, 
    178.7966, 178.7966, 178.7966, 178.7966, 178.7966, 178.7966, 178.7966, 
    178.7966, 178.7966, 178.7967, 178.7967, 178.7967, 178.7967, 178.7967, 
    178.7967, 178.7967, 178.7967, 178.7967, 178.7967,
  179.8221, 179.8221, 179.8221, 179.8221, 179.8221, 179.8221, 179.8221, 
    179.8221, 179.822, 179.822, 179.822, 179.822, 179.822, 179.822, 179.822, 
    179.822, 179.8219, 179.8219, 179.8219, 179.8219, 179.8219, 179.8219, 
    179.8219, 179.8219, 179.8219, 179.8219, 179.8218, 179.8218, 179.8218, 
    179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 
    179.8218, 179.8218, 179.8218, 179.8218, 179.8217, 179.8217, 179.8217, 
    179.8217, 179.8217, 179.8217, 179.8217, 179.8217, 179.8217, 179.8217, 
    179.8217, 179.8217, 179.8217, 179.8217, 179.8217, 179.8217, 179.8218, 
    179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 
    179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8218, 179.8219, 
    179.8219, 179.8219, 179.8219, 179.8219, 179.8219, 179.8219, 179.8219, 
    179.8219, 179.8219, 179.822, 179.822, 179.822, 179.822, 179.822, 179.822, 
    179.822, 179.822, 179.8221, 179.8221, 179.8221, 179.8221, 179.8221, 
    179.8221, 179.8221, 179.8221,
  180.8444, 180.8444, 180.8444, 180.8443, 180.8443, 180.8443, 180.8443, 
    180.8443, 180.8443, 180.8443, 180.8443, 180.8443, 180.8442, 180.8442, 
    180.8442, 180.8442, 180.8442, 180.8442, 180.8442, 180.8441, 180.8441, 
    180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 
    180.8441, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 
    180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 
    180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 
    180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 
    180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.844, 180.8441, 
    180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 180.8441, 
    180.8441, 180.8441, 180.8442, 180.8442, 180.8442, 180.8442, 180.8442, 
    180.8442, 180.8442, 180.8443, 180.8443, 180.8443, 180.8443, 180.8443, 
    180.8443, 180.8443, 180.8443, 180.8443, 180.8444, 180.8444, 180.8444,
  181.8632, 181.8632, 181.8632, 181.8632, 181.8632, 181.8632, 181.8631, 
    181.8631, 181.8631, 181.8631, 181.8631, 181.8631, 181.8631, 181.8631, 
    181.863, 181.863, 181.863, 181.863, 181.863, 181.863, 181.863, 181.8629, 
    181.8629, 181.8629, 181.8629, 181.8629, 181.8629, 181.8629, 181.8629, 
    181.8629, 181.8629, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 
    181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 
    181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 
    181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 
    181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 181.8628, 
    181.8628, 181.8629, 181.8629, 181.8629, 181.8629, 181.8629, 181.8629, 
    181.8629, 181.8629, 181.8629, 181.8629, 181.863, 181.863, 181.863, 
    181.863, 181.863, 181.863, 181.863, 181.8631, 181.8631, 181.8631, 
    181.8631, 181.8631, 181.8631, 181.8631, 181.8631, 181.8632, 181.8632, 
    181.8632, 181.8632, 181.8632, 181.8632,
  182.8783, 182.8783, 182.8783, 182.8783, 182.8783, 182.8783, 182.8783, 
    182.8783, 182.8782, 182.8782, 182.8782, 182.8782, 182.8782, 182.8782, 
    182.8781, 182.8781, 182.8781, 182.8781, 182.8781, 182.8781, 182.8781, 
    182.8781, 182.878, 182.878, 182.878, 182.878, 182.878, 182.878, 182.878, 
    182.878, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 
    182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 
    182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 
    182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 
    182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 182.8779, 
    182.8779, 182.8779, 182.878, 182.878, 182.878, 182.878, 182.878, 182.878, 
    182.878, 182.878, 182.8781, 182.8781, 182.8781, 182.8781, 182.8781, 
    182.8781, 182.8781, 182.8781, 182.8782, 182.8782, 182.8782, 182.8782, 
    182.8782, 182.8782, 182.8783, 182.8783, 182.8783, 182.8783, 182.8783, 
    182.8783, 182.8783, 182.8783,
  183.8895, 183.8895, 183.8895, 183.8894, 183.8894, 183.8894, 183.8894, 
    183.8894, 183.8894, 183.8893, 183.8893, 183.8893, 183.8893, 183.8893, 
    183.8893, 183.8893, 183.8892, 183.8892, 183.8892, 183.8892, 183.8892, 
    183.8892, 183.8892, 183.8891, 183.8891, 183.8891, 183.8891, 183.8891, 
    183.8891, 183.8891, 183.8891, 183.8891, 183.889, 183.889, 183.889, 
    183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 
    183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 
    183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 183.889, 
    183.889, 183.889, 183.889, 183.889, 183.889, 183.8891, 183.8891, 
    183.8891, 183.8891, 183.8891, 183.8891, 183.8891, 183.8891, 183.8891, 
    183.8892, 183.8892, 183.8892, 183.8892, 183.8892, 183.8892, 183.8892, 
    183.8893, 183.8893, 183.8893, 183.8893, 183.8893, 183.8893, 183.8893, 
    183.8894, 183.8894, 183.8894, 183.8894, 183.8894, 183.8894, 183.8895, 
    183.8895, 183.8895,
  184.8964, 184.8963, 184.8963, 184.8963, 184.8963, 184.8963, 184.8963, 
    184.8963, 184.8962, 184.8962, 184.8962, 184.8962, 184.8962, 184.8961, 
    184.8961, 184.8961, 184.8961, 184.8961, 184.8961, 184.8961, 184.896, 
    184.896, 184.896, 184.896, 184.896, 184.896, 184.896, 184.896, 184.8959, 
    184.8959, 184.8959, 184.8959, 184.8959, 184.8959, 184.8959, 184.8959, 
    184.8959, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 
    184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 
    184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 184.8958, 
    184.8958, 184.8958, 184.8959, 184.8959, 184.8959, 184.8959, 184.8959, 
    184.8959, 184.8959, 184.8959, 184.8959, 184.896, 184.896, 184.896, 
    184.896, 184.896, 184.896, 184.896, 184.896, 184.8961, 184.8961, 
    184.8961, 184.8961, 184.8961, 184.8961, 184.8961, 184.8962, 184.8962, 
    184.8962, 184.8962, 184.8962, 184.8963, 184.8963, 184.8963, 184.8963, 
    184.8963, 184.8963, 184.8963, 184.8964,
  185.8987, 185.8987, 185.8987, 185.8987, 185.8987, 185.8986, 185.8986, 
    185.8986, 185.8986, 185.8986, 185.8985, 185.8985, 185.8985, 185.8985, 
    185.8985, 185.8985, 185.8984, 185.8984, 185.8984, 185.8984, 185.8984, 
    185.8984, 185.8983, 185.8983, 185.8983, 185.8983, 185.8983, 185.8983, 
    185.8983, 185.8982, 185.8982, 185.8982, 185.8982, 185.8982, 185.8982, 
    185.8982, 185.8982, 185.8982, 185.8982, 185.8981, 185.8981, 185.8981, 
    185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 
    185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 185.8981, 
    185.8981, 185.8982, 185.8982, 185.8982, 185.8982, 185.8982, 185.8982, 
    185.8982, 185.8982, 185.8982, 185.8982, 185.8983, 185.8983, 185.8983, 
    185.8983, 185.8983, 185.8983, 185.8983, 185.8984, 185.8984, 185.8984, 
    185.8984, 185.8984, 185.8984, 185.8985, 185.8985, 185.8985, 185.8985, 
    185.8985, 185.8985, 185.8986, 185.8986, 185.8986, 185.8986, 185.8986, 
    185.8987, 185.8987, 185.8987, 185.8987, 185.8987,
  186.8963, 186.8963, 186.8963, 186.8962, 186.8962, 186.8962, 186.8962, 
    186.8962, 186.8961, 186.8961, 186.8961, 186.8961, 186.8961, 186.8961, 
    186.896, 186.896, 186.896, 186.896, 186.896, 186.896, 186.8959, 186.8959, 
    186.8959, 186.8959, 186.8959, 186.8958, 186.8958, 186.8958, 186.8958, 
    186.8958, 186.8958, 186.8958, 186.8958, 186.8958, 186.8957, 186.8957, 
    186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 
    186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 
    186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 
    186.8957, 186.8957, 186.8957, 186.8957, 186.8957, 186.8958, 186.8958, 
    186.8958, 186.8958, 186.8958, 186.8958, 186.8958, 186.8958, 186.8958, 
    186.8959, 186.8959, 186.8959, 186.8959, 186.8959, 186.896, 186.896, 
    186.896, 186.896, 186.896, 186.896, 186.8961, 186.8961, 186.8961, 
    186.8961, 186.8961, 186.8961, 186.8962, 186.8962, 186.8962, 186.8962, 
    186.8962, 186.8963, 186.8963, 186.8963,
  187.8888, 187.8888, 187.8888, 187.8888, 187.8888, 187.8887, 187.8887, 
    187.8887, 187.8887, 187.8887, 187.8887, 187.8886, 187.8886, 187.8886, 
    187.8886, 187.8885, 187.8885, 187.8885, 187.8885, 187.8885, 187.8885, 
    187.8884, 187.8884, 187.8884, 187.8884, 187.8884, 187.8884, 187.8884, 
    187.8883, 187.8883, 187.8883, 187.8883, 187.8883, 187.8883, 187.8883, 
    187.8883, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 
    187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 
    187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 187.8882, 
    187.8882, 187.8882, 187.8882, 187.8882, 187.8883, 187.8883, 187.8883, 
    187.8883, 187.8883, 187.8883, 187.8883, 187.8883, 187.8884, 187.8884, 
    187.8884, 187.8884, 187.8884, 187.8884, 187.8884, 187.8885, 187.8885, 
    187.8885, 187.8885, 187.8885, 187.8885, 187.8886, 187.8886, 187.8886, 
    187.8886, 187.8887, 187.8887, 187.8887, 187.8887, 187.8887, 187.8887, 
    187.8888, 187.8888, 187.8888, 187.8888, 187.8888,
  188.8761, 188.8761, 188.8761, 188.8761, 188.8761, 188.8761, 188.876, 
    188.876, 188.876, 188.876, 188.8759, 188.8759, 188.8759, 188.8759, 
    188.8759, 188.8759, 188.8758, 188.8758, 188.8758, 188.8758, 188.8758, 
    188.8757, 188.8757, 188.8757, 188.8757, 188.8757, 188.8757, 188.8756, 
    188.8756, 188.8756, 188.8756, 188.8756, 188.8756, 188.8756, 188.8755, 
    188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 
    188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 
    188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 
    188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8755, 188.8756, 
    188.8756, 188.8756, 188.8756, 188.8756, 188.8756, 188.8756, 188.8757, 
    188.8757, 188.8757, 188.8757, 188.8757, 188.8757, 188.8758, 188.8758, 
    188.8758, 188.8758, 188.8758, 188.8759, 188.8759, 188.8759, 188.8759, 
    188.8759, 188.8759, 188.876, 188.876, 188.876, 188.876, 188.8761, 
    188.8761, 188.8761, 188.8761, 188.8761, 188.8761,
  189.858, 189.858, 189.858, 189.8579, 189.8579, 189.8579, 189.8579, 
    189.8578, 189.8578, 189.8578, 189.8578, 189.8578, 189.8577, 189.8577, 
    189.8577, 189.8577, 189.8577, 189.8577, 189.8576, 189.8576, 189.8576, 
    189.8576, 189.8576, 189.8575, 189.8575, 189.8575, 189.8575, 189.8575, 
    189.8575, 189.8574, 189.8574, 189.8574, 189.8574, 189.8574, 189.8574, 
    189.8574, 189.8574, 189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 
    189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 
    189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 189.8573, 
    189.8573, 189.8573, 189.8573, 189.8574, 189.8574, 189.8574, 189.8574, 
    189.8574, 189.8574, 189.8574, 189.8574, 189.8575, 189.8575, 189.8575, 
    189.8575, 189.8575, 189.8575, 189.8576, 189.8576, 189.8576, 189.8576, 
    189.8576, 189.8577, 189.8577, 189.8577, 189.8577, 189.8577, 189.8577, 
    189.8578, 189.8578, 189.8578, 189.8578, 189.8578, 189.8579, 189.8579, 
    189.8579, 189.8579, 189.858, 189.858, 189.858,
  190.8342, 190.8342, 190.8341, 190.8341, 190.8341, 190.8341, 190.834, 
    190.834, 190.834, 190.834, 190.834, 190.8339, 190.8339, 190.8339, 
    190.8339, 190.8338, 190.8338, 190.8338, 190.8338, 190.8338, 190.8338, 
    190.8337, 190.8337, 190.8337, 190.8337, 190.8337, 190.8336, 190.8336, 
    190.8336, 190.8336, 190.8336, 190.8336, 190.8336, 190.8335, 190.8335, 
    190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 
    190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 
    190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 
    190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 190.8335, 
    190.8336, 190.8336, 190.8336, 190.8336, 190.8336, 190.8336, 190.8336, 
    190.8337, 190.8337, 190.8337, 190.8337, 190.8337, 190.8338, 190.8338, 
    190.8338, 190.8338, 190.8338, 190.8338, 190.8339, 190.8339, 190.8339, 
    190.8339, 190.834, 190.834, 190.834, 190.834, 190.834, 190.8341, 
    190.8341, 190.8341, 190.8341, 190.8342, 190.8342,
  191.8045, 191.8045, 191.8044, 191.8044, 191.8044, 191.8044, 191.8043, 
    191.8043, 191.8043, 191.8043, 191.8043, 191.8042, 191.8042, 191.8042, 
    191.8042, 191.8041, 191.8041, 191.8041, 191.8041, 191.8041, 191.804, 
    191.804, 191.804, 191.804, 191.804, 191.804, 191.8039, 191.8039, 
    191.8039, 191.8039, 191.8039, 191.8038, 191.8038, 191.8038, 191.8038, 
    191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 
    191.8037, 191.8037, 191.8037, 191.8037, 191.8037, 191.8037, 191.8037, 
    191.8037, 191.8037, 191.8037, 191.8037, 191.8037, 191.8038, 191.8038, 
    191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 191.8038, 
    191.8038, 191.8038, 191.8039, 191.8039, 191.8039, 191.8039, 191.8039, 
    191.804, 191.804, 191.804, 191.804, 191.804, 191.804, 191.8041, 191.8041, 
    191.8041, 191.8041, 191.8041, 191.8042, 191.8042, 191.8042, 191.8042, 
    191.8043, 191.8043, 191.8043, 191.8043, 191.8043, 191.8044, 191.8044, 
    191.8044, 191.8044, 191.8045, 191.8045,
  192.7687, 192.7687, 192.7687, 192.7687, 192.7686, 192.7686, 192.7686, 
    192.7686, 192.7686, 192.7685, 192.7685, 192.7685, 192.7685, 192.7684, 
    192.7684, 192.7684, 192.7684, 192.7684, 192.7683, 192.7683, 192.7683, 
    192.7683, 192.7682, 192.7682, 192.7682, 192.7682, 192.7682, 192.7682, 
    192.7681, 192.7681, 192.7681, 192.7681, 192.7681, 192.7681, 192.7681, 
    192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 
    192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 
    192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 192.768, 
    192.768, 192.768, 192.7681, 192.7681, 192.7681, 192.7681, 192.7681, 
    192.7681, 192.7681, 192.7682, 192.7682, 192.7682, 192.7682, 192.7682, 
    192.7682, 192.7683, 192.7683, 192.7683, 192.7683, 192.7684, 192.7684, 
    192.7684, 192.7684, 192.7684, 192.7685, 192.7685, 192.7685, 192.7685, 
    192.7686, 192.7686, 192.7686, 192.7686, 192.7686, 192.7687, 192.7687, 
    192.7687, 192.7687,
  193.7268, 193.7268, 193.7267, 193.7267, 193.7267, 193.7267, 193.7266, 
    193.7266, 193.7266, 193.7266, 193.7265, 193.7265, 193.7265, 193.7265, 
    193.7264, 193.7264, 193.7264, 193.7264, 193.7264, 193.7263, 193.7263, 
    193.7263, 193.7263, 193.7263, 193.7262, 193.7262, 193.7262, 193.7262, 
    193.7262, 193.7262, 193.7261, 193.7261, 193.7261, 193.7261, 193.7261, 
    193.7261, 193.7261, 193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 
    193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 
    193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 193.726, 
    193.7261, 193.7261, 193.7261, 193.7261, 193.7261, 193.7261, 193.7261, 
    193.7262, 193.7262, 193.7262, 193.7262, 193.7262, 193.7262, 193.7263, 
    193.7263, 193.7263, 193.7263, 193.7263, 193.7264, 193.7264, 193.7264, 
    193.7264, 193.7264, 193.7265, 193.7265, 193.7265, 193.7265, 193.7266, 
    193.7266, 193.7266, 193.7266, 193.7267, 193.7267, 193.7267, 193.7267, 
    193.7268, 193.7268,
  194.6784, 194.6784, 194.6784, 194.6784, 194.6783, 194.6783, 194.6783, 
    194.6783, 194.6783, 194.6782, 194.6782, 194.6782, 194.6781, 194.6781, 
    194.6781, 194.6781, 194.6781, 194.678, 194.678, 194.678, 194.678, 
    194.6779, 194.6779, 194.6779, 194.6779, 194.6779, 194.6778, 194.6778, 
    194.6778, 194.6778, 194.6778, 194.6778, 194.6777, 194.6777, 194.6777, 
    194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 
    194.6777, 194.6776, 194.6776, 194.6776, 194.6776, 194.6776, 194.6776, 
    194.6776, 194.6776, 194.6776, 194.6776, 194.6777, 194.6777, 194.6777, 
    194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 194.6777, 
    194.6777, 194.6778, 194.6778, 194.6778, 194.6778, 194.6778, 194.6778, 
    194.6779, 194.6779, 194.6779, 194.6779, 194.6779, 194.678, 194.678, 
    194.678, 194.678, 194.6781, 194.6781, 194.6781, 194.6781, 194.6781, 
    194.6782, 194.6782, 194.6782, 194.6783, 194.6783, 194.6783, 194.6783, 
    194.6783, 194.6784, 194.6784, 194.6784, 194.6784,
  195.6236, 195.6236, 195.6235, 195.6235, 195.6235, 195.6235, 195.6234, 
    195.6234, 195.6234, 195.6234, 195.6233, 195.6233, 195.6233, 195.6233, 
    195.6232, 195.6232, 195.6232, 195.6232, 195.6231, 195.6231, 195.6231, 
    195.6231, 195.623, 195.623, 195.623, 195.623, 195.623, 195.623, 195.6229, 
    195.6229, 195.6229, 195.6229, 195.6229, 195.6229, 195.6228, 195.6228, 
    195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 
    195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 
    195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 
    195.6228, 195.6228, 195.6228, 195.6228, 195.6228, 195.6229, 195.6229, 
    195.6229, 195.6229, 195.6229, 195.6229, 195.623, 195.623, 195.623, 
    195.623, 195.623, 195.623, 195.6231, 195.6231, 195.6231, 195.6231, 
    195.6232, 195.6232, 195.6232, 195.6232, 195.6233, 195.6233, 195.6233, 
    195.6233, 195.6234, 195.6234, 195.6234, 195.6234, 195.6235, 195.6235, 
    195.6235, 195.6235, 195.6236, 195.6236,
  196.5621, 196.562, 196.562, 196.562, 196.562, 196.5619, 196.5619, 196.5619, 
    196.5619, 196.5618, 196.5618, 196.5618, 196.5618, 196.5617, 196.5617, 
    196.5617, 196.5617, 196.5616, 196.5616, 196.5616, 196.5616, 196.5615, 
    196.5615, 196.5615, 196.5615, 196.5615, 196.5614, 196.5614, 196.5614, 
    196.5614, 196.5614, 196.5614, 196.5613, 196.5613, 196.5613, 196.5613, 
    196.5613, 196.5613, 196.5613, 196.5613, 196.5612, 196.5612, 196.5612, 
    196.5612, 196.5612, 196.5612, 196.5612, 196.5612, 196.5612, 196.5612, 
    196.5612, 196.5612, 196.5612, 196.5612, 196.5612, 196.5612, 196.5613, 
    196.5613, 196.5613, 196.5613, 196.5613, 196.5613, 196.5613, 196.5613, 
    196.5614, 196.5614, 196.5614, 196.5614, 196.5614, 196.5614, 196.5615, 
    196.5615, 196.5615, 196.5615, 196.5615, 196.5616, 196.5616, 196.5616, 
    196.5616, 196.5617, 196.5617, 196.5617, 196.5617, 196.5618, 196.5618, 
    196.5618, 196.5618, 196.5619, 196.5619, 196.5619, 196.5619, 196.562, 
    196.562, 196.562, 196.562, 196.5621,
  197.4938, 197.4937, 197.4937, 197.4937, 197.4937, 197.4936, 197.4936, 
    197.4936, 197.4935, 197.4935, 197.4935, 197.4935, 197.4935, 197.4934, 
    197.4934, 197.4934, 197.4933, 197.4933, 197.4933, 197.4933, 197.4933, 
    197.4932, 197.4932, 197.4932, 197.4932, 197.4931, 197.4931, 197.4931, 
    197.4931, 197.4931, 197.4931, 197.493, 197.493, 197.493, 197.493, 
    197.493, 197.493, 197.493, 197.493, 197.493, 197.4929, 197.4929, 
    197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 
    197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 197.4929, 
    197.493, 197.493, 197.493, 197.493, 197.493, 197.493, 197.493, 197.493, 
    197.493, 197.4931, 197.4931, 197.4931, 197.4931, 197.4931, 197.4931, 
    197.4932, 197.4932, 197.4932, 197.4932, 197.4933, 197.4933, 197.4933, 
    197.4933, 197.4933, 197.4934, 197.4934, 197.4934, 197.4935, 197.4935, 
    197.4935, 197.4935, 197.4935, 197.4936, 197.4936, 197.4936, 197.4937, 
    197.4937, 197.4937, 197.4937, 197.4938,
  198.4186, 198.4185, 198.4185, 198.4185, 198.4185, 198.4184, 198.4184, 
    198.4184, 198.4184, 198.4183, 198.4183, 198.4183, 198.4182, 198.4182, 
    198.4182, 198.4182, 198.4182, 198.4181, 198.4181, 198.4181, 198.4181, 
    198.418, 198.418, 198.418, 198.418, 198.418, 198.4179, 198.4179, 
    198.4179, 198.4179, 198.4179, 198.4178, 198.4178, 198.4178, 198.4178, 
    198.4178, 198.4178, 198.4178, 198.4178, 198.4177, 198.4177, 198.4177, 
    198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 
    198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 198.4177, 
    198.4177, 198.4178, 198.4178, 198.4178, 198.4178, 198.4178, 198.4178, 
    198.4178, 198.4178, 198.4179, 198.4179, 198.4179, 198.4179, 198.4179, 
    198.418, 198.418, 198.418, 198.418, 198.418, 198.4181, 198.4181, 
    198.4181, 198.4181, 198.4182, 198.4182, 198.4182, 198.4182, 198.4182, 
    198.4183, 198.4183, 198.4183, 198.4184, 198.4184, 198.4184, 198.4184, 
    198.4185, 198.4185, 198.4185, 198.4185, 198.4186,
  199.3364, 199.3363, 199.3363, 199.3363, 199.3363, 199.3362, 199.3362, 
    199.3362, 199.3362, 199.3361, 199.3361, 199.3361, 199.3361, 199.336, 
    199.336, 199.336, 199.336, 199.3359, 199.3359, 199.3359, 199.3359, 
    199.3358, 199.3358, 199.3358, 199.3358, 199.3358, 199.3357, 199.3357, 
    199.3357, 199.3357, 199.3357, 199.3356, 199.3356, 199.3356, 199.3356, 
    199.3356, 199.3356, 199.3356, 199.3356, 199.3356, 199.3355, 199.3355, 
    199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 
    199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 199.3355, 
    199.3356, 199.3356, 199.3356, 199.3356, 199.3356, 199.3356, 199.3356, 
    199.3356, 199.3356, 199.3357, 199.3357, 199.3357, 199.3357, 199.3357, 
    199.3358, 199.3358, 199.3358, 199.3358, 199.3358, 199.3359, 199.3359, 
    199.3359, 199.3359, 199.336, 199.336, 199.336, 199.336, 199.3361, 
    199.3361, 199.3361, 199.3361, 199.3362, 199.3362, 199.3362, 199.3362, 
    199.3363, 199.3363, 199.3363, 199.3363, 199.3364,
  200.2471, 200.2471, 200.2471, 200.247, 200.247, 200.247, 200.2469, 
    200.2469, 200.2469, 200.2469, 200.2468, 200.2468, 200.2468, 200.2468, 
    200.2467, 200.2467, 200.2467, 200.2467, 200.2466, 200.2466, 200.2466, 
    200.2466, 200.2466, 200.2465, 200.2465, 200.2465, 200.2465, 200.2464, 
    200.2464, 200.2464, 200.2464, 200.2464, 200.2464, 200.2463, 200.2463, 
    200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 
    200.2462, 200.2462, 200.2462, 200.2462, 200.2462, 200.2462, 200.2462, 
    200.2462, 200.2462, 200.2462, 200.2462, 200.2462, 200.2463, 200.2463, 
    200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 200.2463, 
    200.2464, 200.2464, 200.2464, 200.2464, 200.2464, 200.2464, 200.2465, 
    200.2465, 200.2465, 200.2465, 200.2466, 200.2466, 200.2466, 200.2466, 
    200.2466, 200.2467, 200.2467, 200.2467, 200.2467, 200.2468, 200.2468, 
    200.2468, 200.2468, 200.2469, 200.2469, 200.2469, 200.2469, 200.247, 
    200.247, 200.247, 200.2471, 200.2471, 200.2471,
  201.1507, 201.1507, 201.1506, 201.1506, 201.1506, 201.1506, 201.1505, 
    201.1505, 201.1505, 201.1504, 201.1504, 201.1504, 201.1504, 201.1503, 
    201.1503, 201.1503, 201.1503, 201.1502, 201.1502, 201.1502, 201.1502, 
    201.1501, 201.1501, 201.1501, 201.1501, 201.1501, 201.15, 201.15, 201.15, 
    201.15, 201.15, 201.1499, 201.1499, 201.1499, 201.1499, 201.1499, 
    201.1499, 201.1499, 201.1499, 201.1498, 201.1498, 201.1498, 201.1498, 
    201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 
    201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 201.1498, 
    201.1499, 201.1499, 201.1499, 201.1499, 201.1499, 201.1499, 201.1499, 
    201.1499, 201.15, 201.15, 201.15, 201.15, 201.15, 201.1501, 201.1501, 
    201.1501, 201.1501, 201.1501, 201.1502, 201.1502, 201.1502, 201.1502, 
    201.1503, 201.1503, 201.1503, 201.1503, 201.1504, 201.1504, 201.1504, 
    201.1504, 201.1505, 201.1505, 201.1505, 201.1506, 201.1506, 201.1506, 
    201.1506, 201.1507, 201.1507,
  202.047, 202.047, 202.047, 202.047, 202.0469, 202.0469, 202.0469, 202.0468, 
    202.0468, 202.0468, 202.0468, 202.0467, 202.0467, 202.0467, 202.0467, 
    202.0466, 202.0466, 202.0466, 202.0466, 202.0465, 202.0465, 202.0465, 
    202.0465, 202.0464, 202.0464, 202.0464, 202.0464, 202.0464, 202.0463, 
    202.0463, 202.0463, 202.0463, 202.0463, 202.0463, 202.0462, 202.0462, 
    202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 
    202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 
    202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 
    202.0462, 202.0462, 202.0462, 202.0462, 202.0462, 202.0463, 202.0463, 
    202.0463, 202.0463, 202.0463, 202.0463, 202.0464, 202.0464, 202.0464, 
    202.0464, 202.0464, 202.0465, 202.0465, 202.0465, 202.0465, 202.0466, 
    202.0466, 202.0466, 202.0466, 202.0467, 202.0467, 202.0467, 202.0467, 
    202.0468, 202.0468, 202.0468, 202.0468, 202.0469, 202.0469, 202.0469, 
    202.047, 202.047, 202.047, 202.047,
  202.9361, 202.9361, 202.9361, 202.936, 202.936, 202.936, 202.9359, 
    202.9359, 202.9359, 202.9359, 202.9358, 202.9358, 202.9358, 202.9358, 
    202.9357, 202.9357, 202.9357, 202.9357, 202.9356, 202.9356, 202.9356, 
    202.9355, 202.9355, 202.9355, 202.9355, 202.9355, 202.9354, 202.9354, 
    202.9354, 202.9354, 202.9354, 202.9354, 202.9353, 202.9353, 202.9353, 
    202.9353, 202.9353, 202.9353, 202.9353, 202.9353, 202.9353, 202.9352, 
    202.9352, 202.9352, 202.9352, 202.9352, 202.9352, 202.9352, 202.9352, 
    202.9352, 202.9352, 202.9352, 202.9352, 202.9352, 202.9352, 202.9353, 
    202.9353, 202.9353, 202.9353, 202.9353, 202.9353, 202.9353, 202.9353, 
    202.9353, 202.9354, 202.9354, 202.9354, 202.9354, 202.9354, 202.9354, 
    202.9355, 202.9355, 202.9355, 202.9355, 202.9355, 202.9356, 202.9356, 
    202.9356, 202.9357, 202.9357, 202.9357, 202.9357, 202.9358, 202.9358, 
    202.9358, 202.9358, 202.9359, 202.9359, 202.9359, 202.9359, 202.936, 
    202.936, 202.936, 202.9361, 202.9361, 202.9361,
  203.8179, 203.8178, 203.8178, 203.8178, 203.8177, 203.8177, 203.8177, 
    203.8177, 203.8176, 203.8176, 203.8176, 203.8176, 203.8175, 203.8175, 
    203.8175, 203.8174, 203.8174, 203.8174, 203.8174, 203.8173, 203.8173, 
    203.8173, 203.8173, 203.8172, 203.8172, 203.8172, 203.8172, 203.8172, 
    203.8172, 203.8171, 203.8171, 203.8171, 203.8171, 203.8171, 203.8171, 
    203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 
    203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 
    203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 203.817, 
    203.817, 203.817, 203.8171, 203.8171, 203.8171, 203.8171, 203.8171, 
    203.8171, 203.8172, 203.8172, 203.8172, 203.8172, 203.8172, 203.8172, 
    203.8173, 203.8173, 203.8173, 203.8173, 203.8174, 203.8174, 203.8174, 
    203.8174, 203.8175, 203.8175, 203.8175, 203.8176, 203.8176, 203.8176, 
    203.8176, 203.8177, 203.8177, 203.8177, 203.8177, 203.8178, 203.8178, 
    203.8178, 203.8179,
  204.6923, 204.6922, 204.6922, 204.6922, 204.6921, 204.6921, 204.6921, 
    204.692, 204.692, 204.692, 204.692, 204.6919, 204.6919, 204.6919, 
    204.6918, 204.6918, 204.6918, 204.6918, 204.6918, 204.6917, 204.6917, 
    204.6917, 204.6917, 204.6916, 204.6916, 204.6916, 204.6916, 204.6916, 
    204.6915, 204.6915, 204.6915, 204.6915, 204.6915, 204.6915, 204.6914, 
    204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 
    204.6914, 204.6914, 204.6914, 204.6913, 204.6913, 204.6913, 204.6913, 
    204.6913, 204.6913, 204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 
    204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 204.6914, 204.6915, 
    204.6915, 204.6915, 204.6915, 204.6915, 204.6915, 204.6916, 204.6916, 
    204.6916, 204.6916, 204.6916, 204.6917, 204.6917, 204.6917, 204.6917, 
    204.6918, 204.6918, 204.6918, 204.6918, 204.6918, 204.6919, 204.6919, 
    204.6919, 204.692, 204.692, 204.692, 204.692, 204.6921, 204.6921, 
    204.6921, 204.6922, 204.6922, 204.6922, 204.6923,
  205.5592, 205.5592, 205.5592, 205.5592, 205.5591, 205.5591, 205.5591, 
    205.5591, 205.559, 205.559, 205.559, 205.5589, 205.5589, 205.5589, 
    205.5589, 205.5588, 205.5588, 205.5588, 205.5587, 205.5587, 205.5587, 
    205.5587, 205.5587, 205.5586, 205.5586, 205.5586, 205.5586, 205.5585, 
    205.5585, 205.5585, 205.5585, 205.5585, 205.5585, 205.5584, 205.5584, 
    205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 
    205.5584, 205.5583, 205.5583, 205.5583, 205.5583, 205.5583, 205.5583, 
    205.5583, 205.5583, 205.5583, 205.5583, 205.5584, 205.5584, 205.5584, 
    205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 205.5584, 
    205.5585, 205.5585, 205.5585, 205.5585, 205.5585, 205.5585, 205.5586, 
    205.5586, 205.5586, 205.5586, 205.5587, 205.5587, 205.5587, 205.5587, 
    205.5587, 205.5588, 205.5588, 205.5588, 205.5589, 205.5589, 205.5589, 
    205.5589, 205.559, 205.559, 205.559, 205.5591, 205.5591, 205.5591, 
    205.5591, 205.5592, 205.5592, 205.5592, 205.5592,
  206.4188, 206.4188, 206.4188, 206.4187, 206.4187, 206.4187, 206.4187, 
    206.4186, 206.4186, 206.4186, 206.4185, 206.4185, 206.4185, 206.4185, 
    206.4184, 206.4184, 206.4184, 206.4184, 206.4183, 206.4183, 206.4183, 
    206.4183, 206.4182, 206.4182, 206.4182, 206.4182, 206.4182, 206.4181, 
    206.4181, 206.4181, 206.4181, 206.4181, 206.418, 206.418, 206.418, 
    206.418, 206.418, 206.418, 206.418, 206.418, 206.418, 206.418, 206.418, 
    206.4179, 206.4179, 206.4179, 206.4179, 206.4179, 206.4179, 206.4179, 
    206.4179, 206.4179, 206.4179, 206.418, 206.418, 206.418, 206.418, 
    206.418, 206.418, 206.418, 206.418, 206.418, 206.418, 206.418, 206.4181, 
    206.4181, 206.4181, 206.4181, 206.4181, 206.4182, 206.4182, 206.4182, 
    206.4182, 206.4182, 206.4183, 206.4183, 206.4183, 206.4183, 206.4184, 
    206.4184, 206.4184, 206.4184, 206.4185, 206.4185, 206.4185, 206.4185, 
    206.4186, 206.4186, 206.4186, 206.4187, 206.4187, 206.4187, 206.4187, 
    206.4188, 206.4188, 206.4188,
  207.271, 207.271, 207.271, 207.2709, 207.2709, 207.2709, 207.2708, 
    207.2708, 207.2708, 207.2708, 207.2707, 207.2707, 207.2707, 207.2706, 
    207.2706, 207.2706, 207.2706, 207.2705, 207.2705, 207.2705, 207.2705, 
    207.2704, 207.2704, 207.2704, 207.2704, 207.2704, 207.2703, 207.2703, 
    207.2703, 207.2703, 207.2703, 207.2702, 207.2702, 207.2702, 207.2702, 
    207.2702, 207.2702, 207.2702, 207.2702, 207.2701, 207.2701, 207.2701, 
    207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 
    207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 207.2701, 
    207.2701, 207.2702, 207.2702, 207.2702, 207.2702, 207.2702, 207.2702, 
    207.2702, 207.2702, 207.2703, 207.2703, 207.2703, 207.2703, 207.2703, 
    207.2704, 207.2704, 207.2704, 207.2704, 207.2704, 207.2705, 207.2705, 
    207.2705, 207.2705, 207.2706, 207.2706, 207.2706, 207.2706, 207.2707, 
    207.2707, 207.2707, 207.2708, 207.2708, 207.2708, 207.2708, 207.2709, 
    207.2709, 207.2709, 207.271, 207.271, 207.271,
  208.1158, 208.1158, 208.1157, 208.1157, 208.1157, 208.1156, 208.1156, 
    208.1156, 208.1155, 208.1155, 208.1155, 208.1155, 208.1154, 208.1154, 
    208.1154, 208.1154, 208.1153, 208.1153, 208.1153, 208.1152, 208.1152, 
    208.1152, 208.1152, 208.1152, 208.1151, 208.1151, 208.1151, 208.1151, 
    208.1151, 208.115, 208.115, 208.115, 208.115, 208.115, 208.115, 208.115, 
    208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 
    208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 
    208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 208.1149, 
    208.1149, 208.1149, 208.1149, 208.115, 208.115, 208.115, 208.115, 
    208.115, 208.115, 208.115, 208.1151, 208.1151, 208.1151, 208.1151, 
    208.1151, 208.1152, 208.1152, 208.1152, 208.1152, 208.1152, 208.1153, 
    208.1153, 208.1153, 208.1154, 208.1154, 208.1154, 208.1154, 208.1155, 
    208.1155, 208.1155, 208.1155, 208.1156, 208.1156, 208.1156, 208.1157, 
    208.1157, 208.1157, 208.1158, 208.1158,
  208.9531, 208.9531, 208.9531, 208.953, 208.953, 208.953, 208.953, 208.9529, 
    208.9529, 208.9529, 208.9529, 208.9528, 208.9528, 208.9528, 208.9527, 
    208.9527, 208.9527, 208.9527, 208.9526, 208.9526, 208.9526, 208.9526, 
    208.9525, 208.9525, 208.9525, 208.9525, 208.9525, 208.9524, 208.9524, 
    208.9524, 208.9524, 208.9524, 208.9523, 208.9523, 208.9523, 208.9523, 
    208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 
    208.9523, 208.9522, 208.9522, 208.9522, 208.9522, 208.9522, 208.9522, 
    208.9522, 208.9522, 208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 
    208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 208.9523, 
    208.9524, 208.9524, 208.9524, 208.9524, 208.9524, 208.9525, 208.9525, 
    208.9525, 208.9525, 208.9525, 208.9526, 208.9526, 208.9526, 208.9526, 
    208.9527, 208.9527, 208.9527, 208.9527, 208.9528, 208.9528, 208.9528, 
    208.9529, 208.9529, 208.9529, 208.9529, 208.953, 208.953, 208.953, 
    208.953, 208.9531, 208.9531, 208.9531,
  209.7831, 209.7831, 209.7831, 209.783, 209.783, 209.783, 209.7829, 
    209.7829, 209.7829, 209.7828, 209.7828, 209.7828, 209.7828, 209.7827, 
    209.7827, 209.7827, 209.7827, 209.7826, 209.7826, 209.7826, 209.7825, 
    209.7825, 209.7825, 209.7825, 209.7825, 209.7824, 209.7824, 209.7824, 
    209.7824, 209.7824, 209.7823, 209.7823, 209.7823, 209.7823, 209.7823, 
    209.7823, 209.7823, 209.7823, 209.7823, 209.7822, 209.7822, 209.7822, 
    209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 
    209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 209.7822, 
    209.7822, 209.7823, 209.7823, 209.7823, 209.7823, 209.7823, 209.7823, 
    209.7823, 209.7823, 209.7823, 209.7824, 209.7824, 209.7824, 209.7824, 
    209.7824, 209.7825, 209.7825, 209.7825, 209.7825, 209.7825, 209.7826, 
    209.7826, 209.7826, 209.7827, 209.7827, 209.7827, 209.7827, 209.7828, 
    209.7828, 209.7828, 209.7828, 209.7829, 209.7829, 209.7829, 209.783, 
    209.783, 209.783, 209.7831, 209.7831, 209.7831,
  210.6057, 210.6057, 210.6057, 210.6056, 210.6056, 210.6056, 210.6055, 
    210.6055, 210.6055, 210.6054, 210.6054, 210.6054, 210.6054, 210.6053, 
    210.6053, 210.6053, 210.6053, 210.6052, 210.6052, 210.6052, 210.6051, 
    210.6051, 210.6051, 210.6051, 210.6051, 210.605, 210.605, 210.605, 
    210.605, 210.605, 210.6049, 210.6049, 210.6049, 210.6049, 210.6049, 
    210.6049, 210.6049, 210.6049, 210.6049, 210.6048, 210.6048, 210.6048, 
    210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 
    210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 210.6048, 
    210.6048, 210.6049, 210.6049, 210.6049, 210.6049, 210.6049, 210.6049, 
    210.6049, 210.6049, 210.6049, 210.605, 210.605, 210.605, 210.605, 
    210.605, 210.6051, 210.6051, 210.6051, 210.6051, 210.6051, 210.6052, 
    210.6052, 210.6052, 210.6053, 210.6053, 210.6053, 210.6053, 210.6054, 
    210.6054, 210.6054, 210.6054, 210.6055, 210.6055, 210.6055, 210.6056, 
    210.6056, 210.6056, 210.6057, 210.6057, 210.6057,
  211.421, 211.4209, 211.4209, 211.4209, 211.4209, 211.4208, 211.4208, 
    211.4208, 211.4207, 211.4207, 211.4207, 211.4207, 211.4206, 211.4206, 
    211.4206, 211.4205, 211.4205, 211.4205, 211.4205, 211.4204, 211.4204, 
    211.4204, 211.4204, 211.4203, 211.4203, 211.4203, 211.4203, 211.4203, 
    211.4203, 211.4202, 211.4202, 211.4202, 211.4202, 211.4202, 211.4202, 
    211.4202, 211.4202, 211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 
    211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 
    211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 211.4201, 
    211.4201, 211.4201, 211.4201, 211.4202, 211.4202, 211.4202, 211.4202, 
    211.4202, 211.4202, 211.4202, 211.4202, 211.4203, 211.4203, 211.4203, 
    211.4203, 211.4203, 211.4203, 211.4204, 211.4204, 211.4204, 211.4204, 
    211.4205, 211.4205, 211.4205, 211.4205, 211.4206, 211.4206, 211.4206, 
    211.4207, 211.4207, 211.4207, 211.4207, 211.4208, 211.4208, 211.4208, 
    211.4209, 211.4209, 211.4209, 211.4209, 211.421,
  212.2289, 212.2289, 212.2289, 212.2289, 212.2288, 212.2288, 212.2288, 
    212.2287, 212.2287, 212.2287, 212.2286, 212.2286, 212.2286, 212.2286, 
    212.2285, 212.2285, 212.2285, 212.2285, 212.2284, 212.2284, 212.2284, 
    212.2284, 212.2283, 212.2283, 212.2283, 212.2283, 212.2283, 212.2282, 
    212.2282, 212.2282, 212.2282, 212.2282, 212.2282, 212.2281, 212.2281, 
    212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 
    212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.228, 212.228, 
    212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 
    212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 212.2281, 
    212.2282, 212.2282, 212.2282, 212.2282, 212.2282, 212.2282, 212.2283, 
    212.2283, 212.2283, 212.2283, 212.2283, 212.2284, 212.2284, 212.2284, 
    212.2284, 212.2285, 212.2285, 212.2285, 212.2285, 212.2286, 212.2286, 
    212.2286, 212.2286, 212.2287, 212.2287, 212.2287, 212.2288, 212.2288, 
    212.2288, 212.2289, 212.2289, 212.2289, 212.2289,
  213.0296, 213.0296, 213.0296, 213.0296, 213.0295, 213.0295, 213.0295, 
    213.0294, 213.0294, 213.0294, 213.0293, 213.0293, 213.0293, 213.0293, 
    213.0292, 213.0292, 213.0292, 213.0292, 213.0291, 213.0291, 213.0291, 
    213.0291, 213.029, 213.029, 213.029, 213.029, 213.029, 213.0289, 
    213.0289, 213.0289, 213.0289, 213.0289, 213.0289, 213.0289, 213.0288, 
    213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 
    213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 
    213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 
    213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0288, 213.0289, 
    213.0289, 213.0289, 213.0289, 213.0289, 213.0289, 213.0289, 213.029, 
    213.029, 213.029, 213.029, 213.029, 213.0291, 213.0291, 213.0291, 
    213.0291, 213.0292, 213.0292, 213.0292, 213.0292, 213.0293, 213.0293, 
    213.0293, 213.0293, 213.0294, 213.0294, 213.0294, 213.0295, 213.0295, 
    213.0295, 213.0296, 213.0296, 213.0296, 213.0296,
  213.8231, 213.8231, 213.8231, 213.823, 213.823, 213.823, 213.823, 213.8229, 
    213.8229, 213.8229, 213.8228, 213.8228, 213.8228, 213.8228, 213.8227, 
    213.8227, 213.8227, 213.8226, 213.8226, 213.8226, 213.8226, 213.8226, 
    213.8225, 213.8225, 213.8225, 213.8225, 213.8225, 213.8224, 213.8224, 
    213.8224, 213.8224, 213.8224, 213.8224, 213.8224, 213.8223, 213.8223, 
    213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 
    213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 
    213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 
    213.8223, 213.8223, 213.8223, 213.8223, 213.8223, 213.8224, 213.8224, 
    213.8224, 213.8224, 213.8224, 213.8224, 213.8224, 213.8225, 213.8225, 
    213.8225, 213.8225, 213.8225, 213.8226, 213.8226, 213.8226, 213.8226, 
    213.8226, 213.8227, 213.8227, 213.8227, 213.8228, 213.8228, 213.8228, 
    213.8228, 213.8229, 213.8229, 213.8229, 213.823, 213.823, 213.823, 
    213.823, 213.8231, 213.8231, 213.8231,
  214.6095, 214.6095, 214.6094, 214.6094, 214.6094, 214.6093, 214.6093, 
    214.6093, 214.6092, 214.6092, 214.6092, 214.6091, 214.6091, 214.6091, 
    214.6091, 214.609, 214.609, 214.609, 214.609, 214.6089, 214.6089, 
    214.6089, 214.6089, 214.6089, 214.6088, 214.6088, 214.6088, 214.6088, 
    214.6088, 214.6087, 214.6087, 214.6087, 214.6087, 214.6087, 214.6087, 
    214.6087, 214.6087, 214.6087, 214.6086, 214.6086, 214.6086, 214.6086, 
    214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 
    214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 214.6086, 
    214.6086, 214.6086, 214.6087, 214.6087, 214.6087, 214.6087, 214.6087, 
    214.6087, 214.6087, 214.6087, 214.6087, 214.6088, 214.6088, 214.6088, 
    214.6088, 214.6088, 214.6089, 214.6089, 214.6089, 214.6089, 214.6089, 
    214.609, 214.609, 214.609, 214.609, 214.6091, 214.6091, 214.6091, 
    214.6091, 214.6092, 214.6092, 214.6092, 214.6093, 214.6093, 214.6093, 
    214.6094, 214.6094, 214.6094, 214.6095, 214.6095 ;

 grid_latt =
  35.07925, 34.34282, 33.60628, 32.86962, 32.13284, 31.39594, 30.65893, 
    29.92181, 29.18457, 28.44723, 27.70978, 26.97222, 26.23456, 25.4968, 
    24.75893, 24.02097, 23.28291, 22.54476, 21.80651, 21.06818, 20.32976, 
    19.59126, 18.85267, 18.114, 17.37526, 16.63645, 15.89756, 15.15861, 
    14.41959, 13.6805, 12.94136, 12.20216, 11.46291, 10.72361, 9.984256, 
    9.244861, 8.505425, 7.765951, 7.026442, 6.286901, 5.547333, 4.807739, 
    4.068124, 3.32849, 2.588841, 1.849181, 1.109512, 0.3698378, -0.3698378, 
    -1.109512, -1.849181, -2.588841, -3.32849, -4.068124, -4.807739, 
    -5.547333, -6.286901, -7.026442, -7.765951, -8.505425, -9.244861, 
    -9.984256, -10.72361, -11.46291, -12.20216, -12.94136, -13.6805, 
    -14.41959, -15.15861, -15.89756, -16.63645, -17.37526, -18.114, 
    -18.85267, -19.59126, -20.32976, -21.06818, -21.80651, -22.54476, 
    -23.28291, -24.02097, -24.75893, -25.4968, -26.23456, -26.97222, 
    -27.70978, -28.44723, -29.18457, -29.92181, -30.65893, -31.39594, 
    -32.13284, -32.86962, -33.60628, -34.34282, -35.07925,
  35.43988, 34.70005, 33.95987, 33.21932, 32.47842, 31.73718, 30.9956, 
    30.25368, 29.51142, 28.76883, 28.02592, 27.28269, 26.53915, 25.7953, 
    25.05115, 24.3067, 23.56197, 22.81695, 22.07165, 21.32609, 20.58027, 
    19.83419, 19.08786, 18.3413, 17.59451, 16.84749, 16.10026, 15.35282, 
    14.60518, 13.85736, 13.10935, 12.36118, 11.61284, 10.86435, 10.11571, 
    9.366945, 8.618052, 7.869044, 7.119931, 6.370722, 5.621428, 4.872057, 
    4.122622, 3.37313, 2.623593, 1.87402, 1.124422, 0.3748092, -0.3748092, 
    -1.124422, -1.87402, -2.623593, -3.37313, -4.122622, -4.872057, 
    -5.621428, -6.370722, -7.119931, -7.869044, -8.618052, -9.366945, 
    -10.11571, -10.86435, -11.61284, -12.36118, -13.10935, -13.85736, 
    -14.60518, -15.35282, -16.10026, -16.84749, -17.59451, -18.3413, 
    -19.08786, -19.83419, -20.58027, -21.32609, -22.07165, -22.81695, 
    -23.56197, -24.3067, -25.05115, -25.7953, -26.53915, -27.28269, 
    -28.02592, -28.76883, -29.51142, -30.25368, -30.9956, -31.73718, 
    -32.47842, -33.21932, -33.95987, -34.70005, -35.43988,
  35.79544, 35.05236, 34.30869, 33.56442, 32.81957, 32.07414, 31.32814, 
    30.58158, 29.83445, 29.08677, 28.33856, 27.58981, 26.84053, 26.09074, 
    25.34044, 24.58965, 23.83837, 23.08662, 22.33441, 21.58174, 20.82863, 
    20.0751, 19.32115, 18.5668, 17.81206, 17.05695, 16.30147, 15.54564, 
    14.78949, 14.03301, 13.27623, 12.51916, 11.76182, 11.00421, 10.24637, 
    9.488298, 8.730017, 7.971541, 7.212887, 6.454072, 5.695111, 4.936023, 
    4.176824, 3.41753, 2.658159, 1.898728, 1.139254, 0.3797542, -0.3797542, 
    -1.139254, -1.898728, -2.658159, -3.41753, -4.176824, -4.936023, 
    -5.695111, -6.454072, -7.212887, -7.971541, -8.730017, -9.488298, 
    -10.24637, -11.00421, -11.76182, -12.51916, -13.27623, -14.03301, 
    -14.78949, -15.54564, -16.30147, -17.05695, -17.81206, -18.5668, 
    -19.32115, -20.0751, -20.82863, -21.58174, -22.33441, -23.08662, 
    -23.83837, -24.58965, -25.34044, -26.09074, -26.84053, -27.58981, 
    -28.33856, -29.08677, -29.83445, -30.58158, -31.32814, -32.07414, 
    -32.81957, -33.56442, -34.30869, -35.05236, -35.79544,
  36.14578, 35.39962, 34.65261, 33.90479, 33.15614, 32.40669, 31.65643, 
    30.90537, 30.15354, 29.40093, 28.64755, 27.89343, 27.13857, 26.38298, 
    25.62668, 24.86968, 24.112, 23.35365, 22.59464, 21.835, 21.07474, 
    20.31387, 19.55242, 18.79039, 18.02782, 17.26471, 16.50109, 15.73699, 
    14.9724, 14.20737, 13.4419, 12.67602, 11.90976, 11.14313, 10.37615, 
    9.608856, 8.84126, 8.073387, 7.305261, 6.536906, 5.768345, 4.999602, 
    4.230701, 3.461666, 2.692521, 1.92329, 1.153999, 0.3846703, -0.3846703, 
    -1.153999, -1.92329, -2.692521, -3.461666, -4.230701, -4.999602, 
    -5.768345, -6.536906, -7.305261, -8.073387, -8.84126, -9.608856, 
    -10.37615, -11.14313, -11.90976, -12.67602, -13.4419, -14.20737, 
    -14.9724, -15.73699, -16.50109, -17.26471, -18.02782, -18.79039, 
    -19.55242, -20.31387, -21.07474, -21.835, -22.59464, -23.35365, -24.112, 
    -24.86968, -25.62668, -26.38298, -27.13857, -27.89343, -28.64755, 
    -29.40093, -30.15354, -30.90537, -31.65643, -32.40669, -33.15614, 
    -33.90479, -34.65261, -35.39962, -36.14578,
  36.4908, 35.7417, 34.99154, 34.2403, 33.48802, 32.73469, 31.98032, 
    31.22494, 30.46854, 29.71115, 28.95277, 28.19342, 27.43312, 26.67189, 
    25.90973, 25.14667, 24.38272, 23.6179, 22.85224, 22.08575, 21.31846, 
    20.55038, 19.78154, 19.01196, 18.24167, 17.47068, 16.69903, 15.92674, 
    15.15383, 14.38034, 13.60628, 12.83169, 12.05659, 11.28102, 10.505, 
    9.728554, 8.951721, 8.174527, 7.397004, 6.619181, 5.84109, 5.06276, 
    4.284225, 3.505514, 2.72666, 1.947694, 1.168648, 0.3895547, -0.3895547, 
    -1.168648, -1.947694, -2.72666, -3.505514, -4.284225, -5.06276, -5.84109, 
    -6.619181, -7.397004, -8.174527, -8.951721, -9.728554, -10.505, 
    -11.28102, -12.05659, -12.83169, -13.60628, -14.38034, -15.15383, 
    -15.92674, -16.69903, -17.47068, -18.24167, -19.01196, -19.78154, 
    -20.55038, -21.31846, -22.08575, -22.85224, -23.6179, -24.38272, 
    -25.14667, -25.90973, -26.67189, -27.43312, -28.19342, -28.95277, 
    -29.71115, -30.46854, -31.22494, -31.98032, -32.73469, -33.48802, 
    -34.2403, -34.99154, -35.7417, -36.4908,
  36.83038, 36.0785, 35.32531, 34.57083, 33.81506, 33.05801, 32.29969, 
    31.54013, 30.77932, 30.0173, 29.25407, 28.48965, 27.72406, 26.95732, 
    26.18944, 25.42046, 24.65038, 23.87924, 23.10706, 22.33386, 21.55966, 
    20.7845, 20.0084, 19.23139, 18.45349, 17.67474, 16.89517, 16.11481, 
    15.33368, 14.55183, 13.76928, 12.98607, 12.20224, 11.41781, 10.63283, 
    9.847324, 9.061338, 8.274905, 7.488063, 6.70085, 5.913303, 5.125462, 
    4.337364, 3.549049, 2.760556, 1.971925, 1.183195, 0.3944048, -0.3944048, 
    -1.183195, -1.971925, -2.760556, -3.549049, -4.337364, -5.125462, 
    -5.913303, -6.70085, -7.488063, -8.274905, -9.061338, -9.847324, 
    -10.63283, -11.41781, -12.20224, -12.98607, -13.76928, -14.55183, 
    -15.33368, -16.11481, -16.89517, -17.67474, -18.45349, -19.23139, 
    -20.0084, -20.7845, -21.55966, -22.33386, -23.10706, -23.87924, 
    -24.65038, -25.42046, -26.18944, -26.95732, -27.72406, -28.48965, 
    -29.25407, -30.0173, -30.77932, -31.54013, -32.29969, -33.05801, 
    -33.81506, -34.57083, -35.32531, -36.0785, -36.83038,
  37.1644, 36.40988, 35.65382, 34.89624, 34.13713, 33.37651, 32.6144, 
    31.8508, 31.08575, 30.31924, 29.55131, 28.78197, 28.01123, 27.23913, 
    26.46569, 25.69092, 24.91487, 24.13754, 23.35897, 22.57919, 21.79822, 
    21.01611, 20.23287, 19.44855, 18.66317, 17.87678, 17.0894, 16.30107, 
    15.51184, 14.72173, 13.9308, 13.13908, 12.3466, 11.55342, 10.75957, 
    9.965097, 9.170046, 8.37446, 7.578384, 6.781863, 5.984942, 5.187668, 
    4.390087, 3.592245, 2.79419, 1.995969, 1.197629, 0.3992176, -0.3992176, 
    -1.197629, -1.995969, -2.79419, -3.592245, -4.390087, -5.187668, 
    -5.984942, -6.781863, -7.578384, -8.37446, -9.170046, -9.965097, 
    -10.75957, -11.55342, -12.3466, -13.13908, -13.9308, -14.72173, 
    -15.51184, -16.30107, -17.0894, -17.87678, -18.66317, -19.44855, 
    -20.23287, -21.01611, -21.79822, -22.57919, -23.35897, -24.13754, 
    -24.91487, -25.69092, -26.46569, -27.23913, -28.01123, -28.78197, 
    -29.55131, -30.31924, -31.08575, -31.8508, -32.6144, -33.37651, 
    -34.13713, -34.89624, -35.65382, -36.40988, -37.1644,
  37.49273, 36.73572, 35.97694, 35.2164, 34.4541, 33.69006, 32.9243, 
    32.15683, 31.38766, 30.61683, 29.84434, 29.07022, 28.29449, 27.51719, 
    26.73832, 25.95792, 25.17602, 24.39264, 23.60783, 22.8216, 22.034, 
    21.24507, 20.45482, 19.66332, 18.87058, 18.07666, 17.2816, 16.48543, 
    15.6882, 14.88996, 14.09074, 13.29061, 12.4896, 11.68776, 10.88514, 
    10.0818, 9.277779, 8.473132, 7.667912, 6.862171, 6.055964, 5.249342, 
    4.442361, 3.635076, 2.827541, 2.019811, 1.211942, 0.40399, -0.40399, 
    -1.211942, -2.019811, -2.827541, -3.635076, -4.442361, -5.249342, 
    -6.055964, -6.862171, -7.667912, -8.473132, -9.277779, -10.0818, 
    -10.88514, -11.68776, -12.4896, -13.29061, -14.09074, -14.88996, 
    -15.6882, -16.48543, -17.2816, -18.07666, -18.87058, -19.66332, 
    -20.45482, -21.24507, -22.034, -22.8216, -23.60783, -24.39264, -25.17602, 
    -25.95792, -26.73832, -27.51719, -28.29449, -29.07022, -29.84434, 
    -30.61683, -31.38766, -32.15683, -32.9243, -33.69006, -34.4541, -35.2164, 
    -35.97694, -36.73572, -37.49273,
  37.81525, 37.05589, 36.29453, 35.53117, 34.76583, 33.99852, 33.22925, 
    32.45805, 31.68493, 30.90992, 30.13302, 29.35428, 28.5737, 27.79133, 
    27.00718, 26.22129, 25.43369, 24.64441, 23.85349, 23.06096, 22.26687, 
    21.47124, 20.67413, 19.87557, 19.07561, 18.27429, 17.47165, 16.66776, 
    15.86266, 15.05639, 14.24901, 13.44058, 12.63114, 11.82075, 11.00947, 
    10.19736, 9.384465, 8.570855, 7.756588, 6.941722, 6.12632, 5.310442, 
    4.494153, 3.677513, 2.860586, 2.043435, 1.226125, 0.4087191, -0.4087191, 
    -1.226125, -2.043435, -2.860586, -3.677513, -4.494153, -5.310442, 
    -6.12632, -6.941722, -7.756588, -8.570855, -9.384465, -10.19736, 
    -11.00947, -11.82075, -12.63114, -13.44058, -14.24901, -15.05639, 
    -15.86266, -16.66776, -17.47165, -18.27429, -19.07561, -19.87557, 
    -20.67413, -21.47124, -22.26687, -23.06096, -23.85349, -24.64441, 
    -25.43369, -26.22129, -27.00718, -27.79133, -28.5737, -29.35428, 
    -30.13302, -30.90992, -31.68493, -32.45805, -33.22925, -33.99852, 
    -34.76583, -35.53117, -36.29453, -37.05589, -37.81525,
  38.13184, 37.37026, 36.60646, 35.84042, 35.07218, 34.30174, 33.52912, 
    32.75434, 31.97741, 31.19835, 30.4172, 29.63398, 28.84871, 28.06141, 
    27.27213, 26.4809, 25.68774, 24.89271, 24.09582, 23.29713, 22.49667, 
    21.6945, 20.89065, 20.08517, 19.2781, 18.46952, 17.65945, 16.84796, 
    16.0351, 15.22093, 14.4055, 13.58888, 12.77113, 11.9523, 11.13247, 
    10.31169, 9.490034, 8.667565, 7.844352, 7.020462, 6.195964, 5.370928, 
    4.545426, 3.719527, 2.893303, 2.066826, 1.240168, 0.4134014, -0.4134014, 
    -1.240168, -2.066826, -2.893303, -3.719527, -4.545426, -5.370928, 
    -6.195964, -7.020462, -7.844352, -8.667565, -9.490034, -10.31169, 
    -11.13247, -11.9523, -12.77113, -13.58888, -14.4055, -15.22093, -16.0351, 
    -16.84796, -17.65945, -18.46952, -19.2781, -20.08517, -20.89065, 
    -21.6945, -22.49667, -23.29713, -24.09582, -24.89271, -25.68774, 
    -26.4809, -27.27213, -28.06141, -28.84871, -29.63398, -30.4172, 
    -31.19835, -31.97741, -32.75434, -33.52912, -34.30174, -35.07218, 
    -35.84042, -36.60646, -37.37026, -38.13184,
  38.44237, 37.67871, 36.91259, 36.14403, 35.37302, 34.59959, 33.82376, 
    33.04553, 32.26494, 31.482, 30.69673, 29.90917, 29.11935, 28.32729, 
    27.53302, 26.73659, 25.93803, 25.13737, 24.33467, 23.52995, 22.72328, 
    21.91469, 21.10424, 20.29198, 19.47795, 18.66223, 17.84485, 17.02589, 
    16.20541, 15.38346, 14.56011, 13.73542, 12.90947, 12.08233, 11.25405, 
    10.42472, 9.594414, 8.763195, 7.931143, 7.098334, 6.264847, 5.430757, 
    4.596145, 3.761089, 2.925669, 2.089966, 1.254061, 0.4180338, -0.4180338, 
    -1.254061, -2.089966, -2.925669, -3.761089, -4.596145, -5.430757, 
    -6.264847, -7.098334, -7.931143, -8.763195, -9.594414, -10.42472, 
    -11.25405, -12.08233, -12.90947, -13.73542, -14.56011, -15.38346, 
    -16.20541, -17.02589, -17.84485, -18.66223, -19.47795, -20.29198, 
    -21.10424, -21.91469, -22.72328, -23.52995, -24.33467, -25.13737, 
    -25.93803, -26.73659, -27.53302, -28.32729, -29.11935, -29.90917, 
    -30.69673, -31.482, -32.26494, -33.04553, -33.82376, -34.59959, 
    -35.37302, -36.14403, -36.91259, -37.67871, -38.44237,
  38.74672, 37.9811, 37.21281, 36.44184, 35.66821, 34.89193, 34.11302, 
    33.33149, 32.54737, 31.76069, 30.97146, 30.17971, 29.38548, 28.5888, 
    27.78969, 26.98821, 26.18438, 25.37826, 24.56988, 23.75929, 22.94654, 
    22.13168, 21.31477, 20.49586, 19.67501, 18.85229, 18.02774, 17.20144, 
    16.37346, 15.54386, 14.71272, 13.88009, 13.04607, 12.21073, 11.37413, 
    10.53637, 9.697527, 8.857674, 8.016898, 7.175284, 6.332918, 5.489884, 
    4.646272, 3.802168, 2.957661, 2.112839, 1.267794, 0.4226128, -0.4226128, 
    -1.267794, -2.112839, -2.957661, -3.802168, -4.646272, -5.489884, 
    -6.332918, -7.175284, -8.016898, -8.857674, -9.697527, -10.53637, 
    -11.37413, -12.21073, -13.04607, -13.88009, -14.71272, -15.54386, 
    -16.37346, -17.20144, -18.02774, -18.85229, -19.67501, -20.49586, 
    -21.31477, -22.13168, -22.94654, -23.75929, -24.56988, -25.37826, 
    -26.18438, -26.98821, -27.78969, -28.5888, -29.38548, -30.17971, 
    -30.97146, -31.76069, -32.54737, -33.33149, -34.11302, -34.89193, 
    -35.66821, -36.44184, -37.21281, -37.9811, -38.74672,
  39.04476, 38.27731, 37.50697, 36.73372, 35.9576, 35.1786, 34.39675, 
    33.61207, 32.82457, 32.03428, 31.24123, 30.44544, 29.64695, 28.84579, 
    28.04199, 27.2356, 26.42666, 25.61521, 24.8013, 23.98498, 23.1663, 
    22.34532, 21.52209, 20.69669, 19.86915, 19.03956, 18.20799, 17.37449, 
    16.53915, 15.70203, 14.86322, 14.02279, 13.18083, 12.33741, 11.49262, 
    10.64656, 9.799295, 8.95093, 8.101551, 7.251252, 6.400125, 5.548265, 
    4.695769, 3.842732, 2.989253, 2.135427, 1.281355, 0.4271349, -0.4271349, 
    -1.281355, -2.135427, -2.989253, -3.842732, -4.695769, -5.548265, 
    -6.400125, -7.251252, -8.101551, -8.95093, -9.799295, -10.64656, 
    -11.49262, -12.33741, -13.18083, -14.02279, -14.86322, -15.70203, 
    -16.53915, -17.37449, -18.20799, -19.03956, -19.86915, -20.69669, 
    -21.52209, -22.34532, -23.1663, -23.98498, -24.8013, -25.61521, 
    -26.42666, -27.2356, -28.04199, -28.84579, -29.64695, -30.44544, 
    -31.24123, -32.03428, -32.82457, -33.61207, -34.39675, -35.1786, 
    -35.9576, -36.73372, -37.50697, -38.27731, -39.04476,
  39.33637, 38.56721, 37.79493, 37.01954, 36.24105, 35.45947, 34.67482, 
    33.88711, 33.09637, 32.30262, 31.50589, 30.7062, 29.90359, 29.0981, 
    28.28975, 27.47861, 26.6647, 25.84807, 25.02878, 24.20688, 23.38242, 
    22.55546, 21.72607, 20.8943, 20.06023, 19.22392, 18.38545, 17.5449, 
    16.70233, 15.85784, 15.0115, 14.1634, 13.31363, 12.46228, 11.60943, 
    10.75519, 9.899641, 9.042892, 8.185037, 7.326178, 6.466415, 5.605854, 
    4.744597, 3.88275, 3.02042, 2.157712, 1.294735, 0.4315965, -0.4315965, 
    -1.294735, -2.157712, -3.02042, -3.88275, -4.744597, -5.605854, 
    -6.466415, -7.326178, -8.185037, -9.042892, -9.899641, -10.75519, 
    -11.60943, -12.46228, -13.31363, -14.1634, -15.0115, -15.85784, 
    -16.70233, -17.5449, -18.38545, -19.22392, -20.06023, -20.8943, 
    -21.72607, -22.55546, -23.38242, -24.20688, -25.02878, -25.84807, 
    -26.6647, -27.47861, -28.28975, -29.0981, -29.90359, -30.7062, -31.50589, 
    -32.30262, -33.09637, -33.88711, -34.67482, -35.45947, -36.24105, 
    -37.01954, -37.79493, -38.56721, -39.33637,
  39.62142, 38.85067, 38.07658, 37.29916, 36.51843, 35.73439, 34.94707, 
    34.15647, 33.36263, 32.56555, 31.76528, 30.96183, 30.15525, 29.34557, 
    28.53283, 27.71707, 26.89834, 26.07669, 25.25217, 24.42483, 23.59474, 
    22.76195, 21.92654, 21.08856, 20.2481, 19.40522, 18.56001, 17.71254, 
    16.8629, 16.01117, 15.15745, 14.30182, 13.44438, 12.58523, 11.72446, 
    10.86218, 9.998483, 9.133484, 8.267286, 7.4, 6.531734, 5.662601, 
    4.792715, 3.922188, 3.051136, 2.179676, 1.307923, 0.4359938, -0.4359938, 
    -1.307923, -2.179676, -3.051136, -3.922188, -4.792715, -5.662601, 
    -6.531734, -7.4, -8.267286, -9.133484, -9.998483, -10.86218, -11.72446, 
    -12.58523, -13.44438, -14.30182, -15.15745, -16.01117, -16.8629, 
    -17.71254, -18.56001, -19.40522, -20.2481, -21.08856, -21.92654, 
    -22.76195, -23.59474, -24.42483, -25.25217, -26.07669, -26.89834, 
    -27.71707, -28.53283, -29.34557, -30.15525, -30.96183, -31.76528, 
    -32.56555, -33.36263, -34.15647, -34.94707, -35.73439, -36.51843, 
    -37.29916, -38.07658, -38.85067, -39.62142,
  39.89979, 39.12755, 38.35176, 37.57244, 36.78959, 36.00322, 35.21335, 
    34.42, 33.62318, 32.82292, 32.01924, 31.21218, 30.40177, 29.58805, 
    28.77106, 27.95084, 27.12744, 26.30091, 25.4713, 24.63868, 23.8031, 
    22.96464, 22.12335, 21.27932, 20.43262, 19.58332, 18.73152, 17.87728, 
    17.02072, 16.1619, 15.30094, 14.43793, 13.57297, 12.70616, 11.83762, 
    10.96744, 10.09574, 9.222629, 8.34823, 7.472656, 6.596026, 5.718461, 
    4.840082, 3.961012, 3.081377, 2.201299, 1.320906, 0.4403231, -0.4403231, 
    -1.320906, -2.201299, -3.081377, -3.961012, -4.840082, -5.718461, 
    -6.596026, -7.472656, -8.34823, -9.222629, -10.09574, -10.96744, 
    -11.83762, -12.70616, -13.57297, -14.43793, -15.30094, -16.1619, 
    -17.02072, -17.87728, -18.73152, -19.58332, -20.43262, -21.27932, 
    -22.12335, -22.96464, -23.8031, -24.63868, -25.4713, -26.30091, 
    -27.12744, -27.95084, -28.77106, -29.58805, -30.40177, -31.21218, 
    -32.01924, -32.82292, -33.62318, -34.42, -35.21335, -36.00322, -36.78959, 
    -37.57244, -38.35176, -39.12755, -39.89979,
  40.17135, 39.39772, 38.62035, 37.83924, 37.05439, 36.26581, 35.47353, 
    34.67754, 33.87788, 33.07457, 32.26763, 31.45709, 30.643, 29.82537, 
    29.00427, 28.17974, 27.35181, 26.52055, 25.68602, 24.84826, 24.00736, 
    23.16337, 22.31637, 21.46644, 20.61365, 19.75808, 18.89984, 18.03899, 
    17.17565, 16.30991, 15.44186, 14.57162, 13.69929, 12.82498, 11.9488, 
    11.07087, 10.19132, 9.31025, 8.427797, 7.544083, 6.659235, 5.773382, 
    4.886656, 3.999188, 3.111113, 2.222563, 1.333673, 0.4445804, -0.4445804, 
    -1.333673, -2.222563, -3.111113, -3.999188, -4.886656, -5.773382, 
    -6.659235, -7.544083, -8.427797, -9.31025, -10.19132, -11.07087, 
    -11.9488, -12.82498, -13.69929, -14.57162, -15.44186, -16.30991, 
    -17.17565, -18.03899, -18.89984, -19.75808, -20.61365, -21.46644, 
    -22.31637, -23.16337, -24.00736, -24.84826, -25.68602, -26.52055, 
    -27.35181, -28.17974, -29.00427, -29.82537, -30.643, -31.45709, 
    -32.26763, -33.07457, -33.87788, -34.67754, -35.47353, -36.26581, 
    -37.05439, -37.83924, -38.62035, -39.39772, -40.17135,
  40.43598, 39.66107, 38.88222, 38.09942, 37.31269, 36.52202, 35.72744, 
    34.92895, 34.12658, 33.32034, 32.51027, 31.6964, 30.87876, 30.05738, 
    29.23232, 28.40361, 27.57131, 26.73548, 25.89616, 25.05343, 24.20735, 
    23.35799, 22.50543, 21.64975, 20.79103, 19.92936, 19.06483, 18.19754, 
    17.32758, 16.45506, 15.58009, 14.70277, 13.82323, 12.94157, 12.05792, 
    11.1724, 10.28514, 9.396269, 8.505915, 7.614214, 6.721301, 5.827315, 
    4.932395, 4.036681, 3.140318, 2.243447, 1.346213, 0.448762, -0.448762, 
    -1.346213, -2.243447, -3.140318, -4.036681, -4.932395, -5.827315, 
    -6.721301, -7.614214, -8.505915, -9.396269, -10.28514, -11.1724, 
    -12.05792, -12.94157, -13.82323, -14.70277, -15.58009, -16.45506, 
    -17.32758, -18.19754, -19.06483, -19.92936, -20.79103, -21.64975, 
    -22.50543, -23.35799, -24.20735, -25.05343, -25.89616, -26.73548, 
    -27.57131, -28.40361, -29.23232, -30.05738, -30.87876, -31.6964, 
    -32.51027, -33.32034, -34.12658, -34.92895, -35.72744, -36.52202, 
    -37.31269, -38.09942, -38.88222, -39.66107, -40.43598,
  40.69355, 39.91746, 39.13723, 38.35286, 37.56434, 36.7717, 35.97494, 
    35.17407, 34.36911, 33.56009, 32.74702, 31.92994, 31.10889, 30.28391, 
    29.45502, 28.6223, 27.78577, 26.94551, 26.10157, 25.25401, 24.40292, 
    23.54835, 22.69039, 21.82912, 20.96463, 20.09701, 19.22636, 18.35277, 
    17.47636, 16.59723, 15.71549, 14.83126, 13.94467, 13.05583, 12.16487, 
    11.27192, 10.37712, 9.480604, 8.582511, 7.682984, 6.782168, 5.880208, 
    4.977254, 4.073455, 3.168964, 2.263932, 1.358514, 0.4528638, -0.4528638, 
    -1.358514, -2.263932, -3.168964, -4.073455, -4.977254, -5.880208, 
    -6.782168, -7.682984, -8.582511, -9.480604, -10.37712, -11.27192, 
    -12.16487, -13.05583, -13.94467, -14.83126, -15.71549, -16.59723, 
    -17.47636, -18.35277, -19.22636, -20.09701, -20.96463, -21.82912, 
    -22.69039, -23.54835, -24.40292, -25.25401, -26.10157, -26.94551, 
    -27.78577, -28.6223, -29.45502, -30.28391, -31.10889, -31.92994, 
    -32.74702, -33.56009, -34.36911, -35.17407, -35.97494, -36.7717, 
    -37.56434, -38.35286, -39.13723, -39.91746, -40.69355,
  40.94394, 40.16676, 39.38524, 38.5994, 37.80922, 37.01471, 36.21589, 
    35.41275, 34.60533, 33.79364, 32.97771, 32.15757, 31.33325, 30.50479, 
    29.67224, 28.83563, 27.99503, 27.1505, 26.30208, 25.44986, 24.5939, 
    23.73428, 22.87107, 22.00438, 21.13428, 20.26088, 19.38427, 18.50457, 
    17.62187, 16.73629, 15.84795, 14.95698, 14.0635, 13.16765, 12.26954, 
    11.36934, 10.46716, 9.563174, 8.657512, 7.750327, 6.841775, 5.93201, 
    5.02119, 4.109474, 3.197022, 2.283998, 1.370563, 0.4568816, -0.4568816, 
    -1.370563, -2.283998, -3.197022, -4.109474, -5.02119, -5.93201, 
    -6.841775, -7.750327, -8.657512, -9.563174, -10.46716, -11.36934, 
    -12.26954, -13.16765, -14.0635, -14.95698, -15.84795, -16.73629, 
    -17.62187, -18.50457, -19.38427, -20.26088, -21.13428, -22.00438, 
    -22.87107, -23.73428, -24.5939, -25.44986, -26.30208, -27.1505, 
    -27.99503, -28.83563, -29.67224, -30.50479, -31.33325, -32.15757, 
    -32.97771, -33.79364, -34.60533, -35.41275, -36.21589, -37.01471, 
    -37.80922, -38.5994, -39.38524, -40.16676, -40.94394,
  41.18702, 40.40884, 39.62614, 38.83891, 38.04717, 37.2509, 36.45013, 
    35.64485, 34.83509, 34.02087, 33.2022, 32.37912, 31.55167, 30.71988, 
    29.88379, 29.04346, 28.19893, 27.35027, 26.49753, 25.6408, 24.78014, 
    23.91562, 23.04734, 22.17539, 21.29985, 20.42083, 19.53844, 18.65277, 
    17.76396, 16.87211, 15.97735, 15.07981, 14.17962, 13.27692, 12.37185, 
    11.46456, 10.55519, 9.643898, 8.730841, 7.816175, 6.900063, 5.982669, 
    5.064158, 4.144701, 3.224465, 2.303623, 1.382348, 0.4608116, -0.4608116, 
    -1.382348, -2.303623, -3.224465, -4.144701, -5.064158, -5.982669, 
    -6.900063, -7.816175, -8.730841, -9.643898, -10.55519, -11.46456, 
    -12.37185, -13.27692, -14.17962, -15.07981, -15.97735, -16.87211, 
    -17.76396, -18.65277, -19.53844, -20.42083, -21.29985, -22.17539, 
    -23.04734, -23.91562, -24.78014, -25.6408, -26.49753, -27.35027, 
    -28.19893, -29.04346, -29.88379, -30.71988, -31.55167, -32.37912, 
    -33.2022, -34.02087, -34.83509, -35.64485, -36.45013, -37.2509, 
    -38.04717, -38.83891, -39.62614, -40.40884, -41.18702,
  41.42268, 40.64358, 39.85978, 39.07127, 38.27806, 37.48015, 36.67753, 
    35.87022, 35.05824, 34.2416, 33.42032, 32.59444, 31.76398, 30.929, 
    30.08952, 29.2456, 28.3973, 27.54466, 26.68777, 25.82668, 24.96147, 
    24.09223, 23.21904, 22.34199, 21.46118, 20.57672, 19.68871, 18.79726, 
    17.9025, 17.00456, 16.10355, 15.19962, 14.2929, 13.38354, 12.47168, 
    11.55748, 10.6411, 9.722692, 8.802423, 7.880459, 6.956971, 6.032131, 
    5.106114, 4.179099, 3.251263, 2.322789, 1.393856, 0.4646493, -0.4646493, 
    -1.393856, -2.322789, -3.251263, -4.179099, -5.106114, -6.032131, 
    -6.956971, -7.880459, -8.802423, -9.722692, -10.6411, -11.55748, 
    -12.47168, -13.38354, -14.2929, -15.19962, -16.10355, -17.00456, 
    -17.9025, -18.79726, -19.68871, -20.57672, -21.46118, -22.34199, 
    -23.21904, -24.09223, -24.96147, -25.82668, -26.68777, -27.54466, 
    -28.3973, -29.2456, -30.08952, -30.929, -31.76398, -32.59444, -33.42032, 
    -34.2416, -35.05824, -35.87022, -36.67753, -37.48015, -38.27806, 
    -39.07127, -39.85978, -40.64358, -41.42268,
  41.65079, 40.87085, 40.08604, 39.29634, 38.50176, 37.70229, 36.89794, 
    36.08871, 35.27462, 34.45568, 33.63192, 32.80336, 31.97004, 31.132, 
    30.28927, 29.44192, 28.58998, 27.73353, 26.87262, 26.00734, 25.13775, 
    24.26394, 23.386, 22.50403, 21.61812, 20.72838, 19.83493, 18.93789, 
    18.03736, 17.1335, 16.22643, 15.31629, 14.40323, 13.48739, 12.56893, 
    11.64802, 10.72481, 9.799476, 8.872184, 7.943112, 7.012438, 6.080344, 
    5.147013, 4.212631, 3.277388, 2.341473, 1.405076, 0.4683909, -0.4683909, 
    -1.405076, -2.341473, -3.277388, -4.212631, -5.147013, -6.080344, 
    -7.012438, -7.943112, -8.872184, -9.799476, -10.72481, -11.64802, 
    -12.56893, -13.48739, -14.40323, -15.31629, -16.22643, -17.1335, 
    -18.03736, -18.93789, -19.83493, -20.72838, -21.61812, -22.50403, 
    -23.386, -24.26394, -25.13775, -26.00734, -26.87262, -27.73353, 
    -28.58998, -29.44192, -30.28927, -31.132, -31.97004, -32.80336, 
    -33.63192, -34.45568, -35.27462, -36.08871, -36.89794, -37.70229, 
    -38.50176, -39.29634, -40.08604, -40.87085, -41.65079,
  41.87124, 41.09053, 40.30479, 39.51399, 38.71813, 37.9172, 37.11122, 
    36.30017, 35.48409, 34.66297, 33.83684, 33.00574, 32.16968, 31.32872, 
    30.48288, 29.63223, 28.77681, 27.91669, 27.05193, 26.18261, 25.3088, 
    24.43059, 23.54808, 22.66135, 21.77052, 20.87569, 19.97698, 19.07451, 
    18.16841, 17.25882, 16.34587, 15.42971, 14.51049, 13.58837, 12.66351, 
    11.73607, 10.80623, 9.874163, 8.940046, 8.004064, 7.066403, 6.127254, 
    5.186808, 4.245261, 3.30281, 2.359655, 1.415995, 0.472032, -0.472032, 
    -1.415995, -2.359655, -3.30281, -4.245261, -5.186808, -6.127254, 
    -7.066403, -8.004064, -8.940046, -9.874163, -10.80623, -11.73607, 
    -12.66351, -13.58837, -14.51049, -15.42971, -16.34587, -17.25882, 
    -18.16841, -19.07451, -19.97698, -20.87569, -21.77052, -22.66135, 
    -23.54808, -24.43059, -25.3088, -26.18261, -27.05193, -27.91669, 
    -28.77681, -29.63223, -30.48288, -31.32872, -32.16968, -33.00574, 
    -33.83684, -34.66297, -35.48409, -36.30017, -37.11122, -37.9172, 
    -38.71813, -39.51399, -40.30479, -41.09053, -41.87124,
  42.08391, 41.30251, 40.51591, 39.72409, 38.92703, 38.12474, 37.31722, 
    36.50447, 35.68649, 34.86331, 34.03494, 33.20141, 32.36275, 31.519, 
    30.6702, 29.81639, 28.95764, 28.094, 27.22555, 26.35234, 25.47448, 
    24.59204, 23.70512, 22.81381, 21.91823, 21.01848, 20.11469, 19.20699, 
    18.2955, 17.38036, 16.46173, 15.53974, 14.61457, 13.68636, 12.75529, 
    11.82154, 10.88527, 9.946671, 9.005934, 8.063247, 7.118805, 6.172808, 
    5.225454, 4.27695, 3.3275, 2.377314, 1.4266, 0.4755684, -0.4755684, 
    -1.4266, -2.377314, -3.3275, -4.27695, -5.225454, -6.172808, -7.118805, 
    -8.063247, -9.005934, -9.946671, -10.88527, -11.82154, -12.75529, 
    -13.68636, -14.61457, -15.53974, -16.46173, -17.38036, -18.2955, 
    -19.20699, -20.11469, -21.01848, -21.91823, -22.81381, -23.70512, 
    -24.59204, -25.47448, -26.35234, -27.22555, -28.094, -28.95764, 
    -29.81639, -30.6702, -31.519, -32.36275, -33.20141, -34.03494, -34.86331, 
    -35.68649, -36.50447, -37.31722, -38.12474, -38.92703, -39.72409, 
    -40.51591, -41.30251, -42.08391,
  42.28868, 41.50666, 40.71927, 39.9265, 39.12834, 38.32478, 37.51582, 
    36.70145, 35.8817, 35.05656, 34.22607, 33.39024, 32.5491, 31.70269, 
    30.85106, 29.99424, 29.1323, 28.2653, 27.3933, 26.51638, 25.63463, 
    24.74813, 23.85697, 22.96125, 22.0611, 21.15662, 20.24794, 19.33519, 
    18.4185, 17.49802, 16.57389, 15.64629, 14.71535, 13.78126, 12.84419, 
    11.90432, 10.96183, 10.01692, 9.069772, 8.120593, 7.169584, 6.216953, 
    5.262908, 4.307662, 3.35143, 2.394429, 1.436878, 0.478996, -0.478996, 
    -1.436878, -2.394429, -3.35143, -4.307662, -5.262908, -6.216953, 
    -7.169584, -8.120593, -9.069772, -10.01692, -10.96183, -11.90432, 
    -12.84419, -13.78126, -14.71535, -15.64629, -16.57389, -17.49802, 
    -18.4185, -19.33519, -20.24794, -21.15662, -22.0611, -22.96125, 
    -23.85697, -24.74813, -25.63463, -26.51638, -27.3933, -28.2653, -29.1323, 
    -29.99424, -30.85106, -31.70269, -32.5491, -33.39024, -34.22607, 
    -35.05656, -35.8817, -36.70145, -37.51582, -38.32478, -39.12834, 
    -39.9265, -40.71927, -41.50666, -42.28868,
  42.48545, 41.70287, 40.91476, 40.12112, 39.32193, 38.51718, 37.70687, 
    36.891, 36.06956, 35.24258, 34.41008, 33.57207, 32.72858, 31.87964, 
    31.02531, 30.16563, 29.30065, 28.43043, 27.55505, 26.67457, 25.78909, 
    24.89869, 24.00347, 23.10353, 22.19899, 21.28997, 20.37659, 19.45897, 
    18.53728, 17.61165, 16.68224, 15.74921, 14.81272, 13.87296, 12.9301, 
    11.98433, 11.03584, 10.08482, 9.131484, 8.176033, 7.218679, 6.259636, 
    5.299122, 4.337358, 3.374569, 2.41098, 1.446817, 0.4823107, -0.4823107, 
    -1.446817, -2.41098, -3.374569, -4.337358, -5.299122, -6.259636, 
    -7.218679, -8.176033, -9.131484, -10.08482, -11.03584, -11.98433, 
    -12.9301, -13.87296, -14.81272, -15.74921, -16.68224, -17.61165, 
    -18.53728, -19.45897, -20.37659, -21.28997, -22.19899, -23.10353, 
    -24.00347, -24.89869, -25.78909, -26.67457, -27.55505, -28.43043, 
    -29.30065, -30.16563, -31.02531, -31.87964, -32.72858, -33.57207, 
    -34.41008, -35.24258, -36.06956, -36.891, -37.70687, -38.51718, 
    -39.32193, -40.12112, -40.91476, -41.70287, -42.48545,
  42.67411, 41.89101, 41.10225, 40.30781, 39.50767, 38.70182, 37.89024, 
    37.07295, 36.24994, 35.42123, 34.58682, 33.74675, 32.90103, 32.0497, 
    31.19281, 30.3304, 29.46252, 28.58924, 27.71063, 26.82676, 25.93772, 
    25.04359, 24.14449, 23.2405, 22.33176, 21.41838, 20.50048, 19.57821, 
    18.65171, 17.72114, 16.78664, 15.8484, 14.90658, 13.96135, 13.01292, 
    12.06147, 11.10719, 10.1503, 9.190996, 8.229501, 7.266029, 6.300805, 
    5.334054, 4.366004, 3.39689, 2.426945, 1.456406, 0.4855082, -0.4855082, 
    -1.456406, -2.426945, -3.39689, -4.366004, -5.334054, -6.300805, 
    -7.266029, -8.229501, -9.190996, -10.1503, -11.10719, -12.06147, 
    -13.01292, -13.96135, -14.90658, -15.8484, -16.78664, -17.72114, 
    -18.65171, -19.57821, -20.50048, -21.41838, -22.33176, -23.2405, 
    -24.14449, -25.04359, -25.93772, -26.82676, -27.71063, -28.58924, 
    -29.46252, -30.3304, -31.19281, -32.0497, -32.90103, -33.74675, 
    -34.58682, -35.42123, -36.24994, -37.07295, -37.89024, -38.70182, 
    -39.50767, -40.30781, -41.10225, -41.89101, -42.67411,
  42.85454, 42.07099, 41.28164, 40.48646, 39.68544, 38.87856, 38.06581, 
    37.2472, 36.42271, 35.59236, 34.75616, 33.91414, 33.06631, 32.21272, 
    31.3534, 30.4884, 29.61777, 28.74158, 27.8599, 26.9728, 26.08036, 
    25.18268, 24.27987, 23.37202, 22.45926, 21.5417, 20.61949, 19.69276, 
    18.76166, 17.82635, 16.88698, 15.94374, 14.99679, 14.04633, 13.09255, 
    12.13564, 11.17581, 10.21327, 9.248235, 8.280929, 7.311576, 6.340407, 
    5.367657, 4.393563, 3.418365, 2.442306, 1.46563, 0.4885846, -0.4885846, 
    -1.46563, -2.442306, -3.418365, -4.393563, -5.367657, -6.340407, 
    -7.311576, -8.280929, -9.248235, -10.21327, -11.17581, -12.13564, 
    -13.09255, -14.04633, -14.99679, -15.94374, -16.88698, -17.82635, 
    -18.76166, -19.69276, -20.61949, -21.5417, -22.45926, -23.37202, 
    -24.27987, -25.18268, -26.08036, -26.9728, -27.8599, -28.74158, 
    -29.61777, -30.4884, -31.3534, -32.21272, -33.06631, -33.91414, 
    -34.75616, -35.59236, -36.42271, -37.2472, -38.06581, -38.87856, 
    -39.68544, -40.48646, -41.28164, -42.07099, -42.85454,
  43.02665, 42.24269, 41.4528, 40.65696, 39.85512, 39.04729, 38.23346, 
    37.4136, 36.58773, 35.75585, 34.91797, 34.07411, 33.2243, 32.36856, 
    31.50695, 30.6395, 29.76627, 28.88731, 28.00271, 27.11254, 26.21687, 
    25.31582, 24.40947, 23.49794, 22.58134, 21.65982, 20.73348, 19.8025, 
    18.867, 17.92716, 16.98314, 16.03511, 15.08327, 14.1278, 13.16889, 
    12.20676, 11.2416, 10.27365, 9.303126, 8.330251, 7.355261, 6.378393, 
    5.399891, 4.419998, 3.438965, 2.457041, 1.47448, 0.4915359, -0.4915359, 
    -1.47448, -2.457041, -3.438965, -4.419998, -5.399891, -6.378393, 
    -7.355261, -8.330251, -9.303126, -10.27365, -11.2416, -12.20676, 
    -13.16889, -14.1278, -15.08327, -16.03511, -16.98314, -17.92716, -18.867, 
    -19.8025, -20.73348, -21.65982, -22.58134, -23.49794, -24.40947, 
    -25.31582, -26.21687, -27.11254, -28.00271, -28.88731, -29.76627, 
    -30.6395, -31.50695, -32.36856, -33.2243, -34.07411, -34.91797, 
    -35.75585, -36.58773, -37.4136, -38.23346, -39.04729, -39.85512, 
    -40.65696, -41.4528, -42.24269, -43.02665,
  43.19033, 42.40602, 41.61564, 40.81918, 40.0166, 39.20789, 38.39304, 
    37.57203, 36.74487, 35.91155, 35.0721, 34.22652, 33.37484, 32.51709, 
    31.65331, 30.78355, 29.90785, 29.02629, 28.13892, 27.24584, 26.34712, 
    25.44285, 24.53315, 23.61813, 22.69789, 21.77258, 20.84233, 19.90729, 
    18.96761, 18.02345, 17.075, 16.12242, 15.1659, 14.20564, 13.24185, 
    12.27472, 11.30449, 10.33138, 9.355601, 8.377405, 7.397027, 6.414712, 
    5.430711, 4.445276, 3.458663, 2.471131, 1.482942, 0.494358, -0.494358, 
    -1.482942, -2.471131, -3.458663, -4.445276, -5.430711, -6.414712, 
    -7.397027, -8.377405, -9.355601, -10.33138, -11.30449, -12.27472, 
    -13.24185, -14.20564, -15.1659, -16.12242, -17.075, -18.02345, -18.96761, 
    -19.90729, -20.84233, -21.77258, -22.69789, -23.61813, -24.53315, 
    -25.44285, -26.34712, -27.24584, -28.13892, -29.02629, -29.90785, 
    -30.78355, -31.65331, -32.51709, -33.37484, -34.22652, -35.0721, 
    -35.91155, -36.74487, -37.57203, -38.39304, -39.20789, -40.0166, 
    -40.81918, -41.61564, -42.40602, -43.19033,
  43.34549, 42.56086, 41.77005, 40.97303, 40.16977, 39.36025, 38.54446, 
    37.72238, 36.89401, 36.05936, 35.21843, 34.37123, 33.5178, 32.65816, 
    31.79235, 30.92041, 30.04239, 29.15837, 28.2684, 27.37256, 26.47095, 
    25.56366, 24.65079, 23.73245, 22.80877, 21.87987, 20.94591, 20.00702, 
    19.06337, 18.11512, 17.16244, 16.20553, 15.24457, 14.27977, 13.31133, 
    12.33946, 11.3644, 10.38636, 9.40559, 8.422327, 7.436818, 6.449316, 
    5.460076, 4.46936, 3.477432, 2.484558, 1.491006, 0.4970472, -0.4970472, 
    -1.491006, -2.484558, -3.477432, -4.46936, -5.460076, -6.449316, 
    -7.436818, -8.422327, -9.40559, -10.38636, -11.3644, -12.33946, 
    -13.31133, -14.27977, -15.24457, -16.20553, -17.16244, -18.11512, 
    -19.06337, -20.00702, -20.94591, -21.87987, -22.80877, -23.73245, 
    -24.65079, -25.56366, -26.47095, -27.37256, -28.2684, -29.15837, 
    -30.04239, -30.92041, -31.79235, -32.65816, -33.5178, -34.37123, 
    -35.21843, -36.05936, -36.89401, -37.72238, -38.54446, -39.36025, 
    -40.16977, -40.97303, -41.77005, -42.56086, -43.34549,
  43.49203, 42.70713, 41.91592, 41.1184, 40.31451, 39.50425, 38.6876, 
    37.86452, 37.03504, 36.19914, 35.35684, 34.50814, 33.65307, 32.79165, 
    31.92393, 31.04995, 30.16976, 29.28342, 28.391, 27.49258, 26.58825, 
    25.6781, 24.76223, 23.84077, 22.91384, 21.98156, 21.04409, 20.10156, 
    19.15416, 18.20203, 17.24537, 16.28436, 15.3192, 14.35008, 13.37724, 
    12.40088, 11.42123, 10.43853, 9.453025, 8.464956, 7.47458, 6.482156, 
    5.487947, 4.49222, 3.495247, 2.497301, 1.49866, 0.4995998, -0.4995998, 
    -1.49866, -2.497301, -3.495247, -4.49222, -5.487947, -6.482156, -7.47458, 
    -8.464956, -9.453025, -10.43853, -11.42123, -12.40088, -13.37724, 
    -14.35008, -15.3192, -16.28436, -17.24537, -18.20203, -19.15416, 
    -20.10156, -21.04409, -21.98156, -22.91384, -23.84077, -24.76223, 
    -25.6781, -26.58825, -27.49258, -28.391, -29.28342, -30.16976, -31.04995, 
    -31.92393, -32.79165, -33.65307, -34.50814, -35.35684, -36.19914, 
    -37.03504, -37.86452, -38.6876, -39.50425, -40.31451, -41.1184, 
    -41.91592, -42.70713, -43.49203,
  43.62987, 42.84472, 42.05317, 41.25519, 40.45074, 39.63979, 38.82234, 
    37.99836, 37.16784, 36.33079, 35.48721, 34.6371, 33.78051, 32.91744, 
    32.04794, 31.17205, 30.28983, 29.40132, 28.50661, 27.60576, 26.69888, 
    25.78605, 24.86737, 23.94298, 23.01299, 22.07753, 21.13675, 20.19081, 
    19.23986, 18.28409, 17.32367, 16.3588, 15.38967, 14.4165, 13.43949, 
    12.45889, 11.47492, 10.48782, 9.49784, 8.505234, 7.510261, 6.513187, 
    5.514283, 4.513822, 3.512082, 2.509345, 1.505893, 0.502012, -0.502012, 
    -1.505893, -2.509345, -3.512082, -4.513822, -5.514283, -6.513187, 
    -7.510261, -8.505234, -9.49784, -10.48782, -11.47492, -12.45889, 
    -13.43949, -14.4165, -15.38967, -16.3588, -17.32367, -18.28409, 
    -19.23986, -20.19081, -21.13675, -22.07753, -23.01299, -23.94298, 
    -24.86737, -25.78605, -26.69888, -27.60576, -28.50661, -29.40132, 
    -30.28983, -31.17205, -32.04794, -32.91744, -33.78051, -34.6371, 
    -35.48721, -36.33079, -37.16784, -37.99836, -38.82234, -39.63979, 
    -40.45074, -41.25519, -42.05317, -42.84472, -43.62987,
  43.75893, 42.97356, 42.18171, 41.38331, 40.57834, 39.76678, 38.94859, 
    38.12377, 37.2923, 36.45418, 35.60942, 34.75802, 33.90001, 33.03541, 
    32.16426, 31.28659, 30.40247, 29.51195, 28.6151, 27.71199, 26.80272, 
    25.88738, 24.96609, 24.03895, 23.10609, 22.16766, 21.22379, 20.27464, 
    19.32038, 18.36119, 17.39725, 16.42875, 15.4559, 14.47891, 13.49801, 
    12.51342, 11.52539, 10.53416, 9.539974, 8.543103, 7.54381, 6.542367, 
    5.539048, 4.534135, 3.527913, 2.52067, 1.512695, 0.5042805, -0.5042805, 
    -1.512695, -2.52067, -3.527913, -4.534135, -5.539048, -6.542367, 
    -7.54381, -8.543103, -9.539974, -10.53416, -11.52539, -12.51342, 
    -13.49801, -14.47891, -15.4559, -16.42875, -17.39725, -18.36119, 
    -19.32038, -20.27464, -21.22379, -22.16766, -23.10609, -24.03895, 
    -24.96609, -25.88738, -26.80272, -27.71199, -28.6151, -29.51195, 
    -30.40247, -31.28659, -32.16426, -33.03541, -33.90001, -34.75802, 
    -35.60942, -36.45418, -37.2923, -38.12377, -38.94859, -39.76678, 
    -40.57834, -41.38331, -42.18171, -42.97356, -43.75893,
  43.87911, 43.09357, 42.30143, 41.50267, 40.69724, 39.88511, 39.06625, 
    38.24066, 37.40832, 36.56922, 35.72337, 34.87078, 34.01146, 33.14545, 
    32.27277, 31.39346, 30.50758, 29.61518, 28.71634, 27.81114, 26.89966, 
    25.98199, 25.05826, 24.12856, 23.19304, 22.25184, 21.30509, 20.35295, 
    19.39561, 18.43323, 17.466, 16.49412, 15.5178, 14.53725, 13.55271, 
    12.5644, 11.57257, 10.57748, 9.579368, 8.578511, 7.57518, 6.56965, 
    5.562205, 4.55313, 3.542717, 2.53126, 1.519056, 0.5064019, -0.5064019, 
    -1.519056, -2.53126, -3.542717, -4.55313, -5.562205, -6.56965, -7.57518, 
    -8.578511, -9.579368, -10.57748, -11.57257, -12.5644, -13.55271, 
    -14.53725, -15.5178, -16.49412, -17.466, -18.43323, -19.39561, -20.35295, 
    -21.30509, -22.25184, -23.19304, -24.12856, -25.05826, -25.98199, 
    -26.89966, -27.81114, -28.71634, -29.61518, -30.50758, -31.39346, 
    -32.27277, -33.14545, -34.01146, -34.87078, -35.72337, -36.56922, 
    -37.40832, -38.24066, -39.06625, -39.88511, -40.69724, -41.50267, 
    -42.30143, -43.09357, -43.87911,
  43.99035, 43.20465, 42.41228, 41.61318, 40.80733, 39.99469, 39.17523, 
    38.34894, 37.5158, 36.67581, 35.82896, 34.97528, 34.11476, 33.24744, 
    32.37335, 31.49253, 30.60504, 29.71092, 28.81025, 27.90311, 26.98958, 
    26.06977, 25.14377, 24.21172, 23.27374, 22.32997, 21.38055, 20.42565, 
    19.46544, 18.50011, 17.52983, 16.55482, 15.57528, 14.59143, 13.60351, 
    12.61175, 11.6164, 10.61772, 9.615962, 8.611405, 7.604323, 6.594999, 
    5.58372, 4.570779, 3.556473, 2.541101, 1.524966, 0.5083731, -0.5083731, 
    -1.524966, -2.541101, -3.556473, -4.570779, -5.58372, -6.594999, 
    -7.604323, -8.611405, -9.615962, -10.61772, -11.6164, -12.61175, 
    -13.60351, -14.59143, -15.57528, -16.55482, -17.52983, -18.50011, 
    -19.46544, -20.42565, -21.38055, -22.32997, -23.27374, -24.21172, 
    -25.14377, -26.06977, -26.98958, -27.90311, -28.81025, -29.71092, 
    -30.60504, -31.49253, -32.37335, -33.24744, -34.11476, -34.97528, 
    -35.82896, -36.67581, -37.5158, -38.34894, -39.17523, -39.99469, 
    -40.80733, -41.61318, -42.41228, -43.20465, -43.99035,
  44.09258, 43.30674, 42.51416, 41.71477, 40.90854, 40.09544, 39.27544, 
    38.44851, 37.61465, 36.77385, 35.9261, 35.07141, 34.20981, 33.3413, 
    32.46593, 31.58372, 30.69475, 29.79905, 28.89671, 27.98779, 27.07239, 
    26.1506, 25.22254, 24.28832, 23.34808, 22.40195, 21.45008, 20.49264, 
    19.5298, 18.56174, 17.58866, 16.61077, 15.62826, 14.64138, 13.65034, 
    12.6554, 11.65681, 10.65482, 9.649706, 8.641738, 7.631198, 6.618376, 
    5.603562, 4.587056, 3.569159, 2.550177, 1.530417, 0.510191, -0.510191, 
    -1.530417, -2.550177, -3.569159, -4.587056, -5.603562, -6.618376, 
    -7.631198, -8.641738, -9.649706, -10.65482, -11.65681, -12.6554, 
    -13.65034, -14.64138, -15.62826, -16.61077, -17.58866, -18.56174, 
    -19.5298, -20.49264, -21.45008, -22.40195, -23.34808, -24.28832, 
    -25.22254, -26.1506, -27.07239, -27.98779, -28.89671, -29.79905, 
    -30.69475, -31.58372, -32.46593, -33.3413, -34.20981, -35.07141, 
    -35.9261, -36.77385, -37.61465, -38.44851, -39.27544, -40.09544, 
    -40.90854, -41.71477, -42.51416, -43.30674, -44.09258,
  44.18572, 43.39978, 42.60701, 41.80736, 41.0008, 40.18729, 39.3668, 
    38.53931, 37.7048, 36.86326, 36.01469, 35.15911, 34.29651, 33.42693, 
    32.55039, 31.66694, 30.77662, 29.87949, 28.97562, 28.06509, 27.14798, 
    26.2244, 25.29446, 24.35827, 23.41596, 22.46768, 21.51358, 20.55383, 
    19.58859, 18.61805, 17.64242, 16.66188, 15.67667, 14.68701, 13.69314, 
    12.6953, 11.69374, 10.68873, 9.680549, 8.669463, 7.655765, 6.639744, 
    5.6217, 4.601935, 3.580756, 2.558473, 1.535401, 0.511853, -0.511853, 
    -1.535401, -2.558473, -3.580756, -4.601935, -5.6217, -6.639744, 
    -7.655765, -8.669463, -9.680549, -10.68873, -11.69374, -12.6953, 
    -13.69314, -14.68701, -15.67667, -16.66188, -17.64242, -18.61805, 
    -19.58859, -20.55383, -21.51358, -22.46768, -23.41596, -24.35827, 
    -25.29446, -26.2244, -27.14798, -28.06509, -28.97562, -29.87949, 
    -30.77662, -31.66694, -32.55039, -33.42693, -34.29651, -35.15911, 
    -36.01469, -36.86326, -37.7048, -38.53931, -39.3668, -40.18729, -41.0008, 
    -41.80736, -42.60701, -43.39978, -44.18572,
  44.26973, 43.48369, 42.69076, 41.89089, 41.08404, 40.27016, 39.44924, 
    38.62124, 37.78615, 36.94396, 36.09467, 35.23827, 34.37479, 33.50424, 
    32.62666, 31.74208, 30.85055, 29.95214, 29.0469, 28.13491, 27.21628, 
    26.29108, 25.35944, 24.42147, 23.47731, 22.52709, 21.57098, 20.60913, 
    19.64173, 18.66896, 17.69101, 16.7081, 15.72045, 14.72828, 13.73184, 
    12.73137, 11.72714, 10.7194, 9.708443, 8.69454, 7.677984, 6.659072, 
    5.638107, 4.615394, 3.591246, 2.565979, 1.539908, 0.5133564, -0.5133564, 
    -1.539908, -2.565979, -3.591246, -4.615394, -5.638107, -6.659072, 
    -7.677984, -8.69454, -9.708443, -10.7194, -11.72714, -12.73137, 
    -13.73184, -14.72828, -15.72045, -16.7081, -17.69101, -18.66896, 
    -19.64173, -20.60913, -21.57098, -22.52709, -23.47731, -24.42147, 
    -25.35944, -26.29108, -27.21628, -28.13491, -29.0469, -29.95214, 
    -30.85055, -31.74208, -32.62666, -33.50424, -34.37479, -35.23827, 
    -36.09467, -36.94396, -37.78615, -38.62124, -39.44924, -40.27016, 
    -41.08404, -41.89089, -42.69076, -43.48369, -44.26973,
  44.34454, 43.55843, 42.76536, 41.96529, 41.15818, 40.34399, 39.52269, 
    38.69425, 37.85865, 37.01588, 36.16594, 35.30883, 34.44456, 33.57316, 
    32.69466, 31.80908, 30.91648, 30.01692, 29.11047, 28.19719, 27.27719, 
    26.35056, 25.41741, 24.47786, 23.53204, 22.5801, 21.6222, 20.65849, 
    19.68916, 18.71439, 17.73438, 16.74936, 15.75952, 14.76512, 13.76639, 
    12.76358, 11.75696, 10.74679, 9.733348, 8.716929, 7.697824, 6.676331, 
    5.652757, 4.627412, 3.600614, 2.57268, 1.543934, 0.5146989, -0.5146989, 
    -1.543934, -2.57268, -3.600614, -4.627412, -5.652757, -6.676331, 
    -7.697824, -8.716929, -9.733348, -10.74679, -11.75696, -12.76358, 
    -13.76639, -14.76512, -15.75952, -16.74936, -17.73438, -18.71439, 
    -19.68916, -20.65849, -21.6222, -22.5801, -23.53204, -24.47786, 
    -25.41741, -26.35056, -27.27719, -28.19719, -29.11047, -30.01692, 
    -30.91648, -31.80908, -32.69466, -33.57316, -34.44456, -35.30883, 
    -36.16594, -37.01588, -37.85865, -38.69425, -39.52269, -40.34399, 
    -41.15818, -41.96529, -42.76536, -43.55843, -44.34454,
  44.41011, 43.62393, 42.83075, 42.03052, 41.22319, 40.40873, 39.58709, 
    38.75827, 37.92222, 37.07895, 36.22845, 35.37072, 34.50577, 33.63363, 
    32.75431, 31.86786, 30.97433, 30.07377, 29.16625, 28.25185, 27.33065, 
    26.40276, 25.46829, 24.52736, 23.58009, 22.62664, 21.66716, 20.70182, 
    19.7308, 18.75428, 17.77247, 16.78558, 15.79384, 14.79747, 13.79673, 
    12.79187, 11.78315, 10.77084, 9.755226, 8.736598, 7.715252, 6.691492, 
    5.665627, 4.63797, 3.608843, 2.578568, 1.54747, 0.5158784, -0.5158784, 
    -1.54747, -2.578568, -3.608843, -4.63797, -5.665627, -6.691492, 
    -7.715252, -8.736598, -9.755226, -10.77084, -11.78315, -12.79187, 
    -13.79673, -14.79747, -15.79384, -16.78558, -17.77247, -18.75428, 
    -19.7308, -20.70182, -21.66716, -22.62664, -23.58009, -24.52736, 
    -25.46829, -26.40276, -27.33065, -28.25185, -29.16625, -30.07377, 
    -30.97433, -31.86786, -32.75431, -33.63363, -34.50577, -35.37072, 
    -36.22845, -37.07895, -37.92222, -38.75827, -39.58709, -40.40873, 
    -41.22319, -42.03052, -42.83075, -43.62393, -44.41011,
  44.46639, 43.68016, 42.88689, 42.08652, 41.279, 40.46431, 39.6424, 
    38.81324, 37.97682, 37.13312, 36.28214, 35.42388, 34.55835, 33.68556, 
    32.80555, 31.91836, 31.02403, 30.12261, 29.21418, 28.29881, 27.3766, 
    26.44763, 25.51202, 24.5699, 23.62139, 22.66665, 21.70582, 20.73908, 
    19.7666, 18.78858, 17.80522, 16.81673, 15.82335, 14.8253, 13.82283, 
    12.8162, 11.80567, 10.79152, 9.774042, 8.753514, 7.730243, 6.704533, 
    5.676696, 4.647052, 3.615922, 2.583632, 1.550512, 0.5168929, -0.5168929, 
    -1.550512, -2.583632, -3.615922, -4.647052, -5.676696, -6.704533, 
    -7.730243, -8.753514, -9.774042, -10.79152, -11.80567, -12.8162, 
    -13.82283, -14.8253, -15.82335, -16.81673, -17.80522, -18.78858, 
    -19.7666, -20.73908, -21.70582, -22.66665, -23.62139, -24.5699, 
    -25.51202, -26.44763, -27.3766, -28.29881, -29.21418, -30.12261, 
    -31.02403, -31.91836, -32.80555, -33.68556, -34.55835, -35.42388, 
    -36.28214, -37.13312, -37.97682, -38.81324, -39.6424, -40.46431, -41.279, 
    -42.08652, -42.88689, -43.68016, -44.46639,
  44.51335, 43.72708, 42.93373, 42.13324, 41.32558, 40.51069, 39.68855, 
    38.85912, 38.02239, 37.17834, 36.32696, 35.46826, 34.60224, 33.72892, 
    32.84834, 31.96053, 31.06553, 30.1634, 29.25421, 28.33804, 27.41497, 
    26.4851, 25.54855, 24.60544, 23.6559, 22.70007, 21.73811, 20.7702, 
    19.79651, 18.81724, 17.83258, 16.84276, 15.84801, 14.84855, 13.84463, 
    12.83653, 11.8245, 10.80881, 9.789767, 8.767653, 7.742771, 6.715432, 
    5.685948, 4.654643, 3.621838, 2.587865, 1.553055, 0.5177408, -0.5177408, 
    -1.553055, -2.587865, -3.621838, -4.654643, -5.685948, -6.715432, 
    -7.742771, -8.767653, -9.789767, -10.80881, -11.8245, -12.83653, 
    -13.84463, -14.84855, -15.84801, -16.84276, -17.83258, -18.81724, 
    -19.79651, -20.7702, -21.73811, -22.70007, -23.6559, -24.60544, 
    -25.54855, -26.4851, -27.41497, -28.33804, -29.25421, -30.1634, 
    -31.06553, -31.96053, -32.84834, -33.72892, -34.60224, -35.46826, 
    -36.32696, -37.17834, -38.02239, -38.85912, -39.68855, -40.51069, 
    -41.32558, -42.13324, -42.93373, -43.72708, -44.51335,
  44.55096, 43.76466, 42.97124, 42.17067, 41.36288, 40.54784, 39.72552, 
    38.89588, 38.0589, 37.21456, 36.36287, 35.50381, 34.63741, 33.76367, 
    32.88263, 31.99432, 31.09879, 30.19609, 29.28629, 28.36947, 27.44572, 
    26.51514, 25.57783, 24.63392, 23.68355, 22.72686, 21.764, 20.79515, 
    19.82049, 18.84021, 17.85452, 16.86363, 15.86777, 14.86719, 13.86212, 
    12.85283, 11.83959, 10.82268, 9.802377, 8.77899, 7.752818, 6.724172, 
    5.693368, 4.660729, 3.626583, 2.59126, 1.555094, 0.5184209, -0.5184209, 
    -1.555094, -2.59126, -3.626583, -4.660729, -5.693368, -6.724172, 
    -7.752818, -8.77899, -9.802377, -10.82268, -11.83959, -12.85283, 
    -13.86212, -14.86719, -15.86777, -16.86363, -17.85452, -18.84021, 
    -19.82049, -20.79515, -21.764, -22.72686, -23.68355, -24.63392, 
    -25.57783, -26.51514, -27.44572, -28.36947, -29.28629, -30.19609, 
    -31.09879, -31.99432, -32.88263, -33.76367, -34.63741, -35.50381, 
    -36.36287, -37.21456, -38.0589, -38.89588, -39.72552, -40.54784, 
    -41.36288, -42.17067, -42.97124, -43.76466, -44.55096,
  44.57919, 43.79286, 42.9994, 42.19876, 41.39089, 40.57574, 39.75327, 
    38.92347, 38.0863, 37.24176, 36.38982, 35.53051, 34.66381, 33.78976, 
    32.90837, 32.01969, 31.12376, 30.22064, 29.31038, 28.39308, 27.46882, 
    26.5377, 25.59982, 24.65532, 23.70432, 22.74698, 21.78345, 20.81389, 
    19.8385, 18.85747, 17.871, 16.87931, 15.88263, 14.88119, 13.87526, 
    12.86508, 11.85093, 10.83309, 9.811852, 8.787509, 7.760367, 6.73074, 
    5.698944, 4.665304, 3.630148, 2.593811, 1.556626, 0.5189319, -0.5189319, 
    -1.556626, -2.593811, -3.630148, -4.665304, -5.698944, -6.73074, 
    -7.760367, -8.787509, -9.811852, -10.83309, -11.85093, -12.86508, 
    -13.87526, -14.88119, -15.88263, -16.87931, -17.871, -18.85747, -19.8385, 
    -20.81389, -21.78345, -22.74698, -23.70432, -24.65532, -25.59982, 
    -26.5377, -27.46882, -28.39308, -29.31038, -30.22064, -31.12376, 
    -32.01969, -32.90837, -33.78976, -34.66381, -35.53051, -36.38982, 
    -37.24176, -38.0863, -38.92347, -39.75327, -40.57574, -41.39089, 
    -42.19876, -42.9994, -43.79286, -44.57919,
  44.59801, 43.81168, 43.01819, 42.2175, 41.40957, 40.59435, 39.77179, 
    38.94188, 38.10459, 37.2599, 36.40781, 35.54832, 34.68143, 33.80717, 
    32.92555, 32.03662, 31.14043, 30.23702, 29.32646, 28.40884, 27.48424, 
    26.55275, 25.6145, 24.6696, 23.71819, 22.76041, 21.79643, 20.8264, 
    19.85053, 18.86899, 17.882, 16.88978, 15.89254, 14.89054, 13.88403, 
    12.87325, 11.8585, 10.84004, 9.818177, 8.793196, 7.765407, 6.735124, 
    5.702665, 4.668357, 3.632529, 2.595514, 1.557649, 0.519273, -0.519273, 
    -1.557649, -2.595514, -3.632529, -4.668357, -5.702665, -6.735124, 
    -7.765407, -8.793196, -9.818177, -10.84004, -11.8585, -12.87325, 
    -13.88403, -14.89054, -15.89254, -16.88978, -17.882, -18.86899, 
    -19.85053, -20.8264, -21.79643, -22.76041, -23.71819, -24.6696, -25.6145, 
    -26.55275, -27.48424, -28.40884, -29.32646, -30.23702, -31.14043, 
    -32.03662, -32.92555, -33.80717, -34.68143, -35.54832, -36.40781, 
    -37.2599, -38.10459, -38.94188, -39.77179, -40.59435, -41.40957, 
    -42.2175, -43.01819, -43.81168, -44.59801,
  44.60743, 43.82109, 43.02758, 42.22688, 41.41891, 40.60365, 39.78105, 
    38.95109, 38.11374, 37.26898, 36.41681, 35.55723, 34.69025, 33.81588, 
    32.93415, 32.04509, 31.14876, 30.24521, 29.33451, 28.41672, 27.49195, 
    26.56029, 25.62184, 24.67674, 23.72513, 22.76713, 21.80292, 20.83266, 
    19.85655, 18.87476, 17.88751, 16.89501, 15.8975, 14.89522, 13.88841, 
    12.87735, 11.86229, 10.84352, 9.821342, 8.796041, 7.767929, 6.737318, 
    5.704528, 4.669885, 3.63372, 2.596366, 1.55816, 0.5194437, -0.5194437, 
    -1.55816, -2.596366, -3.63372, -4.669885, -5.704528, -6.737318, 
    -7.767929, -8.796041, -9.821342, -10.84352, -11.86229, -12.87735, 
    -13.88841, -14.89522, -15.8975, -16.89501, -17.88751, -18.87476, 
    -19.85655, -20.83266, -21.80292, -22.76713, -23.72513, -24.67674, 
    -25.62184, -26.56029, -27.49195, -28.41672, -29.33451, -30.24521, 
    -31.14876, -32.04509, -32.93415, -33.81588, -34.69025, -35.55723, 
    -36.41681, -37.26898, -38.11374, -38.95109, -39.78105, -40.60365, 
    -41.41891, -42.22688, -43.02758, -43.82109, -44.60743,
  44.60743, 43.82109, 43.02758, 42.22688, 41.41891, 40.60365, 39.78105, 
    38.95109, 38.11374, 37.26898, 36.41681, 35.55723, 34.69025, 33.81588, 
    32.93415, 32.04509, 31.14876, 30.24521, 29.33451, 28.41672, 27.49195, 
    26.56029, 25.62184, 24.67674, 23.72513, 22.76713, 21.80292, 20.83266, 
    19.85655, 18.87476, 17.88751, 16.89501, 15.8975, 14.89522, 13.88841, 
    12.87735, 11.86229, 10.84352, 9.821342, 8.796041, 7.767929, 6.737318, 
    5.704528, 4.669885, 3.63372, 2.596366, 1.55816, 0.5194437, -0.5194437, 
    -1.55816, -2.596366, -3.63372, -4.669885, -5.704528, -6.737318, 
    -7.767929, -8.796041, -9.821342, -10.84352, -11.86229, -12.87735, 
    -13.88841, -14.89522, -15.8975, -16.89501, -17.88751, -18.87476, 
    -19.85655, -20.83266, -21.80292, -22.76713, -23.72513, -24.67674, 
    -25.62184, -26.56029, -27.49195, -28.41672, -29.33451, -30.24521, 
    -31.14876, -32.04509, -32.93415, -33.81588, -34.69025, -35.55723, 
    -36.41681, -37.26898, -38.11374, -38.95109, -39.78105, -40.60365, 
    -41.41891, -42.22688, -43.02758, -43.82109, -44.60743,
  44.59801, 43.81168, 43.01819, 42.2175, 41.40957, 40.59435, 39.77179, 
    38.94188, 38.10459, 37.2599, 36.40781, 35.54832, 34.68143, 33.80717, 
    32.92555, 32.03662, 31.14043, 30.23702, 29.32646, 28.40884, 27.48424, 
    26.55275, 25.6145, 24.6696, 23.71819, 22.76041, 21.79643, 20.8264, 
    19.85053, 18.86899, 17.882, 16.88978, 15.89254, 14.89054, 13.88403, 
    12.87325, 11.8585, 10.84004, 9.818177, 8.793196, 7.765407, 6.735124, 
    5.702665, 4.668357, 3.632529, 2.595514, 1.557649, 0.519273, -0.519273, 
    -1.557649, -2.595514, -3.632529, -4.668357, -5.702665, -6.735124, 
    -7.765407, -8.793196, -9.818177, -10.84004, -11.8585, -12.87325, 
    -13.88403, -14.89054, -15.89254, -16.88978, -17.882, -18.86899, 
    -19.85053, -20.8264, -21.79643, -22.76041, -23.71819, -24.6696, -25.6145, 
    -26.55275, -27.48424, -28.40884, -29.32646, -30.23702, -31.14043, 
    -32.03662, -32.92555, -33.80717, -34.68143, -35.54832, -36.40781, 
    -37.2599, -38.10459, -38.94188, -39.77179, -40.59435, -41.40957, 
    -42.2175, -43.01819, -43.81168, -44.59801,
  44.57919, 43.79286, 42.9994, 42.19876, 41.39089, 40.57574, 39.75327, 
    38.92347, 38.0863, 37.24176, 36.38982, 35.53051, 34.66381, 33.78976, 
    32.90837, 32.01969, 31.12376, 30.22064, 29.31038, 28.39308, 27.46882, 
    26.5377, 25.59982, 24.65532, 23.70432, 22.74698, 21.78345, 20.81389, 
    19.8385, 18.85747, 17.871, 16.87931, 15.88263, 14.88119, 13.87526, 
    12.86508, 11.85093, 10.83309, 9.811852, 8.787509, 7.760367, 6.73074, 
    5.698944, 4.665304, 3.630148, 2.593811, 1.556626, 0.5189319, -0.5189319, 
    -1.556626, -2.593811, -3.630148, -4.665304, -5.698944, -6.73074, 
    -7.760367, -8.787509, -9.811852, -10.83309, -11.85093, -12.86508, 
    -13.87526, -14.88119, -15.88263, -16.87931, -17.871, -18.85747, -19.8385, 
    -20.81389, -21.78345, -22.74698, -23.70432, -24.65532, -25.59982, 
    -26.5377, -27.46882, -28.39308, -29.31038, -30.22064, -31.12376, 
    -32.01969, -32.90837, -33.78976, -34.66381, -35.53051, -36.38982, 
    -37.24176, -38.0863, -38.92347, -39.75327, -40.57574, -41.39089, 
    -42.19876, -42.9994, -43.79286, -44.57919,
  44.55096, 43.76466, 42.97124, 42.17067, 41.36288, 40.54784, 39.72552, 
    38.89588, 38.0589, 37.21456, 36.36287, 35.50381, 34.63741, 33.76367, 
    32.88263, 31.99432, 31.09879, 30.19609, 29.28629, 28.36947, 27.44572, 
    26.51514, 25.57783, 24.63392, 23.68355, 22.72686, 21.764, 20.79515, 
    19.82049, 18.84021, 17.85452, 16.86363, 15.86777, 14.86719, 13.86212, 
    12.85283, 11.83959, 10.82268, 9.802377, 8.77899, 7.752818, 6.724172, 
    5.693368, 4.660729, 3.626583, 2.59126, 1.555094, 0.5184209, -0.5184209, 
    -1.555094, -2.59126, -3.626583, -4.660729, -5.693368, -6.724172, 
    -7.752818, -8.77899, -9.802377, -10.82268, -11.83959, -12.85283, 
    -13.86212, -14.86719, -15.86777, -16.86363, -17.85452, -18.84021, 
    -19.82049, -20.79515, -21.764, -22.72686, -23.68355, -24.63392, 
    -25.57783, -26.51514, -27.44572, -28.36947, -29.28629, -30.19609, 
    -31.09879, -31.99432, -32.88263, -33.76367, -34.63741, -35.50381, 
    -36.36287, -37.21456, -38.0589, -38.89588, -39.72552, -40.54784, 
    -41.36288, -42.17067, -42.97124, -43.76466, -44.55096,
  44.51335, 43.72708, 42.93373, 42.13324, 41.32558, 40.51069, 39.68855, 
    38.85912, 38.02239, 37.17834, 36.32696, 35.46826, 34.60224, 33.72892, 
    32.84834, 31.96053, 31.06553, 30.1634, 29.25421, 28.33804, 27.41497, 
    26.4851, 25.54855, 24.60544, 23.6559, 22.70007, 21.73811, 20.7702, 
    19.79651, 18.81724, 17.83258, 16.84276, 15.84801, 14.84855, 13.84463, 
    12.83653, 11.8245, 10.80881, 9.789767, 8.767653, 7.742771, 6.715432, 
    5.685948, 4.654643, 3.621838, 2.587865, 1.553055, 0.5177408, -0.5177408, 
    -1.553055, -2.587865, -3.621838, -4.654643, -5.685948, -6.715432, 
    -7.742771, -8.767653, -9.789767, -10.80881, -11.8245, -12.83653, 
    -13.84463, -14.84855, -15.84801, -16.84276, -17.83258, -18.81724, 
    -19.79651, -20.7702, -21.73811, -22.70007, -23.6559, -24.60544, 
    -25.54855, -26.4851, -27.41497, -28.33804, -29.25421, -30.1634, 
    -31.06553, -31.96053, -32.84834, -33.72892, -34.60224, -35.46826, 
    -36.32696, -37.17834, -38.02239, -38.85912, -39.68855, -40.51069, 
    -41.32558, -42.13324, -42.93373, -43.72708, -44.51335,
  44.46639, 43.68016, 42.88689, 42.08652, 41.279, 40.46431, 39.6424, 
    38.81324, 37.97682, 37.13312, 36.28214, 35.42388, 34.55835, 33.68556, 
    32.80555, 31.91836, 31.02403, 30.12261, 29.21418, 28.29881, 27.3766, 
    26.44763, 25.51202, 24.5699, 23.62139, 22.66665, 21.70582, 20.73908, 
    19.7666, 18.78858, 17.80522, 16.81673, 15.82335, 14.8253, 13.82283, 
    12.8162, 11.80567, 10.79152, 9.774042, 8.753514, 7.730243, 6.704533, 
    5.676696, 4.647052, 3.615922, 2.583632, 1.550512, 0.5168929, -0.5168929, 
    -1.550512, -2.583632, -3.615922, -4.647052, -5.676696, -6.704533, 
    -7.730243, -8.753514, -9.774042, -10.79152, -11.80567, -12.8162, 
    -13.82283, -14.8253, -15.82335, -16.81673, -17.80522, -18.78858, 
    -19.7666, -20.73908, -21.70582, -22.66665, -23.62139, -24.5699, 
    -25.51202, -26.44763, -27.3766, -28.29881, -29.21418, -30.12261, 
    -31.02403, -31.91836, -32.80555, -33.68556, -34.55835, -35.42388, 
    -36.28214, -37.13312, -37.97682, -38.81324, -39.6424, -40.46431, -41.279, 
    -42.08652, -42.88689, -43.68016, -44.46639,
  44.41011, 43.62393, 42.83075, 42.03052, 41.22319, 40.40873, 39.58709, 
    38.75827, 37.92222, 37.07895, 36.22845, 35.37072, 34.50577, 33.63363, 
    32.75431, 31.86786, 30.97433, 30.07377, 29.16625, 28.25185, 27.33065, 
    26.40276, 25.46829, 24.52736, 23.58009, 22.62664, 21.66716, 20.70182, 
    19.7308, 18.75428, 17.77247, 16.78558, 15.79384, 14.79747, 13.79673, 
    12.79187, 11.78315, 10.77084, 9.755226, 8.736598, 7.715252, 6.691492, 
    5.665627, 4.63797, 3.608843, 2.578568, 1.54747, 0.5158784, -0.5158784, 
    -1.54747, -2.578568, -3.608843, -4.63797, -5.665627, -6.691492, 
    -7.715252, -8.736598, -9.755226, -10.77084, -11.78315, -12.79187, 
    -13.79673, -14.79747, -15.79384, -16.78558, -17.77247, -18.75428, 
    -19.7308, -20.70182, -21.66716, -22.62664, -23.58009, -24.52736, 
    -25.46829, -26.40276, -27.33065, -28.25185, -29.16625, -30.07377, 
    -30.97433, -31.86786, -32.75431, -33.63363, -34.50577, -35.37072, 
    -36.22845, -37.07895, -37.92222, -38.75827, -39.58709, -40.40873, 
    -41.22319, -42.03052, -42.83075, -43.62393, -44.41011,
  44.34454, 43.55843, 42.76536, 41.96529, 41.15818, 40.34399, 39.52269, 
    38.69425, 37.85865, 37.01588, 36.16594, 35.30883, 34.44456, 33.57316, 
    32.69466, 31.80908, 30.91648, 30.01692, 29.11047, 28.19719, 27.27719, 
    26.35056, 25.41741, 24.47786, 23.53204, 22.5801, 21.6222, 20.65849, 
    19.68916, 18.71439, 17.73438, 16.74936, 15.75952, 14.76512, 13.76639, 
    12.76358, 11.75696, 10.74679, 9.733348, 8.716929, 7.697824, 6.676331, 
    5.652757, 4.627412, 3.600614, 2.57268, 1.543934, 0.5146989, -0.5146989, 
    -1.543934, -2.57268, -3.600614, -4.627412, -5.652757, -6.676331, 
    -7.697824, -8.716929, -9.733348, -10.74679, -11.75696, -12.76358, 
    -13.76639, -14.76512, -15.75952, -16.74936, -17.73438, -18.71439, 
    -19.68916, -20.65849, -21.6222, -22.5801, -23.53204, -24.47786, 
    -25.41741, -26.35056, -27.27719, -28.19719, -29.11047, -30.01692, 
    -30.91648, -31.80908, -32.69466, -33.57316, -34.44456, -35.30883, 
    -36.16594, -37.01588, -37.85865, -38.69425, -39.52269, -40.34399, 
    -41.15818, -41.96529, -42.76536, -43.55843, -44.34454,
  44.26973, 43.48369, 42.69076, 41.89089, 41.08404, 40.27016, 39.44924, 
    38.62124, 37.78615, 36.94396, 36.09467, 35.23827, 34.37479, 33.50424, 
    32.62666, 31.74208, 30.85055, 29.95214, 29.0469, 28.13491, 27.21628, 
    26.29108, 25.35944, 24.42147, 23.47731, 22.52709, 21.57098, 20.60913, 
    19.64173, 18.66896, 17.69101, 16.7081, 15.72045, 14.72828, 13.73184, 
    12.73137, 11.72714, 10.7194, 9.708443, 8.69454, 7.677984, 6.659072, 
    5.638107, 4.615394, 3.591246, 2.565979, 1.539908, 0.5133564, -0.5133564, 
    -1.539908, -2.565979, -3.591246, -4.615394, -5.638107, -6.659072, 
    -7.677984, -8.69454, -9.708443, -10.7194, -11.72714, -12.73137, 
    -13.73184, -14.72828, -15.72045, -16.7081, -17.69101, -18.66896, 
    -19.64173, -20.60913, -21.57098, -22.52709, -23.47731, -24.42147, 
    -25.35944, -26.29108, -27.21628, -28.13491, -29.0469, -29.95214, 
    -30.85055, -31.74208, -32.62666, -33.50424, -34.37479, -35.23827, 
    -36.09467, -36.94396, -37.78615, -38.62124, -39.44924, -40.27016, 
    -41.08404, -41.89089, -42.69076, -43.48369, -44.26973,
  44.18572, 43.39978, 42.60701, 41.80736, 41.0008, 40.18729, 39.3668, 
    38.53931, 37.7048, 36.86326, 36.01469, 35.15911, 34.29651, 33.42693, 
    32.55039, 31.66694, 30.77662, 29.87949, 28.97562, 28.06509, 27.14798, 
    26.2244, 25.29446, 24.35827, 23.41596, 22.46768, 21.51358, 20.55383, 
    19.58859, 18.61805, 17.64242, 16.66188, 15.67667, 14.68701, 13.69314, 
    12.6953, 11.69374, 10.68873, 9.680549, 8.669463, 7.655765, 6.639744, 
    5.6217, 4.601935, 3.580756, 2.558473, 1.535401, 0.511853, -0.511853, 
    -1.535401, -2.558473, -3.580756, -4.601935, -5.6217, -6.639744, 
    -7.655765, -8.669463, -9.680549, -10.68873, -11.69374, -12.6953, 
    -13.69314, -14.68701, -15.67667, -16.66188, -17.64242, -18.61805, 
    -19.58859, -20.55383, -21.51358, -22.46768, -23.41596, -24.35827, 
    -25.29446, -26.2244, -27.14798, -28.06509, -28.97562, -29.87949, 
    -30.77662, -31.66694, -32.55039, -33.42693, -34.29651, -35.15911, 
    -36.01469, -36.86326, -37.7048, -38.53931, -39.3668, -40.18729, -41.0008, 
    -41.80736, -42.60701, -43.39978, -44.18572,
  44.09258, 43.30674, 42.51416, 41.71477, 40.90854, 40.09544, 39.27544, 
    38.44851, 37.61465, 36.77385, 35.9261, 35.07141, 34.20981, 33.3413, 
    32.46593, 31.58372, 30.69475, 29.79905, 28.89671, 27.98779, 27.07239, 
    26.1506, 25.22254, 24.28832, 23.34808, 22.40195, 21.45008, 20.49264, 
    19.5298, 18.56174, 17.58866, 16.61077, 15.62826, 14.64138, 13.65034, 
    12.6554, 11.65681, 10.65482, 9.649706, 8.641738, 7.631198, 6.618376, 
    5.603562, 4.587056, 3.569159, 2.550177, 1.530417, 0.510191, -0.510191, 
    -1.530417, -2.550177, -3.569159, -4.587056, -5.603562, -6.618376, 
    -7.631198, -8.641738, -9.649706, -10.65482, -11.65681, -12.6554, 
    -13.65034, -14.64138, -15.62826, -16.61077, -17.58866, -18.56174, 
    -19.5298, -20.49264, -21.45008, -22.40195, -23.34808, -24.28832, 
    -25.22254, -26.1506, -27.07239, -27.98779, -28.89671, -29.79905, 
    -30.69475, -31.58372, -32.46593, -33.3413, -34.20981, -35.07141, 
    -35.9261, -36.77385, -37.61465, -38.44851, -39.27544, -40.09544, 
    -40.90854, -41.71477, -42.51416, -43.30674, -44.09258,
  43.99035, 43.20465, 42.41228, 41.61318, 40.80733, 39.99469, 39.17523, 
    38.34894, 37.5158, 36.67581, 35.82896, 34.97528, 34.11476, 33.24744, 
    32.37335, 31.49253, 30.60504, 29.71092, 28.81025, 27.90311, 26.98958, 
    26.06977, 25.14377, 24.21172, 23.27374, 22.32997, 21.38055, 20.42565, 
    19.46544, 18.50011, 17.52983, 16.55482, 15.57528, 14.59143, 13.60351, 
    12.61175, 11.6164, 10.61772, 9.615962, 8.611405, 7.604323, 6.594999, 
    5.58372, 4.570779, 3.556473, 2.541101, 1.524966, 0.5083731, -0.5083731, 
    -1.524966, -2.541101, -3.556473, -4.570779, -5.58372, -6.594999, 
    -7.604323, -8.611405, -9.615962, -10.61772, -11.6164, -12.61175, 
    -13.60351, -14.59143, -15.57528, -16.55482, -17.52983, -18.50011, 
    -19.46544, -20.42565, -21.38055, -22.32997, -23.27374, -24.21172, 
    -25.14377, -26.06977, -26.98958, -27.90311, -28.81025, -29.71092, 
    -30.60504, -31.49253, -32.37335, -33.24744, -34.11476, -34.97528, 
    -35.82896, -36.67581, -37.5158, -38.34894, -39.17523, -39.99469, 
    -40.80733, -41.61318, -42.41228, -43.20465, -43.99035,
  43.87911, 43.09357, 42.30143, 41.50267, 40.69724, 39.88511, 39.06625, 
    38.24066, 37.40832, 36.56922, 35.72337, 34.87078, 34.01146, 33.14545, 
    32.27277, 31.39346, 30.50758, 29.61518, 28.71634, 27.81114, 26.89966, 
    25.98199, 25.05826, 24.12856, 23.19304, 22.25184, 21.30509, 20.35295, 
    19.39561, 18.43323, 17.466, 16.49412, 15.5178, 14.53725, 13.55271, 
    12.5644, 11.57257, 10.57748, 9.579368, 8.578511, 7.57518, 6.56965, 
    5.562205, 4.55313, 3.542717, 2.53126, 1.519056, 0.5064019, -0.5064019, 
    -1.519056, -2.53126, -3.542717, -4.55313, -5.562205, -6.56965, -7.57518, 
    -8.578511, -9.579368, -10.57748, -11.57257, -12.5644, -13.55271, 
    -14.53725, -15.5178, -16.49412, -17.466, -18.43323, -19.39561, -20.35295, 
    -21.30509, -22.25184, -23.19304, -24.12856, -25.05826, -25.98199, 
    -26.89966, -27.81114, -28.71634, -29.61518, -30.50758, -31.39346, 
    -32.27277, -33.14545, -34.01146, -34.87078, -35.72337, -36.56922, 
    -37.40832, -38.24066, -39.06625, -39.88511, -40.69724, -41.50267, 
    -42.30143, -43.09357, -43.87911,
  43.75893, 42.97356, 42.18171, 41.38331, 40.57834, 39.76678, 38.94859, 
    38.12377, 37.2923, 36.45418, 35.60942, 34.75802, 33.90001, 33.03541, 
    32.16426, 31.28659, 30.40247, 29.51195, 28.6151, 27.71199, 26.80272, 
    25.88738, 24.96609, 24.03895, 23.10609, 22.16766, 21.22379, 20.27464, 
    19.32038, 18.36119, 17.39725, 16.42875, 15.4559, 14.47891, 13.49801, 
    12.51342, 11.52539, 10.53416, 9.539974, 8.543103, 7.54381, 6.542367, 
    5.539048, 4.534135, 3.527913, 2.52067, 1.512695, 0.5042805, -0.5042805, 
    -1.512695, -2.52067, -3.527913, -4.534135, -5.539048, -6.542367, 
    -7.54381, -8.543103, -9.539974, -10.53416, -11.52539, -12.51342, 
    -13.49801, -14.47891, -15.4559, -16.42875, -17.39725, -18.36119, 
    -19.32038, -20.27464, -21.22379, -22.16766, -23.10609, -24.03895, 
    -24.96609, -25.88738, -26.80272, -27.71199, -28.6151, -29.51195, 
    -30.40247, -31.28659, -32.16426, -33.03541, -33.90001, -34.75802, 
    -35.60942, -36.45418, -37.2923, -38.12377, -38.94859, -39.76678, 
    -40.57834, -41.38331, -42.18171, -42.97356, -43.75893,
  43.62987, 42.84472, 42.05317, 41.25519, 40.45074, 39.63979, 38.82234, 
    37.99836, 37.16784, 36.33079, 35.48721, 34.6371, 33.78051, 32.91744, 
    32.04794, 31.17205, 30.28983, 29.40132, 28.50661, 27.60576, 26.69888, 
    25.78605, 24.86737, 23.94298, 23.01299, 22.07753, 21.13675, 20.19081, 
    19.23986, 18.28409, 17.32367, 16.3588, 15.38967, 14.4165, 13.43949, 
    12.45889, 11.47492, 10.48782, 9.49784, 8.505234, 7.510261, 6.513187, 
    5.514283, 4.513822, 3.512082, 2.509345, 1.505893, 0.502012, -0.502012, 
    -1.505893, -2.509345, -3.512082, -4.513822, -5.514283, -6.513187, 
    -7.510261, -8.505234, -9.49784, -10.48782, -11.47492, -12.45889, 
    -13.43949, -14.4165, -15.38967, -16.3588, -17.32367, -18.28409, 
    -19.23986, -20.19081, -21.13675, -22.07753, -23.01299, -23.94298, 
    -24.86737, -25.78605, -26.69888, -27.60576, -28.50661, -29.40132, 
    -30.28983, -31.17205, -32.04794, -32.91744, -33.78051, -34.6371, 
    -35.48721, -36.33079, -37.16784, -37.99836, -38.82234, -39.63979, 
    -40.45074, -41.25519, -42.05317, -42.84472, -43.62987,
  43.49203, 42.70713, 41.91592, 41.1184, 40.31451, 39.50425, 38.6876, 
    37.86452, 37.03504, 36.19914, 35.35684, 34.50814, 33.65307, 32.79165, 
    31.92393, 31.04995, 30.16976, 29.28342, 28.391, 27.49258, 26.58825, 
    25.6781, 24.76223, 23.84077, 22.91384, 21.98156, 21.04409, 20.10156, 
    19.15416, 18.20203, 17.24537, 16.28436, 15.3192, 14.35008, 13.37724, 
    12.40088, 11.42123, 10.43853, 9.453025, 8.464956, 7.47458, 6.482156, 
    5.487947, 4.49222, 3.495247, 2.497301, 1.49866, 0.4995998, -0.4995998, 
    -1.49866, -2.497301, -3.495247, -4.49222, -5.487947, -6.482156, -7.47458, 
    -8.464956, -9.453025, -10.43853, -11.42123, -12.40088, -13.37724, 
    -14.35008, -15.3192, -16.28436, -17.24537, -18.20203, -19.15416, 
    -20.10156, -21.04409, -21.98156, -22.91384, -23.84077, -24.76223, 
    -25.6781, -26.58825, -27.49258, -28.391, -29.28342, -30.16976, -31.04995, 
    -31.92393, -32.79165, -33.65307, -34.50814, -35.35684, -36.19914, 
    -37.03504, -37.86452, -38.6876, -39.50425, -40.31451, -41.1184, 
    -41.91592, -42.70713, -43.49203,
  43.34549, 42.56086, 41.77005, 40.97303, 40.16977, 39.36025, 38.54446, 
    37.72238, 36.89401, 36.05936, 35.21843, 34.37123, 33.5178, 32.65816, 
    31.79235, 30.92041, 30.04239, 29.15837, 28.2684, 27.37256, 26.47095, 
    25.56366, 24.65079, 23.73245, 22.80877, 21.87987, 20.94591, 20.00702, 
    19.06337, 18.11512, 17.16244, 16.20553, 15.24457, 14.27977, 13.31133, 
    12.33946, 11.3644, 10.38636, 9.40559, 8.422327, 7.436818, 6.449316, 
    5.460076, 4.46936, 3.477432, 2.484558, 1.491006, 0.4970472, -0.4970472, 
    -1.491006, -2.484558, -3.477432, -4.46936, -5.460076, -6.449316, 
    -7.436818, -8.422327, -9.40559, -10.38636, -11.3644, -12.33946, 
    -13.31133, -14.27977, -15.24457, -16.20553, -17.16244, -18.11512, 
    -19.06337, -20.00702, -20.94591, -21.87987, -22.80877, -23.73245, 
    -24.65079, -25.56366, -26.47095, -27.37256, -28.2684, -29.15837, 
    -30.04239, -30.92041, -31.79235, -32.65816, -33.5178, -34.37123, 
    -35.21843, -36.05936, -36.89401, -37.72238, -38.54446, -39.36025, 
    -40.16977, -40.97303, -41.77005, -42.56086, -43.34549,
  43.19033, 42.40602, 41.61564, 40.81918, 40.0166, 39.20789, 38.39304, 
    37.57203, 36.74487, 35.91155, 35.0721, 34.22652, 33.37484, 32.51709, 
    31.65331, 30.78355, 29.90785, 29.02629, 28.13892, 27.24584, 26.34712, 
    25.44285, 24.53315, 23.61813, 22.69789, 21.77258, 20.84233, 19.90729, 
    18.96761, 18.02345, 17.075, 16.12242, 15.1659, 14.20564, 13.24185, 
    12.27472, 11.30449, 10.33138, 9.355601, 8.377405, 7.397027, 6.414712, 
    5.430711, 4.445276, 3.458663, 2.471131, 1.482942, 0.494358, -0.494358, 
    -1.482942, -2.471131, -3.458663, -4.445276, -5.430711, -6.414712, 
    -7.397027, -8.377405, -9.355601, -10.33138, -11.30449, -12.27472, 
    -13.24185, -14.20564, -15.1659, -16.12242, -17.075, -18.02345, -18.96761, 
    -19.90729, -20.84233, -21.77258, -22.69789, -23.61813, -24.53315, 
    -25.44285, -26.34712, -27.24584, -28.13892, -29.02629, -29.90785, 
    -30.78355, -31.65331, -32.51709, -33.37484, -34.22652, -35.0721, 
    -35.91155, -36.74487, -37.57203, -38.39304, -39.20789, -40.0166, 
    -40.81918, -41.61564, -42.40602, -43.19033,
  43.02665, 42.24269, 41.4528, 40.65696, 39.85512, 39.04729, 38.23346, 
    37.4136, 36.58773, 35.75585, 34.91797, 34.07411, 33.2243, 32.36856, 
    31.50695, 30.6395, 29.76627, 28.88731, 28.00271, 27.11254, 26.21687, 
    25.31582, 24.40947, 23.49794, 22.58134, 21.65982, 20.73348, 19.8025, 
    18.867, 17.92716, 16.98314, 16.03511, 15.08327, 14.1278, 13.16889, 
    12.20676, 11.2416, 10.27365, 9.303126, 8.330251, 7.355261, 6.378393, 
    5.399891, 4.419998, 3.438965, 2.457041, 1.47448, 0.4915359, -0.4915359, 
    -1.47448, -2.457041, -3.438965, -4.419998, -5.399891, -6.378393, 
    -7.355261, -8.330251, -9.303126, -10.27365, -11.2416, -12.20676, 
    -13.16889, -14.1278, -15.08327, -16.03511, -16.98314, -17.92716, -18.867, 
    -19.8025, -20.73348, -21.65982, -22.58134, -23.49794, -24.40947, 
    -25.31582, -26.21687, -27.11254, -28.00271, -28.88731, -29.76627, 
    -30.6395, -31.50695, -32.36856, -33.2243, -34.07411, -34.91797, 
    -35.75585, -36.58773, -37.4136, -38.23346, -39.04729, -39.85512, 
    -40.65696, -41.4528, -42.24269, -43.02665,
  42.85454, 42.07099, 41.28164, 40.48646, 39.68544, 38.87856, 38.06581, 
    37.2472, 36.42271, 35.59236, 34.75616, 33.91414, 33.06631, 32.21272, 
    31.3534, 30.4884, 29.61777, 28.74158, 27.8599, 26.9728, 26.08036, 
    25.18268, 24.27987, 23.37202, 22.45926, 21.5417, 20.61949, 19.69276, 
    18.76166, 17.82635, 16.88698, 15.94374, 14.99679, 14.04633, 13.09255, 
    12.13564, 11.17581, 10.21327, 9.248235, 8.280929, 7.311576, 6.340407, 
    5.367657, 4.393563, 3.418365, 2.442306, 1.46563, 0.4885846, -0.4885846, 
    -1.46563, -2.442306, -3.418365, -4.393563, -5.367657, -6.340407, 
    -7.311576, -8.280929, -9.248235, -10.21327, -11.17581, -12.13564, 
    -13.09255, -14.04633, -14.99679, -15.94374, -16.88698, -17.82635, 
    -18.76166, -19.69276, -20.61949, -21.5417, -22.45926, -23.37202, 
    -24.27987, -25.18268, -26.08036, -26.9728, -27.8599, -28.74158, 
    -29.61777, -30.4884, -31.3534, -32.21272, -33.06631, -33.91414, 
    -34.75616, -35.59236, -36.42271, -37.2472, -38.06581, -38.87856, 
    -39.68544, -40.48646, -41.28164, -42.07099, -42.85454,
  42.67411, 41.89101, 41.10225, 40.30781, 39.50767, 38.70182, 37.89024, 
    37.07295, 36.24994, 35.42123, 34.58682, 33.74675, 32.90103, 32.0497, 
    31.19281, 30.3304, 29.46252, 28.58924, 27.71063, 26.82676, 25.93772, 
    25.04359, 24.14449, 23.2405, 22.33176, 21.41838, 20.50048, 19.57821, 
    18.65171, 17.72114, 16.78664, 15.8484, 14.90658, 13.96135, 13.01292, 
    12.06147, 11.10719, 10.1503, 9.190996, 8.229501, 7.266029, 6.300805, 
    5.334054, 4.366004, 3.39689, 2.426945, 1.456406, 0.4855082, -0.4855082, 
    -1.456406, -2.426945, -3.39689, -4.366004, -5.334054, -6.300805, 
    -7.266029, -8.229501, -9.190996, -10.1503, -11.10719, -12.06147, 
    -13.01292, -13.96135, -14.90658, -15.8484, -16.78664, -17.72114, 
    -18.65171, -19.57821, -20.50048, -21.41838, -22.33176, -23.2405, 
    -24.14449, -25.04359, -25.93772, -26.82676, -27.71063, -28.58924, 
    -29.46252, -30.3304, -31.19281, -32.0497, -32.90103, -33.74675, 
    -34.58682, -35.42123, -36.24994, -37.07295, -37.89024, -38.70182, 
    -39.50767, -40.30781, -41.10225, -41.89101, -42.67411,
  42.48545, 41.70287, 40.91476, 40.12112, 39.32193, 38.51718, 37.70687, 
    36.891, 36.06956, 35.24258, 34.41008, 33.57207, 32.72858, 31.87964, 
    31.02531, 30.16563, 29.30065, 28.43043, 27.55505, 26.67457, 25.78909, 
    24.89869, 24.00347, 23.10353, 22.19899, 21.28997, 20.37659, 19.45897, 
    18.53728, 17.61165, 16.68224, 15.74921, 14.81272, 13.87296, 12.9301, 
    11.98433, 11.03584, 10.08482, 9.131484, 8.176033, 7.218679, 6.259636, 
    5.299122, 4.337358, 3.374569, 2.41098, 1.446817, 0.4823107, -0.4823107, 
    -1.446817, -2.41098, -3.374569, -4.337358, -5.299122, -6.259636, 
    -7.218679, -8.176033, -9.131484, -10.08482, -11.03584, -11.98433, 
    -12.9301, -13.87296, -14.81272, -15.74921, -16.68224, -17.61165, 
    -18.53728, -19.45897, -20.37659, -21.28997, -22.19899, -23.10353, 
    -24.00347, -24.89869, -25.78909, -26.67457, -27.55505, -28.43043, 
    -29.30065, -30.16563, -31.02531, -31.87964, -32.72858, -33.57207, 
    -34.41008, -35.24258, -36.06956, -36.891, -37.70687, -38.51718, 
    -39.32193, -40.12112, -40.91476, -41.70287, -42.48545,
  42.28868, 41.50666, 40.71927, 39.9265, 39.12834, 38.32478, 37.51582, 
    36.70145, 35.8817, 35.05656, 34.22607, 33.39024, 32.5491, 31.70269, 
    30.85106, 29.99424, 29.1323, 28.2653, 27.3933, 26.51638, 25.63463, 
    24.74813, 23.85697, 22.96125, 22.0611, 21.15662, 20.24794, 19.33519, 
    18.4185, 17.49802, 16.57389, 15.64629, 14.71535, 13.78126, 12.84419, 
    11.90432, 10.96183, 10.01692, 9.069772, 8.120593, 7.169584, 6.216953, 
    5.262908, 4.307662, 3.35143, 2.394429, 1.436878, 0.478996, -0.478996, 
    -1.436878, -2.394429, -3.35143, -4.307662, -5.262908, -6.216953, 
    -7.169584, -8.120593, -9.069772, -10.01692, -10.96183, -11.90432, 
    -12.84419, -13.78126, -14.71535, -15.64629, -16.57389, -17.49802, 
    -18.4185, -19.33519, -20.24794, -21.15662, -22.0611, -22.96125, 
    -23.85697, -24.74813, -25.63463, -26.51638, -27.3933, -28.2653, -29.1323, 
    -29.99424, -30.85106, -31.70269, -32.5491, -33.39024, -34.22607, 
    -35.05656, -35.8817, -36.70145, -37.51582, -38.32478, -39.12834, 
    -39.9265, -40.71927, -41.50666, -42.28868,
  42.08391, 41.30251, 40.51591, 39.72409, 38.92703, 38.12474, 37.31722, 
    36.50447, 35.68649, 34.86331, 34.03494, 33.20141, 32.36275, 31.519, 
    30.6702, 29.81639, 28.95764, 28.094, 27.22555, 26.35234, 25.47448, 
    24.59204, 23.70512, 22.81381, 21.91823, 21.01848, 20.11469, 19.20699, 
    18.2955, 17.38036, 16.46173, 15.53974, 14.61457, 13.68636, 12.75529, 
    11.82154, 10.88527, 9.946671, 9.005934, 8.063247, 7.118805, 6.172808, 
    5.225454, 4.27695, 3.3275, 2.377314, 1.4266, 0.4755684, -0.4755684, 
    -1.4266, -2.377314, -3.3275, -4.27695, -5.225454, -6.172808, -7.118805, 
    -8.063247, -9.005934, -9.946671, -10.88527, -11.82154, -12.75529, 
    -13.68636, -14.61457, -15.53974, -16.46173, -17.38036, -18.2955, 
    -19.20699, -20.11469, -21.01848, -21.91823, -22.81381, -23.70512, 
    -24.59204, -25.47448, -26.35234, -27.22555, -28.094, -28.95764, 
    -29.81639, -30.6702, -31.519, -32.36275, -33.20141, -34.03494, -34.86331, 
    -35.68649, -36.50447, -37.31722, -38.12474, -38.92703, -39.72409, 
    -40.51591, -41.30251, -42.08391,
  41.87124, 41.09053, 40.30479, 39.51399, 38.71813, 37.9172, 37.11122, 
    36.30017, 35.48409, 34.66297, 33.83684, 33.00574, 32.16968, 31.32872, 
    30.48288, 29.63223, 28.77681, 27.91669, 27.05193, 26.18261, 25.3088, 
    24.43059, 23.54808, 22.66135, 21.77052, 20.87569, 19.97698, 19.07451, 
    18.16841, 17.25882, 16.34587, 15.42971, 14.51049, 13.58837, 12.66351, 
    11.73607, 10.80623, 9.874163, 8.940046, 8.004064, 7.066403, 6.127254, 
    5.186808, 4.245261, 3.30281, 2.359655, 1.415995, 0.472032, -0.472032, 
    -1.415995, -2.359655, -3.30281, -4.245261, -5.186808, -6.127254, 
    -7.066403, -8.004064, -8.940046, -9.874163, -10.80623, -11.73607, 
    -12.66351, -13.58837, -14.51049, -15.42971, -16.34587, -17.25882, 
    -18.16841, -19.07451, -19.97698, -20.87569, -21.77052, -22.66135, 
    -23.54808, -24.43059, -25.3088, -26.18261, -27.05193, -27.91669, 
    -28.77681, -29.63223, -30.48288, -31.32872, -32.16968, -33.00574, 
    -33.83684, -34.66297, -35.48409, -36.30017, -37.11122, -37.9172, 
    -38.71813, -39.51399, -40.30479, -41.09053, -41.87124,
  41.65079, 40.87085, 40.08604, 39.29634, 38.50176, 37.70229, 36.89794, 
    36.08871, 35.27462, 34.45568, 33.63192, 32.80336, 31.97004, 31.132, 
    30.28927, 29.44192, 28.58998, 27.73353, 26.87262, 26.00734, 25.13775, 
    24.26394, 23.386, 22.50403, 21.61812, 20.72838, 19.83493, 18.93789, 
    18.03736, 17.1335, 16.22643, 15.31629, 14.40323, 13.48739, 12.56893, 
    11.64802, 10.72481, 9.799476, 8.872184, 7.943112, 7.012438, 6.080344, 
    5.147013, 4.212631, 3.277388, 2.341473, 1.405076, 0.4683909, -0.4683909, 
    -1.405076, -2.341473, -3.277388, -4.212631, -5.147013, -6.080344, 
    -7.012438, -7.943112, -8.872184, -9.799476, -10.72481, -11.64802, 
    -12.56893, -13.48739, -14.40323, -15.31629, -16.22643, -17.1335, 
    -18.03736, -18.93789, -19.83493, -20.72838, -21.61812, -22.50403, 
    -23.386, -24.26394, -25.13775, -26.00734, -26.87262, -27.73353, 
    -28.58998, -29.44192, -30.28927, -31.132, -31.97004, -32.80336, 
    -33.63192, -34.45568, -35.27462, -36.08871, -36.89794, -37.70229, 
    -38.50176, -39.29634, -40.08604, -40.87085, -41.65079,
  41.42268, 40.64358, 39.85978, 39.07127, 38.27806, 37.48015, 36.67753, 
    35.87022, 35.05824, 34.2416, 33.42032, 32.59444, 31.76398, 30.929, 
    30.08952, 29.2456, 28.3973, 27.54466, 26.68777, 25.82668, 24.96147, 
    24.09223, 23.21904, 22.34199, 21.46118, 20.57672, 19.68871, 18.79726, 
    17.9025, 17.00456, 16.10355, 15.19962, 14.2929, 13.38354, 12.47168, 
    11.55748, 10.6411, 9.722692, 8.802423, 7.880459, 6.956971, 6.032131, 
    5.106114, 4.179099, 3.251263, 2.322789, 1.393856, 0.4646493, -0.4646493, 
    -1.393856, -2.322789, -3.251263, -4.179099, -5.106114, -6.032131, 
    -6.956971, -7.880459, -8.802423, -9.722692, -10.6411, -11.55748, 
    -12.47168, -13.38354, -14.2929, -15.19962, -16.10355, -17.00456, 
    -17.9025, -18.79726, -19.68871, -20.57672, -21.46118, -22.34199, 
    -23.21904, -24.09223, -24.96147, -25.82668, -26.68777, -27.54466, 
    -28.3973, -29.2456, -30.08952, -30.929, -31.76398, -32.59444, -33.42032, 
    -34.2416, -35.05824, -35.87022, -36.67753, -37.48015, -38.27806, 
    -39.07127, -39.85978, -40.64358, -41.42268,
  41.18702, 40.40884, 39.62614, 38.83891, 38.04717, 37.2509, 36.45013, 
    35.64485, 34.83509, 34.02087, 33.2022, 32.37912, 31.55167, 30.71988, 
    29.88379, 29.04346, 28.19893, 27.35027, 26.49753, 25.6408, 24.78014, 
    23.91562, 23.04734, 22.17539, 21.29985, 20.42083, 19.53844, 18.65277, 
    17.76396, 16.87211, 15.97735, 15.07981, 14.17962, 13.27692, 12.37185, 
    11.46456, 10.55519, 9.643898, 8.730841, 7.816175, 6.900063, 5.982669, 
    5.064158, 4.144701, 3.224465, 2.303623, 1.382348, 0.4608116, -0.4608116, 
    -1.382348, -2.303623, -3.224465, -4.144701, -5.064158, -5.982669, 
    -6.900063, -7.816175, -8.730841, -9.643898, -10.55519, -11.46456, 
    -12.37185, -13.27692, -14.17962, -15.07981, -15.97735, -16.87211, 
    -17.76396, -18.65277, -19.53844, -20.42083, -21.29985, -22.17539, 
    -23.04734, -23.91562, -24.78014, -25.6408, -26.49753, -27.35027, 
    -28.19893, -29.04346, -29.88379, -30.71988, -31.55167, -32.37912, 
    -33.2022, -34.02087, -34.83509, -35.64485, -36.45013, -37.2509, 
    -38.04717, -38.83891, -39.62614, -40.40884, -41.18702,
  40.94394, 40.16676, 39.38524, 38.5994, 37.80922, 37.01471, 36.21589, 
    35.41275, 34.60533, 33.79364, 32.97771, 32.15757, 31.33325, 30.50479, 
    29.67224, 28.83563, 27.99503, 27.1505, 26.30208, 25.44986, 24.5939, 
    23.73428, 22.87107, 22.00438, 21.13428, 20.26088, 19.38427, 18.50457, 
    17.62187, 16.73629, 15.84795, 14.95698, 14.0635, 13.16765, 12.26954, 
    11.36934, 10.46716, 9.563174, 8.657512, 7.750327, 6.841775, 5.93201, 
    5.02119, 4.109474, 3.197022, 2.283998, 1.370563, 0.4568816, -0.4568816, 
    -1.370563, -2.283998, -3.197022, -4.109474, -5.02119, -5.93201, 
    -6.841775, -7.750327, -8.657512, -9.563174, -10.46716, -11.36934, 
    -12.26954, -13.16765, -14.0635, -14.95698, -15.84795, -16.73629, 
    -17.62187, -18.50457, -19.38427, -20.26088, -21.13428, -22.00438, 
    -22.87107, -23.73428, -24.5939, -25.44986, -26.30208, -27.1505, 
    -27.99503, -28.83563, -29.67224, -30.50479, -31.33325, -32.15757, 
    -32.97771, -33.79364, -34.60533, -35.41275, -36.21589, -37.01471, 
    -37.80922, -38.5994, -39.38524, -40.16676, -40.94394,
  40.69355, 39.91746, 39.13723, 38.35286, 37.56434, 36.7717, 35.97494, 
    35.17407, 34.36911, 33.56009, 32.74702, 31.92994, 31.10889, 30.28391, 
    29.45502, 28.6223, 27.78577, 26.94551, 26.10157, 25.25401, 24.40292, 
    23.54835, 22.69039, 21.82912, 20.96463, 20.09701, 19.22636, 18.35277, 
    17.47636, 16.59723, 15.71549, 14.83126, 13.94467, 13.05583, 12.16487, 
    11.27192, 10.37712, 9.480604, 8.582511, 7.682984, 6.782168, 5.880208, 
    4.977254, 4.073455, 3.168964, 2.263932, 1.358514, 0.4528638, -0.4528638, 
    -1.358514, -2.263932, -3.168964, -4.073455, -4.977254, -5.880208, 
    -6.782168, -7.682984, -8.582511, -9.480604, -10.37712, -11.27192, 
    -12.16487, -13.05583, -13.94467, -14.83126, -15.71549, -16.59723, 
    -17.47636, -18.35277, -19.22636, -20.09701, -20.96463, -21.82912, 
    -22.69039, -23.54835, -24.40292, -25.25401, -26.10157, -26.94551, 
    -27.78577, -28.6223, -29.45502, -30.28391, -31.10889, -31.92994, 
    -32.74702, -33.56009, -34.36911, -35.17407, -35.97494, -36.7717, 
    -37.56434, -38.35286, -39.13723, -39.91746, -40.69355,
  40.43598, 39.66107, 38.88222, 38.09942, 37.31269, 36.52202, 35.72744, 
    34.92895, 34.12658, 33.32034, 32.51027, 31.6964, 30.87876, 30.05738, 
    29.23232, 28.40361, 27.57131, 26.73548, 25.89616, 25.05343, 24.20735, 
    23.35799, 22.50543, 21.64975, 20.79103, 19.92936, 19.06483, 18.19754, 
    17.32758, 16.45506, 15.58009, 14.70277, 13.82323, 12.94157, 12.05792, 
    11.1724, 10.28514, 9.396269, 8.505915, 7.614214, 6.721301, 5.827315, 
    4.932395, 4.036681, 3.140318, 2.243447, 1.346213, 0.448762, -0.448762, 
    -1.346213, -2.243447, -3.140318, -4.036681, -4.932395, -5.827315, 
    -6.721301, -7.614214, -8.505915, -9.396269, -10.28514, -11.1724, 
    -12.05792, -12.94157, -13.82323, -14.70277, -15.58009, -16.45506, 
    -17.32758, -18.19754, -19.06483, -19.92936, -20.79103, -21.64975, 
    -22.50543, -23.35799, -24.20735, -25.05343, -25.89616, -26.73548, 
    -27.57131, -28.40361, -29.23232, -30.05738, -30.87876, -31.6964, 
    -32.51027, -33.32034, -34.12658, -34.92895, -35.72744, -36.52202, 
    -37.31269, -38.09942, -38.88222, -39.66107, -40.43598,
  40.17135, 39.39772, 38.62035, 37.83924, 37.05439, 36.26581, 35.47353, 
    34.67754, 33.87788, 33.07457, 32.26763, 31.45709, 30.643, 29.82537, 
    29.00427, 28.17974, 27.35181, 26.52055, 25.68602, 24.84826, 24.00736, 
    23.16337, 22.31637, 21.46644, 20.61365, 19.75808, 18.89984, 18.03899, 
    17.17565, 16.30991, 15.44186, 14.57162, 13.69929, 12.82498, 11.9488, 
    11.07087, 10.19132, 9.31025, 8.427797, 7.544083, 6.659235, 5.773382, 
    4.886656, 3.999188, 3.111113, 2.222563, 1.333673, 0.4445804, -0.4445804, 
    -1.333673, -2.222563, -3.111113, -3.999188, -4.886656, -5.773382, 
    -6.659235, -7.544083, -8.427797, -9.31025, -10.19132, -11.07087, 
    -11.9488, -12.82498, -13.69929, -14.57162, -15.44186, -16.30991, 
    -17.17565, -18.03899, -18.89984, -19.75808, -20.61365, -21.46644, 
    -22.31637, -23.16337, -24.00736, -24.84826, -25.68602, -26.52055, 
    -27.35181, -28.17974, -29.00427, -29.82537, -30.643, -31.45709, 
    -32.26763, -33.07457, -33.87788, -34.67754, -35.47353, -36.26581, 
    -37.05439, -37.83924, -38.62035, -39.39772, -40.17135,
  39.89979, 39.12755, 38.35176, 37.57244, 36.78959, 36.00322, 35.21335, 
    34.42, 33.62318, 32.82292, 32.01924, 31.21218, 30.40177, 29.58805, 
    28.77106, 27.95084, 27.12744, 26.30091, 25.4713, 24.63868, 23.8031, 
    22.96464, 22.12335, 21.27932, 20.43262, 19.58332, 18.73152, 17.87728, 
    17.02072, 16.1619, 15.30094, 14.43793, 13.57297, 12.70616, 11.83762, 
    10.96744, 10.09574, 9.222629, 8.34823, 7.472656, 6.596026, 5.718461, 
    4.840082, 3.961012, 3.081377, 2.201299, 1.320906, 0.4403231, -0.4403231, 
    -1.320906, -2.201299, -3.081377, -3.961012, -4.840082, -5.718461, 
    -6.596026, -7.472656, -8.34823, -9.222629, -10.09574, -10.96744, 
    -11.83762, -12.70616, -13.57297, -14.43793, -15.30094, -16.1619, 
    -17.02072, -17.87728, -18.73152, -19.58332, -20.43262, -21.27932, 
    -22.12335, -22.96464, -23.8031, -24.63868, -25.4713, -26.30091, 
    -27.12744, -27.95084, -28.77106, -29.58805, -30.40177, -31.21218, 
    -32.01924, -32.82292, -33.62318, -34.42, -35.21335, -36.00322, -36.78959, 
    -37.57244, -38.35176, -39.12755, -39.89979,
  39.62142, 38.85067, 38.07658, 37.29916, 36.51843, 35.73439, 34.94707, 
    34.15647, 33.36263, 32.56555, 31.76528, 30.96183, 30.15525, 29.34557, 
    28.53283, 27.71707, 26.89834, 26.07669, 25.25217, 24.42483, 23.59474, 
    22.76195, 21.92654, 21.08856, 20.2481, 19.40522, 18.56001, 17.71254, 
    16.8629, 16.01117, 15.15745, 14.30182, 13.44438, 12.58523, 11.72446, 
    10.86218, 9.998483, 9.133484, 8.267286, 7.4, 6.531734, 5.662601, 
    4.792715, 3.922188, 3.051136, 2.179676, 1.307923, 0.4359938, -0.4359938, 
    -1.307923, -2.179676, -3.051136, -3.922188, -4.792715, -5.662601, 
    -6.531734, -7.4, -8.267286, -9.133484, -9.998483, -10.86218, -11.72446, 
    -12.58523, -13.44438, -14.30182, -15.15745, -16.01117, -16.8629, 
    -17.71254, -18.56001, -19.40522, -20.2481, -21.08856, -21.92654, 
    -22.76195, -23.59474, -24.42483, -25.25217, -26.07669, -26.89834, 
    -27.71707, -28.53283, -29.34557, -30.15525, -30.96183, -31.76528, 
    -32.56555, -33.36263, -34.15647, -34.94707, -35.73439, -36.51843, 
    -37.29916, -38.07658, -38.85067, -39.62142,
  39.33637, 38.56721, 37.79493, 37.01954, 36.24105, 35.45947, 34.67482, 
    33.88711, 33.09637, 32.30262, 31.50589, 30.7062, 29.90359, 29.0981, 
    28.28975, 27.47861, 26.6647, 25.84807, 25.02878, 24.20688, 23.38242, 
    22.55546, 21.72607, 20.8943, 20.06023, 19.22392, 18.38545, 17.5449, 
    16.70233, 15.85784, 15.0115, 14.1634, 13.31363, 12.46228, 11.60943, 
    10.75519, 9.899641, 9.042892, 8.185037, 7.326178, 6.466415, 5.605854, 
    4.744597, 3.88275, 3.02042, 2.157712, 1.294735, 0.4315965, -0.4315965, 
    -1.294735, -2.157712, -3.02042, -3.88275, -4.744597, -5.605854, 
    -6.466415, -7.326178, -8.185037, -9.042892, -9.899641, -10.75519, 
    -11.60943, -12.46228, -13.31363, -14.1634, -15.0115, -15.85784, 
    -16.70233, -17.5449, -18.38545, -19.22392, -20.06023, -20.8943, 
    -21.72607, -22.55546, -23.38242, -24.20688, -25.02878, -25.84807, 
    -26.6647, -27.47861, -28.28975, -29.0981, -29.90359, -30.7062, -31.50589, 
    -32.30262, -33.09637, -33.88711, -34.67482, -35.45947, -36.24105, 
    -37.01954, -37.79493, -38.56721, -39.33637,
  39.04476, 38.27731, 37.50697, 36.73372, 35.9576, 35.1786, 34.39675, 
    33.61207, 32.82457, 32.03428, 31.24123, 30.44544, 29.64695, 28.84579, 
    28.04199, 27.2356, 26.42666, 25.61521, 24.8013, 23.98498, 23.1663, 
    22.34532, 21.52209, 20.69669, 19.86915, 19.03956, 18.20799, 17.37449, 
    16.53915, 15.70203, 14.86322, 14.02279, 13.18083, 12.33741, 11.49262, 
    10.64656, 9.799295, 8.95093, 8.101551, 7.251252, 6.400125, 5.548265, 
    4.695769, 3.842732, 2.989253, 2.135427, 1.281355, 0.4271349, -0.4271349, 
    -1.281355, -2.135427, -2.989253, -3.842732, -4.695769, -5.548265, 
    -6.400125, -7.251252, -8.101551, -8.95093, -9.799295, -10.64656, 
    -11.49262, -12.33741, -13.18083, -14.02279, -14.86322, -15.70203, 
    -16.53915, -17.37449, -18.20799, -19.03956, -19.86915, -20.69669, 
    -21.52209, -22.34532, -23.1663, -23.98498, -24.8013, -25.61521, 
    -26.42666, -27.2356, -28.04199, -28.84579, -29.64695, -30.44544, 
    -31.24123, -32.03428, -32.82457, -33.61207, -34.39675, -35.1786, 
    -35.9576, -36.73372, -37.50697, -38.27731, -39.04476,
  38.74672, 37.9811, 37.21281, 36.44184, 35.66821, 34.89193, 34.11302, 
    33.33149, 32.54737, 31.76069, 30.97146, 30.17971, 29.38548, 28.5888, 
    27.78969, 26.98821, 26.18438, 25.37826, 24.56988, 23.75929, 22.94654, 
    22.13168, 21.31477, 20.49586, 19.67501, 18.85229, 18.02774, 17.20144, 
    16.37346, 15.54386, 14.71272, 13.88009, 13.04607, 12.21073, 11.37413, 
    10.53637, 9.697527, 8.857674, 8.016898, 7.175284, 6.332918, 5.489884, 
    4.646272, 3.802168, 2.957661, 2.112839, 1.267794, 0.4226128, -0.4226128, 
    -1.267794, -2.112839, -2.957661, -3.802168, -4.646272, -5.489884, 
    -6.332918, -7.175284, -8.016898, -8.857674, -9.697527, -10.53637, 
    -11.37413, -12.21073, -13.04607, -13.88009, -14.71272, -15.54386, 
    -16.37346, -17.20144, -18.02774, -18.85229, -19.67501, -20.49586, 
    -21.31477, -22.13168, -22.94654, -23.75929, -24.56988, -25.37826, 
    -26.18438, -26.98821, -27.78969, -28.5888, -29.38548, -30.17971, 
    -30.97146, -31.76069, -32.54737, -33.33149, -34.11302, -34.89193, 
    -35.66821, -36.44184, -37.21281, -37.9811, -38.74672,
  38.44237, 37.67871, 36.91259, 36.14403, 35.37302, 34.59959, 33.82376, 
    33.04553, 32.26494, 31.482, 30.69673, 29.90917, 29.11935, 28.32729, 
    27.53302, 26.73659, 25.93803, 25.13737, 24.33467, 23.52995, 22.72328, 
    21.91469, 21.10424, 20.29198, 19.47795, 18.66223, 17.84485, 17.02589, 
    16.20541, 15.38346, 14.56011, 13.73542, 12.90947, 12.08233, 11.25405, 
    10.42472, 9.594414, 8.763195, 7.931143, 7.098334, 6.264847, 5.430757, 
    4.596145, 3.761089, 2.925669, 2.089966, 1.254061, 0.4180338, -0.4180338, 
    -1.254061, -2.089966, -2.925669, -3.761089, -4.596145, -5.430757, 
    -6.264847, -7.098334, -7.931143, -8.763195, -9.594414, -10.42472, 
    -11.25405, -12.08233, -12.90947, -13.73542, -14.56011, -15.38346, 
    -16.20541, -17.02589, -17.84485, -18.66223, -19.47795, -20.29198, 
    -21.10424, -21.91469, -22.72328, -23.52995, -24.33467, -25.13737, 
    -25.93803, -26.73659, -27.53302, -28.32729, -29.11935, -29.90917, 
    -30.69673, -31.482, -32.26494, -33.04553, -33.82376, -34.59959, 
    -35.37302, -36.14403, -36.91259, -37.67871, -38.44237,
  38.13184, 37.37026, 36.60646, 35.84042, 35.07218, 34.30174, 33.52912, 
    32.75434, 31.97741, 31.19835, 30.4172, 29.63398, 28.84871, 28.06141, 
    27.27213, 26.4809, 25.68774, 24.89271, 24.09582, 23.29713, 22.49667, 
    21.6945, 20.89065, 20.08517, 19.2781, 18.46952, 17.65945, 16.84796, 
    16.0351, 15.22093, 14.4055, 13.58888, 12.77113, 11.9523, 11.13247, 
    10.31169, 9.490034, 8.667565, 7.844352, 7.020462, 6.195964, 5.370928, 
    4.545426, 3.719527, 2.893303, 2.066826, 1.240168, 0.4134014, -0.4134014, 
    -1.240168, -2.066826, -2.893303, -3.719527, -4.545426, -5.370928, 
    -6.195964, -7.020462, -7.844352, -8.667565, -9.490034, -10.31169, 
    -11.13247, -11.9523, -12.77113, -13.58888, -14.4055, -15.22093, -16.0351, 
    -16.84796, -17.65945, -18.46952, -19.2781, -20.08517, -20.89065, 
    -21.6945, -22.49667, -23.29713, -24.09582, -24.89271, -25.68774, 
    -26.4809, -27.27213, -28.06141, -28.84871, -29.63398, -30.4172, 
    -31.19835, -31.97741, -32.75434, -33.52912, -34.30174, -35.07218, 
    -35.84042, -36.60646, -37.37026, -38.13184,
  37.81525, 37.05589, 36.29453, 35.53117, 34.76583, 33.99852, 33.22925, 
    32.45805, 31.68493, 30.90992, 30.13302, 29.35428, 28.5737, 27.79133, 
    27.00718, 26.22129, 25.43369, 24.64441, 23.85349, 23.06096, 22.26687, 
    21.47124, 20.67413, 19.87557, 19.07561, 18.27429, 17.47165, 16.66776, 
    15.86266, 15.05639, 14.24901, 13.44058, 12.63114, 11.82075, 11.00947, 
    10.19736, 9.384465, 8.570855, 7.756588, 6.941722, 6.12632, 5.310442, 
    4.494153, 3.677513, 2.860586, 2.043435, 1.226125, 0.4087191, -0.4087191, 
    -1.226125, -2.043435, -2.860586, -3.677513, -4.494153, -5.310442, 
    -6.12632, -6.941722, -7.756588, -8.570855, -9.384465, -10.19736, 
    -11.00947, -11.82075, -12.63114, -13.44058, -14.24901, -15.05639, 
    -15.86266, -16.66776, -17.47165, -18.27429, -19.07561, -19.87557, 
    -20.67413, -21.47124, -22.26687, -23.06096, -23.85349, -24.64441, 
    -25.43369, -26.22129, -27.00718, -27.79133, -28.5737, -29.35428, 
    -30.13302, -30.90992, -31.68493, -32.45805, -33.22925, -33.99852, 
    -34.76583, -35.53117, -36.29453, -37.05589, -37.81525,
  37.49273, 36.73572, 35.97694, 35.2164, 34.4541, 33.69006, 32.9243, 
    32.15683, 31.38766, 30.61683, 29.84434, 29.07022, 28.29449, 27.51719, 
    26.73832, 25.95792, 25.17602, 24.39264, 23.60783, 22.8216, 22.034, 
    21.24507, 20.45482, 19.66332, 18.87058, 18.07666, 17.2816, 16.48543, 
    15.6882, 14.88996, 14.09074, 13.29061, 12.4896, 11.68776, 10.88514, 
    10.0818, 9.277779, 8.473132, 7.667912, 6.862171, 6.055964, 5.249342, 
    4.442361, 3.635076, 2.827541, 2.019811, 1.211942, 0.40399, -0.40399, 
    -1.211942, -2.019811, -2.827541, -3.635076, -4.442361, -5.249342, 
    -6.055964, -6.862171, -7.667912, -8.473132, -9.277779, -10.0818, 
    -10.88514, -11.68776, -12.4896, -13.29061, -14.09074, -14.88996, 
    -15.6882, -16.48543, -17.2816, -18.07666, -18.87058, -19.66332, 
    -20.45482, -21.24507, -22.034, -22.8216, -23.60783, -24.39264, -25.17602, 
    -25.95792, -26.73832, -27.51719, -28.29449, -29.07022, -29.84434, 
    -30.61683, -31.38766, -32.15683, -32.9243, -33.69006, -34.4541, -35.2164, 
    -35.97694, -36.73572, -37.49273,
  37.1644, 36.40988, 35.65382, 34.89624, 34.13713, 33.37651, 32.6144, 
    31.8508, 31.08575, 30.31924, 29.55131, 28.78197, 28.01123, 27.23913, 
    26.46569, 25.69092, 24.91487, 24.13754, 23.35897, 22.57919, 21.79822, 
    21.01611, 20.23287, 19.44855, 18.66317, 17.87678, 17.0894, 16.30107, 
    15.51184, 14.72173, 13.9308, 13.13908, 12.3466, 11.55342, 10.75957, 
    9.965097, 9.170046, 8.37446, 7.578384, 6.781863, 5.984942, 5.187668, 
    4.390087, 3.592245, 2.79419, 1.995969, 1.197629, 0.3992176, -0.3992176, 
    -1.197629, -1.995969, -2.79419, -3.592245, -4.390087, -5.187668, 
    -5.984942, -6.781863, -7.578384, -8.37446, -9.170046, -9.965097, 
    -10.75957, -11.55342, -12.3466, -13.13908, -13.9308, -14.72173, 
    -15.51184, -16.30107, -17.0894, -17.87678, -18.66317, -19.44855, 
    -20.23287, -21.01611, -21.79822, -22.57919, -23.35897, -24.13754, 
    -24.91487, -25.69092, -26.46569, -27.23913, -28.01123, -28.78197, 
    -29.55131, -30.31924, -31.08575, -31.8508, -32.6144, -33.37651, 
    -34.13713, -34.89624, -35.65382, -36.40988, -37.1644,
  36.83038, 36.0785, 35.32531, 34.57083, 33.81506, 33.05801, 32.29969, 
    31.54013, 30.77932, 30.0173, 29.25407, 28.48965, 27.72406, 26.95732, 
    26.18944, 25.42046, 24.65038, 23.87924, 23.10706, 22.33386, 21.55966, 
    20.7845, 20.0084, 19.23139, 18.45349, 17.67474, 16.89517, 16.11481, 
    15.33368, 14.55183, 13.76928, 12.98607, 12.20224, 11.41781, 10.63283, 
    9.847324, 9.061338, 8.274905, 7.488063, 6.70085, 5.913303, 5.125462, 
    4.337364, 3.549049, 2.760556, 1.971925, 1.183195, 0.3944048, -0.3944048, 
    -1.183195, -1.971925, -2.760556, -3.549049, -4.337364, -5.125462, 
    -5.913303, -6.70085, -7.488063, -8.274905, -9.061338, -9.847324, 
    -10.63283, -11.41781, -12.20224, -12.98607, -13.76928, -14.55183, 
    -15.33368, -16.11481, -16.89517, -17.67474, -18.45349, -19.23139, 
    -20.0084, -20.7845, -21.55966, -22.33386, -23.10706, -23.87924, 
    -24.65038, -25.42046, -26.18944, -26.95732, -27.72406, -28.48965, 
    -29.25407, -30.0173, -30.77932, -31.54013, -32.29969, -33.05801, 
    -33.81506, -34.57083, -35.32531, -36.0785, -36.83038,
  36.4908, 35.7417, 34.99154, 34.2403, 33.48802, 32.73469, 31.98032, 
    31.22494, 30.46854, 29.71115, 28.95277, 28.19342, 27.43312, 26.67189, 
    25.90973, 25.14667, 24.38272, 23.6179, 22.85224, 22.08575, 21.31846, 
    20.55038, 19.78154, 19.01196, 18.24167, 17.47068, 16.69903, 15.92674, 
    15.15383, 14.38034, 13.60628, 12.83169, 12.05659, 11.28102, 10.505, 
    9.728554, 8.951721, 8.174527, 7.397004, 6.619181, 5.84109, 5.06276, 
    4.284225, 3.505514, 2.72666, 1.947694, 1.168648, 0.3895547, -0.3895547, 
    -1.168648, -1.947694, -2.72666, -3.505514, -4.284225, -5.06276, -5.84109, 
    -6.619181, -7.397004, -8.174527, -8.951721, -9.728554, -10.505, 
    -11.28102, -12.05659, -12.83169, -13.60628, -14.38034, -15.15383, 
    -15.92674, -16.69903, -17.47068, -18.24167, -19.01196, -19.78154, 
    -20.55038, -21.31846, -22.08575, -22.85224, -23.6179, -24.38272, 
    -25.14667, -25.90973, -26.67189, -27.43312, -28.19342, -28.95277, 
    -29.71115, -30.46854, -31.22494, -31.98032, -32.73469, -33.48802, 
    -34.2403, -34.99154, -35.7417, -36.4908,
  36.14578, 35.39962, 34.65261, 33.90479, 33.15614, 32.40669, 31.65643, 
    30.90537, 30.15354, 29.40093, 28.64755, 27.89343, 27.13857, 26.38298, 
    25.62668, 24.86968, 24.112, 23.35365, 22.59464, 21.835, 21.07474, 
    20.31387, 19.55242, 18.79039, 18.02782, 17.26471, 16.50109, 15.73699, 
    14.9724, 14.20737, 13.4419, 12.67602, 11.90976, 11.14313, 10.37615, 
    9.608856, 8.84126, 8.073387, 7.305261, 6.536906, 5.768345, 4.999602, 
    4.230701, 3.461666, 2.692521, 1.92329, 1.153999, 0.3846703, -0.3846703, 
    -1.153999, -1.92329, -2.692521, -3.461666, -4.230701, -4.999602, 
    -5.768345, -6.536906, -7.305261, -8.073387, -8.84126, -9.608856, 
    -10.37615, -11.14313, -11.90976, -12.67602, -13.4419, -14.20737, 
    -14.9724, -15.73699, -16.50109, -17.26471, -18.02782, -18.79039, 
    -19.55242, -20.31387, -21.07474, -21.835, -22.59464, -23.35365, -24.112, 
    -24.86968, -25.62668, -26.38298, -27.13857, -27.89343, -28.64755, 
    -29.40093, -30.15354, -30.90537, -31.65643, -32.40669, -33.15614, 
    -33.90479, -34.65261, -35.39962, -36.14578,
  35.79544, 35.05236, 34.30869, 33.56442, 32.81957, 32.07414, 31.32814, 
    30.58158, 29.83445, 29.08677, 28.33856, 27.58981, 26.84053, 26.09074, 
    25.34044, 24.58965, 23.83837, 23.08662, 22.33441, 21.58174, 20.82863, 
    20.0751, 19.32115, 18.5668, 17.81206, 17.05695, 16.30147, 15.54564, 
    14.78949, 14.03301, 13.27623, 12.51916, 11.76182, 11.00421, 10.24637, 
    9.488298, 8.730017, 7.971541, 7.212887, 6.454072, 5.695111, 4.936023, 
    4.176824, 3.41753, 2.658159, 1.898728, 1.139254, 0.3797542, -0.3797542, 
    -1.139254, -1.898728, -2.658159, -3.41753, -4.176824, -4.936023, 
    -5.695111, -6.454072, -7.212887, -7.971541, -8.730017, -9.488298, 
    -10.24637, -11.00421, -11.76182, -12.51916, -13.27623, -14.03301, 
    -14.78949, -15.54564, -16.30147, -17.05695, -17.81206, -18.5668, 
    -19.32115, -20.0751, -20.82863, -21.58174, -22.33441, -23.08662, 
    -23.83837, -24.58965, -25.34044, -26.09074, -26.84053, -27.58981, 
    -28.33856, -29.08677, -29.83445, -30.58158, -31.32814, -32.07414, 
    -32.81957, -33.56442, -34.30869, -35.05236, -35.79544,
  35.43988, 34.70005, 33.95987, 33.21932, 32.47842, 31.73718, 30.9956, 
    30.25368, 29.51142, 28.76883, 28.02592, 27.28269, 26.53915, 25.7953, 
    25.05115, 24.3067, 23.56197, 22.81695, 22.07165, 21.32609, 20.58027, 
    19.83419, 19.08786, 18.3413, 17.59451, 16.84749, 16.10026, 15.35282, 
    14.60518, 13.85736, 13.10935, 12.36118, 11.61284, 10.86435, 10.11571, 
    9.366945, 8.618052, 7.869044, 7.119931, 6.370722, 5.621428, 4.872057, 
    4.122622, 3.37313, 2.623593, 1.87402, 1.124422, 0.3748092, -0.3748092, 
    -1.124422, -1.87402, -2.623593, -3.37313, -4.122622, -4.872057, 
    -5.621428, -6.370722, -7.119931, -7.869044, -8.618052, -9.366945, 
    -10.11571, -10.86435, -11.61284, -12.36118, -13.10935, -13.85736, 
    -14.60518, -15.35282, -16.10026, -16.84749, -17.59451, -18.3413, 
    -19.08786, -19.83419, -20.58027, -21.32609, -22.07165, -22.81695, 
    -23.56197, -24.3067, -25.05115, -25.7953, -26.53915, -27.28269, 
    -28.02592, -28.76883, -29.51142, -30.25368, -30.9956, -31.73718, 
    -32.47842, -33.21932, -33.95987, -34.70005, -35.43988,
  35.07925, 34.34282, 33.60628, 32.86962, 32.13284, 31.39594, 30.65893, 
    29.92181, 29.18457, 28.44723, 27.70978, 26.97222, 26.23456, 25.4968, 
    24.75893, 24.02097, 23.28291, 22.54476, 21.80651, 21.06818, 20.32976, 
    19.59126, 18.85267, 18.114, 17.37526, 16.63645, 15.89756, 15.15861, 
    14.41959, 13.6805, 12.94136, 12.20216, 11.46291, 10.72361, 9.984256, 
    9.244861, 8.505425, 7.765951, 7.026442, 6.286901, 5.547333, 4.807739, 
    4.068124, 3.32849, 2.588841, 1.849181, 1.109512, 0.3698378, -0.3698378, 
    -1.109512, -1.849181, -2.588841, -3.32849, -4.068124, -4.807739, 
    -5.547333, -6.286901, -7.026442, -7.765951, -8.505425, -9.244861, 
    -9.984256, -10.72361, -11.46291, -12.20216, -12.94136, -13.6805, 
    -14.41959, -15.15861, -15.89756, -16.63645, -17.37526, -18.114, 
    -18.85267, -19.59126, -20.32976, -21.06818, -21.80651, -22.54476, 
    -23.28291, -24.02097, -24.75893, -25.4968, -26.23456, -26.97222, 
    -27.70978, -28.44723, -29.18457, -29.92181, -30.65893, -31.39594, 
    -32.13284, -32.86962, -33.60628, -34.34282, -35.07925 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.500448, 0.6373758, 0.3299181, 0.2709744, 0.3045332, 
    0.9904844, 1, 0.7193916, 0.6372474, 0.08596428, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2001312, 0.4111539, 0, 0, 0, 0, 0, 0, 
    0.3257935, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9846206, 0.1322953, 0, 0, 0,
  0.4213375, 0.7249894, 0.1194391, 0.4090452, 0.0004055478, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1275371, 0.2101071, 0.501195, 0.907451, 0.5348656, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.2795206, 0, 0, 0, 0, 0, 0, 0.4748606, 0.08597825, 0, 
    0, 0, 0, 0, 0.3374754, 0.9515835, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.974499, 0.2595553, 0, 0, 0, 0,
  1, 1, 0.5694539, 0.2257697, 0.07591473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1566211, 0, 0, 0, 0.3620377, 0, 0, 0, 0, 0, 0, 
    0.2321739, 0, 0, 0, 0, 0, 0, 0.6652638, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6224186, 0, 0, 0, 0, 0,
  1, 1, 0.5671622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0328016, 0.3505093, 0.800697, 0.4199587, 0.3645951, 0.2070305, 
    0.1039276, 0.04041792, 0.1039293, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3621618, 0.9914034, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9980344, 0.1799124, 0, 0, 0, 0, 0,
  1, 1, 0.6025393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0554254, 0.07674838, 0.3268177, 0.2018002, 0, 0, 0, 0.2147634, 
    0.246665, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1000221, 0.9995502, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9989821, 
    0.4096552, 0, 0, 0, 0, 0, 0,
  0.628101, 0.6280472, 0.4677134, 0, 0, 0.3171421, 0.0938872, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2612283, 0.06390974, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3284912, 0.3768882, 0.8638445, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7643126, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.05901703, 0.9235198, 0.8531228, 0.7637583, 0.2779488, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0508899, 0.05089059, 0.3887566, 
    0.2545041, 0.2612266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4230824, 0.09009741, 
    0.4622726, 0.9831397, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.3566395, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.3848666, 0.9172006, 1, 1, 0.8194785, 0.02148438, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1404992, 0.4942557, 0, 0, 0.1406009, 0, 
    0, 0, 0, 0.2166595, 0, 0, 0, 0.02490224, 0.9627016, 0.8158007, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9282088, 
    0.03051941, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.5683897, 0.9379957, 0.6364555, 0.2024043, 0.03349722, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.320924, 0.9845472, 0.2649983, 
    0.1140551, 0, 0, 0, 0, 0, 0.01618783, 0, 0, 0, 0.08289424, 0.1259722, 
    0.8170571, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7655389, 0.005966454, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0272528, 0.8907499, 0.9876926, 0.7710279, 0.1670542, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4784564, 1, 0.6486406, 0.6920749, 
    0.2536378, 0, 0, 0, 0, 0, 0, 0, 0, 0.2509409, 0.8028153, 0.9793605, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7416639, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.648589, 1, 0.9992579, 0.2293907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.09293438, 0.9501851, 0.8690677, 1, 0.5762319, 0, 
    0, 0.008900359, 0.003358786, 0, 0, 0, 0, 0.0356602, 0.9891973, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3823546, 
    0.00315241, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.4935699, 1, 0.7489711, 0.1704132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1722069, 0.2898026, 1, 0.8352928, 0.0001595881, 
    0.2050383, 0.6669478, 0.1472481, 0, 0, 0, 0, 0, 0.7378939, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3177179, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.3381471, 0.9340628, 0.9308964, 0.34702, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0710042, 0.01311141, 0.01958092, 0.2182962, 
    0.9644061, 0.2152033, 0.07139239, 0.07196605, 0, 0, 0, 0, 0, 0, 
    0.8858101, 1, 0.933995, 0.8029567, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8098463, 0.2802811, 0.06792729, 0, 0, 0, 0, 0,
  0, 0, 0, 0.062082, 0.4496638, 0.9014636, 1, 0.6371259, 0.0002500278, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07396818, 0.06363945, 0.2273634, 
    0.7217154, 1, 0.4123627, 0, 0, 0, 0, 0, 0, 0, 0.03488547, 0.9638747, 
    0.4518672, 0.2722468, 0.101736, 0.9105512, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8664908, 0.293852, 0.1126182, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0.1481497, 0.8071872, 1, 0.9563567, 0.1187265, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09094947, 0.8744214, 1, 1, 0.6151962, 
    7.862093e-05, 0, 0, 0, 0, 0, 0, 0.05432393, 0.3167762, 0, 0.1943092, 0, 
    0.6416867, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9944282, 0.1187612, 0.2975091, 0.5171648, 0, 0, 0, 0, 0,
  0, 0, 0, 0.006354006, 0.888454, 1, 1, 0.1866042, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2678939, 1, 1, 1, 0.9953833, 0.4038017, 0, 
    0.1863101, 0.1370078, 0, 0, 0, 0, 0, 0, 0, 0, 0.1708246, 0.9664814, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.643471, 
    0.3777492, 0.3611507, 0, 0, 0, 0, 0,
  0, 0, 0, 0.2080797, 0.9673514, 1, 0.8374537, 0.04476063, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01296526, 0.7596481, 1, 1, 1, 
    0.9865646, 0.8895645, 0.9378822, 0.2410906, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01894641, 0.7163382, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9017419, 0.4822293, 0.01936743, 0, 0, 0, 0, 0,
  0.2283506, 0.2283831, 0.3606219, 0.8600088, 1, 1, 0.8187755, 0.09858553, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3482806, 1, 1, 1, 1, 
    1, 1, 0.2386805, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04633646, 0.8615492, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.850582, 0.348906, 
    0.139303, 0, 0, 0, 0,
  0.9058077, 1, 1, 0.9630018, 0.8670257, 0.6587394, 0.3201251, 0.1648381, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1173386, 1, 1, 1, 1, 
    1, 1, 0.7136791, 0.01745822, 0, 0, 0, 0, 0, 0, 0, 0.0606117, 0.3882409, 
    0.9743452, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.784731, 0.03699823, 0, 0, 0,
  0.4231035, 0.9422162, 0.9297223, 0.3348973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01853104, 0.8556062, 1, 1, 1, 1, 1, 
    1, 0.08117965, 0.02060091, 0.04679306, 0.4853819, 0.590209, 0.5901864, 
    0.5901626, 0.5901374, 0.7937525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9957187, 0.1070087, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.5207784, 1, 1, 1, 1, 1, 0.9874919, 0.008527548, 0.2921969, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9391072, 0.1130477, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1617553, 0.9999905, 1, 1, 1, 0.92387, 0.5260675, 0, 0.004612686, 
    0.03066925, 0.3373398, 0.5646344, 0.7950864, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9652795, 
    0.03719426, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01460301, 0.8115592, 1, 1, 1, 0.1636489, 0, 0, 0, 0, 0, 0, 
    0.6152393, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8714985, 0.2261804, 0, 0, 0.3437575, 0.01257803,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2064631, 0.733834, 1, 1, 0.3149392, 0, 0, 0, 0, 0, 0, 
    0.2648452, 0.6866553, 0.7366514, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9174272, 0.1166509, 0, 0.05494488, 
    0.9094183, 0.8397222,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.07105455, 0, 0, 0.1277506, 0.9753432, 1, 0.6722792, 0.08202832, 0, 
    0, 0, 0, 0, 0, 0, 0.04108687, 0.2125929, 0.6796362, 0.8867523, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4437395, 0, 
    0.003395685, 0.9062591, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.06928185, 0, 0, 0, 0.6190757, 0.4693122, 0.9500455, 0.8051443, 
    0.06908886, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5560373, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9714394, 0.4920565, 0.007317367, 0, 
    0.1679957, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1870881, 0.1032061, 0, 0.3068611, 0.901248, 0.525517, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.08475742, 0.9234713, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7293079, 0, 0, 0.4481606, 0.3670389, 
    0.8051461, 0.3047968,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2969156, 0.1804042, 0, 0, 0.6011499, 0.5948403, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3606173, 0.8423501, 0.9566985, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9882501, 0.4393826, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1341057, 0, 0, 0.3335736, 0.2354348, 0, 0, 0.225836, 0.4429893, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7404009, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9729695, 0.7830737, 0.3542824, 0.3088061, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.08371773, 0.6231546, 0.07811955, 0, 0, 0.1299088, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1582873, 0.6573294, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9011589, 0.4768529, 0.2806725, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.4617452, 0.2357396, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.05252013, 0.5075252, 0.9784946, 1, 1, 1, 1, 1, 1, 
    0.9491259, 0.6694556, 0.0476924, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2044773, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1850218, 0.3838319, 0.3948988, 0.6347017, 0.897539, 0.8975486, 
    0.625631, 0.3950224, 0.1931382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.04801759, 0.008659004, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2955928, 0.4134034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2288118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1252723, 0.02888734, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1657154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1331506, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2602637, 
    0.1827536, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.308817, 
    0.1388956, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009059105, 
    0.04102035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1710694,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1561902, 
    0.9037677,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7994146, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02431367, 
    0.5217998, 1, 0.9833409,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03587419, 0.3440025, 
    0.8423416, 1, 0.9747218, 0.3018562,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001283266, 0.05145107, 0, 0, 0, 0, 0, 
    0.4153767, 0.9991337, 1, 0.9749234, 0.6001224, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001449973, 0.7731972, 0.1336049, 0, 0, 
    0.1802618, 0.1813705, 0, 0.8987046, 0.7961607, 0.290663, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3244956, 0.5728012, 0.6642565, 
    0.6642635, 0.7536004, 0.7371183, 0.09692896, 0.2581114, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01432, 0.7955128, 1, 1, 1, 
    0.8594135, 0.4985357, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008547029, 0.6526902, 0.9749812, 
    0.7542722, 0.4022479, 0.04722129, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3207461, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8175688, 0.8197373, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3270165, 0.08929753, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1860417, 
    0.1124855, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2794361, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1755751,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05289424,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2801953, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004320362, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2700683, 0.1831646, 0.1345469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5860988, 0.2863249, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 orog =
  0.05263353, 0.9425675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.210776, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.252779, 74.21071, 95.69428, 
    40.84037, 37.33909, 173.0547, 413.3694, 558.9451, 332.2694, 351.5737, 
    71.52609, 0.03417388, 1.300127, 17.79588, 8.458535, 18.73478, 17.63159, 
    0, 0, 0, 24.16101, 0, 0, 0, 0, 0, 0, 0, 1.372658, 299.2773, 291.463, 0, 
    0, 0, 0, 0, 0.0248737, 34.27986, 188.9342, 329.4237, 350.9251, 251.6835, 
    165.8015, 165.6417, 201.2802, 268.5535, 314.2737, 338.9506, 356.3144, 
    377.6248, 410.6694, 439.9049, 453.2951, 445.0014, 438.5307, 407.9247, 
    339.9653, 265.3149, 224.8092, 190.4008, 158.7892, 103.6094, 19.02374, 0, 
    0, 0,
  9.158454, 18.90683, 3.012916, 53.90588, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2984579, 4.255527, 
    84.79544, 147.7691, 233.7292, 347.7168, 36.84171, 0, 0, 0, 0, 0, 0, 
    0.4999831, 0, 0, 0, 25.2615, 9.891716, 381.2982, 0.7240577, 0, 0, 0, 0, 
    147.3826, 251.5665, 17.10577, 0, 0, 0, 0, 0, 12.48063, 173.854, 367.2847, 
    472.174, 458.6521, 325.3309, 227.1559, 236.9397, 249.4832, 296.6798, 
    348.9885, 370.6396, 368.1631, 393.7355, 411.4686, 451.679, 461.741, 
    457.9003, 439.6093, 391.6231, 291.6416, 227.3665, 205.8765, 180.0435, 
    108.2699, 20.55778, 0, 0, 0, 0,
  146.5898, 178.415, 28.03686, 31.16747, 0, 0, 0, 0, 0, 0, 0, 0, 0.03837012, 
    1.052421, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.03251622, 0.6342183, 0, 0.003365346, 0.1732605, 15.05509, 
    0.627657, 0, 0, 5.064898, 0.5615213, 22.54741, 2.144348, 0, 0, 255.0734, 
    8.867086, 0, 0, 0.008958309, 1.017161, 28.21741, 115.5201, 0, 0, 0, 0, 0, 
    0, 66.54465, 223.7023, 341.7935, 467.8122, 479.3343, 405.95, 344.1333, 
    317.8734, 316.412, 353.7882, 397.7623, 399.601, 410.1562, 420.6944, 
    456.795, 491.1674, 486.9185, 461.8076, 437.4255, 366.8581, 265.5489, 
    220.6245, 207.5233, 145.059, 52.48993, 0.02635965, 0, 0, 0, 0,
  312.5654, 332.0361, 48.98602, 0.01820307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2560336, 10.64937, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6525263, 85.40112, 154.1216, 
    145.2693, 104.7963, 68.44398, 59.66086, 5.658707, 51.90486, 0, 
    0.0002234011, 0.002236324, 0, 4.058273, 2.615149, 0, 0, 0, 0, 0, 0, 0, 
    45.61565, 143.503, 253.2654, 347.6613, 440.0746, 419.2403, 373.5648, 
    356.8692, 343.2001, 372.7208, 395.3455, 415.5849, 430.8153, 461.9744, 
    506.336, 526.5826, 478.6951, 428.0603, 393.4123, 322.4732, 237.9073, 
    211.1528, 175.5259, 95.53486, 5.59942, 0, 0, 0, 0, 0,
  277.1137, 216.7668, 65.78798, 0.01913495, 0, 6.423023, 0.05600383, 0, 0, 0, 
    0.008824782, 0.03805306, 5.421787, 6.542611, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.47252, 
    50.65664, 159.9921, 46.69725, 1.587591, 2.254171, 0.6875598, 155.2946, 
    109.7841, 0, 0, 0, 0, 6.335535, 1.460464, 0, 0, 0, 0, 0, 0, 0, 
    0.001764559, 51.18093, 107.6214, 220.6243, 313.7549, 357.301, 394.333, 
    380.0004, 369.1454, 378.0013, 370.4623, 409.9088, 457.2517, 510.6886, 
    598.5809, 591.0898, 488.7568, 418.8461, 368.6212, 287.8756, 211.7777, 
    183.3996, 128.3429, 26.55859, 0, 0, 0, 0, 0, 0,
  212.3771, 135.9476, 49.42075, 12.49728, 1.597956, 29.35641, 0.7934011, 
    2.107809, 0.008830293, 0.1460706, 1.322528, 19.1708, 1.042597, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1036084, 1.6234, 0.4369082, 1.249874, 151.7508, 
    165.1876, 0.1203202, 0, 0, 0.966633, 12.21299, 9.954236, 0, 0, 0, 0, 0, 
    0, 3.324982, 15.32631, 53.0812, 144.7708, 241.6709, 340.8276, 409.1607, 
    415.9962, 398.8717, 383.6034, 399.2011, 408.1645, 448.2938, 490.6762, 
    554.4016, 678.0546, 651.3043, 520.1175, 420.8705, 346.4621, 250.8538, 
    183.0857, 142.4498, 71.22203, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.2228342, 92.88892, 92.60233, 105.3637, 26.52375, 48.40273, 
    0.01253158, 0.2781332, 0.141384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2986155, 
    21.97212, 8.348226, 29.30048, 39.99499, 130.1351, 0.8950866, 0.01966914, 
    0.1630157, 0, 1.952829, 0.5040591, 0, 0, 0.01611275, 9.610229, 1.459349, 
    12.85996, 65.72018, 116.1776, 128.0019, 182.2513, 290.8639, 369.8836, 
    386.0753, 385.8762, 379.3724, 393.9282, 482.3826, 500.4763, 549.5696, 
    534.1202, 548.6902, 680.6912, 636.6417, 504.3287, 394.722, 296.3079, 
    208.9966, 140.6372, 97.57526, 13.33891, 0, 0, 0, 0, 0, 0, 0,
  3.996322, 0, 0, 0, 50.35525, 185.5548, 442.7651, 434.7867, 141.749, 
    8.424508, 0, 0, 0, 0, 0, 0.1385595, 0, 0.002443571, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001546636, 0, 
    0.01753371, 0.1784294, 55.34111, 40.54953, 0.06547624, 0, 18.5789, 
    0.6467119, 0, 0, 0.177912, 16.41363, 1.020464, 0, 0, 0.602079, 19.27653, 
    21.5851, 68.39326, 126.2266, 171.0694, 149.9013, 169.6777, 212.8275, 
    259.4587, 299.9385, 330.8089, 379.1569, 457.7391, 561.8567, 588.5029, 
    657.3253, 569.2491, 539.7734, 651.1829, 576.2408, 456.6287, 351.4606, 
    268.712, 186.3495, 104.8361, 52.63164, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0005410447, 0, 0, 217.2333, 150.0148, 147.8175, 59.43842, 0.09743718, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.004347128, 0.0005053915, 0, 0, 0, 0, 0, 
    108.7065, 172.8124, 10.6465, 39.72498, 0, 0.7019937, 0.6240747, 
    0.03666175, 3.923619, 11.28015, 0, 0, 0, 3.333197, 1.626409, 22.94781, 
    129.1699, 146.3097, 179.6523, 197.7332, 215.7947, 216.2458, 233.5067, 
    262.7396, 313.8624, 413.2129, 513.4584, 611.7216, 655.2258, 697.314, 
    587.9772, 544.4241, 623.3768, 528.1633, 394.2646, 303.2613, 223.6158, 
    176.0974, 98.5352, 40.67016, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.232757, 299.1098, 203.6477, 310.9305, 75.55457, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.001199378, 0, 0, 0, 0, 0, 424.0066, 651.8306, 74.5641, 
    110.6031, 137.6324, 0, 13.58554, 3.612053, 0, 0, 0, 0, 0, 4.653972, 
    12.98408, 132.1312, 225.6729, 202.1573, 187.3596, 223.9869, 245.0216, 
    232.7687, 241.0014, 265.6889, 318.4467, 431.9607, 541.9741, 643.3138, 
    668.8045, 639.2117, 512.8416, 507.6131, 530.3688, 426.9925, 321.1112, 
    237.3463, 202.2683, 173.7212, 111.4122, 27.88606, 0.0005438055, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 7.312272, 276.3273, 222.199, 363.1713, 12.21931, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90.08727, 874.5997, 248.2439, 134.9055, 
    106.5157, 0.7966748, 0.7750768, 0, 0, 0, 0, 0, 0, 0.2795637, 82.28407, 
    222.2338, 273.5854, 174.7247, 157.3741, 226.9098, 240.163, 230.1125, 
    254.5082, 294.148, 347.3311, 423.4855, 534.6428, 652.4855, 646.5594, 
    522.6107, 419.5539, 415.7138, 385.7757, 312.2747, 240.9982, 187.6149, 
    173.349, 160.6252, 114.4855, 27.0409, 0.0163472, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 160.1758, 213.3217, 235.5445, 48.00871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1112008, 2.781888, 0, 0, 0, 0, 0, 0, 0.003032611, 0.002118202, 
    0.5433614, 129.5313, 49.79841, 273.5827, 358.0385, 0.1867804, 9.040846, 
    16.79832, 2.512043, 0, 0, 0, 0, 0, 35.23597, 159.6615, 147.6077, 
    74.15279, 137.9986, 222.0329, 251.3415, 221.7983, 254.7236, 313.5164, 
    386.5862, 445.4337, 529.6935, 615.8958, 546.6193, 383.2585, 296.0247, 
    296.5038, 254.086, 225.9015, 197.0486, 177.1107, 159.7694, 143.3112, 
    134.4598, 60.69848, 9.276337, 0.07938728, 0.01935789, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 27.43061, 219.741, 182.4642, 145.6093, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14.73238, 8.035018, 0.002533916, 53.32179, 
    714.6627, 33.22498, 0, 0.08153576, 0, 0, 0, 0, 0, 0.1116458, 37.3478, 
    87.57549, 65.60155, 24.98499, 84.27135, 185.5645, 240.6545, 223.1828, 
    218.4679, 277.7992, 354.8269, 407.7614, 464.1208, 475.2428, 366.5284, 
    234.6922, 185.0667, 166.5074, 146.0874, 128.0777, 140.4522, 156.122, 
    159.8683, 152.9146, 170.7601, 142.2226, 55.40218, 25.69629, 0.2789844, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 118.9879, 364.7967, 262.5878, 200.3751, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0001877957, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.174198, 31.60677, 64.70731, 426.1732, 
    1363.807, 80.13299, 0, 0, 0, 0, 0, 0, 0.001290981, 2.815794, 26.87397, 
    19.16058, 8.644664, 1.876151, 39.90991, 143.068, 242.9099, 243.2124, 
    226.8486, 243.0945, 292.6472, 323.9382, 340.012, 310.8246, 220.8903, 
    156.6606, 105.6535, 84.0586, 78.32101, 71.50745, 87.09168, 128.866, 
    135.5459, 129.0692, 191.9514, 186.9409, 94.13192, 30.83496, 1.997563, 0, 
    0, 0, 0, 0,
  0, 0, 0.001936688, 46.618, 536.6373, 662.6491, 249.3386, 9.803163, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0001813781, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.459199, 103.5565, 
    661.9141, 1840.713, 219.5788, 0, 0, 0, 0, 0, 0, 0.1876374, 0.1116077, 
    4.196786, 0.6972661, 4.548798, 0.01515518, 19.67255, 135.7905, 257.0113, 
    277.3361, 253.3402, 236.5977, 238.597, 251.8898, 254.7406, 193.7241, 
    141.234, 99.71603, 61.99655, 29.32073, 13.64046, -0.03668842, 26.70518, 
    81.82543, 91.48897, 122.1683, 146.8756, 124.3265, 10.31211, 9.660895, 
    54.39833, 0.2762197, 0, 0, 0, 0,
  0, 0, 9.334058, 13.71354, 852.7475, 1096.084, 774.6525, 27.61173, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3280411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.112605, 141.024, 
    649.2419, 1983.348, 335.0366, 8.158025, 0.01285483, 1.803418, 2.566564, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.23637, 88.12022, 180.32, 243.7138, 259.6231, 
    232.9355, 205.8438, 203.9321, 192.951, 139.2836, 88.90681, 58.0747, 
    29.76662, 21.18993, 11.34657, 5.685978, 55.80595, 145.4924, 131.7599, 
    161.3288, 202.1818, 105.8592, 47.85705, 21.31422, 9.101623, 0, 0, 0, 0, 0,
  0, 0, 8.083728, 68.44715, 763.899, 819.9758, 573.8215, 67.20765, 0.8818858, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7558494, 202.6879, 
    672.795, 1732.209, 589.0763, 7.808373, 5.980556, 7.959057, 2.644362, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.5032064, 14.71771, 71.34007, 168.8776, 270.6567, 
    303.8179, 249.176, 188.3204, 150.6268, 103.42, 72.58722, 47.76024, 
    32.59775, 32.64248, 32.45184, 44.43424, 191.6641, 289.115, 320.5233, 
    411.2173, 393.0303, 296.0738, 190.0115, 73.94491, 0, 0, 0, 0, 0, 0,
  66.48343, 32.72926, 167.2516, 442.8591, 671.6302, 377.1797, 87.32704, 
    19.9507, 2.892875, 2.136357, 0.122568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003015865, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 80.25523, 370.7058, 1206.437, 775.0638, 72.39935, 
    11.08876, 20.55738, 1.923679, 0, 0, 0, 0, 0, 0, 0, 0, 0.7043098, 
    1.508858, 23.05793, 109.5643, 245.116, 339.6685, 319.9632, 211.4899, 
    138.8699, 98.34061, 73.37244, 64.12723, 38.16045, 37.41049, 28.51176, 
    38.78846, 65.09164, 118.0438, 185.5842, 257.3457, 215.2173, 108.8992, 
    78.36304, 35.72548, 8.264409, 4.238366, 0, 0, 0, 0,
  239.6041, 383.8715, 385.9552, 312.772, 354.1241, 158.2608, 13.44928, 
    4.439478, 0, 0, 0, 0, 0, 0.09766659, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004302262, 0.0009284276, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 65.84852, 257.2979, 725.2047, 976.9874, 203.7428, 
    26.53415, 26.40429, 12.97825, 0.3968416, 0, 0, 0, 0, 0, 0, 0, 0.2833899, 
    4.319847, 22.68953, 64.89889, 145.0534, 252.3569, 284.3854, 198.8476, 
    134.2758, 109.1641, 94.01095, 84.8871, 77.70658, 60.97504, 74.0986, 
    72.99908, 65.58603, 81.69981, 146.6016, 168.7964, 71.73798, 47.58058, 
    76.26965, 85.34253, 80.94412, 51.16417, 1.088907, 0, 0, 0,
  35.46908, 312.2523, 343.7193, 52.41047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1450596, 0.2184766, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.563134, 211.3301, 
    384.9349, 1012.969, 418.6268, 39.3827, 21.14776, 22.11357, 1.319225, 
    0.0001826946, 0.325497, 7.54947, 17.82139, 17.77085, 7.49655, 7.957342, 
    17.79939, 33.27032, 62.76324, 85.09935, 112.5088, 181.6462, 216.9371, 
    186.2492, 155.3895, 145.2876, 116.1752, 123.2312, 99.18019, 108.5044, 
    122.6949, 130.1461, 147.0177, 165.934, 161.3787, 95.41556, 49.94404, 
    50.94572, 86.07488, 121.9567, 174.7541, 113.5709, 7.699672, 0, 0, 0,
  0, 0, 0.5505809, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001916892, 
    0.488546, 0.3526058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01420734, 0, 156.4859, 171.2163, 
    1219.024, 1056.763, 227.3387, 20.19563, 22.60979, 1.255557, 6.144281, 
    45.4059, 62.7279, 97.57623, 101.1371, 78.44479, 56.55574, 70.73415, 
    121.4387, 190.2598, 228.6013, 167.1219, 186.6875, 214.2366, 206.5289, 
    194.4333, 173.067, 148.9911, 138.2063, 137.0002, 114.045, 110.0555, 
    138.2256, 143.1514, 155.9583, 107.2437, 61.62659, 60.00345, 62.52522, 
    75.2979, 158.1422, 252.193, 158.513, 1.751702, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002090689, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.008890191, 0, 67.49846, 202.0233, 1369.146, 1749.797, 
    579.0088, 20.74646, 6.495084, 0.0398635, 0, 0.4435986, 33.07759, 
    104.0203, 126.4093, 121.4114, 170.4067, 174.3627, 297.59, 418.0954, 
    490.278, 321.4501, 244.4302, 235.4262, 221.5576, 202.6546, 203.2396, 
    181.423, 183.7679, 160.8642, 143.6052, 126.7736, 119.1805, 123.6257, 
    103.5322, 71.23041, 75.24308, 72.00915, 65.68742, 95.67825, 220.7509, 
    320.3375, 166.0607, 14.94885, 1.212338, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3.35338, 0, 0, 0, 0, 0.0004769792, 0, 
    0.002373848, 0, 0, 0, 0, 0, 0, 0, 0, 0.01198174, 0, 1.170512, 26.17266, 
    920.9006, 1707.259, 548.358, 20.86545, 0, 0.02919498, 0, 8.295179e-05, 0, 
    0, 35.60873, 140.6726, 286.2187, 453.8871, 521.0576, 613.5406, 659.2684, 
    461.6195, 300.6107, 239.819, 229.6721, 231.9149, 274.6986, 262.3438, 
    217.9245, 185.6427, 156.8371, 124.7931, 111.6993, 114.7953, 105.9933, 
    95.67621, 83.49066, 78.79841, 74.49798, 111.6916, 266.0449, 268.2371, 
    42.25449, 0.02493712, 6.948849, 14.83968, 1.402666,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02394337, 0.2515746, 1.703864, 0.6291896, 0, 0.9544802, 1.295154, 
    1.900995, 1.829548, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003334169, 0.03683696, 0, 0, 61.67533, 497.1606, 1393.26, 921.786, 
    59.75617, 0, 0, 0, 0, 0, 0, 6.670186, 82.0864, 333.7366, 541.2671, 
    570.7663, 536.9034, 532.7047, 394.265, 316.7436, 281.2391, 283.4858, 
    317.4317, 337.6651, 311.4881, 252.3808, 196.0773, 158.135, 125.2839, 
    134.8932, 179.5908, 192.6594, 129.4154, 113.4966, 95.49207, 84.65179, 
    142.4767, 365.9221, 196.9136, 16.26885, 0, 0.993293, 210.9197, 320.5146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02792097, 0.3531507, 0.003153964, 0.09298629, 0, 0, 0, 0, 0, 
    0, 0, 0.0001550621, 0.0009271714, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007608135, 
    3.504901, 0.001191585, 14.31241, 84.53024, 1429.565, 1028.788, 570.2425, 
    25.71225, 0, 0, 0, 0, 0, 0, 0, 0.09222035, 52.24155, 104.2645, 261.9759, 
    312.8363, 286.0649, 269.9135, 332.5363, 391.7218, 436.5949, 425.3459, 
    349.5745, 251.7458, 185.8572, 143.547, 127.1319, 162.576, 240.0095, 
    253.7423, 196.6642, 167.1082, 130.5137, 139.8822, 425.961, 584.0701, 
    310.1891, 38.10512, 0.02188468, 0, 361.8489, 634.4559,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001512036, 0.001056419, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15.89228, 0.001179482, 0, 21.14887, 913.0068, 
    631.769, 1033.281, 837.3952, 31.48905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40.69078, 178.1973, 265.3913, 266.2013, 311.1905, 385.2721, 539.8588, 
    509.8239, 403.6374, 271.508, 176.3666, 138.3279, 123.0365, 145.8404, 
    203.9677, 254.9663, 219.4427, 240.7227, 267.1184, 484.1792, 681.328, 
    560.1155, 64.38747, 0.4352941, 0.003382807, 21.7661, 322.7632, 527.2258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7188078, 0, 0, 61.33807, 32.43402, 0.02485147, 145.2208, 627.1351, 
    287.4496, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.030678, 173.7331, 291.2982, 
    273.0661, 228.335, 327.7041, 474.7168, 494.3539, 377.0089, 256.2113, 
    177.9035, 140.8263, 131.356, 217.1942, 248.0046, 340.0473, 375.9899, 
    423.7958, 646.5859, 890.8132, 866.5603, 245.1126, 0, 0.05396707, 
    15.20921, 54.39197, 211.3136, 100.6684,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004543338, 0.003639919, 0, 
    0, 0, 0, 0, 0, 0, 3.531564, 0, 0, 0.7084563, 78.24866, 42.92502, 0, 0, 
    190.1828, 388.3742, 0, 0, 0, 0, 0, 0, 0.0004599308, 0, 0, 0, 13.8153, 
    130.9336, 144.9227, 177.9052, 219.8537, 376.9983, 361.93, 311.2201, 
    244.8839, 182.8421, 166.0394, 252.0663, 336.3086, 451.3323, 625.0237, 
    672.2084, 702.3406, 778.5399, 890.1186, 667.5145, 73.84701, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005854287, 0.00247674, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.313361, 16.38288, 0, 0, 147.3413, 142.4732, 0, 
    0.01397031, 50.75145, 186.9594, 0.1209901, 0, 0, 0, 0, 0, 0.000225285, 0, 
    0, 0, 0.01659336, 0.8779683, 47.25842, 88.2861, 235.9072, 276.3875, 
    324.9, 309.995, 270.1249, 234.3954, 347.3555, 412.644, 514.5791, 
    475.2197, 635.9094, 686.1741, 527.5653, 319.2344, 137.6655, 58.22589, 
    0.5826872, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001475661, 0.08985677, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0006000945, 5.420241, 14.74992, 9.866526, 369.6528, 
    31.99669, 0, 0.6211213, 22.01926, 26.09454, 0.01676102, 0, 0, 0, 0, 0, 
    0.0003724534, 0.0007511377, 0, 0, 0, 0.01054211, 4.9378, 35.11487, 
    209.5712, 293.8589, 365.6923, 371.3261, 394.2154, 492.1788, 710.024, 
    811.8054, 617.807, 343.5852, 201.6402, 88.6078, 33.18766, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002061675, 0.3639224, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.565544, 67.44887, 210.6318, 174.2347, 0, 0, 
    0.02026485, 0.5374939, 1.169389, 0.06065548, 0, 0, 0, 0, 0, 0.0005888037, 
    0, 0, 0, 0, 0, 0, 0.1444359, 50.93018, 158.3956, 294.5731, 366.2896, 
    503.3458, 626.3784, 834.7375, 746.9637, 477.1703, 102.5894, 2.179536, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0016285, 0.005161504, 
    0, 0, 0, 0, 0, 0, 0, 0.1744462, 11.87143, 189.9295, 0, 0, 0, 0, 3.378064, 
    2.925041, 6.432992, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001116622, 
    2.862813, 19.07391, 72.97668, 86.10835, 181.0871, 146.8998, 161.6484, 
    63.05329, 18.52388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.587682e-05, 0.0007486434, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003512555, 0, 0, 0.004746107, 0, 0, 0, 0, 0, 0, 0, 0, 0.001910802, 
    1.540883, 1.139802, 0, 0, 0, 0.00339965, 0, 5.067101, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7.394003e-05, 0, 0, 0, 0, 0, 0, 0, 0.1596736, 0.01119117, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002488717, 0, 0, 0, 
    0.00192382, 0, 0.0008238192, 0, 0, 0, 0, 0.004534618, 0.01042992, 
    128.6895, 111.6004, 0.9109875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 51.51996, 6.180326, 1.820795, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001911541, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009544371, 0, 24.92486, 51.07422, 23.80963, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.353347, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.248243, 20.32495, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.077861e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.002998321, 0.00326913, 0, 30.07554, 20.11271, 3.618359, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1637487, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001798506, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.00186227, 0, 0.03316185, 16.06968, 162.5954, 0, 
    3.422852, 0, 0, 0, 0, 0, 0, 0, 0.01038289, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001204468, 0, 0, 0.002527093, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66.34259, 22.89227, 15.44103, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001601016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06553058, 0.5628351, 51.22266, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9606495, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002309131, 
    0.6115905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.192964, 73.24959, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00447468, 0, 0, 0.001755983, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002103772, 1.21489, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 87.1916, 75.72276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.003544959, 0, 0, 0, 0, 0, 0, 0.0002654338, 0.001121242, 
    0.004204868, 0.001509032, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.04547353, 5.79191, 1.342976, 0.6890895, 0.2234796, 61.70195, 
    24.68652, 0, 0, 0, 0, 1.058887, 146.1155, 5.113419, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001511727, 0.00117502, 0.001633006, 
    0.007605216, 0, 0, 0, 0, 0, 0, 0, 0, 0.04061029, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1014451, 0, 1.253367, 0.0007692035, 16.09134, 27.76863, 48.46694, 
    11.74502, 0, 0, 0, 4.819854, 6.666916, 2.695935, 0, 0, 0, 0, 0, 0, 
    0.01972353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202.3895,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0006035659, 0, 0, 0, 0, 0, 0, 0.01408904, 0, 
    0.003578367, 0.004032353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03354037, 0, 0, 7.591219, 30.95796, 10.42947, 11.57776, 0, 0, 0, 
    2.446361, 0.008315299, 0, 0, 0, 0, 0, 0, 0.5451445, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 120.6041, 854.0955,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001588834, 0, 0, 0, 0.005239161, 0.009033938, 
    0.0005203752, 0.001356567, 0.001431737, 0.006111554, 0, 0, 0, 0, 0, 
    0.02182276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007873155, 0, 0, 0, 0, 0, 0, 
    18.8254, 15.31145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.272007, 709.054, 928.3032,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002614032, 0, 0.007351434, 
    0.003707968, 6.454103e-05, 0.001235135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0002616841, 0, 0, 0, 0, 0, 0, 0, 0.2473145, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    463.5101, 849.1191, 684.9581,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004843049, 0.002349587, 
    0.01799333, 0.00371025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004212329, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.004271484, 0, 0, 0, 0, 0, 0, 0, 0, 57.22657, 460.95, 639.7565, 
    519.5239, 33.79907,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001354043, 0, 
    0.006613636, 0.007528742, 0.02743311, 0.01341464, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003410095, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05400946, 4.694293, 0.3870355, 0, 0, 0, 0, 0, 141.1749, 
    601.933, 831.244, 543.7769, 58.66973, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01415738, 0.04210776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.679655, 
    105.733, 8.447727, 0, 0, 27.24204, 24.39606, 7.753161, 352.5742, 
    608.2495, 37.65978, 0.09178872, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01123114, 0.01882986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29.1145, 27.4687, 
    38.2424, 74.43308, 193.5007, 196.5712, 7.365326, 66.00092, 2.113855, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01327394, 0.003187717, 0, 0, 0.002941251, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.80582, 
    74.16306, 226.1258, 582.3444, 525.9813, 293.4045, 129.4705, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0153161, 0.005200402, 0, 0, 0, 0.003570459, 0.002388353, 0, 0, 0, 0, 
    0.1976552, 0, 0, 0, 0.1872808, 0.7276393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3034186, 214.9815, 492.9658, 326.6951, 
    73.56389, 0.05476749, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002162333, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9388899, 
    193.1229, 6.378803, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 258.6678, 289.7753, 3.976977, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.009249282, 0.001536941, 0, 0, 0, 0, 0, 0, 0, 40.0586, 
    32.99025, 2.803985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.30081, 1.451902, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0009401445, 0.0004037078, 0, 0, 0, 0, 
    0.1391184, 50.75321, 3.125369, 1.116508, 0.2084151, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933637, 0.05200977, 
    1.095076, 0.4746633, 0, 0.0152259, 0.00121065, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003794074, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.873821, 0, 0, 0, 
    0.0909774, 0.106935, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04739007, 0.5167308, 
    0.02355359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005289078, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0004078763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.796603,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.600741e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008196245, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2539265, 0, 
    0.1848694, 0, 0, 0, 0, 0, 0, 0.02119472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.612157,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009860342, 0, 0, 0, 
    0.5821458, 1.014729, 1.475074, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007580966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00020889, 0.003413063, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.08453731, 0, 0.6124651, 0.0904895, 0.04531468, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.060883, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006160314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0004963353, 0, 0.002697561, 0, 0, 0, 
    0.002501344, 0.003084639, 0, 0, 0, 60.34301, 23.29774, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001295554, 0.002088146, 0, 0, 0, 0, 0.003850434, 0, 0.003216584, 
    0, 0, 6.297387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2759891, 0, 0, 0, 0, 1.456678, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002685973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.603688, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.042054e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003275427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001260254, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004184085, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001634963, 0, 0, 0, 0, 
    0.00182365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004781314, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002623971, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1032847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02264775, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01294437, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45.58595, 
    19.94605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01843011, 0, 0, 0, 0, 0.0006814443, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05284531, 0, 0.2416257, 0.6087035, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01169867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009131898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006104111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002335767, 39.18405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0105723, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01319931, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1318502, 0, 0, 0.3468482, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45.02456, 0.7059237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0927918, 0.01668262, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0472814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    140.8308, 155.7868, 125.8311, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02154752, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    749.9999, 457.7867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.01483413, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.498203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002601753, 
    0.002704989, 0, 0, 0, 0, 0, 0, 0.001969324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003557655, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02448131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00550229, 0, 0, 0, 0, 0.0046798, 
    1.793624, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.448954, 0, 
    0.00866163, 0, 0, 0, 0, 0.4479904, 0.01966327, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005507405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.460738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03048245, 
    61.25506, 0, 0, 0, 0, 0, 0, 0.3824942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02183831, 
    0.2123545, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04637172, 
    0.008339238, 0, 0, 0.03448581, 0, 0, 0, 0, 0, 0, 0, 0.196157, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005239569, 
    0.0212123, 0.0003524371, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02602657, 
    0.02576878, 0.0369913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01774269, 
    0.006849611, 0.01812511, 0.007378699, 0.04169989, 0, 0, 0, 0.0002408772, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.500448, 0.6373758, 0.3299181, 0.2709744, 0.3045332, 
    0.9904844, 1, 0.7193916, 0.6372474, 0.08596428, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2001312, 0.4111539, 0, 0, 0, 0, 0, 0, 
    0.3257935, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9846206, 0.1322953, 0, 0, 0,
  0.4213375, 0.7249894, 0.1194391, 0.4090452, 0.0004055478, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1275371, 0.2101071, 0.501195, 0.907451, 0.5348656, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.2795206, 0, 0, 0, 0, 0, 0, 0.4748606, 0.08597825, 0, 
    0, 0, 0, 0, 0.3374754, 0.9515835, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.974499, 0.2595553, 0, 0, 0, 0,
  1, 1, 0.5694539, 0.2257697, 0.07591473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1566211, 0, 0, 0, 0.3620377, 0, 0, 0, 0, 0, 0, 
    0.2321739, 0, 0, 0, 0, 0, 0, 0.6652638, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6224186, 0, 0, 0, 0, 0,
  1, 1, 0.5671622, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0328016, 0.3505093, 0.800697, 0.4199587, 0.3645951, 0.2070305, 
    0.1039276, 0.04041792, 0.1039293, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3621618, 0.9914034, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.9980344, 0.1799124, 0, 0, 0, 0, 0,
  1, 1, 0.6025393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0554254, 0.07674838, 0.3268177, 0.2018002, 0, 0, 0, 0.2147634, 
    0.246665, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1000221, 0.9995502, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9989821, 
    0.4096552, 0, 0, 0, 0, 0, 0,
  0.628101, 0.6280472, 0.4677134, 0, 0, 0.3171421, 0.0938872, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2612283, 0.06390974, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3284912, 0.3768882, 0.8638445, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7643126, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.05901703, 0.9235198, 0.8531228, 0.7637583, 0.2779488, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0508899, 0.05089059, 0.3887566, 
    0.2545041, 0.2612266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4230824, 0.09009741, 
    0.4622726, 0.9831397, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.3566395, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.3848666, 0.9172006, 1, 1, 0.8194785, 0.02148438, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1404992, 0.4942557, 0, 0, 0.1406009, 0, 
    0, 0, 0, 0.2166595, 0, 0, 0, 0.02490224, 0.9627016, 0.8158007, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9282088, 
    0.03051941, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.5683897, 0.9379957, 0.6364555, 0.2024043, 0.03349722, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.320924, 0.9845472, 0.2649983, 
    0.1140551, 0, 0, 0, 0, 0, 0.01618783, 0, 0, 0, 0.08289424, 0.1259722, 
    0.8170571, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7655389, 0.005966454, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0272528, 0.8907499, 0.9876926, 0.7710279, 0.1670542, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4784564, 1, 0.6486406, 0.6920749, 
    0.2536378, 0, 0, 0, 0, 0, 0, 0, 0, 0.2509409, 0.8028153, 0.9793605, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7416639, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.648589, 1, 0.9992579, 0.2293907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.09293438, 0.9501851, 0.8690677, 1, 0.5762319, 0, 
    0, 0.008900359, 0.003358786, 0, 0, 0, 0, 0.0356602, 0.9891973, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3823546, 
    0.00315241, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.4935699, 1, 0.7489711, 0.1704132, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1722069, 0.2898026, 1, 0.8352928, 0.0001595881, 
    0.2050383, 0.6669478, 0.1472481, 0, 0, 0, 0, 0, 0.7378939, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.3177179, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.3381471, 0.9340628, 0.9308964, 0.34702, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0710042, 0.01311141, 0.01958092, 0.2182962, 
    0.9644061, 0.2152033, 0.07139239, 0.07196605, 0, 0, 0, 0, 0, 0, 
    0.8858101, 1, 0.933995, 0.8029567, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8098463, 0.2802811, 0.06792729, 0, 0, 0, 0, 0,
  0, 0, 0, 0.062082, 0.4496638, 0.9014636, 1, 0.6371259, 0.0002500278, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07396818, 0.06363945, 0.2273634, 
    0.7217154, 1, 0.4123627, 0, 0, 0, 0, 0, 0, 0, 0.03488547, 0.9638747, 
    0.4518672, 0.2722468, 0.101736, 0.9105512, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.8664908, 0.293852, 0.1126182, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0.1481497, 0.8071872, 1, 0.9563567, 0.1187265, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09094947, 0.8744214, 1, 1, 0.6151962, 
    7.862093e-05, 0, 0, 0, 0, 0, 0, 0.05432393, 0.3167762, 0, 0.1943092, 0, 
    0.6416867, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9944282, 0.1187612, 0.2975091, 0.5171648, 0, 0, 0, 0, 0,
  0, 0, 0, 0.006354006, 0.888454, 1, 1, 0.1866042, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2678939, 1, 1, 1, 0.9953833, 0.4038017, 0, 
    0.1863101, 0.1370078, 0, 0, 0, 0, 0, 0, 0, 0, 0.1708246, 0.9664814, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.643471, 
    0.3777492, 0.3611507, 0, 0, 0, 0, 0,
  0, 0, 0, 0.2080797, 0.9673514, 1, 0.8374537, 0.04476063, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01296526, 0.7596481, 1, 1, 1, 
    0.9865646, 0.8895645, 0.9378822, 0.2410906, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01894641, 0.7163382, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9017419, 0.4822293, 0.01936743, 0, 0, 0, 0, 0,
  0.2283506, 0.2283831, 0.3606219, 0.8600088, 1, 1, 0.8187755, 0.09858553, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3482806, 1, 1, 1, 1, 
    1, 1, 0.2386805, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04633646, 0.8615492, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.850582, 0.348906, 
    0.139303, 0, 0, 0, 0,
  0.9058077, 1, 1, 0.9630018, 0.8670257, 0.6587394, 0.3201251, 0.1648381, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1173386, 1, 1, 1, 1, 
    1, 1, 0.7136791, 0.01745822, 0, 0, 0, 0, 0, 0, 0, 0.0606117, 0.3882409, 
    0.9743452, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.784731, 0.03699823, 0, 0, 0,
  0.4231035, 0.9422162, 0.9297223, 0.3348973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01853104, 0.8556062, 1, 1, 1, 1, 1, 
    1, 0.08117965, 0.02060091, 0.04679306, 0.4853819, 0.590209, 0.5901864, 
    0.5901626, 0.5901374, 0.7937525, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9957187, 0.1070087, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.5207784, 1, 1, 1, 1, 1, 0.9874919, 0.008527548, 0.2921969, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.9391072, 0.1130477, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1617553, 0.9999905, 1, 1, 1, 0.92387, 0.5260675, 0, 0.004612686, 
    0.03066925, 0.3373398, 0.5646344, 0.7950864, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9652795, 
    0.03719426, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01460301, 0.8115592, 1, 1, 1, 0.1636489, 0, 0, 0, 0, 0, 0, 
    0.6152393, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8714985, 0.2261804, 0, 0, 0.3437575, 0.01257803,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2064631, 0.733834, 1, 1, 0.3149392, 0, 0, 0, 0, 0, 0, 
    0.2648452, 0.6866553, 0.7366514, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9174272, 0.1166509, 0, 0.05494488, 
    0.9094183, 0.8397222,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.07105455, 0, 0, 0.1277506, 0.9753432, 1, 0.6722792, 0.08202832, 0, 
    0, 0, 0, 0, 0, 0, 0.04108687, 0.2125929, 0.6796362, 0.8867523, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4437395, 0, 
    0.003395685, 0.9062591, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.06928185, 0, 0, 0, 0.6190757, 0.4693122, 0.9500455, 0.8051443, 
    0.06908886, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5560373, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9714394, 0.4920565, 0.007317367, 0, 
    0.1679957, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1870881, 0.1032061, 0, 0.3068611, 0.901248, 0.525517, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.08475742, 0.9234713, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7293079, 0, 0, 0.4481606, 0.3670389, 
    0.8051461, 0.3047968,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2969156, 0.1804042, 0, 0, 0.6011499, 0.5948403, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.3606173, 0.8423501, 0.9566985, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9882501, 0.4393826, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1341057, 0, 0, 0.3335736, 0.2354348, 0, 0, 0.225836, 0.4429893, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7404009, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.9729695, 0.7830737, 0.3542824, 0.3088061, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.08371773, 0.6231546, 0.07811955, 0, 0, 0.1299088, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1582873, 0.6573294, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9011589, 0.4768529, 0.2806725, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.4617452, 0.2357396, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.05252013, 0.5075252, 0.9784946, 1, 1, 1, 1, 1, 1, 
    0.9491259, 0.6694556, 0.0476924, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2044773, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1850218, 0.3838319, 0.3948988, 0.6347017, 0.897539, 0.8975486, 
    0.625631, 0.3950224, 0.1931382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.04801759, 0.008659004, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.2955928, 0.4134034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2288118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1252723, 0.02888734, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1657154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1331506, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2602637, 
    0.1827536, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.308817, 
    0.1388956, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009059105, 
    0.04102035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1710694,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1561902, 
    0.9037677,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7994146, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02431367, 
    0.5217998, 1, 0.9833409,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03587419, 0.3440025, 
    0.8423416, 1, 0.9747218, 0.3018562,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001283266, 0.05145107, 0, 0, 0, 0, 0, 
    0.4153767, 0.9991337, 1, 0.9749234, 0.6001224, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001449973, 0.7731972, 0.1336049, 0, 0, 
    0.1802618, 0.1813705, 0, 0.8987046, 0.7961607, 0.290663, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3244956, 0.5728012, 0.6642565, 
    0.6642635, 0.7536004, 0.7371183, 0.09692896, 0.2581114, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01432, 0.7955128, 1, 1, 1, 
    0.8594135, 0.4985357, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008547029, 0.6526902, 0.9749812, 
    0.7542722, 0.4022479, 0.04722129, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3207461, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8175688, 0.8197373, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3270165, 0.08929753, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1860417, 
    0.1124855, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2794361, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1755751,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05289424,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2801953, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004320362, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2700683, 0.1831646, 0.1345469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5860988, 0.2863249, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 zsurf =
  0.05263353, 0.9425675, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.210776, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.252779, 74.21071, 95.69428, 
    40.84037, 37.33909, 173.0547, 413.3694, 558.9451, 332.2694, 351.5737, 
    71.52609, 0.03417388, 1.300127, 17.79588, 8.458535, 18.73478, 17.63159, 
    0, 0, 0, 24.16101, 0, 0, 0, 0, 0, 0, 0, 1.372658, 299.2773, 291.463, 0, 
    0, 0, 0, 0, 0.0248737, 34.27986, 188.9342, 329.4237, 350.9251, 251.6835, 
    165.8015, 165.6417, 201.2802, 268.5535, 314.2737, 338.9506, 356.3144, 
    377.6248, 410.6694, 439.9049, 453.2951, 445.0014, 438.5307, 407.9247, 
    339.9653, 265.3149, 224.8092, 190.4008, 158.7892, 103.6094, 19.02374, 0, 
    0, 0,
  9.158454, 18.90683, 3.012916, 53.90588, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2984579, 4.255527, 
    84.79544, 147.7691, 233.7292, 347.7168, 36.84171, 0, 0, 0, 0, 0, 0, 
    0.4999831, 0, 0, 0, 25.2615, 9.891716, 381.2982, 0.7240577, 0, 0, 0, 0, 
    147.3826, 251.5665, 17.10577, 0, 0, 0, 0, 0, 12.48063, 173.854, 367.2847, 
    472.174, 458.6521, 325.3309, 227.1559, 236.9397, 249.4832, 296.6798, 
    348.9885, 370.6396, 368.1631, 393.7355, 411.4686, 451.679, 461.741, 
    457.9003, 439.6093, 391.6231, 291.6416, 227.3665, 205.8765, 180.0435, 
    108.2699, 20.55778, 0, 0, 0, 0,
  146.5898, 178.415, 28.03686, 31.16747, 0, 0, 0, 0, 0, 0, 0, 0, 0.03837012, 
    1.052421, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.03251622, 0.6342183, 0, 0.003365346, 0.1732605, 15.05509, 
    0.627657, 0, 0, 5.064898, 0.5615213, 22.54741, 2.144348, 0, 0, 255.0734, 
    8.867086, 0, 0, 0.008958309, 1.017161, 28.21741, 115.5201, 0, 0, 0, 0, 0, 
    0, 66.54465, 223.7023, 341.7935, 467.8122, 479.3343, 405.95, 344.1333, 
    317.8734, 316.412, 353.7882, 397.7623, 399.601, 410.1562, 420.6944, 
    456.795, 491.1674, 486.9185, 461.8076, 437.4255, 366.8581, 265.5489, 
    220.6245, 207.5233, 145.059, 52.48993, 0.02635965, 0, 0, 0, 0,
  312.5654, 332.0361, 48.98602, 0.01820307, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2560336, 10.64937, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6525263, 85.40112, 154.1216, 
    145.2693, 104.7963, 68.44398, 59.66086, 5.658707, 51.90486, 0, 
    0.0002234011, 0.002236324, 0, 4.058273, 2.615149, 0, 0, 0, 0, 0, 0, 0, 
    45.61565, 143.503, 253.2654, 347.6613, 440.0746, 419.2403, 373.5648, 
    356.8692, 343.2001, 372.7208, 395.3455, 415.5849, 430.8153, 461.9744, 
    506.336, 526.5826, 478.6951, 428.0603, 393.4123, 322.4732, 237.9073, 
    211.1528, 175.5259, 95.53486, 5.59942, 0, 0, 0, 0, 0,
  277.1137, 216.7668, 65.78798, 0.01913495, 0, 6.423023, 0.05600383, 0, 0, 0, 
    0.008824782, 0.03805306, 5.421787, 6.542611, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.47252, 
    50.65664, 159.9921, 46.69725, 1.587591, 2.254171, 0.6875598, 155.2946, 
    109.7841, 0, 0, 0, 0, 6.335535, 1.460464, 0, 0, 0, 0, 0, 0, 0, 
    0.001764559, 51.18093, 107.6214, 220.6243, 313.7549, 357.301, 394.333, 
    380.0004, 369.1454, 378.0013, 370.4623, 409.9088, 457.2517, 510.6886, 
    598.5809, 591.0898, 488.7568, 418.8461, 368.6212, 287.8756, 211.7777, 
    183.3996, 128.3429, 26.55859, 0, 0, 0, 0, 0, 0,
  212.3771, 135.9476, 49.42075, 12.49728, 1.597956, 29.35641, 0.7934011, 
    2.107809, 0.008830293, 0.1460706, 1.322528, 19.1708, 1.042597, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1036084, 1.6234, 0.4369082, 1.249874, 151.7508, 
    165.1876, 0.1203202, 0, 0, 0.966633, 12.21299, 9.954236, 0, 0, 0, 0, 0, 
    0, 3.324982, 15.32631, 53.0812, 144.7708, 241.6709, 340.8276, 409.1607, 
    415.9962, 398.8717, 383.6034, 399.2011, 408.1645, 448.2938, 490.6762, 
    554.4016, 678.0546, 651.3043, 520.1175, 420.8705, 346.4621, 250.8538, 
    183.0857, 142.4498, 71.22203, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.2228342, 92.88892, 92.60233, 105.3637, 26.52375, 48.40273, 
    0.01253158, 0.2781332, 0.141384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2986155, 
    21.97212, 8.348226, 29.30048, 39.99499, 130.1351, 0.8950866, 0.01966914, 
    0.1630157, 0, 1.952829, 0.5040591, 0, 0, 0.01611275, 9.610229, 1.459349, 
    12.85996, 65.72018, 116.1776, 128.0019, 182.2513, 290.8639, 369.8836, 
    386.0753, 385.8762, 379.3724, 393.9282, 482.3826, 500.4763, 549.5696, 
    534.1202, 548.6902, 680.6912, 636.6417, 504.3287, 394.722, 296.3079, 
    208.9966, 140.6372, 97.57526, 13.33891, 0, 0, 0, 0, 0, 0, 0,
  3.996322, 0, 0, 0, 50.35525, 185.5548, 442.7651, 434.7867, 141.749, 
    8.424508, 0, 0, 0, 0, 0, 0.1385595, 0, 0.002443571, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001546636, 0, 
    0.01753371, 0.1784294, 55.34111, 40.54953, 0.06547624, 0, 18.5789, 
    0.6467119, 0, 0, 0.177912, 16.41363, 1.020464, 0, 0, 0.602079, 19.27653, 
    21.5851, 68.39326, 126.2266, 171.0694, 149.9013, 169.6777, 212.8275, 
    259.4587, 299.9385, 330.8089, 379.1569, 457.7391, 561.8567, 588.5029, 
    657.3253, 569.2491, 539.7734, 651.1829, 576.2408, 456.6287, 351.4606, 
    268.712, 186.3495, 104.8361, 52.63164, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0005410447, 0, 0, 217.2333, 150.0148, 147.8175, 59.43842, 0.09743718, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.004347128, 0.0005053915, 0, 0, 0, 0, 0, 
    108.7065, 172.8124, 10.6465, 39.72498, 0, 0.7019937, 0.6240747, 
    0.03666175, 3.923619, 11.28015, 0, 0, 0, 3.333197, 1.626409, 22.94781, 
    129.1699, 146.3097, 179.6523, 197.7332, 215.7947, 216.2458, 233.5067, 
    262.7396, 313.8624, 413.2129, 513.4584, 611.7216, 655.2258, 697.314, 
    587.9772, 544.4241, 623.3768, 528.1633, 394.2646, 303.2613, 223.6158, 
    176.0974, 98.5352, 40.67016, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3.232757, 299.1098, 203.6477, 310.9305, 75.55457, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.001199378, 0, 0, 0, 0, 0, 424.0066, 651.8306, 74.5641, 
    110.6031, 137.6324, 0, 13.58554, 3.612053, 0, 0, 0, 0, 0, 4.653972, 
    12.98408, 132.1312, 225.6729, 202.1573, 187.3596, 223.9869, 245.0216, 
    232.7687, 241.0014, 265.6889, 318.4467, 431.9607, 541.9741, 643.3138, 
    668.8045, 639.2117, 512.8416, 507.6131, 530.3688, 426.9925, 321.1112, 
    237.3463, 202.2683, 173.7212, 111.4122, 27.88606, 0.0005438055, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 7.312272, 276.3273, 222.199, 363.1713, 12.21931, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90.08727, 874.5997, 248.2439, 134.9055, 
    106.5157, 0.7966748, 0.7750768, 0, 0, 0, 0, 0, 0, 0.2795637, 82.28407, 
    222.2338, 273.5854, 174.7247, 157.3741, 226.9098, 240.163, 230.1125, 
    254.5082, 294.148, 347.3311, 423.4855, 534.6428, 652.4855, 646.5594, 
    522.6107, 419.5539, 415.7138, 385.7757, 312.2747, 240.9982, 187.6149, 
    173.349, 160.6252, 114.4855, 27.0409, 0.0163472, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 160.1758, 213.3217, 235.5445, 48.00871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1112008, 2.781888, 0, 0, 0, 0, 0, 0, 0.003032611, 0.002118202, 
    0.5433614, 129.5313, 49.79841, 273.5827, 358.0385, 0.1867804, 9.040846, 
    16.79832, 2.512043, 0, 0, 0, 0, 0, 35.23597, 159.6615, 147.6077, 
    74.15279, 137.9986, 222.0329, 251.3415, 221.7983, 254.7236, 313.5164, 
    386.5862, 445.4337, 529.6935, 615.8958, 546.6193, 383.2585, 296.0247, 
    296.5038, 254.086, 225.9015, 197.0486, 177.1107, 159.7694, 143.3112, 
    134.4598, 60.69848, 9.276337, 0.07938728, 0.01935789, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 27.43061, 219.741, 182.4642, 145.6093, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14.73238, 8.035018, 0.002533916, 53.32179, 
    714.6627, 33.22498, 0, 0.08153576, 0, 0, 0, 0, 0, 0.1116458, 37.3478, 
    87.57549, 65.60155, 24.98499, 84.27135, 185.5645, 240.6545, 223.1828, 
    218.4679, 277.7992, 354.8269, 407.7614, 464.1208, 475.2428, 366.5284, 
    234.6922, 185.0667, 166.5074, 146.0874, 128.0777, 140.4522, 156.122, 
    159.8683, 152.9146, 170.7601, 142.2226, 55.40218, 25.69629, 0.2789844, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 118.9879, 364.7967, 262.5878, 200.3751, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0001877957, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.174198, 31.60677, 64.70731, 426.1732, 
    1363.807, 80.13299, 0, 0, 0, 0, 0, 0, 0.001290981, 2.815794, 26.87397, 
    19.16058, 8.644664, 1.876151, 39.90991, 143.068, 242.9099, 243.2124, 
    226.8486, 243.0945, 292.6472, 323.9382, 340.012, 310.8246, 220.8903, 
    156.6606, 105.6535, 84.0586, 78.32101, 71.50745, 87.09168, 128.866, 
    135.5459, 129.0692, 191.9514, 186.9409, 94.13192, 30.83496, 1.997563, 0, 
    0, 0, 0, 0,
  0, 0, 0.001936688, 46.618, 536.6373, 662.6491, 249.3386, 9.803163, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0001813781, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.459199, 103.5565, 
    661.9141, 1840.713, 219.5788, 0, 0, 0, 0, 0, 0, 0.1876374, 0.1116077, 
    4.196786, 0.6972661, 4.548798, 0.01515518, 19.67255, 135.7905, 257.0113, 
    277.3361, 253.3402, 236.5977, 238.597, 251.8898, 254.7406, 193.7241, 
    141.234, 99.71603, 61.99655, 29.32073, 13.64046, -0.03668842, 26.70518, 
    81.82543, 91.48897, 122.1683, 146.8756, 124.3265, 10.31211, 9.660895, 
    54.39833, 0.2762197, 0, 0, 0, 0,
  0, 0, 9.334058, 13.71354, 852.7475, 1096.084, 774.6525, 27.61173, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3280411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.112605, 141.024, 
    649.2419, 1983.348, 335.0366, 8.158025, 0.01285483, 1.803418, 2.566564, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.23637, 88.12022, 180.32, 243.7138, 259.6231, 
    232.9355, 205.8438, 203.9321, 192.951, 139.2836, 88.90681, 58.0747, 
    29.76662, 21.18993, 11.34657, 5.685978, 55.80595, 145.4924, 131.7599, 
    161.3288, 202.1818, 105.8592, 47.85705, 21.31422, 9.101623, 0, 0, 0, 0, 0,
  0, 0, 8.083728, 68.44715, 763.899, 819.9758, 573.8215, 67.20765, 0.8818858, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7558494, 202.6879, 
    672.795, 1732.209, 589.0763, 7.808373, 5.980556, 7.959057, 2.644362, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.5032064, 14.71771, 71.34007, 168.8776, 270.6567, 
    303.8179, 249.176, 188.3204, 150.6268, 103.42, 72.58722, 47.76024, 
    32.59775, 32.64248, 32.45184, 44.43424, 191.6641, 289.115, 320.5233, 
    411.2173, 393.0303, 296.0738, 190.0115, 73.94491, 0, 0, 0, 0, 0, 0,
  66.48343, 32.72926, 167.2516, 442.8591, 671.6302, 377.1797, 87.32704, 
    19.9507, 2.892875, 2.136357, 0.122568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003015865, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 80.25523, 370.7058, 1206.437, 775.0638, 72.39935, 
    11.08876, 20.55738, 1.923679, 0, 0, 0, 0, 0, 0, 0, 0, 0.7043098, 
    1.508858, 23.05793, 109.5643, 245.116, 339.6685, 319.9632, 211.4899, 
    138.8699, 98.34061, 73.37244, 64.12723, 38.16045, 37.41049, 28.51176, 
    38.78846, 65.09164, 118.0438, 185.5842, 257.3457, 215.2173, 108.8992, 
    78.36304, 35.72548, 8.264409, 4.238366, 0, 0, 0, 0,
  239.6041, 383.8715, 385.9552, 312.772, 354.1241, 158.2608, 13.44928, 
    4.439478, 0, 0, 0, 0, 0, 0.09766659, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004302262, 0.0009284276, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 65.84852, 257.2979, 725.2047, 976.9874, 203.7428, 
    26.53415, 26.40429, 12.97825, 0.3968416, 0, 0, 0, 0, 0, 0, 0, 0.2833899, 
    4.319847, 22.68953, 64.89889, 145.0534, 252.3569, 284.3854, 198.8476, 
    134.2758, 109.1641, 94.01095, 84.8871, 77.70658, 60.97504, 74.0986, 
    72.99908, 65.58603, 81.69981, 146.6016, 168.7964, 71.73798, 47.58058, 
    76.26965, 85.34253, 80.94412, 51.16417, 1.088907, 0, 0, 0,
  35.46908, 312.2523, 343.7193, 52.41047, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1450596, 0.2184766, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.563134, 211.3301, 
    384.9349, 1012.969, 418.6268, 39.3827, 21.14776, 22.11357, 1.319225, 
    0.0001826946, 0.325497, 7.54947, 17.82139, 17.77085, 7.49655, 7.957342, 
    17.79939, 33.27032, 62.76324, 85.09935, 112.5088, 181.6462, 216.9371, 
    186.2492, 155.3895, 145.2876, 116.1752, 123.2312, 99.18019, 108.5044, 
    122.6949, 130.1461, 147.0177, 165.934, 161.3787, 95.41556, 49.94404, 
    50.94572, 86.07488, 121.9567, 174.7541, 113.5709, 7.699672, 0, 0, 0,
  0, 0, 0.5505809, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001916892, 
    0.488546, 0.3526058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01420734, 0, 156.4859, 171.2163, 
    1219.024, 1056.763, 227.3387, 20.19563, 22.60979, 1.255557, 6.144281, 
    45.4059, 62.7279, 97.57623, 101.1371, 78.44479, 56.55574, 70.73415, 
    121.4387, 190.2598, 228.6013, 167.1219, 186.6875, 214.2366, 206.5289, 
    194.4333, 173.067, 148.9911, 138.2063, 137.0002, 114.045, 110.0555, 
    138.2256, 143.1514, 155.9583, 107.2437, 61.62659, 60.00345, 62.52522, 
    75.2979, 158.1422, 252.193, 158.513, 1.751702, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002090689, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.008890191, 0, 67.49846, 202.0233, 1369.146, 1749.797, 
    579.0088, 20.74646, 6.495084, 0.0398635, 0, 0.4435986, 33.07759, 
    104.0203, 126.4093, 121.4114, 170.4067, 174.3627, 297.59, 418.0954, 
    490.278, 321.4501, 244.4302, 235.4262, 221.5576, 202.6546, 203.2396, 
    181.423, 183.7679, 160.8642, 143.6052, 126.7736, 119.1805, 123.6257, 
    103.5322, 71.23041, 75.24308, 72.00915, 65.68742, 95.67825, 220.7509, 
    320.3375, 166.0607, 14.94885, 1.212338, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3.35338, 0, 0, 0, 0, 0.0004769792, 0, 
    0.002373848, 0, 0, 0, 0, 0, 0, 0, 0, 0.01198174, 0, 1.170512, 26.17266, 
    920.9006, 1707.259, 548.358, 20.86545, 0, 0.02919498, 0, 8.295179e-05, 0, 
    0, 35.60873, 140.6726, 286.2187, 453.8871, 521.0576, 613.5406, 659.2684, 
    461.6195, 300.6107, 239.819, 229.6721, 231.9149, 274.6986, 262.3438, 
    217.9245, 185.6427, 156.8371, 124.7931, 111.6993, 114.7953, 105.9933, 
    95.67621, 83.49066, 78.79841, 74.49798, 111.6916, 266.0449, 268.2371, 
    42.25449, 0.02493712, 6.948849, 14.83968, 1.402666,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02394337, 0.2515746, 1.703864, 0.6291896, 0, 0.9544802, 1.295154, 
    1.900995, 1.829548, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003334169, 0.03683696, 0, 0, 61.67533, 497.1606, 1393.26, 921.786, 
    59.75617, 0, 0, 0, 0, 0, 0, 6.670186, 82.0864, 333.7366, 541.2671, 
    570.7663, 536.9034, 532.7047, 394.265, 316.7436, 281.2391, 283.4858, 
    317.4317, 337.6651, 311.4881, 252.3808, 196.0773, 158.135, 125.2839, 
    134.8932, 179.5908, 192.6594, 129.4154, 113.4966, 95.49207, 84.65179, 
    142.4767, 365.9221, 196.9136, 16.26885, 0, 0.993293, 210.9197, 320.5146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02792097, 0.3531507, 0.003153964, 0.09298629, 0, 0, 0, 0, 0, 
    0, 0, 0.0001550621, 0.0009271714, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007608135, 
    3.504901, 0.001191585, 14.31241, 84.53024, 1429.565, 1028.788, 570.2425, 
    25.71225, 0, 0, 0, 0, 0, 0, 0, 0.09222035, 52.24155, 104.2645, 261.9759, 
    312.8363, 286.0649, 269.9135, 332.5363, 391.7218, 436.5949, 425.3459, 
    349.5745, 251.7458, 185.8572, 143.547, 127.1319, 162.576, 240.0095, 
    253.7423, 196.6642, 167.1082, 130.5137, 139.8822, 425.961, 584.0701, 
    310.1891, 38.10512, 0.02188468, 0, 361.8489, 634.4559,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001512036, 0.001056419, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15.89228, 0.001179482, 0, 21.14887, 913.0068, 
    631.769, 1033.281, 837.3952, 31.48905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    40.69078, 178.1973, 265.3913, 266.2013, 311.1905, 385.2721, 539.8588, 
    509.8239, 403.6374, 271.508, 176.3666, 138.3279, 123.0365, 145.8404, 
    203.9677, 254.9663, 219.4427, 240.7227, 267.1184, 484.1792, 681.328, 
    560.1155, 64.38747, 0.4352941, 0.003382807, 21.7661, 322.7632, 527.2258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7188078, 0, 0, 61.33807, 32.43402, 0.02485147, 145.2208, 627.1351, 
    287.4496, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.030678, 173.7331, 291.2982, 
    273.0661, 228.335, 327.7041, 474.7168, 494.3539, 377.0089, 256.2113, 
    177.9035, 140.8263, 131.356, 217.1942, 248.0046, 340.0473, 375.9899, 
    423.7958, 646.5859, 890.8132, 866.5603, 245.1126, 0, 0.05396707, 
    15.20921, 54.39197, 211.3136, 100.6684,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004543338, 0.003639919, 0, 
    0, 0, 0, 0, 0, 0, 3.531564, 0, 0, 0.7084563, 78.24866, 42.92502, 0, 0, 
    190.1828, 388.3742, 0, 0, 0, 0, 0, 0, 0.0004599308, 0, 0, 0, 13.8153, 
    130.9336, 144.9227, 177.9052, 219.8537, 376.9983, 361.93, 311.2201, 
    244.8839, 182.8421, 166.0394, 252.0663, 336.3086, 451.3323, 625.0237, 
    672.2084, 702.3406, 778.5399, 890.1186, 667.5145, 73.84701, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005854287, 0.00247674, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.313361, 16.38288, 0, 0, 147.3413, 142.4732, 0, 
    0.01397031, 50.75145, 186.9594, 0.1209901, 0, 0, 0, 0, 0, 0.000225285, 0, 
    0, 0, 0.01659336, 0.8779683, 47.25842, 88.2861, 235.9072, 276.3875, 
    324.9, 309.995, 270.1249, 234.3954, 347.3555, 412.644, 514.5791, 
    475.2197, 635.9094, 686.1741, 527.5653, 319.2344, 137.6655, 58.22589, 
    0.5826872, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001475661, 0.08985677, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0006000945, 5.420241, 14.74992, 9.866526, 369.6528, 
    31.99669, 0, 0.6211213, 22.01926, 26.09454, 0.01676102, 0, 0, 0, 0, 0, 
    0.0003724534, 0.0007511377, 0, 0, 0, 0.01054211, 4.9378, 35.11487, 
    209.5712, 293.8589, 365.6923, 371.3261, 394.2154, 492.1788, 710.024, 
    811.8054, 617.807, 343.5852, 201.6402, 88.6078, 33.18766, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002061675, 0.3639224, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.565544, 67.44887, 210.6318, 174.2347, 0, 0, 
    0.02026485, 0.5374939, 1.169389, 0.06065548, 0, 0, 0, 0, 0, 0.0005888037, 
    0, 0, 0, 0, 0, 0, 0.1444359, 50.93018, 158.3956, 294.5731, 366.2896, 
    503.3458, 626.3784, 834.7375, 746.9637, 477.1703, 102.5894, 2.179536, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0016285, 0.005161504, 
    0, 0, 0, 0, 0, 0, 0, 0.1744462, 11.87143, 189.9295, 0, 0, 0, 0, 3.378064, 
    2.925041, 6.432992, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001116622, 
    2.862813, 19.07391, 72.97668, 86.10835, 181.0871, 146.8998, 161.6484, 
    63.05329, 18.52388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.587682e-05, 0.0007486434, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003512555, 0, 0, 0.004746107, 0, 0, 0, 0, 0, 0, 0, 0, 0.001910802, 
    1.540883, 1.139802, 0, 0, 0, 0.00339965, 0, 5.067101, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7.394003e-05, 0, 0, 0, 0, 0, 0, 0, 0.1596736, 0.01119117, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002488717, 0, 0, 0, 
    0.00192382, 0, 0.0008238192, 0, 0, 0, 0, 0.004534618, 0.01042992, 
    128.6895, 111.6004, 0.9109875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 51.51996, 6.180326, 1.820795, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001911541, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009544371, 0, 24.92486, 51.07422, 23.80963, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.353347, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 4.248243, 20.32495, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.077861e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.002998321, 0.00326913, 0, 30.07554, 20.11271, 3.618359, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1637487, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001798506, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.00186227, 0, 0.03316185, 16.06968, 162.5954, 0, 
    3.422852, 0, 0, 0, 0, 0, 0, 0, 0.01038289, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001204468, 0, 0, 0.002527093, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 66.34259, 22.89227, 15.44103, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001601016, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06553058, 0.5628351, 51.22266, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9606495, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002309131, 
    0.6115905, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.192964, 73.24959, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00447468, 0, 0, 0.001755983, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002103772, 1.21489, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 87.1916, 75.72276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.003544959, 0, 0, 0, 0, 0, 0, 0.0002654338, 0.001121242, 
    0.004204868, 0.001509032, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.04547353, 5.79191, 1.342976, 0.6890895, 0.2234796, 61.70195, 
    24.68652, 0, 0, 0, 0, 1.058887, 146.1155, 5.113419, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001511727, 0.00117502, 0.001633006, 
    0.007605216, 0, 0, 0, 0, 0, 0, 0, 0, 0.04061029, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1014451, 0, 1.253367, 0.0007692035, 16.09134, 27.76863, 48.46694, 
    11.74502, 0, 0, 0, 4.819854, 6.666916, 2.695935, 0, 0, 0, 0, 0, 0, 
    0.01972353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 202.3895,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0006035659, 0, 0, 0, 0, 0, 0, 0.01408904, 0, 
    0.003578367, 0.004032353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03354037, 0, 0, 7.591219, 30.95796, 10.42947, 11.57776, 0, 0, 0, 
    2.446361, 0.008315299, 0, 0, 0, 0, 0, 0, 0.5451445, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 120.6041, 854.0955,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001588834, 0, 0, 0, 0.005239161, 0.009033938, 
    0.0005203752, 0.001356567, 0.001431737, 0.006111554, 0, 0, 0, 0, 0, 
    0.02182276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007873155, 0, 0, 0, 0, 0, 0, 
    18.8254, 15.31145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.272007, 709.054, 928.3032,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002614032, 0, 0.007351434, 
    0.003707968, 6.454103e-05, 0.001235135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0002616841, 0, 0, 0, 0, 0, 0, 0, 0.2473145, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    463.5101, 849.1191, 684.9581,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004843049, 0.002349587, 
    0.01799333, 0.00371025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004212329, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.004271484, 0, 0, 0, 0, 0, 0, 0, 0, 57.22657, 460.95, 639.7565, 
    519.5239, 33.79907,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001354043, 0, 
    0.006613636, 0.007528742, 0.02743311, 0.01341464, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003410095, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.05400946, 4.694293, 0.3870355, 0, 0, 0, 0, 0, 141.1749, 
    601.933, 831.244, 543.7769, 58.66973, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01415738, 0.04210776, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.679655, 
    105.733, 8.447727, 0, 0, 27.24204, 24.39606, 7.753161, 352.5742, 
    608.2495, 37.65978, 0.09178872, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01123114, 0.01882986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29.1145, 27.4687, 
    38.2424, 74.43308, 193.5007, 196.5712, 7.365326, 66.00092, 2.113855, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01327394, 0.003187717, 0, 0, 0.002941251, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.80582, 
    74.16306, 226.1258, 582.3444, 525.9813, 293.4045, 129.4705, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0153161, 0.005200402, 0, 0, 0, 0.003570459, 0.002388353, 0, 0, 0, 0, 
    0.1976552, 0, 0, 0, 0.1872808, 0.7276393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3034186, 214.9815, 492.9658, 326.6951, 
    73.56389, 0.05476749, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002162333, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9388899, 
    193.1229, 6.378803, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 258.6678, 289.7753, 3.976977, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.009249282, 0.001536941, 0, 0, 0, 0, 0, 0, 0, 40.0586, 
    32.99025, 2.803985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.30081, 1.451902, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0009401445, 0.0004037078, 0, 0, 0, 0, 
    0.1391184, 50.75321, 3.125369, 1.116508, 0.2084151, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001933637, 0.05200977, 
    1.095076, 0.4746633, 0, 0.0152259, 0.00121065, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003794074, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.873821, 0, 0, 0, 
    0.0909774, 0.106935, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04739007, 0.5167308, 
    0.02355359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005289078, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0004078763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.796603,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.600741e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008196245, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2539265, 0, 
    0.1848694, 0, 0, 0, 0, 0, 0, 0.02119472, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.612157,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009860342, 0, 0, 0, 
    0.5821458, 1.014729, 1.475074, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007580966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00020889, 0.003413063, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.08453731, 0, 0.6124651, 0.0904895, 0.04531468, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.060883, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006160314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0004963353, 0, 0.002697561, 0, 0, 0, 
    0.002501344, 0.003084639, 0, 0, 0, 60.34301, 23.29774, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001295554, 0.002088146, 0, 0, 0, 0, 0.003850434, 0, 0.003216584, 
    0, 0, 6.297387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2759891, 0, 0, 0, 0, 1.456678, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002685973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.603688, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.042054e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003275427, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001260254, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004184085, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001634963, 0, 0, 0, 0, 
    0.00182365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004781314, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002623971, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1032847, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02264775, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01294437, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45.58595, 
    19.94605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01843011, 0, 0, 0, 0, 0.0006814443, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05284531, 0, 0.2416257, 0.6087035, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01169867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.009131898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006104111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002335767, 39.18405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0105723, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01319931, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1318502, 0, 0, 0.3468482, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45.02456, 0.7059237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0927918, 0.01668262, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0472814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    140.8308, 155.7868, 125.8311, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02154752, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    749.9999, 457.7867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.01483413, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.498203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002601753, 
    0.002704989, 0, 0, 0, 0, 0, 0, 0.001969324, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003557655, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02448131, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00550229, 0, 0, 0, 0, 0.0046798, 
    1.793624, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.448954, 0, 
    0.00866163, 0, 0, 0, 0, 0.4479904, 0.01966327, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005507405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.460738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03048245, 
    61.25506, 0, 0, 0, 0, 0, 0, 0.3824942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02183831, 
    0.2123545, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04637172, 
    0.008339238, 0, 0, 0.03448581, 0, 0, 0, 0, 0, 0, 0, 0.196157, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005239569, 
    0.0212123, 0.0003524371, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02602657, 
    0.02576878, 0.0369913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01774269, 
    0.006849611, 0.01812511, 0.007378699, 0.04169989, 0, 0, 0, 0.0002408772, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
