netcdf \00010101.ocean_static.dxCv {
dimensions:
	time = UNLIMITED ; // (1 currently)
	yq = 10 ;
	xh = 15 ;
	xq = 15 ;
	yh = 10 ;
variables:
	float dxCv(yq, xh) ;
		dxCv:_FillValue = 1.e+20f ;
		dxCv:missing_value = 1.e+20f ;
		dxCv:units = "m" ;
		dxCv:long_name = "Delta(x) at v points (meter)" ;
		dxCv:cell_methods = "time: point" ;
		dxCv:interp_method = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Jun 13 14:06:58 2025: ncks -d xh,532,546 -d yh,526,535 -d xq,532,546 -d yq,526,535 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.ocean_static.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.ocean_static.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 dxCv =
  26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 
    26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 
    26917.07,
  26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 
    26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 
    26946.19,
  26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 
    26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 
    26974.86,
  27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 
    27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 
    27003.08,
  27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 
    27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 
    27030.83,
  27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 
    27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 
    27058.13,
  27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 
    27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 
    27084.97,
  27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 
    27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 
    27111.35,
  27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 
    27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 
    27137.26,
  27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 
    27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 
    27162.71 ;

 time = 0 ;

 xh = -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 xq = -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 yh = -14.3476556382336, -14.1053228834302, -13.862732304759, 
    -13.6198879813569, -13.3767940148509, -13.1334545290505, 
    -12.889873669635, -12.6460556038367, -12.4020045201193, -12.1577246278516 ;

 yq = -14.4687240631789, -14.2265217428746, -13.9840595676627, 
    -13.7413416053212, -13.4983719462701, -13.2551547032665, 
    -13.011694011094, -12.7679940262485, -12.5240589266184, -12.279892911161 ;
}
