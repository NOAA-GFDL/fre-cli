netcdf atmos.1980-1981.aliq.01 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:15 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.01.nc reduced/atmos.1980-1981.aliq.01.nc\n",
			"Mon Aug 25 14:40:28 2025: cdo -O -s -select,month=1 merged_output.nc monthly_nc_files/all_years.1.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -7.363828e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0003468938, 0, 0, 0, 0, 0, 0, 0, 0, -1.015621e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -4.429732e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.763149e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.278249e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.003568112, 7.887879e-05, 0, 0, 0, 0, -1.502017e-05, 
    -9.671434e-06, 6.770824e-05, -3.427417e-05, 0, 0, -2.848659e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, -9.360258e-06, 0, 0, 0, 0,
  0, 0, -4.732072e-06, 0, 0, 0.0001513866, -5.289447e-05, 0, 0, 0, 
    -3.729734e-10, 0, 0, -2.19673e-05, -1.757202e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.946535e-05, 0, 0, 1.989067e-06, 
    7.168793e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.374052e-06, -2.769679e-06, 2.868807e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001124487, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, -8.622322e-08, 0.006046799, 0.0002231596, 0.000192132, 0, 0, 0, 
    -5.395369e-06, -7.618359e-06, 0.001193236, -1.329224e-05, 0, 0, 
    -5.082234e-05, 0, 0, 0, 0, 0, 0, 0, -8.987858e-08, 0.0009678213, 
    0.0001483564, 0, 0, 0,
  0, 0, 0.0006829959, 0, 6.047575e-05, 0.0004150458, -7.038817e-05, 
    -4.719004e-06, 0, 0, 0.0002128184, 0, 0, -3.969223e-05, -4.471886e-05, 0, 
    -8.935053e-06, 0, 0, 0, 0, 0, 0, -2.115818e-07, -1.787316e-10, 
    -3.214496e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001251601, 0, 0, -1.196803e-05, 0.00015682, 0, 
    -1.575303e-06, 7.070886e-06, 1.173033e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.235307e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001700451, 0.0003045442, 0.0001117172, 
    -1.571246e-06, 0, 0, 0.0001225012, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0002069101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4.963325e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.393176e-05, 0, 0, 0.002528994, 0, 0, 0.0003199948, 0, 
    0, 0, -3.229594e-05, 0, 0, 0, 0, 0, 0, 0, -1.182716e-05, 0, 
    -3.139127e-05, 0, 0,
  0, 0, -2.321002e-06, 0.01013409, 0.0006137282, 0.0005167123, -5.787579e-06, 
    0, 0, 0.0003318985, 0.0006363702, 0.002296257, 0.0006888872, 0, 0, 
    0.0003382304, -4.22391e-05, 2.848217e-06, 0, 0, 0, 0, 0, -2.696357e-07, 
    0.002563883, 0.0003047311, 0, 0, 0,
  0, 0, 0.0009373818, -1.787363e-05, 0.000108785, 0.001488058, -0.0001374804, 
    -8.223637e-05, 0, 0, 0.0004235709, 0, 0, 0.0009883444, -4.58297e-05, 
    0.0009350691, 0.0001705676, 0, 0, 0, 0, 0, 0, -2.547138e-07, 
    6.356565e-05, 0.0004062194, 0, 0, 0,
  0, 0, 0, 0, -1.402646e-10, -1.530469e-05, 0.0008158231, 0, 0, 
    -3.232031e-05, 0.0008343049, 0, 0.000326232, 0.001703776, 0.001953145, 0, 
    -8.089992e-06, 0, 0, 0, 0, 0, 0, 0, -3.837726e-06, -3.548382e-05, 0, 0, 0,
  0, 0, 0, 0, 0, -1.152974e-05, 0, -3.051627e-06, 0, 0.0003390776, 
    0.0003756555, 0.0008293684, 0.0009214346, -1.10305e-05, 0, 0, 
    0.001130976, 0, 0, 0, 0.0005184304, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.00199725, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008817194, -3.826602e-06, 0.0008132577, 0, 0,
  0, 0, -9.666323e-07, -2.400689e-06, 0, 0, -4.665617e-05, 0, 0, 0.003927528, 
    0, 0, 0.0007978121, -4.431036e-06, 0, 0, 0.000702787, 0.001156713, 
    -4.828374e-08, 0, 0, 0, 0, 0, 5.27481e-05, -2.153833e-06, 0.0001126413, 
    0, 0,
  0, -2.920995e-05, 5.338054e-05, 0.01184445, 0.0007747919, 0.002268009, 
    0.001001507, 0, 0, 0.001849305, 0.001288586, 0.00319184, 0.001964029, 
    0.0003786287, 0, 0.001722791, 0.0004279665, 0.0004207391, 0, 0, 0, 0, 0, 
    -2.986008e-06, 0.005601919, 0.001302016, 0, 0, 0,
  0, 0, 0.002123553, -5.376404e-05, 0.0001731613, 0.002991819, 0.0003858407, 
    -0.0002085071, 0, 0.0003325184, 0.001742656, 0.0002579924, -1.965447e-05, 
    0.002617273, 5.976149e-05, 0.001693348, 0.0009333555, 2.089505e-05, 0, 0, 
    0, 0, 0, -6.728231e-06, 0.001016685, 0.002270084, 0, 0, 0,
  0, 0, 0, 0, -3.19703e-10, -4.649825e-05, 0.002818835, 0, -8.180113e-06, 
    0.000231508, 0.001814359, 0, 0.003749661, 0.007861725, 0.008525283, 
    7.207104e-05, -2.53004e-05, 0, 0, 0, 0, 0, 0, -1.928245e-06, 
    7.754003e-05, 0.0004553747, 0, 0, 0,
  0, 0, 0, 0, 0, -4.058285e-05, 0, 0.0007014206, 0, 0.000675004, 
    0.0008600135, 0.002141407, 0.002157426, 0.001859099, 0, -3.261727e-05, 
    0.002270703, 0, -1.178809e-05, 0, 0.002302204, -1.921128e-05, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.389488e-06, 0, 0, 0,
  0, 0, 0, 0.005597793, 0.0004557264, 0.0006469226, 0, 0, 0, 0, 0, 0, 
    5.932737e-05, 0, 0, 0, -9.95197e-06, -9.82077e-07, 7.914577e-05, 
    -9.838413e-06, 0, 0, 0, 0, 0.001656214, 0.0008312016, 0.002270857, 0, 0,
  0, 0, -1.700663e-06, 0.0007984373, -3.725525e-05, -9.926032e-06, 
    0.002917385, 0, 0, 0.005295489, 0, 0, 0.001142852, -1.550863e-05, 
    -4.614825e-06, -9.7571e-05, 0.003277591, 0.003097947, -9.88366e-07, 0, 0, 
    0, 0, 0, 0.0001335976, -2.301468e-05, 0.0008439922, 0, 0,
  0, 0.0006595507, 0.0001256985, 0.0172606, 0.002429031, 0.004938448, 
    0.00146689, 0, 0, 0.004881167, 0.002610792, 0.006603616, 0.004202751, 
    0.0008606157, -1.021467e-05, 0.002467264, 0.0009008423, 0.001963713, 
    0.0005992454, 0, 0, 0, 0, -1.340549e-05, 0.009736534, 0.00386131, 
    0.0003141004, 0, 0,
  0, 0, 0.00465352, 0.0001797527, 0.002113543, 0.004013491, 0.0008106963, 
    -9.982745e-05, -7.495759e-06, 0.001494612, 0.003723009, 0.001112406, 
    -6.828645e-06, 0.003211215, 0.001124431, 0.002775689, 0.002879745, 
    4.865911e-05, 0, 0, 0, 0, 0, 2.950077e-06, 0.002990948, 0.003281872, 
    9.949968e-05, 0, 0,
  0, 0, 0, 0, 1.33027e-05, 0.0002379751, 0.007269307, 3.319753e-06, 
    0.0002124923, 0.00245001, 0.005283603, 0.000213335, 0.006571532, 
    0.01612738, 0.01339556, 0.001426343, -3.8621e-05, 0, 7.179433e-05, 0, 
    -1.028143e-05, 0, 0, -1.928245e-06, 0.000283097, 0.003553868, 
    -8.445634e-06, 0, 0,
  0, 0, 0, 0, 0, -0.0001103674, 0, 0.00100146, 0, 0.0007924786, 0.004844656, 
    0.005290551, 0.00434326, 0.003626761, -2.220837e-07, -0.0001309093, 
    0.004720834, -1.85161e-05, -5.774866e-05, -4.702264e-05, 0.005721793, 
    1.41119e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -2.390274e-06, 0, 0, 0, 0, 0, 0, 0, 0, -7.872414e-05, 
    -5.887881e-06, 0, 0, -1.693163e-05, 0, 0, 0, 0, 0, 0, 0, -2.218284e-05, 
    -2.200381e-05, 0, 0,
  0, 0, 0, 0.008799365, 0.006159117, 0.004396006, -1.909977e-05, 0.001149741, 
    0, 6.007154e-05, 0, 0.0009088502, 0.002814545, 0.0001919991, 
    -6.663022e-07, 0, 3.200075e-05, 0.000591276, 0.001719561, -0.000179826, 
    0, 0, 0, 0, 0.002777288, 0.00366555, 0.006712748, 0.0006813456, 0,
  0, 0, -9.242537e-06, 0.003332648, 0.0002176759, -0.0003034646, 0.006001565, 
    0, 0, 0.006093781, 0, -5.891067e-06, 0.00252047, -4.900837e-05, 
    -0.0001118976, 0.000847741, 0.007361409, 0.00662106, -1.067203e-05, 0, 0, 
    0, 0, 0, 0.0005522493, 0.0004619156, 0.002976233, 0, 0,
  0, 0.002107489, 0.0001728124, 0.02428266, 0.00914899, 0.008797932, 
    0.005174937, 0, 0, 0.01020808, 0.004488002, 0.01310519, 0.00936108, 
    0.001116405, 0.0007504203, 0.01268706, 0.0055054, 0.005009706, 
    0.002733892, 0, 0, 0, 0, -3.188773e-05, 0.0157695, 0.005852027, 
    0.001693417, 0, 0,
  0, 0.0002322066, 0.008308734, 0.0004423383, 0.004081899, 0.004973883, 
    0.002320526, 0.0004445713, 0.0001499184, 0.005659968, 0.005618632, 
    0.002376017, 0.0003356724, 0.004721674, 0.004418676, 0.003818574, 
    0.006651992, 0.0001667552, 0, 0, 0, 0, 0, -4.096237e-05, 0.006630517, 
    0.005466895, 0.0003398354, 0, 0,
  0, 0, 0, 0.0001270712, 0.0005868991, 0.002004822, 0.01727506, 0.0002414046, 
    0.001915593, 0.007482093, 0.009087131, 0.0007285787, 0.00949965, 
    0.02510638, 0.02100114, 0.003215773, 9.631445e-05, -2.403638e-05, 
    0.0007701347, 0, -1.434231e-05, 0, 0, 0.0001784717, 0.0002952538, 
    0.01033398, 0.001699082, 0, 0,
  0, 0, 0, 0, -1.700727e-06, -6.085856e-05, 0, 0.00210834, 0, 0.001851091, 
    0.006980861, 0.008608033, 0.007395587, 0.00567356, -1.577238e-05, 
    0.0002305305, 0.01003598, -8.20393e-05, 0.0006473598, -8.201694e-05, 
    0.01186063, 0.001304529, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0001979469, 0, 0, 0, 0, 0.001676462, 0, 0, 0, 0, 0, 
    0, -9.146282e-06, 0, -2.885683e-05, 0, 0, 4.676857e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.535969e-07, 0, 
    0.0005790186, 0, -1.752291e-05, 0, 0, 0, 0, -2.202491e-06, 2.795208e-05, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.26666e-05, 2.925535e-05, 0.0004111773, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.063926e-06, 0, -2.877666e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.435464e-05, 0.0002013601, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0004288905, 0.001309462, 0.002350187, -1.39765e-05, 0.001901275, 
    0.0009352251, 0, 0, 0, 0, 0.004055185, 0.001013167, 3.759666e-05, 0, 
    0.0002124368, 0.000851781, 0.0007544663, 0, -6.334013e-07, 0, 0, 0, 
    6.584295e-05, 0.003555404, 0.0001488428, -8.480972e-07,
  0, 0, 0, 0.01291051, 0.0118, 0.008277914, -7.988459e-05, 0.002282832, 0, 
    0.001621236, 0, 0.00353805, 0.005957454, 0.001885002, -6.642054e-06, 
    -2.503222e-05, 0.003038786, 0.002283092, 0.01173666, -0.0002643683, 0, 
    -5.391511e-06, 0, 0, 0.006194122, 0.01564369, 0.01370825, 0.001595638, 
    0.0005618859,
  0, 0, 0.0002515629, 0.007660474, 0.004404311, 0.003701776, 0.01049482, 0, 
    0, 0.006817032, -1.096249e-05, 2.352893e-06, 0.01143608, 0.0002186215, 
    -4.218977e-05, 0.004671329, 0.01896391, 0.01448526, 0.0009912279, 0, 0, 
    0, 0, 0, 0.005753408, 0.005938749, 0.01522681, 0, 0,
  0, 0.004060008, 0.001524845, 0.03195173, 0.02478782, 0.01126469, 
    0.01468937, -3.817516e-06, 0, 0.02608612, 0.009733162, 0.02770602, 
    0.02249338, 0.004246153, 0.002540812, 0.0394203, 0.0184706, 0.01157512, 
    0.004760633, 0, 0, 0, 0, 0.001230321, 0.02993653, 0.01422851, 
    0.005861097, 0, 0,
  0, 0.0008920152, 0.01688166, 0.003931677, 0.01759309, 0.0130573, 
    0.01448352, 0.002855443, 0.00164686, 0.01154009, 0.008888641, 
    0.005667158, 0.003624117, 0.01252668, 0.01214778, 0.008533034, 
    0.01530576, 0.001025702, 0, 0, 0, 0, 0, 0.0007823122, 0.0136766, 
    0.01749676, 0.00229054, 0, 0,
  0, 0, 0, 0.0002235279, 0.003137773, 0.008499213, 0.04070725, 0.001861471, 
    0.002765811, 0.01607794, 0.01448523, 0.001614236, 0.0143179, 0.04112271, 
    0.03288089, 0.006545304, 0.0009808616, 6.170331e-05, 0.002330611, 0, 
    0.000443328, 0, -3.167048e-06, 0.0008587094, 0.0007761889, 0.02261324, 
    0.004774569, 0, 0,
  0, 0, 0, 0, -5.208502e-05, 0.000305724, -3.471439e-05, 0.006974578, 0, 
    0.002949034, 0.01312773, 0.01651449, 0.01416429, 0.01116141, 
    -0.0001445699, 0.001817385, 0.01599235, 0.002568282, 0.002683438, 
    0.001003487, 0.02240447, 0.002654123, 0, -7.748087e-07, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -7.032821e-10, 0.001420722, 0, 0, 3.634102e-05, 
    -1.063763e-05, 0.003318012, 0, 0, 0, -1.334631e-09, -3.042314e-06, 0, 
    0.000290718, 3.926469e-05, 0.0002325321, 0, 0, 0.0004391529, 
    -1.847406e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.28314e-06, 6.552266e-05, -2.19275e-09, 
    -3.13811e-06, 0, 0.0004402956, 2.933839e-05, 0.00291027, 0, 0.001208002, 
    0, 0, -1.274065e-05, 3.240932e-05, -4.616169e-05, 0.001217858, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.018551e-07, 0, 0.0005245823, 
    0.0002819446, 0.0001108126, -1.982711e-05, -1.609767e-05, 0, 0, 
    0.0003476821, -3.813735e-05, 0.002497325, 0.004546024, 4.443499e-05, 
    -8.084766e-06, -1.310791e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.575638e-06, 
    -2.636101e-06, 0, 0, 0, 0, 0, 0, 0.0001978852, 0.0008492544, 
    -2.295522e-05, 0.0003140819, -6.044327e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.203366e-10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -5.033492e-07, 0, 0, 0, -4.559039e-05, -1.431388e-05, 6.531667e-06, 
    0, -3.756159e-10, 0, -6.149552e-05, 0.003165124, 0.001563917, 
    3.927744e-06, 0, 0, 0, 0, 0, 0, -1.086994e-05, 0, 0, 0, -1.024639e-05, 0, 0,
  0.00188791, -1.214084e-05, -1.119997e-06, 0.000607691, 0.002286286, 
    0.006530093, -2.339476e-05, 0.002302676, 0.001983813, -1.297806e-06, 0, 
    -6.639202e-06, -6.106782e-06, 0.01590675, 0.00179717, 0.001280956, 
    -2.141584e-05, 0.002631821, 0.002182493, 0.002624875, 0.0008556225, 
    0.0002026056, -3.734986e-05, 0, 0.0002381313, 0.003176087, 0.01213867, 
    0.001551016, 0.001417568,
  -1.272196e-05, -9.134666e-06, -2.574806e-08, 0.01717869, 0.01621988, 
    0.0172693, 0.0008246354, 0.002638177, -1.368142e-06, 0.002797607, 
    -1.447551e-05, 0.00677767, 0.01067174, 0.005379904, 0.0004746295, 
    0.0008781806, 0.009269753, 0.00659386, 0.0380741, 0.005548884, 
    0.0002295577, 0.0003158493, 0, -7.331432e-06, 0.01402885, 0.03653747, 
    0.02539841, 0.002665297, 0.001303855,
  0, -6.761459e-07, 0.004300587, 0.01620743, 0.0131489, 0.03602235, 
    0.01494452, 5.455871e-05, -2.313185e-06, 0.007822813, 0.0003808359, 
    0.001488909, 0.02495853, 0.0004939489, 0.0007085892, 0.01548787, 
    0.02650461, 0.02865112, 0.01094651, -2.077551e-09, 0, 0, 0, 0, 
    0.01186294, 0.01676278, 0.04063754, 2.694851e-05, 0,
  0, 0.008221603, 0.008075677, 0.04260761, 0.04358185, 0.02591865, 
    0.03128107, -6.553076e-05, 0, 0.0436923, 0.0225311, 0.06374897, 
    0.04930611, 0.01451654, 0.006669693, 0.06287394, 0.04460896, 0.02149856, 
    0.007624072, 0, 0, -3.414575e-09, 2.188752e-07, 0.006622558, 0.07618755, 
    0.02920797, 0.01172381, 2.459115e-05, 0,
  0, 0.001968135, 0.0410899, 0.01213883, 0.04418617, 0.0272984, 0.03102343, 
    0.01668715, 0.009160494, 0.02304175, 0.01547701, 0.01366172, 0.01720015, 
    0.0317632, 0.04893946, 0.02040784, 0.02998321, 0.001722667, 
    -9.326763e-06, 0, 0, 0, -3.100153e-07, 0.01705568, 0.06041917, 
    0.03346419, 0.006739568, -5.095661e-10, 0,
  0, 0, 2.713305e-06, 0.0002779756, 0.01309681, 0.02274185, 0.0827126, 
    0.003860528, 0.008320999, 0.03667165, 0.02197314, 0.006584266, 
    0.03414353, 0.06435549, 0.05250769, 0.0101376, 0.002070946, 0.001671073, 
    0.004475679, -3.651543e-08, 0.003258094, -7.06663e-08, 0.000432825, 
    0.00401489, 0.002741714, 0.03855168, 0.009472364, -1.193373e-09, 
    -2.811552e-11,
  -3.719376e-10, 0, 0, 0, 0.001023703, 0.00317339, -6.808838e-05, 0.0167546, 
    -1.903902e-05, 0.003939449, 0.02781136, 0.03998166, 0.03545783, 
    0.01518598, -3.138775e-05, 0.002899046, 0.02644938, 0.01099012, 
    0.005449621, 0.006150124, 0.03528051, 0.004894046, 1.166943e-06, 
    -7.061622e-06, 7.422087e-10, 5.803029e-10, -9.199943e-09, -1.932743e-07, 
    -1.419027e-07,
  0, 0, 0, 0, 0, 0, 2.769583e-05, 0.003284464, 4.652442e-07, 0, 0.0004003473, 
    0.0007296901, 0.005268937, 0, 0, -1.838574e-08, 2.743901e-05, 
    0.001673598, 0.0002759735, 0.008242704, 0.004653784, 0.003285551, 
    -8.39374e-05, 4.288099e-09, 0.002647221, 6.816295e-05, 6.999794e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001316631, 0.0007930074, -4.728162e-05, 
    -4.0098e-05, 0.0002620381, 0.001770798, 0.005816514, 0.004957795, 
    0.0001064483, 0.00315181, 0, 0, 0.0005131187, 0.0001225484, 0.0008394819, 
    0.001969537, 0, 0,
  0.0005223778, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.120952e-05, 0.0008655902, 
    0.0003674998, 0.002034194, 0.001220577, 0.004021717, 0.003300464, 
    0.00059609, 0, -7.130092e-06, 0.001448565, 0.000872827, 0.007284674, 
    0.01200688, 0.002186904, -4.063599e-05, 0.002592757,
  4.634277e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006726474, 
    0.00133906, -1.287994e-05, -1.230323e-05, 0, 0, 0, -3.671121e-05, 
    0.001036416, 0.001740289, 0.00107387, 0.002982258, 0.001213497,
  0, -1.014022e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0009471958, -6.427023e-06, -7.513584e-06, 0, 0, -6.876646e-06, 
    0.001884265, 0.001576885, 0.001700105, 1.329634e-09, 2.561414e-05, 0, 
    0.000472904, 0.005446059, 0.003895383, 0.0002607964, -8.964251e-05, 
    0.001377806, 0, -5.942783e-06, -2.208756e-05, 0, -3.003725e-05, 
    -2.856407e-05, 4.913288e-06, -7.154569e-06, 0.001347899, 0, -6.037531e-06,
  0.006256233, 0.002729879, -1.925045e-05, 0.003077442, 0.006156206, 
    0.02250919, 0.006269827, 0.00572917, 0.002948351, 0.00414324, 
    1.712975e-08, 0.000143901, 0.001115752, 0.03691888, 0.009285406, 
    0.003253025, 0.001354098, 0.01028166, 0.006734345, 0.01038897, 
    0.006529666, 0.0005370149, 0.0007418901, 4.826718e-06, 0.00223055, 
    0.008858554, 0.01964253, 0.01101734, 0.01353479,
  2.715114e-05, 0.001096595, 0.0001563805, 0.02524484, 0.02745131, 
    0.02915035, 0.008346973, 0.003568372, 0.0005049725, 0.004602478, 
    0.0006997266, 0.01308617, 0.02322404, 0.01353621, 0.003412774, 
    0.004465615, 0.01764099, 0.01229853, 0.06248029, 0.0199532, 0.001508894, 
    0.0006393534, 0.001113706, -1.877746e-05, 0.02270375, 0.06164753, 
    0.0482904, 0.0161912, 0.002508074,
  4.010976e-10, 4.522981e-05, 0.01271263, 0.04613801, 0.03412648, 0.06460659, 
    0.02145966, -4.138818e-05, 0.0003245437, 0.01531032, 0.0153675, 
    0.003279734, 0.03933674, 0.005361534, 0.002075593, 0.02789375, 
    0.04363402, 0.05519388, 0.03877128, 0.0001691224, -3.489269e-05, 0, 0, 
    6.024018e-05, 0.04279283, 0.04486388, 0.07637952, 0.0001529095, 
    1.929693e-05,
  0.0002886714, 0.0323687, 0.04163257, 0.09358516, 0.08102733, 0.09089021, 
    0.06720141, 0.00304821, 0.000614342, 0.07918452, 0.1245744, 0.1902409, 
    0.186048, 0.1063229, 0.03627665, 0.1458589, 0.1365699, 0.0409823, 
    0.01348407, 0.0005757593, 2.690589e-07, 0.0002710439, 0.00169743, 
    0.1222184, 0.3289421, 0.05024547, 0.01522701, 0.0001096268, -7.31107e-09,
  1.073939e-05, 0.004251658, 0.08181123, 0.03458502, 0.09296998, 0.07784823, 
    0.06522873, 0.07415938, 0.04517638, 0.1503089, 0.08577977, 0.1217666, 
    0.1659401, 0.1216394, 0.1809303, 0.13786, 0.07068841, 0.002665454, 
    0.0006942449, 3.79595e-05, 0, 7.752262e-07, 0.009291851, 0.1244161, 
    0.2688979, 0.0839016, 0.017748, 0.0006260531, -1.754799e-08,
  1.347913e-06, 2.496997e-06, 0.0002034639, 0.0006512611, 0.01893885, 
    0.03797341, 0.1401755, 0.03479271, 0.03042937, 0.1034123, 0.06138936, 
    0.1123767, 0.1487229, 0.1579317, 0.1196513, 0.03581021, 0.002197, 
    0.007600519, 0.007824407, 1.155389e-05, 0.008166974, -9.83248e-07, 
    0.004159718, 0.03708261, 0.02047454, 0.06378637, 0.01565097, 
    0.0005256005, 8.141821e-07,
  -9.92879e-08, 0, 1.565583e-06, 0, 0.001890573, 0.007229572, 0.0003727242, 
    0.02994307, 0.0004658431, 0.01723977, 0.07570474, 0.09567214, 0.1381414, 
    0.04499653, 0.00696663, 0.003620686, 0.03733719, 0.02813025, 0.01205452, 
    0.01903238, 0.04791149, 0.008714895, -1.393793e-05, -2.467677e-05, 
    0.001038319, 0.0004630347, 3.979263e-06, 0.0002876333, 0.0001502035,
  -1.134409e-08, -2.258256e-06, 0, 1.433293e-08, 0, -1.452074e-08, 
    0.0005057755, 0.00452818, 1.362122e-05, 1.947733e-07, 0.0005710463, 
    0.01512128, 0.01964078, 8.42487e-06, 3.122377e-07, 1.343964e-06, 
    0.002796723, 0.01018328, 0.006389828, 0.02127879, 0.01919933, 0.02086694, 
    0.001853333, 6.774614e-06, 0.004067716, 0.002195976, 1.174423e-07, 
    4.827692e-05, -9.416162e-06,
  0, 0, -4.095626e-09, -2.743774e-12, 0, -2.285931e-11, -1.857506e-05, 0, 0, 
    4.506017e-09, 3.782384e-09, 0.004791297, 0.004814559, 0.002612155, 
    0.002083324, 0.007237266, 0.006414196, 0.02740832, 0.0105211, 
    0.003652391, 0.007437212, 0.005542523, 0.004527877, 0.001951542, 
    0.004398938, 0.01445628, 0.007764956, -5.558812e-06, 0,
  0.002115848, 0, 0, 0.0001374153, 0, 8.936191e-05, 0, 0, 0, 0, 0, 
    -4.283215e-06, 0.0007571002, 0.002735747, 0.003942533, 0.005752774, 
    0.003785014, 0.02201899, 0.007192052, 0.001849515, -2.588595e-05, 
    0.0006112481, 0.004844327, 0.005242415, 0.01312883, 0.0322785, 
    0.01701964, 0.003071898, 0.004995045,
  2.538158e-05, 0.0002340322, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.061986e-06, 
    0, 6.177595e-06, 0.003413268, 0.002359205, 0.0003738367, -6.636724e-06, 
    -4.533502e-09, 0, 0, -2.130328e-05, 0.003700576, 0.003102654, 
    0.003553787, 0.006356281, 0.004335555,
  0, 0.00134468, -2.112188e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005358549, -6.683946e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.000997258, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0001199418, 0, 0, 0, 0, 0, -5.311483e-06, -2.215619e-05, -1.963213e-11, 
    0, 0, 0, -6.550339e-05, 0, 0, -8.787697e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0009216329, 0.00190932,
  0.003375014, 0.0007291378, 1.98828e-05, 0, 0.00223299, 0.004981244, 
    0.01637407, 0.01239625, 0.008015514, 0.0003100034, 0.000782292, 0, 
    0.002622253, 0.008371696, 0.01643549, 0.004000307, 0.0008738641, 
    0.004702229, 0.0004752304, -0.0001781599, -6.912409e-05, 0, 0.001955597, 
    0.001088444, 0.002121716, 0.000293292, 0.002824618, 0.001389146, 
    0.0006160659,
  0.0133168, 0.007339987, 0.001506114, 0.009851512, 0.01835279, 0.05187973, 
    0.02854934, 0.03138807, 0.009912244, 0.0142956, 0.001048844, 
    0.0004306328, 0.009990805, 0.07306478, 0.03312182, 0.01225997, 
    0.01412344, 0.02280393, 0.02143044, 0.01857488, 0.02912308, 0.00929046, 
    0.008285934, 0.004035871, 0.007234339, 0.01617297, 0.02620247, 
    0.02517242, 0.02218344,
  0.008704777, 0.006317859, 0.007404099, 0.04549472, 0.05233592, 0.0757601, 
    0.0415123, 0.0201163, 0.004726769, 0.02005781, 0.02666514, 0.05181832, 
    0.05831423, 0.04863738, 0.008140372, 0.01751011, 0.04550337, 0.03528022, 
    0.1082981, 0.05189817, 0.02086193, 0.002568241, 0.002804319, 
    -4.364269e-05, 0.03102881, 0.09249233, 0.0820928, 0.06763879, 0.02527635,
  0.001947212, 0.004499737, 0.08308093, 0.08236634, 0.1073781, 0.1289135, 
    0.06663036, 0.03795868, 0.01944477, 0.02976254, 0.0705282, 0.03969714, 
    0.07584533, 0.07585388, 0.06471739, 0.0735368, 0.1402916, 0.1950899, 
    0.1963969, 0.02411109, 0.001147513, -4.80042e-06, 4.630513e-06, 
    0.004658292, 0.1059997, 0.1832298, 0.1914588, 0.01772809, 0.001133311,
  0.002687396, 0.1146839, 0.1956196, 0.1067159, 0.1154917, 0.1573832, 
    0.1377623, 0.01156905, 0.000288618, 0.06037692, 0.1385062, 0.1977267, 
    0.2111434, 0.1811671, 0.07529492, 0.1780163, 0.2240902, 0.1729099, 
    0.1569968, 0.01338119, 0.0004769176, 0.0002039586, 0.01219348, 0.122711, 
    0.3089781, 0.2032854, 0.08083265, 0.03017577, 0.006638217,
  0.002132878, 0.04577326, 0.4221116, 0.2017719, 0.199355, 0.1807576, 
    0.1478525, 0.08838469, 0.05859619, 0.147349, 0.09727162, 0.1026422, 
    0.1316231, 0.1050197, 0.1565071, 0.1326364, 0.1140696, 0.01866388, 
    0.02297446, 0.00596379, -9.740726e-06, 1.182217e-05, 0.03404658, 
    0.4377522, 0.4104794, 0.3030963, 0.1697582, 0.01503223, 0.01128281,
  0.0001779015, 0.01034575, 0.03354757, 0.03263598, 0.0943784, 0.1363139, 
    0.262906, 0.1260363, 0.1737905, 0.3276539, 0.1100295, 0.1541058, 
    0.1545636, 0.1527393, 0.1230688, 0.04047669, 0.0008962749, 0.007832065, 
    0.01759075, 0.0003315854, 0.007076874, 3.242826e-05, 0.01240777, 
    0.3030446, 0.2836206, 0.2071944, 0.07175671, 0.01739367, 0.02136024,
  2.834942e-05, -1.289819e-05, 6.983487e-05, -2.966803e-06, 0.003326783, 
    0.02379945, 0.02007337, 0.05921026, 0.003528422, 0.08454019, 0.09344787, 
    0.1038669, 0.1309367, 0.04398722, 0.00411418, 0.01396133, 0.06054679, 
    0.04768109, 0.03586548, 0.1139297, 0.1393469, 0.01884073, 0.002455839, 
    0.00819089, 0.007716572, 0.0007329757, 0.002981514, 0.02122492, 
    0.001482272,
  0.001070985, 2.037733e-05, 5.615251e-07, 2.271474e-06, 1.464511e-05, 
    2.86162e-05, 0.001065404, 0.005774167, 0.0006176637, 3.952619e-06, 
    0.004023747, 0.01455884, 0.02427716, -1.306965e-05, 8.459724e-07, 
    0.0003074897, 0.01411747, 0.05443445, 0.04238234, 0.06380294, 0.1861721, 
    0.07790311, 0.02018164, 0.0008584389, 0.013213, 0.006899842, 
    6.696806e-06, 0.003302317, -5.325795e-05,
  0, -1.132546e-06, 0.0001088122, 7.297826e-05, 2.959738e-05, 0.0001241949, 
    -0.0001045731, 0, 0, 1.714915e-07, 1.076569e-05, 0.01066657, 0.02731106, 
    0.01341423, 0.007534636, 0.01376035, 0.01769948, 0.0555061, 0.02506317, 
    0.01234377, 0.02185007, 0.01788435, 0.01307316, 0.01135148, 0.0174829, 
    0.03882445, 0.01903943, 6.500313e-05, 0.0001786385,
  0.006269428, 0.0007840529, 9.525343e-08, 0.0009378352, -0.0001446128, 
    0.0007102559, 0, 0, 0, 0, 0, 0.001408218, 0.003054325, 0.007823321, 
    0.01033054, 0.01127218, 0.03039812, 0.04049686, 0.02078179, 0.006174399, 
    0.001063313, 0.002767914, 0.008307541, 0.01311743, 0.02160737, 
    0.06274127, 0.05095809, 0.01177819, 0.009008515,
  0.002101424, 0.001258917, 9.372061e-05, -4.421062e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.485212e-05, 0, 0.002183987, 0.009030178, 0.007454195, 
    0.004911348, 0.0006090308, -3.756178e-05, 0, 0, 0.000796715, 0.006013726, 
    0.009183504, 0.009604692, 0.01355145, 0.01381881,
  0.0006652151, 0.002401232, 1.197897e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -5.398118e-06, 0, 0, 0, 0, 0, 0, 1.111379e-05, 0.001711095, 0, 
    0.002171072, 0.0004816722,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005060422, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.342868e-06, -5.222323e-07, 
    -6.453587e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.004430693, 0.0005479861, 0, 0, -1.266481e-09, 0, 0.003236752, 
    -0.0001346003, -1.532055e-05, 0, 0, 0, 0.0004890886, 0.0003722121, 
    0.0001231043, 0.003650929, 0.002321318, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002138227, 0.003158528, 0.002863511,
  0.007209599, 0.004109026, 0.001254328, 9.967558e-06, 0.00731212, 0.0139764, 
    0.02644116, 0.02065018, 0.02420028, 0.008631475, 0.001694541, 
    0.0001286107, 0.005352406, 0.01211887, 0.04450588, 0.03597797, 
    0.02317183, 0.01582115, 0.005588198, 0.002970822, 7.426888e-05, 
    -2.001701e-05, 0.00439673, 0.007975184, 0.003846204, 0.001340401, 
    0.008328276, 0.006544347, 0.005537989,
  0.0436681, 0.02617557, 0.0193359, 0.03841215, 0.08420749, 0.09280263, 
    0.07432471, 0.05669152, 0.04272824, 0.03272229, 0.004976822, 0.001960161, 
    0.02879699, 0.1405609, 0.1000019, 0.06463315, 0.05230381, 0.0717196, 
    0.05553071, 0.04794563, 0.0728426, 0.07157601, 0.0370783, 0.01810477, 
    0.01547947, 0.03281774, 0.04415475, 0.05576305, 0.06297401,
  0.03399134, 0.02873229, 0.03102423, 0.07914808, 0.09454804, 0.1023248, 
    0.06334942, 0.03987255, 0.05292287, 0.04756116, 0.06550229, 0.119159, 
    0.1330502, 0.1328706, 0.05110174, 0.04991601, 0.1122042, 0.08248508, 
    0.164377, 0.1571657, 0.08974653, 0.04313264, 0.04395597, 0.002041748, 
    0.05715948, 0.1369531, 0.1387528, 0.1525732, 0.07246195,
  0.001518088, 0.00443065, 0.1148195, 0.07840942, 0.1059475, 0.1502604, 
    0.1245799, 0.04309022, 0.02194395, 0.04584453, 0.078146, 0.04722638, 
    0.1043962, 0.1046121, 0.08406641, 0.08557395, 0.1364999, 0.1897222, 
    0.2399849, 0.1206634, 0.06281021, 0.01314697, 2.966687e-05, 0.005825187, 
    0.09818245, 0.1781203, 0.2378997, 0.048466, 0.0172487,
  0.0008498117, 0.08863771, 0.1598721, 0.0960336, 0.09677615, 0.129979, 
    0.1132719, 0.007754366, 0.0001001746, 0.05032725, 0.1248729, 0.1699728, 
    0.18422, 0.1361405, 0.06143617, 0.1558712, 0.1872237, 0.14419, 0.1358438, 
    0.04962311, 0.03364092, 1.557104e-06, 0.001977327, 0.1036953, 0.2633385, 
    0.182545, 0.07289284, 0.04120146, 0.02555897,
  0.0002181464, 0.0333558, 0.3857112, 0.1498656, 0.1700985, 0.1294376, 
    0.1141185, 0.06290544, 0.043284, 0.1258984, 0.06809701, 0.07786931, 
    0.08322112, 0.08384769, 0.1247319, 0.09590554, 0.09089333, 0.01183434, 
    0.01669133, 0.01015509, -2.661699e-05, 2.878233e-06, 0.02002313, 
    0.4102502, 0.3723972, 0.2728509, 0.1322675, 0.01366403, 0.009714358,
  0.0002634172, 0.004099643, 0.007102196, 0.02803793, 0.0552854, 0.09315444, 
    0.2327495, 0.09963238, 0.1243376, 0.2734051, 0.08811762, 0.1187927, 
    0.1213913, 0.1196584, 0.1029574, 0.03306621, 0.000419843, 0.001174839, 
    0.01098627, 0.0001870442, 0.006196529, 0.002116713, 0.007253203, 
    0.1966617, 0.223187, 0.1826456, 0.04788091, 0.02777375, 0.0193013,
  0.008126521, 1.43973e-05, 2.00141e-05, 1.202397e-05, 0.0008951396, 
    0.01433455, 0.01423256, 0.04702499, 0.001817613, 0.06312099, 0.07347358, 
    0.07568518, 0.1055243, 0.03149614, 0.002621862, 0.01056404, 0.05076384, 
    0.0401838, 0.02258805, 0.07945494, 0.1043891, 0.01562235, 0.000453466, 
    0.005627022, 0.00262557, 8.011824e-05, 0.00493632, 0.04460274, 0.1296141,
  0.250131, 0.01049199, 0.0001548362, 2.144135e-07, 1.766986e-06, 
    4.343626e-06, 0.0006396047, 0.007555921, 0.008954842, 0.0002751619, 
    0.004103308, 0.01104054, 0.02272168, 1.740006e-05, 1.321033e-05, 
    0.0005324734, 0.03388581, 0.08963034, 0.04486811, 0.1136909, 0.1792896, 
    0.08106708, 0.01124065, 0.00678244, 0.02717548, 0.01838112, 0.01700608, 
    0.023554, 0.09293951,
  4.654201e-05, 0.0159054, 0.01594088, 0.003409169, 0.001282404, 
    0.0004792451, 0.001907458, -6.621352e-07, 1.651863e-07, 0.008385498, 
    0.005312202, 0.01691411, 0.05104389, 0.02410524, 0.02497673, 0.0287141, 
    0.0387802, 0.1090179, 0.09370622, 0.03795646, 0.04430027, 0.07469909, 
    0.04899503, 0.05165808, 0.09143131, 0.1017167, 0.09138137, 0.005844979, 
    0.001502011,
  0.01381768, 0.006098577, 0.0006765461, 0.003737005, 0.0001379947, 
    0.001132932, 5.898153e-05, 0, 0, 0, 0, 0.00194421, 0.009718604, 
    0.01714838, 0.02520961, 0.03308769, 0.07267911, 0.07243662, 0.05241084, 
    0.01904103, 0.00202663, 0.006861218, 0.02335125, 0.03092427, 0.03763115, 
    0.09037925, 0.1016182, 0.04381663, 0.01589143,
  0.01199942, 0.00259218, 0.002776006, -9.775947e-06, -7.024351e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0003365543, -5.17838e-05, 0.004013315, 0.01758737, 
    0.01676235, 0.01521643, 0.001432276, 0.0002825548, 0, -1.185466e-05, 
    0.001612067, 0.0116604, 0.02033586, 0.0251875, 0.03460424, 0.03429183,
  0.003862982, 0.003150466, 0.0006123242, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.862867e-07, 1.066617e-06, -1.838148e-05, 0.0007872349, 9.04966e-05, 
    -6.407411e-05, -1.117654e-05, 0, 0, 0, 0.000761393, 0.006910449, 
    0.001987529, 0.003341721, 0.002748604,
  -2.710382e-05, -1.193523e-05, -4.646286e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007683344, 0.0006897768,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007302415, -0.0001392451, 
    -3.871563e-05, 6.456384e-05, -4.910383e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01210244, 0.01102981, 0.007069195, 0.001675786, -2.014871e-07, 
    -3.539316e-07, 0.005042214, 0.001020172, -0.0001552666, -1.07015e-12, 0, 
    -8.905467e-06, 0.002738291, 0.009313652, 0.01476789, 0.01781639, 
    0.02003431, 0.01073941, 0.01133157, 0.00647369, 0.004887525, 
    -1.638708e-10, 0, 0, 0, -5.023886e-06, 0.00024749, 0.004413195, 
    0.005326705,
  0.01641976, 0.02779694, 0.02276953, 0.005418681, 0.01071628, 0.02501645, 
    0.04446141, 0.06412858, 0.05805043, 0.03385475, 0.01068252, 0.002433592, 
    0.01428798, 0.03119918, 0.07239348, 0.07464819, 0.07204019, 0.04011942, 
    0.04291866, 0.02781289, 0.01962162, 0.0184565, 0.01576619, 0.03307177, 
    0.03965972, 0.04057226, 0.03632551, 0.02859424, 0.02786299,
  0.1055011, 0.08715148, 0.07688738, 0.1133807, 0.1558496, 0.1491517, 
    0.1004844, 0.09169494, 0.1058227, 0.07448889, 0.05828517, 0.05470954, 
    0.08967637, 0.2048917, 0.1635021, 0.1128292, 0.09618071, 0.1267569, 
    0.1162552, 0.1037068, 0.1281653, 0.1360012, 0.1438559, 0.07014941, 
    0.07056904, 0.1021488, 0.102314, 0.1018842, 0.1167966,
  0.0371541, 0.03873677, 0.03219718, 0.08537544, 0.09032533, 0.1154754, 
    0.07923624, 0.06334455, 0.06485707, 0.05370761, 0.07609765, 0.12519, 
    0.1349739, 0.135432, 0.07208859, 0.0496829, 0.1124526, 0.09494826, 
    0.1692342, 0.1655996, 0.09162057, 0.08914136, 0.06443742, 0.01810444, 
    0.08168344, 0.150532, 0.1429265, 0.1482863, 0.07139573,
  0.004848952, 0.001406082, 0.1059092, 0.06684043, 0.1023767, 0.1411658, 
    0.1069524, 0.03538136, 0.01688582, 0.04671003, 0.07457799, 0.04616086, 
    0.101126, 0.1070632, 0.05904081, 0.06272937, 0.1185611, 0.1622202, 
    0.2166754, 0.1214115, 0.04481447, 0.01450379, 2.913485e-06, 0.01501743, 
    0.07927923, 0.1616339, 0.1996939, 0.03566743, 0.007279592,
  0.002717518, 0.06980328, 0.136991, 0.09279628, 0.09101917, 0.1067312, 
    0.1057035, 0.004584638, 0.0001820227, 0.04467771, 0.1246727, 0.1580346, 
    0.1721175, 0.1104581, 0.04865745, 0.146127, 0.1678278, 0.1378607, 
    0.1105763, 0.0233052, 0.0277063, 0.0001114835, 0.0007048876, 0.08641426, 
    0.2187815, 0.1698626, 0.05222715, 0.02940149, 0.00411705,
  7.491359e-05, 0.02919666, 0.3226813, 0.1310119, 0.1470707, 0.1027609, 
    0.1015159, 0.0495524, 0.03922381, 0.1051731, 0.05647274, 0.06494076, 
    0.06513344, 0.07443771, 0.1161099, 0.08909079, 0.08626609, 0.01597014, 
    0.006722552, 0.00434737, -2.50413e-07, 9.732411e-07, 0.004386619, 
    0.392905, 0.3417191, 0.2416702, 0.08354063, 0.01193937, 0.00167918,
  0.0009154282, 0.002410824, 0.002850605, 0.01186861, 0.03614991, 0.07242931, 
    0.2201117, 0.0873002, 0.1061947, 0.2486227, 0.07820483, 0.09853759, 
    0.1152578, 0.1113519, 0.09785004, 0.02889829, 0.000364713, 0.0001776593, 
    0.007944246, 6.344516e-05, 0.00888002, 0.0003276507, 0.006872943, 
    0.1412688, 0.1860245, 0.1790531, 0.04507266, 0.03529733, 0.006347786,
  0.004768163, 4.80661e-06, 4.499195e-06, 5.385364e-05, 0.0006047416, 
    0.0100111, 0.005148359, 0.0423268, 0.002154404, 0.05597988, 0.06799027, 
    0.06697385, 0.09063066, 0.02451118, 0.001920485, 0.007755122, 0.04087553, 
    0.04100891, 0.02262826, 0.06047327, 0.09043197, 0.01521338, 0.0003111918, 
    0.005824578, 0.0008160661, 0.00204642, 0.01015858, 0.05961733, 0.1195118,
  0.1802443, 0.003993591, 0.004067689, 1.424977e-06, 2.629797e-07, 
    8.821006e-07, 0.003745466, 0.009015123, 0.01804259, 0.003933232, 
    0.004609079, 0.009171305, 0.01761756, 1.536196e-05, -4.421859e-06, 
    0.002463285, 0.04038173, 0.07953256, 0.04777493, 0.1266752, 0.1404451, 
    0.05657061, 0.006387809, 0.009339051, 0.01814788, 0.02601727, 0.03298822, 
    0.03199157, 0.1246598,
  0.03519456, 0.06215919, 0.01864969, 0.03361183, 0.01118042, 0.01662905, 
    0.04059708, -0.0001586574, 6.897452e-06, 0.02249849, 0.01483753, 
    0.02585174, 0.07930601, 0.04069863, 0.05872811, 0.06345117, 0.08724695, 
    0.1962848, 0.1722981, 0.09544933, 0.06448013, 0.08615416, 0.06335944, 
    0.05633992, 0.1084089, 0.1472002, 0.1530309, 0.04039278, 0.03695005,
  0.03187227, 0.01977035, 0.0101906, 0.01486784, 0.005125335, 0.002213672, 
    0.00076301, 0, 0, 0, -1.150365e-05, 0.003217372, 0.01554911, 0.03230888, 
    0.05402622, 0.06469237, 0.1315964, 0.1291832, 0.1030182, 0.04871257, 
    0.007591841, 0.02562481, 0.07098976, 0.08129483, 0.09585931, 0.1565004, 
    0.1845618, 0.161079, 0.05322814,
  0.04548373, 0.006359924, 0.008144526, 0.0003556274, 0.0006415281, 0, 0, 0, 
    0, 0, 0, 0, -1.762624e-05, 0.009992684, 0.004779255, 0.008247282, 
    0.04486174, 0.06247768, 0.04873509, 0.003851262, 0.002105089, 
    -9.322084e-05, 0.0003489812, 0.004082576, 0.02321654, 0.04204534, 
    0.06027322, 0.07431919, 0.07480966,
  0.009076861, 0.005681868, 0.00163847, 7.114282e-05, 0.0008775722, 
    -5.59943e-06, 0, 0, 0, 0, 0, 0, 0, 0, 5.029995e-06, 0.001441732, 
    0.00391219, 0.01304878, 0.002659386, 0.003135137, 0.001467956, 0, 0, 0, 
    0.001930071, 0.01648489, 0.01542037, 0.007078445, 0.01065162,
  0.0006585651, 0.001009616, 0.0009194739, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00025871, -2.565893e-05, 0, 0.0003806091, -9.718388e-06, 0, 0, 0, 0, 0, 
    2.204132e-05, 8.989769e-05, -1.055725e-06, 0.009857247, 0.001395676,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.339966e-08, 0.009476444, 
    -0.0004266347, 0.00223779, 0.003953456, 0.00323166, 0.0002058153, 0, 0, 
    0, 0, 0, -1.526223e-07, -5.8479e-05, -6.641745e-06, 0, 0,
  0.03391937, 0.02578122, 0.006595714, 0.00868353, -8.032991e-05, 
    -0.001296165, 0.01976256, 0.003960165, 0.0004768381, -0.0002461578, 
    -8.35e-09, -0.000154918, 0.007722995, 0.06273349, 0.05326939, 0.03803363, 
    0.03256843, 0.03483567, 0.01684935, 0.01528448, 0.02374914, 0.01137584, 
    0.002607635, 0.01029055, 0.007702705, -6.146754e-05, 0.005454029, 
    0.01595251, 0.036985,
  0.0571454, 0.06916954, 0.04079404, 0.02405743, 0.02092793, 0.04728875, 
    0.08997573, 0.09392685, 0.08651549, 0.08146639, 0.05409858, 0.02558156, 
    0.08158546, 0.07451468, 0.08924088, 0.1401332, 0.1161207, 0.09980224, 
    0.08947186, 0.08366585, 0.06913009, 0.07622281, 0.07570295, 0.09316428, 
    0.08837714, 0.1261206, 0.08848663, 0.0816313, 0.08187343,
  0.1401763, 0.1180214, 0.1394193, 0.161173, 0.1797485, 0.1699685, 0.1273983, 
    0.1374909, 0.1376651, 0.1297724, 0.1326807, 0.1216094, 0.1290265, 
    0.2341242, 0.1631581, 0.1041784, 0.09975767, 0.1405538, 0.1293778, 
    0.1251142, 0.1391627, 0.1745971, 0.20382, 0.1254397, 0.123004, 0.1295084, 
    0.1212555, 0.118877, 0.1547095,
  0.03268552, 0.03323144, 0.02985225, 0.08065248, 0.07689923, 0.1052109, 
    0.06964412, 0.05883809, 0.05716425, 0.04490199, 0.07718654, 0.1157395, 
    0.1126951, 0.1097497, 0.06667256, 0.0321838, 0.09506726, 0.08641197, 
    0.1542929, 0.167981, 0.08663659, 0.07315166, 0.06149062, 0.02231574, 
    0.08145075, 0.1248258, 0.1253848, 0.1283524, 0.06242368,
  0.00127014, 0.0006968852, 0.09333569, 0.05291674, 0.101752, 0.1213335, 
    0.09500112, 0.03163104, 0.012594, 0.05209241, 0.075518, 0.04413555, 
    0.09583861, 0.09384936, 0.04326653, 0.05173423, 0.1124386, 0.1361328, 
    0.201677, 0.1261401, 0.03800497, 0.01148623, 2.4572e-07, 0.007773572, 
    0.06840585, 0.1473029, 0.1724792, 0.02919268, 0.0005261892,
  0.0009152408, 0.05449783, 0.1129049, 0.07415606, 0.08254775, 0.08922901, 
    0.1010129, 0.003707962, 0.0001567489, 0.03804513, 0.1128801, 0.1364886, 
    0.1633814, 0.09102964, 0.04314911, 0.1382036, 0.1481741, 0.1362386, 
    0.09630743, 0.01515057, 0.01359044, 6.742945e-06, 0.008011782, 
    0.07230067, 0.1701493, 0.1753094, 0.04350217, 0.01236781, 7.999398e-05,
  1.14932e-05, 0.02828655, 0.2612796, 0.09976513, 0.1115816, 0.07719497, 
    0.08786444, 0.04219232, 0.03148766, 0.09095211, 0.05361809, 0.0561465, 
    0.05129031, 0.05957611, 0.1048936, 0.07646192, 0.07297708, 0.01704918, 
    0.005722786, 0.002070971, 5.825997e-08, 4.740867e-07, 0.001418513, 
    0.3303706, 0.3088515, 0.2077199, 0.05401104, 0.007903195, 2.520068e-05,
  0.0006966391, 0.004566985, 0.002392567, 0.002698981, 0.03348133, 
    0.05848889, 0.216341, 0.07145882, 0.08833034, 0.2130718, 0.06769564, 
    0.08051064, 0.1039161, 0.1055171, 0.08890976, 0.02765266, 0.0002881758, 
    -7.850739e-05, 0.00397982, -1.312256e-05, 0.01181524, -1.730211e-05, 
    0.006009474, 0.1034249, 0.1445759, 0.2136554, 0.04267434, 0.02933664, 
    0.0009444364,
  0.0001103636, 3.873207e-06, 2.905955e-06, 2.225065e-05, 0.0007486361, 
    0.00491492, 0.001607173, 0.04244878, 0.003341973, 0.04827549, 0.06540106, 
    0.06531437, 0.08138251, 0.02306418, 0.006709585, 0.01375585, 0.03592012, 
    0.03917544, 0.0332738, 0.05574866, 0.07737613, 0.01591966, 0.0003955991, 
    0.002347659, 0.001406001, 0.004807701, 0.01339348, 0.04817309, 0.09657235,
  0.09964331, 0.001413695, 0.000418489, -1.986283e-06, 2.330096e-07, 
    4.618016e-07, 0.009250535, 0.01015398, 0.02977581, 0.004258407, 
    0.01823374, 0.01417949, 0.02281297, 0.001225822, -5.474318e-06, 
    0.003305975, 0.03585302, 0.06155044, 0.02804821, 0.1097107, 0.1128571, 
    0.03694059, 0.00563485, 0.009132432, 0.01173141, 0.02610422, 0.01587958, 
    0.0582198, 0.106135,
  0.05646566, 0.05994414, 0.01684699, 0.02121979, 0.01921411, 0.01499586, 
    0.03352826, -0.000102586, 0.0005913083, 0.03663099, 0.02488227, 
    0.04743914, 0.09754923, 0.08091551, 0.08808801, 0.08077005, 0.09391905, 
    0.2000675, 0.1473048, 0.06385581, 0.07260114, 0.07732216, 0.04601723, 
    0.04384077, 0.1095854, 0.1302719, 0.1227741, 0.03846958, 0.07772347,
  0.09778674, 0.05962093, 0.05373621, 0.03997516, 0.02011886, 0.02492016, 
    0.001225529, 0.0002342987, 2.055747e-05, -1.740234e-07, 0.0001600392, 
    0.008703765, 0.02897599, 0.06448943, 0.08808328, 0.1094689, 0.1965524, 
    0.1901967, 0.1555247, 0.1109696, 0.01622951, 0.05648596, 0.1197122, 
    0.1547044, 0.1494597, 0.2226247, 0.2122438, 0.1924213, 0.1389564,
  0.1365693, 0.05366202, 0.02295073, 0.008012237, 0.006249289, 0.003800593, 
    -2.419228e-06, 0, 0, 0, 0, -5.41477e-06, 0.002919856, 0.02455393, 
    0.01780185, 0.04752412, 0.1150622, 0.1065868, 0.07440929, 0.01877881, 
    0.009409403, 0.01822649, 0.01176511, 0.01846993, 0.0539794, 0.08414248, 
    0.1329809, 0.1605235, 0.1878903,
  0.05697247, 0.01290955, 0.01005218, 0.006082614, 0.00601061, -4.923086e-05, 
    0.0001022875, 0.001505641, 0, 0, 0, 0, 0, 0.0003541916, 0.008493127, 
    0.01569765, 0.03587536, 0.06674715, 0.01563885, 0.01215561, 0.0100827, 
    0.003442388, 0.0001191111, 0.0002674123, 0.004373953, 0.02466985, 
    0.04915818, 0.04737322, 0.0477676,
  0.008661246, 0.007586571, 0.00572291, 0.002989822, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.280022e-06, 0.005889037, -0.0001190856, 0.00125189, 0.0090012, 
    0.01302157, 0.001361107, -1.030558e-05, -5.340244e-06, -5.135567e-08, 0, 
    0.001652655, 0.002196139, -3.790145e-06, 0.01273673, 0.004741399,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.237105e-06, 
    1.091237e-06, -5.256646e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001356449, 0.01483385, 0.006528482, 
    0.007417846, 0.009875877, 0.006107758, 0.001673685, -2.292589e-06, 
    -8.675137e-08, -1.292121e-10, 0.001800745, 0.02124237, 0.004983074, 
    -0.001008619, -0.0003840189, -5.138222e-05, 0,
  0.04071791, 0.02568392, 0.01429065, 0.009039256, -0.0003181102, 
    0.007811655, 0.06406096, 0.009796592, 0.00534498, -0.0003394354, 
    2.836342e-05, 0.003258782, 0.0164318, 0.1673915, 0.1450562, 0.09408784, 
    0.09176858, 0.07662718, 0.04184649, 0.07474127, 0.09713255, 0.07700734, 
    0.07548621, 0.05090914, 0.07608992, 0.08205096, 0.03700156, 0.03694197, 
    0.07580681,
  0.1099695, 0.1137586, 0.1027714, 0.1062083, 0.08749799, 0.112273, 
    0.1314838, 0.1354902, 0.1139627, 0.1390562, 0.1199222, 0.1079192, 
    0.1597758, 0.1592761, 0.1430389, 0.2016003, 0.1461594, 0.1194721, 
    0.1295957, 0.1175096, 0.1157301, 0.1183939, 0.1632787, 0.2067649, 
    0.2012368, 0.2174352, 0.1735341, 0.1460438, 0.153484,
  0.1589193, 0.1421752, 0.1514478, 0.1740122, 0.1833404, 0.1748794, 
    0.1289503, 0.1435884, 0.1523823, 0.1296543, 0.1370308, 0.1207252, 
    0.1105085, 0.232262, 0.1660775, 0.1154413, 0.09971376, 0.1344554, 
    0.122434, 0.1179817, 0.1408421, 0.1836657, 0.213172, 0.1521617, 
    0.1389283, 0.139494, 0.1387706, 0.1077935, 0.1712599,
  0.03109584, 0.02998301, 0.02643983, 0.08086912, 0.07341564, 0.09656431, 
    0.05378812, 0.05034916, 0.04049363, 0.03601513, 0.06353433, 0.09730828, 
    0.09993635, 0.09417439, 0.05691599, 0.02565478, 0.08479369, 0.08143534, 
    0.1344735, 0.164822, 0.07340842, 0.05223972, 0.04689229, 0.01919475, 
    0.07996958, 0.1032711, 0.1222837, 0.1210773, 0.05937009,
  0.000333039, 0.0006704705, 0.08104366, 0.04486322, 0.09497955, 0.0916681, 
    0.06303729, 0.02810615, 0.007129756, 0.05438686, 0.07037576, 0.04346097, 
    0.08683744, 0.07781885, 0.03145386, 0.04698084, 0.110308, 0.1227868, 
    0.2039345, 0.1293249, 0.03711498, 0.002857072, -6.713236e-08, 
    0.0007786201, 0.05575351, 0.1306246, 0.1544074, 0.02402188, 2.19888e-05,
  0.0001812925, 0.04429841, 0.1009765, 0.06681966, 0.07343176, 0.06358334, 
    0.09267835, 0.005896181, 9.577328e-05, 0.0329947, 0.09638464, 0.1175653, 
    0.1485289, 0.07200491, 0.03836727, 0.1329051, 0.139453, 0.1334362, 
    0.07705828, 0.008891291, 0.001720768, 8.466375e-07, 0.008546325, 
    0.05694606, 0.1333296, 0.1600112, 0.0277159, 0.002248096, 2.366155e-05,
  3.491449e-06, 0.02669042, 0.1997748, 0.07374336, 0.07663058, 0.05193407, 
    0.07765615, 0.03555708, 0.02619291, 0.07421851, 0.04828261, 0.04213045, 
    0.03586205, 0.04707881, 0.09593156, 0.06923379, 0.06113534, 0.01775247, 
    0.005186849, 9.911244e-05, 6.950962e-09, 3.552694e-07, 0.000983505, 
    0.2368432, 0.2887168, 0.1688053, 0.03942152, 0.002558781, 2.598437e-06,
  0.0004073725, 0.006586117, 0.002421076, 0.001247419, 0.02555895, 0.0550908, 
    0.1878269, 0.05556151, 0.07587273, 0.187332, 0.05481724, 0.0550281, 
    0.09573036, 0.09966503, 0.07390934, 0.03499316, 0.0001723147, 
    0.0004572364, 0.0002588134, -4.742462e-05, 0.008321183, 0.0004771035, 
    0.006529015, 0.07798263, 0.115198, 0.2429133, 0.03515928, 0.01823544, 
    0.0004546912,
  1.652174e-05, 2.811521e-06, 4.297922e-06, 8.796198e-06, 0.001036034, 
    0.004313455, 0.003350592, 0.04367312, 0.00450646, 0.03861669, 0.06238203, 
    0.0687746, 0.07904886, 0.0209557, 0.005277392, 0.01521301, 0.03961055, 
    0.03317478, 0.04419657, 0.0551276, 0.06590718, 0.01723714, 0.0003781613, 
    0.001201065, 0.001733889, 0.01313714, 0.0233017, 0.02196757, 0.07299699,
  0.05711968, 0.0001388971, 3.011384e-05, -3.052976e-06, 8.186895e-08, 
    5.07772e-07, 0.01166254, 0.01024416, 0.03526634, 0.0053066, 0.03770934, 
    0.01491376, 0.02292731, 0.008481303, 0.0001251699, 0.00235438, 
    0.03351295, 0.03419396, 0.02612764, 0.1046134, 0.09353013, 0.02767578, 
    0.004334752, 0.007629421, 0.00618647, 0.02829121, 0.008016201, 
    0.04844109, 0.0740832,
  0.0503739, 0.04665105, 0.02368345, 0.02149005, 0.02401201, 0.005388489, 
    0.01211918, 0.003264996, 0.004973896, 0.07206935, 0.03477244, 0.06278415, 
    0.1121116, 0.1016626, 0.08425787, 0.09397162, 0.0951761, 0.1843577, 
    0.1223118, 0.03344294, 0.07663594, 0.07296097, 0.03609391, 0.03967087, 
    0.09718746, 0.09996125, 0.07463118, 0.02889877, 0.06992218,
  0.1298072, 0.09803779, 0.1072118, 0.08333418, 0.07024141, 0.09492498, 
    0.005192971, 0.03509785, 0.002965314, 8.897472e-06, 0.00765466, 
    0.02311765, 0.04743841, 0.08137028, 0.123747, 0.1330805, 0.2239077, 
    0.2140792, 0.1769546, 0.1627126, 0.05587387, 0.08828259, 0.1492807, 
    0.1516603, 0.158429, 0.23114, 0.2039448, 0.1713135, 0.1429088,
  0.193394, 0.1359804, 0.07456618, 0.07164237, 0.08461659, 0.08476782, 
    0.02885893, 0, -4.018258e-06, -3.721889e-07, 0, 0.001609142, 0.01889926, 
    0.05683011, 0.0882784, 0.09371983, 0.1487132, 0.1201956, 0.1111187, 
    0.0452195, 0.0388774, 0.05468136, 0.04513171, 0.04887889, 0.09466776, 
    0.1320107, 0.1592073, 0.2049607, 0.2456789,
  0.114792, 0.0674228, 0.04733182, 0.02895144, 0.01322735, 0.008764211, 
    0.02389365, 0.02371884, 0.001877821, 4.605616e-05, 0, -4.339521e-08, 
    -0.0004325284, 0.02992018, 0.07065265, 0.1033826, 0.1039935, 0.1362864, 
    0.05358038, 0.04272958, 0.03130323, 0.01811971, 0.011221, 0.01640233, 
    0.01805448, 0.04936458, 0.1029409, 0.1179382, 0.1111711,
  0.01762462, 0.0248345, 0.01249988, 0.005407447, 0.0002053147, 2.835807e-05, 
    0, 0, 0, 0, -2.737148e-09, 0, -1.121206e-06, 0.01332245, 0.0255898, 
    0.014896, 0.04243423, 0.03170536, 0.03789771, 0.04499033, 0.01555771, 
    0.007340341, 0.004426945, -5.014299e-05, 0.003725332, 0.003653191, 
    -1.358197e-05, 0.01728549, 0.009515721,
  -9.942556e-08, 3.594539e-05, -9.526087e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.869868e-05, 0.003432505, 0.003310885, 0.004605932, 0.007670173, 
    0.004657683, 1.485379e-05, -1.695306e-05, -1.681324e-06, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001092149, 0.002571091, 0.003235067, 
    0.01528176, 0.01965584, 0.1052285, 0.1362143, 0.08420543, 0.03600416, 
    0.009116905, -0.0003902226, -5.646205e-05, 0.01924059, 0.1025404, 
    0.05992985, 0.009396583, 0.01715384, -8.856218e-05, 0,
  0.1164333, 0.1323015, 0.08161372, 0.08032405, 7.867349e-05, 0.02528206, 
    0.1149158, 0.02270767, 0.0131669, -0.0007068003, 0.006735818, 0.00967571, 
    0.06807992, 0.2570063, 0.2046655, 0.1539282, 0.142582, 0.1324632, 
    0.1149283, 0.1762691, 0.1754342, 0.1477685, 0.2039665, 0.1319802, 
    0.1743123, 0.1644923, 0.08324458, 0.08902727, 0.1705706,
  0.1705891, 0.1752525, 0.197632, 0.1867362, 0.1437131, 0.1495005, 0.1592761, 
    0.1869779, 0.1865071, 0.1904019, 0.1711214, 0.1697507, 0.23716, 
    0.1975863, 0.1506221, 0.2023172, 0.1801054, 0.1272683, 0.151721, 
    0.1367021, 0.1435433, 0.1858211, 0.205026, 0.2250152, 0.2295346, 
    0.2363076, 0.1999077, 0.2057431, 0.2237946,
  0.1646508, 0.1548728, 0.1484845, 0.1765644, 0.1787907, 0.1850158, 
    0.1331291, 0.1411424, 0.1566415, 0.1385959, 0.1354111, 0.1096035, 
    0.1010412, 0.2161234, 0.1537986, 0.1107236, 0.1046347, 0.1302904, 
    0.1039732, 0.1152101, 0.1555282, 0.1824559, 0.223046, 0.1598182, 
    0.1334496, 0.1353801, 0.1293467, 0.102402, 0.1754757,
  0.03692352, 0.02790363, 0.02865899, 0.07813925, 0.06440504, 0.07656519, 
    0.05164436, 0.04433459, 0.02924179, 0.03177656, 0.05515036, 0.08201723, 
    0.09195286, 0.08633275, 0.05389395, 0.02257307, 0.0856267, 0.07825059, 
    0.1197548, 0.1679497, 0.08777265, 0.04338191, 0.0333422, 0.02067523, 
    0.0783067, 0.08607092, 0.1135581, 0.1283366, 0.05539791,
  0.0001602023, 0.0001005555, 0.07608193, 0.03473325, 0.0755745, 0.07683547, 
    0.03476216, 0.02379244, 0.003482181, 0.05057064, 0.05850804, 0.03899187, 
    0.07565919, 0.05321126, 0.02348206, 0.04736534, 0.1027714, 0.1071272, 
    0.1744585, 0.1093293, 0.03179545, 3.583898e-05, -4.473029e-08, 
    0.0001178855, 0.04865417, 0.1122077, 0.1339811, 0.01735262, 3.482382e-05,
  0.001819193, 0.04183813, 0.08592609, 0.05556443, 0.06677903, 0.04137725, 
    0.07891617, 0.005864725, 0.0001091545, 0.04127865, 0.08044197, 0.1080034, 
    0.1331729, 0.04887716, 0.02570841, 0.1242448, 0.131424, 0.1270186, 
    0.06037638, 0.005155939, 2.398064e-05, 1.155765e-07, 0.00766299, 
    0.04528374, 0.1161459, 0.1275105, 0.02559219, 0.0001472713, 9.852806e-05,
  3.37076e-05, 0.02322793, 0.1765873, 0.05680221, 0.06666453, 0.03851905, 
    0.06719966, 0.02915623, 0.0239642, 0.06746343, 0.04409357, 0.03306129, 
    0.02843262, 0.03863927, 0.09335235, 0.06535689, 0.04583662, 0.01908703, 
    0.005445017, 7.81939e-05, -1.544071e-09, 4.206915e-07, 0.0002670725, 
    0.1782561, 0.2661882, 0.1435368, 0.03238909, -4.930964e-05, 1.375985e-06,
  0.002736079, 0.00442377, 0.002194889, 0.002355207, 0.0243775, 0.05617867, 
    0.1753193, 0.05042118, 0.06769019, 0.1589981, 0.04856326, 0.04450482, 
    0.08053303, 0.09425093, 0.06784686, 0.02432722, 0.00102163, 0.004504053, 
    -7.479775e-05, -3.662447e-05, 0.006482331, 0.000718054, 0.01526864, 
    0.06041284, 0.1149518, 0.2549154, 0.02984004, 0.004711799, 0.000233093,
  0.0006809711, 1.727961e-06, 2.370577e-06, 3.117546e-06, 0.003353298, 
    0.006213484, 0.007406383, 0.0553269, 0.002837578, 0.03248166, 0.06460603, 
    0.07663751, 0.07658291, 0.01768898, 0.003954178, 0.01072198, 0.04058024, 
    0.03695036, 0.04439545, 0.0521425, 0.06170969, 0.01875621, 0.0005936449, 
    0.0008204496, 0.009104115, 0.02287664, 0.01583842, 0.003665187, 0.05559922,
  0.03457508, 1.282226e-05, 2.950057e-07, 6.794297e-06, 1.638325e-07, 
    1.52095e-07, 0.01563088, 0.01064904, 0.03075369, 0.01111345, 0.0447911, 
    0.02483778, 0.02552709, 0.02004419, 0.008759498, 0.0004121594, 
    0.03452931, 0.02416325, 0.008648827, 0.1127516, 0.07557117, 0.02491746, 
    0.002385593, 0.00543312, 0.005572725, 0.02169507, 0.003622902, 
    0.03136387, 0.05171259,
  0.02543184, 0.03032841, 0.03206501, 0.0200837, 0.02061748, 0.001457642, 
    0.01382727, 0.006875935, 0.01496308, 0.1057957, 0.04238322, 0.07105987, 
    0.1143192, 0.1377442, 0.1126741, 0.09956415, 0.0901577, 0.1567671, 
    0.08828615, 0.01696722, 0.07607506, 0.06576814, 0.04655974, 0.04132716, 
    0.08194036, 0.08074571, 0.07077657, 0.02524738, 0.05184246,
  0.1305736, 0.09992707, 0.1412926, 0.1522804, 0.1087186, 0.1510717, 
    0.02869786, 0.07986932, 0.02227823, 0.004101846, 0.03724263, 0.07502484, 
    0.08583416, 0.1184847, 0.1606838, 0.1594049, 0.2288518, 0.2283597, 
    0.1704255, 0.1652975, 0.1059102, 0.08977796, 0.1662348, 0.1473568, 
    0.1682139, 0.2271889, 0.1955184, 0.1457013, 0.1388153,
  0.2206719, 0.16528, 0.1245449, 0.1449107, 0.2104963, 0.2255909, 0.09792799, 
    -0.000150418, 0.0003169173, 8.447102e-05, 0.004812092, 0.006433393, 
    0.04963037, 0.1074857, 0.1499666, 0.1204275, 0.1575872, 0.1344617, 
    0.1305828, 0.09599577, 0.06309909, 0.1070187, 0.1076279, 0.0942369, 
    0.1319421, 0.1462146, 0.1732202, 0.2199074, 0.2444583,
  0.1671859, 0.1088641, 0.1000916, 0.09097508, 0.06782184, 0.1089146, 
    0.1771638, 0.1240307, 0.04952312, 0.01339451, 1.372273e-06, 
    -3.414581e-05, 0.007720843, 0.07443008, 0.1456903, 0.1687292, 0.1492938, 
    0.1909888, 0.1218389, 0.07659651, 0.06152767, 0.06064125, 0.05045931, 
    0.02528751, 0.04672783, 0.1250877, 0.1793196, 0.1975788, 0.1665486,
  0.03970169, 0.06401198, 0.04115869, 0.03952894, 0.01751278, 0.005738832, 
    0.004565778, 0.00923615, 0.004961052, 0.003229019, 0.0001577548, 
    -6.230768e-05, 0.02191746, 0.0301514, 0.05760315, 0.06640224, 0.1005247, 
    0.06658333, 0.07202747, 0.0974711, 0.06983371, 0.02035653, 0.01932197, 
    0.004232321, 0.01189642, 0.005498549, -0.0001596249, 0.02633236, 
    0.02306549,
  5.815824e-05, 0.002735541, 5.998997e-07, -7.060493e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, -5.729517e-05, 0.00645761, 0.01279786, 0.01437603, 0.01703925, 
    0.01538816, 0.01224822, 0.004825721, 0.0001813544, -6.642781e-06, 0, 0, 
    0, 0, -1.850079e-08, -1.799705e-05, -0.0001119163,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -9.515882e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004416703, 0.005397001, 
    0.00708212, 0.04661752, 0.0806194, 0.1671988, 0.204235, 0.1753612, 
    0.1160651, 0.03459512, 0.03463272, 0.007796701, 0.08174478, 0.1242073, 
    0.0869575, 0.03999884, 0.06026884, 0.01665705, 0.0006821856,
  0.1637407, 0.2264057, 0.1545059, 0.1577782, 0.003300602, 0.05699975, 
    0.173909, 0.0473959, 0.05281723, 0.01662293, 0.01378085, 0.007306824, 
    0.1449629, 0.2798861, 0.2514321, 0.1680856, 0.1408881, 0.1451926, 
    0.1282195, 0.2234322, 0.2380581, 0.1953436, 0.2442411, 0.1977189, 
    0.2222244, 0.1921363, 0.113027, 0.101221, 0.2752422,
  0.1904526, 0.2048401, 0.2553531, 0.2319942, 0.1756005, 0.1745372, 0.176657, 
    0.1949581, 0.2194892, 0.2109407, 0.1955556, 0.1854759, 0.2403627, 
    0.2144108, 0.1643266, 0.1999521, 0.1829264, 0.1445781, 0.1617301, 
    0.1499799, 0.18133, 0.2139341, 0.2347927, 0.2174256, 0.235556, 0.2368338, 
    0.2024359, 0.2226587, 0.26141,
  0.1635633, 0.1675295, 0.1486142, 0.1748101, 0.1683056, 0.1884481, 
    0.1334834, 0.1347276, 0.1600837, 0.1375075, 0.1479282, 0.1009548, 
    0.1099081, 0.2027832, 0.1527819, 0.1011861, 0.1211524, 0.1124205, 
    0.09675834, 0.1194226, 0.150934, 0.175977, 0.202617, 0.1631372, 
    0.1257544, 0.1304791, 0.1246857, 0.1004806, 0.1747846,
  0.03942686, 0.02715279, 0.02037622, 0.08028446, 0.05541811, 0.0615348, 
    0.04833419, 0.04071613, 0.0345061, 0.01925852, 0.05102208, 0.07196429, 
    0.08879232, 0.06856026, 0.04927473, 0.01927779, 0.08722511, 0.07794912, 
    0.1267077, 0.154588, 0.05989932, 0.0377719, 0.03534797, 0.02039998, 
    0.08249471, 0.07526474, 0.101538, 0.1100798, 0.06247713,
  0.0001230013, -9.065703e-06, 0.07639269, 0.03391622, 0.06222428, 
    0.08270165, 0.03139959, 0.02023801, 0.002183445, 0.05039288, 0.05087281, 
    0.03662086, 0.0690148, 0.03988617, 0.02239187, 0.03845191, 0.07992038, 
    0.1061114, 0.162857, 0.08863588, 0.02308934, -9.452208e-05, 
    -2.644029e-07, 0.0001012467, 0.04330552, 0.09180626, 0.1119836, 
    0.008499081, 2.884109e-05,
  0.002280142, 0.041169, 0.06307177, 0.05427063, 0.06258087, 0.02849872, 
    0.06364989, 0.002768584, 9.901477e-05, 0.05383892, 0.06740586, 0.1001443, 
    0.1338137, 0.04823314, 0.02488615, 0.1193735, 0.1285834, 0.1152396, 
    0.04950025, 0.004480481, 8.902358e-06, 4.067274e-08, 0.0002749379, 
    0.03023422, 0.1062459, 0.1030929, 0.01907604, 7.918859e-06, 0.008350223,
  0.001765307, 0.02756152, 0.1703627, 0.05114689, 0.05953556, 0.03077244, 
    0.05400303, 0.02433259, 0.01890508, 0.06537288, 0.04144496, 0.02889441, 
    0.0234687, 0.03504722, 0.09131052, 0.05807832, 0.04050814, 0.02393711, 
    0.007240724, 4.559804e-05, 1.010733e-08, 1.251738e-06, 7.285306e-05, 
    0.1302306, 0.2548709, 0.1278784, 0.02163666, -3.776844e-06, 1.310255e-06,
  0.01274815, 0.003808105, 0.00289868, 0.006526635, 0.03128658, 0.05686649, 
    0.1521813, 0.04459415, 0.06339224, 0.1528975, 0.04657029, 0.03775543, 
    0.07147339, 0.08755207, 0.06959993, 0.01138619, 0.003032405, 0.003035994, 
    -1.765194e-05, -2.193732e-05, 0.005991628, 0.00113886, 0.02781751, 
    0.04863953, 0.1433658, 0.2410628, 0.0270494, 0.002727408, 0.0008587879,
  0.003963564, 3.805719e-06, 1.066643e-06, 2.201191e-06, 0.007681534, 
    0.01076019, 0.01926177, 0.06242342, 0.002502162, 0.04493767, 0.08027359, 
    0.08304667, 0.07611387, 0.02108107, 0.007422911, 0.01068859, 0.0404649, 
    0.03170192, 0.05026288, 0.0591977, 0.062016, 0.01865672, 0.0005690003, 
    0.0006716307, 0.002489264, 0.01336771, 0.01875018, 0.003451956, 0.04704918,
  0.03319424, 3.947773e-06, 3.386701e-07, 1.760617e-06, 2.731306e-07, 
    5.044347e-06, 0.01556064, 0.01114603, 0.02416582, 0.01788077, 0.05708906, 
    0.03937384, 0.03130078, 0.006656667, 0.001577795, 0.002336295, 
    0.03741403, 0.02340766, 0.002196495, 0.09736498, 0.05544107, 0.0221555, 
    0.001520771, 0.004253353, 0.00459567, 0.02387855, 0.004590518, 
    0.02978177, 0.04375526,
  0.009508858, 0.01521319, 0.024498, 0.02435048, 0.0189517, 0.004362902, 
    0.0183983, 0.01783628, 0.02072073, 0.1314679, 0.05332262, 0.08569756, 
    0.09357196, 0.1317101, 0.1291667, 0.09775261, 0.09171457, 0.1386469, 
    0.06997135, 0.009081411, 0.06887513, 0.05717955, 0.05110952, 0.0510924, 
    0.06782026, 0.08146673, 0.05697151, 0.02436741, 0.03805472,
  0.1240242, 0.08825863, 0.1449164, 0.211439, 0.1261478, 0.1447783, 
    0.06903769, 0.1213342, 0.06418024, 0.03350127, 0.05454176, 0.09069199, 
    0.1087777, 0.1309889, 0.1607145, 0.1919626, 0.2353157, 0.2257908, 
    0.165322, 0.1661404, 0.1198566, 0.1008768, 0.1651042, 0.1440509, 
    0.1795176, 0.2229066, 0.1845451, 0.1235454, 0.1309226,
  0.2268765, 0.2011883, 0.1491518, 0.1759845, 0.2254723, 0.2554072, 
    0.1544763, 0.008743894, 0.003582697, 0.02276252, 0.03906991, 0.04872796, 
    0.09695721, 0.1951355, 0.2016912, 0.1728189, 0.1754588, 0.1629564, 
    0.1473813, 0.117066, 0.07739353, 0.161024, 0.1804565, 0.1719558, 
    0.189629, 0.1577072, 0.18078, 0.2066377, 0.230406,
  0.2175279, 0.1498133, 0.1532273, 0.1536792, 0.1198294, 0.2209348, 
    0.2996392, 0.2552538, 0.1880849, 0.1024955, 0.003887673, 0.004328888, 
    0.03272676, 0.1328014, 0.176465, 0.1909358, 0.1947952, 0.2513766, 
    0.1604377, 0.1028481, 0.1098247, 0.109236, 0.06389021, 0.04568246, 
    0.123666, 0.2028472, 0.2251594, 0.2283391, 0.1734898,
  0.09173161, 0.1241139, 0.07777748, 0.08479142, 0.08704541, 0.05812575, 
    0.06102053, 0.0601664, 0.02944147, 0.03160327, 0.01244431, 0.01880939, 
    0.06071182, 0.06422555, 0.09279874, 0.08459098, 0.139612, 0.1704213, 
    0.1533058, 0.1617891, 0.09918839, 0.04879627, 0.02771446, 0.01772249, 
    0.04989266, 0.007713088, -0.0002474309, 0.06628651, 0.06983026,
  0.03860375, 0.04038617, 0.03810197, 0.03341144, 0.01634354, 0.003278785, 
    0.002380151, 0.003547242, 0.000262516, 5.918501e-06, 0, -7.92063e-05, 
    0.004407182, 0.01151132, 0.01736182, 0.01857797, 0.01949095, 0.01894901, 
    0.01849254, 0.009100329, 0.005287327, 0.0002319641, -1.51862e-05, 
    -1.080281e-06, -1.986762e-08, 0, -6.688255e-06, -0.00429738, 0.03356687,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -0.0001626298, -0.0001626298, -0.0001626298, -0.0001626298, 
    -0.0001626298, -0.0001626298, -0.0001626298, 0,
  0.006054895, 0.004080682, 0.002378028, -4.988973e-05, 0, -8.809185e-05, 0, 
    0, 0, 0.003345293, 0.006581978, 0.008572697, 0.004738943, 0.1202681, 
    0.1283388, 0.223663, 0.2681596, 0.2410845, 0.1845541, 0.1226661, 
    0.1057127, 0.06333551, 0.1300344, 0.1064728, 0.07497638, 0.03697752, 
    0.07876252, 0.08866321, 0.01704648,
  0.1592276, 0.2274643, 0.1314783, 0.1555283, 0.05123201, 0.1260861, 
    0.1962646, 0.09138012, 0.07994172, 0.06443116, 0.04111223, 0.0646036, 
    0.1718922, 0.2713533, 0.2464075, 0.1801131, 0.1487224, 0.1678731, 
    0.1512346, 0.2276252, 0.2541997, 0.177634, 0.2692459, 0.2105979, 
    0.2302456, 0.1898937, 0.1272973, 0.118017, 0.270564,
  0.2039716, 0.1954809, 0.2659625, 0.2361045, 0.1779782, 0.1973025, 
    0.1817327, 0.2023585, 0.2215202, 0.2259193, 0.2199287, 0.1953062, 
    0.2290474, 0.237596, 0.1710301, 0.2107264, 0.1875185, 0.1486498, 
    0.1687516, 0.1773282, 0.1985682, 0.243374, 0.248875, 0.2211187, 
    0.2391398, 0.2349634, 0.217909, 0.2331747, 0.2693264,
  0.1594032, 0.1673146, 0.1535313, 0.171405, 0.1731372, 0.1883138, 0.1453606, 
    0.1343565, 0.1392291, 0.1393797, 0.1399257, 0.1044329, 0.1105219, 
    0.2014373, 0.1557559, 0.1003518, 0.1197628, 0.1049989, 0.09724526, 
    0.1273654, 0.1459428, 0.1927305, 0.2098429, 0.155062, 0.1104358, 
    0.1227745, 0.1139752, 0.09613346, 0.1648879,
  0.03807758, 0.02988921, 0.01541355, 0.07785714, 0.05293126, 0.0509412, 
    0.0498589, 0.039038, 0.02701904, 0.009422378, 0.04716073, 0.06999855, 
    0.08462422, 0.06230145, 0.04034558, 0.01588665, 0.06775498, 0.07394287, 
    0.1199594, 0.1478624, 0.06086844, 0.03770068, 0.03426245, 0.01556952, 
    0.08109007, 0.07056779, 0.0885096, 0.09889729, 0.05706599,
  0.0001495244, 4.822325e-05, 0.08431502, 0.0298935, 0.04593531, 0.07863738, 
    0.02387095, 0.01869427, 0.001208401, 0.05141419, 0.04546667, 0.03266614, 
    0.06293686, 0.02304809, 0.02835762, 0.03974142, 0.05779071, 0.0968163, 
    0.1362888, 0.09091422, 0.01582551, -0.0001106901, -7.597015e-07, 
    2.283424e-05, 0.03748569, 0.06946959, 0.1051072, 0.004126173, 0.000145671,
  0.005062426, 0.03470675, 0.05540974, 0.05632628, 0.06268305, 0.02688483, 
    0.05662895, 0.001846413, 6.820987e-05, 0.05182242, 0.0542913, 0.08873588, 
    0.1248346, 0.03615544, 0.02450898, 0.1133915, 0.1325528, 0.1078411, 
    0.04256136, 0.00479305, 2.719775e-07, -7.801316e-09, -1.313358e-05, 
    0.01745993, 0.1089674, 0.09901981, 0.01715614, 0.0005748567, 0.00199266,
  0.0005239808, 0.051971, 0.1871391, 0.05512647, 0.05591292, 0.03072694, 
    0.04397716, 0.02245548, 0.01357912, 0.06347829, 0.0449397, 0.03017701, 
    0.02749122, 0.03326787, 0.08709989, 0.05936011, 0.0354557, 0.02658092, 
    0.003130404, 0.0001074346, 4.104486e-08, 1.592604e-06, 7.157559e-05, 
    0.09585185, 0.2527806, 0.1217269, 0.01750445, 0.0001003778, 3.806136e-07,
  0.04271316, 0.02840097, 0.008673371, 0.01322686, 0.02828922, 0.0598818, 
    0.1411563, 0.03591494, 0.0593279, 0.1537452, 0.04267043, 0.03544866, 
    0.06704596, 0.08388676, 0.06356522, 0.009752127, 0.007947008, 
    0.005177933, 3.435655e-06, -2.297073e-05, 0.005449622, 0.01256252, 
    0.04203064, 0.04618413, 0.1397294, 0.2181104, 0.02611568, 0.003684824, 
    0.004833675,
  0.002170583, 4.321656e-06, 8.022864e-07, 1.583264e-06, 0.01067407, 
    0.01898391, 0.01961705, 0.06049424, 0.002270621, 0.04383427, 0.07906522, 
    0.08350505, 0.073917, 0.02309025, 0.008275812, 0.009026967, 0.0419221, 
    0.0291306, 0.04615412, 0.0528935, 0.06380916, 0.0210446, 0.001076637, 
    0.001077844, 0.006010851, 0.009609523, 0.01562604, 0.001169989, 0.03562053,
  0.03729611, 6.652835e-06, 1.221409e-06, 4.571343e-07, 1.140067e-06, 
    0.0002267358, 0.0135038, 0.01162337, 0.01954467, 0.01691877, 0.05841079, 
    0.05713929, 0.02720098, 0.009995883, 1.70165e-05, 0.0003847809, 
    0.03618603, 0.01906012, 0.001145049, 0.07297841, 0.0380478, 0.01797507, 
    0.003706055, 0.0009314318, 0.004743197, 0.02520013, 0.004127378, 
    0.0211461, 0.02721719,
  0.002560629, 0.007570184, 0.01628507, 0.02246426, 0.02203322, 0.003362164, 
    0.0204952, 0.0213125, 0.02733981, 0.1432775, 0.05798732, 0.08304884, 
    0.06805512, 0.1183224, 0.1330825, 0.09143858, 0.1035685, 0.1369549, 
    0.05294186, 0.008881366, 0.06546661, 0.0540209, 0.06131615, 0.05590011, 
    0.06014699, 0.07569005, 0.04946465, 0.02548748, 0.02592797,
  0.1083908, 0.07020488, 0.1591872, 0.2636234, 0.1108654, 0.1370998, 
    0.1503965, 0.1176089, 0.08381005, 0.06423532, 0.05548432, 0.112363, 
    0.1206979, 0.1368981, 0.1690735, 0.204269, 0.2327793, 0.2225484, 
    0.1377129, 0.1767557, 0.1388504, 0.09566507, 0.1689519, 0.143431, 
    0.1815917, 0.2170109, 0.1769481, 0.1014677, 0.1246724,
  0.2325224, 0.2257501, 0.140246, 0.2036638, 0.2193489, 0.2557566, 0.1600768, 
    0.03760476, 0.04215766, 0.05754764, 0.06233681, 0.1088561, 0.1620322, 
    0.2245736, 0.2240986, 0.192863, 0.1776962, 0.1656446, 0.1571833, 
    0.134663, 0.08887643, 0.1726498, 0.217925, 0.2294462, 0.2090256, 
    0.1805608, 0.18318, 0.2071785, 0.2248949,
  0.2415639, 0.1592842, 0.1975985, 0.204599, 0.1593525, 0.2548713, 0.3482215, 
    0.3058872, 0.2397597, 0.1826973, 0.06108619, 0.03188298, 0.06885274, 
    0.1711272, 0.2025883, 0.1879485, 0.204429, 0.282384, 0.1970424, 
    0.1169728, 0.1497613, 0.1317974, 0.1001095, 0.1372093, 0.1709851, 
    0.2388951, 0.2423456, 0.2680581, 0.2079051,
  0.1771683, 0.1487595, 0.1237862, 0.1436534, 0.1608403, 0.1225666, 
    0.1583246, 0.1685775, 0.1191452, 0.09692183, 0.06340063, 0.06640226, 
    0.1007537, 0.1174967, 0.1059816, 0.09683473, 0.1712703, 0.2367359, 
    0.2283995, 0.2067778, 0.1383189, 0.08559977, 0.05248945, 0.02404233, 
    0.09635182, 0.009781275, 0.0007245869, 0.1145863, 0.1181562,
  0.113822, 0.1265402, 0.1052709, 0.08590253, 0.03158053, 0.005755039, 
    0.008731985, 0.01197851, 0.02606824, 0.04147053, 0.02910485, 0.01809144, 
    0.02348166, 0.04156121, 0.04650262, 0.03600617, 0.03029356, 0.0313984, 
    0.032144, 0.01389937, 0.01892279, 0.02643816, 0.002637326, 0.001732436, 
    -0.0004938119, -2.299707e-05, -0.001478009, 0.0296126, 0.1222018,
  0.01148348, 0.01084707, 0.01021065, 0.009574234, 0.008937817, 0.0083014, 
    0.007664983, 0.009919872, 0.01008539, 0.0102509, 0.01041641, 0.01058193, 
    0.01074744, 0.01091296, 0.01099973, 0.01195054, 0.01290135, 0.01385215, 
    0.01480296, 0.01575377, 0.01670458, 0.01447431, 0.01399441, 0.01351451, 
    0.0130346, 0.0125547, 0.01207479, 0.01159489, 0.01199262,
  0.03299177, 0.01067059, 0.006971766, 0.002198238, 0.0001564488, 
    0.0005511909, -0.0002052186, -2.077182e-05, 0.0001629186, 0.00735247, 
    0.008045964, 0.00765242, 0.00713843, 0.1440597, 0.1359539, 0.216781, 
    0.2729087, 0.2637413, 0.2187427, 0.1775541, 0.145515, 0.1114813, 
    0.1624877, 0.08710975, 0.05805559, 0.03383469, 0.07924269, 0.1356549, 
    0.0664878,
  0.1754701, 0.2198712, 0.1240297, 0.1498454, 0.1706925, 0.1792395, 
    0.1920996, 0.1568677, 0.129507, 0.1214382, 0.08565357, 0.1260315, 
    0.1762466, 0.2712752, 0.247927, 0.190944, 0.1534963, 0.2283228, 
    0.1686182, 0.2351212, 0.2734725, 0.2097168, 0.3165017, 0.2344975, 
    0.2397872, 0.1861376, 0.1226803, 0.1222135, 0.2651469,
  0.2085195, 0.1897567, 0.2636276, 0.2287344, 0.1907293, 0.2139717, 
    0.2024626, 0.2285704, 0.2442843, 0.2550581, 0.2311536, 0.2166933, 
    0.2320687, 0.2459752, 0.1994011, 0.1948239, 0.1794183, 0.1515035, 
    0.1708049, 0.2141497, 0.2063373, 0.2640043, 0.2515636, 0.2260007, 
    0.239879, 0.2322613, 0.2200016, 0.2397767, 0.270768,
  0.1601744, 0.1696905, 0.1548041, 0.1737029, 0.1767206, 0.1925288, 
    0.1563125, 0.1320073, 0.1405621, 0.1530012, 0.16106, 0.1144539, 
    0.1299584, 0.2148651, 0.1688591, 0.087854, 0.1171137, 0.104165, 
    0.08017207, 0.1354391, 0.1402871, 0.1955613, 0.188981, 0.1500822, 
    0.1022718, 0.1222266, 0.1154405, 0.09756559, 0.156202,
  0.0394396, 0.02493536, 0.01262932, 0.07642798, 0.05533287, 0.04417873, 
    0.0453956, 0.04110011, 0.03511723, 0.009391136, 0.03920792, 0.07111765, 
    0.08255239, 0.05933802, 0.03528465, 0.0139335, 0.07575022, 0.08591814, 
    0.1326288, 0.1363207, 0.05792666, 0.037351, 0.02507683, 0.01365087, 
    0.07869612, 0.06963263, 0.07839934, 0.09219442, 0.05173656,
  0.0007870634, 0.001137973, 0.0988059, 0.03321844, 0.04314109, 0.07571819, 
    0.02199543, 0.01858189, 0.0001595851, 0.04769949, 0.03980028, 0.06122306, 
    0.06737615, 0.0114912, 0.02913054, 0.04407863, 0.06296266, 0.08416194, 
    0.108361, 0.08865574, 0.0115691, -0.0001127335, -2.211962e-07, 
    6.352721e-05, 0.03254917, 0.0643177, 0.11319, 0.002766334, 0.0002152914,
  0.001432372, 0.03964371, 0.06498201, 0.05827906, 0.07426377, 0.0340056, 
    0.04933485, -0.0001720854, 0.0007996886, 0.06375186, 0.05595139, 
    0.0848294, 0.1237133, 0.04480634, 0.03064746, 0.132053, 0.1439168, 
    0.1115914, 0.03347839, 0.004884005, -1.783862e-06, 4.968014e-09, 
    1.083409e-05, 0.01196702, 0.1222823, 0.09942365, 0.01801713, 0.006099707, 
    -0.000125278,
  0.004106004, 0.07109368, 0.2068311, 0.07211356, 0.06529069, 0.03152171, 
    0.04206904, 0.02532201, 0.01166003, 0.06858657, 0.05232995, 0.03469633, 
    0.03697456, 0.03263611, 0.08120114, 0.06929886, 0.04381299, 0.02749976, 
    0.002723227, 0.0003714165, 2.258208e-08, 1.661633e-06, 0.0002431728, 
    0.08594004, 0.2734838, 0.1228926, 0.0152086, 6.486343e-05, 1.080466e-05,
  0.07701528, 0.03797206, 0.03670583, 0.01912971, 0.02506029, 0.05750867, 
    0.1363134, 0.03132379, 0.04955726, 0.1628665, 0.04948875, 0.04001439, 
    0.06665666, 0.0831778, 0.06603926, 0.009883557, 0.006115698, 0.003242685, 
    0.0008756993, 0.0001998996, 0.00534929, 0.02330712, 0.0455133, 
    0.04594085, 0.137809, 0.186658, 0.02795074, 0.004656931, 0.02178822,
  -0.0001836997, 3.088935e-06, 7.257445e-07, 9.122909e-06, 0.01586071, 
    0.01846246, 0.02331835, 0.05737633, 0.001856547, 0.04940958, 0.08559138, 
    0.08513565, 0.07631355, 0.02384973, 0.00657073, 0.01533542, 0.04133564, 
    0.03110201, 0.04022384, 0.05102812, 0.06343662, 0.02192917, 0.003024179, 
    0.002449979, 0.006034041, 0.01266449, 0.004649759, 5.730077e-05, 
    0.02585008,
  0.02621205, -2.674194e-06, 1.004289e-06, 7.229545e-06, 1.294096e-06, 
    0.0006174613, 0.01081446, 0.004261745, 0.01771726, 0.02398053, 
    0.05797849, 0.06671988, 0.03161547, 0.002359, 2.026361e-06, 0.000466326, 
    0.03063532, 0.01215235, 0.003042747, 0.05015796, 0.02990671, 0.0157338, 
    0.01399859, 0.0004003388, 0.008388474, 0.02784275, 0.003815194, 
    0.008904736, 0.0230452,
  0.001146031, 0.004561693, 0.01352249, 0.02013539, 0.02773834, 0.002592017, 
    0.01946158, 0.02247049, 0.04461545, 0.141794, 0.06133053, 0.06550358, 
    0.05500742, 0.1105677, 0.127322, 0.08564201, 0.1050134, 0.1270723, 
    0.03903198, 0.003162025, 0.06406317, 0.04713114, 0.06674259, 0.05218272, 
    0.05840268, 0.07073282, 0.04887053, 0.02795419, 0.01782071,
  0.09776167, 0.0684008, 0.1786643, 0.2919958, 0.09856673, 0.1159571, 
    0.2234559, 0.09941402, 0.07657077, 0.06898059, 0.05616269, 0.1208866, 
    0.1267768, 0.1440281, 0.1782975, 0.187305, 0.221752, 0.2174607, 
    0.1255524, 0.1848238, 0.1539693, 0.08615431, 0.1529962, 0.1441935, 
    0.1740407, 0.2059964, 0.158612, 0.09021474, 0.1093525,
  0.2074292, 0.2147984, 0.1467971, 0.2095408, 0.2208343, 0.2511233, 
    0.1747195, 0.1003075, 0.09439665, 0.08216259, 0.07244429, 0.162655, 
    0.1838746, 0.229746, 0.2310344, 0.1942955, 0.171519, 0.1631384, 
    0.1358566, 0.1562543, 0.1028861, 0.1883202, 0.247181, 0.2665979, 
    0.2245895, 0.1932623, 0.1813242, 0.1915862, 0.2135458,
  0.2357862, 0.1694634, 0.2017376, 0.2322056, 0.1989859, 0.321992, 0.3597621, 
    0.3265167, 0.2563258, 0.22198, 0.1228854, 0.07140446, 0.09857292, 
    0.2112505, 0.217137, 0.2134111, 0.224807, 0.2956786, 0.2349637, 0.128427, 
    0.1549535, 0.1522876, 0.1342156, 0.1679769, 0.1839594, 0.2947657, 
    0.2553675, 0.2538448, 0.1983496,
  0.2067496, 0.2100583, 0.1606645, 0.2117955, 0.1701771, 0.1588372, 
    0.2275031, 0.2377463, 0.1785445, 0.1468288, 0.0936083, 0.1156301, 
    0.1414226, 0.1728108, 0.1404699, 0.1133888, 0.2136181, 0.2839905, 
    0.3019959, 0.225736, 0.1321269, 0.09300208, 0.08456852, 0.07617912, 
    0.165152, 0.02494347, 0.00551026, 0.1482674, 0.1329422,
  0.1863671, 0.2100021, 0.1634428, 0.1136129, 0.07119134, 0.07212947, 
    0.06546219, 0.07225963, 0.0817211, 0.08091538, 0.0489205, 0.03538568, 
    0.06381378, 0.09967716, 0.1199267, 0.1238175, 0.1016457, 0.06093057, 
    0.06516902, 0.05958632, 0.04370208, 0.04878989, 0.01679549, 0.0004201932, 
    0.0008576869, -1.16084e-05, -0.0100381, 0.09361554, 0.2027184,
  0.01904568, 0.01898508, 0.01892448, 0.01886388, 0.01880327, 0.01874267, 
    0.01868207, 0.02189944, 0.02224447, 0.02258949, 0.02293452, 0.02327955, 
    0.02362457, 0.0239696, 0.02389471, 0.02384642, 0.02379812, 0.02374983, 
    0.02370153, 0.02365324, 0.02360495, 0.02154131, 0.02130518, 0.02106906, 
    0.02083293, 0.0205968, 0.02036067, 0.02012454, 0.01909417,
  0.1049126, 0.04149325, 0.01474444, 0.01629763, 0.01252931, 0.007054068, 
    0.008510007, 0.00352569, 0.006646234, 0.01017048, 0.007129486, 
    0.01707035, 0.02975081, 0.1400236, 0.1546413, 0.2142356, 0.2631974, 
    0.2909117, 0.2235021, 0.2396763, 0.2019867, 0.1779379, 0.1775461, 
    0.06406161, 0.04269731, 0.03003873, 0.08409899, 0.1483038, 0.1536228,
  0.1890748, 0.2111221, 0.1305604, 0.1446592, 0.2139082, 0.222876, 0.2002559, 
    0.2065875, 0.1891167, 0.1594861, 0.1988028, 0.1898505, 0.1800737, 
    0.272061, 0.24729, 0.2247412, 0.1710652, 0.2425363, 0.1947095, 0.237791, 
    0.2905989, 0.2306052, 0.3390667, 0.2612231, 0.2600795, 0.2023457, 
    0.1265075, 0.1449569, 0.2759496,
  0.2313931, 0.2233999, 0.2799427, 0.2649921, 0.2220896, 0.2443812, 
    0.2260143, 0.2581242, 0.265782, 0.2745729, 0.2414782, 0.2320388, 
    0.2554101, 0.2433315, 0.2032712, 0.1921791, 0.188051, 0.1946018, 
    0.2045984, 0.2211089, 0.2476425, 0.2781207, 0.2421446, 0.2230633, 
    0.2323931, 0.224531, 0.2170106, 0.265579, 0.2837085,
  0.1608867, 0.1631839, 0.1853819, 0.1979931, 0.1967284, 0.2022829, 
    0.1594834, 0.1271785, 0.1402552, 0.1628524, 0.169146, 0.1284967, 
    0.1364565, 0.210622, 0.1838125, 0.09478433, 0.1143387, 0.1040009, 
    0.09136839, 0.1258179, 0.1468145, 0.1898718, 0.1980754, 0.1433302, 
    0.1035254, 0.1253677, 0.1239063, 0.1100286, 0.1733701,
  0.0443522, 0.02242914, 0.011762, 0.07529983, 0.05430831, 0.04313522, 
    0.05020999, 0.03832633, 0.03187136, 0.008768789, 0.02783738, 0.06774272, 
    0.08163725, 0.05920026, 0.03035634, 0.01321741, 0.06012659, 0.07901132, 
    0.1406134, 0.141122, 0.04512724, 0.03616688, 0.02321626, 0.01372566, 
    0.07652164, 0.06953017, 0.07541387, 0.07952943, 0.05241151,
  0.001507404, 0.0001088014, 0.1155848, 0.0394088, 0.04096057, 0.07301126, 
    0.01893743, 0.02141423, 2.558691e-06, 0.0495209, 0.04965128, 0.04489094, 
    0.07070417, 0.008565194, 0.03095619, 0.04160551, 0.05986456, 0.07614838, 
    0.09291111, 0.09172927, 0.01246645, -7.815619e-05, -1.532535e-08, 
    0.0002480724, 0.02977567, 0.06788664, 0.1223363, 0.004137083, 6.122201e-05,
  2.8536e-05, 0.05189998, 0.07809118, 0.06047444, 0.09096429, 0.04289777, 
    0.05674207, -2.658553e-05, 0.004672711, 0.08598965, 0.07990769, 
    0.09114972, 0.137778, 0.05194964, 0.04006229, 0.1752709, 0.1636558, 
    0.1280817, 0.02989605, 0.005633198, 6.302403e-06, 4.229425e-08, 
    2.532735e-05, 0.009180138, 0.150909, 0.1050913, 0.01943134, 4.005117e-05, 
    -2.343117e-05,
  0.01593148, 0.1111404, 0.2429576, 0.1065891, 0.08507048, 0.03931964, 
    0.05133881, 0.02805401, 0.01743692, 0.08902004, 0.06107321, 0.04935142, 
    0.05874363, 0.04165124, 0.09598193, 0.08430016, 0.05686165, 0.02670597, 
    0.003362959, 0.0005713461, 3.690554e-07, 5.32855e-06, 0.0001016479, 
    0.09820387, 0.3280831, 0.1343958, 0.01775429, 0.0001617934, 0.002995082,
  0.1098894, 0.04844059, 0.04688537, 0.02153377, 0.02428185, 0.05754101, 
    0.1349051, 0.03300863, 0.04922026, 0.1934097, 0.05682785, 0.04634556, 
    0.07667488, 0.09226911, 0.06786496, 0.01112089, 0.006030938, 0.001016587, 
    0.0001660404, 0.001020944, 0.01524212, 0.04712105, 0.05919892, 
    0.04750685, 0.1368207, 0.1794953, 0.03458974, 0.004057286, 0.03020487,
  -0.000112544, 1.078456e-06, 5.548826e-05, 9.606106e-05, 0.020441, 
    0.02332621, 0.0284696, 0.06353813, 0.002340239, 0.06454074, 0.1069154, 
    0.0984426, 0.08337122, 0.02951014, 0.007503385, 0.01709178, 0.04087922, 
    0.02285281, 0.04041324, 0.05293049, 0.06719175, 0.02336167, 0.003997164, 
    0.002480487, 0.004618309, 0.00394439, -0.0002967978, -5.004551e-05, 
    0.02299049,
  0.01464648, 7.667414e-07, 1.6345e-06, 8.465254e-05, 1.362029e-06, 
    0.0005737987, 0.008282263, 0.002063762, 0.01510391, 0.01569722, 
    0.05985725, 0.06604972, 0.03624276, 0.0002890535, -7.955031e-06, 
    0.0005839164, 0.03021595, 0.007683965, 0.001055195, 0.04079899, 
    0.03306777, 0.01868667, 0.03031251, 0.0006793452, 0.01247266, 0.02850896, 
    0.002894673, 0.001787781, 0.03719058,
  0.0006173832, 0.007832245, 0.01683483, 0.01404533, 0.03208986, 0.006164211, 
    0.01657737, 0.02809685, 0.07892045, 0.137257, 0.0706545, 0.05986376, 
    0.06040059, 0.1109621, 0.1310126, 0.102822, 0.1036616, 0.1166377, 
    0.0305783, 0.003038174, 0.06114623, 0.0503143, 0.06975636, 0.05534814, 
    0.05884135, 0.07039314, 0.04815378, 0.02237024, 0.01287248,
  0.08315824, 0.07216101, 0.1872003, 0.2970633, 0.09431961, 0.09722494, 
    0.2565162, 0.08061596, 0.06690364, 0.05974423, 0.0592456, 0.1194784, 
    0.1291867, 0.1440903, 0.1887597, 0.1994582, 0.2301921, 0.2212126, 
    0.1222607, 0.1825544, 0.1732565, 0.08452389, 0.1496105, 0.146965, 
    0.1753334, 0.1915258, 0.1487051, 0.08580188, 0.1081711,
  0.1903565, 0.2095529, 0.1597869, 0.2180853, 0.2136678, 0.23562, 0.1711998, 
    0.1296005, 0.1286006, 0.08046051, 0.07380112, 0.1953932, 0.189147, 
    0.2197338, 0.2375269, 0.18313, 0.1477957, 0.1478195, 0.1270642, 
    0.1710088, 0.116684, 0.1796332, 0.2518377, 0.2955228, 0.2217337, 
    0.2009041, 0.1811214, 0.1787771, 0.2161673,
  0.2186895, 0.1754695, 0.1988313, 0.2763752, 0.2116182, 0.3187429, 
    0.3511314, 0.3494738, 0.2833569, 0.2636508, 0.1763273, 0.1154058, 
    0.1427885, 0.219875, 0.2471177, 0.2097912, 0.234613, 0.3002555, 
    0.2436489, 0.1799316, 0.1703065, 0.1675339, 0.1638412, 0.2363609, 
    0.2042723, 0.3136022, 0.2418067, 0.2467894, 0.2112162,
  0.2190998, 0.2103181, 0.2199504, 0.2541224, 0.187195, 0.2183325, 0.2689848, 
    0.2935475, 0.2357515, 0.2221468, 0.1509293, 0.1700349, 0.1910942, 
    0.2163936, 0.1885609, 0.1443994, 0.2520107, 0.3079169, 0.330208, 
    0.2370291, 0.1504222, 0.1113004, 0.09157678, 0.1090664, 0.2186158, 
    0.05810253, 0.0129523, 0.1584749, 0.136278,
  0.2316949, 0.2605951, 0.1847143, 0.1556765, 0.1245208, 0.1266825, 
    0.1407191, 0.1265021, 0.1018322, 0.108089, 0.08710889, 0.08641488, 
    0.1007287, 0.1229802, 0.1712107, 0.1676077, 0.1285186, 0.08980867, 
    0.08000895, 0.08281392, 0.08419864, 0.0936672, 0.0577824, 0.01684794, 
    0.02051697, 0.003674378, 0.00923533, 0.178513, 0.2466534,
  0.03891264, 0.03889621, 0.03887978, 0.03886335, 0.03884692, 0.03883049, 
    0.03881406, 0.04079556, 0.04095547, 0.04111537, 0.04127528, 0.04143519, 
    0.04159509, 0.041755, 0.03099877, 0.03221276, 0.03342675, 0.03464073, 
    0.03585472, 0.03706871, 0.0382827, 0.04756962, 0.04621216, 0.0448547, 
    0.04349723, 0.04213977, 0.04078231, 0.03942484, 0.03892579,
  0.2106388, 0.11329, 0.02016304, 0.01933945, 0.02170233, 0.01654405, 
    0.01467285, 0.01333711, 0.01030625, 0.01109948, 0.02035518, 0.02505407, 
    0.06856512, 0.1566496, 0.1819866, 0.2557654, 0.275002, 0.2894351, 
    0.2241338, 0.2630449, 0.2105266, 0.1988454, 0.159103, 0.03996059, 
    0.03556804, 0.02973454, 0.09656505, 0.1710184, 0.1530281,
  0.2037833, 0.2173391, 0.1601488, 0.1467938, 0.227515, 0.2458337, 0.2057652, 
    0.2411592, 0.2170717, 0.2114127, 0.2680973, 0.2111836, 0.1740334, 
    0.2860371, 0.2469024, 0.2403947, 0.2011138, 0.2522556, 0.1681589, 
    0.266115, 0.2747712, 0.2618349, 0.3008527, 0.2659944, 0.2640253, 
    0.2120909, 0.1504427, 0.1818945, 0.2920422,
  0.2666222, 0.2797279, 0.2819447, 0.3258684, 0.2860134, 0.2864687, 
    0.2548013, 0.3150563, 0.2934246, 0.2966284, 0.2428176, 0.2552988, 
    0.2526571, 0.2203067, 0.2034458, 0.1769296, 0.2000152, 0.1942227, 
    0.2213145, 0.232142, 0.2596954, 0.2757457, 0.2756249, 0.2516747, 
    0.2460232, 0.2484493, 0.220098, 0.2646943, 0.2902093,
  0.1607803, 0.181174, 0.195888, 0.2016734, 0.1955389, 0.2060373, 0.1701571, 
    0.1375359, 0.1426033, 0.1675147, 0.161378, 0.1454274, 0.1483006, 
    0.2186591, 0.1861487, 0.1112354, 0.1005287, 0.1080233, 0.1013075, 
    0.1354673, 0.153808, 0.206498, 0.1793082, 0.1385257, 0.1054755, 
    0.1222723, 0.1182203, 0.1250921, 0.1578115,
  0.0471523, 0.01951052, 0.01531332, 0.07922739, 0.05302051, 0.04950792, 
    0.05380978, 0.04154422, 0.03893411, 0.00800867, 0.02324626, 0.0666781, 
    0.08381303, 0.06210323, 0.03644583, 0.01392736, 0.05178529, 0.07672894, 
    0.1526744, 0.146898, 0.04734291, 0.04206247, 0.01474441, 0.02311006, 
    0.07329445, 0.08330343, 0.07960714, 0.07679363, 0.0580044,
  0.002713626, 0.0002564263, 0.1255968, 0.03848125, 0.03884075, 0.06400224, 
    0.01731885, 0.02141605, -3.340358e-05, 0.05109114, 0.0532153, 0.05686431, 
    0.07736997, 0.007073202, 0.03343874, 0.03924978, 0.0620483, 0.09506446, 
    0.08896132, 0.09146349, 0.01570187, 0.0001242826, 5.545193e-08, 
    0.0006826849, 0.03766985, 0.07527218, 0.1415368, 0.01132462, 0.0001300757,
  2.082177e-06, 0.08479437, 0.0966875, 0.06584098, 0.107596, 0.05434879, 
    0.06852293, 2.96791e-05, 0.005922603, 0.09085634, 0.08835769, 0.1074525, 
    0.1373666, 0.05204334, 0.03967794, 0.2074998, 0.1854682, 0.1635975, 
    0.03185419, 0.009381209, 4.378741e-05, 5.639311e-08, 1.580228e-05, 
    0.006036702, 0.1861067, 0.1251281, 0.01932554, 1.82717e-05, -5.528535e-06,
  0.01298102, 0.08930556, 0.3090372, 0.1502007, 0.08882123, 0.05148899, 
    0.06433603, 0.03287561, 0.02000545, 0.1108905, 0.07683061, 0.05733088, 
    0.08266951, 0.04759197, 0.09881385, 0.1001531, 0.06139482, 0.02492072, 
    0.003355471, 0.0003877811, 2.278054e-07, 2.815191e-05, 0.0001432407, 
    0.125709, 0.397595, 0.1676351, 0.01755723, 9.745824e-05, 0.000445049,
  0.1370217, 0.0575203, 0.05357446, 0.02340709, 0.02224521, 0.05562468, 
    0.1379845, 0.04033077, 0.06785776, 0.2304582, 0.06852729, 0.05631727, 
    0.08020329, 0.0946668, 0.07760868, 0.01054263, 0.008868206, 0.0002105165, 
    5.674357e-05, 0.0009379532, 0.005538797, 0.05207732, 0.0864925, 
    0.06245112, 0.1652887, 0.1841868, 0.03967372, 0.003297281, 0.04453504,
  -6.107587e-06, 6.529136e-06, 0.0004678597, 0.002573418, 0.02323324, 
    0.02695203, 0.02912701, 0.07333523, 0.004124898, 0.06783341, 0.1253994, 
    0.1059938, 0.08434963, 0.03611513, 0.01595015, 0.02152088, 0.04849721, 
    0.02255024, 0.04110825, 0.05302146, 0.06912431, 0.02509989, 0.006301481, 
    0.003886922, 0.006746395, 0.001868323, -0.0003968222, 0.0004513122, 
    0.01664851,
  0.004669103, 7.293687e-07, 1.15407e-06, 0.001037897, 7.285564e-07, 
    0.002297821, 0.008518772, 0.01017733, 0.01159394, 0.01528617, 0.0694719, 
    0.06990715, 0.04390378, 0.0008867495, 0.0002723596, 0.0007618601, 
    0.03447857, 0.006713401, 0.002004434, 0.04237691, 0.04011223, 0.03006429, 
    0.04068696, 0.00282474, 0.01849855, 0.03684346, 0.001635216, 0.001927372, 
    0.05032307,
  0.00221648, 0.01782319, 0.02099095, 0.01354362, 0.03722752, 0.01091794, 
    0.01329181, 0.02204922, 0.1161651, 0.1397404, 0.06640045, 0.05856602, 
    0.06254852, 0.1179882, 0.1280568, 0.1139476, 0.09943588, 0.1081656, 
    0.03181662, 0.007548612, 0.05868979, 0.05950449, 0.07009435, 0.05809622, 
    0.06199151, 0.07559128, 0.05038058, 0.01442994, 0.02301786,
  0.06504592, 0.07509985, 0.1906849, 0.3110239, 0.0904608, 0.08067933, 
    0.2650362, 0.05887866, 0.05891825, 0.04563661, 0.06013925, 0.1072508, 
    0.1233169, 0.1428666, 0.2082781, 0.2044459, 0.2250613, 0.2143345, 
    0.1188109, 0.1787755, 0.1789747, 0.08672609, 0.139501, 0.127355, 
    0.1750509, 0.182225, 0.1475306, 0.07845533, 0.1020987,
  0.2023272, 0.2154733, 0.1412634, 0.2110185, 0.1991048, 0.2176468, 
    0.1585768, 0.1445382, 0.1268773, 0.07061659, 0.07144897, 0.202953, 
    0.1831188, 0.2215938, 0.2427111, 0.1764134, 0.1416919, 0.1470759, 
    0.1212491, 0.1828482, 0.1232074, 0.1648937, 0.2646954, 0.3373699, 
    0.2399653, 0.1864924, 0.1846142, 0.1716742, 0.2062998,
  0.2155248, 0.1717704, 0.2059799, 0.3099162, 0.2285055, 0.3135114, 
    0.3438784, 0.3424845, 0.2855931, 0.3047984, 0.2030463, 0.1395041, 
    0.1603429, 0.2261986, 0.2609336, 0.2128959, 0.2250635, 0.3092806, 
    0.2482404, 0.1974884, 0.1853664, 0.1727579, 0.1778706, 0.2817441, 
    0.2171506, 0.3347486, 0.2471612, 0.2648219, 0.2155512,
  0.2110611, 0.1906535, 0.2269685, 0.2657447, 0.2529628, 0.2796251, 
    0.2666152, 0.334517, 0.260036, 0.2525482, 0.1714602, 0.2031191, 0.200021, 
    0.2294652, 0.1870827, 0.1373136, 0.273232, 0.3203533, 0.3268351, 
    0.2523783, 0.1762139, 0.1333912, 0.1221045, 0.1504623, 0.2286613, 
    0.1329075, 0.03281054, 0.1744022, 0.1494756,
  0.2262275, 0.2631178, 0.221701, 0.1855351, 0.1851633, 0.1749035, 0.1899498, 
    0.1737367, 0.1525566, 0.154942, 0.1603507, 0.1426074, 0.126007, 
    0.1645913, 0.2242074, 0.2191068, 0.1780045, 0.1313348, 0.118523, 
    0.1096191, 0.1193948, 0.1672215, 0.1156256, 0.04393728, 0.06630433, 
    0.01000429, 0.06665596, 0.2413312, 0.2462616,
  0.06072867, 0.06006814, 0.05940761, 0.05874708, 0.05808656, 0.05742603, 
    0.0567655, 0.0571702, 0.06203046, 0.06689072, 0.07175098, 0.07661124, 
    0.08147149, 0.08633175, 0.09052213, 0.09012004, 0.08971795, 0.08931586, 
    0.08891377, 0.08851169, 0.0881096, 0.0888679, 0.08507025, 0.08127262, 
    0.07747497, 0.07367733, 0.0698797, 0.06608205, 0.06125709,
  0.2102692, 0.1796487, 0.08086099, 0.02384726, 0.03101099, 0.02704925, 
    0.01303085, 0.01698169, 0.01792557, 0.05481141, 0.03033827, 0.07845104, 
    0.1218798, 0.1583936, 0.179069, 0.2127394, 0.2715108, 0.3100536, 
    0.2352102, 0.2869848, 0.2125191, 0.207839, 0.1537741, 0.02326836, 
    0.04985666, 0.02716279, 0.1102555, 0.1852256, 0.1594143,
  0.2335084, 0.2336587, 0.1918712, 0.1653459, 0.2463964, 0.2406893, 
    0.2194254, 0.2561872, 0.2580751, 0.2342227, 0.2684928, 0.2073933, 
    0.1940394, 0.2922777, 0.2810972, 0.2422445, 0.2661856, 0.3141918, 
    0.2141995, 0.3296415, 0.2879508, 0.2875753, 0.297951, 0.2801419, 
    0.2461048, 0.1664115, 0.1308726, 0.180584, 0.28849,
  0.2792555, 0.329867, 0.3151578, 0.3531658, 0.2940529, 0.2650297, 0.2755976, 
    0.3257652, 0.30046, 0.3031304, 0.2601645, 0.2659735, 0.2459435, 
    0.2330439, 0.2130966, 0.1986935, 0.2325879, 0.2134036, 0.254523, 
    0.2414593, 0.2387869, 0.2585335, 0.2453083, 0.2290877, 0.2278768, 
    0.2270849, 0.2037471, 0.2636667, 0.2860893,
  0.2030962, 0.1853454, 0.2173193, 0.2109875, 0.2081707, 0.216635, 0.1741495, 
    0.1486655, 0.1490644, 0.1583187, 0.170365, 0.1510006, 0.1571167, 
    0.2176981, 0.1800565, 0.1251128, 0.09815328, 0.1072734, 0.1090236, 
    0.1284948, 0.1606643, 0.2107978, 0.1756783, 0.1427275, 0.1143351, 
    0.1160797, 0.1230895, 0.1355548, 0.1750341,
  0.05271239, 0.01843768, 0.01954096, 0.07068171, 0.06197153, 0.05474711, 
    0.05863437, 0.04522454, 0.04630841, 0.008094497, 0.02186601, 0.06401968, 
    0.08327711, 0.06243775, 0.04634653, 0.01412964, 0.05843268, 0.08319347, 
    0.1654123, 0.1496703, 0.0517754, 0.04058042, 0.01220402, 0.02440946, 
    0.06274489, 0.08884341, 0.09054422, 0.09337141, 0.06783158,
  0.003511361, 0.002400449, 0.1322135, 0.03825381, 0.03402477, 0.05826791, 
    0.0215074, 0.02733072, -5.409219e-06, 0.03321799, 0.02920097, 0.04017639, 
    0.09093787, 0.005097139, 0.03929711, 0.05303659, 0.0775457, 0.1117388, 
    0.09413982, 0.09386955, 0.01860796, 0.0003158704, 3.64977e-07, 
    0.001056295, 0.04824902, 0.08694584, 0.1498971, 0.01423458, 0.0006459106,
  0.0009671124, 0.1158045, 0.1343273, 0.05412763, 0.1074966, 0.04356823, 
    0.06647299, 0.001704834, 0.001222919, 0.06383767, 0.08047586, 0.1145457, 
    0.1167148, 0.03673977, 0.04012883, 0.2041357, 0.1607724, 0.1588893, 
    0.03316431, 0.01141287, 0.0007276304, 9.489364e-08, 4.138476e-06, 
    0.001611388, 0.1686101, 0.1386492, 0.01950425, 0.0002454816, -4.030248e-06,
  0.001134851, 0.032267, 0.3654505, 0.1620139, 0.07913937, 0.05290084, 
    0.06106122, 0.03847653, 0.01379984, 0.08880658, 0.07352151, 0.03705214, 
    0.06801435, 0.03967281, 0.0744766, 0.09232134, 0.06042831, 0.02416404, 
    0.004465044, 0.0003928256, 6.887429e-08, 3.878705e-06, 6.379405e-05, 
    0.1313705, 0.3796542, 0.1895833, 0.01817307, 0.0002360107, 0.003328523,
  0.08495417, 0.08096617, 0.04224023, 0.02364374, 0.02472511, 0.05804189, 
    0.1363789, 0.03443133, 0.08334795, 0.2678005, 0.06407856, 0.04633466, 
    0.0629371, 0.08365202, 0.07689382, 0.008693945, 0.006745365, 
    0.0001080764, 0.00033994, 0.002265996, 0.002309696, 0.07350244, 
    0.1097933, 0.07511806, 0.1553132, 0.1764752, 0.04288218, 0.005243167, 
    0.03539415,
  -7.830514e-07, 4.04095e-05, 0.0003272698, 0.03201629, 0.02216133, 
    0.02283153, 0.02599568, 0.0752894, 0.007810755, 0.068111, 0.1376039, 
    0.09943514, 0.07055305, 0.03496436, 0.02630667, 0.02253909, 0.05434789, 
    0.02249227, 0.0427928, 0.05321489, 0.06761354, 0.02459719, 0.01321164, 
    0.006807699, 0.008003536, 0.004997733, -0.0001178805, 0.0001952793, 
    0.01486495,
  6.860706e-05, 3.020967e-06, 6.443022e-07, 0.001489186, 1.925219e-06, 
    0.00334415, 0.01383451, 0.0139958, 0.007861924, 0.02370603, 0.08024056, 
    0.07902263, 0.0400896, 0.0002354144, 0.0006711126, 0.00123832, 
    0.03801376, 0.008882338, 0.001169993, 0.06137821, 0.04270018, 0.04641514, 
    0.04514528, 0.0100051, 0.02376087, 0.04295696, 0.002297323, 0.006875994, 
    0.04257021,
  0.003527299, 0.01894638, 0.01688115, 0.01079658, 0.04848114, 0.0148704, 
    0.01088562, 0.01611885, 0.1367828, 0.1485138, 0.07118479, 0.05951456, 
    0.06787921, 0.1364926, 0.1188523, 0.1162226, 0.09234074, 0.1029415, 
    0.03507855, 0.01409174, 0.05494053, 0.06438992, 0.07439582, 0.05226669, 
    0.06546214, 0.08460873, 0.05641749, 0.014448, 0.02390674,
  0.05730102, 0.0713068, 0.1816231, 0.3265368, 0.1045056, 0.06730305, 
    0.2763313, 0.04332682, 0.04655249, 0.03979207, 0.06555641, 0.1005168, 
    0.131063, 0.1545303, 0.208287, 0.2102973, 0.2118438, 0.2056172, 
    0.1104172, 0.18547, 0.1789438, 0.0854249, 0.160827, 0.1328087, 0.1688794, 
    0.1772086, 0.1516541, 0.07341986, 0.09181784,
  0.188303, 0.2040866, 0.1751364, 0.2059724, 0.1909026, 0.2185762, 0.1478522, 
    0.1450786, 0.1328089, 0.0645079, 0.06807632, 0.1892271, 0.1832204, 
    0.2199264, 0.2410669, 0.1726579, 0.130259, 0.1421573, 0.1165815, 
    0.1729953, 0.1407808, 0.177145, 0.2644385, 0.3179301, 0.2619296, 
    0.1878839, 0.1752584, 0.1694574, 0.2041015,
  0.2126917, 0.1803681, 0.2277033, 0.33097, 0.2262794, 0.315073, 0.3305873, 
    0.3305048, 0.2737159, 0.3035619, 0.2075684, 0.1626222, 0.1636377, 
    0.2300322, 0.2571212, 0.2055201, 0.2227671, 0.3094877, 0.2539698, 
    0.1844876, 0.1943253, 0.1820402, 0.2307378, 0.3222439, 0.2155765, 
    0.3368441, 0.2667812, 0.285749, 0.2169599,
  0.215263, 0.1871156, 0.240357, 0.2851777, 0.2709115, 0.3000754, 0.2860516, 
    0.3688563, 0.2763247, 0.2698105, 0.2039122, 0.2202544, 0.2414903, 
    0.2185298, 0.1869055, 0.1433384, 0.2822834, 0.3278638, 0.3045242, 
    0.2798356, 0.1843211, 0.1567335, 0.1303644, 0.17635, 0.2223008, 
    0.2196346, 0.06667665, 0.1866715, 0.1518314,
  0.2062817, 0.2422684, 0.2229096, 0.1946633, 0.1894218, 0.1830821, 0.178086, 
    0.1791883, 0.1789423, 0.167125, 0.1938781, 0.1778952, 0.1586696, 
    0.1998594, 0.2470886, 0.2619295, 0.2206519, 0.15621, 0.1367302, 
    0.1147374, 0.1510605, 0.1853389, 0.1603819, 0.05311124, 0.09950916, 
    0.03960974, 0.1120569, 0.2502472, 0.2428133,
  0.0585931, 0.06032073, 0.06204838, 0.06377602, 0.06550366, 0.06723129, 
    0.06895893, 0.06817141, 0.07381804, 0.07946469, 0.08511133, 0.09075797, 
    0.0964046, 0.1020512, 0.1258442, 0.123817, 0.1217898, 0.1197626, 
    0.1177354, 0.1157082, 0.113681, 0.09835062, 0.09300354, 0.08765647, 
    0.0823094, 0.07696231, 0.07161523, 0.06626816, 0.05721099,
  0.2062344, 0.1941845, 0.1433106, 0.08314151, 0.05580033, 0.05701768, 
    0.06401756, 0.06235341, 0.1009283, 0.1121776, 0.1280145, 0.08529896, 
    0.1284606, 0.2008358, 0.2034204, 0.2881756, 0.2453885, 0.3304929, 
    0.2050551, 0.2955313, 0.2424506, 0.2366192, 0.1543467, 0.03171689, 
    0.04264559, 0.05085519, 0.0948639, 0.1697598, 0.1504663,
  0.1992127, 0.1850953, 0.1808221, 0.1939893, 0.2403073, 0.2337344, 
    0.2277794, 0.2561337, 0.2573217, 0.2647219, 0.251686, 0.2019175, 
    0.2318857, 0.2710645, 0.2752712, 0.2404339, 0.2409129, 0.317234, 
    0.2422882, 0.3358848, 0.348989, 0.3438508, 0.307821, 0.2909106, 
    0.2333821, 0.1613982, 0.1825343, 0.2715688, 0.2985445,
  0.295896, 0.3493574, 0.3285069, 0.3695018, 0.3247463, 0.3328688, 0.3367052, 
    0.3132055, 0.3271325, 0.3389595, 0.2931318, 0.292353, 0.2723345, 
    0.258284, 0.228347, 0.2096656, 0.2118275, 0.1816992, 0.2450022, 
    0.2442115, 0.2383776, 0.2746753, 0.2374782, 0.2356589, 0.2576453, 
    0.22802, 0.2204613, 0.2714102, 0.2969706,
  0.2150572, 0.2229251, 0.2095723, 0.2181781, 0.1952155, 0.2219858, 
    0.1657267, 0.1475396, 0.1501072, 0.1654408, 0.1672471, 0.1631042, 
    0.164997, 0.2244862, 0.1836991, 0.1220722, 0.09729181, 0.1170001, 
    0.1103859, 0.1275352, 0.1885615, 0.2101132, 0.1852244, 0.1527411, 
    0.1145884, 0.1224643, 0.1404067, 0.1416437, 0.1706619,
  0.05380207, 0.02102172, 0.01999593, 0.06488977, 0.07262041, 0.05556495, 
    0.06252731, 0.06003103, 0.03598529, 0.008848022, 0.02209485, 0.05682325, 
    0.07909214, 0.0717441, 0.06066696, 0.02288442, 0.0662994, 0.08120408, 
    0.1667187, 0.1491319, 0.06278034, 0.04707934, 0.02002117, 0.03472658, 
    0.05427054, 0.09373929, 0.1001115, 0.1042217, 0.08372155,
  0.00601786, 0.003033482, 0.1404917, 0.03773762, 0.02215731, 0.04642201, 
    0.02547843, 0.01432294, 5.865447e-06, 0.01781772, 0.01001416, 0.0158291, 
    0.09423198, 0.009818874, 0.03784711, 0.05072057, 0.06688719, 0.112803, 
    0.09271795, 0.08981472, 0.02039649, 0.000898472, 3.372708e-07, 
    0.002552907, 0.04554001, 0.0658869, 0.1431508, 0.02156017, 0.002108436,
  0.0003978106, 0.101924, 0.1440392, 0.04862881, 0.09486882, 0.03970241, 
    0.05344113, 0.0006180803, 0.0005894142, 0.05509095, 0.06476462, 
    0.09600234, 0.1154444, 0.02828493, 0.03871439, 0.1959911, 0.1349207, 
    0.1298325, 0.03396538, 0.01589984, 0.003182345, 3.479595e-09, 
    1.686885e-06, 0.0004415005, 0.146616, 0.1526229, 0.02498912, 
    0.0009997585, -1.762614e-07,
  -1.853636e-05, 0.008111499, 0.3986464, 0.1120203, 0.07477543, 0.04308932, 
    0.04778763, 0.04270492, 0.01116958, 0.07490007, 0.06393587, 0.02838491, 
    0.05949698, 0.03756566, 0.07241315, 0.08968647, 0.0614998, 0.02597624, 
    0.007479875, 0.0008886643, 9.854567e-08, 1.333533e-06, 1.708823e-05, 
    0.0784343, 0.2578895, 0.1439949, 0.0221539, 0.0005637223, 9.976375e-05,
  0.03033713, 0.03808703, 0.03418661, 0.02587065, 0.02178612, 0.0640277, 
    0.1182904, 0.03492621, 0.07711742, 0.2380872, 0.06303654, 0.0359546, 
    0.0513791, 0.06643607, 0.06353997, 0.009452321, 0.01075781, 0.0001265414, 
    0.002240689, 0.005128063, 0.003689695, 0.04446666, 0.1283981, 0.05305748, 
    0.1214527, 0.1576049, 0.05027961, 0.006608478, 0.01740235,
  3.845226e-07, 2.803948e-06, 8.613578e-06, 0.1027488, 0.01992016, 
    0.03020358, 0.02019925, 0.06865962, 0.01385682, 0.05768506, 0.1529699, 
    0.09011446, 0.06129958, 0.03073898, 0.03305805, 0.02765283, 0.04905987, 
    0.02177889, 0.03615107, 0.05161422, 0.06197803, 0.02838354, 0.02492972, 
    0.01013449, 0.01132309, 0.001537091, 0.0002418159, -7.461147e-05, 
    0.0209554,
  6.852309e-06, 1.484966e-06, 2.392535e-07, 0.0022481, 0.01320047, 
    0.005018588, 0.02057523, 0.02167279, 0.009999733, 0.02076701, 0.07651163, 
    0.06180122, 0.04073384, 7.749481e-05, 0.001741359, 0.002183159, 
    0.02862006, 0.008628319, 0.001545304, 0.05573902, 0.03168543, 0.05550941, 
    0.03772471, 0.02477852, 0.02750134, 0.04717854, 0.002266493, 0.003848775, 
    0.0227142,
  0.007813468, 0.01649292, 0.0152668, 0.01042286, 0.06184432, 0.01763471, 
    0.01098699, 0.0174791, 0.1516399, 0.1577122, 0.0574515, 0.0622353, 
    0.09023869, 0.151022, 0.1186856, 0.1228589, 0.0907287, 0.09544353, 
    0.04068329, 0.01441498, 0.04505162, 0.0608168, 0.08102491, 0.05944792, 
    0.08360155, 0.09435365, 0.05945729, 0.01780471, 0.02886902,
  0.05364673, 0.06468847, 0.1811121, 0.3445622, 0.1226609, 0.05752336, 
    0.2791, 0.0363831, 0.03024867, 0.03955784, 0.06306119, 0.1012942, 
    0.1454577, 0.1587836, 0.2061263, 0.2137195, 0.198781, 0.207669, 0.122834, 
    0.1847436, 0.1838613, 0.08765172, 0.1605505, 0.1437272, 0.1792296, 
    0.1821347, 0.1708404, 0.07817758, 0.08261351,
  0.1924597, 0.2176152, 0.1838838, 0.2553084, 0.1817524, 0.2040521, 
    0.1454625, 0.1424967, 0.1362323, 0.05861834, 0.06367826, 0.1737303, 
    0.1862758, 0.234587, 0.2873564, 0.1910023, 0.1333372, 0.1462262, 
    0.1175755, 0.18264, 0.1663069, 0.1874367, 0.2634457, 0.3333939, 
    0.2727249, 0.1839636, 0.1877923, 0.1748075, 0.2091433,
  0.2332366, 0.1898276, 0.2358813, 0.3352351, 0.2476633, 0.3099115, 
    0.3297384, 0.3308028, 0.2671795, 0.2935077, 0.2047084, 0.1616655, 
    0.1723132, 0.2598381, 0.2924035, 0.2134634, 0.2320809, 0.315936, 
    0.2602818, 0.1835566, 0.1881767, 0.1953903, 0.2405409, 0.3220763, 
    0.2291355, 0.3208609, 0.2849051, 0.3009402, 0.2170579,
  0.2266667, 0.197327, 0.250386, 0.286111, 0.2747977, 0.3052946, 0.2983992, 
    0.3881045, 0.2857214, 0.2605232, 0.2170337, 0.2411266, 0.2728944, 
    0.2158273, 0.1907848, 0.1605065, 0.2968299, 0.3239073, 0.2965433, 
    0.2949028, 0.1759191, 0.1597247, 0.1664066, 0.2121292, 0.2140136, 
    0.2980812, 0.0919648, 0.2009691, 0.1621917,
  0.2052282, 0.234489, 0.2029262, 0.178778, 0.1809253, 0.1820244, 0.1802506, 
    0.2044683, 0.208778, 0.1825058, 0.2237175, 0.1975791, 0.1986235, 
    0.264012, 0.3095235, 0.3144659, 0.2604198, 0.1744077, 0.1419242, 
    0.1355271, 0.1803125, 0.2002312, 0.1593819, 0.07192487, 0.1066538, 
    0.05094521, 0.160816, 0.2380053, 0.2407746,
  0.05507351, 0.05676989, 0.05846627, 0.06016265, 0.06185903, 0.06355541, 
    0.0652518, 0.07894661, 0.08461692, 0.09028724, 0.09595755, 0.1016279, 
    0.1072982, 0.1129685, 0.1260854, 0.1245795, 0.1230737, 0.1215678, 
    0.1200619, 0.1185561, 0.1170502, 0.105474, 0.09961312, 0.09375229, 
    0.08789147, 0.08203065, 0.07616982, 0.07030899, 0.0537164,
  0.1880603, 0.1919041, 0.1762494, 0.1539585, 0.1046647, 0.1110864, 
    0.1341274, 0.1413385, 0.1034622, 0.1809304, 0.1207051, 0.09031618, 
    0.15149, 0.1587392, 0.1368158, 0.244796, 0.2804201, 0.2946615, 0.2317716, 
    0.2807907, 0.2488029, 0.2435253, 0.146835, 0.03446467, 0.04618335, 
    0.06025461, 0.08519785, 0.1417137, 0.1405503,
  0.2742921, 0.2690038, 0.1496675, 0.1897432, 0.2429021, 0.2608764, 
    0.2149297, 0.2606637, 0.2534164, 0.2743861, 0.2579433, 0.1914327, 
    0.2527979, 0.2676215, 0.2770731, 0.2878722, 0.2299942, 0.2851877, 
    0.2438027, 0.3482955, 0.3757152, 0.3493514, 0.3581481, 0.3469202, 
    0.2720756, 0.198852, 0.1882767, 0.2711636, 0.2880072,
  0.2962304, 0.3979157, 0.4192673, 0.4135737, 0.4026982, 0.3470729, 
    0.3110801, 0.3595352, 0.3247228, 0.3897575, 0.3420061, 0.3065271, 
    0.2847302, 0.267986, 0.2782398, 0.225307, 0.2777557, 0.2216791, 
    0.2834308, 0.2719454, 0.2634315, 0.2812925, 0.2727728, 0.2528009, 
    0.2562308, 0.2059636, 0.2422614, 0.2870462, 0.2918826,
  0.2326421, 0.2112666, 0.2457437, 0.250683, 0.2142271, 0.2383911, 0.1814911, 
    0.1480745, 0.1609011, 0.1849823, 0.1866795, 0.1672457, 0.1890847, 
    0.2192889, 0.197447, 0.1544346, 0.1141977, 0.1302044, 0.1432672, 
    0.1314059, 0.216555, 0.2082089, 0.1977131, 0.162862, 0.1067566, 
    0.1140362, 0.1455703, 0.1601951, 0.1868375,
  0.05783437, 0.02909673, 0.03009336, 0.07515573, 0.07162807, 0.05495366, 
    0.07918374, 0.09397592, 0.03533959, 0.01281717, 0.02855804, 0.04310047, 
    0.07593928, 0.07019867, 0.07607335, 0.04789893, 0.0756035, 0.08576527, 
    0.1487754, 0.1423843, 0.06392787, 0.05117572, 0.02900756, 0.03403697, 
    0.04878299, 0.09664536, 0.1037933, 0.1021049, 0.08644986,
  0.006864815, 0.00477449, 0.1414328, 0.03247019, 0.02432211, 0.03816465, 
    0.02906647, 0.02569853, 3.511332e-06, 0.00748045, 0.003705984, 
    0.004868968, 0.08644857, 0.01270938, 0.03973659, 0.04145616, 0.0720024, 
    0.1169596, 0.07096229, 0.0612696, 0.01603902, 0.003504364, -5.133945e-07, 
    0.001994754, 0.04317844, 0.05672577, 0.1405792, 0.02690605, 0.004090013,
  0.0002531741, 0.07925681, 0.1286393, 0.04811467, 0.09156661, 0.0398773, 
    0.04425739, 0.001278681, 0.0002225755, 0.04507839, 0.05849475, 0.0977533, 
    0.1218155, 0.02854277, 0.03851588, 0.1871966, 0.1219294, 0.1093784, 
    0.03652705, 0.03770526, 0.0100121, 8.958237e-05, 6.224028e-07, 
    -6.082996e-05, 0.1508827, 0.1280867, 0.03451457, 0.004608485, 9.615154e-07,
  -4.432397e-06, 0.007940708, 0.3375914, 0.08314575, 0.06829593, 0.03763685, 
    0.04270621, 0.04691246, 0.01413612, 0.06538157, 0.05390448, 0.02277624, 
    0.05284486, 0.03369293, 0.07151604, 0.09430129, 0.06353121, 0.03406685, 
    0.01689395, 0.004459176, 6.556299e-06, 3.255345e-07, 4.469508e-06, 
    0.07249077, 0.2102765, 0.1118027, 0.03301371, 0.0009624353, 5.593308e-06,
  0.01433103, 0.01248933, 0.02762453, 0.04924506, 0.02356387, 0.0676333, 
    0.1127366, 0.03334534, 0.09104346, 0.225619, 0.0600826, 0.03102219, 
    0.04806983, 0.05869075, 0.05382529, 0.01196601, 0.01151829, 5.777771e-05, 
    0.005330376, 0.006479631, 0.004900452, 0.03029838, 0.1124747, 0.05412387, 
    0.1113278, 0.1471917, 0.0534067, 0.01337432, 0.01333046,
  1.989709e-07, 1.1566e-06, 1.017072e-05, 0.1302587, 0.02207524, 0.04329669, 
    0.021733, 0.06610155, 0.02647894, 0.07210556, 0.1598963, 0.0906854, 
    0.05778274, 0.03223466, 0.03572597, 0.03191652, 0.04096052, 0.01795436, 
    0.02790371, 0.04909878, 0.05778503, 0.03007193, 0.04370666, 0.01759127, 
    0.02691904, 0.001205041, 0.0001621588, 1.717655e-05, 0.0195825,
  4.018557e-06, 6.94331e-07, 1.083234e-07, 0.005663037, 0.01984685, 
    0.004993026, 0.0246845, 0.0306864, 0.01390724, 0.01658547, 0.07203916, 
    0.05976622, 0.04149401, 0.001170727, 0.005721646, 0.004099539, 
    0.02627419, 0.006008917, 0.001895838, 0.04883477, 0.02055613, 0.06869341, 
    0.03386085, 0.05509192, 0.03419369, 0.04983259, 0.00255642, 0.001359827, 
    0.01731472,
  0.01130911, 0.01825157, 0.02077738, 0.01799021, 0.07236838, 0.02158894, 
    0.00972903, 0.02142519, 0.1515653, 0.1547516, 0.04907501, 0.0856148, 
    0.1009433, 0.1439156, 0.1130986, 0.1480019, 0.09390213, 0.0987391, 
    0.05063055, 0.01873409, 0.03966066, 0.06079105, 0.09003405, 0.07054047, 
    0.1029731, 0.1014655, 0.06615624, 0.02459562, 0.03011263,
  0.05737427, 0.06288701, 0.1753522, 0.3643868, 0.1345922, 0.05194299, 
    0.280631, 0.03111344, 0.01719869, 0.03363717, 0.05904951, 0.10901, 
    0.1551837, 0.1801808, 0.2096138, 0.2173923, 0.1999291, 0.2091071, 
    0.141062, 0.1917829, 0.1929045, 0.08576194, 0.1574507, 0.1474482, 
    0.1917911, 0.1852672, 0.1825655, 0.10204, 0.08408873,
  0.2063472, 0.2246018, 0.1784941, 0.2508522, 0.1759771, 0.2008252, 
    0.1358155, 0.1383895, 0.1285443, 0.05043697, 0.05231685, 0.1742465, 
    0.1921736, 0.2448995, 0.2906428, 0.2059045, 0.1544619, 0.147289, 
    0.122337, 0.1965521, 0.1473452, 0.1864514, 0.268804, 0.3269864, 
    0.2561044, 0.1919433, 0.1878847, 0.176145, 0.2050935,
  0.2282174, 0.1893594, 0.2599252, 0.345011, 0.2808617, 0.3016484, 0.3595511, 
    0.3254358, 0.2795074, 0.3263747, 0.2123578, 0.1543672, 0.1897014, 
    0.2472795, 0.3152657, 0.2043868, 0.2537548, 0.3408902, 0.269443, 
    0.1977303, 0.2028517, 0.170909, 0.2300183, 0.3043991, 0.2489848, 
    0.3305418, 0.3017626, 0.2987627, 0.2235068,
  0.2494897, 0.2469137, 0.2576125, 0.2667766, 0.269223, 0.3370608, 0.2959158, 
    0.4188668, 0.2928834, 0.2523627, 0.2104652, 0.2608206, 0.2643886, 
    0.2051282, 0.1919718, 0.1494743, 0.29427, 0.3386157, 0.2737174, 0.289049, 
    0.2157629, 0.1847745, 0.1901498, 0.2042071, 0.1997167, 0.347068, 
    0.1184259, 0.2182723, 0.1917094,
  0.1965577, 0.2477432, 0.2116805, 0.2106968, 0.1851083, 0.1795774, 
    0.1940835, 0.2085294, 0.1995699, 0.1911565, 0.2451654, 0.2004384, 
    0.2167422, 0.2656918, 0.335009, 0.3423926, 0.2661839, 0.1570902, 
    0.144303, 0.1382567, 0.192824, 0.2089022, 0.1553212, 0.07133471, 
    0.1048343, 0.08797328, 0.1955092, 0.2296528, 0.243732,
  0.07063024, 0.07186922, 0.0731082, 0.07434718, 0.07558617, 0.07682514, 
    0.07806413, 0.08975758, 0.09452108, 0.09928457, 0.1040481, 0.1088116, 
    0.1135751, 0.1183386, 0.1381873, 0.1387293, 0.1392714, 0.1398135, 
    0.1403556, 0.1408977, 0.1414398, 0.1243464, 0.1178018, 0.1112573, 
    0.1047127, 0.09816812, 0.09162355, 0.08507898, 0.06963906,
  0.1885164, 0.1828577, 0.1708737, 0.1741126, 0.1596946, 0.1842122, 
    0.2159217, 0.1922243, 0.1598626, 0.2245309, 0.1214755, 0.1131081, 
    0.164493, 0.1273623, 0.1103211, 0.2285462, 0.250079, 0.2407761, 0.238851, 
    0.2598571, 0.2301687, 0.2521805, 0.1351557, 0.05784683, 0.08294596, 
    0.09694898, 0.05963591, 0.1126747, 0.148323,
  0.2149846, 0.2475992, 0.1565274, 0.1704955, 0.2308763, 0.3034375, 
    0.2023066, 0.2658588, 0.2414473, 0.2696008, 0.2655419, 0.1837359, 
    0.2202301, 0.2534932, 0.2571821, 0.3192424, 0.1893605, 0.2879192, 
    0.277443, 0.2869586, 0.2953454, 0.337851, 0.3257232, 0.3874508, 
    0.2288913, 0.1765311, 0.1691849, 0.2482999, 0.2694762,
  0.329843, 0.3859303, 0.3682566, 0.409528, 0.4399304, 0.4287531, 0.32862, 
    0.3372033, 0.3516958, 0.328775, 0.3583198, 0.3532516, 0.3170046, 
    0.2773377, 0.2678211, 0.2443536, 0.2836554, 0.2518613, 0.286671, 
    0.2884113, 0.2572013, 0.2554939, 0.2528849, 0.269962, 0.2700689, 
    0.2108892, 0.2388085, 0.3106317, 0.3190642,
  0.2416804, 0.2430525, 0.2471741, 0.2381833, 0.2270044, 0.2372918, 
    0.1828865, 0.1810473, 0.1877583, 0.1727558, 0.2082299, 0.1951734, 
    0.2133803, 0.2249564, 0.2033369, 0.1562759, 0.128724, 0.1340789, 
    0.1664077, 0.1536688, 0.2053761, 0.2374049, 0.2230249, 0.1768523, 
    0.09173495, 0.1010696, 0.1545932, 0.1571117, 0.2094709,
  0.05919874, 0.04136188, 0.03920296, 0.08797455, 0.08282591, 0.054277, 
    0.09417309, 0.1116461, 0.04877861, 0.01587244, 0.02777561, 0.03832315, 
    0.07701707, 0.07753734, 0.08797985, 0.053512, 0.08989856, 0.09828319, 
    0.1391574, 0.1347166, 0.06926529, 0.04804907, 0.03869034, 0.03876002, 
    0.04201166, 0.09221782, 0.1046169, 0.09996897, 0.08822098,
  0.006968145, 0.004785631, 0.1248263, 0.02887273, 0.03423189, 0.04147198, 
    0.03563765, 0.02972708, 0.0001375314, 0.005386075, 0.001007872, 
    0.00180555, 0.07852469, 0.01643198, 0.04452884, 0.03475554, 0.07003062, 
    0.1154154, 0.06042206, 0.05314298, 0.01873565, 0.01182871, 1.481094e-05, 
    0.0003168537, 0.0483219, 0.05528377, 0.130739, 0.03627004, 0.01052792,
  0.001951423, 0.05907486, 0.1423884, 0.05233067, 0.08935922, 0.04853534, 
    0.05079352, 0.005656243, 0.0002772567, 0.03752589, 0.04895011, 
    0.09139189, 0.1225506, 0.02934696, 0.039169, 0.1713684, 0.1032087, 
    0.09981325, 0.03257565, 0.04626945, 0.04614308, 0.005802156, 
    3.120092e-07, -0.000112586, 0.1576528, 0.1228896, 0.05323603, 0.03322708, 
    0.001410144,
  2.428496e-06, 0.008681445, 0.3224296, 0.06278799, 0.05717827, 0.03571487, 
    0.04391437, 0.04835663, 0.01903019, 0.06210612, 0.05039233, 0.02025669, 
    0.05441907, 0.02936507, 0.0641021, 0.0794605, 0.06059295, 0.03710041, 
    0.02398305, 0.007453924, 0.000380908, 1.225857e-05, 1.776244e-05, 
    0.07245123, 0.1754165, 0.09640144, 0.03687892, 0.002006771, 7.873497e-05,
  0.008685841, 0.006769489, 0.0167544, 0.05887974, 0.02786795, 0.07557244, 
    0.1137335, 0.03291043, 0.1219867, 0.2157357, 0.0546035, 0.02865683, 
    0.04453103, 0.06053839, 0.0487553, 0.01397876, 0.01329743, 0.002078852, 
    0.009519882, 0.01273254, 0.007256371, 0.03207168, 0.09953449, 0.05649982, 
    0.1045633, 0.1354365, 0.05042254, 0.02297875, 0.01433045,
  7.550081e-08, 4.726625e-07, -2.3307e-06, 0.08645178, 0.03081727, 0.0494937, 
    0.03050793, 0.05932277, 0.03724574, 0.08896187, 0.1729799, 0.09261766, 
    0.05728026, 0.03835767, 0.03691436, 0.03716252, 0.03494349, 0.01757487, 
    0.0324608, 0.04783607, 0.05665651, 0.03513915, 0.06847731, 0.02538132, 
    0.03838209, 0.002710308, 0.0001703476, -5.655221e-06, 0.01560608,
  2.877232e-06, 3.013313e-07, -3.620297e-07, 0.01366376, 0.0006280976, 
    0.003864592, 0.02218705, 0.04217887, 0.02438035, 0.02485721, 0.08254854, 
    0.06352286, 0.05679915, 0.003897997, 0.01327075, 0.00856911, 0.03347083, 
    0.009929997, 0.003614282, 0.04637265, 0.01132111, 0.1039007, 0.03439164, 
    0.07805455, 0.04427945, 0.04682471, 0.006743725, 0.001475899, 0.01241626,
  0.005720179, 0.003435227, 0.02298038, 0.02220487, 0.07219666, 0.02312771, 
    0.005303039, 0.02118771, 0.148673, 0.1267658, 0.0452971, 0.1233826, 
    0.1135696, 0.1419938, 0.1128555, 0.153835, 0.1020103, 0.09845395, 
    0.06086162, 0.02680184, 0.04094369, 0.06101573, 0.0940998, 0.07600197, 
    0.1026166, 0.1010693, 0.06439992, 0.03230079, 0.02173639,
  0.05394094, 0.07178102, 0.1653197, 0.3799989, 0.145744, 0.06473802, 
    0.2779898, 0.02595611, 0.01086512, 0.02486292, 0.0538976, 0.1354104, 
    0.1630195, 0.1955723, 0.2322428, 0.2244351, 0.2154774, 0.2062458, 
    0.1536988, 0.2033992, 0.1872999, 0.07283787, 0.1419569, 0.143596, 
    0.2273832, 0.1865536, 0.195748, 0.1180244, 0.1005927,
  0.2204274, 0.235578, 0.1975906, 0.2442567, 0.1710346, 0.1899409, 0.1231147, 
    0.1409839, 0.1170813, 0.04007668, 0.04448136, 0.1851748, 0.2252243, 
    0.2873888, 0.3189036, 0.2398929, 0.1527601, 0.1672219, 0.123644, 
    0.208068, 0.137904, 0.1790131, 0.2632122, 0.3036509, 0.2456632, 
    0.2112768, 0.214248, 0.1855659, 0.2128806,
  0.2488018, 0.2017359, 0.2294951, 0.3295673, 0.2712059, 0.3234961, 
    0.3617908, 0.3204455, 0.2810445, 0.3414444, 0.2391143, 0.1401209, 
    0.2094419, 0.2434589, 0.3164209, 0.1919684, 0.2590258, 0.3557929, 
    0.2642585, 0.1809855, 0.1892555, 0.1751065, 0.214496, 0.2862013, 
    0.2297303, 0.3457491, 0.3172941, 0.3031945, 0.2614139,
  0.2560236, 0.2964432, 0.2449785, 0.3313259, 0.2989048, 0.3244812, 
    0.3194277, 0.4316089, 0.2975883, 0.2570834, 0.227001, 0.2811974, 
    0.2728152, 0.2195612, 0.1954731, 0.149552, 0.2727693, 0.3540181, 
    0.2728115, 0.2460313, 0.2528111, 0.1770725, 0.1903208, 0.1638058, 
    0.2055477, 0.4069258, 0.1297678, 0.2295569, 0.2130733,
  0.1958748, 0.2391278, 0.203843, 0.2058152, 0.1834047, 0.1984574, 0.1997195, 
    0.2312422, 0.1895227, 0.1974711, 0.2376776, 0.2054238, 0.2252808, 
    0.2697943, 0.3195605, 0.3392972, 0.2546763, 0.1396419, 0.1532362, 
    0.1683775, 0.2018802, 0.2062348, 0.165015, 0.07832222, 0.1000929, 
    0.1027908, 0.1842084, 0.2215886, 0.2376652,
  0.07756125, 0.07892063, 0.08027999, 0.08163936, 0.08299874, 0.0843581, 
    0.08571748, 0.1025454, 0.1059368, 0.1093282, 0.1127196, 0.116111, 
    0.1195024, 0.1228938, 0.1289995, 0.1288216, 0.1286436, 0.1284657, 
    0.1282877, 0.1281098, 0.1279318, 0.112446, 0.1078732, 0.1033003, 
    0.09872752, 0.09415469, 0.08958185, 0.08500903, 0.07647376,
  0.1969301, 0.1781384, 0.1861036, 0.1729915, 0.1623851, 0.2141434, 
    0.2649475, 0.2659005, 0.1530878, 0.240103, 0.133879, 0.1080882, 
    0.1890809, 0.06756324, 0.07435203, 0.1403405, 0.1789874, 0.1767524, 
    0.2013719, 0.224244, 0.2378453, 0.2365764, 0.1152594, 0.05399625, 
    0.1070088, 0.1735752, 0.1252552, 0.1097862, 0.1779886,
  0.1759762, 0.173325, 0.169129, 0.1688088, 0.210343, 0.3341773, 0.195691, 
    0.2748697, 0.234423, 0.2526891, 0.2584201, 0.1742061, 0.243603, 0.22081, 
    0.2378767, 0.2476008, 0.2162304, 0.2625333, 0.2437242, 0.3077757, 
    0.2132913, 0.2501348, 0.3200125, 0.3719279, 0.1744482, 0.1567709, 
    0.1837687, 0.2685302, 0.2711928,
  0.3276001, 0.39336, 0.3324373, 0.3698798, 0.3698794, 0.3420593, 0.316951, 
    0.3011129, 0.33565, 0.3400896, 0.3320581, 0.3209723, 0.2801814, 
    0.2653364, 0.2370964, 0.2346876, 0.2612958, 0.2323375, 0.26261, 
    0.2835625, 0.2366907, 0.2406314, 0.2534537, 0.2660724, 0.2537794, 
    0.2052877, 0.2365877, 0.2780527, 0.3098216,
  0.2301359, 0.2414265, 0.2381935, 0.2268472, 0.2445364, 0.2373807, 
    0.2002448, 0.1998437, 0.213373, 0.1859866, 0.233915, 0.2218721, 
    0.2375394, 0.2289018, 0.1954295, 0.1591772, 0.1261731, 0.1469136, 
    0.149308, 0.1732519, 0.2095126, 0.2265379, 0.2484361, 0.1772104, 
    0.09093638, 0.1033625, 0.1409028, 0.1456343, 0.2057208,
  0.07361671, 0.0681165, 0.06074379, 0.1054547, 0.1075235, 0.06195016, 
    0.09957723, 0.1014156, 0.0599515, 0.01709549, 0.02633458, 0.04325348, 
    0.08059649, 0.08750718, 0.1057701, 0.06636856, 0.1167983, 0.1045027, 
    0.1342559, 0.1442427, 0.09020742, 0.05547203, 0.06410259, 0.04605159, 
    0.03274381, 0.08810988, 0.1207003, 0.09443696, 0.09655182,
  0.009062937, 0.004681489, 0.1113362, 0.03606282, 0.0320303, 0.04935593, 
    0.04677079, 0.04848509, 0.0008040535, 0.004236262, 0.0001300772, 
    0.0003569853, 0.06511469, 0.01998401, 0.05352326, 0.04761922, 0.07195569, 
    0.1199084, 0.05850522, 0.05708544, 0.03163736, 0.02952407, 0.001883986, 
    8.514319e-05, 0.049448, 0.05375104, 0.123303, 0.04752686, 0.01971301,
  0.001863506, 0.03779427, 0.1603097, 0.05381346, 0.07693158, 0.05097435, 
    0.05866064, 0.01644277, 0.00275113, 0.03855854, 0.03862222, 0.07596371, 
    0.1199132, 0.03324369, 0.03965208, 0.1520783, 0.08958703, 0.0846166, 
    0.02643317, 0.03903693, 0.07779795, 0.04233678, -5.200184e-06, 
    6.203083e-06, 0.1605256, 0.111389, 0.03863549, 0.08030573, 0.01612387,
  0.0004461783, 0.01002292, 0.3060247, 0.05356232, 0.04651822, 0.03143445, 
    0.04412724, 0.04922283, 0.02153497, 0.05698334, 0.05337574, 0.01756812, 
    0.05006547, 0.0266456, 0.05064663, 0.06422494, 0.05301657, 0.03037365, 
    0.02493904, 0.01521294, 0.001422074, 0.0003021313, 8.359603e-05, 
    0.06811947, 0.1447769, 0.08230014, 0.03625051, 0.004614646, 0.002527591,
  0.005308207, 0.007748675, 0.008244097, 0.04237524, 0.03524648, 0.07794083, 
    0.1069303, 0.02638575, 0.1558833, 0.2159968, 0.05289855, 0.02580136, 
    0.0365819, 0.05370637, 0.04462192, 0.01648582, 0.01957414, 0.01131988, 
    0.01211746, 0.01498748, 0.01777758, 0.03075802, 0.07590609, 0.05764236, 
    0.109904, 0.1201074, 0.04423032, 0.02604523, 0.01433276,
  2.532936e-08, 9.198961e-08, 2.031705e-09, 0.03807316, 0.04071039, 
    0.07324136, 0.0404203, 0.05450009, 0.04019376, 0.09746628, 0.1841695, 
    0.08803512, 0.05808036, 0.04750704, 0.0392228, 0.03926384, 0.03445046, 
    0.02054641, 0.03957038, 0.04721562, 0.05441146, 0.03526661, 0.09821592, 
    0.02955574, 0.03293556, 0.006592939, 0.0005315684, 7.325533e-05, 
    0.01270505,
  2.154317e-06, 2.062807e-07, -4.586241e-05, 0.03544738, -1.589988e-07, 
    0.00544245, 0.03588447, 0.04779686, 0.03681761, 0.08198288, 0.08254436, 
    0.06906404, 0.06042349, 0.01220331, 0.03393061, 0.01444975, 0.03724517, 
    0.0211221, 0.006155321, 0.04497414, 0.006040387, 0.1528714, 0.04116936, 
    0.09364422, 0.0451612, 0.06092705, 0.02030906, 0.003947348, 0.006064294,
  0.01113623, 0.005638443, 0.03760892, 0.02584603, 0.0665179, 0.02008023, 
    0.004259293, 0.01654099, 0.1351193, 0.08880401, 0.06604788, 0.1769537, 
    0.1265602, 0.1434868, 0.1202914, 0.1626665, 0.1102398, 0.09561702, 
    0.07648773, 0.02523787, 0.05034374, 0.06188781, 0.09485052, 0.107879, 
    0.1059851, 0.1048588, 0.07080483, 0.03972185, 0.01914925,
  0.05378395, 0.09512732, 0.1587929, 0.4052167, 0.1649314, 0.06274316, 
    0.264716, 0.02268014, 0.00548723, 0.02127486, 0.04890822, 0.1797214, 
    0.1994147, 0.2200531, 0.2470819, 0.2415564, 0.222206, 0.2048174, 
    0.1745085, 0.2151118, 0.180699, 0.08201325, 0.1517096, 0.1541929, 
    0.2533481, 0.1977497, 0.1983074, 0.1241219, 0.1154662,
  0.2134503, 0.2555167, 0.2100517, 0.2137466, 0.1703241, 0.1856823, 
    0.1144872, 0.1448835, 0.1041657, 0.02998942, 0.04207374, 0.1992326, 
    0.2817809, 0.3437023, 0.3449514, 0.2465963, 0.1559856, 0.1878847, 
    0.1302626, 0.2243959, 0.1538925, 0.1897459, 0.2616316, 0.2915274, 
    0.2540711, 0.2354159, 0.2316883, 0.2140693, 0.2183427,
  0.2716778, 0.2039053, 0.2156217, 0.3165648, 0.3126442, 0.3215852, 
    0.3472434, 0.3225046, 0.2896096, 0.3412376, 0.258, 0.1242939, 0.2114947, 
    0.2468403, 0.3285189, 0.161636, 0.2358363, 0.3671395, 0.2730772, 
    0.1562053, 0.1773067, 0.1900369, 0.2429075, 0.2553635, 0.2214137, 
    0.34458, 0.3301613, 0.3176329, 0.2554862,
  0.2840129, 0.3377894, 0.2576062, 0.3505348, 0.2752805, 0.348423, 0.3414563, 
    0.4617503, 0.3135374, 0.2672337, 0.2426768, 0.2786874, 0.2908004, 
    0.23444, 0.2310028, 0.1382296, 0.2788805, 0.3840399, 0.2852387, 
    0.2404897, 0.2642761, 0.1952822, 0.2217564, 0.126279, 0.2160996, 
    0.4675737, 0.1348711, 0.2228189, 0.2215622,
  0.2170984, 0.212305, 0.2390421, 0.2123658, 0.2190626, 0.2347994, 0.2104911, 
    0.219753, 0.1825397, 0.211995, 0.2218154, 0.2267924, 0.2533583, 
    0.2893982, 0.317716, 0.3313791, 0.2585874, 0.1452245, 0.1602286, 
    0.2009668, 0.2140926, 0.2316817, 0.1838389, 0.08212442, 0.09762961, 
    0.1048731, 0.1918048, 0.2473738, 0.2831947,
  0.07177738, 0.07374607, 0.07571475, 0.07768343, 0.07965212, 0.08162081, 
    0.08358949, 0.1028914, 0.1048308, 0.1067702, 0.1087097, 0.1106491, 
    0.1125885, 0.1145279, 0.1307912, 0.1304261, 0.130061, 0.1296958, 
    0.1293307, 0.1289655, 0.1286004, 0.1094469, 0.1059039, 0.1023609, 
    0.09881797, 0.09527501, 0.09173205, 0.08818909, 0.07020244,
  0.1991549, 0.1729981, 0.1823778, 0.1760529, 0.1747032, 0.22306, 0.3012792, 
    0.2727414, 0.1547663, 0.2187124, 0.1704121, 0.1228874, 0.2073361, 
    0.05105985, 0.1140422, 0.1480189, 0.1884384, 0.1632211, 0.2025188, 
    0.2231172, 0.284156, 0.2202855, 0.1270158, 0.06228419, 0.159888, 
    0.1372804, 0.05176094, 0.08790512, 0.1940029,
  0.1855603, 0.1948401, 0.1654953, 0.114062, 0.2069466, 0.3418957, 0.1513609, 
    0.275341, 0.2335432, 0.246666, 0.2606984, 0.1793725, 0.2323539, 
    0.2277541, 0.2608104, 0.2922668, 0.2602293, 0.304203, 0.2730995, 
    0.3182649, 0.2889219, 0.2544797, 0.2792223, 0.3637032, 0.1781292, 
    0.1941399, 0.2435258, 0.3386311, 0.2854862,
  0.3599409, 0.3938628, 0.3667728, 0.3583918, 0.3478388, 0.3751264, 
    0.3538289, 0.3397142, 0.3804079, 0.3697892, 0.3858998, 0.3195828, 
    0.2674225, 0.2906128, 0.2552825, 0.2601035, 0.2769893, 0.2576816, 
    0.2878181, 0.313537, 0.2844521, 0.2892179, 0.2989652, 0.2972019, 
    0.2722467, 0.2159816, 0.2485878, 0.3102385, 0.3419653,
  0.2643935, 0.2631836, 0.2551584, 0.2530677, 0.2756747, 0.2609109, 
    0.2262912, 0.2501, 0.218384, 0.2191827, 0.2599172, 0.2454628, 0.2596008, 
    0.2439299, 0.1888632, 0.1580762, 0.1480566, 0.1837746, 0.168883, 
    0.2242923, 0.2251926, 0.2566988, 0.2786165, 0.1750696, 0.08835417, 
    0.1111853, 0.1505524, 0.1638306, 0.2342403,
  0.1080342, 0.1041758, 0.1102329, 0.1534852, 0.1359596, 0.09232381, 
    0.1318851, 0.1242075, 0.09542558, 0.03161843, 0.04102593, 0.06661321, 
    0.08786858, 0.09114663, 0.1257555, 0.09296314, 0.1365167, 0.124594, 
    0.1567495, 0.1700611, 0.1113667, 0.08385252, 0.1228727, 0.05485884, 
    0.02939179, 0.09289541, 0.1412937, 0.09734602, 0.1090793,
  0.02752213, 0.02835215, 0.1140131, 0.05701641, 0.03489635, 0.06466109, 
    0.06107396, 0.05227632, 0.007805334, 0.002601676, 3.284885e-05, 
    -2.839198e-06, 0.06027784, 0.05117114, 0.06395846, 0.06245505, 
    0.08474663, 0.1365128, 0.05413968, 0.05817804, 0.04830899, 0.05646795, 
    0.02354527, 1.908904e-05, 0.0556559, 0.06400656, 0.1130806, 0.04801208, 
    0.04181071,
  0.01229669, 0.03233982, 0.159945, 0.05577642, 0.06738614, 0.04779532, 
    0.05431397, 0.02634654, 0.007934254, 0.05293768, 0.03282881, 0.06607091, 
    0.1079568, 0.03000507, 0.04175595, 0.1390493, 0.08136576, 0.07079503, 
    0.02380499, 0.02832124, 0.06146685, 0.1151802, 0.001564917, 0.0002463174, 
    0.1703525, 0.1139528, 0.02918475, 0.06831248, 0.06920234,
  0.005243808, 0.007996164, 0.2725869, 0.05012213, 0.03849404, 0.02831959, 
    0.04067513, 0.05048361, 0.02498325, 0.04950141, 0.06562485, 0.0157009, 
    0.0493374, 0.02358226, 0.03886451, 0.04541354, 0.04490409, 0.02678851, 
    0.02530962, 0.03511277, 0.01482524, 0.003942169, 0.0003083406, 
    0.06500177, 0.1149733, 0.06988701, 0.04115722, 0.009993114, 0.01217531,
  0.005464268, 0.009746258, 0.008132596, 0.02868435, 0.03445054, 0.06749163, 
    0.09306173, 0.02195093, 0.16098, 0.2314924, 0.05195874, 0.02181398, 
    0.03013392, 0.04636548, 0.04350552, 0.01949322, 0.02256332, 0.01484835, 
    0.01406326, 0.01994715, 0.02746806, 0.038544, 0.05365063, 0.05693216, 
    0.1047207, 0.1022269, 0.03810386, 0.0236931, 0.01184267,
  9.264275e-09, 2.663665e-08, 4.082895e-08, 0.01429612, 0.07368299, 
    0.08629566, 0.04479733, 0.05081002, 0.05478854, 0.09529205, 0.1856278, 
    0.07822891, 0.05712548, 0.05255651, 0.04389524, 0.03974493, 0.03285017, 
    0.02557956, 0.04525636, 0.04346769, 0.04840962, 0.02866706, 0.1282616, 
    0.03508719, 0.03047909, 0.01440951, 0.004212094, 4.945949e-05, 0.01002206,
  1.036187e-06, 1.646142e-07, 0.0004628999, 0.0424123, -9.884328e-06, 
    0.05969144, 0.04993434, 0.04668783, 0.06816496, 0.1741051, 0.09759824, 
    0.1135539, 0.07543223, 0.037128, 0.06540856, 0.03469129, 0.03838166, 
    0.03132236, 0.02322083, 0.04368296, 0.003690798, 0.1783223, 0.04537463, 
    0.1039635, 0.04284891, 0.05781173, 0.05915419, 0.01247508, 0.0008279458,
  0.002579359, 0.007734504, 0.06399792, 0.02970086, 0.06524523, 0.01393953, 
    0.01319417, 0.01319551, 0.1197988, 0.07273196, 0.184405, 0.2349278, 
    0.1529945, 0.1573074, 0.1514286, 0.1797162, 0.1261333, 0.09909804, 
    0.0999874, 0.03508107, 0.06158227, 0.07969914, 0.08677322, 0.1528895, 
    0.1277968, 0.1114864, 0.07967141, 0.05109973, 0.0162567,
  0.05103441, 0.1000903, 0.1537358, 0.4141365, 0.1575812, 0.06424592, 
    0.2275818, 0.01638625, 0.005383232, 0.02099687, 0.04570806, 0.2738684, 
    0.2642636, 0.2311627, 0.2503522, 0.2645875, 0.2444922, 0.2132986, 
    0.2274397, 0.2467405, 0.1962232, 0.1018657, 0.1830252, 0.1955535, 
    0.291157, 0.2037149, 0.229405, 0.1537485, 0.1349008,
  0.2526704, 0.268826, 0.2260363, 0.2148712, 0.1634592, 0.2131425, 0.127093, 
    0.1542884, 0.09877212, 0.02469247, 0.04835953, 0.2057657, 0.3392794, 
    0.4248243, 0.3826507, 0.3098802, 0.2138635, 0.2397596, 0.180218, 
    0.2244172, 0.1615559, 0.2112516, 0.2818637, 0.2976879, 0.2763766, 
    0.3014501, 0.2725008, 0.2251514, 0.2381303,
  0.2889962, 0.1842097, 0.2372937, 0.3103325, 0.3282414, 0.2995462, 
    0.3976163, 0.349923, 0.297824, 0.3622882, 0.2827623, 0.1102727, 
    0.2069141, 0.2721703, 0.3450542, 0.1562482, 0.2505594, 0.3804567, 
    0.2841651, 0.1486751, 0.1936366, 0.2229703, 0.2329464, 0.2483186, 
    0.2665521, 0.3201719, 0.3202224, 0.34233, 0.2620014,
  0.3770165, 0.330017, 0.299314, 0.3200104, 0.2983944, 0.3820589, 0.3808196, 
    0.4911512, 0.34038, 0.3107595, 0.2473948, 0.2771403, 0.2820841, 
    0.2694632, 0.2579285, 0.145909, 0.3215059, 0.4210272, 0.2958125, 
    0.2276349, 0.2674731, 0.2097237, 0.2264613, 0.1027743, 0.2013452, 
    0.4974819, 0.1432499, 0.2092406, 0.3177264,
  0.2400765, 0.2024216, 0.2690099, 0.2500435, 0.2294389, 0.2576038, 
    0.2270053, 0.2405083, 0.2066694, 0.2205156, 0.225161, 0.2418002, 
    0.2678147, 0.3084102, 0.3273087, 0.3273743, 0.2838347, 0.1573666, 
    0.2028611, 0.2392534, 0.2240318, 0.2443569, 0.1809487, 0.08097078, 
    0.09873452, 0.1167171, 0.2032586, 0.2861124, 0.3668998,
  0.1004651, 0.1026717, 0.1048782, 0.1070848, 0.1092914, 0.1114979, 
    0.1137045, 0.1319584, 0.131978, 0.1319976, 0.1320172, 0.1320369, 
    0.1320565, 0.1320761, 0.123794, 0.1224717, 0.1211495, 0.1198272, 
    0.1185049, 0.1171826, 0.1158603, 0.1028088, 0.1019049, 0.1010009, 
    0.100097, 0.09919313, 0.09828922, 0.09738532, 0.09869987,
  0.1996403, 0.1758333, 0.1904247, 0.1667487, 0.2026823, 0.2430759, 
    0.3138554, 0.2879211, 0.1719327, 0.2279047, 0.1826965, 0.130158, 
    0.2139291, 0.05463694, 0.1189097, 0.1992507, 0.20196, 0.2065703, 
    0.2173043, 0.2056393, 0.2876555, 0.2533562, 0.1756549, 0.1116238, 
    0.1774259, 0.113344, 0.1358432, 0.1419035, 0.2057894,
  0.2314472, 0.2000553, 0.1613334, 0.111806, 0.2028545, 0.3608537, 0.1246676, 
    0.2639224, 0.2497888, 0.2379784, 0.252051, 0.1852799, 0.245398, 0.233892, 
    0.3121507, 0.3328328, 0.3179775, 0.4246018, 0.3178639, 0.3378372, 
    0.3233291, 0.3461571, 0.3348624, 0.3793549, 0.1979026, 0.231034, 
    0.3161912, 0.401437, 0.3463486,
  0.4337018, 0.4052368, 0.3833297, 0.4386269, 0.3918735, 0.4241797, 
    0.3948628, 0.3945121, 0.4170676, 0.404942, 0.4120272, 0.4189023, 
    0.3531669, 0.3586879, 0.3439925, 0.3195873, 0.333437, 0.3178196, 
    0.3514133, 0.3880751, 0.3438093, 0.3480112, 0.3841909, 0.3747407, 
    0.3935019, 0.334868, 0.3019947, 0.3440234, 0.419818,
  0.327311, 0.3047533, 0.3245318, 0.3100753, 0.3206269, 0.3003439, 0.2652289, 
    0.3090374, 0.2338096, 0.2575741, 0.3075522, 0.2990085, 0.3041246, 
    0.2704023, 0.1776328, 0.195727, 0.1673482, 0.2199542, 0.1979001, 
    0.2543781, 0.2786545, 0.2908592, 0.3125479, 0.162414, 0.07659961, 
    0.1156516, 0.192285, 0.2160216, 0.272419,
  0.156739, 0.1487535, 0.2082424, 0.2197855, 0.1891064, 0.1693208, 0.1914054, 
    0.1792902, 0.1213345, 0.07325782, 0.08344789, 0.1050563, 0.09343047, 
    0.1283437, 0.1571067, 0.1107152, 0.1853793, 0.1579251, 0.2080966, 
    0.2099499, 0.1439253, 0.149239, 0.1689314, 0.06973644, 0.03637291, 
    0.1207173, 0.1774375, 0.133474, 0.1441663,
  0.1110721, 0.03308049, 0.1149771, 0.08767679, 0.04255571, 0.09029428, 
    0.08052593, 0.08958185, 0.04336766, 0.002653235, -3.473713e-05, 
    1.724599e-05, 0.04959157, 0.06115761, 0.09174173, 0.095171, 0.1130577, 
    0.1412392, 0.06444011, 0.05509523, 0.04989516, 0.07997011, 0.09419118, 
    -1.759522e-06, 0.07031989, 0.06754411, 0.1135695, 0.05035448, 0.07825287,
  0.09959187, 0.02162617, 0.1382003, 0.05285191, 0.05779812, 0.04709151, 
    0.0501549, 0.05381035, 0.02961555, 0.05637462, 0.03600056, 0.05396771, 
    0.09971188, 0.02958531, 0.04488068, 0.1312134, 0.07734217, 0.06097101, 
    0.02636028, 0.03065137, 0.04435501, 0.1587616, 0.04941503, 0.0003203357, 
    0.1826258, 0.1275736, 0.03158822, 0.06455534, 0.1203822,
  0.01155564, 0.007044189, 0.2340138, 0.05196911, 0.03317957, 0.02869007, 
    0.03802095, 0.05176207, 0.03357369, 0.04564068, 0.0698674, 0.0181426, 
    0.04976706, 0.02447531, 0.03241329, 0.03901483, 0.04291175, 0.02932809, 
    0.02753149, 0.03026662, 0.04345087, 0.03000213, 0.00781719, 0.05997044, 
    0.09230819, 0.06265479, 0.05051921, 0.03047703, 0.0308056,
  0.01956628, 0.02210601, 0.004524016, 0.02052965, 0.03438834, 0.05679921, 
    0.07920136, 0.02336333, 0.1614146, 0.2215357, 0.05031688, 0.02024117, 
    0.0269568, 0.04295023, 0.04207287, 0.02203964, 0.02466078, 0.01097101, 
    0.01669717, 0.02238476, 0.04436092, 0.03463591, 0.03912115, 0.05532191, 
    0.1007729, 0.08512293, 0.03567838, 0.02552984, 0.01580546,
  5.069507e-09, 1.02991e-08, 1.329628e-08, 0.005870801, 0.1313287, 0.1097654, 
    0.03699206, 0.08371939, 0.07814619, 0.09533129, 0.1742087, 0.06981514, 
    0.05159377, 0.05405042, 0.05275682, 0.03951509, 0.03243978, 0.03347987, 
    0.05145106, 0.04035984, 0.04452064, 0.03003637, 0.1368022, 0.04834656, 
    0.03597354, 0.0282557, 0.01131955, -3.666195e-05, 0.007663086,
  4.189981e-07, 7.464039e-08, 0.0005337175, 0.03804546, 5.767886e-07, 
    0.08842903, 0.05005502, 0.08017723, 0.04756146, 0.2119018, 0.1913961, 
    0.1914799, 0.1429465, 0.09205781, 0.1569333, 0.1019502, 0.05227114, 
    0.03960821, 0.04921282, 0.08309115, 0.005374436, 0.2275229, 0.09408981, 
    0.1068835, 0.061196, 0.07482523, 0.1085902, 0.02194129, -2.441665e-05,
  0.003815975, 0.02779422, 0.1132933, 0.04113807, 0.07304354, 0.009859612, 
    0.01204808, 0.009013187, 0.09478872, 0.07504998, 0.332636, 0.1865346, 
    0.1256826, 0.1612821, 0.1434517, 0.1712592, 0.1412436, 0.1727487, 
    0.1125501, 0.08524951, 0.06394763, 0.1057103, 0.07308017, 0.1803523, 
    0.1183744, 0.1473934, 0.09920762, 0.06804402, 0.01645759,
  0.04503657, 0.1007394, 0.170854, 0.4149054, 0.1599987, 0.07622387, 
    0.1951955, 0.01030007, 0.002048314, 0.02110137, 0.05975058, 0.365474, 
    0.3009086, 0.2128668, 0.2219309, 0.2647118, 0.2583112, 0.2315924, 
    0.2597665, 0.2703335, 0.2148291, 0.09414905, 0.2168017, 0.2144901, 
    0.3211913, 0.2344888, 0.2258515, 0.193612, 0.1676942,
  0.2802026, 0.320419, 0.252672, 0.2890696, 0.2134314, 0.2793693, 0.1318641, 
    0.1646207, 0.09099888, 0.02315369, 0.06265467, 0.2299781, 0.3896872, 
    0.3784675, 0.3645972, 0.3446723, 0.2767188, 0.2962195, 0.1920729, 
    0.2422082, 0.1708637, 0.2424976, 0.307668, 0.3024389, 0.3198365, 
    0.3447728, 0.2892312, 0.235981, 0.265842,
  0.3394893, 0.1821341, 0.2408461, 0.3108334, 0.3376181, 0.3181736, 0.445005, 
    0.3892537, 0.3325853, 0.3960759, 0.2957978, 0.1127927, 0.2053609, 
    0.3279609, 0.4406741, 0.1745656, 0.3108756, 0.3981749, 0.2879035, 
    0.1572812, 0.2150514, 0.2259097, 0.2245648, 0.2510787, 0.3738441, 
    0.2988245, 0.3226571, 0.3179141, 0.2882458,
  0.3703192, 0.3048421, 0.3157767, 0.3334541, 0.3309593, 0.4087595, 
    0.3981647, 0.5200198, 0.3734217, 0.3543942, 0.2671398, 0.2781627, 
    0.2919785, 0.2861205, 0.2893866, 0.1769155, 0.3739291, 0.4500185, 
    0.2965789, 0.2463774, 0.2709173, 0.2219616, 0.2253855, 0.09854059, 
    0.1886863, 0.5050979, 0.1475908, 0.1922425, 0.3989843,
  0.2440605, 0.2220331, 0.2969181, 0.2593498, 0.2293969, 0.2792766, 0.264048, 
    0.2579025, 0.2441199, 0.2585242, 0.2609379, 0.2582428, 0.2805758, 
    0.3250264, 0.353653, 0.3513996, 0.2878314, 0.1503806, 0.1844678, 
    0.2744858, 0.2331191, 0.2544084, 0.1861654, 0.08076268, 0.0982402, 
    0.1141233, 0.2212199, 0.3180485, 0.3673283,
  0.1566395, 0.1573331, 0.1580267, 0.1587202, 0.1594138, 0.1601074, 
    0.1608009, 0.1706757, 0.170166, 0.1696564, 0.1691468, 0.1686371, 
    0.1681275, 0.1676178, 0.1459947, 0.1441618, 0.1423288, 0.1404958, 
    0.1386628, 0.1368298, 0.1349969, 0.1121781, 0.1138272, 0.1154763, 
    0.1171253, 0.1187744, 0.1204234, 0.1220725, 0.1560847,
  0.2438885, 0.1787127, 0.2108183, 0.1732268, 0.2272893, 0.2607077, 
    0.3144073, 0.2772256, 0.1620593, 0.2498132, 0.2184614, 0.1723068, 
    0.2481121, 0.04797612, 0.1449985, 0.1750598, 0.1965169, 0.204966, 
    0.2126811, 0.2332719, 0.3321746, 0.2727605, 0.2246664, 0.1481977, 
    0.1702632, 0.153987, 0.1110515, 0.2017663, 0.2503371,
  0.2680483, 0.1927864, 0.1680439, 0.111678, 0.2197834, 0.4117394, 0.1003503, 
    0.2509379, 0.2702884, 0.2645592, 0.2592883, 0.2520164, 0.2440203, 
    0.2541229, 0.3540066, 0.4286997, 0.4339809, 0.5018978, 0.3440653, 
    0.4120452, 0.3996732, 0.4225238, 0.4014142, 0.3870392, 0.2263055, 
    0.370573, 0.5026637, 0.4061979, 0.4218117,
  0.4630283, 0.4301504, 0.4141735, 0.5100102, 0.454957, 0.4801038, 0.436365, 
    0.4790096, 0.4904942, 0.428899, 0.4737488, 0.4710087, 0.4516402, 
    0.4599753, 0.3924145, 0.3910595, 0.3970557, 0.3837312, 0.453159, 
    0.4080013, 0.4054448, 0.3994575, 0.4113336, 0.4116966, 0.4417846, 
    0.4186906, 0.3852264, 0.4355152, 0.4636422,
  0.3784615, 0.3799152, 0.4353657, 0.3617443, 0.3544714, 0.3292845, 
    0.3080423, 0.3409056, 0.2813881, 0.3259102, 0.3639681, 0.3563793, 
    0.2994419, 0.2515345, 0.156025, 0.2088325, 0.1725554, 0.2333361, 
    0.2683704, 0.2607414, 0.2894211, 0.3139735, 0.343435, 0.155362, 
    0.06492797, 0.1483287, 0.2590926, 0.2964505, 0.3041558,
  0.1983176, 0.2125988, 0.2193201, 0.2279017, 0.2291522, 0.2469288, 
    0.2315758, 0.2324258, 0.2016309, 0.1521738, 0.2074326, 0.1336438, 
    0.08926547, 0.1670656, 0.189411, 0.1916464, 0.2981403, 0.2504219, 
    0.2539986, 0.2567993, 0.1447949, 0.2154545, 0.2177263, 0.08612543, 
    0.05433446, 0.1415471, 0.2442462, 0.2065925, 0.2265716,
  0.1432197, 0.04315274, 0.1006749, 0.1346003, 0.05675261, 0.08640645, 
    0.1505772, 0.1890068, 0.2120956, 0.007762956, 0.0004954685, 9.095662e-06, 
    0.03763352, 0.06906883, 0.1374171, 0.1298566, 0.2039855, 0.1696494, 
    0.1118311, 0.08055007, 0.05562823, 0.1094994, 0.2241403, -1.551987e-06, 
    0.06422567, 0.09659802, 0.1209114, 0.0522344, 0.1211668,
  0.2365946, 0.02118609, 0.1119277, 0.0611729, 0.06104632, 0.05518041, 
    0.0607205, 0.09221381, 0.0971193, 0.06709974, 0.03226288, 0.04014831, 
    0.09247859, 0.04419443, 0.07192025, 0.1203822, 0.09097879, 0.06309342, 
    0.03596007, 0.04210299, 0.04789975, 0.1843203, 0.3514513, 0.0008980334, 
    0.1565434, 0.1263198, 0.04457146, 0.0573357, 0.1301481,
  0.05073747, 0.01167894, 0.1956373, 0.05379686, 0.0337343, 0.03253026, 
    0.04030035, 0.05350109, 0.04270298, 0.04706538, 0.0609058, 0.02707743, 
    0.04696836, 0.03461954, 0.04447062, 0.042781, 0.06659238, 0.05153442, 
    0.05538862, 0.05317689, 0.06835535, 0.07643957, 0.04608938, 0.04850512, 
    0.07841086, 0.04347198, 0.0872467, 0.06381261, 0.07976979,
  0.01304233, 0.017083, 0.001567481, 0.01300887, 0.04537904, 0.06651258, 
    0.0837653, 0.03156782, 0.1537119, 0.1979657, 0.04919566, 0.0238379, 
    0.029797, 0.04590497, 0.05422922, 0.04345524, 0.02926396, 0.01472992, 
    0.02155234, 0.02676026, 0.04585477, 0.04822522, 0.03847935, 0.04301926, 
    0.0888631, 0.07051214, 0.03934302, 0.03280829, 0.02000054,
  3.548333e-09, 5.138406e-09, 3.88818e-09, 0.0001849835, 0.1564875, 
    0.1329755, 0.01524338, 0.1377285, 0.108792, 0.07759997, 0.1694398, 
    0.07127045, 0.04948694, 0.05617285, 0.06169382, 0.0743288, 0.05765457, 
    0.04460396, 0.05765268, 0.04469329, 0.04976716, 0.04559736, 0.1734994, 
    0.05513176, 0.05847016, 0.08180889, 0.2022588, 0.009449132, 0.008032215,
  1.715289e-07, -2.787863e-08, 0.0001460534, 0.01949304, -5.900646e-08, 
    0.054109, 0.03491741, 0.06895985, 0.0374335, 0.308756, 0.2001259, 
    0.2461997, 0.1794631, 0.1478033, 0.1354423, 0.1316537, 0.1065224, 
    0.05115189, 0.1095669, 0.174702, 0.01345942, 0.2698481, 0.1367816, 
    0.1100598, 0.09862965, 0.08518668, 0.1484441, 0.01685217, -6.594123e-06,
  0.004202363, 0.06220856, 0.1220331, 0.06360418, 0.0807783, 0.00773428, 
    0.005007822, 0.005655666, 0.07207458, 0.07375321, 0.2701255, 0.1023324, 
    0.08683077, 0.1101118, 0.1048644, 0.1521856, 0.1314666, 0.1711844, 
    0.09726261, 0.09361695, 0.0739302, 0.1484428, 0.1081218, 0.1539405, 
    0.09947546, 0.1386396, 0.1452122, 0.09464188, 0.01614606,
  0.0403964, 0.1238498, 0.1798082, 0.4153139, 0.1489247, 0.06809916, 
    0.1689497, 0.007164896, 0.0008332973, 0.02004977, 0.07328379, 0.2892644, 
    0.2134376, 0.1539741, 0.1972617, 0.2514833, 0.2791519, 0.277357, 
    0.2375869, 0.2918316, 0.2262952, 0.1066738, 0.2502188, 0.2201706, 
    0.3123201, 0.2162575, 0.1993795, 0.2185521, 0.190588,
  0.3182553, 0.3553693, 0.2847632, 0.3078063, 0.273718, 0.3166443, 0.1633989, 
    0.1741175, 0.08703892, 0.02721077, 0.07017485, 0.2639569, 0.377449, 
    0.2868895, 0.3262295, 0.3326616, 0.3208802, 0.2871472, 0.1852327, 
    0.2650878, 0.1993838, 0.2774741, 0.3411638, 0.3264908, 0.3515668, 
    0.318049, 0.2338735, 0.2265158, 0.3074211,
  0.291416, 0.155328, 0.2826667, 0.3770149, 0.3889391, 0.3345815, 0.4598645, 
    0.41506, 0.3529751, 0.4388548, 0.3675779, 0.1268159, 0.2009772, 
    0.3206494, 0.5644627, 0.2510937, 0.3717691, 0.413619, 0.3127052, 
    0.1756986, 0.2329371, 0.2233764, 0.2142618, 0.2453339, 0.5501697, 
    0.2196694, 0.2694122, 0.2611139, 0.2365803,
  0.2870576, 0.1979858, 0.2791478, 0.2990038, 0.373341, 0.4279606, 0.4177774, 
    0.5651989, 0.3893551, 0.4072464, 0.3042587, 0.2746203, 0.3251367, 
    0.3246972, 0.3306153, 0.1927602, 0.3994981, 0.481932, 0.3154012, 
    0.3112109, 0.2755656, 0.2308284, 0.2234824, 0.09734072, 0.1655345, 
    0.5171972, 0.14961, 0.1579475, 0.4412608,
  0.224504, 0.2168309, 0.2862285, 0.2509914, 0.2364857, 0.3080851, 0.3508409, 
    0.3391095, 0.2969672, 0.311076, 0.2887279, 0.2781694, 0.3002055, 
    0.3736871, 0.3583533, 0.3731737, 0.2765608, 0.1528046, 0.2096442, 
    0.2866296, 0.2641073, 0.2512986, 0.1919353, 0.08496875, 0.1007585, 
    0.1267551, 0.235909, 0.3293248, 0.3799539,
  0.1817484, 0.1840956, 0.1864428, 0.1887901, 0.1911373, 0.1934845, 
    0.1958318, 0.2095396, 0.2072039, 0.2048682, 0.2025324, 0.2001968, 
    0.1978611, 0.1955253, 0.1829255, 0.1814949, 0.1800642, 0.1786336, 
    0.1772029, 0.1757723, 0.1743417, 0.1568877, 0.1583068, 0.1597259, 
    0.161145, 0.1625641, 0.1639832, 0.1654023, 0.1798706,
  0.3031531, 0.2240513, 0.2549827, 0.194872, 0.2517972, 0.2808021, 0.3257743, 
    0.2702516, 0.182025, 0.3132783, 0.2893526, 0.255739, 0.2869729, 
    0.03438993, 0.1588206, 0.1894409, 0.209118, 0.2565867, 0.2137727, 
    0.2348837, 0.3700337, 0.3437512, 0.2412119, 0.1676399, 0.1152035, 
    0.2959384, 0.09474089, 0.1466069, 0.2415916,
  0.2631764, 0.259062, 0.2043389, 0.1313171, 0.1964954, 0.4499576, 
    0.09539254, 0.2431849, 0.276797, 0.291097, 0.2735163, 0.3393711, 
    0.2118316, 0.3092141, 0.478425, 0.5713874, 0.5149198, 0.5673895, 
    0.3918922, 0.403377, 0.4407787, 0.4423532, 0.4233812, 0.4174761, 
    0.2183923, 0.4489912, 0.4916124, 0.4177064, 0.37614,
  0.523725, 0.4636297, 0.4479968, 0.5160466, 0.5324846, 0.5201598, 0.4634234, 
    0.4956807, 0.5168597, 0.4647013, 0.4783164, 0.4823202, 0.4945955, 
    0.4671479, 0.3957436, 0.4369711, 0.474703, 0.4847535, 0.5120771, 0.42766, 
    0.3977026, 0.3935178, 0.3981849, 0.4200343, 0.4291924, 0.4698754, 
    0.4942711, 0.5249581, 0.5428705,
  0.3996886, 0.4261588, 0.4773311, 0.3492683, 0.4018682, 0.3875193, 
    0.3439168, 0.3575166, 0.3307911, 0.3503316, 0.3627879, 0.3353739, 
    0.2830169, 0.2562194, 0.1585219, 0.2289117, 0.2495465, 0.2809635, 
    0.3378187, 0.3065062, 0.3311161, 0.3609961, 0.3440224, 0.1549186, 
    0.08738789, 0.1584689, 0.3210941, 0.3492914, 0.3261421,
  0.2630006, 0.2630028, 0.1585208, 0.2345527, 0.2260404, 0.2465748, 
    0.2393618, 0.3088939, 0.3275971, 0.2983638, 0.3210226, 0.1204444, 
    0.0911755, 0.1786005, 0.1992568, 0.21701, 0.3006757, 0.3218557, 
    0.2920588, 0.3018102, 0.2804728, 0.2786484, 0.2220929, 0.1061831, 
    0.0510264, 0.167371, 0.2561396, 0.2823249, 0.2556739,
  0.1380108, 0.1243589, 0.07607315, 0.1282459, 0.06206869, 0.1069857, 
    0.1507266, 0.207869, 0.2758573, 0.01356626, 0.0002028604, 2.659147e-06, 
    0.02787772, 0.121907, 0.1539024, 0.1036603, 0.2388192, 0.220945, 
    0.1477334, 0.1121645, 0.1013103, 0.121805, 0.2861113, 0.004370279, 
    0.06500877, 0.07907779, 0.1244838, 0.1009152, 0.1415669,
  0.3384438, 0.02952924, 0.0902175, 0.07733551, 0.06035808, 0.06623837, 
    0.0663229, 0.1127285, 0.3460321, 0.08600266, 0.03083816, 0.02980522, 
    0.0970494, 0.06827872, 0.06581405, 0.1109487, 0.1023282, 0.06458177, 
    0.04519114, 0.03847262, 0.04038201, 0.1148769, 0.5720022, 0.006847052, 
    0.1265253, 0.1067754, 0.072526, 0.03762973, 0.08705854,
  0.1704841, 0.04098625, 0.1521934, 0.05670134, 0.04118683, 0.05806604, 
    0.08150353, 0.08729151, 0.1008169, 0.06368755, 0.04211966, 0.06936442, 
    0.05006707, 0.1080508, 0.07508858, 0.07155873, 0.05915218, 0.0797144, 
    0.04854137, 0.0761383, 0.1381687, 0.2384286, 0.184927, 0.03208823, 
    0.06079487, 0.02931553, 0.08262615, 0.1456822, 0.1709472,
  0.02253099, 0.01084301, 0.0006973983, 0.009265831, 0.07548781, 0.1363256, 
    0.09931386, 0.05698504, 0.1534138, 0.1704421, 0.06315994, 0.08160254, 
    0.04726559, 0.06897796, 0.0773925, 0.07005168, 0.04418239, 0.03151693, 
    0.036172, 0.05793954, 0.08269713, 0.07623975, 0.05306591, 0.02228641, 
    0.05499095, 0.06970698, 0.05213879, 0.06953676, 0.03863704,
  3.024129e-09, 3.025679e-09, 1.099389e-09, -0.003579624, 0.1793811, 
    0.1202196, 0.005004856, 0.1184741, 0.07993229, 0.08168426, 0.1498463, 
    0.08080791, 0.05344959, 0.05108992, 0.06386948, 0.08757286, 0.07807549, 
    0.0729741, 0.08186557, 0.05464996, 0.06496198, 0.06333031, 0.2594847, 
    0.06952775, 0.04006829, 0.05367796, 0.1229645, 0.02128251, 0.007470491,
  6.644805e-08, -4.920481e-06, 0.0001620449, 0.01224561, 7.240423e-09, 
    0.0118832, 0.02179667, 0.04352682, 0.0222852, 0.3125673, 0.1065297, 
    0.1560527, 0.1279852, 0.1147799, 0.08602905, 0.08249015, 0.1407883, 
    0.06157137, 0.1121256, 0.2640961, 0.01559205, 0.2836293, 0.1261469, 
    0.06946129, 0.06861609, 0.08101142, 0.0897103, 0.01131351, -2.617627e-07,
  0.0007692945, 0.05772534, 0.07441655, 0.04254595, 0.08933122, 0.004976418, 
    0.006967309, 0.004383754, 0.0516765, 0.06870983, 0.1693506, 0.06086271, 
    0.05549517, 0.08381993, 0.07681629, 0.1463479, 0.1390195, 0.132359, 
    0.1657503, 0.1040746, 0.08866816, 0.1627335, 0.1253038, 0.1163389, 
    0.08340587, 0.1096255, 0.1478989, 0.1392351, 0.01756159,
  0.03966093, 0.09716365, 0.1437639, 0.4191813, 0.1074021, 0.09284136, 
    0.1517383, 0.006693783, 0.0002245351, 0.01492667, 0.08103488, 0.1275349, 
    0.1342422, 0.1207775, 0.1580558, 0.1982593, 0.236347, 0.2521041, 
    0.2224802, 0.3150474, 0.2240921, 0.1101627, 0.2808369, 0.2249882, 
    0.2355323, 0.1983336, 0.1833108, 0.1944856, 0.2236944,
  0.3397749, 0.3516663, 0.2834615, 0.3125835, 0.300476, 0.3129572, 0.1814395, 
    0.1837116, 0.08378994, 0.04191935, 0.08461726, 0.2747037, 0.2804201, 
    0.202163, 0.2953233, 0.345052, 0.3394594, 0.2864028, 0.201205, 0.2899839, 
    0.2117545, 0.296709, 0.3559181, 0.3875098, 0.4067697, 0.2533212, 
    0.2247539, 0.2145667, 0.2900448,
  0.2266658, 0.1552894, 0.3161725, 0.4322407, 0.4366984, 0.3883106, 
    0.5446943, 0.4941452, 0.416977, 0.4733005, 0.4460721, 0.147849, 
    0.2036739, 0.2663231, 0.5811508, 0.3318493, 0.4058484, 0.4405725, 
    0.3499158, 0.1973178, 0.2820182, 0.2701338, 0.2179583, 0.2333852, 
    0.6459177, 0.1569112, 0.2166514, 0.2088504, 0.2067883,
  0.185441, 0.1335954, 0.2234133, 0.2555335, 0.4157337, 0.3873104, 0.4541551, 
    0.6184369, 0.3792124, 0.4597141, 0.3511838, 0.2826437, 0.3631962, 
    0.3427902, 0.38107, 0.2131548, 0.420756, 0.4988353, 0.3282773, 0.3862593, 
    0.286638, 0.2368796, 0.2368637, 0.1033537, 0.1441038, 0.5025944, 
    0.1555129, 0.1349116, 0.3140671,
  0.2062432, 0.2436966, 0.3150989, 0.2927735, 0.2802392, 0.3620168, 
    0.4121611, 0.3945981, 0.3386852, 0.3348692, 0.318552, 0.3198241, 
    0.3384499, 0.4349321, 0.3748463, 0.4000996, 0.2977254, 0.1915494, 
    0.2574871, 0.3477217, 0.2987399, 0.2679376, 0.1844105, 0.09186491, 
    0.1052828, 0.1367089, 0.2414654, 0.3373206, 0.4427853,
  0.1974759, 0.2031698, 0.2088636, 0.2145575, 0.2202514, 0.2259453, 
    0.2316392, 0.2502146, 0.2463658, 0.2425171, 0.2386684, 0.2348197, 
    0.2309709, 0.2271222, 0.219476, 0.2186177, 0.2177594, 0.2169011, 
    0.2160428, 0.2151844, 0.2143261, 0.1926672, 0.1916804, 0.1906935, 
    0.1897067, 0.1887199, 0.187733, 0.1867462, 0.1929208,
  0.2958975, 0.2346792, 0.2698095, 0.249582, 0.2856941, 0.253442, 0.2831317, 
    0.2507038, 0.2183918, 0.3399493, 0.3187335, 0.2472755, 0.285133, 
    0.03905363, 0.1607305, 0.203906, 0.1824185, 0.2544671, 0.2189671, 
    0.1415332, 0.3012302, 0.3507779, 0.2132575, 0.1292191, 0.1040593, 
    0.2279998, 0.179082, 0.1160706, 0.20296,
  0.2227649, 0.2167116, 0.2380435, 0.1137411, 0.12494, 0.3908572, 0.08934059, 
    0.1906395, 0.2167857, 0.2207359, 0.2470312, 0.3031427, 0.1531676, 
    0.3236152, 0.5672042, 0.556968, 0.4856485, 0.5455487, 0.4188926, 
    0.4885502, 0.4721363, 0.4957627, 0.5152053, 0.4447546, 0.2464606, 
    0.426324, 0.3851303, 0.3260307, 0.3075607,
  0.5405105, 0.4664601, 0.4112562, 0.4763838, 0.5501149, 0.5372881, 0.506723, 
    0.4625372, 0.5094568, 0.4736611, 0.4638487, 0.472225, 0.4702039, 
    0.4231413, 0.3739707, 0.4480855, 0.537763, 0.5440236, 0.5187572, 
    0.4192733, 0.3639354, 0.3607008, 0.3580778, 0.3876183, 0.4279405, 
    0.4316002, 0.5106409, 0.5260665, 0.4964044,
  0.4097773, 0.4118659, 0.4341848, 0.3413451, 0.4166834, 0.3886577, 
    0.3486239, 0.3814679, 0.4008167, 0.3670536, 0.3190672, 0.2529321, 
    0.2410259, 0.2317978, 0.1697605, 0.23528, 0.3124652, 0.3747494, 
    0.3716341, 0.3525217, 0.3504871, 0.3426467, 0.314407, 0.1506485, 
    0.06159478, 0.1747791, 0.3499405, 0.3787965, 0.3724492,
  0.2415744, 0.2090723, 0.106488, 0.1801994, 0.1960372, 0.2349847, 0.2331353, 
    0.3050598, 0.3200399, 0.3017476, 0.2244006, 0.08066801, 0.0715455, 
    0.1385411, 0.2080723, 0.1986998, 0.2064231, 0.2477071, 0.3100812, 
    0.3224449, 0.3017889, 0.2544579, 0.1846469, 0.1298975, 0.0400727, 
    0.194488, 0.2538331, 0.3125426, 0.2236924,
  0.1115937, 0.1465504, 0.06462997, 0.08807321, 0.07495826, 0.06150344, 
    0.06867604, 0.09619851, 0.2076359, 0.01372384, 8.230587e-05, 
    3.005828e-07, 0.02565392, 0.09334894, 0.1092084, 0.06308107, 0.1786704, 
    0.2268798, 0.1397994, 0.06813951, 0.08517981, 0.05830423, 0.1289117, 
    0.02402809, 0.05766118, 0.07121491, 0.1201692, 0.05096367, 0.06915367,
  0.1568614, 0.05384595, 0.0640647, 0.08644035, 0.02564656, 0.03405321, 
    0.03770792, 0.04408605, 0.2320221, 0.1301784, 0.02871123, 0.02095491, 
    0.07104709, 0.03664106, 0.05803587, 0.07959746, 0.06987671, 0.04798351, 
    0.01406679, 0.007269261, 0.01441085, 0.03030782, 0.2798612, 0.2014921, 
    0.1103804, 0.08910547, 0.01740199, 0.007124186, 0.03167034,
  0.3457349, 0.1674593, 0.1228815, 0.06291138, 0.04416688, 0.07927693, 
    0.046092, 0.04577316, 0.0478005, 0.03996494, 0.02652841, 0.03592505, 
    0.03876076, 0.02482904, 0.02509867, 0.02041359, 0.02488091, 0.01792222, 
    0.01036436, 0.017429, 0.03815739, 0.1264321, 0.3306325, 0.0190955, 
    0.04462657, 0.01893912, 0.01840623, 0.04884355, 0.1638084,
  0.02290493, 0.006805738, 0.0003163048, 0.005571354, 0.04915657, 0.09516388, 
    0.07658017, 0.0565102, 0.09637292, 0.1239135, 0.07486778, 0.1111019, 
    0.04339323, 0.03797794, 0.03860947, 0.0407262, 0.03559536, 0.01900459, 
    0.02105542, 0.05302645, 0.1330434, 0.1424394, 0.1105769, 0.01058447, 
    0.02871785, 0.06249637, 0.02399226, 0.03962861, 0.07033528,
  2.749898e-09, 2.358293e-09, 4.784164e-10, -0.00481047, 0.1320463, 
    0.04093023, -0.003243398, 0.05847986, 0.02021855, 0.04397345, 0.1183264, 
    0.05975154, 0.03163739, 0.02119743, 0.02090347, 0.03428464, 0.04361939, 
    0.03390836, 0.06129526, 0.06355764, 0.04570193, 0.03308671, 0.3731316, 
    0.1190187, 0.006978923, 0.01805837, 0.03622718, 0.004962949, 0.006681667,
  2.07036e-08, -1.328765e-05, 0.002713312, 0.002328164, 4.394796e-10, 
    0.003684379, 0.01382634, 0.02187087, 0.01548815, 0.2631747, 0.05966505, 
    0.0755367, 0.068626, 0.05990863, 0.05539062, 0.02977521, 0.06092761, 
    0.0415202, 0.07642774, 0.1470996, 0.0283048, 0.2588981, 0.03261498, 
    0.03097894, 0.03807444, 0.0283371, 0.02724304, 0.00234405, 5.935395e-08,
  0.0008598529, 0.04505378, 0.03253905, 0.02940204, 0.08924252, 0.002376095, 
    0.003702416, 0.005409147, 0.03518409, 0.09089798, 0.1086654, 0.0436565, 
    0.03792901, 0.07239078, 0.07109693, 0.1290109, 0.1280912, 0.09953254, 
    0.1359124, 0.08838412, 0.09423632, 0.1740582, 0.1096588, 0.1080128, 
    0.07068904, 0.09544824, 0.09788388, 0.1073854, 0.02174266,
  0.03988228, 0.0532709, 0.1027172, 0.4124056, 0.06230973, 0.08819485, 
    0.1330344, 0.008428062, 0.0001441427, 0.01347445, 0.08560389, 0.05950813, 
    0.09029794, 0.09889045, 0.1203219, 0.1665373, 0.1970447, 0.2139523, 
    0.1923419, 0.3282954, 0.203994, 0.09737319, 0.3010856, 0.1890409, 
    0.1667272, 0.1696595, 0.1921739, 0.2240147, 0.2523656,
  0.319459, 0.3546227, 0.2782909, 0.3739219, 0.3370652, 0.3427917, 0.1708146, 
    0.1862166, 0.07898092, 0.05421851, 0.08407529, 0.2822102, 0.200162, 
    0.156243, 0.269319, 0.3321723, 0.336493, 0.294414, 0.2182919, 0.3142689, 
    0.2340529, 0.295823, 0.3531464, 0.4380288, 0.4207036, 0.2043035, 
    0.2060124, 0.192871, 0.2427127,
  0.1842813, 0.174251, 0.3588397, 0.4980555, 0.5078447, 0.3899218, 0.6344795, 
    0.527131, 0.4315469, 0.5189819, 0.4952983, 0.1861686, 0.2055281, 
    0.2290881, 0.4874811, 0.3075341, 0.4230194, 0.4273835, 0.3727679, 
    0.2144231, 0.3521186, 0.2941741, 0.2384828, 0.2419778, 0.5812473, 
    0.1126493, 0.1868214, 0.1654862, 0.1771224,
  0.1158523, 0.09230827, 0.2075138, 0.2133489, 0.4848628, 0.4400475, 
    0.5303617, 0.653226, 0.355401, 0.4714533, 0.4139961, 0.3031611, 
    0.4195805, 0.3802383, 0.4155062, 0.25274, 0.4654814, 0.5039691, 
    0.3488045, 0.432285, 0.3025319, 0.2502083, 0.2785353, 0.1126429, 
    0.1224975, 0.4956228, 0.1667765, 0.115549, 0.2199777,
  0.2445391, 0.2984149, 0.3792489, 0.3294459, 0.3054595, 0.4010175, 
    0.4622118, 0.4497333, 0.3825229, 0.3958564, 0.3802468, 0.3684774, 
    0.3874872, 0.4585047, 0.4153026, 0.4302416, 0.3160658, 0.2403393, 
    0.2987241, 0.3900389, 0.3444351, 0.276312, 0.1832049, 0.1140794, 
    0.1247655, 0.1432214, 0.2288782, 0.3362927, 0.5326229,
  0.2514531, 0.2578727, 0.2642923, 0.270712, 0.2771316, 0.2835512, 0.2899708, 
    0.2740163, 0.2699565, 0.2658967, 0.2618369, 0.2577772, 0.2537174, 
    0.2496576, 0.3011893, 0.3004899, 0.2997904, 0.299091, 0.2983916, 
    0.2976921, 0.2969927, 0.2594882, 0.2578278, 0.2561674, 0.254507, 
    0.2528466, 0.2511862, 0.2495258, 0.2463174,
  0.2497503, 0.2561477, 0.2512917, 0.2356944, 0.2412724, 0.1901587, 
    0.2359693, 0.2300338, 0.2057028, 0.3171934, 0.2698497, 0.1775041, 
    0.2285921, 0.0297199, 0.1582593, 0.2367424, 0.1507906, 0.2531572, 
    0.1795683, 0.09096424, 0.215848, 0.2620587, 0.1978411, 0.08250866, 
    0.1674351, 0.1688307, 0.1818829, 0.06629787, 0.1684542,
  0.198997, 0.1506669, 0.2064878, 0.1105066, 0.07197915, 0.3073944, 
    0.08615547, 0.1404251, 0.1515773, 0.1648934, 0.1775288, 0.2189288, 
    0.09957846, 0.2975578, 0.4907838, 0.4765736, 0.4495186, 0.4660092, 
    0.4125801, 0.5227186, 0.5167333, 0.5062626, 0.5698695, 0.4634796, 
    0.2894638, 0.3800998, 0.3055124, 0.2572382, 0.2602256,
  0.4515688, 0.4668985, 0.3763812, 0.4172847, 0.5171174, 0.5274486, 
    0.4969198, 0.4195599, 0.482307, 0.4431689, 0.427187, 0.4505436, 
    0.4588588, 0.4009243, 0.3760499, 0.4255491, 0.5318745, 0.5089978, 
    0.4656305, 0.3823336, 0.3048357, 0.3240753, 0.3225131, 0.3550442, 
    0.3786192, 0.4168578, 0.4836294, 0.4780261, 0.4391392,
  0.4140542, 0.3933963, 0.4010388, 0.3380591, 0.406399, 0.3622546, 0.3393273, 
    0.3374321, 0.3680654, 0.3542309, 0.2690199, 0.196547, 0.2096628, 
    0.2361408, 0.1631968, 0.2792945, 0.3330613, 0.3720509, 0.3532666, 
    0.3642197, 0.3339871, 0.3131737, 0.2872101, 0.1284512, 0.06190272, 
    0.2249547, 0.3944865, 0.4067, 0.3787016,
  0.213233, 0.151276, 0.07836363, 0.1502918, 0.1832747, 0.1864882, 0.2055077, 
    0.2406902, 0.2314779, 0.1671969, 0.1098898, 0.04407894, 0.06203098, 
    0.1494307, 0.2046034, 0.1232307, 0.1429564, 0.1761645, 0.2983312, 
    0.3331168, 0.2690574, 0.184553, 0.1312951, 0.13674, 0.0337982, 0.1794519, 
    0.2771415, 0.3222911, 0.2403956,
  0.04564805, 0.0713672, 0.05228656, 0.05664391, 0.05130758, 0.03914439, 
    0.03376625, 0.04700059, 0.09020705, 0.02004373, -1.217049e-05, 
    -2.786455e-07, 0.02266267, 0.04220412, 0.06849548, 0.03330744, 0.1484568, 
    0.2407407, 0.09400731, 0.02911331, 0.02562581, 0.01672693, 0.04513532, 
    0.05106345, 0.04759875, 0.05199372, 0.07552018, 0.01325337, 0.01973797,
  0.0451817, 0.09139181, 0.05021014, 0.02213482, 0.003678056, 0.01898871, 
    0.02928362, 0.007897422, 0.08484225, 0.1193478, 0.02323133, 0.01591699, 
    0.03594734, 0.009535091, 0.01566431, 0.051392, 0.03820087, 0.02387288, 
    0.001044779, 0.000429049, 0.001189037, 0.005729982, 0.09080987, 
    0.1618166, 0.09057058, 0.08092673, 0.003858366, 0.0003090388, 0.00516483,
  0.1141354, 0.07665696, 0.1058196, 0.05846415, 0.01407639, 0.0132921, 
    0.01396426, 0.01532749, 0.01062354, 0.01062364, 0.01440181, 0.004804203, 
    0.01152409, 0.005177901, 0.006936624, 0.005214144, 0.007476733, 
    0.005004322, 0.001513509, 0.003361944, 0.009354251, 0.03111353, 
    0.07897718, 0.01445586, 0.03803908, 0.01403831, 0.002089564, 0.01120789, 
    0.04339536,
  0.002877665, 0.005500195, 0.0001642653, 0.003868826, 0.01567796, 0.0255063, 
    0.04999145, 0.01014889, 0.06150441, 0.07733528, 0.02326526, 0.01727371, 
    0.01563009, 0.02030382, 0.0149666, 0.009137824, 0.01691175, 0.008529752, 
    0.00778574, 0.02055485, 0.07490876, 0.2134419, 0.3159299, 0.007286632, 
    0.01644133, 0.04869096, 0.005738514, 0.003978944, 0.01506849,
  2.627232e-09, 2.15245e-09, 3.412639e-10, -0.00231927, 0.06302223, 
    0.01040981, -0.004844478, 0.01132299, 0.003885149, 0.01785305, 
    0.06933158, 0.03071447, 0.01947122, 0.009831525, 0.003805936, 0.01056652, 
    0.01539436, 0.01191902, 0.02602817, 0.03214674, 0.01698056, 0.01095591, 
    0.4051377, 0.1252075, 0.0004472449, 0.004063093, 0.01116682, 0.001976916, 
    0.007565236,
  5.971208e-09, -4.723447e-06, 0.001858599, 0.0002062571, -1.567565e-08, 
    0.001629105, 0.01168541, 0.01134435, 0.01703503, 0.1957104, 0.029767, 
    0.03971159, 0.02685652, 0.01876416, 0.01160641, 0.008537292, 0.01730742, 
    0.0155882, 0.04615311, 0.08784042, 0.03412897, 0.1939707, 0.01051692, 
    0.008390073, 0.01021429, 0.006966095, 0.008706726, 0.0006794668, 
    -9.093038e-08,
  0.00213417, 0.03158517, 0.01980473, 0.02221432, 0.08456941, 0.0004619711, 
    0.001986555, 0.0047568, 0.02595519, 0.07189323, 0.07758999, 0.03156662, 
    0.02856408, 0.06056324, 0.05873989, 0.1115092, 0.1190614, 0.08359754, 
    0.1055549, 0.09174717, 0.08760625, 0.1826657, 0.08169857, 0.07368194, 
    0.05482782, 0.06903973, 0.04055605, 0.05021903, 0.0213398,
  0.03202527, 0.03974572, 0.0639364, 0.3792316, 0.03274129, 0.09345295, 
    0.1166953, 0.007906977, -3.444495e-05, 0.01085891, 0.08200017, 
    0.03455182, 0.06403741, 0.07904902, 0.09189042, 0.1475009, 0.1838385, 
    0.1810651, 0.1690118, 0.3240774, 0.1847927, 0.08522341, 0.2739406, 
    0.1584142, 0.1217598, 0.1269545, 0.1617729, 0.224622, 0.2424959,
  0.2901027, 0.3315141, 0.2811134, 0.3986787, 0.3083356, 0.3460345, 
    0.1402322, 0.1821186, 0.08247004, 0.06074584, 0.07958821, 0.3186223, 
    0.1449968, 0.1226846, 0.2236718, 0.2841823, 0.326712, 0.2472178, 
    0.2285429, 0.3433559, 0.2283191, 0.3193264, 0.3728426, 0.4710443, 
    0.3693046, 0.1719985, 0.1708558, 0.152048, 0.2266673,
  0.1517108, 0.2018015, 0.3792624, 0.561567, 0.5689034, 0.4225561, 0.6613029, 
    0.5723263, 0.4664768, 0.5630785, 0.5319602, 0.2413795, 0.2194131, 
    0.2106342, 0.4098902, 0.2615744, 0.4671555, 0.3939869, 0.377239, 
    0.2446307, 0.4694435, 0.3073539, 0.2961048, 0.2281648, 0.5041742, 
    0.08508254, 0.1567636, 0.1294413, 0.133214,
  0.0794639, 0.06802793, 0.1819637, 0.1718514, 0.4787232, 0.5097504, 
    0.5906305, 0.6289103, 0.3257375, 0.4653155, 0.4949642, 0.3445278, 
    0.4406602, 0.405018, 0.423165, 0.2874797, 0.5086228, 0.4922457, 
    0.3652921, 0.4846283, 0.3225186, 0.2948745, 0.3468755, 0.1268439, 
    0.1166389, 0.4797677, 0.1834205, 0.09454099, 0.1659841,
  0.3260558, 0.3352467, 0.4693394, 0.3740274, 0.3663927, 0.4873881, 0.531741, 
    0.4841294, 0.4272297, 0.4918182, 0.4475165, 0.415322, 0.4291819, 
    0.4937221, 0.4550038, 0.4557477, 0.3500856, 0.2785545, 0.3458179, 
    0.4358035, 0.4032281, 0.2802426, 0.1901889, 0.1569578, 0.1445709, 
    0.150608, 0.2107883, 0.3207015, 0.6193337,
  0.2536884, 0.2625101, 0.2713318, 0.2801535, 0.2889752, 0.2977969, 
    0.3066186, 0.3199387, 0.3169076, 0.3138765, 0.3108454, 0.3078143, 
    0.3047832, 0.3017521, 0.3335117, 0.3298189, 0.3261262, 0.3224334, 
    0.3187406, 0.3150479, 0.3113551, 0.3119568, 0.309859, 0.3077611, 
    0.3056633, 0.3035655, 0.3014677, 0.2993699, 0.2466311,
  0.1949793, 0.2187735, 0.1896527, 0.1715942, 0.1803179, 0.1401722, 
    0.1868592, 0.2159881, 0.1846049, 0.250976, 0.168198, 0.0980401, 
    0.1651051, 0.02325855, 0.1172182, 0.1880957, 0.126596, 0.2144506, 
    0.1212678, 0.0575919, 0.1484421, 0.182211, 0.1555101, 0.05233975, 
    0.14033, 0.1296121, 0.1372677, 0.05305175, 0.1194589,
  0.1547548, 0.1222894, 0.1312942, 0.07865107, 0.04077827, 0.2394329, 
    0.08281113, 0.09558548, 0.1047723, 0.1132889, 0.1166103, 0.1664803, 
    0.07402216, 0.2550264, 0.3992261, 0.4140058, 0.4008605, 0.4027121, 
    0.3456774, 0.4977771, 0.5122849, 0.4637246, 0.5346009, 0.480333, 
    0.3119913, 0.3240933, 0.2804947, 0.1990407, 0.1938172,
  0.3936362, 0.4163586, 0.3113052, 0.3645603, 0.4449884, 0.4716218, 
    0.4516816, 0.3474868, 0.4171771, 0.3854891, 0.3941637, 0.4130597, 
    0.4730161, 0.3731092, 0.3486946, 0.3913441, 0.483895, 0.4965463, 
    0.434112, 0.3163713, 0.2581781, 0.2736992, 0.2564351, 0.2955902, 
    0.3305735, 0.3941264, 0.4567619, 0.4156502, 0.4008431,
  0.3658577, 0.3550189, 0.367578, 0.3316288, 0.3968542, 0.3482223, 0.3182079, 
    0.2861384, 0.2964723, 0.3043573, 0.2094065, 0.161244, 0.1761647, 
    0.2300675, 0.1895837, 0.3001819, 0.3042853, 0.3085929, 0.292724, 
    0.3341572, 0.2901543, 0.2727683, 0.2605484, 0.09976506, 0.07762974, 
    0.2717643, 0.4043462, 0.3841794, 0.3633562,
  0.1610788, 0.09543158, 0.04735848, 0.1368358, 0.1780149, 0.1355524, 
    0.1625677, 0.1957766, 0.1939189, 0.08765439, 0.04971291, 0.02407928, 
    0.05159318, 0.1379757, 0.2011595, 0.07196615, 0.1182425, 0.142295, 
    0.2242431, 0.29116, 0.2058811, 0.1215738, 0.07518138, 0.14065, 
    0.04295262, 0.1397066, 0.290143, 0.2952604, 0.1925821,
  0.01470862, 0.03041565, 0.04051569, 0.03298392, 0.0393323, 0.01156496, 
    0.017674, 0.02512161, 0.0432148, 0.01050725, -3.800494e-05, 
    -9.620006e-08, 0.01912318, 0.016001, 0.04613077, 0.01593954, 0.1059547, 
    0.1712653, 0.05474789, 0.007630756, 0.008730069, 0.004400083, 0.01611607, 
    0.05279607, 0.03811486, 0.04837144, 0.04413103, 0.002987707, 0.005490294,
  0.01340723, 0.1039254, 0.03608262, 0.004822562, -0.002828935, 0.005698185, 
    0.007056867, 0.003139924, 0.03443562, 0.04786661, 0.01906596, 0.01554881, 
    0.01232245, 0.002851873, 0.002776217, 0.03161973, 0.01196977, 0.01301104, 
    0.0001276539, 8.317964e-05, 0.0004150078, 0.001793513, 0.02938643, 
    0.05986558, 0.07298058, 0.07713974, 0.001297883, 5.741612e-05, 0.00093735,
  0.04343237, 0.02136053, 0.09890874, 0.04070746, 0.005506014, 0.002204446, 
    0.002806732, 0.003074104, 0.002176187, 0.001831719, 0.007655224, 
    0.0008197018, 0.001859591, 0.001074529, 0.001992955, 0.001592453, 
    0.004215624, 0.002169729, 0.0003927255, 0.001442142, 0.003471763, 
    0.01198289, 0.03103632, 0.01140919, 0.03516341, 0.01169674, 0.000241572, 
    0.004331002, 0.01546588,
  0.0004810888, 0.005748174, 0.0001072012, 0.004130821, 0.005069328, 
    0.01311986, 0.0283829, 0.00122935, 0.04305748, 0.06228432, 0.00786426, 
    0.005146603, 0.005822583, 0.01201572, 0.00898953, 0.001614927, 
    0.005093846, 0.00195534, 0.001607874, 0.003492439, 0.01924263, 
    0.06576531, 0.09786929, 0.006040086, 0.01008819, 0.03596996, 0.001372923, 
    0.001099009, 0.005287243,
  2.553276e-09, 2.083089e-09, 3.07794e-10, 9.568583e-05, 0.03054313, 
    0.002719318, -0.004052206, 0.003377993, 0.001228645, 0.00477147, 
    0.02916498, 0.01023092, 0.008075319, 0.005164828, 0.0008168257, 
    0.002204457, 0.006152868, 0.002933893, 0.007041288, 0.008748197, 
    0.009281813, 0.005302363, 0.3376071, 0.1027567, 0.0001407385, 
    0.001707462, 0.004890293, 0.001036603, 0.007857486,
  2.553551e-09, -1.921734e-06, 0.0004731294, 6.384484e-05, 4.742756e-09, 
    0.000969769, 0.01078685, 0.004816793, 0.02169875, 0.1228274, 0.01309029, 
    0.02035037, 0.0110232, 0.004858066, 0.003255601, 0.003651786, 
    0.006411479, 0.009661823, 0.02897262, 0.04194529, 0.01375521, 0.1520674, 
    0.004705498, 0.0007059266, 0.002976883, 0.002408074, 0.004290512, 
    0.0002166862, -1.684593e-05,
  0.0009851534, 0.0194767, 0.01373725, 0.01662908, 0.07897273, -0.0003650115, 
    0.001334865, 0.004938737, 0.01855221, 0.062728, 0.05918906, 0.01981793, 
    0.023078, 0.04365957, 0.03952384, 0.09542376, 0.09312339, 0.05215874, 
    0.07455996, 0.05024246, 0.07639144, 0.1605745, 0.07306949, 0.03861601, 
    0.03907717, 0.0499749, 0.01841214, 0.0184137, 0.01594738,
  0.02343141, 0.05240304, 0.04262345, 0.3415418, 0.01726213, 0.09462225, 
    0.106473, 0.0060074, -0.0001008515, 0.008690326, 0.07945763, 0.02256152, 
    0.04826377, 0.06599393, 0.06811476, 0.1289162, 0.1753754, 0.1484143, 
    0.1250305, 0.3020411, 0.1700923, 0.07615265, 0.2302661, 0.1360935, 
    0.08135612, 0.1003578, 0.1194845, 0.1533597, 0.1984363,
  0.2391078, 0.2906691, 0.2473386, 0.3715919, 0.2801132, 0.3253014, 
    0.1125319, 0.1651935, 0.0782493, 0.06514079, 0.07269891, 0.3602928, 
    0.1129253, 0.09374107, 0.1874138, 0.2425802, 0.2887461, 0.2024742, 
    0.1730964, 0.3619522, 0.1995489, 0.2933421, 0.3565795, 0.4924096, 
    0.2867436, 0.1434104, 0.136204, 0.1046365, 0.1933261,
  0.1121184, 0.2120421, 0.4237967, 0.585606, 0.6010963, 0.4493214, 0.6316298, 
    0.5744478, 0.5104143, 0.5761687, 0.5768749, 0.3266889, 0.2332265, 
    0.1984702, 0.3529329, 0.2840418, 0.5182511, 0.3641468, 0.375548, 
    0.2706745, 0.5845637, 0.2807383, 0.3254145, 0.241744, 0.4465213, 
    0.06443219, 0.1307486, 0.09278475, 0.1017035,
  0.05741236, 0.05360517, 0.1673698, 0.1257063, 0.4192911, 0.5570871, 
    0.7108527, 0.5843636, 0.2832929, 0.4866633, 0.5346802, 0.4092719, 
    0.5039126, 0.4373443, 0.4476522, 0.3135854, 0.538053, 0.475017, 
    0.3931633, 0.4952393, 0.2991782, 0.3736982, 0.3988809, 0.1622278, 
    0.1136331, 0.4268917, 0.2010034, 0.07769167, 0.1340293,
  0.4529053, 0.3955057, 0.5157622, 0.449497, 0.4303896, 0.5466928, 0.5760503, 
    0.5451746, 0.5597475, 0.5908099, 0.5080217, 0.4801794, 0.5186751, 
    0.5408918, 0.4925359, 0.4871478, 0.4146823, 0.3475587, 0.4165491, 
    0.5115117, 0.4800504, 0.2703778, 0.2306089, 0.2236591, 0.1392694, 
    0.1414717, 0.1755045, 0.3003565, 0.6374703,
  0.2592213, 0.268535, 0.2778487, 0.2871624, 0.2964761, 0.3057898, 0.3151035, 
    0.2939279, 0.2922776, 0.2906272, 0.2889769, 0.2873266, 0.2856763, 
    0.284026, 0.3274534, 0.3209032, 0.314353, 0.3078029, 0.3012527, 
    0.2947025, 0.2881523, 0.3005286, 0.2994155, 0.2983023, 0.2971891, 
    0.2960759, 0.2949627, 0.2938495, 0.2517703,
  0.1368654, 0.1647114, 0.1338, 0.1340621, 0.1287189, 0.1010629, 0.1424503, 
    0.1728002, 0.1471555, 0.1827763, 0.1019382, 0.06098276, 0.1063533, 
    0.02294389, 0.09499449, 0.1315207, 0.1052254, 0.1747339, 0.07997862, 
    0.0332953, 0.1072772, 0.1429807, 0.1122472, 0.04360251, 0.1420134, 
    0.1063414, 0.1058943, 0.03684676, 0.08234207,
  0.1114323, 0.09584293, 0.08924607, 0.05484293, 0.02364691, 0.185947, 
    0.07833945, 0.06430091, 0.07522008, 0.08229971, 0.08036155, 0.1292882, 
    0.05592185, 0.2022952, 0.3221031, 0.3493292, 0.3099416, 0.3332735, 
    0.2818542, 0.433207, 0.4396792, 0.4351508, 0.4816661, 0.4611339, 
    0.2834837, 0.2913642, 0.2398474, 0.1491595, 0.1459189,
  0.3373397, 0.3446528, 0.2521034, 0.2975829, 0.3494734, 0.3840209, 
    0.3762645, 0.2716609, 0.3344622, 0.3292292, 0.3435919, 0.3648609, 
    0.4437106, 0.3214256, 0.2919562, 0.3383292, 0.42862, 0.4530987, 
    0.3883651, 0.2604567, 0.2094503, 0.2068738, 0.1866529, 0.2263891, 
    0.29194, 0.3567115, 0.4207363, 0.3482904, 0.3350359,
  0.3034128, 0.2780791, 0.3036667, 0.292906, 0.3519667, 0.3033719, 0.2703372, 
    0.230135, 0.231225, 0.23419, 0.1541052, 0.1138218, 0.1416752, 0.1934564, 
    0.1814157, 0.2702783, 0.2427917, 0.2477573, 0.220818, 0.2738205, 
    0.2311577, 0.2142123, 0.2141344, 0.07518931, 0.07057483, 0.2822602, 
    0.3627924, 0.3289675, 0.3134753,
  0.1121423, 0.05568544, 0.03104667, 0.1163475, 0.1515329, 0.09583759, 
    0.1258899, 0.1634016, 0.1537475, 0.05075858, 0.0291684, 0.01586896, 
    0.04179941, 0.09843998, 0.1808225, 0.04047259, 0.08867136, 0.1082051, 
    0.1862852, 0.239711, 0.1371628, 0.07653734, 0.03865336, 0.1354069, 
    0.04352497, 0.1014036, 0.2550676, 0.2399383, 0.1374701,
  0.006726057, 0.01432313, 0.02655945, 0.01498189, 0.02120781, 0.002378236, 
    0.006605986, 0.01573396, 0.01921837, 0.007280114, -1.723392e-05, 
    -3.798311e-09, 0.01461428, 0.005563318, 0.02262292, 0.00664302, 
    0.07478274, 0.10303, 0.0413686, 0.002668449, 0.003307229, 0.002221894, 
    0.00889216, 0.0319014, 0.02777269, 0.0326865, 0.02509703, 0.001583863, 
    0.002878549,
  0.005860194, 0.0842469, 0.02340347, 0.001641098, -0.002898327, 0.001694951, 
    0.003006027, 0.001783555, 0.01781353, 0.01943086, 0.01180361, 0.0102049, 
    0.003648373, 0.0009156014, 0.001062176, 0.01609082, 0.003583263, 
    0.007206396, 5.66146e-05, 4.063332e-05, 0.0002362719, 0.0008601247, 
    0.01255476, 0.03263857, 0.06012036, 0.06282651, 0.0005365846, 
    2.348164e-05, 0.0004370346,
  0.02241969, 0.009276308, 0.09177661, 0.02533309, 0.002910547, 0.0007643519, 
    0.0008624797, 0.000922858, 0.0009820913, 0.0002636819, 0.003443229, 
    0.000362428, 0.0001779313, 0.0003682568, 0.0009700722, 0.0005667856, 
    0.00249943, 0.001177397, 0.0002131043, 0.0008446752, 0.00195214, 
    0.006603251, 0.01682937, 0.009458497, 0.03971647, 0.009860434, 
    0.0001839225, 0.002390305, 0.00794165,
  0.0002076328, 0.003757966, 5.261816e-05, 0.005854626, 0.0009659025, 
    0.007473576, 0.01231105, 0.0003955951, 0.04352751, 0.0621731, 
    0.003483715, 0.002218408, 0.003497381, 0.007140625, 0.006647191, 
    0.0006022978, 0.002582126, 0.0005552315, 0.0004708895, 0.001053115, 
    0.004269311, 0.02092643, 0.04175518, 0.005949504, 0.006378981, 
    0.02026115, 0.0004789623, 0.0005215774, 0.002775001,
  2.544688e-09, 2.058791e-09, 3.044158e-10, 0.001691984, 0.01695262, 
    0.001036102, -0.003302926, 0.00175562, 0.0007494849, 0.0007488384, 
    0.01156049, 0.002855516, 0.003258609, 0.002518686, 0.0003649741, 
    0.0006959662, 0.002492348, 0.00122863, 0.002535987, 0.003447919, 
    0.005500752, 0.003647872, 0.2497781, 0.08007941, 6.780543e-05, 
    0.0009541953, 0.002782098, 0.0006626672, 0.008009718,
  1.309768e-09, -9.993747e-07, 0.0001674791, 5.807994e-05, 1.261098e-08, 
    0.0006711065, 0.01041409, 0.002203953, 0.03159825, 0.07106911, 
    0.005668645, 0.01062042, 0.005222302, 0.002158861, 0.001654064, 
    0.001870645, 0.002798263, 0.004084043, 0.01976336, 0.01854275, 
    0.007663942, 0.1144909, 0.002730862, -0.001056885, 0.001333794, 
    0.001093712, 0.002649251, 0.0001220285, -1.168224e-05,
  0.0003669357, 0.01397256, 0.009350991, 0.01149199, 0.07004367, 
    -0.0005223413, 0.0007441804, 0.006517274, 0.01314288, 0.0503557, 
    0.04749476, 0.01133664, 0.0133921, 0.0284533, 0.02474604, 0.06992249, 
    0.06547249, 0.02964536, 0.04106348, 0.02999025, 0.06598331, 0.1425488, 
    0.06721684, 0.01884052, 0.0243255, 0.03089785, 0.008423185, 0.009838128, 
    0.01093349,
  0.01473019, 0.03934795, 0.03044934, 0.3052179, 0.01039104, 0.07746057, 
    0.09818099, 0.004416741, -0.0001004498, 0.008048595, 0.07173036, 
    0.01685508, 0.03719444, 0.05416181, 0.04574607, 0.1030387, 0.1487536, 
    0.1160289, 0.08349798, 0.2800588, 0.1561031, 0.06837574, 0.1918788, 
    0.1155884, 0.05345801, 0.0729591, 0.07791001, 0.08645315, 0.1437232,
  0.176686, 0.2573365, 0.1863239, 0.3275009, 0.2456501, 0.280857, 0.09108973, 
    0.1465187, 0.06677756, 0.07241627, 0.05600591, 0.4040199, 0.09017674, 
    0.07334487, 0.1553852, 0.2073312, 0.2510162, 0.1515993, 0.1178465, 
    0.3741647, 0.1714075, 0.214563, 0.3054898, 0.5139518, 0.2263941, 
    0.1184701, 0.1061827, 0.07658285, 0.1512969,
  0.07119755, 0.2261485, 0.4044608, 0.5581993, 0.5945297, 0.4108865, 
    0.559572, 0.5063362, 0.5024325, 0.5415617, 0.6113597, 0.4048072, 
    0.2443451, 0.2191631, 0.2986774, 0.2937591, 0.5501906, 0.3227296, 
    0.3415552, 0.3053823, 0.6576406, 0.2728996, 0.3004649, 0.2393816, 
    0.4052505, 0.04811446, 0.1078574, 0.06446069, 0.072947,
  0.04382493, 0.04204669, 0.1786416, 0.09198251, 0.3807225, 0.5681355, 
    0.7189896, 0.5392497, 0.2629639, 0.5345521, 0.598839, 0.4370015, 
    0.6701343, 0.4614206, 0.4446969, 0.3118989, 0.4953461, 0.4243622, 
    0.3700405, 0.4571023, 0.3237397, 0.4616559, 0.4803228, 0.2237199, 
    0.1604153, 0.3686774, 0.2197104, 0.07282104, 0.103267,
  0.4928001, 0.4202574, 0.5362493, 0.4907686, 0.517794, 0.6038891, 0.5891665, 
    0.6007534, 0.6653339, 0.6601412, 0.5738786, 0.5973524, 0.6122004, 
    0.5656086, 0.5008293, 0.4872251, 0.4901966, 0.4359174, 0.4974105, 
    0.549027, 0.495777, 0.2774852, 0.2512555, 0.2991177, 0.1136514, 
    0.1366446, 0.1464693, 0.2488719, 0.6219578,
  0.205179, 0.2146974, 0.2242157, 0.2337341, 0.2432524, 0.2527707, 0.2622891, 
    0.219348, 0.2199554, 0.2205628, 0.2211702, 0.2217776, 0.2223849, 
    0.2229923, 0.2872248, 0.2789463, 0.2706679, 0.2623895, 0.254111, 
    0.2458326, 0.2375541, 0.2358609, 0.2340136, 0.2321663, 0.2303191, 
    0.2284718, 0.2266245, 0.2247772, 0.1975644,
  0.09926781, 0.1124239, 0.0969225, 0.1073858, 0.1113435, 0.07104945, 
    0.1080507, 0.1346556, 0.1221099, 0.1336375, 0.06974246, 0.03576645, 
    0.06104307, 0.01953409, 0.07075977, 0.07863445, 0.07744497, 0.136908, 
    0.05983263, 0.01990745, 0.07942799, 0.1100037, 0.08255985, 0.0379023, 
    0.1293496, 0.08953454, 0.08019353, 0.02736265, 0.0578571,
  0.0731295, 0.06869669, 0.06320189, 0.03934713, 0.01529002, 0.1470695, 
    0.06329645, 0.04441103, 0.05592768, 0.0687834, 0.05565286, 0.1031125, 
    0.04286831, 0.1533133, 0.2537922, 0.2776791, 0.2435051, 0.2587734, 
    0.2094162, 0.3202177, 0.3475267, 0.3781253, 0.4344377, 0.398175, 
    0.2395727, 0.2464985, 0.1928601, 0.1067824, 0.1092417,
  0.2606877, 0.2573261, 0.1822732, 0.2256136, 0.2617234, 0.2890595, 
    0.2867336, 0.2062434, 0.2598984, 0.2712768, 0.2759036, 0.2897485, 
    0.3707398, 0.2441864, 0.2171767, 0.266818, 0.3521253, 0.38766, 0.320527, 
    0.1962937, 0.1522065, 0.143073, 0.1255873, 0.1505019, 0.2371882, 
    0.2977241, 0.3402208, 0.2702813, 0.2517658,
  0.2391792, 0.2066005, 0.2256339, 0.2314755, 0.2853834, 0.2486863, 
    0.2121046, 0.1721309, 0.1756012, 0.1619871, 0.09639071, 0.06786978, 
    0.101745, 0.1404138, 0.1481163, 0.1997811, 0.171728, 0.1782434, 
    0.1571715, 0.2027946, 0.1596193, 0.1499573, 0.1543735, 0.05736557, 
    0.05276083, 0.2565978, 0.3071111, 0.2682265, 0.2539166,
  0.07269754, 0.03080521, 0.02048839, 0.08455519, 0.1105355, 0.05823007, 
    0.08653174, 0.125581, 0.1129007, 0.03218745, 0.01941262, 0.009893101, 
    0.0335974, 0.06465763, 0.1578179, 0.02248276, 0.05679493, 0.07942909, 
    0.152945, 0.1815553, 0.08634321, 0.04042757, 0.0193352, 0.1236966, 
    0.03863512, 0.07148007, 0.1875318, 0.1582479, 0.08835308,
  0.004166952, 0.00715645, 0.01444345, 0.006463503, 0.01021398, 0.001071375, 
    0.002671774, 0.009868528, 0.01118913, 0.004317867, -1.127066e-05, 
    1.565665e-08, 0.009951252, 0.002484143, 0.01015924, 0.003274594, 
    0.04524103, 0.06447323, 0.01954928, 0.001392562, 0.002018622, 
    0.001482429, 0.006041174, 0.02103034, 0.01850493, 0.01543719, 0.01037129, 
    0.001024029, 0.001928042,
  0.003486601, 0.05407507, 0.01371916, 0.0009031215, -0.002217371, 
    0.0006552068, 0.001123331, 0.001193121, 0.01117629, 0.01020513, 
    0.007124713, 0.00502922, 0.001416554, 0.0005131271, 0.0006423516, 
    0.005990322, 0.001140829, 0.002958189, 3.601149e-05, 2.714347e-05, 
    0.0001613966, 0.0005184336, 0.006995118, 0.02161768, 0.04418892, 
    0.04854951, 0.0002980359, 1.276279e-05, 0.0002677486,
  0.0144975, 0.005494251, 0.08399136, 0.01880096, 0.001479828, 0.0004259076, 
    0.0004575846, 0.0003131428, 0.0006423782, 0.0001064589, 0.001527151, 
    0.0002248047, 6.93952e-05, 0.0002202359, 0.0004589965, 0.0002826605, 
    0.001203678, 0.0007475551, 0.0001379204, 0.0005740492, 0.001294664, 
    0.004377785, 0.01110433, 0.008157399, 0.03348646, 0.006925186, 
    0.0001143545, 0.001567571, 0.005057802,
  0.0001170111, 0.003106534, 3.28053e-05, 0.005212445, 0.0003973968, 
    0.003810693, 0.005180046, 0.0002363076, 0.04689842, 0.05740205, 
    0.001681181, 0.001217782, 0.001620914, 0.003128942, 0.003844246, 
    0.0003483785, 0.0009358774, 0.0003526817, 0.0002544178, 0.000548392, 
    0.002039404, 0.0109268, 0.02360645, 0.005637196, 0.004505264, 
    0.009876692, 0.0001748732, 0.0003134474, 0.001691685,
  2.634219e-09, 2.061034e-09, 3.086545e-10, 0.002059387, 0.009234235, 
    0.0006242352, -0.002195988, 0.001140155, 0.0004685404, 0.0001738611, 
    0.004697284, 0.001034482, 0.001259255, 0.001159337, 0.0002400459, 
    0.0003790009, 0.0009620728, 0.000429424, 0.001150567, 0.00146603, 
    0.002618555, 0.001917323, 0.1926041, 0.0622299, 5.301559e-05, 
    0.0006260001, 0.001856453, 0.0004755651, 0.007244234,
  2.123595e-09, -6.051563e-07, 9.893092e-05, 6.517291e-05, -3.073962e-08, 
    0.0005106855, 0.009246325, 0.001234913, 0.03190507, 0.04402295, 
    0.002792709, 0.006406594, 0.002579625, 0.001417481, 0.001081838, 
    0.001279023, 0.001647371, 0.001112341, 0.01390296, 0.01035698, 
    0.005242371, 0.08837334, 0.001892528, -0.001255363, 0.0009100524, 
    0.000663834, 0.001869206, 8.190496e-05, -7.905294e-06,
  0.0002266037, 0.01059354, 0.005748907, 0.006367262, 0.06146424, 
    -0.000503137, 0.001540718, 0.01063988, 0.01173911, 0.0356486, 0.03635353, 
    0.006384895, 0.007180612, 0.01565791, 0.01354966, 0.04431286, 0.03836879, 
    0.01592617, 0.01945379, 0.01527069, 0.05360045, 0.1210223, 0.05843628, 
    0.009914425, 0.01295164, 0.01705886, 0.00419817, 0.00607132, 0.007422413,
  0.01017702, 0.03220239, 0.02237065, 0.2722244, 0.007054697, 0.06102643, 
    0.0890111, 0.003949258, -0.0001027478, 0.01026241, 0.05982862, 
    0.01294674, 0.02774259, 0.04038535, 0.02872096, 0.07385651, 0.1057201, 
    0.08314851, 0.05218626, 0.2551761, 0.1395961, 0.0568801, 0.1627509, 
    0.09729032, 0.03560284, 0.05005008, 0.04797769, 0.04541682, 0.09475937,
  0.1294334, 0.2230209, 0.1488723, 0.2795237, 0.2020347, 0.2351416, 
    0.07552835, 0.1326063, 0.06937022, 0.07910701, 0.04035083, 0.4190227, 
    0.07657292, 0.05894267, 0.1252434, 0.1669668, 0.1997798, 0.105325, 
    0.07737009, 0.3599298, 0.1321459, 0.1508847, 0.2463817, 0.5035851, 
    0.1809348, 0.09862526, 0.07937077, 0.05038145, 0.1051312,
  0.04094379, 0.2526487, 0.3722513, 0.4948523, 0.5681466, 0.3514476, 
    0.4723992, 0.3931419, 0.4511447, 0.4511316, 0.5437455, 0.4848644, 
    0.2776753, 0.2334063, 0.2547867, 0.2900612, 0.56407, 0.2929758, 
    0.3130152, 0.2961445, 0.6618838, 0.3219115, 0.2502406, 0.2461821, 
    0.3737814, 0.03595051, 0.08186267, 0.04705602, 0.05088973,
  0.03391021, 0.03253721, 0.2107244, 0.07210853, 0.3374093, 0.4990838, 
    0.6828372, 0.4988067, 0.3288135, 0.5880042, 0.6294672, 0.3890021, 
    0.697306, 0.418422, 0.3928913, 0.2696024, 0.4390789, 0.3609589, 
    0.2917844, 0.379171, 0.2803102, 0.4633755, 0.5429958, 0.3247894, 
    0.1879358, 0.3143445, 0.2498603, 0.06231071, 0.0805883,
  0.5150365, 0.4287205, 0.494777, 0.475116, 0.5438295, 0.5654393, 0.5115182, 
    0.5256301, 0.5743338, 0.6045482, 0.5372393, 0.6116063, 0.6280143, 
    0.5660309, 0.4830001, 0.451636, 0.4803477, 0.4570196, 0.4745633, 
    0.5186555, 0.5116649, 0.2739977, 0.2502803, 0.3600592, 0.08469029, 
    0.1232385, 0.1337036, 0.2360692, 0.5385273,
  0.1280798, 0.1349047, 0.1417295, 0.1485544, 0.1553793, 0.1622041, 0.169029, 
    0.1441011, 0.1461674, 0.1482337, 0.1503, 0.1523664, 0.1544327, 0.156499, 
    0.2075291, 0.201029, 0.1945289, 0.1880288, 0.1815287, 0.1750287, 
    0.1685286, 0.1638061, 0.161415, 0.1590239, 0.1566328, 0.1542417, 
    0.1518506, 0.1494595, 0.1226199,
  0.07581176, 0.08558665, 0.07363965, 0.09560151, 0.09889228, 0.05390116, 
    0.07617884, 0.1164697, 0.1011024, 0.1036815, 0.05651842, 0.02445537, 
    0.04079669, 0.01585031, 0.05747084, 0.05196247, 0.05482586, 0.1153634, 
    0.05012497, 0.01514536, 0.06294859, 0.09241745, 0.06106263, 0.0357739, 
    0.1189393, 0.07953518, 0.0695686, 0.02355593, 0.04767495,
  0.05239005, 0.05282725, 0.04744016, 0.0322744, 0.01223981, 0.1221233, 
    0.05361958, 0.03537526, 0.04549562, 0.06242901, 0.04093766, 0.08677974, 
    0.03623955, 0.120272, 0.1932418, 0.2135982, 0.1908041, 0.2033116, 
    0.1644337, 0.2412395, 0.2738399, 0.3062915, 0.353515, 0.3364107, 
    0.2035107, 0.2029707, 0.1516824, 0.08429143, 0.07928991,
  0.2062209, 0.1981324, 0.1383141, 0.1783549, 0.2051195, 0.2294825, 
    0.2279272, 0.1598968, 0.207082, 0.2229145, 0.2196207, 0.2296896, 
    0.3004377, 0.1854753, 0.1594299, 0.2048881, 0.2806253, 0.3188519, 
    0.2553979, 0.1470824, 0.1128755, 0.09919478, 0.08922506, 0.0999738, 
    0.1826707, 0.2334689, 0.2684937, 0.21148, 0.1961728,
  0.1893855, 0.1611429, 0.1724218, 0.1853402, 0.2377826, 0.2170977, 
    0.1758046, 0.1367696, 0.13849, 0.1200327, 0.06305019, 0.04453961, 
    0.07170751, 0.09723005, 0.1161206, 0.1456287, 0.1196439, 0.1233805, 
    0.1175606, 0.1553179, 0.1138474, 0.1110145, 0.1152059, 0.04769466, 
    0.03865339, 0.2129222, 0.2562405, 0.2215313, 0.2143564,
  0.04920758, 0.01901172, 0.01405391, 0.05549666, 0.07642769, 0.0352376, 
    0.05637272, 0.09406745, 0.07624871, 0.02196882, 0.01235083, 0.005878428, 
    0.02780791, 0.04118951, 0.1373262, 0.01419674, 0.03427338, 0.05477588, 
    0.1117241, 0.1286139, 0.05538379, 0.02146197, 0.01185285, 0.1142874, 
    0.02922596, 0.05031659, 0.1274385, 0.1075933, 0.05832858,
  0.003035091, 0.00448798, 0.009342537, 0.003545547, 0.006084024, 
    0.0007334017, 0.001655641, 0.006117017, 0.008197564, 0.003132664, 
    -8.673891e-06, 2.012772e-08, 0.007824126, 0.001586006, 0.005576766, 
    0.002107009, 0.02825089, 0.03782324, 0.009961769, 0.0009648607, 
    0.001467852, 0.001124347, 0.004630326, 0.0159245, 0.01308289, 
    0.007424725, 0.005179503, 0.0007519793, 0.001463306,
  0.002454907, 0.03844538, 0.007661967, 0.0006449014, -0.001612525, 
    0.0003513205, 0.0005714754, 0.0008901032, 0.00807356, 0.006885108, 
    0.004064719, 0.002520606, 0.0007285997, 0.0003450315, 0.0004581615, 
    0.002673673, 0.0004991796, 0.001255527, 2.632919e-05, 2.039543e-05, 
    0.0001239266, 0.0003642004, 0.00469391, 0.016341, 0.02845092, 0.04037175, 
    0.0002086265, 7.947524e-06, 0.0001908774,
  0.01071737, 0.003844338, 0.07216355, 0.02547343, 0.0008415638, 
    0.0002997592, 0.0003298294, 0.0001531345, 0.0004779455, 0.0001434366, 
    0.0009566178, 0.0001621538, 7.369411e-05, 0.0001623166, 0.0002529786, 
    0.0001930719, 0.0006090397, 0.0005183337, 0.0001009768, 0.0004363719, 
    0.0009709012, 0.003279772, 0.008306669, 0.01081633, 0.02325852, 
    0.005851236, 4.323652e-05, 0.001164831, 0.003687798,
  7.876154e-05, 0.003744517, 0.0001851757, 0.004476049, 0.0002549353, 
    0.002068565, 0.002508035, 0.0001712377, 0.0488898, 0.06393039, 
    0.0009706656, 0.0008153801, 0.0008418546, 0.001480059, 0.001903236, 
    0.0002415625, 0.000425776, 0.0002552894, 0.0001652913, 0.0003584573, 
    0.001307679, 0.007202539, 0.01574315, 0.006176271, 0.003918801, 
    0.004796837, 0.0001103696, 0.0002192208, 0.001212543,
  2.783038e-09, 2.090162e-09, 3.161135e-10, 0.003784936, 0.005925314, 
    0.0004525592, -0.001429358, 0.0008670634, 0.0002270779, 0.0001048495, 
    0.002400407, 0.0005147489, 0.0005711884, 0.0005226892, 0.0001808831, 
    0.0002819921, 0.0005195232, 0.0002116149, 0.0006629003, 0.000737428, 
    0.001211805, 0.0009485252, 0.1439034, 0.04465713, 4.421566e-05, 
    0.0004652589, 0.001393289, 0.000375197, 0.0052003,
  2.518273e-09, -4.227364e-07, 7.237867e-05, 6.111981e-05, -1.001054e-06, 
    0.0004179125, 0.008088279, 0.0009169835, 0.02987184, 0.03116892, 
    0.001852628, 0.003849702, 0.00143613, 0.001105887, 0.0008079709, 
    0.001003371, 0.001203537, 0.0006829753, 0.008630985, 0.00728544, 
    0.003695971, 0.07328855, 0.001465922, -0.001152466, 0.0006486638, 
    0.0004912459, 0.001458635, 6.218254e-05, -1.202783e-05,
  0.000164005, 0.008841101, 0.003931305, 0.004348515, 0.05572545, 
    -0.0004546254, 0.002834156, 0.01817033, 0.01199751, 0.02565989, 
    0.02879786, 0.003899931, 0.00398444, 0.007034717, 0.007305022, 
    0.02676494, 0.02512269, 0.008790108, 0.0116889, 0.009969343, 0.04863261, 
    0.09950403, 0.04968132, 0.006399958, 0.007408005, 0.009426446, 
    0.002767508, 0.00440804, 0.005864284,
  0.007556377, 0.02896076, 0.01704008, 0.2500888, 0.005601109, 0.05064097, 
    0.08119808, 0.004749564, -0.0001203807, 0.01706933, 0.05931484, 
    0.01067578, 0.02161977, 0.03156801, 0.02039096, 0.05298954, 0.07066061, 
    0.05960941, 0.03407921, 0.2315924, 0.131016, 0.05092108, 0.1489147, 
    0.08918241, 0.02624718, 0.03389861, 0.0316647, 0.02646697, 0.06578402,
  0.09645738, 0.2065234, 0.1434536, 0.2548544, 0.1771731, 0.2026042, 
    0.06777175, 0.1460289, 0.1141503, 0.07576665, 0.03313962, 0.4043522, 
    0.06760533, 0.04888449, 0.09684359, 0.1328015, 0.1568731, 0.08072869, 
    0.05702173, 0.3503452, 0.1099148, 0.1208832, 0.2094371, 0.471762, 
    0.1555772, 0.08403534, 0.06095645, 0.03426035, 0.07202348,
  0.02749714, 0.2891639, 0.3527533, 0.4413709, 0.5260563, 0.3064304, 
    0.3921088, 0.3230312, 0.371089, 0.377582, 0.4747163, 0.5694089, 
    0.3371334, 0.2577637, 0.2248314, 0.2850159, 0.5563264, 0.2761148, 
    0.3357764, 0.302228, 0.6071366, 0.3604581, 0.1874185, 0.2190479, 
    0.3523826, 0.02932821, 0.06277242, 0.03622617, 0.03681323,
  0.02812163, 0.02610879, 0.2903067, 0.06104568, 0.3076029, 0.3929377, 
    0.6366181, 0.4517502, 0.418005, 0.5891129, 0.6705371, 0.3692319, 
    0.5777879, 0.2982794, 0.3115926, 0.2433324, 0.3827317, 0.2982786, 
    0.2440016, 0.2561641, 0.2395885, 0.3999963, 0.4545449, 0.3350139, 
    0.1918209, 0.2422575, 0.3218993, 0.06186986, 0.06805703,
  0.5045267, 0.4286029, 0.436143, 0.3668942, 0.4300033, 0.4402534, 0.3291502, 
    0.2757971, 0.3992252, 0.3964219, 0.330214, 0.3972755, 0.4080541, 
    0.3583299, 0.3315454, 0.3076576, 0.3706087, 0.4051112, 0.2989962, 
    0.3365735, 0.3439315, 0.2529713, 0.2796953, 0.4244444, 0.1112572, 
    0.09976387, 0.1258474, 0.2163888, 0.4188606,
  0.08229835, 0.08714278, 0.09198721, 0.09683163, 0.1016761, 0.1065205, 
    0.1113649, 0.09544677, 0.09801844, 0.1005901, 0.1031618, 0.1057335, 
    0.1083051, 0.1108768, 0.1522639, 0.146855, 0.1414461, 0.1360372, 
    0.1306284, 0.1252195, 0.1198106, 0.1096476, 0.1076404, 0.1056332, 
    0.1036259, 0.1016187, 0.09961152, 0.0976043, 0.07842281,
  0.07103452, 0.07896355, 0.07284175, 0.113088, 0.132664, 0.04448023, 
    0.06416783, 0.1226584, 0.1184096, 0.1001848, 0.05011158, 0.01964358, 
    0.03172742, 0.01352851, 0.05768443, 0.04462408, 0.04459564, 0.1048396, 
    0.04576419, 0.01641565, 0.05484528, 0.08106421, 0.04991084, 0.03500421, 
    0.1155174, 0.07315388, 0.06361893, 0.02175984, 0.05028401,
  0.04504492, 0.04506553, 0.04050805, 0.03351189, 0.0103937, 0.1121359, 
    0.05459694, 0.03451482, 0.04754312, 0.05860652, 0.03530362, 0.08545913, 
    0.03430784, 0.10829, 0.1593035, 0.1780617, 0.1562271, 0.173051, 
    0.1411184, 0.2051461, 0.2328754, 0.2559127, 0.3096252, 0.29606, 
    0.1838648, 0.1728433, 0.1248132, 0.06842886, 0.06295833,
  0.173661, 0.1668966, 0.1099122, 0.1484315, 0.1737421, 0.1916478, 0.19337, 
    0.1322166, 0.1760199, 0.1889673, 0.1816715, 0.1845202, 0.2535819, 
    0.146877, 0.1215572, 0.1663036, 0.2279236, 0.2674287, 0.213066, 
    0.1188344, 0.09228379, 0.0760095, 0.07038425, 0.07561551, 0.1395975, 
    0.1905988, 0.2279802, 0.1743158, 0.167426,
  0.160123, 0.135922, 0.1431549, 0.1498849, 0.1941811, 0.1768397, 0.1459109, 
    0.1137344, 0.1159728, 0.09853758, 0.04760965, 0.03337712, 0.05421558, 
    0.06935487, 0.09025604, 0.1172, 0.08491846, 0.09075903, 0.09123196, 
    0.1227996, 0.08965435, 0.08342866, 0.08974849, 0.04989092, 0.03121044, 
    0.1750763, 0.2081988, 0.1899302, 0.1827977,
  0.03697362, 0.01385895, 0.009324593, 0.03794055, 0.05598338, 0.02438173, 
    0.03803413, 0.07040421, 0.05305453, 0.01762233, 0.008998352, 0.004518178, 
    0.02186368, 0.02859661, 0.1359642, 0.009147419, 0.02195571, 0.03756616, 
    0.07679932, 0.08635094, 0.03894107, 0.01324939, 0.008536939, 0.1158503, 
    0.02288476, 0.03500519, 0.09558453, 0.07937846, 0.04244658,
  0.00249697, 0.003376821, 0.01098935, 0.002541916, 0.004286084, 
    0.0005912328, 0.001303688, 0.003932873, 0.006822037, 0.002552489, 
    -6.796043e-06, 2.218022e-08, 0.01030303, 0.001229267, 0.003786359, 
    0.001657476, 0.01948018, 0.02466455, 0.006389606, 0.0007590398, 
    0.001202033, 0.0009389292, 0.003876826, 0.01336772, 0.01847039, 
    0.004040756, 0.003257624, 0.0006202051, 0.001227038,
  0.00199827, 0.03060498, 0.005733823, 0.0005231763, -0.001435985, 
    0.0002455613, 0.0003865069, 0.0007460889, 0.00661719, 0.005409119, 
    0.002667763, 0.002180401, 0.000461237, 0.000277046, 0.0003723267, 
    0.001626275, 0.0003429848, 0.0007090251, 2.154495e-05, 1.707992e-05, 
    0.0001043546, 0.0002916561, 0.003709459, 0.01326949, 0.03731859, 
    0.09331492, 0.0001676054, 6.326332e-06, 0.0001554814,
  0.008813329, 0.003021456, 0.104368, 0.08607456, 0.0005680131, 0.0002364616, 
    0.0002721047, 0.0001140111, 0.0003958581, 0.0001111361, 0.000747769, 
    0.0001292591, 7.049255e-05, 0.0001315707, 0.0001850801, 0.0001501424, 
    0.0004087838, 0.0004191047, 8.259187e-05, 0.0003679978, 0.0008133958, 
    0.002732253, 0.006878773, 0.1222079, 0.0663238, 0.04580519, 6.01861e-05, 
    0.0009716422, 0.003019812,
  5.602051e-05, 0.02087948, 0.003291655, 0.005180391, 0.0001928146, 
    0.001433261, 0.001733996, 0.0001382659, 0.0840304, 0.112305, 
    0.0007217299, 0.0006378493, 0.0006068844, 0.0009022283, 0.001257659, 
    0.0001960661, 0.0002701505, 0.000210923, 0.0001290515, 0.0002789098, 
    0.001005032, 0.005504403, 0.0122447, 0.0464327, 0.03000004, 0.002922605, 
    8.930289e-05, 0.0001745108, 0.0009961366,
  2.892327e-09, 2.139248e-09, 3.250243e-10, 0.00535962, 0.004491711, 
    0.0003768916, -0.0009639867, 0.0007315568, -0.0001068299, 7.979079e-05, 
    0.001537124, 0.0003544338, 0.0003838118, 0.0003299247, 0.0001503124, 
    0.0002379973, 0.0003987871, 0.0001567645, 0.0004733179, 0.0004950177, 
    0.0006711294, 0.0006240795, 0.1503181, 0.03759378, 3.917055e-05, 
    0.0003956294, 0.001184002, 0.000324676, 0.003711408,
  3.04962e-09, -3.459838e-07, 5.636689e-05, 5.705114e-05, -1.325488e-07, 
    0.0003676525, 0.006800889, 0.0007383875, 0.03145495, 0.02348546, 
    0.001446358, 0.002630587, 0.00106811, 0.0009315931, 0.0006757543, 
    0.0008641621, 0.0009935156, 0.0005200171, 0.00583799, 0.005957263, 
    0.002562678, 0.06593294, 0.001253429, -0.001195468, 0.0005420121, 
    0.0004075678, 0.001249855, 5.312265e-05, -8.092386e-06,
  0.0001328417, 0.007553572, 0.003022664, 0.003968502, 0.05332475, 
    -0.0004182862, 0.002350328, 0.05904754, 0.01881612, 0.02205745, 
    0.02389692, 0.002996747, 0.002694804, 0.00413194, 0.004767567, 
    0.01828127, 0.01754648, 0.005649257, 0.008486723, 0.00760533, 0.04363346, 
    0.09010652, 0.05532606, 0.004905703, 0.004843009, 0.006256507, 
    0.002219599, 0.003662412, 0.00510788,
  0.006657932, 0.02677203, 0.01436324, 0.2524452, 0.004999268, 0.04431697, 
    0.07731526, 0.007451997, -0.000190506, 0.02625334, 0.07194079, 
    0.009748943, 0.01877185, 0.0257736, 0.01704923, 0.04151003, 0.05409348, 
    0.04610667, 0.0258503, 0.2296115, 0.1406157, 0.05085345, 0.1489007, 
    0.08439858, 0.02217009, 0.02509198, 0.02377874, 0.01765148, 0.05478143,
  0.08034253, 0.2201353, 0.1677528, 0.2401531, 0.1629493, 0.1858269, 
    0.06594315, 0.2578296, 0.2221679, 0.09381512, 0.0532519, 0.4369355, 
    0.06356053, 0.0416146, 0.08043499, 0.1108684, 0.1290462, 0.0678943, 
    0.04631786, 0.3697694, 0.1056113, 0.1242628, 0.2189641, 0.469164, 
    0.1518464, 0.07501744, 0.05153375, 0.02607167, 0.05339959,
  0.02185907, 0.4088458, 0.3555756, 0.4201289, 0.5447454, 0.3358525, 
    0.3752497, 0.3357601, 0.4618537, 0.4230668, 0.4680983, 0.5979261, 
    0.4314725, 0.2967711, 0.213871, 0.2828559, 0.56673, 0.2903566, 0.4050012, 
    0.3710156, 0.5807757, 0.4122257, 0.1642001, 0.2472602, 0.3432155, 
    0.0293445, 0.05237206, 0.03021479, 0.0297723,
  0.02505656, 0.0226255, 0.380894, 0.05350953, 0.2933379, 0.3361753, 
    0.5638272, 0.4277098, 0.5127143, 0.5444542, 0.6632278, 0.4386871, 
    0.4286199, 0.2578885, 0.2541279, 0.215197, 0.3640927, 0.2998199, 
    0.2180675, 0.1999581, 0.2023803, 0.3524405, 0.3688365, 0.3527653, 
    0.1636901, 0.2039453, 0.4282491, 0.06305875, 0.06246687,
  0.4827552, 0.4285725, 0.4072319, 0.30822, 0.3288798, 0.3795512, 0.2651968, 
    0.2144923, 0.310955, 0.2906811, 0.2337494, 0.2842383, 0.2934392, 
    0.2725927, 0.2577922, 0.2446215, 0.2958433, 0.2762636, 0.1750425, 
    0.2225945, 0.2722601, 0.1998066, 0.3248446, 0.4525406, 0.1192192, 
    0.09429353, 0.1221411, 0.2292351, 0.3569252 ;

 average_DT = 732 ;

 average_T1 = 14.5 ;

 average_T2 = 746.5 ;

 climatology_bounds =
  14.5, 746.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
