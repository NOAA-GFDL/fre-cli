netcdf atmos_level_cmip.185001-185412.cl.SECOND_TRY_W_NCKS_lat01_lon01 {
dimensions:
	lev = 49 ;
	bnds = 2 ;
	time = UNLIMITED ; // (60 currently)
	lat = 2 ;
	lon = 2 ;
variables:
	double ap(lev) ;
		ap:long_name = "vertical coordinate formula term: ap(k)" ;
		ap:units = "Pa" ;
		ap:missing_value = 1.e+20 ;
		ap:_FillValue = 1.e+20 ;
		ap:cell_methods = "time: point" ;
	double ap_bnds(lev, bnds) ;
		ap_bnds:long_name = "vertical coordinate formula term: ap(k+1/2)" ;
		ap_bnds:units = "Pa" ;
		ap_bnds:missing_value = 1.e+20 ;
		ap_bnds:_FillValue = 1.e+20 ;
		ap_bnds:cell_methods = "time: point" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	double b(lev) ;
		b:long_name = "vertical coordinate formula term: b(k)" ;
		b:units = "1.0" ;
		b:missing_value = 1.e+20 ;
		b:_FillValue = 1.e+20 ;
		b:cell_methods = "time: point" ;
	double b_bnds(lev, bnds) ;
		b_bnds:long_name = "vertical coordinate formula term: b(k+1/2)" ;
		b_bnds:units = "1.0" ;
		b_bnds:missing_value = 1.e+20 ;
		b_bnds:_FillValue = 1.e+20 ;
		b_bnds:cell_methods = "time: point" ;
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	float cl(time, lev, lat, lon) ;
		cl:long_name = "Percentage Cloud Cover" ;
		cl:units = "%" ;
		cl:missing_value = 1.e+20f ;
		cl:_FillValue = 1.e+20f ;
		cl:cell_methods = "time: mean" ;
		cl:cell_measures = "area: area" ;
		cl:time_avg_info = "average_T1,average_T2,average_DT" ;
		cl:standard_name = "cloud_area_fraction_in_atmosphere_layer" ;
		cl:interp_method = "conserve_order1" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lev(lev) ;
		lev:long_name = "hybrid sigma pressure coordinate" ;
		lev:units = "1.0" ;
		lev:axis = "Z" ;
		lev:positive = "down" ;
		lev:formula = "p(n,k,j,i) = ap(k) + b(k)*ps(n,j,i)" ;
		lev:formula_terms = "ap: ap b: b ps: ps" ;
		lev:bounds = "lev_bnds" ;
		lev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
	double lev_bnds(lev, bnds) ;
		lev_bnds:long_name = "hybrid sigma pressure coordinate" ;
		lev_bnds:units = "1.0" ;
		lev_bnds:missing_value = 1.e+20 ;
		lev_bnds:_FillValue = 1.e+20 ;
		lev_bnds:cell_methods = "time: point" ;
		lev_bnds:formula = "p(n,k+1/2,j,i) = ap(k+1/2) + b(k+1/2)*ps(n,j,i)" ;
		lev_bnds:formula_terms = "ap: ap_bnds b: b_bnds ps: ps" ;
		lev_bnds:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;

// global attributes:
		:filename = "atmos_level_cmip.185001-185412.cl.nc" ;
		:title = "ESM4_historical_D1" ;
		:associated_files = "area: 18540101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Mon Jul 21 16:30:54 2025: ncks -d lon,0,1 fre/tests/test_files/ascii_files/mock_archive/cm6/ESM4/DECK/ESM4_historical_D1/gfdl.ncrc4-intel16-prod-openmp/pp/atmos_level_cmip/ts/monthly/5yr/atmos_level_cmip.185001-185412.cl.SECOND_TRY_W_NCKS_lat01.nc fre/tests/test_files/ascii_files/mock_archive/cm6/ESM4/DECK/ESM4_historical_D1/gfdl.ncrc4-intel16-prod-openmp/pp/atmos_level_cmip/ts/monthly/5yr/atmos_level_cmip.185001-185412.cl.SECOND_TRY_W_NCKS_lat01_lon01.nc\n",
			"Mon Jul 21 16:29:56 2025: ncks -d lat,0,1 /archive/cm6/ESM4/DECK/ESM4_historical_D1/gfdl.ncrc4-intel16-prod-openmp/pp/atmos_level_cmip/ts/monthly/5yr/atmos_level_cmip.185001-185412.cl.nc fre/tests/test_files/ascii_files/mock_archive/cm6/ESM4/DECK/ESM4_historical_D1/gfdl.ncrc4-intel16-prod-openmp/pp/atmos_level_cmip/ts/monthly/5yr/atmos_level_cmip.185001-185412.cl.SECOND_TRY_W_NCKS_lat01.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 18540101.atmos_level_cmip --interp_method conserve_order2 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field ap,b,ap_bnds,b_bnds,lev_bnds,ps,cl,clw,cli,mc,pfull,phalf,tntrl,tntrs,tntrlcs,tntrscs,tntpbl,tntscp,tnhuspbl,tnhusscp,ec550aer,rsu,rsd,rsucs,rsdcs,rsuaf,rsdaf,rsucsaf,rsdcsaf,time_bnds --output_file out.nc" ;
		:code_version = "$Name: bronx-10_performance_z1l $" ;
		:external_variables = "area ps" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 ap = 5, 117.5, 421.739915, 893.90957, 1524.99281, 2319.624475, 3287.104845, 
    4440.89285, 5800.305335, 7387.967285, 9221.47223, 11308.18362, 
    13637.394975, 16168.74996, 18812.38506, 21393.82351, 23624.90421, 
    25140.26087, 25599.435575, 24747.49219, 22371.578655, 18888.51393, 
    15409.188855, 12483.56931, 10040.876315, 8016.256785, 6350.800645, 
    4991.46627, 3890.9233, 3007.32337, 2304.010415, 1749.18294, 1315.52082, 
    979.788985, 722.42975, 527.15454, 380.54455, 271.66834, 191.72284, 
    133.702575, 92.10024, 62.640445, 42.046895, 27.8422, 18.159735, 
    11.571225, 7.032955, 3.93429, 1.84861 ;

 ap_bnds =
  0, 10,
  10, 225,
  225, 618.47983,
  618.47983, 1169.33931,
  1169.33931, 1880.64631,
  1880.64631, 2758.60264,
  2758.60264, 3815.60705,
  3815.60705, 5066.17865,
  5066.17865, 6534.43202,
  6534.43202, 8241.50255,
  8241.50255, 10201.44191,
  10201.44191, 12414.92533,
  12414.92533, 14859.86462,
  14859.86462, 17477.6353,
  17477.6353, 20147.13482,
  20147.13482, 22640.5122,
  22640.5122, 24609.29622,
  24609.29622, 25671.22552,
  25671.22552, 25527.64563,
  25527.64563, 23967.33875,
  23967.33875, 20775.81856,
  20775.81856, 17001.2093,
  17001.2093, 13817.16841,
  13817.16841, 11149.97021,
  11149.97021, 8931.78242,
  8931.78242, 7100.73115,
  7100.73115, 5600.87014,
  5600.87014, 4382.0624,
  4382.0624, 3399.7842,
  3399.7842, 2614.86254,
  2614.86254, 1993.15829,
  1993.15829, 1505.20759,
  1505.20759, 1125.83405,
  1125.83405, 833.74392,
  833.74392, 611.11558,
  611.11558, 443.1935,
  443.1935, 317.8956,
  317.8956, 225.44108,
  225.44108, 158.0046,
  158.0046, 109.40055,
  109.40055, 74.79993,
  74.79993, 50.48096,
  50.48096, 33.61283,
  33.61283, 22.07157,
  22.07157, 14.2479,
  14.2479, 8.89455,
  8.89455, 5.17136,
  5.17136, 2.69722,
  2.69722, 1 ;

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 
    30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 
    396, 424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 
    820, 850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 
    1215, 1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 
    1580, 1611, 1641, 1672, 1703, 1733, 1764, 1794 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 
    424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 
    850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 1215, 
    1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 1580, 
    1611, 1641, 1672, 1703, 1733, 1764, 1794, 1825 ;

 b = 0.9979, 0.991615, 0.98119, 0.96672, 0.948075, 0.92488, 0.896675, 
    0.86289, 0.822815, 0.77563, 0.720575, 0.65702, 0.58464, 0.50363, 
    0.415085, 0.321875, 0.22958, 0.145895, 0.078055, 0.0307, 0.006265, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 b_bnds =
  1, 0.9958,
  0.9958, 0.98743,
  0.98743, 0.97495,
  0.97495, 0.95849,
  0.95849, 0.93766,
  0.93766, 0.9121,
  0.9121, 0.88125,
  0.88125, 0.84453,
  0.84453, 0.8011,
  0.8011, 0.75016,
  0.75016, 0.69099,
  0.69099, 0.62305,
  0.62305, 0.54623,
  0.54623, 0.46103,
  0.46103, 0.36914,
  0.36914, 0.27461,
  0.27461, 0.18455,
  0.18455, 0.10724,
  0.10724, 0.04887,
  0.04887, 0.01253,
  0.01253, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0 ;

 bnds = 1, 2 ;

 cl =
  27.85148, 27.85148,
  12.73434, 12.87011,
  38.67724, 38.67724,
  18.09217, 18.27705,
  55.41908, 55.41908,
  32.66186, 32.86625,
  58.72105, 58.72105,
  43.27279, 43.41153,
  55.50704, 55.50704,
  45.11281, 45.20617,
  54.92191, 54.92191,
  40.67747, 40.80541,
  54.26905, 54.26905,
  39.1628, 39.29848,
  49.87909, 49.87909,
  32.2811, 32.43915,
  40.19349, 40.19349,
  25.45548, 25.58785,
  32.5076, 32.5076,
  22.14293, 22.23602,
  27.28093, 27.28093,
  19.91741, 19.98354,
  29.98196, 29.98196,
  22.16932, 22.23949,
  25.85976, 25.85976,
  17.54006, 17.61478,
  19.52938, 19.52938,
  12.98143, 13.04024,
  17.40876, 17.40876,
  11.57389, 11.6263,
  16.32877, 16.32877,
  12.98447, 13.01451,
  12.19973, 12.19973,
  10.64583, 10.65978,
  8.309202, 8.309202,
  6.060558, 6.080754,
  3.042281, 3.042281,
  2.477646, 2.482717,
  0.1005351, 0.1005351,
  0.06708267, 0.06738311,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  33.0099, 33.0099,
  23.73979, 23.82304,
  38.41985, 38.41985,
  27.48684, 27.58503,
  51.3399, 51.3399,
  28.13884, 28.34722,
  58.64093, 58.64093,
  40.13245, 40.29868,
  54.19417, 54.19417,
  41.58451, 41.69776,
  49.21782, 49.21782,
  41.42955, 41.4995,
  44.66877, 44.66877,
  39.34883, 39.39661,
  34.44837, 34.44837,
  31.39874, 31.42612,
  27.90295, 27.90295,
  22.78058, 22.82658,
  24.11592, 24.11592,
  16.41889, 16.48802,
  18.63088, 18.63088,
  13.87077, 13.91352,
  18.91646, 18.91646,
  10.68683, 10.76074,
  19.23944, 19.23944,
  11.32769, 11.39875,
  19.33073, 19.33073,
  12.55065, 12.61155,
  18.20393, 18.20393,
  14.14947, 14.18588,
  15.71866, 15.71866,
  12.54174, 12.57027,
  11.05948, 11.05948,
  11.14073, 11.14,
  7.368762, 7.368762,
  9.441517, 9.422901,
  1.444367, 1.444367,
  5.056911, 5.024466,
  0.05909855, 0.05909855,
  0.5828446, 0.5781407,
  0, 0,
  0.0009941104, 0.000985182,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  75.95712, 75.95712,
  57.38451, 57.55131,
  78.12782, 78.12782,
  60.37099, 60.53047,
  77.48823, 77.48823,
  66.1749, 66.2765,
  73.51383, 73.51383,
  57.44607, 57.59038,
  69.02752, 69.02752,
  56.66345, 56.77449,
  67.23795, 67.23795,
  56.66991, 56.76482,
  64.79355, 64.79355,
  55.12547, 55.2123,
  58.87162, 58.87162,
  50.67424, 50.74786,
  55.58938, 55.58938,
  49.53196, 49.58636,
  56.07236, 56.07236,
  48.75732, 48.82301,
  52.25702, 52.25702,
  45.8217, 45.8795,
  47.99851, 47.99851,
  43.03007, 43.07469,
  44.53238, 44.53238,
  39.34657, 39.39314,
  41.15305, 41.15305,
  35.0128, 35.06795,
  36.58344, 36.58344,
  32.32814, 32.36636,
  33.14792, 33.14792,
  31.13007, 31.1482,
  30.99298, 30.99298,
  29.19408, 29.21023,
  30.09105, 30.09105,
  28.626, 28.63916,
  21.23617, 21.23617,
  21.29935, 21.29878,
  4.057632, 4.057632,
  3.817808, 3.819962,
  0.03776565, 0.03776565,
  0.02217093, 0.02231099,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  91.0776, 91.0776,
  67.38197, 67.59478,
  91.14924, 91.14924,
  68.77433, 68.97528,
  84.90218, 84.90218,
  61.82907, 62.03629,
  79.55137, 79.55137,
  52.23996, 52.48524,
  75.47091, 75.47091,
  48.48681, 48.72916,
  68.74878, 68.74878,
  49.53168, 49.70427,
  65.45902, 65.45902,
  45.80873, 45.98522,
  61.7374, 61.7374,
  38.22552, 38.43669,
  57.68725, 57.68725,
  36.88497, 37.0718,
  53.71977, 53.71977,
  35.69449, 35.85638,
  49.75279, 49.75279,
  32.08895, 32.24759,
  46.66859, 46.66859,
  28.84737, 29.00742,
  46.72389, 46.72389,
  28.77671, 28.9379,
  46.0657, 46.0657,
  29.85096, 29.99659,
  45.9656, 45.9656,
  30.15489, 30.29689,
  46.46061, 46.46061,
  30.88661, 31.02648,
  44.47289, 44.47289,
  30.93209, 31.0537,
  40.85146, 40.85146,
  29.02374, 29.12996,
  34.55372, 34.55372,
  25.00076, 25.08656,
  21.56639, 21.56639,
  16.60826, 16.65279,
  5.810819, 5.810819,
  3.310213, 3.332672,
  0.09695192, 0.09695192,
  0.009173589, 0.009961947,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  82.36574, 82.36574,
  57.01478, 57.24247,
  84.69451, 84.69451,
  57.38116, 57.62647,
  76.16801, 76.16801,
  60.14574, 60.28964,
  66.31133, 66.31133,
  43.25971, 43.46674,
  64.43953, 64.43953,
  39.01301, 39.24137,
  58.31358, 58.31358,
  36.56245, 36.7578,
  56.4133, 56.4133,
  36.83033, 37.00621,
  49.67712, 49.67712,
  31.18184, 31.34795,
  44.3818, 44.3818,
  27.05942, 27.215,
  38.34169, 38.34169,
  24.41472, 24.5398,
  36.66898, 36.66898,
  22.34451, 22.47316,
  33.6657, 33.6657,
  22.29036, 22.39253,
  33.75163, 33.75163,
  22.29708, 22.39995,
  33.57313, 33.57313,
  23.42899, 23.52009,
  32.49377, 32.49377,
  23.65401, 23.7334,
  33.07833, 33.07833,
  24.77794, 24.85248,
  33.32863, 33.32863,
  25.58429, 25.65385,
  29.17925, 29.17925,
  23.94832, 23.9953,
  27.01131, 27.01131,
  21.93313, 21.97874,
  24.35997, 24.35997,
  19.15182, 19.19859,
  9.268961, 9.268961,
  8.518264, 8.525005,
  0.8297518, 0.8297518,
  0.7395716, 0.7403816,
  0.000717256, 0.000717256,
  0.0005819697, 0.0005831847,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  86.18253, 86.18253,
  72.24055, 72.36578,
  85.204, 85.204,
  72.12112, 72.23862,
  78.31268, 78.31268,
  72.97943, 73.02734,
  70.92127, 70.92127,
  59.52374, 59.62611,
  70.6129, 70.6129,
  59.34283, 59.44405,
  58.85361, 58.85361,
  55.58355, 55.61292,
  56.54573, 56.54573,
  51.25243, 51.29997,
  50.67115, 50.67115,
  44.95353, 45.00488,
  43.88674, 43.88674,
  40.72234, 40.75076,
  41.65145, 41.65145,
  38.88433, 38.90919,
  36.69619, 36.69619,
  35.11242, 35.12665,
  35.58663, 35.58663,
  30.83768, 30.88033,
  33.44549, 33.44549,
  27.92631, 27.97588,
  31.41978, 31.41978,
  26.08587, 26.13377,
  28.29036, 28.29036,
  25.44368, 25.46925,
  25.30692, 25.30692,
  23.82336, 23.83669,
  23.16894, 23.16894,
  21.64002, 21.65376,
  19.31705, 19.31705,
  17.28086, 17.29915,
  13.47898, 13.47898,
  14.18256, 14.17624,
  10.13065, 10.13065,
  9.474202, 9.480098,
  6.261026, 6.261026,
  4.373269, 4.390224,
  1.946118, 1.946118,
  0.8044162, 0.8146701,
  0.07344403, 0.07344403,
  0.009772204, 0.01034406,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  83.60775, 83.60775,
  64.07918, 64.25457,
  84.62437, 84.62437,
  65.37153, 65.54444,
  75.3931, 75.3931,
  67.43545, 67.50691,
  69.94276, 69.94276,
  48.6241, 48.81556,
  63.05647, 63.05647,
  49.0743, 49.19987,
  63.76386, 63.76386,
  49.29998, 49.42989,
  54.73239, 54.73239,
  48.97493, 49.02664,
  47.16717, 47.16717,
  39.94339, 40.00827,
  43.39661, 43.39661,
  36.47509, 36.53726,
  43.6961, 43.6961,
  34.24856, 34.33341,
  41.12586, 41.12586,
  33.4893, 33.55788,
  39.41077, 39.41077,
  32.76638, 32.82605,
  36.87906, 36.87906,
  31.56076, 31.60852,
  35.27384, 35.27384,
  30.73241, 30.7732,
  34.79221, 34.79221,
  30.58564, 30.62342,
  33.1995, 33.1995,
  29.85908, 29.88908,
  26.65848, 26.65848,
  27.75535, 27.7455,
  15.77363, 15.77363,
  16.32709, 16.32211,
  16.80542, 16.80542,
  20.14971, 20.11968,
  14.64305, 14.64305,
  15.23681, 15.23148,
  13.28204, 13.28204,
  13.22374, 13.22426,
  14.30448, 14.30448,
  12.34219, 12.35981,
  7.163228, 7.163228,
  5.970452, 5.981165,
  0.3783171, 0.3783171,
  0.4046365, 0.4044002,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.8148125, 0.8148125,
  0.2531647, 0.258209,
  0.8461053, 0.8461053,
  0.1419454, 0.1482697,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  87.69922, 87.69922,
  71.08559, 71.2348,
  87.21751, 87.21751,
  67.97785, 68.15065,
  73.85736, 73.85736,
  59.5816, 59.70981,
  73.15524, 73.15524,
  48.32474, 48.54774,
  66.22725, 66.22725,
  51.8307, 51.96,
  57.73967, 57.73967,
  47.92585, 48.01399,
  51.77511, 51.77511,
  44.98016, 45.04119,
  43.65107, 43.65107,
  40.2463, 40.27688,
  37.45925, 37.45925,
  33.47801, 33.51377,
  33.27981, 33.27981,
  29.79948, 29.83074,
  29.38867, 29.38867,
  27.30948, 27.32815,
  27.15902, 27.15902,
  25.29218, 25.30895,
  26.2178, 26.2178,
  24.50603, 24.52141,
  23.64171, 23.64171,
  21.673, 21.69068,
  22.64807, 22.64807,
  20.41923, 20.43925,
  21.22153, 21.22153,
  19.24845, 19.26617,
  20.33834, 20.33834,
  17.71302, 17.7366,
  17.26342, 17.26342,
  13.26269, 13.29862,
  19.41961, 19.41961,
  16.83152, 16.85476,
  16.45845, 16.45845,
  13.49654, 13.52314,
  15.21401, 15.21401,
  11.59475, 11.62726,
  13.23087, 13.23087,
  10.41926, 10.44451,
  9.176882, 9.176882,
  8.561828, 8.567351,
  4.602982, 4.602982,
  4.570874, 4.571162,
  2.332996, 2.332996,
  1.246696, 1.256452,
  2.74172, 2.74172,
  1.240687, 1.254169,
  4.585376, 4.585376,
  2.492507, 2.511304,
  3.643159, 3.643159,
  0.8920868, 0.9167948,
  1.128492, 1.128492,
  0.2674411, 0.2751744,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  88.60856, 88.60856,
  70.87464, 71.03392,
  87.65398, 87.65398,
  71.95767, 72.09864,
  83.93428, 83.93428,
  58.46349, 58.69225,
  68.731, 68.731,
  46.06889, 46.27243,
  63.3314, 63.3314,
  39.92346, 40.13369,
  55.77443, 55.77443,
  43.026, 43.1405,
  51.08231, 51.08231,
  34.35034, 34.50061,
  42.2154, 42.2154,
  28.34123, 28.46584,
  32.75753, 32.75753,
  25.00379, 25.07343,
  27.93323, 27.93323,
  22.06142, 22.11416,
  23.02752, 23.02752,
  18.83795, 18.87558,
  20.57451, 20.57451,
  16.1633, 16.20292,
  17.17031, 17.17031,
  12.3079, 12.35157,
  15.44964, 15.44964,
  11.21398, 11.25202,
  13.86632, 13.86632,
  10.01645, 10.05103,
  12.88282, 12.88282,
  8.320961, 8.361933,
  12.32004, 12.32004,
  7.738605, 7.779752,
  10.56006, 10.56006,
  6.729684, 6.764085,
  7.87149, 7.87149,
  4.706281, 4.734708,
  9.808927, 9.808927,
  5.264897, 5.305708,
  8.959722, 8.959722,
  5.00068, 5.036238,
  6.847228, 6.847228,
  2.897586, 2.933059,
  3.12221, 3.12221,
  0.8599946, 0.8803122,
  1.665695, 1.665695,
  0.9051223, 0.9119532,
  1.889747, 1.889747,
  1.037393, 1.045049,
  1.357957, 1.357957,
  0.7005038, 0.7064086,
  0.5413536, 0.5413536,
  0.1912674, 0.1944116,
  0.05902348, 0.05902348,
  0.005229237, 0.005712376,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  60.28604, 60.28604,
  44.50106, 44.64283,
  65.13776, 65.13776,
  39.89321, 40.11994,
  56.5442, 56.5442,
  45.67058, 45.76824,
  55.19204, 55.19204,
  39.08491, 39.22957,
  50.2137, 50.2137,
  38.65057, 38.75443,
  45.30199, 45.30199,
  40.48684, 40.53009,
  39.71307, 39.71307,
  34.44616, 34.49346,
  35.36015, 35.36015,
  27.60796, 27.67759,
  31.10368, 31.10368,
  22.1196, 22.20029,
  26.0524, 26.0524,
  18.52843, 18.59601,
  25.22886, 25.22886,
  17.86715, 17.93327,
  24.68988, 24.68988,
  15.98495, 16.06313,
  22.56774, 22.56774,
  14.42622, 14.49934,
  21.05914, 21.05914,
  14.01578, 14.07904,
  19.37714, 19.37714,
  13.40715, 13.46076,
  17.94027, 17.94027,
  12.70532, 12.75234,
  15.73155, 15.73155,
  10.5796, 10.62587,
  16.04595, 16.04595,
  11.67714, 11.71638,
  13.12858, 13.12858,
  10.12949, 10.15642,
  9.314322, 9.314322,
  7.720235, 7.734551,
  3.154539, 3.154539,
  3.07175, 3.072494,
  0.4674128, 0.4674128,
  0.7032006, 0.7010829,
  0.002243446, 0.002243446,
  0.005477278, 0.005448234,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  41.04879, 41.04879,
  29.32367, 29.42898,
  50.78015, 50.78015,
  31.39756, 31.57164,
  57.30561, 57.30561,
  44.57119, 44.68556,
  65.69215, 65.69215,
  49.64815, 49.79224,
  58.33223, 58.33223,
  48.81319, 48.89869,
  53.47593, 53.47593,
  48.46997, 48.51493,
  48.00808, 48.00808,
  46.52162, 46.53497,
  44.82268, 44.82268,
  38.2453, 38.30437,
  42.58523, 42.58523,
  37.34234, 37.38943,
  42.90445, 42.90445,
  36.47087, 36.52865,
  42.01976, 42.01976,
  36.02472, 36.07856,
  41.29137, 41.29137,
  36.43649, 36.48009,
  38.5184, 38.5184,
  34.82958, 34.86271,
  38.11272, 38.11272,
  36.12147, 36.13935,
  34.52104, 34.52104,
  33.83583, 33.84199,
  33.28193, 33.28193,
  34.11216, 34.1047,
  29.0212, 29.0212,
  30.34693, 30.33502,
  22.69158, 22.69158,
  24.69324, 24.67527,
  23.33706, 23.33706,
  23.16289, 23.16446,
  16.47484, 16.47484,
  15.56931, 15.57745,
  11.68597, 11.68597,
  10.31775, 10.33004,
  3.745219, 3.745219,
  2.163064, 2.177274,
  0.06905304, 0.06905304,
  0.01437885, 0.01486989,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  18.36902, 18.36902,
  7.787469, 7.882504,
  22.42304, 22.42304,
  11.39631, 11.49534,
  34.66896, 34.66896,
  19.24629, 19.38481,
  39.09616, 39.09616,
  25.62749, 25.74845,
  35.97769, 35.97769,
  27.86979, 27.94261,
  31.89813, 31.89813,
  22.78843, 22.87025,
  30.75087, 30.75087,
  21.20797, 21.29368,
  28.67646, 28.67646,
  20.80708, 20.87776,
  26.44823, 26.44823,
  17.98232, 18.05836,
  22.96865, 22.96865,
  15.1504, 15.22062,
  23.10245, 23.10245,
  13.82704, 13.91034,
  23.55371, 23.55371,
  13.14872, 13.24217,
  23.16136, 23.16136,
  12.79831, 12.89138,
  23.30759, 23.30759,
  14.27833, 14.35943,
  21.54025, 21.54025,
  15.4502, 15.50489,
  18.45222, 18.45222,
  14.92026, 14.95198,
  13.6558, 13.6558,
  13.31536, 13.31842,
  10.65237, 10.65237,
  9.118917, 9.132689,
  4.901077, 4.901077,
  3.728601, 3.739131,
  3.060575, 3.060575,
  1.131379, 1.148705,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  33.84033, 33.84033,
  27.2863, 27.34516,
  46.56712, 46.56712,
  36.41655, 36.50772,
  58.99448, 58.99448,
  49.93821, 50.01955,
  69.31546, 69.31546,
  63.21351, 63.26831,
  68.45028, 68.45028,
  61.05843, 61.12482,
  64.75687, 64.75687,
  61.81873, 61.84512,
  58.06006, 58.06006,
  55.38262, 55.40667,
  54.4766, 54.4766,
  53.34429, 53.35446,
  49.5568, 49.5568,
  49.90364, 49.90052,
  44.10765, 44.10765,
  40.78618, 40.81601,
  38.28327, 38.28327,
  33.9332, 33.97227,
  37.51474, 37.51474,
  30.8276, 30.88766,
  35.07786, 35.07786,
  28.97018, 29.02504,
  33.70816, 33.70816,
  26.59732, 26.66118,
  30.5865, 30.5865,
  24.95137, 25.00198,
  26.53994, 26.53994,
  22.88749, 22.9203,
  21.34949, 21.34949,
  20.36502, 20.37386,
  12.75331, 12.75331,
  13.94264, 13.93196,
  9.993784, 9.993784,
  10.93214, 10.92371,
  4.374573, 4.374573,
  4.701332, 4.698397,
  0.06031336, 0.06031336,
  0.1038093, 0.1034186,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  29.65408, 29.65408,
  15.10975, 15.24038,
  34.32711, 34.32711,
  17.89237, 18.03998,
  44.65901, 44.65901,
  27.08773, 27.24554,
  47.19104, 47.19104,
  36.82177, 36.9149,
  48.41227, 48.41227,
  41.74208, 41.80199,
  43.74643, 43.74643,
  43.25352, 43.25794,
  34.85738, 34.85738,
  35.6727, 35.66537,
  30.50502, 30.50502,
  27.4644, 27.49171,
  28.0655, 28.0655,
  26.69365, 26.70597,
  24.10934, 24.10934,
  23.93903, 23.94056,
  22.9411, 22.9411,
  22.14451, 22.15166,
  20.4796, 20.4796,
  21.64696, 21.63647,
  17.33268, 17.33268,
  18.26295, 18.2546,
  16.04115, 16.04115,
  16.85567, 16.84836,
  15.2565, 15.2565,
  14.94815, 14.95092,
  14.94616, 14.94616,
  11.45837, 11.4897,
  16.35825, 16.35825,
  11.73182, 11.77337,
  7.212742, 7.212742,
  5.338599, 5.355432,
  1.403314, 1.403314,
  0.4351376, 0.4438331,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  72.69177, 72.69177,
  55.43908, 55.59403,
  75.66699, 75.66699,
  59.81784, 59.96018,
  69.40527, 69.40527,
  59.48939, 59.57844,
  67.45607, 67.45607,
  54.9846, 55.09661,
  60.85008, 60.85008,
  53.36108, 53.42834,
  59.20927, 59.20927,
  50.14109, 50.22253,
  55.69727, 55.69727,
  47.2944, 47.36987,
  49.65295, 49.65295,
  40.22675, 40.31141,
  43.43752, 43.43752,
  36.37317, 36.43661,
  42.55772, 42.55772,
  32.03513, 32.12963,
  40.16559, 40.16559,
  26.94563, 27.06436,
  38.60447, 38.60447,
  27.11471, 27.2179,
  38.28672, 38.28672,
  29.43429, 29.51379,
  37.47762, 37.47762,
  30.64664, 30.70799,
  35.8486, 35.8486,
  25.25717, 25.35229,
  35.25663, 35.25663,
  22.79612, 22.90803,
  32.52319, 32.52319,
  22.14123, 22.23447,
  28.09079, 28.09079,
  20.00234, 20.07499,
  20.40389, 20.40389,
  15.20357, 15.25028,
  5.999115, 5.999115,
  5.828499, 5.830031,
  0.01715261, 0.01715261,
  0.03539596, 0.03523212,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  80.43752, 80.43752,
  63.22637, 63.38095,
  81.38194, 81.38194,
  65.48329, 65.62608,
  73.4452, 73.4452,
  62.45115, 62.54989,
  64.45582, 64.45582,
  50.98948, 51.11042,
  56.28338, 56.28338,
  48.5307, 48.60033,
  53.64651, 53.64651,
  48.26631, 48.31463,
  50.26707, 50.26707,
  44.75055, 44.80009,
  44.29041, 44.29041,
  40.67047, 40.70298,
  41.88541, 41.88541,
  38.12044, 38.15425,
  40.88935, 40.88935,
  36.47017, 36.50986,
  39.19927, 39.19927,
  35.91332, 35.94284,
  37.03757, 37.03757,
  35.09685, 35.11428,
  37.4533, 37.4533,
  33.99301, 34.02409,
  35.74662, 35.74662,
  33.96606, 33.98205,
  32.24739, 32.24739,
  29.69457, 29.71749,
  30.55599, 30.55599,
  26.89007, 26.923,
  28.10254, 28.10254,
  21.16537, 21.22767,
  24.85092, 24.85092,
  15.9024, 15.98277,
  19.3036, 19.3036,
  10.74576, 10.82262,
  11.43656, 11.43656,
  6.16103, 6.208411,
  0.7646336, 0.7646336,
  0.4329328, 0.4359119,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  91.07148, 91.07148,
  76.38961, 76.52147,
  92.55285, 92.55285,
  78.81962, 78.94296,
  91.42081, 91.42081,
  81.82219, 81.9084,
  79.05412, 79.05412,
  64.97026, 65.09675,
  75.2737, 75.2737,
  63.89119, 63.99342,
  69.52408, 69.52408,
  62.64622, 62.708,
  65.1014, 65.1014,
  52.47869, 52.59205,
  58.40356, 58.40356,
  50.96869, 51.03547,
  58.86279, 58.86279,
  51.6371, 51.702,
  54.91489, 54.91489,
  47.15028, 47.22002,
  52.82702, 52.82702,
  42.43481, 42.52814,
  51.67241, 51.67241,
  41.12812, 41.22282,
  52.7272, 52.7272,
  40.04153, 40.15546,
  53.74435, 53.74435,
  41.21182, 41.32438,
  53.65279, 53.65279,
  42.71864, 42.81684,
  51.355, 51.355,
  44.09439, 44.1596,
  51.55342, 51.55342,
  44.57055, 44.63327,
  50.92412, 50.92412,
  42.08414, 42.16353,
  48.15841, 48.15841,
  41.4864, 41.54632,
  44.79505, 44.79505,
  38.8558, 38.90915,
  22.25142, 22.25142,
  19.19169, 19.21917,
  1.012282, 1.012282,
  0.7884501, 0.7904603,
  0.0009267638, 0.0009267638,
  8.210744e-05, 8.969351e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  91.24292, 91.24292,
  77.69407, 77.81576,
  89.26237, 89.26237,
  79.08054, 79.17198,
  89.7021, 89.7021,
  73.10731, 73.25636,
  84.26292, 84.26292,
  70.69861, 70.82043,
  81.51834, 81.51834,
  66.23811, 66.37534,
  72.15055, 72.15055,
  63.97031, 64.04379,
  66.94313, 66.94313,
  57.64417, 57.72768,
  60.84529, 60.84529,
  54.39739, 54.4553,
  57.5248, 57.5248,
  52.39037, 52.43648,
  55.30743, 55.30743,
  48.75763, 48.81646,
  51.16525, 51.16525,
  46.98395, 47.0215,
  49.09942, 49.09942,
  44.4086, 44.45073,
  47.24413, 47.24413,
  42.57239, 42.61435,
  44.82894, 44.82894,
  38.28224, 38.34104,
  38.15202, 38.15202,
  35.78122, 35.80251,
  35.09396, 35.09396,
  32.30602, 32.33106,
  34.68427, 34.68427,
  31.38581, 31.41543,
  29.14944, 29.14944,
  28.39794, 28.40469,
  29.03428, 29.03428,
  28.01397, 28.02313,
  26.18208, 26.18208,
  26.18678, 26.18673,
  17.37171, 17.37171,
  19.34364, 19.32593,
  1.854022, 1.854022,
  2.878694, 2.869491,
  0, 0,
  0.008304689, 0.008230103,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  75.21869, 75.21869,
  61.76374, 61.88459,
  76.06578, 76.06578,
  64.45177, 64.55608,
  76.47005, 76.47005,
  58.52828, 58.68941,
  72.32109, 72.32109,
  58.84317, 58.96422,
  68.48396, 68.48396,
  52.2369, 52.38282,
  63.02151, 63.02151,
  47.93088, 48.06641,
  56.77206, 56.77206,
  46.29016, 46.3843,
  53.72889, 53.72889,
  43.3747, 43.46769,
  50.589, 50.589,
  40.87509, 40.96233,
  46.96298, 46.96298,
  39.2509, 39.32016,
  48.69425, 48.69425,
  39.68483, 39.76575,
  48.20253, 48.20253,
  41.63576, 41.69474,
  47.3098, 47.3098,
  43.59694, 43.63029,
  44.75171, 44.75171,
  44.06405, 44.07022,
  39.66209, 39.66209,
  40.48475, 40.47736,
  36.52698, 36.52698,
  36.71202, 36.71035,
  39.5498, 39.5498,
  40.6244, 40.61475,
  27.93516, 27.93516,
  33.3862, 33.33725,
  20.19409, 20.19409,
  26.19165, 26.13779,
  12.88982, 12.88982,
  14.49226, 14.47787,
  10.76949, 10.76949,
  11.12687, 11.12366,
  7.541388, 7.541388,
  7.580519, 7.580168,
  4.866945, 4.866945,
  5.016397, 5.015054,
  1.943356, 1.943356,
  2.509125, 2.504044,
  0.18086, 0.18086,
  0.4784748, 0.4758019,
  0, 0,
  0.05198649, 0.05151959,
  0.01503994, 0.01503994,
  0.1526891, 0.1514529,
  0.02989021, 0.02989021,
  0.1239897, 0.1231446,
  0.01131836, 0.01131836,
  0.006866139, 0.006906126,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  84.61886, 84.61886,
  66.17895, 66.34456,
  83.3917, 83.3917,
  68.79189, 68.92302,
  76.35095, 76.35095,
  59.77974, 59.92857,
  73.62038, 73.62038,
  50.70363, 50.90945,
  65.26362, 65.26362,
  53.37563, 53.4824,
  64.34101, 64.34101,
  49.91254, 50.04212,
  58.84681, 58.84681,
  49.16481, 49.25177,
  55.9709, 55.9709,
  46.64351, 46.72728,
  50.90992, 50.90992,
  43.81835, 43.88204,
  46.80626, 46.80626,
  42.904, 42.93904,
  43.18971, 43.18971,
  40.17949, 40.20652,
  40.01971, 40.01971,
  39.28183, 39.28846,
  37.82498, 37.82498,
  36.9709, 36.97857,
  33.52654, 33.52654,
  31.98517, 31.99902,
  31.79138, 31.79138,
  30.33396, 30.34705,
  30.51748, 30.51748,
  27.50603, 27.53308,
  29.13795, 29.13795,
  24.67879, 24.71884,
  27.54419, 27.54419,
  23.5176, 23.55376,
  24.86397, 24.86397,
  20.53463, 20.57351,
  18.61643, 18.61643,
  14.0685, 14.10935,
  16.09585, 16.09585,
  10.68491, 10.7335,
  12.82015, 12.82015,
  8.25979, 8.300748,
  11.70037, 11.70037,
  6.695739, 6.740687,
  11.18384, 11.18384,
  6.107756, 6.153345,
  10.96967, 10.96967,
  4.339327, 4.398876,
  9.948685, 9.948685,
  3.549235, 3.60671,
  8.697188, 8.697188,
  2.371389, 2.428202,
  5.435771, 5.435771,
  1.116733, 1.155524,
  2.097258, 2.097258,
  0.2627517, 0.2792279,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  86.84027, 86.84027,
  76.63775, 76.72938,
  88.07008, 88.07008,
  77.97308, 78.06377,
  82.9573, 82.9573,
  73.86852, 73.95016,
  74.34325, 74.34325,
  70.27624, 70.31276,
  70.57412, 70.57412,
  64.77266, 64.82476,
  63.07999, 63.07999,
  62.28955, 62.29665,
  57.01578, 57.01578,
  59.04842, 59.03016,
  50.70815, 50.70815,
  51.90926, 51.89848,
  43.70774, 43.70774,
  48.04795, 48.00897,
  39.88729, 39.88729,
  42.22672, 42.20571,
  38.45871, 38.45871,
  37.70174, 37.70854,
  36.95009, 36.95009,
  35.53875, 35.55143,
  33.35974, 33.35974,
  33.36399, 33.36395,
  30.73524, 30.73524,
  30.53143, 30.53326,
  29.37552, 29.37552,
  28.21528, 28.22571,
  28.91315, 28.91315,
  26.66242, 26.68263,
  25.94025, 25.94025,
  24.14255, 24.1587,
  28.15064, 28.15064,
  27.14162, 27.15068,
  25.71218, 25.71218,
  24.35399, 24.36619,
  22.00871, 22.00871,
  22.55729, 22.55236,
  18.34512, 18.34512,
  18.53923, 18.53749,
  10.58983, 10.58983,
  10.48666, 10.48759,
  7.888262, 7.888262,
  7.252894, 7.2586,
  4.366797, 4.366797,
  4.693205, 4.690274,
  2.709329, 2.709329,
  1.085347, 1.099932,
  1.626017, 1.626017,
  0.3665031, 0.377815,
  0.1477631, 0.1477631,
  0.0130912, 0.01430072,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  67.47005, 67.47005,
  49.01247, 49.17824,
  70.04877, 70.04877,
  51.63755, 51.80291,
  65.77728, 65.77728,
  49.35382, 49.50132,
  63.70708, 63.70708,
  47.95997, 48.1014,
  57.88197, 57.88197,
  44.36944, 44.4908,
  55.26914, 55.26914,
  45.98282, 46.06622,
  53.84293, 53.84293,
  45.99737, 46.06783,
  50.26569, 50.26569,
  40.82062, 40.90545,
  49.06453, 49.06453,
  38.43606, 38.53152,
  48.06089, 48.06089,
  36.81169, 36.91272,
  47.60706, 47.60706,
  37.0014, 37.09665,
  47.81564, 47.81564,
  37.97055, 38.05898,
  47.98672, 47.98672,
  39.24986, 39.32833,
  45.32954, 45.32954,
  38.62781, 38.688,
  44.55975, 44.55975,
  36.929, 36.99754,
  45.75008, 45.75008,
  35.73799, 35.82792,
  43.29406, 43.29406,
  35.75914, 35.82681,
  38.65184, 38.65184,
  31.40356, 31.46866,
  34.31614, 34.31614,
  30.07471, 30.1128,
  29.02463, 29.02463,
  25.5811, 25.61203,
  21.8947, 21.8947,
  17.13733, 17.18006,
  8.692136, 8.692136,
  6.760091, 6.777443,
  0.3421859, 0.3421859,
  0.2281468, 0.229171,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  40.16953, 40.16953,
  21.79098, 21.95604,
  51.5576, 51.5576,
  27.06559, 27.28556,
  61.83241, 61.83241,
  34.63529, 34.87955,
  69.31725, 69.31725,
  42.05862, 42.30344,
  63.88956, 63.88956,
  44.22694, 44.40354,
  54.3316, 54.3316,
  40.44492, 40.56964,
  48.39622, 48.39622,
  34.31178, 34.43827,
  41.34971, 41.34971,
  30.33134, 30.4303,
  39.03883, 39.03883,
  28.27273, 28.36942,
  37.212, 37.212,
  28.06952, 28.15163,
  36.37587, 36.37587,
  27.48089, 27.56078,
  33.93891, 33.93891,
  26.24201, 26.31114,
  29.85873, 29.85873,
  26.13869, 26.1721,
  27.21823, 27.21823,
  26.05152, 26.062,
  23.69759, 23.69759,
  24.42499, 24.41846,
  19.8083, 19.8083,
  22.48247, 22.45845,
  17.75429, 17.75429,
  20.83263, 20.80498,
  15.50017, 15.50017,
  18.44424, 18.4178,
  13.13509, 13.13509,
  16.34904, 16.32018,
  10.859, 10.859,
  13.06167, 13.04189,
  5.538041, 5.538041,
  7.696838, 7.677449,
  0.5690635, 0.5690635,
  0.9084936, 0.9054451,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  17.52904, 17.52904,
  7.127599, 7.221017,
  25.60023, 25.60023,
  9.029312, 9.17814,
  30.05016, 30.05016,
  14.69126, 14.8292,
  39.57146, 39.57146,
  19.6902, 19.86875,
  30.30638, 30.30638,
  19.38338, 19.48148,
  22.48365, 22.48365,
  17.20796, 17.25534,
  17.74803, 17.74803,
  9.202535, 9.279284,
  17.52551, 17.52551,
  9.964564, 10.03247,
  21.23277, 21.23277,
  11.99004, 12.07306,
  21.29769, 21.29769,
  14.05051, 14.11559,
  22.14792, 22.14792,
  15.24981, 15.31176,
  20.44595, 20.44595,
  16.00714, 16.047,
  20.35946, 20.35946,
  16.54547, 16.57973,
  18.7437, 18.7437,
  14.90865, 14.94309,
  17.20442, 17.20442,
  14.07716, 14.10525,
  16.90276, 16.90276,
  12.57154, 12.61044,
  15.15893, 15.15893,
  12.18588, 12.21258,
  8.617671, 8.617671,
  5.566706, 5.594108,
  4.736269, 4.736269,
  4.170672, 4.175752,
  1.476027, 1.476027,
  1.930797, 1.926713,
  0.01615722, 0.01615722,
  0.03728047, 0.03709076,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  10.81064, 10.81064,
  5.867019, 5.911418,
  15.45317, 15.45317,
  8.066678, 8.133018,
  34.19195, 34.19195,
  21.32741, 21.44295,
  47.69416, 47.69416,
  27.38854, 27.57091,
  43.05161, 43.05161,
  30.16816, 30.28387,
  36.89909, 36.89909,
  27.22395, 27.31084,
  31.75538, 31.75538,
  24.45585, 24.52141,
  27.94718, 27.94718,
  19.47024, 19.54638,
  24.87759, 24.87759,
  17.33325, 17.401,
  21.75636, 21.75636,
  16.20465, 16.25451,
  18.31926, 18.31926,
  17.17071, 17.18102,
  18.79663, 18.79663,
  17.3411, 17.35417,
  20.16318, 20.16318,
  18.64443, 18.65807,
  22.92964, 22.92964,
  20.32375, 20.34715,
  21.39393, 21.39393,
  20.4346, 20.44322,
  16.2913, 16.2913,
  19.12927, 19.10378,
  12.32457, 12.32457,
  15.13138, 15.10617,
  8.22173, 8.22173,
  8.871326, 8.865492,
  0.1869356, 0.1869356,
  0.2663672, 0.2656538,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  30.028, 30.028,
  16.97302, 17.09027,
  37.61171, 37.61171,
  20.13409, 20.29106,
  52.79651, 52.79651,
  32.60755, 32.78887,
  62.39805, 62.39805,
  38.72001, 38.93267,
  60.14057, 60.14057,
  36.83656, 37.04585,
  49.11794, 49.11794,
  37.42228, 37.52732,
  40.28808, 40.28808,
  30.56243, 30.64978,
  34.61011, 34.61011,
  26.02754, 26.10462,
  31.24658, 31.24658,
  23.89301, 23.95905,
  29.61551, 29.61551,
  23.04136, 23.1004,
  26.3269, 26.3269,
  21.88353, 21.92343,
  23.12608, 23.12608,
  19.90937, 19.93826,
  20.14623, 20.14623,
  17.96568, 17.98526,
  17.83187, 17.83187,
  17.21615, 17.22168,
  16.50222, 16.50222,
  16.06968, 16.07356,
  14.86554, 14.86554,
  14.45632, 14.45999,
  14.7194, 14.7194,
  13.5628, 13.57319,
  13.01081, 13.01081,
  12.48756, 12.49226,
  6.546091, 6.546091,
  6.90749, 6.904244,
  0.4843011, 0.4843011,
  0.2562916, 0.2583394,
  0.000726262, 0.000726262,
  6.434382e-05, 7.028866e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  76.18258, 76.18258,
  55.792, 55.97514,
  79.70839, 79.70839,
  59.88235, 60.06041,
  82.34193, 82.34193,
  55.62024, 55.86024,
  77.06115, 77.06115,
  56.37587, 56.56165,
  74.77445, 74.77445,
  53.48367, 53.67488,
  63.2865, 63.2865,
  50.11274, 50.23106,
  57.58793, 57.58793,
  42.73286, 42.86628,
  53.27625, 53.27625,
  40.10105, 40.21938,
  50.69118, 50.69118,
  37.11646, 37.23838,
  46.68024, 46.68024,
  34.02298, 34.13666,
  41.46693, 41.46693,
  30.91038, 31.00519,
  38.30272, 38.30272,
  27.51413, 27.61102,
  36.21748, 36.21748,
  26.76281, 26.84773,
  31.04323, 31.04323,
  22.99087, 23.06319,
  28.90704, 28.90704,
  19.93822, 20.01877,
  28.70416, 28.70416,
  19.43212, 19.5154,
  28.73874, 28.73874,
  18.80142, 18.89067,
  27.27501, 27.27501,
  18.26928, 18.35016,
  20.23475, 20.23475,
  13.53599, 13.59615,
  2.39466, 2.39466,
  0.8321598, 0.846193,
  0.02810951, 0.02810951,
  0.003604388, 0.003824475,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  79.54731, 79.54731,
  62.45577, 62.60927,
  84.77292, 84.77292,
  64.0456, 64.23176,
  75.25787, 75.25787,
  65.35848, 65.44739,
  68.76734, 68.76734,
  54.44142, 54.57008,
  67.16058, 67.16058,
  59.74152, 59.80816,
  64.36774, 64.36774,
  59.26051, 59.30638,
  58.24414, 58.24414,
  56.89751, 56.9096,
  52.97651, 52.97651,
  47.0073, 47.06091,
  48.39702, 48.39702,
  44.56824, 44.60262,
  41.63731, 41.63731,
  37.82932, 37.86352,
  43.94361, 43.94361,
  38.007, 38.06032,
  39.38363, 39.38363,
  34.56459, 34.60787,
  37.64906, 37.64906,
  33.70855, 33.74394,
  33.83582, 33.83582,
  30.29144, 30.32327,
  30.44156, 30.44156,
  26.42394, 26.46002,
  28.70564, 28.70564,
  24.40618, 24.44479,
  24.60176, 24.60176,
  23.04972, 23.06366,
  16.00137, 16.00137,
  18.03611, 18.01783,
  5.537753, 5.537753,
  7.09766, 7.08365,
  0.1397303, 0.1397303,
  0.2325259, 0.2316925,
  3.18525e-05, 3.18525e-05,
  4.623621e-05, 4.610703e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  88.63386, 88.63386,
  75.69227, 75.8085,
  89.34067, 89.34067,
  77.66756, 77.77241,
  81.54593, 81.54593,
  74.54582, 74.6087,
  74.88578, 74.88578,
  59.99479, 60.12853,
  70.72366, 70.72366,
  60.78084, 60.87014,
  65.50259, 65.50259,
  63.40592, 63.42475,
  62.7384, 62.7384,
  57.83884, 57.88285,
  56.95292, 56.95292,
  52.11766, 52.16109,
  48.54087, 48.54087,
  45.18047, 45.21065,
  42.89141, 42.89141,
  37.44188, 37.49082,
  35.96813, 35.96813,
  31.49961, 31.53974,
  31.24824, 31.24824,
  27.81101, 27.84188,
  29.5803, 29.5803,
  25.16737, 25.207,
  29.38462, 29.38462,
  23.45258, 23.50585,
  27.21396, 27.21396,
  22.39841, 22.44166,
  21.79621, 21.79621,
  20.38035, 20.39306,
  22.46325, 22.46325,
  20.30913, 20.32847,
  18.36586, 18.36586,
  18.57017, 18.56833,
  15.98176, 15.98176,
  14.39044, 14.40473,
  11.24217, 11.24217,
  10.92882, 10.93163,
  4.068458, 4.068458,
  4.627243, 4.622224,
  0.08648864, 0.08648864,
  0.2035335, 0.2024823,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  86.62928, 86.62928,
  65.73692, 65.92457,
  84.08295, 84.08295,
  67.79131, 67.93762,
  71.91749, 71.91749,
  62.47082, 62.55566,
  65.26395, 65.26395,
  47.68043, 47.83835,
  54.45742, 54.45742,
  47.29594, 47.36025,
  48.22163, 48.22163,
  42.21669, 42.27062,
  42.34187, 42.34187,
  36.63821, 36.68943,
  35.19902, 35.19902,
  29.7449, 29.79388,
  27.87762, 27.87762,
  26.35059, 26.36431,
  24.53527, 24.53527,
  22.29431, 22.31443,
  21.07539, 21.07539,
  20.97315, 20.97407,
  18.79482, 18.79482,
  17.29833, 17.31177,
  16.10358, 16.10358,
  12.63207, 12.66325,
  14.56567, 14.56567,
  9.823259, 9.865851,
  15.09603, 15.09603,
  9.746312, 9.794359,
  15.53017, 15.53017,
  9.833385, 9.884549,
  15.80779, 15.80779,
  10.97083, 11.01427,
  19.61478, 19.61478,
  12.79227, 12.85355,
  13.5673, 13.5673,
  10.61241, 10.63895,
  9.250558, 9.250558,
  6.304818, 6.331274,
  1.825499, 1.825499,
  1.137465, 1.143645,
  0.03778417, 0.03778417,
  0.005461728, 0.005752024,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  82.25242, 82.25242,
  68.12205, 68.24895,
  81.41699, 81.41699,
  70.00395, 70.10646,
  83.69369, 83.69369,
  65.93298, 66.09249,
  68.71919, 68.71919,
  64.47299, 64.51113,
  68.96155, 68.96155,
  53.13868, 53.28079,
  61.53284, 61.53284,
  53.98596, 54.05374,
  57.74524, 57.74524,
  51.33428, 51.39186,
  46.1486, 46.1486,
  43.88787, 43.90818,
  40.03127, 40.03127,
  40.56861, 40.56379,
  35.70294, 35.70294,
  36.5998, 36.59175,
  32.25544, 32.25544,
  33.61382, 33.60162,
  30.84151, 30.84151,
  31.83216, 31.82326,
  27.20778, 27.20778,
  30.10418, 30.07817,
  24.70153, 24.70153,
  27.3058, 27.28241,
  24.37851, 24.37851,
  25.29958, 25.29131,
  23.68178, 23.68178,
  22.85977, 22.86716,
  22.38335, 22.38335,
  21.20689, 21.21746,
  21.50411, 21.50411,
  20.29176, 20.30265,
  20.50905, 20.50905,
  20.25431, 20.2566,
  17.5701, 17.5701,
  16.58217, 16.59105,
  15.73302, 15.73302,
  14.7588, 14.76755,
  8.764238, 8.764238,
  8.18434, 8.189548,
  1.657494, 1.657494,
  1.832403, 1.830832,
  0.01736214, 0.01736214,
  0.02609199, 0.02601358,
  0, 0,
  0, 0,
  0, 0,
  0.009173715, 0.009091323,
  0.08719734, 0.08719734,
  0.3586452, 0.3562073,
  0.7842461, 0.7842461,
  1.010594, 1.008561,
  0.06510743, 0.06510743,
  0.1725552, 0.1715902,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  81.30362, 81.30362,
  55.85831, 56.08684,
  79.80363, 79.80363,
  58.63059, 58.82075,
  74.79266, 74.79266,
  54.01315, 54.19978,
  63.16971, 63.16971,
  52.1753, 52.27405,
  55.88431, 55.88431,
  39.69559, 39.84098,
  48.80812, 48.80812,
  44.00201, 44.04518,
  42.19798, 42.19798,
  41.20203, 41.21098,
  33.65993, 33.65993,
  29.86595, 29.90003,
  28.99355, 28.99355,
  24.69155, 24.73018,
  26.87388, 26.87388,
  23.61724, 23.64649,
  26.99927, 26.99927,
  23.56284, 23.5937,
  26.88212, 26.88212,
  23.14068, 23.17428,
  26.07437, 26.07437,
  22.78506, 22.8146,
  26.44845, 26.44845,
  23.3922, 23.41965,
  24.30231, 24.30231,
  22.60077, 22.61606,
  22.60131, 22.60131,
  20.36318, 20.38329,
  17.45304, 17.45304,
  16.96045, 16.96488,
  10.80139, 10.80139,
  12.09931, 12.08765,
  6.485567, 6.485567,
  7.513194, 7.503964,
  4.352758, 4.352758,
  4.167194, 4.16886,
  3.379382, 3.379382,
  2.03993, 2.05196,
  0.9859016, 0.9859016,
  0.3453183, 0.3510715,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0487478, 0.0487478,
  0.005476018, 0.005864653,
  0.1600363, 0.1600363,
  0.02159171, 0.02283512,
  0.01516616, 0.01516616,
  0.001343659, 0.001467803,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  89.06666, 89.06666,
  58.31568, 58.59186,
  86.85265, 86.85265,
  59.7725, 60.01572,
  73.05346, 73.05346,
  63.21812, 63.30645,
  62.15367, 62.15367,
  35.00862, 35.25242,
  53.51307, 53.51307,
  36.57105, 36.72321,
  44.27382, 44.27382,
  33.88681, 33.98009,
  40.18012, 40.18012,
  31.34474, 31.42409,
  35.1348, 35.1348,
  26.13741, 26.21821,
  32.95485, 32.95485,
  24.7568, 24.83043,
  26.28286, 26.28286,
  22.52315, 22.55692,
  22.81212, 22.81212,
  18.77444, 18.81071,
  22.24076, 22.24076,
  18.06356, 18.10108,
  22.06899, 22.06899,
  15.79049, 15.84688,
  21.30525, 21.30525,
  15.75172, 15.8016,
  20.72294, 20.72294,
  15.34273, 15.39105,
  18.08024, 18.08024,
  13.516, 13.55699,
  16.75351, 16.75351,
  11.98464, 12.02747,
  13.77077, 13.77077,
  9.787292, 9.823069,
  10.95989, 10.95989,
  7.121408, 7.155882,
  7.369947, 7.369947,
  3.62472, 3.658357,
  5.257377, 5.257377,
  3.179593, 3.198254,
  3.216109, 3.216109,
  2.984017, 2.986102,
  2.609965, 2.609965,
  3.14715, 3.142326,
  2.5467, 2.5467,
  1.409359, 1.419573,
  0.1321896, 0.1321896,
  0.0532343, 0.05394341,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  79.91679, 79.91679,
  55.38636, 55.60668,
  80.86201, 80.86201,
  58.49819, 58.69904,
  77.20976, 77.20976,
  50.37524, 50.61625,
  69.98296, 69.98296,
  53.05875, 53.21075,
  64.14995, 64.14995,
  45.56811, 45.735,
  64.24861, 64.24861,
  46.34573, 46.50652,
  61.20833, 61.20833,
  44.50655, 44.65655,
  58.62381, 58.62381,
  40.12804, 40.29416,
  52.97514, 52.97514,
  37.18856, 37.33034,
  45.37001, 45.37001,
  33.69802, 33.80285,
  39.91879, 39.91879,
  30.04397, 30.13266,
  39.96268, 39.96268,
  29.11174, 29.20919,
  36.33958, 36.33958,
  26.80166, 26.88732,
  35.49271, 35.49271,
  25.98291, 26.06832,
  35.08326, 35.08326,
  25.48951, 25.57568,
  33.45935, 33.45935,
  25.0409, 25.1165,
  31.22209, 31.22209,
  24.23234, 24.29511,
  27.78898, 27.78898,
  22.0968, 22.14792,
  23.04955, 23.04955,
  18.23051, 18.27379,
  20.32435, 20.32435,
  13.8912, 13.94897,
  16.31941, 16.31941,
  8.684522, 8.753093,
  6.754183, 6.754183,
  3.601439, 3.629755,
  0.3241685, 0.3241685,
  0.2059964, 0.2070577,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  33.62373, 33.62373,
  17.49222, 17.6371,
  38.73801, 38.73801,
  21.24877, 21.40584,
  37.94302, 37.94302,
  25.08826, 25.20371,
  37.39295, 37.39295,
  26.52502, 26.62263,
  35.2679, 35.2679,
  26.46796, 26.547,
  32.18398, 32.18398,
  23.13135, 23.21265,
  32.55042, 32.55042,
  21.17723, 21.27937,
  32.60008, 32.60008,
  22.13146, 22.22548,
  30.79644, 30.79644,
  21.52221, 21.6055,
  30.93982, 30.93982,
  20.75346, 20.84495,
  27.78126, 27.78126,
  18.77025, 18.85118,
  26.63289, 26.63289,
  18.67578, 18.74724,
  25.11158, 25.11158,
  18.22897, 18.29079,
  24.63388, 24.63388,
  18.79956, 18.85196,
  24.25712, 24.25712,
  19.39597, 19.43962,
  23.10967, 23.10967,
  19.07997, 19.11616,
  21.96367, 21.96367,
  18.61431, 18.64439,
  20.47152, 20.47152,
  17.38178, 17.40953,
  16.72561, 16.72561,
  14.24363, 14.26592,
  8.5326, 8.5326,
  8.239841, 8.242471,
  2.900849, 2.900849,
  3.059468, 3.058043,
  0.07384977, 0.07384977,
  0.06864223, 0.068689,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  5.966227, 5.966227,
  1.371689, 1.412954,
  9.262882, 9.262882,
  2.551268, 2.611547,
  18.1924, 18.1924,
  10.30554, 10.37637,
  25.7967, 25.7967,
  9.216871, 9.365779,
  24.17033, 24.17033,
  15.84277, 15.91756,
  23.12196, 23.12196,
  17.53243, 17.58263,
  23.01181, 23.01181,
  15.48402, 15.55163,
  16.80652, 16.80652,
  7.988311, 8.06751,
  11.12956, 11.12956,
  6.251781, 6.29559,
  8.170634, 8.170634,
  3.128414, 3.1737,
  7.095222, 7.095222,
  1.968541, 2.014585,
  6.031737, 6.031737,
  1.664112, 1.703339,
  7.229155, 7.229155,
  2.906313, 2.945138,
  4.807169, 4.807169,
  2.595167, 2.615034,
  3.718016, 3.718016,
  2.341126, 2.353493,
  2.748447, 2.748447,
  1.719498, 1.728739,
  1.18523, 1.18523,
  0.6926696, 0.6970934,
  0.3559631, 0.3559631,
  0.05273092, 0.05545432,
  0.006463509, 0.006463509,
  0.0005726402, 0.0006255475,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  23.22158, 23.22158,
  15.70272, 15.77025,
  32.62326, 32.62326,
  22.51619, 22.60697,
  48.68129, 48.68129,
  35.03176, 35.15435,
  54.85059, 54.85059,
  40.39695, 40.52677,
  56.29134, 56.29134,
  46.24766, 46.33786,
  50.72787, 50.72787,
  41.40687, 41.49058,
  41.53741, 41.53741,
  32.79535, 32.87386,
  37.59119, 37.59119,
  30.20838, 30.27468,
  31.91895, 31.91895,
  28.95024, 28.9769,
  32.91797, 32.91797,
  29.11134, 29.14552,
  33.80388, 33.80388,
  30.58267, 30.6116,
  33.64843, 33.64843,
  32.05956, 32.07383,
  27.61408, 27.61408,
  29.05504, 29.0421,
  25.85921, 25.85921,
  29.62929, 29.59543,
  25.50407, 25.50407,
  28.20168, 28.17745,
  26.18268, 26.18268,
  28.48476, 28.46408,
  21.89878, 21.89878,
  23.22819, 23.21626,
  17.15549, 17.15549,
  19.4968, 19.47577,
  8.820042, 8.820042,
  8.945402, 8.944276,
  0.1518927, 0.1518927,
  0.1773327, 0.1771042,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  38.64006, 38.64006,
  19.92671, 20.09478,
  41.74013, 41.74013,
  19.59987, 19.79872,
  50.46775, 50.46775,
  25.52979, 25.75377,
  58.68349, 58.68349,
  30.02803, 30.28539,
  53.60434, 53.60434,
  36.46402, 36.61795,
  55.2436, 55.2436,
  35.72738, 35.90266,
  46.4294, 46.4294,
  33.59615, 33.71141,
  37.90416, 37.90416,
  22.68382, 22.82051,
  39.71423, 39.71423,
  23.6056, 23.75027,
  41.19454, 41.19454,
  24.58506, 24.73423,
  39.3755, 39.3755,
  26.17235, 26.29094,
  39.18819, 39.18819,
  30.07731, 30.15914,
  36.0661, 36.0661,
  30.66088, 30.70943,
  35.76655, 35.76655,
  31.20955, 31.25048,
  33.90644, 33.90644,
  29.42942, 29.46963,
  29.54941, 29.54941,
  27.30506, 27.32521,
  28.73625, 28.73625,
  25.20052, 25.23228,
  25.85544, 25.85544,
  24.28, 24.29415,
  17.84716, 17.84716,
  16.78932, 16.79882,
  5.026426, 5.026426,
  5.810385, 5.803344,
  0.2105996, 0.2105996,
  0.2533927, 0.2530084,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  79.24601, 79.24601,
  57.79538, 57.98804,
  80.13828, 80.13828,
  60.29278, 60.47102,
  71.92309, 71.92309,
  61.51707, 61.61053,
  70.8017, 70.8017,
  54.70915, 54.85368,
  71.30772, 71.30772,
  55.41657, 55.55929,
  67.68161, 67.68161,
  52.92781, 53.06032,
  65.96368, 65.96368,
  53.37241, 53.48549,
  63.02182, 63.02182,
  49.53392, 49.65506,
  57.71815, 57.71815,
  47.82159, 47.91048,
  56.73235, 56.73235,
  46.35308, 46.4463,
  56.59931, 56.59931,
  45.34956, 45.45059,
  53.62693, 53.62693,
  43.42262, 43.51426,
  51.66898, 51.66898,
  42.19343, 42.27853,
  50.97385, 50.97385,
  40.47538, 40.56967,
  49.23113, 49.23113,
  39.55446, 39.64137,
  48.46596, 48.46596,
  39.60046, 39.68008,
  43.52379, 43.52379,
  36.95488, 37.01387,
  33.31086, 33.31086,
  27.82812, 27.87737,
  19.21383, 19.21383,
  12.41443, 12.4755,
  3.550111, 3.550111,
  3.176987, 3.180338,
  0.01524834, 0.01524834,
  0.0617557, 0.06133801,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  82.98531, 82.98531,
  56.51059, 56.74836,
  83.43565, 83.43565,
  60.13165, 60.34095,
  72.18361, 72.18361,
  52.24447, 52.42355,
  66.66711, 66.66711,
  44.38539, 44.58551,
  54.19216, 54.19216,
  41.2583, 41.37446,
  49.55851, 49.55851,
  40.22667, 40.31048,
  46.75474, 46.75474,
  39.98617, 40.04696,
  45.01972, 45.01972,
  36.68518, 36.76003,
  47.07398, 47.07398,
  35.99305, 36.09257,
  50.94254, 50.94254,
  36.48938, 36.61919,
  53.37182, 53.37182,
  38.25715, 38.3929,
  58.64065, 58.64065,
  41.63197, 41.78473,
  63.17636, 63.17636,
  46.49513, 46.64495,
  67.88692, 67.88692,
  55.36922, 55.48165,
  70.39029, 70.39029,
  59.29605, 59.39569,
  72.55582, 72.55582,
  62.79049, 62.8782,
  71.87102, 71.87102,
  65.6245, 65.6806,
  70.98444, 70.98444,
  67.16101, 67.19535,
  60.29814, 60.29814,
  61.28705, 61.27817,
  44.52695, 44.52695,
  47.5003, 47.47359,
  7.470063, 7.470063,
  9.498391, 9.480175,
  0.3658519, 0.3658519,
  0.3793402, 0.3792191,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  86.37715, 86.37715,
  74.68766, 74.79265,
  85.74915, 85.74915,
  76.72147, 76.80254,
  80.18251, 80.18251,
  68.57805, 68.68227,
  76.13127, 76.13127,
  63.38472, 63.4992,
  73.64953, 73.64953,
  63.41899, 63.51088,
  66.72651, 66.72651,
  63.04871, 63.08175,
  61.82658, 61.82658,
  61.77855, 61.77898,
  57.29843, 57.29843,
  54.61814, 54.64221,
  53.03938, 53.03938,
  50.65366, 50.67509,
  52.66277, 52.66277,
  43.8299, 43.90923,
  50.35103, 50.35103,
  40.63107, 40.71837,
  47.81311, 47.81311,
  38.60198, 38.6847,
  46.84927, 46.84927,
  37.13326, 37.22052,
  45.30422, 45.30422,
  37.83006, 37.89719,
  43.73293, 43.73293,
  37.83511, 37.88808,
  42.87513, 42.87513,
  37.53225, 37.58024,
  36.46911, 36.46911,
  33.95288, 33.97548,
  37.22033, 37.22033,
  33.95038, 33.97975,
  33.62799, 33.62799,
  30.03415, 30.06642,
  32.04847, 32.04847,
  24.62745, 24.6941,
  22.74569, 22.74569,
  16.08619, 16.14601,
  1.812045, 1.812045,
  2.071178, 2.068851,
  0.002842642, 0.002842642,
  0.008052452, 0.008005661,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  91.08011, 91.08011,
  81.60759, 81.69267,
  92.49055, 92.49055,
  82.55821, 82.64742,
  87.23602, 87.23602,
  83.98425, 84.01346,
  87.65124, 87.65124,
  74.73445, 74.85046,
  88.59489, 88.59489,
  78.76695, 78.85522,
  83.46328, 83.46328,
  80.65579, 80.68101,
  80.66483, 80.66483,
  77.02431, 77.05701,
  75.53438, 75.53438,
  69.19285, 69.2498,
  69.49114, 69.49114,
  63.08727, 63.14479,
  62.99983, 62.99983,
  58.28503, 58.32737,
  59.56868, 59.56868,
  57.01996, 57.04285,
  59.82357, 59.82357,
  58.48628, 58.49829,
  57.04403, 57.04403,
  54.8001, 54.82025,
  54.78952, 54.78952,
  52.70399, 52.72273,
  51.26512, 51.26512,
  49.23371, 49.25196,
  43.18177, 43.18177,
  41.70538, 41.71864,
  43.20277, 43.20277,
  43.85312, 43.84727,
  39.99153, 39.99153,
  41.62403, 41.60936,
  33.4043, 33.4043,
  34.7673, 34.75506,
  32.01302, 32.01302,
  33.29556, 33.28405,
  29.19212, 29.19212,
  30.48406, 30.47246,
  21.21286, 21.21286,
  21.37792, 21.37644,
  5.876729, 5.876729,
  5.733111, 5.734401,
  0.4897031, 0.4897031,
  0.2256521, 0.2280236,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  81.93231, 81.93231,
  46.8837, 47.19848,
  79.13785, 79.13785,
  48.64889, 48.92272,
  67.50829, 67.50829,
  49.4568, 49.61893,
  50.57817, 50.57817,
  39.46181, 39.56165,
  42.74279, 42.74279,
  27.65261, 27.78814,
  40.10505, 40.10505,
  27.16477, 27.28099,
  35.04682, 35.04682,
  25.51322, 25.59884,
  33.321, 33.321,
  23.77823, 23.86394,
  29.83331, 29.83331,
  22.36566, 22.43273,
  27.21341, 27.21341,
  20.03868, 20.10312,
  26.75628, 26.75628,
  19.18929, 19.25725,
  26.57255, 26.57255,
  18.78698, 18.8569,
  26.65866, 26.65866,
  18.60005, 18.67243,
  26.9758, 26.9758,
  18.51313, 18.58913,
  26.8036, 26.8036,
  18.10427, 18.1824,
  22.41191, 22.41191,
  13.34075, 13.42222,
  24.31982, 24.31982,
  17.30991, 17.37287,
  20.99974, 20.99974,
  14.79717, 14.85288,
  16.38126, 16.38126,
  13.05725, 13.08711,
  11.71942, 11.71942,
  10.72891, 10.73781,
  8.019305, 8.019305,
  8.036815, 8.036657,
  7.411441, 7.411441,
  5.82711, 5.84134,
  5.549763, 5.549763,
  2.497121, 2.524537,
  4.639157, 4.639157,
  2.43635, 2.456134,
  4.362528, 4.362528,
  3.069443, 3.081057,
  5.927238, 5.927238,
  4.330632, 4.344972,
  6.956077, 6.956077,
  3.606621, 3.636703,
  6.01419, 6.01419,
  2.190705, 2.225044,
  1.046177, 1.046177,
  0.1962575, 0.2038908,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  89.53651, 89.53651,
  75.57757, 75.70294,
  87.93845, 87.93845,
  75.87868, 75.98698,
  84.4379, 84.4379,
  71.63428, 71.74928,
  80.86108, 80.86108,
  69.10352, 69.20912,
  75.52479, 75.52479,
  64.11156, 64.21407,
  69.31435, 69.31435,
  62.12513, 62.1897,
  63.49043, 63.49043,
  56.38983, 56.45361,
  59.41845, 59.41845,
  55.17508, 55.21318,
  54.47862, 54.47862,
  51.89628, 51.91947,
  52.8354, 52.8354,
  50.92566, 50.94281,
  51.27205, 51.27205,
  48.73533, 48.75811,
  51.36393, 51.36393,
  47.23969, 47.27673,
  48.74008, 48.74008,
  44.45314, 44.49164,
  45.41788, 45.41788,
  42.73772, 42.76179,
  41.38969, 41.38969,
  40.89532, 40.89976,
  38.1203, 38.1203,
  38.05639, 38.05696,
  36.7743, 36.7743,
  35.57874, 35.58948,
  34.46813, 34.46813,
  33.41225, 33.42173,
  39.00342, 39.00342,
  38.06905, 38.07744,
  36.49532, 36.49532,
  35.56026, 35.56865,
  36.87576, 36.87576,
  36.36149, 36.36611,
  32.75834, 32.75834,
  31.27015, 31.28352,
  28.98593, 28.98593,
  28.82929, 28.83069,
  24.28461, 24.28461,
  20.82015, 20.85127,
  23.50908, 23.50908,
  19.00391, 19.04437,
  21.93133, 21.93133,
  16.16083, 16.21265,
  19.64911, 19.64911,
  11.74323, 11.81423,
  15.55542, 15.55542,
  7.670301, 7.741119,
  5.641857, 5.641857,
  2.189613, 2.220618,
  0.003149982, 0.003149982,
  0.0002790754, 0.0003048597,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  92.88332, 92.88332,
  84.91631, 84.98786,
  92.28134, 92.28134,
  85.93388, 85.99088,
  91.74674, 91.74674,
  79.11253, 79.226,
  91.51745, 91.51745,
  82.95531, 83.03222,
  89.71323, 89.71323,
  80.71497, 80.79579,
  84.17126, 84.17126,
  76.66644, 76.73384,
  80.66576, 80.66576,
  72.57384, 72.64652,
  74.03139, 74.03139,
  71.2684, 71.29322,
  68.72276, 68.72276,
  65.16676, 65.19869,
  64.70107, 64.70107,
  60.00916, 60.0513,
  60.02988, 60.02988,
  58.864, 58.87447,
  56.41476, 56.41476,
  56.43779, 56.43758,
  52.404, 52.404,
  54.47493, 54.45633,
  49.1163, 49.1163,
  50.60777, 50.59437,
  44.90831, 44.90831,
  47.79296, 47.76705,
  40.15885, 40.15885,
  42.57464, 42.55294,
  32.73796, 32.73796,
  35.91246, 35.88395,
  27.95528, 27.95528,
  33.22482, 33.17749,
  26.04338, 26.04338,
  31.10746, 31.06198,
  23.80121, 23.80121,
  27.54609, 27.51246,
  17.92188, 17.92188,
  19.2907, 19.27841,
  9.065582, 9.065582,
  11.26693, 11.24716,
  4.833261, 4.833261,
  5.166615, 5.163621,
  2.102767, 2.102767,
  1.833233, 1.835653,
  0.7490259, 0.7490259,
  0.5905836, 0.5920066,
  0.2657282, 0.2657282,
  0.05110688, 0.05303444,
  0.1847846, 0.1847846,
  0.02078627, 0.02225918,
  0.1135055, 0.1135055,
  0.01005612, 0.01098522,
  0.0188782, 0.0188782,
  0.00167253, 0.001827059,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  67.64062, 67.64062,
  43.92253, 44.13555,
  73.49737, 73.49737,
  47.19931, 47.4355,
  58.58291, 58.58291,
  42.60692, 42.7504,
  50.37034, 50.37034,
  31.82479, 31.99135,
  46.17822, 46.17822,
  31.6362, 31.76681,
  42.48708, 42.48708,
  29.92547, 30.03829,
  38.80738, 38.80738,
  24.56724, 24.69514,
  32.52196, 32.52196,
  22.42224, 22.51295,
  32.20818, 32.20818,
  21.05396, 21.15414,
  32.24512, 32.24512,
  23.17947, 23.26089,
  30.02928, 30.02928,
  28.81191, 28.82284,
  26.85967, 26.85967,
  28.31903, 28.30593,
  25.48123, 25.48123,
  24.56207, 24.57033,
  21.82909, 21.82909,
  21.54375, 21.54631,
  20.64343, 20.64343,
  18.3887, 18.40895,
  20.26807, 20.26807,
  17.40103, 17.42678,
  19.42604, 19.42604,
  15.91812, 15.94963,
  18.2561, 18.2561,
  13.86737, 13.90679,
  16.31524, 16.31524,
  12.04527, 12.08362,
  10.53387, 10.53387,
  5.798255, 5.840786,
  7.927471, 7.927471,
  2.696069, 2.743054,
  5.004031, 5.004031,
  1.299726, 1.332995,
  0.8532029, 0.8532029,
  0.4299779, 0.433779,
  0.01034765, 0.01034765,
  0.003009786, 0.003075689,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  37.38588, 37.38588,
  23.07253, 23.20108,
  42.64875, 42.64875,
  25.912, 26.06232,
  48.06854, 48.06854,
  25.95955, 26.15812,
  48.9556, 48.9556,
  33.47476, 33.6138,
  49.77634, 49.77634,
  33.09949, 33.24927,
  47.407, 47.407,
  34.22712, 34.34549,
  38.2331, 38.2331,
  29.60768, 29.68515,
  34.43695, 34.43695,
  25.6662, 25.74497,
  33.27904, 33.27904,
  24.95403, 25.0288,
  30.66352, 30.66352,
  24.58885, 24.64341,
  30.17347, 30.17347,
  23.50724, 23.56711,
  29.82155, 29.82155,
  22.82473, 22.88757,
  31.01112, 31.01112,
  21.8663, 21.94843,
  32.16736, 32.16736,
  21.42139, 21.5179,
  32.41002, 32.41002,
  20.81855, 20.92265,
  32.62226, 32.62226,
  19.5011, 19.61895,
  32.06128, 32.06128,
  21.68447, 21.77767,
  27.46659, 27.46659,
  20.76477, 20.82496,
  19.37686, 19.37686,
  15.92974, 15.9607,
  11.02466, 11.02466,
  12.32843, 12.31672,
  1.48027, 1.48027,
  2.966478, 2.95313,
  0.0008728448, 0.0008728448,
  0.03587349, 0.03555914,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  13.3155, 13.3155,
  6.520794, 6.581819,
  20.50767, 20.50767,
  9.103213, 9.205639,
  24.96583, 24.96583,
  13.56547, 13.66786,
  31.26238, 31.26238,
  16.33848, 16.47252,
  27.35124, 27.35124,
  17.58262, 17.67035,
  25.00159, 25.00159,
  15.80691, 15.88949,
  22.43082, 22.43082,
  14.16291, 14.23717,
  22.07308, 22.07308,
  14.16936, 14.24035,
  23.10789, 23.10789,
  15.54108, 15.60904,
  24.12961, 24.12961,
  14.653, 14.73811,
  21.36971, 21.36971,
  17.95808, 17.98872,
  17.94203, 17.94203,
  16.48577, 16.49885,
  18.03988, 18.03988,
  15.87168, 15.89115,
  16.70758, 16.70758,
  15.25877, 15.27179,
  17.67567, 17.67567,
  14.78924, 14.81517,
  17.5211, 17.5211,
  15.73663, 15.75266,
  14.88671, 14.88671,
  14.92414, 14.9238,
  11.73866, 11.73866,
  12.40322, 12.39725,
  5.053337, 5.053337,
  6.659327, 6.644904,
  0.3875833, 0.3875833,
  0.3124668, 0.3131414,
  0.0006404052, 0.0006404052,
  0.0002255228, 0.0002292489,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  6.305695, 6.305695,
  4.104105, 4.123878,
  9.619361, 9.619361,
  5.300735, 5.339522,
  15.11261, 15.11261,
  9.843261, 9.890586,
  15.53289, 15.53289,
  9.788972, 9.84056,
  15.78795, 15.78795,
  10.63405, 10.68034,
  12.50484, 12.50484,
  10.44198, 10.4605,
  8.311556, 8.311556,
  7.58878, 7.595272,
  11.4758, 11.4758,
  7.975823, 8.007257,
  12.6149, 12.6149,
  8.363544, 8.401727,
  11.99652, 11.99652,
  8.17718, 8.211483,
  12.32582, 12.32582,
  12.48102, 12.47963,
  10.90409, 10.90409,
  8.795409, 8.814348,
  8.110285, 8.110285,
  9.376361, 9.364989,
  6.87991, 6.87991,
  7.505955, 7.500333,
  5.004357, 5.004357,
  6.470951, 6.457779,
  5.39528, 5.39528,
  5.321359, 5.322023,
  5.812306, 5.812306,
  3.678902, 3.698063,
  3.029098, 3.029098,
  0.8521963, 0.8717476,
  0.3302004, 0.3302004,
  0.03827901, 0.04090083,
  0.0003269068, 0.0003269068,
  2.896259e-05, 3.16385e-05,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  52.78875, 52.78875,
  29.44508, 29.65474,
  62.90112, 62.90112,
  35.70272, 35.94699,
  67.95486, 67.95486,
  42.00377, 42.23684,
  74.44737, 74.44737,
  45.38539, 45.6464,
  72.80553, 72.80553,
  47.43408, 47.66195,
  66.05341, 66.05341,
  48.60946, 48.76612,
  52.11737, 52.11737,
  37.65244, 37.78235,
  43.23641, 43.23641,
  31.64022, 31.74437,
  40.23101, 40.23101,
  27.49651, 27.61089,
  35.4647, 35.4647,
  24.02641, 24.12914,
  28.60297, 28.60297,
  21.35393, 21.41903,
  26.35934, 26.35934,
  19.16726, 19.23185,
  23.30768, 23.30768,
  19.56248, 19.59612,
  22.39705, 22.39705,
  16.40843, 16.46221,
  20.8924, 20.8924,
  15.89114, 15.93606,
  20.37545, 20.37545,
  15.04084, 15.08875,
  14.29356, 14.29356,
  14.06448, 14.06654,
  12.53311, 12.53311,
  11.62007, 11.62827,
  11.37377, 11.37377,
  11.27065, 11.27157,
  2.527729, 2.527729,
  4.128578, 4.114201,
  0.00144631, 0.00144631,
  0.01579883, 0.01566993,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  78.25938, 78.25938,
  55.71166, 55.91417,
  77.79131, 77.79131,
  55.80183, 55.99932,
  70.49044, 70.49044,
  49.66177, 49.84883,
  72.14246, 72.14246,
  52.70153, 52.87614,
  70.18784, 70.18784,
  51.74885, 51.91445,
  63.91494, 63.91494,
  51.95892, 52.0663,
  53.02873, 53.02873,
  49.13683, 49.17179,
  46.77215, 46.77215,
  46.32254, 46.32658,
  45.71366, 45.71366,
  42.7886, 42.81488,
  46.00961, 46.00961,
  41.46438, 41.5052,
  41.39309, 41.39309,
  38.53631, 38.56197,
  38.12512, 38.12512,
  34.77702, 34.80709,
  38.54844, 38.54844,
  35.21801, 35.24792,
  37.32542, 37.32542,
  32.14968, 32.19617,
  33.03171, 33.03171,
  28.47952, 28.5204,
  32.97549, 32.97549,
  28.30342, 28.34538,
  30.70425, 30.70425,
  26.68898, 26.72504,
  27.28682, 27.28682,
  22.63087, 22.67269,
  18.55352, 18.55352,
  13.23132, 13.27912,
  10.06217, 10.06217,
  7.522776, 7.545583,
  0.2771406, 0.2771406,
  0.1235882, 0.1249673,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  90.34143, 90.34143,
  84.88987, 84.93883,
  92.25782, 92.25782,
  85.04118, 85.10599,
  92.46198, 92.46198,
  87.67979, 87.72275,
  92.9602, 92.9602,
  81.43403, 81.53754,
  89.92547, 89.92547,
  82.40402, 82.47157,
  86.29021, 86.29021,
  82.97136, 83.00117,
  85.49364, 85.49364,
  82.41571, 82.44335,
  83.46843, 83.46843,
  83.60523, 83.604,
  79.06779, 79.06779,
  78.00068, 78.01027,
  77.09541, 77.09541,
  74.40504, 74.42921,
  72.33126, 72.33126,
  72.34224, 72.34214,
  67.31396, 67.31396,
  68.51383, 68.50306,
  65.54859, 65.54859,
  64.02675, 64.04041,
  64.63265, 64.63265,
  61.90753, 61.932,
  63.3524, 63.3524,
  61.17812, 61.19764,
  62.15071, 62.15071,
  60.14611, 60.16412,
  58.88877, 58.88877,
  56.30418, 56.3274,
  52.84317, 52.84317,
  51.05177, 51.06786,
  46.24502, 46.24502,
  44.43304, 44.44932,
  29.9822, 29.9822,
  30.04417, 30.04361,
  3.414676, 3.414676,
  4.429391, 4.420278,
  0.005693896, 0.005693896,
  0.02146333, 0.0213217,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  82.07555, 82.07555,
  66.60013, 66.73912,
  82.00278, 82.00278,
  69.00137, 69.11814,
  75.74184, 75.74184,
  64.89709, 64.99448,
  70.5143, 70.5143,
  54.16298, 54.30984,
  67.87514, 67.87514,
  53.47395, 53.60329,
  63.19024, 63.19024,
  54.58491, 54.6622,
  56.56672, 56.56672,
  53.20623, 53.23641,
  54.2597, 54.2597,
  47.8769, 47.93422,
  46.62695, 46.62695,
  42.96897, 43.00183,
  43.87945, 43.87945,
  40.04974, 40.08414,
  43.85063, 43.85063,
  38.52614, 38.57396,
  43.65066, 43.65066,
  36.79166, 36.85326,
  42.34803, 42.34803,
  36.01804, 36.07489,
  39.31591, 39.31591,
  34.72325, 34.7645,
  38.09743, 38.09743,
  34.08432, 34.12037,
  37.17603, 37.17603,
  32.92831, 32.96646,
  37.9944, 37.9944,
  33.44738, 33.48822,
  42.14789, 42.14789,
  34.9526, 35.01722,
  41.21495, 41.21495,
  33.10981, 33.1826,
  38.56582, 38.56582,
  32.08443, 32.14264,
  24.24236, 24.24236,
  21.28824, 21.31477,
  1.679659, 1.679659,
  1.612889, 1.613489,
  9.447462e-06, 9.447462e-06,
  0.0004018998, 0.0003983751,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  75.57242, 75.57242,
  61.86242, 61.98555,
  77.92242, 77.92242,
  59.18376, 59.35206,
  70.1525, 70.1525,
  59.28236, 59.37999,
  66.78737, 66.78737,
  45.81137, 45.99977,
  56.52939, 56.52939,
  48.8796, 48.9483,
  53.07075, 53.07075,
  42.90758, 42.99886,
  48.54192, 48.54192,
  38.23595, 38.32851,
  43.00229, 43.00229,
  31.73748, 31.83865,
  41.95842, 41.95842,
  31.99343, 32.08292,
  35.44351, 35.44351,
  29.31606, 29.37109,
  31.63778, 31.63778,
  25.93102, 25.98228,
  30.0705, 30.0705,
  25.43577, 25.4774,
  29.29236, 29.29236,
  24.63131, 24.67317,
  26.73204, 26.73204,
  22.71109, 22.7472,
  24.88805, 24.88805,
  21.42374, 21.45486,
  25.23137, 25.23137,
  20.08922, 20.1354,
  27.22157, 27.22157,
  20.97085, 21.02699,
  22.09079, 22.09079,
  18.7704, 18.80022,
  25.38029, 25.38029,
  19.37717, 19.43109,
  20.74439, 20.74439,
  13.8392, 13.90122,
  16.07204, 16.07204,
  9.729834, 9.786795,
  5.756322, 5.756322,
  3.100231, 3.124086,
  1.94941, 1.94941,
  0.4256229, 0.4393084,
  0.08133447, 0.08133447,
  0.01130016, 0.01192916,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  85.31528, 85.31528,
  64.4229, 64.61054,
  80.38901, 80.38901,
  67.32265, 67.44,
  70.02403, 70.02403,
  54.43231, 54.57234,
  67.64642, 67.64642,
  38.93146, 39.18935,
  64.14961, 64.14961,
  37.92901, 38.1645,
  59.32875, 59.32875,
  38.6173, 38.80331,
  50.71839, 50.71839,
  40.14064, 40.23564,
  42.64672, 42.64672,
  33.30913, 33.39299,
  34.75709, 34.75709,
  30.42414, 30.46306,
  30.59479, 30.59479,
  23.80723, 23.86819,
  25.8657, 25.8657,
  19.71703, 19.77225,
  24.11697, 24.11697,
  17.63501, 17.69323,
  20.70873, 20.70873,
  16.52056, 16.55817,
  19.19666, 19.19666,
  15.52788, 15.56083,
  18.10356, 18.10356,
  14.71966, 14.75005,
  15.12522, 15.12522,
  13.05223, 13.07085,
  15.09255, 15.09255,
  11.32769, 11.3615,
  12.57122, 12.57122,
  7.992382, 8.033505,
  11.63809, 11.63809,
  8.030373, 8.062774,
  11.49622, 11.49622,
  8.499177, 8.526093,
  11.97542, 11.97542,
  8.251622, 8.285067,
  8.411666, 8.411666,
  7.367039, 7.37642,
  3.226112, 3.226112,
  2.283622, 2.292087,
  0.2270149, 0.2270149,
  0.02620136, 0.02800491,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  85.03723, 85.03723,
  69.98151, 70.11672,
  86.09824, 86.09824,
  71.15895, 71.29313,
  82.83266, 82.83266,
  74.89445, 74.96574,
  74.31833, 74.31833,
  61.47178, 61.58715,
  63.00635, 63.00635,
  62.71317, 62.7158,
  53.64307, 53.64307,
  54.52642, 54.51849,
  50.97019, 50.97019,
  42.01061, 42.09108,
  47.37215, 47.37215,
  37.54349, 37.63176,
  42.65371, 42.65371,
  37.32167, 37.36956,
  39.60907, 39.60907,
  36.27053, 36.30052,
  31.97943, 31.97943,
  30.43582, 30.44969,
  31.36078, 31.36078,
  27.99077, 28.02104,
  30.62183, 30.62183,
  26.93032, 26.96347,
  30.42588, 30.42588,
  25.81332, 25.85475,
  30.29451, 30.29451,
  24.74087, 24.79075,
  27.81119, 27.81119,
  24.63252, 24.66107,
  24.75825, 24.75825,
  22.12754, 22.15117,
  23.25025, 23.25025,
  19.53045, 19.56386,
  20.37233, 20.37233,
  18.01965, 18.04078,
  19.54182, 19.54182,
  18.0434, 18.05686,
  19.41059, 19.41059,
  18.18313, 18.19416,
  17.36652, 17.36652,
  16.52367, 16.53124,
  12.8668, 12.8668,
  11.42169, 11.43467,
  8.598517, 8.598517,
  8.016893, 8.022117,
  6.430734, 6.430734,
  6.529112, 6.528229,
  8.801474, 8.801474,
  7.962327, 7.969864,
  12.13899, 12.13899,
  8.730135, 8.760751,
  9.342519, 9.342519,
  6.678372, 6.702299,
  3.141517, 3.141517,
  2.251501, 2.259494,
  0.0207718, 0.0207718,
  0.001840296, 0.002010324,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  82.60934, 82.60934,
  72.70028, 72.78928,
  84.21429, 84.21429,
  74.55608, 74.64282,
  82.75797, 82.75797,
  75.81718, 75.87952,
  77.01313, 77.01313,
  66.11024, 66.20815,
  78.98689, 78.98689,
  62.76892, 62.91457,
  73.35776, 73.35776,
  65.57955, 65.64941,
  62.18752, 62.18752,
  58.99772, 59.02637,
  55.50527, 55.50527,
  51.0866, 51.12629,
  49.92838, 49.92838,
  44.05367, 44.10643,
  48.179, 48.179,
  41.31121, 41.37289,
  46.5518, 46.5518,
  40.62423, 40.67746,
  45.5034, 45.5034,
  40.82119, 40.86324,
  43.62707, 43.62707,
  39.62011, 39.65609,
  40.55501, 40.55501,
  37.90501, 37.92881,
  34.99547, 34.99547,
  34.1201, 34.12796,
  31.20151, 31.20151,
  30.55139, 30.55723,
  24.57554, 24.57554,
  24.59276, 24.59261,
  19.68936, 19.68936,
  17.74133, 17.75883,
  18.83914, 18.83914,
  15.81509, 15.84225,
  14.72225, 14.72225,
  13.29542, 13.30824,
  10.40821, 10.40821,
  8.842506, 8.856568,
  6.340128, 6.340128,
  5.768337, 5.773472,
  3.56518, 3.56518,
  3.826853, 3.824502,
  2.118745, 2.118745,
  3.001197, 2.993272,
  0.8323127, 0.8323127,
  1.302154, 1.297935,
  0.04298011, 0.04298011,
  0.1871182, 0.1858237,
  0.01688335, 0.01688335,
  0.001914187, 0.002048628,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  70.97849, 70.97849,
  52.80009, 52.96336,
  72.83981, 72.83981,
  55.71019, 55.86404,
  73.89983, 73.89983,
  55.46131, 55.62691,
  79.26441, 79.26441,
  52.06144, 52.30576,
  76.82455, 76.82455,
  62.69462, 62.82153,
  73.82509, 73.82509,
  57.68683, 57.83178,
  64.85822, 64.85822,
  53.97697, 54.0747,
  54.44579, 54.44579,
  51.72076, 51.74523,
  40.64886, 40.64886,
  42.33951, 42.32433,
  33.94129, 33.94129,
  39.21353, 39.16618,
  31.5133, 31.5133,
  33.67567, 33.65625,
  29.16374, 29.16374,
  31.15042, 31.13258,
  29.01032, 29.01032,
  30.68007, 30.66508,
  28.86435, 28.86435,
  27.54799, 27.55981,
  26.40376, 26.40376,
  25.29453, 25.30449,
  24.66853, 24.66853,
  23.59821, 23.60782,
  21.80454, 21.80454,
  22.41611, 22.41062,
  17.00998, 17.00998,
  19.22733, 19.20742,
  13.58867, 13.58867,
  14.93714, 14.92502,
  13.58361, 13.58361,
  13.39033, 13.39207,
  7.873963, 7.873963,
  8.251403, 8.248013,
  0.6397788, 0.6397788,
  0.5380676, 0.5389811,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  29.47814, 29.47814,
  17.63503, 17.7414,
  36.06388, 36.06388,
  21.95141, 22.07816,
  46.82228, 46.82228,
  31.43551, 31.5737,
  53.9309, 53.9309,
  43.53775, 43.6311,
  57.79251, 57.79251,
  51.27372, 51.33227,
  54.46742, 54.46742,
  47.63, 47.69141,
  43.97896, 43.97896,
  32.72979, 32.83082,
  36.17587, 36.17587,
  28.48501, 28.55409,
  31.61798, 31.61798,
  26.53037, 26.57607,
  28.81577, 28.81577,
  25.16603, 25.1988,
  26.14541, 26.14541,
  23.31073, 23.33619,
  22.99272, 22.99272,
  21.72667, 21.73804,
  20.60434, 20.60434,
  18.82668, 18.84265,
  19.70421, 19.70421,
  18.95456, 18.96129,
  18.31168, 18.31168,
  18.32328, 18.32318,
  12.55419, 12.55419,
  13.33557, 13.32855,
  8.78577, 8.78577,
  9.86748, 9.857765,
  5.064898, 5.064898,
  6.223226, 6.212822,
  1.608376, 1.608376,
  4.042251, 4.020392,
  0.1179678, 0.1179678,
  1.762088, 1.747322,
  0.002788691, 0.002788691,
  0.0002470665, 0.0002698935,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  6.984023, 6.984023,
  3.515866, 3.547014,
  9.97495, 9.97495,
  6.759108, 6.78799,
  21.77545, 21.77545,
  11.48474, 11.57716,
  20.32658, 20.32658,
  10.64229, 10.72926,
  12.24531, 12.24531,
  7.71451, 7.755202,
  8.728997, 8.728997,
  5.91965, 5.944881,
  6.558224, 6.558224,
  5.320841, 5.331954,
  3.923496, 3.923496,
  3.153401, 3.160317,
  4.36447, 4.36447,
  3.476101, 3.48408,
  5.520906, 5.520906,
  4.614528, 4.622669,
  6.644382, 6.644382,
  5.95359, 5.959794,
  8.878189, 8.878189,
  8.136605, 8.143266,
  12.65983, 12.65983,
  9.234739, 9.265501,
  14.76682, 14.76682,
  9.195086, 9.245127,
  14.47866, 14.47866,
  11.65589, 11.68125,
  14.34762, 14.34762,
  11.18871, 11.21708,
  14.58594, 14.58594,
  10.63648, 10.67195,
  10.93098, 10.93098,
  10.27124, 10.27717,
  2.089658, 2.089658,
  1.732257, 1.735467,
  0.006255088, 0.006255088,
  0.009104982, 0.009079386,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0 ;

 lat = -89.5, -88.5 ;

 lat_bnds =
  -90, -89,
  -89, -88 ;

 lev = 0.99795, 0.99279, 0.98540739915, 0.9756590957, 0.9633249281, 
    0.94807624475, 0.92954604845, 0.9072989285, 0.88081805335, 0.84950967285, 
    0.8127897223, 0.7701018362, 0.72101394975, 0.6653174996, 0.6032088506, 
    0.5358132351, 0.4658290421, 0.3972976087, 0.33404935575, 0.2781749219, 
    0.22998078655, 0.1888851393, 0.15409188855, 0.1248356931, 0.10040876315, 
    0.08016256785, 0.06350800645, 0.0499146627, 0.038909233, 0.0300732337, 
    0.02304010415, 0.0174918294, 0.0131552082, 0.00979788985, 0.0072242975, 
    0.0052715454, 0.0038054455, 0.0027166834, 0.0019172284, 0.00133702575, 
    0.0009210024, 0.00062640445, 0.00042046895, 0.000278422, 0.00018159735, 
    0.00011571225, 7.032955e-05, 3.93429e-05, 1.84861e-05 ;

 lev_bnds =
  1, 0.9959,
  0.9959, 0.98968,
  0.98968, 0.9811347983,
  0.9811347983, 0.9701833931,
  0.9701833931, 0.9564664631,
  0.9564664631, 0.9396860264,
  0.9396860264, 0.9194060705,
  0.9194060705, 0.8951917865,
  0.8951917865, 0.8664443202,
  0.8664443202, 0.8325750255,
  0.8325750255, 0.7930044191,
  0.7930044191, 0.7471992533,
  0.7471992533, 0.6948286462,
  0.6948286462, 0.635806353,
  0.635806353, 0.5706113482,
  0.5706113482, 0.501015122,
  0.501015122, 0.4306429622,
  0.4306429622, 0.3639522552,
  0.3639522552, 0.3041464563,
  0.3041464563, 0.2522033875,
  0.2522033875, 0.2077581856,
  0.2077581856, 0.170012093,
  0.170012093, 0.1381716841,
  0.1381716841, 0.1114997021,
  0.1114997021, 0.0893178242,
  0.0893178242, 0.0710073115,
  0.0710073115, 0.0560087014,
  0.0560087014, 0.043820624,
  0.043820624, 0.033997842,
  0.033997842, 0.0261486254,
  0.0261486254, 0.0199315829,
  0.0199315829, 0.0150520759,
  0.0150520759, 0.0112583405,
  0.0112583405, 0.0083374392,
  0.0083374392, 0.0061111558,
  0.0061111558, 0.004431935,
  0.004431935, 0.003178956,
  0.003178956, 0.0022544108,
  0.0022544108, 0.001580046,
  0.001580046, 0.0010940055,
  0.0010940055, 0.0007479993,
  0.0007479993, 0.0005048096,
  0.0005048096, 0.0003361283,
  0.0003361283, 0.0002207157,
  0.0002207157, 0.000142479,
  0.000142479, 8.89455e-05,
  8.89455e-05, 5.17136e-05,
  5.17136e-05, 2.69722e-05,
  2.69722e-05, 1e-05 ;

 lon = 0.625, 1.875 ;

 lon_bnds =
  0, 1.25,
  1.25, 2.5 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825 ;
}
