netcdf ocean_monthly.200001-200412.sos {
dimensions:
	time = UNLIMITED ; // (60 currently)
	nv = 2 ;
	yh = 576 ;
	xh = 720 ;
variables:
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:_FillValue = 1.e+20 ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1850-01-01 00:00:00" ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:_FillValue = 1.e+20 ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1850-01-01 00:00:00" ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:_FillValue = 1.e+20 ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	float sos(time, yh, xh) ;
		sos:long_name = "Sea Surface Salinity" ;
		sos:units = "psu" ;
		sos:missing_value = 1.e+20f ;
		sos:_FillValue = 1.e+20f ;
		sos:cell_methods = "area:mean yh:mean xh:mean time: mean" ;
		sos:cell_measures = "area: areacello" ;
		sos:time_avg_info = "average_T1,average_T2,average_DT" ;
		sos:standard_name = "sea_surface_salinity" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1850-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 1850-01-01 00:00:00" ;
		time_bnds:missing_value = 1.e+20 ;
		time_bnds:_FillValue = 1.e+20 ;
	double xh(xh) ;
		xh:long_name = "h point nominal longitude" ;
		xh:units = "degrees_east" ;
		xh:axis = "X" ;
	double yh(yh) ;
		yh:long_name = "h point nominal latitude" ;
		yh:units = "degrees_north" ;
		yh:axis = "Y" ;

// global attributes:
		:filename = "ocean_monthly.200001-200412.sos.nc" ;
		:title = "ESM4_historical_D151" ;
		:associated_files = "areacello: 20000101.ocean_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:external_variables = "areacello" ;
data:

 nv = 1, 2 ;

 time = 54765.5, 54795, 54824.5, 54855, 54885.5, 54916, 54946.5, 54977.5, 
    55008, 55038.5, 55069, 55099.5, 55130.5, 55160, 55189.5, 55220, 55250.5, 
    55281, 55311.5, 55342.5, 55373, 55403.5, 55434, 55464.5, 55495.5, 55525, 
    55554.5, 55585, 55615.5, 55646, 55676.5, 55707.5, 55738, 55768.5, 55799, 
    55829.5, 55860.5, 55890, 55919.5, 55950, 55980.5, 56011, 56041.5, 
    56072.5, 56103, 56133.5, 56164, 56194.5, 56225.5, 56255, 56284.5, 56315, 
    56345.5, 56376, 56406.5, 56437.5, 56468, 56498.5, 56529, 56559.5 ;

 xh = -299.75, -299.25, -298.75, -298.25, -297.75, -297.25, -296.75, -296.25, 
    -295.75, -295.25, -294.75, -294.25, -293.75, -293.25, -292.75, -292.25, 
    -291.75, -291.25, -290.75, -290.25, -289.75, -289.25, -288.75, -288.25, 
    -287.75, -287.25, -286.75, -286.25, -285.75, -285.25, -284.75, -284.25, 
    -283.75, -283.25, -282.75, -282.25, -281.75, -281.25, -280.75, -280.25, 
    -279.75, -279.25, -278.75, -278.25, -277.75, -277.25, -276.75, -276.25, 
    -275.75, -275.25, -274.75, -274.25, -273.75, -273.25, -272.75, -272.25, 
    -271.75, -271.25, -270.75, -270.25, -269.75, -269.25, -268.75, -268.25, 
    -267.75, -267.25, -266.75, -266.25, -265.75, -265.25, -264.75, -264.25, 
    -263.75, -263.25, -262.75, -262.25, -261.75, -261.25, -260.75, -260.25, 
    -259.75, -259.25, -258.75, -258.25, -257.75, -257.25, -256.75, -256.25, 
    -255.75, -255.25, -254.75, -254.25, -253.75, -253.25, -252.75, -252.25, 
    -251.75, -251.25, -250.75, -250.25, -249.75, -249.25, -248.75, -248.25, 
    -247.75, -247.25, -246.75, -246.25, -245.75, -245.25, -244.75, -244.25, 
    -243.75, -243.25, -242.75, -242.25, -241.75, -241.25, -240.75, -240.25, 
    -239.75, -239.25, -238.75, -238.25, -237.75, -237.25, -236.75, -236.25, 
    -235.75, -235.25, -234.75, -234.25, -233.75, -233.25, -232.75, -232.25, 
    -231.75, -231.25, -230.75, -230.25, -229.75, -229.25, -228.75, -228.25, 
    -227.75, -227.25, -226.75, -226.25, -225.75, -225.25, -224.75, -224.25, 
    -223.75, -223.25, -222.75, -222.25, -221.75, -221.25, -220.75, -220.25, 
    -219.75, -219.25, -218.75, -218.25, -217.75, -217.25, -216.75, -216.25, 
    -215.75, -215.25, -214.75, -214.25, -213.75, -213.25, -212.75, -212.25, 
    -211.75, -211.25, -210.75, -210.25, -209.75, -209.25, -208.75, -208.25, 
    -207.75, -207.25, -206.75, -206.25, -205.75, -205.25, -204.75, -204.25, 
    -203.75, -203.25, -202.75, -202.25, -201.75, -201.25, -200.75, -200.25, 
    -199.75, -199.25, -198.75, -198.25, -197.75, -197.25, -196.75, -196.25, 
    -195.75, -195.25, -194.75, -194.25, -193.75, -193.25, -192.75, -192.25, 
    -191.75, -191.25, -190.75, -190.25, -189.75, -189.25, -188.75, -188.25, 
    -187.75, -187.25, -186.75, -186.25, -185.75, -185.25, -184.75, -184.25, 
    -183.75, -183.25, -182.75, -182.25, -181.75, -181.25, -180.75, -180.25, 
    -179.75, -179.25, -178.75, -178.25, -177.75, -177.25, -176.75, -176.25, 
    -175.75, -175.25, -174.75, -174.25, -173.75, -173.25, -172.75, -172.25, 
    -171.75, -171.25, -170.75, -170.25, -169.75, -169.25, -168.75, -168.25, 
    -167.75, -167.25, -166.75, -166.25, -165.75, -165.25, -164.75, -164.25, 
    -163.75, -163.25, -162.75, -162.25, -161.75, -161.25, -160.75, -160.25, 
    -159.75, -159.25, -158.75, -158.25, -157.75, -157.25, -156.75, -156.25, 
    -155.75, -155.25, -154.75, -154.25, -153.75, -153.25, -152.75, -152.25, 
    -151.75, -151.25, -150.75, -150.25, -149.75, -149.25, -148.75, -148.25, 
    -147.75, -147.25, -146.75, -146.25, -145.75, -145.25, -144.75, -144.25, 
    -143.75, -143.25, -142.75, -142.25, -141.75, -141.25, -140.75, -140.25, 
    -139.75, -139.25, -138.75, -138.25, -137.75, -137.25, -136.75, -136.25, 
    -135.75, -135.25, -134.75, -134.25, -133.75, -133.25, -132.75, -132.25, 
    -131.75, -131.25, -130.75, -130.25, -129.75, -129.25, -128.75, -128.25, 
    -127.75, -127.25, -126.75, -126.25, -125.75, -125.25, -124.75, -124.25, 
    -123.75, -123.25, -122.75, -122.25, -121.75, -121.25, -120.75, -120.25, 
    -119.75, -119.25, -118.75, -118.25, -117.75, -117.25, -116.75, -116.25, 
    -115.75, -115.25, -114.75, -114.25, -113.75, -113.25, -112.75, -112.25, 
    -111.75, -111.25, -110.75, -110.25, -109.75, -109.25, -108.75, -108.25, 
    -107.75, -107.25, -106.75, -106.25, -105.75, -105.25, -104.75, -104.25, 
    -103.75, -103.25, -102.75, -102.25, -101.75, -101.25, -100.75, -100.25, 
    -99.75, -99.25, -98.75, -98.25, -97.75, -97.25, -96.75, -96.25, -95.75, 
    -95.25, -94.75, -94.25, -93.75, -93.25, -92.75, -92.25, -91.75, -91.25, 
    -90.75, -90.25, -89.75, -89.25, -88.75, -88.25, -87.75, -87.25, -86.75, 
    -86.25, -85.75, -85.25, -84.75, -84.25, -83.75, -83.25, -82.75, -82.25, 
    -81.75, -81.25, -80.75, -80.25, -79.75, -79.25, -78.75, -78.25, -77.75, 
    -77.25, -76.75, -76.25, -75.75, -75.25, -74.75, -74.25, -73.75, -73.25, 
    -72.75, -72.25, -71.75, -71.25, -70.75, -70.25, -69.75, -69.25, -68.75, 
    -68.25, -67.75, -67.25, -66.75, -66.25, -65.75, -65.25, -64.75, -64.25, 
    -63.75, -63.25, -62.75, -62.25, -61.75, -61.25, -60.75, -60.25, -59.75, 
    -59.25, -58.75, -58.25, -57.75, -57.25, -56.75, -56.25, -55.75, -55.25, 
    -54.75, -54.25, -53.75, -53.25, -52.75, -52.25, -51.75, -51.25, -50.75, 
    -50.25, -49.75, -49.25, -48.75, -48.25, -47.75, -47.25, -46.75, -46.25, 
    -45.75, -45.25, -44.75, -44.25, -43.75, -43.25, -42.75, -42.25, -41.75, 
    -41.25, -40.75, -40.25, -39.75, -39.25, -38.75, -38.25, -37.75, -37.25, 
    -36.75, -36.25, -35.75, -35.25, -34.75, -34.25, -33.75, -33.25, -32.75, 
    -32.25, -31.75, -31.25, -30.75, -30.25, -29.75, -29.25, -28.75, -28.25, 
    -27.75, -27.25, -26.75, -26.25, -25.75, -25.25, -24.75, -24.25, -23.75, 
    -23.25, -22.75, -22.25, -21.75, -21.25, -20.75, -20.25, -19.75, -19.25, 
    -18.75, -18.25, -17.75, -17.25, -16.75, -16.25, -15.75, -15.25, -14.75, 
    -14.25, -13.75, -13.25, -12.75, -12.25, -11.75, -11.25, -10.75, -10.25, 
    -9.75, -9.25, -8.75, -8.25, -7.75, -7.25, -6.75, -6.25, -5.75, -5.25, 
    -4.75, -4.25, -3.75, -3.25, -2.75, -2.25, -1.75, -1.25, -0.75, -0.25, 
    0.25, 0.75, 1.25, 1.75, 2.25, 2.75, 3.25, 3.75, 4.25, 4.75, 5.25, 5.75, 
    6.25, 6.75, 7.25, 7.75, 8.25, 8.75, 9.25, 9.75, 10.25, 10.75, 11.25, 
    11.75, 12.25, 12.75, 13.25, 13.75, 14.25, 14.75, 15.25, 15.75, 16.25, 
    16.75, 17.25, 17.75, 18.25, 18.75, 19.25, 19.75, 20.25, 20.75, 21.25, 
    21.75, 22.25, 22.75, 23.25, 23.75, 24.25, 24.75, 25.25, 25.75, 26.25, 
    26.75, 27.25, 27.75, 28.25, 28.75, 29.25, 29.75, 30.25, 30.75, 31.25, 
    31.75, 32.25, 32.75, 33.25, 33.75, 34.25, 34.75, 35.25, 35.75, 36.25, 
    36.75, 37.25, 37.75, 38.25, 38.75, 39.25, 39.75, 40.25, 40.75, 41.25, 
    41.75, 42.25, 42.75, 43.25, 43.75, 44.25, 44.75, 45.25, 45.75, 46.25, 
    46.75, 47.25, 47.75, 48.25, 48.75, 49.25, 49.75, 50.25, 50.75, 51.25, 
    51.75, 52.25, 52.75, 53.25, 53.75, 54.25, 54.75, 55.25, 55.75, 56.25, 
    56.75, 57.25, 57.75, 58.25, 58.75, 59.25, 59.75 ;

 yh = -77.9079375348705, -77.7238126046114, -77.5396876743523, 
    -77.3555627440933, -77.1714378138342, -76.9873128835751, 
    -76.8031879533161, -76.619063023057, -76.4349380927979, 
    -76.2508131625389, -76.0666882322798, -75.8825633020207, 
    -75.6984383717617, -75.5143134415026, -75.3301885112435, 
    -75.1460635809845, -74.9619386507254, -74.7778137204664, 
    -74.5936887902073, -74.4095638599482, -74.2254389296892, 
    -74.0413139994301, -73.857189069171, -73.673064138912, -73.4889392086529, 
    -73.3048142783938, -73.1206893481348, -72.9365644178757, 
    -72.7524394876166, -72.5683145573576, -72.3841896270985, 
    -72.2000646968394, -72.0159397665804, -71.8318148363213, 
    -71.6476899060622, -71.4635649758032, -71.2794400455441, 
    -71.095315115285, -70.911190185026, -70.7270652547669, -70.5429403245078, 
    -70.3588153942488, -70.1746904639897, -69.9905655337306, 
    -69.8064406034716, -69.6223156732125, -69.4381907429535, 
    -69.2540658126944, -69.0699408824353, -68.8858159521763, 
    -68.7016910219172, -68.5175660916581, -68.3334411613991, -68.14931623114, 
    -67.9636445304209, -67.7752866505205, -67.5854009965385, 
    -67.3939772792524, -67.2010051944971, -67.0064744247379, 
    -66.8103746406885, -66.6126955029787, -66.4134266638701, 
    -66.2125577690213, -66.0100784593041, -65.8059783726705, 
    -65.6002471460721, -65.3928744174328, -65.1838498276744, 
    -64.9731630227985, -64.760803656022, -64.5467613899703, 
    -64.3310258989275, -64.1135868711439, -63.894434011203, 
    -63.6735570424482, -63.4509457094688, -63.2265897806486, 
    -63.0004790507758, -62.7726033437149, -62.5429525151436, 
    -62.3115164553525, -62.0782850921101, -61.8432483935938, 
    -61.6063963713863, -61.3677190835396, -61.1272066377062, 
    -60.884849194338, -60.6406369699546, -60.3945602404801, -60.14660934465, 
    -59.8967746874882, -59.6450467438542, -59.3914160620619, 
    -59.1358732675693, -58.8784090667402, -58.6190142506776, 
    -58.3576796991292, -58.0943963844658, -57.8291553757318, 
    -57.5619478427679, -57.2927650604075, -57.0215984127446, 
    -56.7484393974749, -56.4732796303085, -56.1961108494559, 
    -55.9169249201846, -55.6357138394475, -55.3524697405834, 
    -55.0671848980862, -54.7798517324457, -54.4904628150566, 
    -54.199010873197, -53.9054887950733, -53.6098896349336, 
    -53.3122066182453, -53.0124331469381, -52.7105628047106, 
    -52.4065893623985, -52.1005067834039, -51.7923092291839, 
    -51.4819910647963, -51.1695468645014, -50.8549714174182, 
    -50.5382597332318, -50.2194070479511, -49.8984088297146, 
    -49.5752607846407, -49.2499588627218, -48.9224992637582, 
    -48.5928784433296, -48.2610931188013, -47.9271402753627, 
    -47.5910171720938, -47.2527213480571, -46.9122506284122, 
    -46.5696031305474, -46.2247772702279, -45.8777717677532, 
    -45.5285856541224, -45.1772182772023, -44.8236693078935, 
    -44.4679387462917, -44.1100269278373, -43.7499345294513, 
    -43.3876625756504, -43.0232124446377, -42.6565858743633, 
    -42.2877849685499, -41.9168122026777, -41.5436704299229, 
    -41.1683628870455, -40.790893200218, -40.4112653907925, 
    -40.0294838809968, -39.6455534995561, -39.2594794872318, 
    -38.8712675022735, -38.4809236257751, -38.0884543669302, 
    -37.6938666681796, -37.2971679102448, -36.8983659170386, 
    -36.4974689604493, -36.0944857649878, -35.6894255122942, 
    -35.2822978454935, -34.8731128733961, -34.461881174534, 
    -34.0486138010269, -33.6333222822699, -33.2160186284369, 
    -32.7967153337909, -32.3754253797966, -31.952162238025, 
    -31.5269398728455, -31.0997727438981, -30.6706758083373, 
    -30.2396645228428, -29.8067548453888, -29.3722350905309, 
    -28.9369844818468, -28.5011135682704, -28.0647328987354, 
    -27.6279530221758, -27.1908844875253, -26.7536378437177, 
    -26.316323639687, -25.8790524243669, -25.4419347466912, 
    -25.0050811555939, -24.5686022000086, -24.1326084288694, 
    -23.6972103911098, -23.2625186356639, -22.8286437114655, 
    -22.3956961674483, -21.9637865525462, -21.533025415693, 
    -21.1035233058226, -20.6753907718688, -20.2487383627654, 
    -19.8236766274463, -19.4003161148452, -18.9787673738961, 
    -18.5591409535327, -18.1415474026888, -17.7260972702984, 
    -17.3129011052952, -16.9020694566131, -16.4937128731858, 
    -16.0879419039473, -15.6848670978313, -15.2845990037717, 
    -14.8872481707024, -14.492925147557, -14.1017404832696, 
    -13.7138047267738, -13.3292284270036, -12.9481221328927, 
    -12.5705963933751, -12.1967617573844, -11.8267287738547, 
    -11.4606079917196, -11.098509959913, -10.7405452273687, 
    -10.3868243430207, -10.0374578558026, -9.6925563146484, 
    -9.35223026849184, -9.01659026626678, -8.68574685690705, 
    -8.35981058934647, -8.03889201251887, -7.7231016753581, 
    -7.41255012679797, -7.10734791577232, -6.80760559121498, 
    -6.51343370205977, -6.22494279724053, -5.94224342569109, 
    -5.66544613634527, -5.39466147813692, -5.12999999999985, 
    -4.87179487179475, -4.6153846153845, -4.35897435897425, -4.102564102564, 
    -3.84615384615375, -3.5897435897435, -3.33333333333325, -3.076923076923, 
    -2.82051282051275, -2.5641025641025, -2.30769230769225, -2.051282051282, 
    -1.79487179487175, -1.5384615384615, -1.28205128205125, -1.025641025641, 
    -0.76923076923075, -0.5128205128205, -0.25641025641025, -0, 
    0.25641025641025, 0.5128205128205, 0.76923076923075, 1.025641025641, 
    1.28205128205125, 1.5384615384615, 1.79487179487175, 2.051282051282, 
    2.30769230769225, 2.5641025641025, 2.82051282051275, 3.076923076923, 
    3.33333333333325, 3.5897435897435, 3.84615384615375, 4.102564102564, 
    4.35897435897425, 4.6153846153845, 4.87179487179475, 5.12999999999985, 
    5.39466147813692, 5.66544613634527, 5.94224342569109, 6.22494279724053, 
    6.51343370205977, 6.80760559121498, 7.10734791577232, 7.41255012679797, 
    7.7231016753581, 8.03889201251887, 8.35981058934647, 8.68574685690705, 
    9.01659026626678, 9.35223026849184, 9.6925563146484, 10.0374578558026, 
    10.3868243430207, 10.7405452273687, 11.098509959913, 11.4606079917196, 
    11.8267287738547, 12.1967617573844, 12.5705963933751, 12.9481221328927, 
    13.3292284270036, 13.7138047267738, 14.1017404832696, 14.492925147557, 
    14.8872481707024, 15.2845990037717, 15.6848670978313, 16.0879419039473, 
    16.4937128731858, 16.9020694566131, 17.3129011052952, 17.7260972702984, 
    18.1415474026888, 18.5591409535327, 18.9787673738961, 19.4003161148452, 
    19.8236766274463, 20.2487383627654, 20.6753907718688, 21.1035233058226, 
    21.533025415693, 21.9637865525462, 22.3956961674483, 22.8286437114655, 
    23.2625186356639, 23.6972103911098, 24.1326084288694, 24.5686022000086, 
    25.0050811555939, 25.4419347466912, 25.8790524243669, 26.316323639687, 
    26.7536378437177, 27.1908844875253, 27.6279530221758, 28.0647328987354, 
    28.5011135682704, 28.9369844818468, 29.3722350905309, 29.8067548453888, 
    30.2396645228428, 30.6706758083373, 31.0997727438981, 31.5269398728455, 
    31.952162238025, 32.3754253797966, 32.7967153337909, 33.2160186284369, 
    33.6333222822699, 34.0486138010269, 34.461881174534, 34.8731128733961, 
    35.2822978454935, 35.6894255122942, 36.0944857649878, 36.4974689604493, 
    36.8983659170386, 37.2971679102448, 37.6938666681796, 38.0884543669302, 
    38.4809236257751, 38.8712675022735, 39.2594794872318, 39.6455534995561, 
    40.0294838809968, 40.4112653907925, 40.790893200218, 41.1683628870455, 
    41.5436704299229, 41.9168122026777, 42.2877849685499, 42.6565858743633, 
    43.0232124446377, 43.3876625756504, 43.7499345294513, 44.1100269278373, 
    44.4679387462917, 44.8236693078935, 45.1772182772023, 45.5285856541224, 
    45.8777717677532, 46.2247772702279, 46.5696031305474, 46.9122506284122, 
    47.2527213480571, 47.5910171720938, 47.9271402753627, 48.2610931188013, 
    48.5928784433296, 48.9224992637582, 49.2499588627218, 49.5752607846407, 
    49.8984088297146, 50.2194070479511, 50.5382597332318, 50.8549714174182, 
    51.1695468645014, 51.4819910647963, 51.7923092291839, 52.1005067834039, 
    52.4065893623985, 52.7105628047106, 53.0124331469381, 53.3122066182453, 
    53.6098896349336, 53.9054887950733, 54.199010873197, 54.4904628150566, 
    54.7798517324457, 55.0671848980862, 55.3524697405834, 55.6357138394475, 
    55.9169249201846, 56.1961108494559, 56.4732796303085, 56.7484393974749, 
    57.0215984127446, 57.2927650604075, 57.5619478427679, 57.8291553757318, 
    58.0943963844658, 58.3576796991292, 58.6190142506776, 58.8784090667402, 
    59.1358732675693, 59.3914160620619, 59.6450467438542, 59.8967746874882, 
    60.14660934465, 60.3945602404801, 60.6406369699546, 60.884849194338, 
    61.1272066377062, 61.3677190835396, 61.6063963713863, 61.8432483935938, 
    62.0782850921101, 62.3115164553525, 62.5429525151436, 62.7726033437149, 
    63.0004790507758, 63.2265897806486, 63.4509457094688, 63.6735570424482, 
    63.894434011203, 64.1135868711439, 64.3310258989275, 64.5467613899703, 
    64.760803656022, 64.9727930851569, 65.18399314351, 65.3951932018631, 
    65.6063932602162, 65.8175933185693, 66.0287933769224, 66.2399934352755, 
    66.4511934936286, 66.6623935519817, 66.8735936103349, 67.084793668688, 
    67.2959937270411, 67.5071937853942, 67.7183938437473, 67.9295939021004, 
    68.1407939604535, 68.3519940188066, 68.5631940771597, 68.7743941355128, 
    68.9855941938659, 69.196794252219, 69.4079943105721, 69.6191943689252, 
    69.8303944272783, 70.0415944856315, 70.2527945439845, 70.4639946023377, 
    70.6751946606908, 70.8863947190439, 71.097594777397, 71.3087948357501, 
    71.5199948941032, 71.7311949524563, 71.9423950108094, 72.1535950691625, 
    72.3647951275156, 72.5759951858687, 72.7871952442218, 72.9983953025749, 
    73.209595360928, 73.4207954192811, 73.6319954776342, 73.8431955359874, 
    74.0543955943405, 74.2655956526936, 74.4767957110467, 74.6879957693998, 
    74.8991958277529, 75.110395886106, 75.3215959444591, 75.5327960028122, 
    75.7439960611653, 75.9551961195184, 76.1663961778715, 76.3775962362246, 
    76.5887962945777, 76.7999963529308, 77.011196411284, 77.2223964696371, 
    77.4335965279902, 77.6447965863433, 77.8559966446964, 78.0671967030495, 
    78.2783967614026, 78.4895968197557, 78.7007968781088, 78.9119969364619, 
    79.123196994815, 79.3343970531681, 79.5455971115212, 79.7567971698743, 
    79.9679972282274, 80.1791972865805, 80.3903973449337, 80.6015974032868, 
    80.8127974616399, 81.023997519993, 81.2351975783461, 81.4463976366992, 
    81.6575976950523, 81.8687977534054, 82.0799978117585, 82.2911978701116, 
    82.5023979284647, 82.7135979868178, 82.9247980451709, 83.135998103524, 
    83.3471981618771, 83.5583982202303, 83.7695982785834, 83.9807983369365, 
    84.1919983952896, 84.4031984536427, 84.6143985119958, 84.8255985703489, 
    85.036798628702, 85.2479986870551, 85.4591987454082, 85.6703988037613, 
    85.8815988621144, 86.0927989204675, 86.3039989788206, 86.5151990371737, 
    86.7263990955269, 86.93759915388, 87.1487992122331, 87.3599992705862, 
    87.5711993289393, 87.7823993872924, 87.9935994456455, 88.2047995039986, 
    88.4159995623517, 88.6271996207048, 88.8383996790579, 89.049599737411, 
    89.2607997957641, 89.4719998541172, 89.6831999124703, 89.8943999708235 ;
}
