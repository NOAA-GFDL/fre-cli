netcdf \00010101.atmos_daily.tile3.rlut {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float rlut(time, grid_yt, grid_xt) ;
		rlut:_FillValue = 1.e+20f ;
		rlut:missing_value = 1.e+20f ;
		rlut:units = "W m-2" ;
		rlut:long_name = "TOA Outgoing Longwave Radiation" ;
		rlut:cell_methods = "time: mean" ;
		rlut:cell_measures = "area: area" ;
		rlut:time_avg_info = "average_T1,average_T2,average_DT" ;
		rlut:standard_name = "toa_outgoing_longwave_flux" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 rlut =
  186.7222, 194.2757, 192.7097, 204.8557, 198.6682, 190.0629, 195.1854, 
    191.2768, 191.5528, 171.4344, 170.7977, 171.6754, 164.1939, 168.8092, 
    158.8546,
  188.569, 199.0868, 195.0602, 191.7088, 181.9433, 179.9996, 189.8094, 
    194.9452, 195.5129, 190.2661, 178.1034, 177.6634, 174.888, 163.1884, 
    156.7982,
  193.3486, 200.4762, 196.3385, 189.6511, 183.9561, 169.8442, 185.0716, 
    196.8983, 203.4032, 199.4102, 192.038, 180.4719, 175.3746, 171.045, 
    163.5138,
  190.5482, 197.5287, 194.6769, 197.7034, 193.525, 190.0928, 167.2314, 
    191.3926, 197.0063, 197.2567, 192.7287, 184.7601, 180.4041, 172.0914, 
    169.2234,
  192.428, 201.084, 203.5893, 202.3525, 199.8602, 197.9088, 196.4487, 
    164.582, 171.6045, 186.5409, 189.5247, 182.4898, 178.1878, 175.7353, 
    172.4164,
  198.1227, 199.3893, 200.0807, 206.8369, 208.3036, 210.6583, 201.5773, 
    197.7393, 198.9808, 189.6227, 179.2669, 175.1239, 174.4442, 166.9892, 
    170.521,
  205.4943, 208.1395, 198.7731, 194.4453, 196.5861, 208.0246, 196.0914, 
    193.8118, 195.6661, 187.9236, 179.3095, 173.8251, 169.6132, 169.3038, 
    172.2475,
  215.1657, 204.3699, 198.1151, 200.5763, 199.3142, 206.8559, 199.336, 
    195.6741, 191.0237, 177.6417, 178.0886, 169.8724, 167.5806, 163.5483, 
    169.0258,
  201.2531, 199.6181, 199.9539, 204.4133, 203.1487, 205.023, 201.4388, 
    196.647, 187.41, 188.539, 178.0096, 170.9474, 166.5488, 166.2778, 171.542,
  201.4429, 205.7095, 200.5584, 205.5298, 196.558, 200.9058, 194.6199, 
    198.8224, 189.6818, 182.9379, 179.0433, 176.0473, 166.2269, 167.8445, 
    167.78,
  184.7233, 195.8312, 191.2898, 205.2937, 203.5549, 190.8419, 176.6682, 
    166.258, 163.1609, 163.4114, 162.5, 155.1787, 151.9681, 154.7532, 158.0946,
  200.022, 193.3197, 195.9277, 202.2185, 196.451, 189.8699, 181.7442, 
    172.3282, 167.4415, 167.909, 159.9196, 163.2513, 155.8603, 157.4274, 
    158.1145,
  201.2159, 198.2912, 203.312, 197.6499, 201.1906, 170.627, 185.5983, 
    174.022, 172.6525, 171.4199, 167.3178, 159.9857, 163.6272, 163.937, 
    163.6401,
  210.726, 202.0393, 209.5648, 205.1411, 203.255, 204.7584, 169.032, 178.09, 
    178.5542, 173.3483, 167.4994, 164.3115, 165.7402, 162.9797, 164.9045,
  216.2454, 212.5307, 199.1647, 203.931, 206.988, 209.2002, 204.23, 171.1328, 
    164.2349, 172.6315, 170.6471, 170.0926, 167.533, 168.3033, 169.2719,
  211.3516, 209.5372, 202.0083, 203.5089, 190.5234, 198.7406, 199.4697, 
    201.1189, 187.692, 178.8015, 173.9836, 172.0318, 169.8255, 170.5081, 
    171.135,
  210.6067, 205.5921, 208.4576, 206.919, 199.6504, 192.5153, 196.7047, 
    194.6034, 196.2474, 190.4058, 185.8932, 175.952, 176.5656, 173.8887, 
    174.6303,
  215.4309, 210.3895, 201.1946, 202.4957, 200.5618, 202.9854, 198.5481, 
    196.2984, 189.4414, 189.1752, 184.6711, 179.7362, 179.278, 176.5906, 
    179.7525,
  213.7549, 212.1475, 206.0556, 204.1759, 199.4206, 199.6671, 200.9135, 
    194.9045, 189.8655, 197.6914, 188.2903, 178.6505, 178.0285, 178.926, 
    178.8849,
  217.2834, 210.082, 208.3664, 204.8511, 199.734, 195.168, 194.8864, 
    196.0617, 198.2664, 186.7502, 186.24, 180.73, 180.5617, 183.3732, 184.4637,
  189.6529, 196.1631, 195.0582, 202.9131, 196.1674, 183.4075, 183.5612, 
    189.7891, 190.1398, 176.9493, 178.3311, 183.3206, 180.3806, 178.702, 
    168.7405,
  192.0303, 204.6477, 202.7372, 196.7122, 183.9797, 177.4079, 173.6509, 
    186.49, 189.1751, 182.0827, 180.9524, 186.2009, 186.3264, 173.3558, 
    172.2489,
  193.5036, 198.8956, 205.4256, 199.5666, 182.3115, 167.3545, 177.3315, 
    179.7782, 181.0047, 179.0688, 186.0652, 184.5729, 182.8174, 182.6535, 
    182.8483,
  192.5618, 203.5035, 206.7883, 198.4347, 186.7669, 178.7205, 167.3269, 
    176.7122, 175.3115, 177.5633, 182.7944, 184.0048, 181.6175, 180.6633, 
    185.6208,
  191.9871, 202.7338, 205.5755, 203.6465, 197.3231, 190.5532, 175.9481, 
    170.1742, 176.0128, 177.5989, 180.6221, 181.9673, 178.3699, 181.3714, 
    184.5762,
  188.7365, 194.889, 202.9477, 205.0181, 200.4332, 189.939, 174.4878, 
    168.9975, 181.8043, 187.5904, 181.6445, 179.0583, 176.2176, 176.8677, 
    183.0909,
  191.852, 191.8294, 198.1012, 205.9717, 201.8825, 189.0352, 181.4689, 
    170.9267, 173.006, 182.1028, 183.6269, 173.4653, 174.6311, 178.6035, 
    187.5443,
  196.8191, 200.2873, 198.2163, 200.2031, 196.425, 190.5728, 177.0167, 
    177.9075, 171.4627, 172.7506, 178.0359, 173.8857, 173.3276, 178.2831, 
    184.1537,
  195.8696, 199.3202, 201.0211, 196.7089, 192.886, 182.4494, 183.0689, 
    180.098, 173.5388, 172.5543, 172.9055, 166.4972, 168.6031, 171.1896, 
    175.5643,
  193.8489, 198.014, 201.3718, 199.5975, 191.0545, 187.8248, 180.3439, 
    182.5317, 180.0779, 176.3932, 171.9, 164.298, 160.4768, 166.2088, 171.9181,
  178.21, 189.6674, 193.4578, 190.1511, 186.7158, 178.1618, 184.3498, 
    191.1536, 191.4254, 177.2012, 178.1212, 179.4348, 173.3155, 174.8007, 
    162.3042,
  185.5631, 196.5712, 201.0572, 200.3667, 181.3515, 179.0037, 189.1129, 
    192.302, 193.1843, 189.1101, 182.0591, 185.0364, 187.4249, 169.6404, 
    164.0162,
  193.2972, 204.9, 212.5006, 201.6777, 187.9576, 172.5871, 191.0068, 
    191.9142, 192.4579, 188.8043, 188.8459, 186.595, 185.9883, 189.9301, 
    180.7668,
  206.7185, 212.9506, 214.8423, 210.1007, 199.5133, 192.1976, 180.6362, 
    195.2039, 194.4796, 187.8724, 187.6271, 186.9634, 186.7268, 187.7769, 
    186.713,
  208.4145, 216.6991, 208.2877, 211.8591, 211.0705, 204.2927, 199.106, 
    182.32, 181.3149, 186.5441, 188.1573, 187.9528, 188.7668, 190.919, 
    190.6857,
  212.7972, 214.187, 209.9382, 204.509, 210.2691, 208.455, 205.8527, 
    204.3872, 204.2013, 203.823, 191.3185, 189.576, 191.0996, 192.2801, 
    192.5249,
  213.585, 209.2566, 210.0099, 211.2687, 210.9932, 203.2493, 203.4936, 
    192.1752, 189.966, 187.8583, 199.4037, 193.064, 193.5826, 194.106, 
    195.1924,
  214.3189, 208.6735, 208.989, 206.1106, 210.7313, 205.0695, 202.3956, 
    182.2422, 181.2571, 187.5807, 199.9992, 195.6059, 195.5839, 196.2396, 
    196.5947,
  212.9668, 213.5696, 207.2896, 199.1766, 198.5658, 201.7014, 201.9837, 
    185.3644, 190.3381, 184.8422, 203.6237, 197.211, 197.2937, 195.6932, 
    196.8702,
  214.7295, 211.0367, 199.7714, 189.9033, 194.6543, 200.6186, 199.0499, 
    192.5262, 192.3605, 204.7978, 201.9819, 198.5388, 197.8454, 195.8987, 
    197.4881,
  183.8251, 184.5343, 185.6517, 182.2028, 185.2313, 185.8823, 192.1637, 
    189.0338, 186.1033, 176.9804, 173.1203, 176.1617, 168.8056, 168.8001, 
    159.3069,
  183.2041, 187.2525, 183.7998, 178.0948, 183.782, 193.5636, 193.6224, 
    191.0232, 188.1986, 184.6943, 177.2116, 182.8356, 184.6137, 165.2372, 
    157.7709,
  179.8858, 191.1798, 188.2583, 189.8261, 196.5146, 188.3292, 191.7613, 
    188.5183, 187.4629, 186.8656, 186.8172, 184.3006, 182.9824, 184.021, 
    173.2089,
  185.2762, 190.5429, 194.0299, 195.6798, 205.7625, 204.2292, 183.4012, 
    188.7171, 187.6075, 186.5285, 185.3798, 182.3423, 182.3359, 183.1618, 
    180.7804,
  192.4728, 189.3161, 192.6808, 195.5852, 205.5567, 207.6953, 208.2173, 
    179.2886, 176.6615, 182.9436, 184.477, 182.7782, 184.4384, 185.9309, 
    188.8512,
  190.6599, 193.4204, 201.6325, 207.1298, 206.4667, 206.5201, 209.3751, 
    213.3174, 201.2946, 198.39, 185.79, 184.5507, 185.1239, 188.2639, 190.2789,
  197.3387, 200.5914, 208.646, 210.0501, 206.5598, 201.4171, 208.5033, 
    208.4221, 194.0596, 182.8011, 192.4233, 185.4347, 187.6548, 190.7095, 
    191.9543,
  200.726, 203.6435, 212.7498, 208.8255, 210.5148, 202.947, 208.6291, 
    196.7516, 181.062, 180.3868, 190.2836, 187.4228, 190.1459, 192.426, 
    193.6748,
  196.3068, 210.7412, 215.6006, 210.2402, 207.7432, 201.9706, 206.0927, 
    194.6734, 180.1466, 179.0952, 193.2456, 190.0428, 192.7361, 193.9766, 
    194.1563,
  202.5395, 218.167, 212.6049, 210.0103, 204.8958, 208.571, 209.6059, 
    200.3778, 187.3386, 200.6711, 193.5994, 191.4284, 194.4434, 193.7843, 
    194.4785,
  174.8817, 179.179, 184.5674, 201.6878, 191.7131, 191.0393, 190.244, 
    185.993, 186.3615, 174.7225, 169.1858, 175.9149, 169.1531, 169.7152, 
    160.6719,
  186.1062, 182.6237, 190.2538, 198.4079, 191.7784, 192.8273, 189.9063, 
    189.7682, 188.7966, 185.2857, 174.2711, 184.7956, 186.6108, 166.05, 
    160.6142,
  189.5703, 185.3344, 199.7036, 203.1022, 190.5415, 187.7236, 192.1384, 
    190.1754, 189.0283, 188.0257, 189.0256, 188.5426, 186.096, 183.9939, 
    171.4182,
  193.7685, 196.7892, 201.871, 198.9587, 195.3203, 203.2772, 183.6691, 
    188.7187, 188.3186, 188.2539, 188.1181, 188.5257, 189.469, 187.2016, 
    180.6187,
  194.1763, 200.2747, 202.2044, 199.0602, 190.0157, 199.1076, 210.1085, 
    177.4644, 171.3307, 180.1859, 186.8474, 190.0231, 191.1842, 190.6071, 
    192.1458,
  190.4062, 205.7716, 202.8627, 194.291, 195.3471, 204.1333, 205.1304, 
    215.9129, 201.5482, 195.912, 187.2534, 191.6686, 192.7213, 192.9477, 
    190.2757,
  206.3174, 197.7324, 198.4649, 193.6992, 201.7589, 207.0463, 207.3078, 
    195.9633, 197.5324, 201.4737, 198.8005, 193.6389, 193.7423, 194.7128, 
    193.3201,
  209.7284, 198.1629, 196.9394, 194.0919, 200.5297, 211.1079, 209.5643, 
    212.9722, 191.923, 199.0704, 196.3184, 194.4492, 195.3504, 195.1813, 
    196.5733,
  206.5737, 199.5023, 194.3421, 196.5642, 201.8413, 209.2943, 213.4621, 
    211.9773, 185.4158, 193.9403, 195.4361, 194.786, 195.5128, 195.6523, 
    195.4365,
  201.3146, 197.7581, 194.9565, 197.9901, 199.4324, 209.8519, 208.6528, 
    208.4963, 197.4283, 196.1465, 194.9733, 194.8639, 195.4819, 196.2189, 
    195.1501,
  201.7088, 202.6943, 202.6483, 215.489, 195.8579, 189.8722, 192.7155, 
    189.0985, 181.0121, 165.3829, 162.0921, 158.5541, 158.9541, 160.5423, 
    156.686,
  197.6376, 202.911, 211.3022, 208.5738, 194.6554, 190.103, 193.2992, 
    189.5504, 181.3312, 173.0132, 163.4924, 165.4354, 167.8232, 159.7534, 
    158.4227,
  191.8219, 197.687, 197.4951, 191.5084, 202.3217, 186.0701, 193.2486, 
    190.1486, 182.838, 174.7247, 166.8676, 164.1086, 166.2188, 167.7323, 
    163.6642,
  182.0518, 198.2945, 197.1869, 191.0258, 195.9575, 202.5276, 184.3849, 
    185.6718, 183.7984, 173.6453, 166.6696, 166.9883, 167.4416, 176.4176, 
    172.5551,
  173.4191, 191.4585, 202.5588, 213.7998, 204.6155, 195.2953, 203.0484, 
    177.9341, 166.6492, 169.2371, 165.8742, 170.9322, 176.7742, 182.6738, 
    189.6656,
  169.7825, 178.2912, 192.2476, 213.0121, 210.2611, 197.866, 197.747, 
    201.2321, 189.1348, 179.0758, 173.6582, 176.9107, 181.7083, 185.5632, 
    192.8004,
  187.0834, 175.131, 182.3041, 209.444, 212.1446, 216.1978, 197.5943, 
    197.4542, 193.0072, 198.2351, 185.4937, 183.5379, 184.1958, 188.7384, 
    192.6646,
  193.9768, 184.5837, 183.5229, 202.2667, 213.6675, 215.1996, 208.9732, 
    202.4516, 195.9422, 188.9591, 187.6601, 184.8729, 186.9081, 189.4638, 
    194.0591,
  192.7118, 189.9535, 189.1092, 195.5499, 210.8157, 214.0344, 212.6297, 
    196.36, 201.9595, 194.3313, 191.6078, 190.0383, 188.0192, 187.7234, 
    191.2823,
  199.4868, 191.9271, 188.1425, 192.9143, 209.2627, 211.5701, 213.4476, 
    211.7982, 205.6748, 198.4872, 194.69, 191.7188, 192.1942, 190.0605, 
    191.2882,
  166.076, 184.9417, 188.6756, 206.9754, 193.3423, 182.0441, 180.8298, 
    177.7563, 178.0731, 170.7606, 169.3409, 172.1099, 167.9636, 170.9668, 
    166.2264,
  157.3606, 170.229, 190.9027, 194.6674, 190.2905, 181.2477, 184.5648, 
    174.7771, 176.5346, 176.937, 171.9126, 176.5008, 178.1026, 165.2915, 
    161.0782,
  161.5049, 166.1855, 180.222, 192.276, 199.2684, 180.388, 184.6894, 
    174.3119, 175.9337, 176.2188, 180.1569, 180.4059, 180.2237, 178.2646, 
    170.4398,
  161.9946, 159.9536, 177.5155, 188.1383, 195.1164, 199.9819, 171.9908, 
    174.0584, 174.1649, 172.5758, 176.6618, 179.9837, 179.0603, 181.2479, 
    177.5644,
  157.6088, 158.2175, 172.2316, 205.6689, 197.1091, 191.7651, 193.7255, 
    170.5627, 168.0935, 169.9499, 175.5994, 183.4982, 184.2977, 184.7478, 
    184.4049,
  164.2867, 159.3405, 173.7874, 211.0625, 193.44, 193.9403, 186.731, 
    175.4471, 171.7916, 174.3836, 178.7774, 186.2961, 188.4492, 186.1325, 
    188.307,
  196.1517, 167.1112, 177.6304, 209.1248, 214.1675, 192.6037, 187.5827, 
    175.9857, 174.5636, 176.0134, 181.7739, 183.5895, 186.7948, 185.6145, 
    182.9503,
  214.2456, 196.2383, 185.8192, 208.3351, 211.5965, 213.7927, 186.642, 
    177.4766, 169.4874, 171.4282, 180.9191, 183.4135, 186.4716, 183.5255, 
    183.9451,
  198.9928, 208.7713, 203.7015, 212.4762, 212.0638, 214.5126, 209.9119, 
    179.7587, 168.8001, 174.8251, 178.7294, 179.1827, 182.1116, 182.7077, 
    177.1404,
  182.6478, 194.3455, 208.2619, 208.5341, 207.5265, 212.2813, 207.3, 
    184.5354, 170.9606, 172.0572, 177.7166, 178.1848, 176.4654, 175.5421, 
    176.2809,
  173.2276, 161.3723, 163.0906, 186.7729, 183.1713, 179.2021, 183.9904, 
    181.3428, 182.7025, 168.8303, 168.565, 174.4652, 169.1282, 172.1268, 
    163.6497,
  182.9226, 165.5657, 167.0094, 182.0475, 180.4076, 176.1895, 183.5619, 
    186.3634, 184.8493, 184.1581, 173.3033, 185.637, 187.863, 164.2473, 
    160.6998,
  188.0504, 167.3659, 167.2691, 179.2697, 192.1143, 170.6736, 183.8467, 
    185.1459, 187.4739, 188.4836, 189.0277, 189.6186, 189.2434, 185.0499, 
    173.403,
  187.9035, 185.7293, 168.2432, 174.7856, 195.6918, 190.5326, 173.6239, 
    182.5948, 187.02, 187.3914, 187.8515, 188.5096, 186.4774, 184.2864, 
    176.346,
  190.1111, 183.7605, 176.854, 183.707, 187.0469, 189.8557, 193.5996, 
    175.6428, 173.6584, 180.2408, 186.7348, 186.6415, 181.9238, 182.8264, 
    183.3579,
  188.1999, 188.1763, 186.0405, 190.7193, 190.3402, 195.6658, 188.3818, 
    197.1132, 191.8534, 190.3849, 186.5618, 186.987, 183.0535, 186.3058, 
    185.0368,
  192.4191, 187.8146, 188.3535, 196.3148, 204.3493, 183.4546, 192.8885, 
    188.9318, 196.0884, 200.6286, 192.3218, 188.0825, 186.3844, 186.454, 
    183.5217,
  196.5435, 187.4131, 191.7962, 201.4636, 208.1957, 193.8644, 184.3074, 
    189.3703, 193.5583, 196.6341, 190.9362, 189.6597, 188.7623, 188.3534, 
    183.0527,
  205.3039, 196.6926, 200.926, 209.3853, 209.3591, 197.0709, 190.7253, 
    190.9836, 194.0313, 190.3247, 189.8556, 188.5905, 189.8682, 187.0935, 
    181.0382,
  204.9118, 204.2001, 207.2708, 210.8457, 210.3475, 207.9162, 195.489, 
    188.1134, 192.5571, 190.9594, 191.0692, 187.8173, 189.2667, 185.3636, 
    178.4503,
  188.934, 200.821, 187.4682, 188.3904, 180.5279, 177.7551, 183.7192, 
    183.4645, 185.1236, 175.8962, 175.3545, 175.9209, 172.4807, 171.9983, 
    165.5004,
  185.6548, 188.0735, 188.186, 186.9599, 178.8437, 175.9348, 185.044, 
    186.1467, 186.9168, 185.7652, 177.1852, 183.4397, 184.6355, 170.3863, 
    170.2388,
  189.6214, 182.3493, 186.935, 179.7603, 193.1126, 173.6465, 180.8497, 
    187.037, 185.3866, 186.3601, 185.8911, 183.614, 183.4504, 182.4693, 
    174.1892,
  204.325, 188.732, 180.4052, 182.8837, 188.1198, 198.7395, 175.5086, 
    180.3053, 186.7526, 184.7734, 184.1062, 183.3428, 183.4613, 184.7524, 
    179.8795,
  207.0408, 199.9482, 194.4389, 188.7801, 190.7837, 190.9457, 197.147, 
    173.9213, 170.3479, 176.6638, 182.4624, 184.2108, 182.2973, 181.6445, 
    180.6794,
  216.063, 208.2541, 208.0411, 205.847, 186.679, 193.1036, 191.6099, 
    199.6998, 195.131, 188.4659, 179.993, 186.4297, 184.4947, 182.995, 
    183.3602,
  209.2601, 211.9514, 213.3434, 214.3397, 211.5965, 200.2002, 193.0322, 
    192.9276, 195.49, 197.8728, 188.7867, 187.9631, 184.3412, 184.2043, 
    183.6076,
  219.4777, 217.632, 217.629, 211.1228, 210.0728, 205.7138, 206.6063, 
    191.665, 194.28, 195.976, 192.7955, 188.0094, 185.2325, 184.7254, 184.886,
  221.87, 217.9739, 214.9557, 208.5705, 211.2607, 201.9245, 206.2405, 
    209.702, 195.4254, 194.3584, 193.1107, 188.1396, 186.2349, 184.2061, 
    184.8286,
  193.0493, 217.2848, 213.7271, 211.1086, 205.2314, 198.696, 196.8908, 
    203.8765, 209.0978, 200.2059, 197.3472, 189.5519, 186.5868, 185.7033, 
    181.9763,
  191.539, 208.6926, 191.2934, 199.0369, 189.3, 182.183, 184.4153, 180.8613, 
    178.3468, 174.7244, 174.1073, 174.4007, 170.3137, 172.5731, 168.9137,
  191.4263, 200.5252, 204.6564, 207.5146, 182.6718, 179.0712, 188.1112, 
    183.3826, 180.7789, 177.5035, 172.105, 171.9558, 174.4845, 169.558, 
    167.9124,
  193.5044, 192.5537, 195.9114, 197.5862, 197.2098, 177.3335, 185.3286, 
    182.1664, 175.4053, 174.2233, 173.2455, 172.927, 172.3201, 171.3065, 
    166.4761,
  192.0758, 187.5826, 186.6785, 192.3, 198.9267, 200.576, 177.7638, 178.8467, 
    176.5012, 172.1426, 173.5802, 175.1517, 170.4685, 169.0404, 164.9067,
  194.0689, 193.2643, 186.9946, 187.5069, 191.2813, 198.9488, 198.717, 
    176.8536, 176.7901, 176.5642, 173.4284, 177.785, 175.0312, 176.6739, 
    168.1625,
  211.1549, 197.4732, 191.3837, 187.108, 187.3987, 191.5348, 198.3495, 
    197.0457, 184.6314, 176.1112, 174.074, 180.471, 182.4063, 182.3427, 
    176.337,
  217.2793, 215.8339, 203.0276, 210.2057, 211.3779, 196.0707, 199.542, 
    199.4352, 188.9895, 184.4576, 183.0769, 176.8983, 177.9009, 181.0144, 
    176.3956,
  200.0313, 198.7886, 201.3724, 203.3671, 208.6075, 212.3199, 211.5008, 
    201.5463, 189.8024, 187.4907, 183.9646, 179.164, 178.1839, 181.7654, 
    179.4436,
  173.2891, 174.6065, 181.6508, 193.154, 200.5069, 211.9413, 211.7699, 
    209.5006, 199.6327, 182.8431, 186.8041, 184.3533, 182.9286, 180.0809, 
    182.4582,
  173.8513, 172.1703, 180.5692, 185.2931, 190.5521, 205.7306, 211.4211, 
    211.3106, 202.129, 187.1164, 189.0537, 184.7108, 185.2221, 182.9504, 
    184.4198,
  190.2779, 206.9267, 191.9235, 198.3234, 189.8681, 179.9279, 184.1884, 
    184.4073, 183.0509, 176.7965, 171.0303, 168.1196, 164.9808, 164.3602, 
    162.6673,
  203.1012, 191.0945, 197.7007, 198.6754, 185.8931, 177.5896, 181.0383, 
    185.2747, 188.1756, 183.0195, 173.3847, 166.9397, 166.1354, 163.3392, 
    158.3423,
  193.5648, 189.0574, 194.1327, 196.0754, 193.8328, 180.3467, 180.3545, 
    183.4409, 184.9285, 184.7803, 180.0012, 173.9763, 167.3802, 166.1703, 
    162.1734,
  196.099, 189.8256, 188.8339, 193.5038, 201.4222, 196.3123, 172.3728, 
    179.2793, 184.1731, 184.6138, 181.6742, 175.1756, 171.5051, 166.0675, 
    157.3137,
  197.7281, 196.0939, 192.6023, 195.0307, 195.5399, 204.0678, 195.2647, 
    174.4324, 178.3878, 182.2867, 184.9639, 180.8918, 173.4573, 170.7905, 
    164.5887,
  179.1168, 177.528, 194.418, 199.8675, 202.9964, 203.3924, 196.2744, 
    202.1637, 190.0349, 187.472, 183.6829, 186.4576, 181.1109, 177.8504, 
    169.9155,
  177.3992, 178.0928, 173.5652, 186.4276, 203.5207, 213.2989, 208.1127, 
    194.1243, 205.2435, 193.1502, 192.5308, 189.2345, 186.8977, 181.6392, 
    175.2123,
  173.2111, 177.4987, 182.2862, 186.6988, 198.5153, 209.9547, 214.8831, 
    204.888, 192.6885, 194.421, 192.9108, 190.9265, 187.7727, 182.1708, 
    179.3132,
  195.7237, 203.7303, 197.272, 195.8132, 195.0307, 197.0305, 214.6418, 
    206.6343, 201.8808, 191.7219, 193.4454, 191.7779, 188.814, 186.5283, 
    184.8577,
  197.7352, 209.2023, 203.3156, 207.5623, 200.9688, 186.7694, 207.5675, 
    212.5427, 206.7309, 197.7148, 195.0233, 193.4537, 190.8465, 190.7657, 
    187.9041,
  189.1118, 202.6919, 191.2866, 196.9572, 192.7179, 185.1651, 191.1037, 
    191.1155, 186.4114, 176.1277, 168.8121, 165.7881, 161.5901, 167.7887, 
    167.8637,
  207.9876, 208.238, 200.9083, 201.2402, 188.4911, 183.5559, 189.7091, 
    191.1924, 188.0278, 183.9507, 171.5903, 171.1809, 164.9429, 163.6056, 
    169.2648,
  195.2335, 200.6788, 206.5734, 208.3878, 194.6127, 183.441, 188.8175, 
    190.1809, 188.7024, 187.4935, 180.8628, 173.1349, 165.51, 166.6562, 
    167.1033,
  202.9236, 198.7798, 198.6815, 214.0885, 207.8145, 193.9601, 185.9942, 
    184.9595, 189.5082, 188.6744, 186.0479, 179.3066, 170.8574, 166.3533, 
    163.9173,
  198.3771, 196.8521, 214.4223, 205.1841, 210.991, 215.3413, 201.7614, 
    179.8303, 178.5747, 187.5612, 189.6694, 184.1885, 175.774, 166.4607, 
    167.7899,
  203.1481, 195.9865, 216.1398, 215.1722, 213.4606, 213.3652, 205.2635, 
    210.0112, 194.218, 188.8678, 190.1746, 188.9659, 179.8946, 173.1909, 
    167.7636,
  214.9069, 216.7763, 202.1035, 200.5341, 211.5348, 215.7548, 207.3631, 
    205.3095, 202.3671, 198.5458, 193.8876, 190.8078, 187.234, 181.9306, 
    170.2581,
  206.0312, 215.9694, 203.3045, 207.0577, 216.7719, 216.5951, 211.1518, 
    204.3382, 205.6378, 194.9829, 192.2779, 191.1115, 189.7112, 184.6546, 
    180.631,
  212.9707, 210.7908, 221.9066, 219.5805, 218.6066, 217.9916, 214.9345, 
    212.5769, 204.237, 194.5401, 192.9726, 192.7673, 191.4551, 188.9988, 
    188.8947,
  190.3286, 199.8, 203.3082, 211.4465, 212.346, 217.4321, 214.3662, 214.9485, 
    211.8521, 196.6359, 195.3888, 194.658, 192.8974, 191.8474, 190.0191,
  165.2533, 178.4529, 177.2005, 181.4824, 181.7382, 182.6407, 186.3513, 
    189.8624, 190.8417, 187.8826, 186.1933, 184.4137, 179.7713, 173.6317, 
    166.946,
  175.509, 176.0062, 181.4209, 181.4068, 181.4524, 181.4847, 187.7519, 
    193.1375, 192.3437, 189.6066, 186.5142, 185.7233, 181.1935, 174.7439, 
    164.9356,
  187.9284, 190.0651, 188.3955, 189.7057, 185.6272, 179.5002, 191.8866, 
    192.9891, 192.0276, 191.0057, 190.7862, 186.4778, 180.1253, 174.0546, 
    164.8372,
  192.0261, 200.6218, 195.1545, 196.8809, 203.0953, 193.537, 189.1175, 
    193.379, 195.1037, 190.6804, 192.5102, 188.4762, 182.5804, 173.1547, 
    164.2885,
  206.6716, 204.9406, 204.091, 210.9838, 210.9729, 202.9218, 202.0164, 
    192.525, 189.4348, 189.1668, 190.9154, 187.522, 182.063, 176.5793, 
    168.8369,
  213.782, 207.8969, 212.7731, 214.654, 213.713, 216.1317, 213.8341, 
    210.5972, 203.0097, 189.767, 188.4258, 187.3327, 183.4897, 177.148, 
    167.7473,
  216.0424, 214.6789, 212.421, 215.6198, 216.2265, 214.869, 215.0583, 
    213.1655, 211.4482, 188.7411, 188.312, 187.4764, 182.8526, 176.1702, 
    173.6766,
  219.6542, 215.0727, 213.6823, 212.2219, 217.0063, 217.6018, 215.9996, 
    216.858, 216.4377, 198.8608, 188.7064, 188.224, 183.8566, 177.6899, 
    174.8143,
  216.0741, 219.6943, 219.4004, 218.9009, 214.6531, 218.4779, 218.6609, 
    217.8375, 217.5972, 209.9975, 198.9702, 196.4576, 188.4718, 176.656, 
    179.6082,
  219.1145, 218.3588, 219.5549, 221.2919, 218.4946, 218.156, 219.0985, 
    218.3952, 215.0217, 204.7028, 198.7357, 196.4281, 190.3377, 175.849, 
    172.676,
  169.2758, 165.2463, 162.6013, 163.7714, 165.0899, 169.1855, 173.6555, 
    183.9417, 189.3531, 187.2271, 186.282, 184.5567, 177.6854, 177.3265, 
    170.1574,
  174.0717, 167.1447, 165.6304, 164.1332, 164.2652, 165.5533, 172.9399, 
    183.6012, 190.4371, 193.1544, 189.9911, 187.0189, 180.6231, 176.817, 
    174.9484,
  180.8024, 169.2946, 164.2207, 164.7915, 166.3336, 163.7399, 171.4155, 
    181.7446, 190.1767, 192.5861, 188.0089, 184.1148, 179.9477, 176.2458, 
    177.2515,
  180.7212, 171.6034, 162.4245, 158.3489, 169.0285, 170.977, 167.5759, 
    175.1742, 184.8063, 187.1844, 184.9518, 181.3437, 172.6017, 172.3905, 
    178.8779,
  176.3234, 166.6619, 163.6437, 163.7082, 162.2913, 175.6711, 179.9435, 
    177.3138, 182.9214, 184.5158, 184.5133, 182.0537, 172.879, 169.7491, 
    180.0712,
  171.5766, 167.5782, 163.2173, 168.4171, 168.6897, 174.0273, 179.982, 
    194.973, 192.7306, 185.3004, 185.8874, 183.1784, 173.0467, 163.035, 
    172.3277,
  175.5389, 170.4462, 172.7724, 174.7863, 174.2304, 184.7669, 182.8113, 
    192.9625, 200.8519, 187.1605, 187.0488, 185.5979, 176.1782, 164.6527, 
    169.9735,
  184.2969, 180.6272, 181.4081, 185.0746, 184.0093, 188.5266, 197.3014, 
    202.1012, 208.9711, 208.9369, 200.5926, 193.5981, 182.9159, 164.9072, 
    166.6589,
  196.3732, 191.4736, 192.3886, 193.2507, 197.9694, 200.6913, 206.6003, 
    208.4176, 213.4786, 211.4764, 201.1225, 193.8455, 188.5177, 172.2649, 
    168.471,
  206.0662, 206.4526, 206.6734, 206.3634, 206.8135, 211.7848, 214.6548, 
    214.1902, 214.0784, 201.4858, 200.1131, 191.9208, 191.8499, 183.8163, 
    175.184,
  186.2418, 186.2841, 183.6533, 182.6848, 177.4935, 178.5286, 186.3084, 
    189.4813, 188.7428, 187.8136, 185.9529, 189.6053, 179.688, 172.3625, 
    157.814,
  196.2221, 196.816, 195.3049, 181.4514, 171.1182, 172.009, 181.5841, 
    187.355, 190.3468, 187.5449, 184.6568, 187.8333, 188.6687, 174.3643, 
    161.7683,
  202.1295, 195.6837, 179.8632, 172.5015, 174.6628, 165.9041, 173.3671, 
    176.2865, 186.3928, 185.028, 183.8764, 183.8559, 187.4793, 183.0415, 
    163.4868,
  194.6346, 187.0524, 173.8048, 170.1725, 171.652, 174.7365, 165.1047, 
    169.6508, 183.3181, 181.9808, 183.7155, 183.9138, 183.5579, 186.8924, 
    167.364,
  196.2689, 191.8822, 181.0731, 170.6799, 166.5229, 172.5234, 180.8582, 
    166.11, 179.7921, 176.493, 182.9961, 183.8551, 183.8965, 192.7905, 
    177.7161,
  201.0526, 192.847, 185.8321, 175.8838, 172.4556, 170.0161, 172.4615, 
    179.8232, 172.7159, 168.438, 179.1637, 183.6331, 184.3034, 192.5748, 
    182.206,
  211.3275, 200.0469, 184.5618, 171.5271, 168.4639, 168.4126, 169.4649, 
    177.5485, 174.387, 169.0289, 176.8016, 183.1974, 189.6668, 190.3488, 
    187.6776,
  203.4536, 195.3213, 182.404, 175.1599, 168.6779, 161.2367, 162.1138, 
    164.7289, 166.0221, 177.8747, 182.0099, 184.7293, 189.1575, 187.8921, 
    186.9809,
  194.2136, 191.8772, 185.8458, 171.7708, 167.0375, 161.8872, 163.3751, 
    164.9324, 168.2198, 179.0144, 188.7, 198.9432, 191.8923, 192.7713, 
    185.7705,
  193.3021, 184.7134, 179.7683, 170.3887, 167.1714, 159.6148, 165.2173, 
    166.7761, 173.555, 178.8953, 193.8543, 201.718, 199.077, 188.4205, 182.887,
  194.8262, 200.4311, 195.0319, 195.8924, 190.0945, 185.5752, 186.8303, 
    187.9595, 186.145, 181.1482, 181.1306, 180.4779, 181.0514, 170.5244, 
    166.1931,
  211.9855, 212.4895, 206.3439, 199.3666, 181.5332, 177.8288, 184.8847, 
    184.2905, 185.6841, 182.3524, 182.1743, 182.4543, 177.306, 177.3772, 
    167.542,
  212.8447, 213.2739, 200.5416, 199.4122, 190.2845, 168.1677, 177.3422, 
    178.2285, 180.4905, 181.6264, 183.1907, 183.668, 178.3122, 176.7221, 
    168.6892,
  212.2586, 203.4768, 188.5104, 183.0762, 189.4041, 188.3934, 170.5299, 
    166.6823, 175.9231, 179.1574, 181.3671, 182.6392, 179.6454, 176.489, 
    176.9953,
  204.0921, 192.088, 184.3533, 184.4099, 179.7171, 174.1815, 182.4747, 
    170.8789, 171.4262, 172.4639, 178.7619, 188.6771, 182.2159, 175.8059, 
    176.1615,
  192.868, 185.6618, 180.6396, 182.4153, 177.4951, 176.0919, 174.7869, 
    175.5098, 170.4958, 168.4687, 176.8392, 186.8061, 185.9138, 176.6085, 
    173.9448,
  187.9469, 182.9293, 189.7625, 182.4494, 179.0619, 178.9165, 177.9902, 
    172.704, 170.5662, 176.6267, 175.0379, 183.5256, 188.4028, 175.1901, 
    174.3503,
  186.7109, 184.7137, 176.9147, 178.0262, 179.0817, 173.8292, 175.9043, 
    173.5556, 173.6007, 168.0305, 170.0645, 177.0175, 191.1975, 184.6884, 
    171.8362,
  185.7611, 182.8329, 178.6387, 179.9008, 180.6966, 179.199, 176.5831, 
    175.6449, 171.9264, 168.3266, 169.0205, 171.7658, 187.2198, 197.5059, 
    174.3906,
  206.1961, 201.9148, 196.7274, 193.1594, 187.7871, 186.4101, 178.1886, 
    170.3633, 170.6319, 163.3091, 171.2311, 168.624, 178.6277, 197.2972, 
    173.9022,
  198.4365, 202.33, 197.3578, 196.6746, 190.6805, 184.2547, 190.6456, 
    187.7199, 186.4632, 182.2782, 184.6362, 184.0091, 173.506, 169.2287, 
    159.429,
  208.5546, 201.2317, 202.8913, 199.7446, 180.8575, 178.9517, 182.6068, 
    185.2363, 181.6768, 186.3224, 185.7745, 187.9847, 183.61, 164.275, 
    157.1149,
  204.0539, 197.5654, 196.9797, 198.3163, 196.074, 180.299, 178.021, 
    171.7178, 172.6866, 179.7681, 188.0078, 188.421, 185.7224, 181.0636, 
    169.165,
  196.9866, 198.0177, 196.3371, 194.5579, 194.9428, 189.3194, 180.8293, 
    169.1816, 173.1808, 176.8346, 185.056, 189.9918, 185.6719, 182.272, 
    175.9344,
  198.0096, 200.6001, 193.9093, 193.9494, 187.8861, 183.6682, 178.1486, 
    172.6183, 182.5368, 173.905, 180.1117, 190.7641, 184.595, 184.2305, 
    181.5503,
  197.1755, 193.4578, 193.0074, 185.2733, 185.91, 182.7886, 172.7478, 
    175.0358, 177.5299, 173.6591, 175.8212, 187.5528, 184.7809, 184.169, 
    183.0905,
  214.7843, 196.9034, 196.5821, 187.4521, 178.35, 177.3399, 175.3113, 
    179.7416, 179.805, 182.0367, 176.4297, 183.7932, 185.6361, 183.8808, 
    183.1911,
  191.6417, 184.0259, 182.0909, 176.5012, 172.7036, 176.6303, 181.3334, 
    186.3817, 193.1479, 186.8362, 178.1542, 182.8472, 185.5318, 182.0379, 
    180.9657,
  178.7415, 172.9741, 171.5943, 171.2801, 184.2493, 193.7505, 197.2864, 
    196.4104, 193.8369, 192.1252, 183.849, 179.2492, 186.3297, 182.757, 
    179.8451,
  175.7146, 178.2124, 189.5334, 199.4802, 206.5596, 206.6257, 204.4745, 
    200.8259, 190.8041, 189.206, 192.2515, 181.153, 184.6692, 188.1195, 
    179.6614,
  198.3133, 202.3608, 192.853, 197.0658, 193.6001, 188.8903, 187.6415, 
    188.9239, 186.8085, 170.7703, 166.9621, 168.8718, 162.7319, 162.7355, 
    155.4132,
  199.9964, 201.9128, 211.3546, 202.4641, 189.1576, 186.6713, 185.414, 
    187.2579, 189.8794, 183.3739, 173.1267, 178.877, 176.9809, 159.8787, 
    156.1708,
  194.9319, 197.8029, 202.7699, 208.2709, 197.2042, 187.6537, 183.5554, 
    176.7893, 185.6271, 188.4052, 185.6494, 182.4368, 179.3593, 175.2784, 
    162.7216,
  195.051, 194.8905, 199.6693, 195.8272, 205.8271, 192.2855, 179.9698, 
    182.3951, 188.7271, 189.9846, 186.8913, 184.0161, 180.9351, 175.839, 
    167.5706,
  193.4557, 196.4745, 195.5321, 189.2719, 194.4339, 190.4945, 191.0637, 
    184.0028, 188.941, 190.9426, 188.6937, 185.9256, 182.0762, 178.2221, 
    168.841,
  192.2419, 195.1391, 188.7382, 196.3601, 194.5855, 194.0226, 191.3609, 
    200.6403, 196.4115, 195.0711, 189.119, 188.2584, 184.0555, 179.6807, 
    171.2893,
  213.6053, 216.6031, 201.7092, 189.5748, 189.4432, 194.5253, 204.1782, 
    206.5475, 204.8182, 201.0106, 193.6968, 190.0038, 186.6519, 181.4342, 
    176.4589,
  220.7885, 211.7127, 190.6715, 184.2857, 187.3717, 196.774, 207.9901, 
    211.061, 206.8722, 200.0683, 193.6272, 191.7737, 189.7828, 185.3368, 
    177.5756,
  213.5569, 201.3064, 184.4688, 181.5368, 187.1048, 201.7882, 207.8099, 
    205.0501, 195.293, 193.3549, 193.2062, 192.5366, 192.5255, 189.3771, 
    179.4742,
  202.9296, 185.6923, 180.0671, 180.4313, 191.4523, 196.5375, 205.3776, 
    192.9335, 189.7696, 186.5182, 197.0189, 192.6759, 192.2541, 190.5428, 
    186.8102,
  189.4944, 197.8191, 192.874, 197.9619, 197.2111, 193.9381, 193.8143, 
    196.4439, 193.6008, 191.4528, 183.5755, 177.5059, 166.4829, 164.3737, 
    160.0684,
  202.0676, 202.2384, 205.4062, 203.5286, 194.3508, 193.8628, 194.9048, 
    198.1333, 195.7691, 197.541, 185.1947, 179.9506, 171.5597, 162.2416, 
    160.6941,
  194.0029, 195.8513, 192.6258, 194.4584, 200.1541, 192.2019, 193.9623, 
    192.1482, 189.1429, 189.6903, 187.7087, 182.6432, 174.6563, 163.1245, 
    159.8253,
  189.4022, 199.6018, 194.6466, 188.2378, 196.894, 193.9406, 188.7021, 
    189.1441, 189.9941, 184.7584, 183.68, 181.3032, 177.9266, 165.6406, 
    159.9864,
  196.4259, 199.7608, 196.2785, 187.0576, 193.0667, 184.8748, 187.8812, 
    188.3107, 192.6352, 184.4912, 181.8309, 181.0989, 178.6995, 163.827, 
    157.4989,
  212.087, 207.5476, 203.3911, 198.8126, 190.4983, 185.7838, 182.2111, 
    189.6783, 187.7343, 182.1647, 179.8853, 183.5388, 182.1395, 167.7111, 
    159.2271,
  216.8755, 214.4136, 210.9103, 200.9534, 189.8396, 184.5159, 186.511, 
    183.7677, 184.9241, 181.7896, 183.2433, 185.2811, 187.864, 175.5894, 
    162.3388,
  220.9754, 219.2921, 215.0511, 205.4892, 198.0127, 188.4801, 190.0009, 
    191.7361, 186.2218, 178.8327, 183.1956, 188.1859, 189.4162, 176.0858, 
    163.216,
  219.5797, 220.0316, 219.4546, 209.0383, 200.9991, 197.4437, 188.0664, 
    180.178, 175.6636, 176.4205, 184.0927, 189.9131, 192.2658, 184.9361, 
    163.044,
  222.7669, 216.103, 211.3195, 208.8976, 193.2335, 189.5139, 182.3237, 
    178.9765, 174.3038, 169.4682, 185.4081, 192.1393, 193.6432, 185.2891, 
    169.0737,
  153.3472, 162.5296, 164.9339, 170.3727, 173.1503, 170.8525, 170.516, 
    176.2973, 171.9738, 173.389, 173.8581, 176.4021, 168.9418, 165.4267, 
    160.2303,
  178.1378, 180.2607, 177.6008, 174.9805, 169.8706, 170.9018, 176.8314, 
    176.363, 177.059, 179.2044, 174.8219, 177.962, 168.7903, 165.2242, 
    159.1773,
  197.7071, 182.8584, 182.8479, 184.0473, 181.3797, 175.7322, 180.3107, 
    173.8244, 177.3938, 181.6133, 181.3444, 178.5832, 172.8096, 168.2126, 
    156.4176,
  191.4079, 183.7307, 186.3373, 196.3289, 196.8625, 195.2593, 179.9218, 
    184.3219, 180.3711, 176.1037, 184.1617, 180.4128, 171.4518, 166.3307, 
    155.315,
  193.9382, 200.3034, 207.1947, 203.6073, 203.5979, 196.033, 189.696, 
    182.198, 185.3183, 183.909, 181.3298, 178.1342, 172.097, 166.4096, 
    155.6296,
  206.5, 210.3633, 213.9089, 210.4296, 202.6017, 197.1974, 186.4321, 
    183.8294, 184.7466, 180.5215, 180.4179, 175.1759, 169.5288, 161.9444, 
    156.2621,
  207.5664, 212.5146, 210.1103, 199.6134, 189.1614, 191.4791, 185.9259, 
    185.1052, 183.4617, 183.0018, 175.7289, 170.1607, 165.5104, 160.9487, 
    157.0114,
  203.5136, 201.3331, 201.9566, 196.0707, 189.4582, 184.9046, 185.5128, 
    188.1687, 184.8209, 180.8178, 178.4627, 164.7238, 160.6022, 161.3341, 
    159.1743,
  201.5272, 193.7462, 190.299, 189.7858, 187.5457, 181.7655, 187.0465, 
    190.2728, 192.9836, 185.9024, 172.0347, 165.2719, 160.1821, 164.1456, 
    161.1334,
  185.2352, 184.3079, 179.3137, 186.6869, 184.5291, 188.7864, 191.4946, 
    189.9297, 191.7534, 179.4854, 174.2086, 165.3855, 164.9781, 167.0766, 
    161.816,
  193.9835, 195.4347, 193.9062, 193.0161, 191.3153, 191.4431, 191.1877, 
    190.057, 186.2222, 178.5727, 171.8582, 166.5643, 164.4466, 162.5044, 
    157.7741,
  211.1569, 211.9404, 213.9922, 203.1856, 191.1732, 192.7339, 196.1349, 
    190.9007, 184.4232, 173.1083, 163.8551, 163.8621, 163.6621, 161.2274, 
    155.0986,
  209.1981, 208.8561, 204.6883, 201.4523, 205.3879, 194.4271, 199.7494, 
    178.7084, 164.9818, 160.9671, 157.3644, 158.0455, 163.071, 163.533, 
    158.9816,
  204.6537, 200.3432, 200.6742, 197.8432, 203.5007, 206.9757, 188.8759, 
    173.3499, 155.1075, 150.8471, 151.2596, 154.9707, 163.5273, 165.1442, 
    163.5807,
  204.004, 205.6955, 199.6323, 204.5704, 198.5276, 192.5081, 184.6078, 
    172.3479, 162.1083, 150.6903, 148.1582, 159.2293, 169.892, 170.054, 
    163.2526,
  200.8267, 201.5223, 198.4015, 197.4085, 190.0678, 175.315, 166.8175, 
    153.8752, 153.3762, 155.2252, 157.5341, 175.231, 176.0594, 170.5038, 
    163.328,
  198.4407, 194.0272, 184.7698, 185.1655, 178.8489, 164.5555, 161.5624, 
    158.0942, 155.3404, 158.2511, 174.4962, 186.7164, 180.2653, 168.0059, 
    168.2823,
  190.8552, 176.5267, 176.1805, 167.9453, 168.393, 161.6864, 161.6671, 
    160.513, 167.3493, 176.8013, 186.577, 192.3339, 178.7278, 171.7121, 
    170.0065,
  181.7217, 172.0506, 170.6438, 157.8166, 163.8315, 160.6148, 159.0227, 
    164.9082, 175.2626, 183.2996, 188.8611, 190.3459, 186.4523, 177.4098, 
    169.6212,
  181.1813, 173.4784, 162.2457, 161.1062, 160.7365, 161.6879, 163.0975, 
    165.1094, 176.998, 179.414, 190.2444, 194.8649, 190.6905, 180.7194, 
    172.2895,
  189.1165, 199.1396, 198.1536, 196.8206, 191.2343, 191.877, 194.2181, 
    190.7916, 188.9005, 183.9791, 174.0448, 160.3396, 152.2369, 147.4534, 
    160.6581,
  188.8595, 200.1219, 207.6391, 204.7547, 190.9577, 197.1172, 199.2335, 
    193.7983, 191.6195, 184.0676, 171.5411, 162.0963, 151.741, 150.2903, 
    173.3407,
  176.9414, 184.774, 191.2454, 194.2811, 198.2547, 190.4045, 204.0444, 
    196.2632, 190.3715, 184.3643, 172.4596, 160.479, 152.6097, 164.5542, 
    183.6097,
  175.6193, 177.9324, 180.5417, 183.2904, 187.1977, 196.0927, 189.2478, 
    195.5163, 193.932, 185.6738, 171.5308, 163.637, 157.0104, 167.2382, 
    186.9925,
  170.2421, 169.8405, 170.1984, 174.1335, 179.0401, 178.3079, 184.7817, 
    180.0565, 187.3179, 178.4003, 168.5792, 163.3335, 165.2236, 177.4098, 
    185.827,
  173.4674, 170.3157, 171.0112, 168.1058, 168.6876, 165.5007, 171.7928, 
    174.1299, 173.177, 170.8677, 168.1661, 166.5713, 164.4486, 183.0667, 
    184.2491,
  174.3835, 172.8481, 170.7845, 173.4449, 173.9176, 171.645, 166.3259, 
    161.0625, 165.3654, 164.931, 167.783, 160.8358, 170.0369, 177.9919, 
    188.9279,
  179.8237, 180.9603, 184.6557, 186.8017, 184.3945, 184.7178, 173.8145, 
    168.8472, 164.1461, 165.686, 161.6862, 163.49, 171.5238, 177.5186, 
    184.1923,
  196.8211, 207.9463, 215.2351, 207.9642, 200.3037, 189.1441, 184.5355, 
    177.6167, 170.9522, 168.6292, 164.3853, 161.5715, 170.6037, 181.3272, 
    179.1474,
  213.9892, 219.8231, 213.9325, 203.8914, 191.2803, 185.9542, 181.4257, 
    176.5075, 174.2416, 169.7009, 165.6408, 161.8992, 171.9443, 182.2398, 
    180.3065,
  173.0043, 171.7373, 180.0117, 193.9452, 191.0222, 191.271, 194.7402, 
    189.5405, 186.5872, 177.1851, 176.1414, 166.2379, 158.1705, 151.8894, 
    163.7258,
  171.9753, 171.8735, 174.9962, 186.883, 189.8127, 197.3239, 198.9882, 
    192.3161, 189.8513, 184.768, 179.719, 171.5167, 161.4599, 151.8815, 
    166.6584,
  175.3174, 172.3201, 168.1729, 179.2893, 190.8561, 187.8643, 204.2561, 
    196.269, 192.2754, 188.1845, 185.5211, 175.1786, 166.985, 160.9124, 
    177.5961,
  176.8101, 172.4795, 166.7232, 168.0827, 179.6427, 197.4194, 186.2313, 
    198.3932, 196.4805, 191.6503, 184.8075, 180.1965, 170.1374, 165.5132, 
    182.9863,
  176.8221, 167.4477, 164.5184, 162.0576, 162.8466, 177.9813, 196.6335, 
    183.1945, 188.1461, 193.9529, 191.4148, 186.3446, 179.5371, 170.4291, 
    186.6782,
  191.5152, 171.8565, 165.1173, 162.8769, 164.3685, 167.2734, 169.5338, 
    189.297, 187.6538, 185.0505, 184.2298, 187.5463, 183.7334, 178.4741, 
    187.7953,
  209.1904, 189.2918, 168.4385, 160.198, 159.0061, 159.9008, 163.4924, 
    167.9121, 173.2945, 182.1081, 181.3336, 184.9075, 180.0045, 179.5552, 
    188.1044,
  223.4055, 210.0673, 187.9349, 172.2579, 165.1919, 162.4435, 163.843, 
    161.8414, 166.3418, 170.1346, 171.0543, 176.5931, 179.0768, 182.072, 
    187.9223,
  218.3782, 217.4454, 208.5655, 194.7637, 187.9887, 185.0271, 176.655, 
    175.8318, 168.238, 168.4006, 167.1225, 165.9649, 176.4486, 178.8705, 
    184.8378,
  213.0721, 214.5636, 204.4108, 202.9416, 196.6358, 193.7866, 190.3804, 
    189.3169, 182.5971, 174.866, 167.6769, 160.908, 172.3004, 174.9701, 
    184.6366,
  174.226, 173.7092, 175.3793, 187.8489, 186.7557, 190.4792, 193.5173, 
    186.2728, 183.4426, 174.4716, 170.4035, 171.2718, 165.827, 165.6843, 
    161.3136,
  174.3027, 180.8568, 185.5477, 191.7577, 186.5282, 195.6215, 195.2847, 
    188.1021, 185.7478, 181.5081, 174.1823, 179.3985, 176.1113, 162.2484, 
    159.8541,
  182.9073, 182.2676, 198.9533, 203.5592, 198.0123, 188.122, 197.3589, 
    190.1315, 186.9606, 184.0933, 183.463, 178.6331, 177.4741, 174.5299, 
    168.5569,
  173.2727, 180.2356, 191.7766, 195.0783, 217.364, 209.0488, 187.7279, 
    192.4384, 189.7396, 184.7529, 182.5898, 181.0487, 180.4701, 178.5933, 
    176.0029,
  174.3616, 174.981, 183.975, 190.6678, 198.2263, 218.0876, 216.7689, 
    185.3404, 182.7288, 188.6602, 187.767, 186.193, 180.4914, 180.7072, 
    184.1138,
  171.1583, 170.7266, 177.8987, 187.1908, 190.536, 201.0586, 215.8463, 
    218.0311, 200.3532, 193.1721, 191.5662, 191.5871, 184.3368, 183.1961, 
    183.7815,
  177.0586, 165.4442, 170.0357, 176.9415, 186.8708, 193.5122, 204.6136, 
    210.7657, 213.4549, 202.8059, 196.2174, 191.0216, 186.0342, 186.0749, 
    185.2253,
  186.9747, 172.6884, 167.8805, 168.2531, 178.7767, 184.8073, 190.7353, 
    198.327, 199.1413, 201.6906, 196.0451, 191.5428, 190.038, 186.7048, 
    184.6086,
  193.7421, 181.5769, 174.5547, 170.4774, 172.0788, 176.0258, 180.7731, 
    183.8956, 189.6388, 200.2272, 192.223, 191.6749, 191.4616, 187.3901, 
    183.7181,
  198.8093, 199.1425, 189.3396, 177.7165, 173.972, 173.1108, 176.6228, 
    180.585, 183.5295, 188.7572, 193.2247, 191.2735, 192.2253, 190.0414, 
    186.3558,
  191.4523, 194.877, 188.9674, 188.8836, 186.9893, 187.7108, 191.8572, 
    182.987, 183.3859, 172.4389, 168.858, 171.173, 166.7355, 168.9818, 
    165.3349,
  200.4228, 197.008, 196.7599, 192.8029, 186.7012, 190.5902, 189.0764, 
    184.3944, 182.3049, 180.5838, 174.6865, 179.7727, 180.1466, 164.9603, 
    162.2336,
  211.6138, 204.1566, 205.0653, 199.2075, 196.9643, 181.0085, 187.3661, 
    183.8012, 182.8223, 182.4568, 184.4734, 180.247, 178.4912, 178.1351, 
    169.1747,
  205.2451, 201.1271, 206.0682, 212.6165, 214.3631, 203.6098, 178.3907, 
    183.0455, 183.1804, 182.6989, 182.0114, 180.3459, 179.0313, 178.6443, 
    176.5701,
  190.6794, 195.5198, 203.6477, 208.2529, 215.0573, 214.3768, 212.0152, 
    178.653, 173.2293, 179.5543, 184.2051, 183.6625, 181.1855, 182.1426, 
    182.9749,
  188.7524, 188.026, 199.8544, 201.8757, 214.9886, 211.9271, 215.0909, 
    211.9131, 197.8357, 189.7394, 186.2969, 188.4028, 183.8386, 182.696, 
    181.3596,
  179.5586, 183.3569, 197.1217, 204.3035, 211.6056, 208.6309, 209.0157, 
    214.9004, 211.7189, 200.6723, 194.2259, 189.7124, 186.3906, 184.5111, 
    182.1139,
  179.7699, 182.4229, 197.9197, 211.2712, 212.9184, 212.8874, 205.2758, 
    201.1329, 200.8494, 200.8281, 193.0845, 189.5054, 188.4359, 184.8657, 
    182.0146,
  172.2781, 180.0896, 196.5966, 210.1201, 206.4706, 204.8093, 211.0178, 
    208.5628, 203.2354, 199.9059, 193.5956, 191.1036, 190.0223, 185.9972, 
    182.0577,
  172.7432, 180.9424, 195.1625, 205.847, 196.9971, 205.0667, 200.0922, 
    197.488, 205.2673, 197.5632, 199.2826, 193.4229, 191.5241, 188.4516, 
    185.6316,
  183.6155, 186.883, 178.7236, 179.7959, 184.1502, 184.3273, 187.4774, 
    181.9222, 184.4205, 175.6584, 174.1519, 178.798, 175.7397, 174.7343, 
    171.6342,
  189.4834, 186.0762, 183.2206, 183.6286, 184.4469, 183.0422, 183.8428, 
    181.3985, 180.887, 184.5557, 178.9971, 184.1733, 186.1787, 172.496, 
    169.2006,
  200.5318, 193.1449, 191.9442, 195.5059, 196.7336, 174.9945, 181.4867, 
    177.9786, 178.0687, 183.3763, 185.753, 183.9774, 184.7134, 183.3227, 
    173.896,
  201.7761, 194.4471, 192.7186, 210.5842, 214.1496, 199.495, 171.3894, 
    176.0189, 176.7251, 181.4928, 182.951, 183.0216, 183.3402, 183.1775, 
    178.4046,
  193.3799, 188.6629, 199.8605, 212.2552, 218.7214, 206.5946, 194.2186, 
    173.2717, 167.5683, 177.2692, 184.0219, 185.1105, 182.4613, 185.0729, 
    183.6841,
  194.3347, 196.7087, 193.5658, 213.9323, 219.6339, 208.7191, 194.9735, 
    194.4725, 192.3898, 189.5458, 184.2537, 187.9522, 185.3064, 184.7746, 
    182.8128,
  203.8227, 212.8628, 213.3336, 210.2157, 209.5909, 205.7026, 205.4434, 
    205.8891, 207.2284, 200.0319, 192.9757, 189.3607, 186.847, 185.8918, 
    185.3273,
  215.6507, 215.4161, 218.2705, 217.9305, 207.7403, 195.4014, 202.7187, 
    207.7191, 209.8561, 197.497, 191.8386, 189.9294, 189.0816, 185.6151, 
    184.0702,
  215.5389, 219.2113, 217.6764, 214.8607, 210.4617, 201.0638, 202.6569, 
    212.0387, 208.5573, 195.2643, 192.2273, 192.2111, 191.6046, 187.7214, 
    185.9819,
  214.351, 216.5083, 215.0208, 212.5471, 209.419, 204.7521, 200.6383, 
    201.3004, 200.2381, 191.7247, 196.9601, 194.6843, 192.9724, 190.856, 
    187.9057,
  181.7213, 195.8928, 193.1602, 194.5111, 188.1861, 185.1388, 188.748, 
    185.7639, 186.8969, 177.8025, 174.481, 174.8196, 171.4453, 173.725, 
    174.3334,
  184.2675, 201.5151, 203.5131, 194.6415, 184.9451, 182.3143, 185.9649, 
    183.7809, 183.1386, 181.4378, 174.905, 174.0084, 175.9677, 173.0198, 
    174.09,
  189.0346, 204.7656, 210.7811, 200.2444, 197.8706, 174.0996, 185.3045, 
    182.3377, 178.4605, 176.3711, 175.3629, 172.7123, 174.3217, 177.5799, 
    178.3447,
  188.9248, 202.2532, 215.7323, 211.9905, 212.0578, 201.0593, 173.1058, 
    182.1985, 179.6736, 174.2623, 171.2354, 169.8906, 172.5474, 176.1421, 
    179.618,
  183.7342, 194.2949, 211.3244, 211.1665, 214.4812, 208.505, 205.6532, 
    176.1261, 178.106, 177.3061, 173.1408, 171.8656, 173.9899, 177.7859, 
    180.4816,
  177.5148, 193.8829, 206.3459, 207.157, 213.1353, 209.5508, 205.7912, 
    200.7652, 184.891, 184.7812, 175.576, 175.7761, 173.4363, 175.4045, 
    178.705,
  176.6763, 185.5393, 189.023, 204.1786, 206.5079, 204.7169, 206.7396, 
    201.0054, 198.9392, 192.5531, 182.2859, 178.2471, 175.2876, 175.6396, 
    177.6632,
  172.7525, 190.1222, 198.2178, 199.5094, 199.5536, 196.4691, 199.084, 
    208.2099, 205.7448, 194.0135, 188.2792, 183.6326, 181.7716, 178.3152, 
    177.0345,
  172.4729, 185.8739, 205.8303, 208.3937, 198.1143, 190.0565, 197.4044, 
    204.8541, 208.8704, 198.084, 195.3475, 190.8644, 185.6201, 181.4451, 
    180.4616,
  178.6779, 188.0746, 206.7685, 211.9832, 206.5609, 188.8045, 196.005, 
    202.2576, 200.4702, 196.1644, 199.2428, 195.3363, 190.7352, 186.2399, 
    184.2978,
  193.6615, 198.046, 191.3411, 193.7809, 188.0198, 184.74, 187.4393, 
    186.8427, 187.475, 177.315, 174.6763, 177.4551, 176.6796, 177.3021, 
    172.4327,
  204.8925, 202.5065, 201.1731, 193.8773, 185.2501, 181.8757, 185.4863, 
    186.558, 184.9431, 184.8285, 178.7294, 183.0846, 183.7694, 173.3228, 
    168.6955,
  205.0101, 202.185, 203.0231, 196.5565, 192.4316, 173.7433, 182.5883, 
    181.1636, 182.1831, 182.8658, 183.7023, 184.2014, 183.47, 180.6591, 
    175.3649,
  200.6576, 200.3941, 198.207, 192.1689, 185.2926, 175.9664, 173.0143, 
    176.6536, 180.5058, 181.7962, 183.4835, 184.5518, 183.7963, 184.1476, 
    181.5623,
  197.0143, 194.1781, 190.5018, 184.6711, 178.6877, 169.2953, 171.1375, 
    172.9538, 177.8391, 181.9554, 184.4601, 188.9794, 187.095, 188.3465, 
    185.7906,
  196.3148, 192.0714, 187.8259, 182.62, 179.017, 180.5146, 177.7933, 
    179.3923, 184.4324, 186.9946, 187.3797, 192.1851, 191.6176, 188.1638, 
    185.5548,
  202.933, 196.7691, 192.3923, 184.5956, 179.6826, 179.3493, 180.4668, 
    180.5308, 185.0113, 185.9227, 189.9478, 192.9423, 192.6573, 187.5946, 
    184.2321,
  208.7392, 197.175, 192.9355, 189.9849, 187.7627, 184.3719, 184.3187, 
    184.1891, 186.8693, 185.7943, 187.1693, 190.1848, 190.8249, 188.1092, 
    190.444,
  213.3862, 209.6021, 215.9852, 192.5348, 191.3121, 190.4923, 190.2818, 
    189.8109, 186.6438, 185.2873, 185.0495, 184.6613, 179.2652, 185.2687, 
    184.0035,
  206.2672, 209.3208, 211.471, 197.9399, 195.0805, 193.9385, 192.9729, 
    195.4935, 187.392, 190.7573, 187.3557, 183.9469, 180.8974, 179.1785, 
    178.3268,
  189.7838, 192.4921, 184.0575, 189.058, 184.1556, 181.7685, 184.4979, 
    187.2234, 188.6491, 192.1171, 191.5202, 190.4724, 180.867, 178.4074, 
    174.4711,
  199.7157, 197.9028, 194.1885, 187.7502, 178.2681, 178.5197, 181.3391, 
    184.5654, 187.1655, 190.0006, 184.2255, 180.3544, 177.4215, 173.8859, 
    172.7713,
  199.1261, 203.4028, 202.4711, 193.5291, 188.8161, 171.2806, 177.5103, 
    177.2629, 181.325, 177.6391, 172.5046, 174.3574, 175.4242, 174.5335, 
    175.7656,
  195.0494, 200.2965, 194.1044, 196.0038, 193.4257, 186.0077, 170.7738, 
    176.29, 175.9639, 171.0777, 170.7299, 172.2955, 170.7483, 176.6958, 
    176.2381,
  192.1901, 189.9599, 186.5612, 188.5769, 194.5298, 189.2774, 190.5614, 
    175.122, 166.6527, 166.4098, 166.8294, 167.9368, 168.8698, 176.7465, 
    181.8684,
  191.4094, 184.9544, 182.7028, 183.4969, 186.6073, 189.7722, 188.2233, 
    183.0965, 176.2375, 171.6458, 166.0624, 167.9887, 170.3061, 175.4221, 
    185.8347,
  177.6781, 183.1834, 185.2181, 185.0586, 188.0355, 190.5729, 192.111, 
    182.171, 177.2255, 172.0433, 168.6484, 168.9583, 172.802, 179.7758, 
    188.2496,
  178.5495, 177.8623, 180.0632, 189.6208, 192.7448, 198.0733, 189.8246, 
    183.3239, 179.9694, 176.6782, 168.088, 168.2183, 174.3936, 184.8563, 
    189.0553,
  180.4996, 177.3455, 182.4762, 189.3645, 194.5961, 196.5651, 192.6966, 
    186.4068, 181.4233, 172.6552, 169.5232, 170.128, 173.9651, 185.3082, 
    190.5813,
  190.3352, 191.0338, 194.2709, 192.6325, 195.1435, 196.3162, 193.3251, 
    184.4517, 179.9957, 173.8134, 173.0538, 172.4844, 178.2707, 186.4831, 
    192.058,
  184.0011, 190.1458, 185.5066, 192.0797, 185.5515, 187.5529, 189.1314, 
    188.4082, 190.2542, 184.8807, 186.7612, 190.2979, 187.5332, 184.2947, 
    179.891,
  194.5829, 195.151, 194.4393, 192.16, 184.3461, 187.5128, 189.7784, 
    189.1936, 188.2545, 188.0604, 184.5069, 188.639, 189.7836, 180.0554, 
    178.34,
  194.8192, 194.3008, 198.621, 196.1927, 191.698, 187.7841, 190.0387, 
    187.1541, 185.3528, 184.7411, 188.746, 189.419, 190.3109, 191.3601, 
    184.6953,
  186.8414, 187.134, 189.1374, 191.4109, 189.866, 191.3793, 187.6022, 
    185.5372, 179.111, 180.588, 182.1594, 185.416, 187.9262, 189.2903, 
    189.3836,
  180.1524, 186.292, 181.8226, 183.4068, 186.8555, 187.8641, 192.5138, 
    178.5129, 172.8776, 176.2587, 180.3398, 184.4538, 187.9694, 190.5872, 
    190.7588,
  186.945, 185.9155, 186.4963, 180.184, 184.2965, 188.1466, 182.1671, 
    175.9793, 175.0591, 178.1543, 178.5147, 184.4614, 189.6466, 190.3737, 
    190.7692,
  197.1106, 184.2548, 181.775, 176.8723, 182.6404, 185.286, 179.543, 
    167.5047, 170.8187, 175.5381, 180.9978, 186.4739, 190.2431, 189.767, 
    190.1047,
  193.3516, 190.8282, 180.6833, 182.2506, 182.0594, 178.241, 171.458, 
    165.6688, 168.5853, 176.9563, 179.6596, 186.0811, 189.9815, 189.8238, 
    190.1864,
  186.4531, 195.1767, 182.679, 185.3985, 182.8993, 178.2176, 169.7039, 
    164.8071, 164.5462, 169.3711, 171.4186, 184.396, 189.2061, 189.5989, 
    190.6674,
  190.7117, 191.5193, 187.8814, 185.4689, 183.1621, 182.3788, 170.2858, 
    163.6579, 161.4396, 162.7649, 172.3977, 179.3494, 187.8633, 190.2466, 
    191.9059,
  183.81, 192.2092, 179.4305, 176.2797, 170.0126, 170.5082, 177.2402, 
    183.5609, 189.8173, 189.5783, 187.6196, 186.4028, 182.6086, 178.6495, 
    173.3182,
  199.5395, 198.8638, 195.3278, 180.8607, 169.2387, 170.3681, 176.4356, 
    185.1772, 190.7498, 191.7815, 189.5671, 190.4663, 190.5412, 176.3493, 
    173.5064,
  216.1432, 202.662, 202.8724, 187.8491, 178.7561, 169.4633, 177.2818, 
    185.9002, 190.8141, 190.9365, 191.8882, 189.213, 188.8994, 189.5668, 
    181.4555,
  205.5648, 198.5452, 196.2006, 192.9586, 180.4125, 176.6387, 174.3305, 
    182.3283, 189.9989, 190.4409, 188.1295, 185.4015, 185.4718, 185.5125, 
    186.5947,
  201.5891, 214.4656, 211.1084, 195.0356, 184.4937, 179.0104, 185.202, 
    176.1729, 178.397, 184.8009, 185.9049, 184.4273, 184.5133, 186.1711, 
    187.4643,
  195.9348, 210.4459, 208.1397, 203.946, 192.2815, 179.7162, 181.0757, 
    196.4434, 197.3809, 194.6633, 185.9625, 184.5714, 184.3345, 185.1022, 
    185.9084,
  199.3089, 209.1952, 212.8332, 213.8449, 209.1742, 186.851, 179.1143, 
    190.1855, 195.2004, 193.1187, 189.2471, 185.4999, 184.7785, 184.2248, 
    185.0802,
  206.3103, 198.8073, 210.074, 209.437, 206.5927, 183.4142, 175.1222, 
    185.1892, 194.6791, 190.4868, 186.8972, 185.0007, 184.1116, 182.8951, 
    184.0399,
  201.4758, 192.5716, 201.3339, 208.5398, 204.9791, 188.8174, 176.989, 
    177.972, 189.7123, 187.4151, 185.9045, 184.8194, 182.9433, 182.9662, 
    184.1239,
  199.001, 184.7259, 188.4149, 202.0248, 205.1451, 188.186, 175.6545, 
    178.7069, 185.5152, 187.7138, 189.7325, 186.1385, 184.0986, 183.804, 
    183.3752,
  185.2715, 192.6319, 186.0857, 185.2472, 177.3334, 175.7768, 182.5788, 
    183.3665, 183.0627, 172.0358, 170.942, 179.5115, 180.8765, 172.6329, 
    165.6677,
  191.8002, 197.9002, 196.536, 188.527, 174.7984, 173.004, 181.765, 184.8028, 
    182.7025, 182.4227, 175.521, 182.9742, 186.2656, 170.4446, 165.881,
  199.4068, 205.3376, 207.2247, 196.7202, 181.6298, 169.6892, 178.2972, 
    183.6144, 183.6794, 183.9042, 183.516, 183.8793, 185.6754, 185.6741, 
    177.0113,
  187.4877, 196.952, 201.6185, 197.2723, 193.7216, 184.3435, 171.1503, 
    181.5565, 185.4904, 184.5421, 182.2552, 181.5976, 183.1473, 184.5173, 
    182.5516,
  177.299, 187.2764, 209.6947, 210.3493, 198.4312, 188.9372, 188.2046, 
    174.9776, 173.1912, 182.6593, 182.1205, 181.2908, 182.3511, 183.9216, 
    184.5588,
  166.8648, 189.2411, 202.6355, 213.2393, 215.2116, 195.8716, 188.3834, 
    196.1351, 193.6355, 193.7698, 186.3372, 183.078, 182.2228, 181.9905, 
    183.0242,
  165.2561, 189.2827, 202.1444, 206.4252, 215.1063, 203.8137, 194.1149, 
    188.2348, 189.9771, 192.5319, 189.039, 184.0099, 182.9106, 181.8342, 
    182.8427,
  179.3326, 186.5064, 195.9398, 200.7243, 205.1757, 207.9202, 194.1519, 
    186.5748, 188.0854, 187.9611, 187.1273, 184.3461, 182.9546, 181.6173, 
    181.7536,
  182.7208, 187.2477, 191.9195, 196.2721, 200.2917, 204.6595, 199.8637, 
    189.8464, 185.8597, 183.8984, 185.1208, 184.3305, 182.8548, 181.4494, 
    182.2802,
  182.4231, 184.7164, 184.0787, 191.0428, 199.0865, 200.7153, 195.7757, 
    187.9166, 183.8364, 182.4843, 187.3459, 184.7582, 183.4005, 183.4628, 
    182.9584,
  160.7696, 168.2033, 174.7543, 184.5515, 187.6063, 183.6973, 180.9739, 
    179.9174, 178.0426, 165.0125, 164.6252, 169.9594, 169.318, 165.9119, 
    159.9372,
  161.1606, 162.7562, 173.5098, 180.1268, 183.3852, 180.773, 181.0321, 
    179.4662, 176.8211, 174.9496, 168.4965, 176.3308, 179.9657, 162.9606, 
    159.9603,
  160.6807, 158.2667, 168.7054, 177.0484, 186.5096, 174.1678, 179.9176, 
    179.05, 176.2417, 176.2727, 176.9124, 178.198, 179.2894, 178.0894, 
    168.7063,
  159.6525, 157.2713, 163.305, 172.9014, 191.7647, 194.4458, 172.2727, 
    177.6585, 177.4691, 175.2641, 176.2605, 177.5812, 178.9767, 177.7379, 
    172.6407,
  161.082, 157.4058, 159.5945, 169.708, 188.3278, 198.2341, 202.0635, 
    171.8451, 167.9776, 175.3985, 175.5549, 177.9821, 181.3066, 180.8059, 
    175.2428,
  163.8017, 160.2509, 160.4445, 163.7538, 178.4066, 195.9815, 195.8282, 
    201.5042, 192.3412, 190.3525, 182.9935, 180.1291, 179.6023, 179.0416, 
    175.7888,
  180.8083, 174.5976, 167.3491, 160.1775, 176.4186, 193.7973, 202.1306, 
    196.8275, 193.1261, 192.5486, 187.4941, 180.7532, 179.4657, 179.8012, 
    177.3868,
  174.3613, 171.3915, 164.9117, 164.3994, 169.3242, 191.0569, 201.0918, 
    201.8215, 198.0089, 190.5064, 186.7572, 182.9666, 179.7763, 178.814, 
    177.3264,
  178.2391, 172.6751, 169.4738, 163.0239, 166.5253, 176.1024, 192.0115, 
    201.4451, 198.6069, 195.2388, 190.4303, 187.0963, 182.2645, 177.9681, 
    177.2734,
  180.1445, 171.8622, 168.9377, 165.4529, 164.4344, 168.858, 175.8394, 
    186.6412, 188.6385, 194.1017, 192.5347, 189.5122, 186.0781, 183.5708, 
    178.9665,
  172.7105, 171.013, 168.1794, 167.8967, 163.4906, 169.0422, 176.4349, 
    178.5678, 176.3661, 163.7409, 162.6645, 168.3547, 165.8123, 165.247, 
    157.4241,
  172.9319, 171.0119, 170.8714, 168.799, 162.9783, 167.9005, 177.1131, 
    177.7816, 173.8795, 167.7878, 166.1994, 174.5796, 175.8729, 161.7503, 
    157.8817,
  173.1839, 170.7466, 179.8717, 171.0692, 166.1791, 163.8876, 176.2432, 
    176.9522, 171.7772, 168.8341, 170.9987, 174.3366, 176.0363, 176.0501, 
    169.5111,
  175.3279, 176.2291, 174.8303, 183.4836, 174.0567, 178.1009, 168.7421, 
    174.355, 171.6029, 163.4464, 167.1507, 169.1012, 172.9753, 174.2393, 
    171.6865,
  177.4659, 177.274, 175.0711, 171.4964, 176.5712, 187.0158, 191.7296, 
    170.3708, 165.7416, 165.9286, 164.4967, 168.2312, 171.0267, 174.0667, 
    173.3419,
  182.1756, 178.0024, 187.2613, 186.7654, 174.8166, 179.9364, 203.5338, 
    199.9397, 189.1569, 178.9454, 170.5795, 170.0508, 171.9428, 170.9724, 
    170.0706,
  182.6353, 179.546, 183.438, 183.7675, 180.8604, 176.552, 203.6301, 
    201.7583, 195.3739, 185.1497, 175.1388, 169.1233, 170.8676, 170.2886, 
    171.7896,
  189.6633, 176.854, 177.9618, 188.6273, 190.4259, 178.8497, 185.3236, 
    202.5344, 199.422, 185.4647, 175.5232, 169.9192, 169.7804, 170.9393, 
    169.7312,
  190.1446, 177.1702, 174.2009, 182.2984, 185.8141, 187.6646, 180.5325, 
    188.544, 195.4005, 186.9103, 181.4668, 174.0757, 171.9969, 169.8589, 
    169.4613,
  196.5093, 180.4438, 176.5299, 180.9852, 183.9937, 192.9175, 188.472, 
    200.8427, 192.5629, 189.521, 189.4718, 181.3754, 177.0409, 174.57, 
    172.8329,
  191.1314, 186.0858, 178.2341, 171.78, 169.3315, 168.35, 172.7629, 172.4496, 
    172.8654, 162.974, 162.344, 163.9885, 160.448, 160.6003, 155.4696,
  191.3018, 188.4957, 180.8428, 173.2546, 168.7653, 169.4185, 172.077, 
    173.9566, 172.6877, 169.519, 165.0847, 171.2766, 171.2203, 157.3017, 
    154.1853,
  193.4494, 189.4702, 181.43, 171.9501, 173.1947, 169.3873, 174.5515, 175.47, 
    172.4792, 169.3426, 172.4804, 172.8482, 172.5421, 170.7704, 164.1956,
  194.7932, 193.1214, 182.4025, 178.6543, 172.2573, 177.1042, 168.1005, 
    173.2547, 170.9781, 168.4058, 170.5358, 172.2842, 171.7785, 170.3385, 
    167.9155,
  197.3885, 195.6236, 187.7349, 180.6966, 185.9074, 175.4245, 192.182, 
    167.6088, 162.4939, 166.0145, 170.4191, 172.8645, 171.7757, 170.0492, 
    169.183,
  204.2597, 196.6863, 188.6802, 178.229, 183.6552, 182.311, 195.4764, 
    197.0228, 185.8171, 178.866, 175.0182, 175.3308, 172.9148, 168.8975, 
    165.3789,
  208.326, 205.1787, 192.4909, 174.5362, 190.7074, 183.7381, 196.2157, 
    199.4155, 187.3912, 182.0283, 179.0285, 175.8509, 173.6871, 167.434, 
    164.1853,
  222.7256, 212.4416, 188.4799, 179.4864, 185.0863, 190.9214, 182.3547, 
    209.5815, 195.7054, 179.4009, 175.6127, 175.1866, 172.5941, 168.2175, 
    163.0484,
  224.1189, 210.8874, 188.6246, 172.3206, 180.0033, 194.3289, 188.9953, 
    202.7226, 189.148, 179.9143, 174.1509, 172.6102, 171.1512, 166.1735, 
    163.3572,
  220.4164, 209.6077, 178.6585, 176.6035, 184.4393, 190.468, 201.4509, 
    199.7828, 186.8988, 180.292, 179.2207, 173.0174, 171.7145, 166.1812, 
    163.7532,
  166.478, 168.3862, 169.8067, 175.9836, 176.5101, 174.7259, 177.251, 
    175.5779, 171.1313, 164.6014, 163.6918, 164.2197, 158.4053, 158.2165, 
    152.872,
  166.3453, 167.4509, 170.938, 175.3896, 176.7599, 175.5866, 177.1751, 
    177.6281, 170.6422, 167.9009, 166.8473, 171.292, 169.5581, 154.6752, 
    151.4978,
  167.1715, 170.1705, 172.8959, 173.2699, 175.7718, 178.1778, 174.6215, 
    176.3746, 172.8412, 169.3549, 170.9169, 171.6648, 171.1552, 168.618, 
    162.0596,
  166.9486, 167.0254, 172.278, 176.586, 176.3252, 181.4615, 173.6335, 
    172.795, 172.9247, 170.9401, 169.8536, 170.4418, 169.6595, 168.8453, 
    166.7471,
  164.2107, 166.6663, 170.2965, 173.6707, 179.1263, 178.1682, 180.2076, 
    169.8504, 164.7814, 168.3439, 170.6266, 170.6496, 169.9096, 169.636, 
    168.8548,
  172.5625, 169.7837, 176.4495, 176.6185, 179.5857, 178.1681, 175.0277, 
    188.685, 187.5836, 185.2083, 176.127, 172.5782, 170.742, 168.873, 168.3482,
  207.748, 186.4121, 182.7258, 181.3929, 178.6824, 186.4522, 186.3622, 
    186.029, 182.2762, 184.7952, 180.039, 173.2177, 171.2159, 168.6822, 
    168.0824,
  224.4503, 212.0718, 196.5245, 179.3752, 178.8491, 191.0355, 195.6415, 
    191.4267, 190.9167, 178.1439, 176.0505, 172.8553, 170.7317, 168.2554, 
    167.9697,
  215.6465, 214.8938, 195.6672, 182.2483, 180.881, 194.1808, 196.2609, 
    192.6431, 186.2635, 177.5661, 174.3692, 172.4847, 170.634, 167.2253, 
    166.7652,
  216.1772, 204.2723, 186.8994, 179.3907, 187.6693, 193.1129, 192.6436, 
    195.8208, 179.6184, 177.1568, 179.8493, 173.58, 171.067, 168.4861, 167.578,
  181.4006, 177.7977, 170.0664, 167.6595, 166.7792, 164.2089, 162.3689, 
    163.2138, 165.8722, 166.4436, 164.9159, 167.6619, 162.2676, 160.0512, 
    155.9764,
  170.7948, 170.4935, 167.2454, 164.5576, 163.0405, 165.4556, 164.4396, 
    166.7002, 166.6079, 167.8258, 165.9678, 172.1952, 172.9225, 157.0754, 
    152.9166,
  174.7279, 175.446, 173.7182, 170.4279, 167.8543, 165.6625, 163.322, 
    163.6646, 165.3363, 170.076, 169.3496, 172.6266, 174.3069, 172.233, 
    161.9637,
  192.6327, 191.8683, 183.5416, 173.6685, 169.6862, 170.2331, 165.3626, 
    163.1304, 165.8917, 169.2088, 171.884, 172.4113, 172.683, 171.1699, 
    167.9096,
  205.8485, 200.4671, 188.4624, 176.7874, 171.393, 169.3466, 175.4502, 
    168.0029, 169.8813, 169.0382, 171.7255, 172.701, 172.1432, 171.7009, 
    171.9468,
  210.0247, 206.9654, 197.1485, 186.0815, 177.5789, 177.9721, 176.2605, 
    186.9721, 182.1529, 182.0581, 178.8422, 175.013, 172.6799, 170.366, 
    169.9454,
  221.623, 213.7257, 199.0602, 186.5241, 176.5657, 180.1266, 195.7169, 
    186.3241, 183.0362, 187.5292, 182.7426, 175.054, 172.7569, 169.4143, 
    168.8446,
  220.8308, 212.7672, 190.6584, 182.2237, 170.1011, 174.2356, 194.1763, 
    191.7615, 187.6423, 180.7034, 177.8784, 174.5887, 172.0444, 168.6006, 
    167.7076,
  212.2419, 201.0372, 188.2444, 171.725, 165.0232, 174.9545, 183.4708, 
    183.6317, 182.6427, 177.2662, 174.9308, 173.2552, 170.817, 168.2425, 
    166.745,
  216.0289, 208.2375, 193.3187, 178.4707, 174.0358, 183.5513, 183.8379, 
    187.9964, 177.0219, 175.6666, 178.2328, 173.3955, 171.4536, 169.5648, 
    168.562,
  185.9361, 184.4274, 184.1617, 183.1974, 181.4623, 179.8279, 178.2845, 
    172.8754, 171.5522, 170.6972, 168.1136, 168.8416, 165.3358, 161.4097, 
    159.9989,
  178.5915, 177.119, 170.7689, 175.3925, 180.229, 181.2983, 176.4449, 
    177.0169, 171.9814, 169.0875, 167.8306, 167.1469, 168.3191, 162.4476, 
    160.4049,
  190.8187, 184.378, 175.3083, 167.825, 167.8108, 174.5708, 172.5, 171.5925, 
    174.3074, 170.0639, 171.661, 168.9249, 165.5687, 165.9458, 164.2476,
  214.3379, 203.3923, 194.4197, 182.1098, 173.034, 175.7978, 170.189, 
    171.045, 171.0753, 172.3801, 171.6471, 169.6376, 168.7343, 165.7007, 
    165.1032,
  219.1346, 214.8444, 204.4563, 198.2721, 181.3595, 175.2894, 179.45, 
    175.1653, 179.8508, 169.7688, 169.8957, 169.153, 168.1687, 167.8366, 
    168.1967,
  223.2824, 216.0713, 204.5733, 195.9732, 180.5418, 174.6087, 179.8774, 
    181.3522, 178.1612, 175.8398, 172.8416, 171.8243, 169.5244, 168.642, 
    168.7205,
  224.9825, 215.9173, 207.1808, 194.4066, 179.79, 183.7701, 189.974, 
    178.6213, 182.139, 183.0663, 175.862, 171.0129, 169.1711, 167.1716, 
    168.9124,
  222.8335, 216.1134, 212.9346, 202.4344, 183.7906, 192.569, 183.3448, 
    183.0964, 181.9746, 178.2222, 175.2475, 172.023, 170.3252, 168.074, 
    168.5882,
  220.1729, 217.8751, 212.8803, 198.5538, 190.181, 189.497, 183.0446, 
    184.8053, 182.4112, 177.9495, 174.1245, 173.2157, 171.0472, 168.8431, 
    168.3259,
  222.1404, 215.1173, 210.426, 199.0352, 186.9793, 184.6302, 180.9359, 
    188.6669, 179.8921, 176.6857, 178.0779, 173.7811, 172.5935, 170.4701, 
    169.2114,
  201.137, 200.598, 197.7709, 195.1946, 191.07, 189.1099, 188.3615, 188.4368, 
    186.9038, 177.2177, 176.1898, 175.7781, 175.2661, 173.0575, 170.8612,
  204.6354, 203.6681, 201.2054, 196.7982, 189.3214, 186.8484, 186.854, 
    187.7634, 185.8832, 184.6823, 180.1917, 180.1934, 180.8129, 173.4452, 
    171.8294,
  218.9124, 215.113, 208.6862, 200.3769, 194.062, 183.5244, 178.0446, 
    177.9584, 180.8443, 182.474, 182.6483, 182.6546, 179.4995, 177.375, 
    174.9554,
  220.3008, 221.6018, 219.3554, 208.8725, 199.479, 190.2938, 177.1996, 
    171.5239, 172.6688, 177.7074, 178.5134, 178.5735, 179.6869, 177.7137, 
    175.9337,
  222.6054, 221.6855, 213.3962, 218.2912, 203.3975, 186.7951, 183.3094, 
    175.2561, 170.4503, 164.0727, 169.0855, 174.4894, 175.4616, 176.326, 
    175.9172,
  223.0204, 220.0336, 214.4631, 215.946, 204.9157, 185.8612, 177.6879, 
    171.9068, 163.6384, 161.201, 166.2855, 173.0065, 172.8644, 171.9967, 
    171.5938,
  221.4343, 221.9093, 216.0124, 207.9754, 202.5792, 200.5546, 189.9064, 
    178.9131, 170.5401, 169.2531, 169.168, 169.4072, 170.0011, 168.9229, 
    171.1932,
  223.5081, 223.2796, 218.5562, 212.4082, 211.1415, 205.6401, 191.8141, 
    190.2662, 189.0375, 177.2652, 168.8704, 168.4955, 167.5969, 167.3934, 
    171.2308,
  222.9599, 217.2496, 216.5479, 217.7561, 212.9341, 199.1613, 192.4662, 
    186.1935, 184.1102, 176.6313, 168.2029, 166.5806, 164.4353, 166.7077, 
    168.2617,
  218.0827, 219.0242, 216.8354, 210.4279, 211.8744, 190.5135, 184.6609, 
    185.3878, 180.9941, 175.7982, 172.5324, 165.5814, 163.4525, 165.2198, 
    167.3323,
  198.939, 200.4755, 201.2559, 195.9594, 194.5145, 191.8964, 191.0119, 
    183.6259, 181.5524, 176.84, 169.8398, 164.7493, 164.1519, 166.0679, 
    167.644,
  204.4088, 204.2846, 204.301, 200.1799, 195.0274, 195.1188, 188.2293, 
    188.5228, 186.6232, 184.6713, 181.0763, 178.8566, 171.4597, 166.9815, 
    167.7378,
  205.2804, 217.3899, 212.8153, 202.8078, 199.3296, 190.6413, 188.9784, 
    185.2427, 186.6859, 184.898, 182.7755, 184.8805, 178.4239, 172.678, 
    171.6138,
  214.7155, 220.7104, 215.3476, 213.5023, 204.3632, 200.0417, 190.6676, 
    191.5457, 189.2368, 188.8189, 186.197, 186.0777, 183.5424, 180.1349, 
    175.5511,
  216.7589, 221.4525, 216.5313, 217.0653, 209.6936, 210.4752, 201.8719, 
    187.39, 186.8803, 180.205, 178.9237, 179.7358, 181.5675, 180.2549, 
    177.7995,
  208.8435, 222.1394, 213.649, 208.644, 206.8466, 204.8896, 194.3791, 
    196.5057, 193.6647, 188.3182, 178.4833, 173.4153, 174.6557, 175.7855, 
    173.4257,
  213.9571, 225.0484, 212.1274, 201.9658, 200.428, 188.2744, 191.5245, 
    193.9815, 196.364, 192.4842, 179.888, 170.6204, 172.0434, 168.6493, 
    171.9727,
  222.0314, 224.4347, 209.8405, 194.7057, 193.8001, 198.0221, 190.1376, 
    192.0837, 193.2535, 189.7954, 180.3781, 168.6829, 168.1433, 167.8034, 
    166.4569,
  225.8037, 212.5829, 189.6076, 185.7094, 187.9337, 182.7154, 188.747, 
    189.5729, 189.61, 185.6216, 177.9126, 168.9242, 165.1539, 163.5357, 
    166.6832,
  210.1907, 196.6497, 175.9524, 174.5143, 183.2454, 182.1584, 188.9381, 
    186.3952, 183.6035, 178.3698, 177.8573, 166.5419, 161.9963, 161.2855, 
    172.1433,
  201.3077, 206.9236, 199.1504, 200.8688, 197.2352, 194.3553, 187.0318, 
    181.707, 179.6975, 180.8202, 182.3737, 183.5744, 181.1294, 176.8055, 
    174.016,
  208.7455, 204.8034, 200.7045, 200.3814, 195.2201, 189.8144, 182.3432, 
    176.4996, 179.0598, 180.827, 183.721, 186.6646, 185.8595, 177.636, 
    172.6492,
  210.9603, 211.2, 210.6733, 199.338, 188.4558, 175.935, 179.6363, 169.0557, 
    173.8833, 181.5927, 186.0819, 188.7775, 187.0974, 180.554, 172.6246,
  210.323, 215.5924, 199.9531, 193.6235, 169.2417, 164.6452, 162.9282, 
    173.6653, 176.143, 179.3794, 186.2676, 188.9195, 187.9163, 183.1179, 
    175.159,
  221.3375, 214.7017, 196.2718, 169.9489, 154.6029, 157.1804, 165.5013, 
    169.4212, 177.8594, 181.4758, 188.1699, 189.3836, 187.4433, 183.9132, 
    180.7028,
  206.2656, 203.5202, 177.3271, 154.6332, 153.0301, 165.1969, 169.5224, 
    178.4566, 187.6683, 190.3321, 189.6664, 188.4615, 186.3886, 184.8781, 
    181.8454,
  202.1028, 188.7193, 156.3155, 153.0055, 155.6083, 173.3039, 181.2402, 
    185.8304, 186.4222, 189.0144, 189.7861, 185.5667, 183.3308, 180.1756, 
    179.682,
  196.9222, 164.4534, 149.7614, 148.3932, 159.7646, 181.1273, 190.8602, 
    193.8705, 188.3065, 184.2405, 184.2908, 182.5663, 181.8146, 176.757, 
    177.1372,
  186.9677, 156.4128, 143.8653, 151.5721, 162.6754, 185.3759, 196.259, 
    195.6034, 184.2768, 183.8835, 182.7102, 181.8069, 179.593, 173.3635, 
    173.6883,
  170.5959, 155.8853, 148.7005, 157.2275, 177.7543, 191.084, 193.8798, 
    194.0478, 184.4082, 180.5956, 179.7107, 182.0059, 176.9849, 172.695, 
    170.8642,
  202.229, 207.7352, 199.7722, 200.0305, 178.258, 167.9727, 171.8902, 
    174.5194, 174.3485, 173.67, 176.3847, 176.4626, 177.6967, 180.3743, 
    180.0861,
  209.692, 205.4255, 202.285, 183.504, 165.4036, 168.7363, 171.9462, 
    175.9943, 181.0437, 184.0869, 181.6712, 178.2309, 179.7339, 178.4809, 
    180.3243,
  212.6818, 206.4642, 199.6864, 170.7939, 161.1975, 167.659, 183.7512, 
    184.3246, 184.2103, 187.7095, 182.1074, 175.687, 176.2946, 179.8106, 
    183.955,
  205.1552, 204.4346, 177.9214, 166.353, 164.4437, 179.5303, 186.5881, 
    196.0936, 193.6555, 185.3309, 178.5414, 179.5888, 184.3356, 186.7566, 
    187.5929,
  207.7267, 199.3423, 172.8016, 168.349, 171.3702, 188.1026, 199.9558, 
    191.7853, 185.5161, 187.1343, 184.366, 186.8019, 188.8631, 188.718, 
    185.7857,
  205.7931, 193.2303, 176.9594, 169.4131, 169.4384, 185.6118, 196.4596, 
    189.5744, 193.5157, 192.2303, 186.6828, 187.6247, 187.5094, 185.9406, 
    186.8201,
  202.2805, 192.4953, 182.9661, 174.6081, 170.0408, 174.9957, 185.5143, 
    187.1301, 188.3983, 190.6951, 186.8669, 186.0805, 187.4975, 185.5372, 
    181.8047,
  203.4386, 194.6193, 185.8916, 180.3146, 168.8974, 165.273, 174.3004, 
    181.9896, 181.029, 183.6129, 182.7975, 184.0866, 182.307, 180.696, 
    179.4954,
  204.3684, 197.5087, 189.776, 178.8448, 165.6551, 166.0237, 165.437, 
    172.1369, 174.8944, 176.4722, 177.8181, 179.2517, 179.6257, 178.1369, 
    177.9933,
  202.291, 196.5675, 190.6381, 188.9395, 172.8465, 166.3956, 164.3654, 
    165.6178, 167.8132, 170.2978, 172.5614, 177.3634, 178.7883, 177.8752, 
    177.5699,
  204.3727, 205.5432, 199.3987, 198.9084, 193.8961, 192.6417, 192.5794, 
    183.1397, 177.3069, 181.0682, 187.8699, 188.6855, 184.3013, 183.8764, 
    180.2226,
  207.5947, 204.7762, 200.3936, 197.3153, 190.2737, 193.1381, 194.1724, 
    181.4731, 173.5026, 181.1958, 185.42, 192.2168, 189.6246, 180.7171, 
    178.1054,
  215.2231, 216.1561, 208.3902, 197.3712, 190.7881, 186.937, 187.9907, 
    169.6847, 167.3338, 171.829, 183.2462, 191.8826, 192.0362, 188.0683, 
    181.5404,
  211.6674, 201.018, 200.0387, 199.7684, 194.7812, 192.5815, 185.5556, 
    175.3914, 172.2125, 168.5348, 175.9574, 188.866, 192.1782, 188.6927, 
    185.2937,
  204.2196, 201.9737, 198.8891, 196.0486, 194.2234, 194.4142, 194.1829, 
    188.4, 172.6079, 166.0823, 167.6786, 183.4937, 187.7873, 189.3134, 188.219,
  214.3451, 218.6251, 203.0727, 197.956, 199.788, 197.7984, 185.9522, 
    177.9344, 168.7334, 165.0383, 165.6364, 176.9911, 183.9811, 185.7419, 
    185.0041,
  219.4479, 205.6696, 208.705, 215.0612, 201.0552, 197.6209, 187.2055, 
    175.0476, 170.7408, 170.0706, 169.5007, 172.2345, 180.5729, 181.9111, 
    180.3616,
  210.5738, 217.401, 212.567, 216.581, 200.4428, 197.1111, 186.4124, 180.507, 
    181.767, 177.2554, 170.9701, 172.705, 177.4881, 181.7496, 177.5605,
  209.698, 209.2333, 202.8481, 214.1317, 196.703, 194.0285, 190.3497, 
    186.2864, 182.9395, 181.927, 178.0585, 176.2387, 177.434, 175.8529, 
    176.841,
  202.8332, 202.9368, 205.486, 208.5965, 204.7287, 201.9749, 193.7406, 
    193.1904, 192.0376, 189.1043, 185.0792, 178.5037, 176.8747, 179.0568, 
    177.8408,
  175.2228, 187.9012, 199.4427, 202.8709, 201.0859, 201.243, 201.117, 
    198.5177, 193.4387, 180.7805, 184.1809, 188.3084, 184.9035, 178.4158, 
    176.7191,
  180.8177, 195.5332, 201.7409, 202.7208, 200.9991, 201.2199, 201.0866, 
    203.3819, 197.7207, 190.9062, 181.575, 188.6385, 187.1126, 176.2471, 
    174.2617,
  199.4154, 199.6942, 201.122, 201.374, 203.6178, 200.2581, 203.4118, 
    197.6539, 193.4328, 192.4292, 189.5847, 187.593, 188.1203, 187.4241, 
    185.0393,
  202.9856, 201.5832, 202.8405, 203.3266, 203.4547, 203.193, 199.2478, 
    206.0317, 199.7365, 193.7758, 190.7253, 187.7478, 183.7887, 185.9355, 
    186.8797,
  202.9508, 202.4919, 202.9273, 203.0552, 203.1005, 201.3, 199.0299, 
    194.7399, 192.5831, 193.4093, 191.316, 190.5727, 186.5332, 184.0633, 
    188.6682,
  203.0346, 204.4895, 203.5004, 202.9516, 201.9325, 199.3391, 191.577, 
    190.2457, 192.2038, 192.986, 193.0688, 193.6853, 189.0792, 185.6307, 
    183.9385,
  200.5421, 209.4431, 202.6678, 204.719, 199.9878, 194.8788, 189.0722, 
    186.5546, 189.4042, 190.1202, 194.4409, 195.579, 193.1849, 187.5262, 
    184.7669,
  209.5017, 214.1681, 210.0848, 202.4665, 193.6355, 190.9653, 187.7468, 
    187.3191, 190.6036, 192.3267, 193.9281, 196.555, 195.3041, 192.0236, 
    186.1132,
  212.9641, 212.6061, 210.7861, 200.2177, 196.9084, 190.7924, 190.5083, 
    186.0294, 193.236, 194.9742, 195.0412, 199.3432, 196.3987, 193.3738, 
    189.6475,
  211.8967, 209.1337, 207.1206, 190.0883, 186.3555, 188.077, 187.0372, 
    193.7527, 192.7626, 195.1213, 196.451, 195.7617, 195.502, 194.8823, 
    191.3828,
  180.5681, 197.4022, 202.8646, 205.2315, 200.6681, 198.2383, 196.1381, 
    190.4534, 186.1688, 187.789, 181.6593, 185.4892, 175.3155, 178.5193, 
    179.6768,
  193.4261, 200.9077, 204.8512, 206.325, 201.7239, 198.7204, 195.6855, 
    189.1102, 182.2368, 185.87, 183.6016, 184.5618, 185.2551, 183.1731, 
    181.3422,
  199.9434, 204.8558, 207.0419, 204.7372, 202.0381, 198.4895, 199.144, 
    183.1518, 178.6062, 179.9622, 185.0804, 180.9255, 184.7184, 184.611, 
    179.2007,
  205.6835, 208.2839, 206.2828, 205.3035, 203.5209, 201.899, 195.7424, 
    184.8091, 182.9083, 179.9218, 180.7608, 178.5344, 178.1389, 175.5392, 
    177.0741,
  209.7725, 210.6791, 208.097, 207.0191, 204.3085, 200.0119, 192.8599, 
    188.0676, 186.7369, 179.4064, 178.2937, 175.7941, 174.5933, 173.1417, 
    174.3118,
  212.9328, 213.0701, 213.1094, 209.8327, 208.7395, 197.0592, 184.8454, 
    181.6285, 176.9969, 169.0521, 170.1604, 174.007, 171.2271, 171.1843, 
    171.2754,
  216.3716, 212.2275, 211.2487, 211.6117, 210.0223, 191.7839, 175.2406, 
    168.5055, 167.9942, 167.3295, 167.7045, 170.8378, 168.7739, 167.1587, 
    166.608,
  217.3408, 212.1824, 211.6674, 211.7829, 195.1115, 186.458, 172.9527, 
    166.6086, 162.4677, 159.8269, 163.2548, 162.4606, 164.9411, 161.734, 
    166.3529,
  215.849, 211.6161, 204.9158, 196.1373, 193.8128, 182.7525, 170.9818, 
    161.9824, 160.8105, 155.2305, 159.7045, 156.8757, 158.2725, 161.5821, 
    163.2784,
  204.4634, 193.6946, 187.5359, 185.9227, 185.8037, 182.2688, 173.2864, 
    164.7658, 160.7758, 157.7911, 155.5839, 157.878, 154.6056, 155.4387, 
    160.9957,
  195.1595, 208.9485, 206.2002, 201.516, 194.9736, 194.6325, 197.1393, 
    189.4294, 184.9838, 178.838, 177.5581, 173.2391, 172.0721, 177.2769, 
    169.7825,
  199.7376, 206.7042, 208.0409, 202.2363, 195.9175, 196.1006, 195.9254, 
    195.8199, 193.74, 183.4486, 176.0206, 171.5843, 173.3012, 175.5407, 
    176.5692,
  206.2942, 209.5781, 211.9361, 206.3188, 200.4786, 191.2077, 202.2846, 
    192.4264, 185.4487, 190.4058, 187.384, 176.2435, 174.6687, 175.4193, 
    177.5896,
  215.2034, 216.5201, 219.4892, 216.9355, 210.6898, 203.2328, 199.0992, 
    189.8642, 175.9258, 170.9038, 182.4126, 180.3271, 176.3693, 174.1982, 
    177.2271,
  214.9829, 218.7109, 220.7153, 220.0223, 214.8723, 209.5607, 195.8073, 
    190.9946, 183.7964, 174.774, 173.7272, 178.9706, 181.161, 185.8334, 
    178.9015,
  214.9785, 216.341, 218.3452, 220.1233, 218.6875, 209.5947, 199.0288, 
    193.7593, 183.7805, 180.7762, 186.8007, 190.6015, 186.4295, 189.9576, 
    188.6447,
  214.162, 213.5255, 216.9039, 217.4697, 217.4894, 204.8481, 199.3594, 
    188.9763, 187.5625, 195.3712, 196.5189, 196.7485, 199.5254, 194.7963, 
    192.7882,
  215.8695, 215.2139, 218.06, 219.3787, 210.5606, 203.5757, 199.2202, 
    193.6647, 202.8627, 203.8951, 201.635, 204.1803, 202.0417, 198.9839, 
    194.488,
  218.153, 218.1477, 212.7593, 205.4177, 196.3853, 200.1575, 197.9361, 
    203.5179, 205.2466, 209.4538, 209.926, 208.4253, 200.5834, 196.0922, 
    193.2495,
  215.2352, 209.2097, 202.705, 189.4467, 190.3101, 197.1825, 204.411, 
    206.7478, 210.7153, 208.396, 211.2988, 206.5797, 199.3755, 196.8396, 
    191.1571,
  199.3675, 201.1226, 205.6254, 205.941, 203.6208, 201.4194, 203.0839, 
    196.8361, 193.4968, 189.1066, 189.6252, 191.409, 189.5607, 189.2242, 
    186.7863,
  198.1215, 197.5201, 204.0715, 204.9231, 202.3248, 200.7848, 203.187, 
    198.8969, 197.0233, 193.7061, 193.1524, 194.2577, 194.6769, 196.7068, 
    192.155,
  191.4934, 193.6052, 197.0729, 198.1019, 203.1504, 200.6148, 205.0927, 
    201.3496, 202.6083, 200.5159, 199.7475, 193.6334, 194.6892, 198.05, 
    193.0619,
  191.9844, 189.1718, 190.9985, 191.6094, 193.0647, 196.3823, 197.3743, 
    195.7983, 200.6351, 198.7643, 198.9138, 195.3037, 194.6776, 195.8422, 
    194.123,
  187.0397, 185.6533, 187.6708, 180.1113, 185.5917, 186.6537, 185.9754, 
    192.9188, 196.7262, 192.7933, 195.9791, 192.6514, 191.6884, 191.1816, 
    188.3362,
  193.832, 189.9705, 186.9846, 184.2106, 182.2473, 180.6964, 184.7343, 
    184.9767, 191.1676, 191.1402, 190.5094, 188.8005, 190.4292, 186.9472, 
    184.0062,
  197.6391, 193.0078, 189.6459, 185.701, 182.0988, 187.7043, 185.1615, 
    187.702, 185.4539, 188.537, 184.0391, 184.6243, 188.2104, 186.1781, 
    182.6918,
  200.5696, 193.4866, 195.1906, 192.8872, 193.7604, 195.3397, 201.3712, 
    206.2444, 201.4651, 191.3162, 187.7361, 187.9473, 186.8998, 185.3306, 
    184.7978,
  202.1246, 199.4647, 200.6838, 201.0996, 210.3558, 210.8041, 212.4534, 
    204.6093, 196.4145, 191.2971, 190.7847, 189.1697, 187.8546, 183.2923, 
    178.8963,
  207.0369, 214.2264, 212.1416, 216.2019, 215.1626, 207.341, 197.7375, 
    194.6712, 189.4048, 188.9298, 187.5429, 186.7601, 184.3527, 177.8828, 
    176.936,
  186.362, 199.4793, 204.4702, 201.5064, 200.9714, 198.0721, 197.2128, 
    191.3372, 186.1103, 180.7702, 177.5011, 177.1512, 177.032, 174.6706, 
    177.3747,
  198.9951, 208.3084, 204.928, 201.9433, 198.3788, 195.7711, 193.3657, 
    189.4035, 190.3139, 180.7467, 173.2765, 173.6443, 172.2686, 171.9184, 
    173.7342,
  208.3218, 207.1472, 205.8305, 200.477, 194.9472, 191.8591, 189.5906, 
    182.7503, 182.7979, 174.8036, 169.4035, 167.3845, 170.3148, 175.5756, 
    178.6121,
  211.4587, 208.8453, 201.3408, 196.66, 192.9271, 192.1318, 187.2817, 
    185.3737, 176.5682, 169.3788, 165.625, 167.7254, 171.9588, 176.3671, 
    177.5774,
  212.6144, 206.0544, 201.8606, 200.7211, 196.0599, 189.3698, 186.0064, 
    184.7909, 179.0144, 166.0368, 168.0686, 174.5596, 178.9288, 181.0039, 
    181.012,
  210.4932, 211.0325, 206.5338, 202.2629, 198.7729, 194.9131, 189.5288, 
    181.8054, 181.213, 179.1825, 175.6949, 181.6176, 179.8876, 182.4542, 
    183.66,
  212.5768, 213.3143, 210.4922, 204.1836, 202.3413, 191.6201, 194.6022, 
    185.5224, 185.6086, 179.5456, 180.3904, 181.6888, 182.6557, 183.3702, 
    187.0869,
  210.0654, 210.2057, 208.9992, 207.6762, 204.8127, 198.8187, 199.2979, 
    197.7268, 185.0305, 183.9921, 182.5292, 184.6395, 182.7209, 183.4508, 
    185.7516,
  217.0168, 210.9196, 211.1508, 206.816, 203.9684, 204.7011, 207.6609, 
    188.7431, 188.9583, 185.7445, 188.0872, 181.944, 181.5333, 180.5652, 
    181.7822,
  219.5653, 213.1706, 206.275, 203.5226, 206.5217, 203.1616, 192.1717, 
    190.0592, 186.2073, 184.2043, 182.0421, 181.5229, 178.2556, 177.5312, 
    178.4748,
  188.1551, 199.5356, 210.9589, 212.2143, 205.8541, 197.4967, 196.0619, 
    194.8857, 197.1316, 192.7615, 193.874, 186.9998, 184.1326, 181.1009, 
    177.6371,
  193.5579, 203.9705, 213.9953, 210.2984, 204.2813, 199.4047, 193.8535, 
    195.0812, 200.8097, 199.6451, 196.5206, 190.0514, 184.8982, 181.1631, 
    180.0778,
  209.0441, 216.5441, 217.0527, 207.4774, 203.1293, 199.1783, 204.5163, 
    195.4631, 197.0341, 198.7757, 196.5691, 194.3801, 187.6492, 185.0584, 
    180.9437,
  218.3556, 220.5432, 218.5039, 206.1816, 199.313, 202.1966, 201.5242, 
    207.4261, 201.4429, 195.5987, 195.0572, 193.8889, 190.0438, 185.2631, 
    186.2272,
  222.7526, 218.9823, 216.5507, 208.0488, 205.0717, 201.4885, 198.3603, 
    200.2304, 198.5838, 197.257, 195.4655, 193.645, 190.8728, 188.6018, 
    182.8673,
  222.1099, 220.2137, 216.4978, 210.8326, 210.036, 202.8661, 194.303, 
    196.872, 196.9413, 196.795, 195.4931, 189.0912, 189.0091, 188.0452, 
    183.6048,
  220.0483, 218.3685, 216.6132, 214.2702, 213.0801, 203.7045, 196.4167, 
    193.0627, 191.0088, 190.3575, 189.8581, 187.7747, 190.4066, 186.8241, 
    187.4658,
  225.8829, 220.6426, 216.2462, 214.022, 210.948, 200.2318, 194.0554, 
    193.0922, 187.0437, 183.5318, 181.9597, 185.6269, 184.9256, 186.3759, 
    184.0785,
  226.9079, 221.7666, 218.354, 212.527, 203.7512, 195.1725, 191.9288, 
    187.9048, 184.0441, 180.1928, 181.0595, 184.6977, 185.4875, 180.4512, 
    179.3387,
  226.2915, 222.0146, 211.9372, 199.5522, 189.097, 187.0114, 188.011, 
    178.7499, 176.3721, 177.513, 179.159, 180.4532, 180.5079, 178.5222, 
    179.251,
  185.9149, 188.3181, 199.3785, 210.5087, 210.395, 212.3794, 212.0359, 
    208.886, 199.2099, 198.5671, 198.2734, 196.7849, 194.15, 181.9129, 
    175.3031,
  187.7746, 192.6179, 204.3523, 206.7214, 213.4958, 217.6848, 215.1716, 
    209.6732, 209.3009, 199.589, 194.2669, 191.1259, 185.0802, 180.769, 
    176.0489,
  202.8151, 204.829, 211.2661, 213.43, 216.2475, 215.2336, 214.1919, 
    193.4666, 184.5062, 188.7486, 186.9967, 188.7548, 180.3971, 172.3213, 
    171.8293,
  207.7875, 215.682, 218.4554, 220.1885, 218.5678, 218.0806, 208.1086, 
    197.1832, 185.8992, 178.8485, 188.45, 184.189, 175.3887, 178.9883, 
    176.5416,
  216.1966, 218.3795, 220.6631, 221.7017, 220.093, 217.6751, 213.8169, 
    201.3846, 196.9154, 192.8242, 184.3258, 187.4557, 180.0593, 177.9717, 
    173.393,
  217.8552, 222.2033, 221.0446, 223.0901, 220.0845, 219.04, 213.0298, 
    203.3393, 201.4414, 191.5633, 188.7326, 190.3646, 184.772, 178.2007, 
    175.171,
  220.6161, 220.7248, 221.0257, 219.7534, 220.9865, 215.8641, 211.5527, 
    202.1963, 195.4531, 195.9601, 188.3924, 189.3708, 184.065, 175.176, 
    171.4156,
  220.2152, 220.8093, 220.712, 220.1187, 219.5198, 214.3557, 213.1702, 
    206.5105, 203.2709, 198.9028, 193.9539, 189.1464, 177.3031, 171.926, 
    171.4735,
  221.4151, 220.1815, 221.0228, 221.0107, 217.2341, 214.086, 214.6173, 
    209.7948, 203.3855, 196.9648, 195.5969, 184.2618, 174.4667, 174.3918, 
    164.8985,
  219.0371, 218.5253, 218.734, 216.261, 209.3667, 207.6123, 212.1129, 
    208.5496, 201.3807, 196.8587, 191.5772, 177.5129, 173.7161, 168.7015, 
    168.2911,
  185.263, 189.3972, 184.8334, 188.2115, 189.9402, 193.9083, 199.182, 
    204.6864, 204.3806, 203.1179, 202.3388, 204.4013, 204.1433, 203.9069, 
    198.6311,
  188.7037, 193.7925, 190.3229, 192.3455, 192.8994, 199.8355, 194.5164, 
    203.6855, 209.5079, 205.6751, 201.8598, 205.1437, 203.918, 203.0058, 
    200.1215,
  197.0851, 203.4668, 201.6777, 199.301, 198.8813, 200.8195, 204.9384, 
    196.4906, 203.0505, 207.86, 206.6772, 202.1154, 201.8179, 200.7634, 
    201.6575,
  201.8477, 208.0236, 203.3499, 207.2957, 201.8767, 201.1818, 199.702, 
    202.9147, 203.475, 204.6156, 204.9855, 200.9662, 202.9842, 197.1034, 
    198.6453,
  203.0317, 201.4774, 202.471, 201.8698, 201.1205, 198.2115, 193.5309, 
    200.2123, 202.5489, 207.5608, 201.3658, 199.985, 199.9132, 197.8718, 
    195.7849,
  201.6191, 199.2109, 199.2513, 199.6915, 197.9969, 195.262, 195.3896, 
    194.2996, 197.7719, 197.5937, 198.877, 199.3745, 198.8498, 197.9802, 
    193.4639,
  203.9602, 201.154, 200.3845, 202.477, 200.2919, 196.2676, 197.3933, 
    191.9687, 192.8766, 194.7937, 198.4357, 199.1927, 197.0148, 195.1748, 
    188.6887,
  206.2727, 201.5273, 205.0945, 198.8967, 198.1327, 192.8392, 192.4631, 
    191.7218, 192.3332, 193.7006, 196.0991, 200.4682, 195.2203, 190.6307, 
    184.0941,
  199.5171, 197.4179, 193.1552, 195.7651, 194.9076, 192.8708, 196.2324, 
    193.4482, 192.9446, 192.7763, 194.7507, 198.1013, 192.28, 187.8305, 
    174.7474,
  185.0881, 179.587, 183.4568, 184.689, 188.4131, 185.7643, 190.2995, 
    195.9391, 191.3693, 194.7953, 195.9634, 192.6451, 185.1119, 180.6057, 
    169.7119,
  189.1532, 199.0325, 189.6304, 182.3546, 175.6521, 174.9652, 174.4733, 
    173.4325, 176.7643, 181.2953, 179.9637, 183.8737, 184.9358, 189.0773, 
    186.827,
  173.6711, 182.6187, 178.3466, 171.832, 173.5172, 175.9695, 171.443, 
    172.7857, 179.2971, 181.3095, 179.9008, 180.8605, 182.4645, 190.0738, 
    185.1553,
  166.3784, 176.1279, 177.085, 171.5612, 165.6576, 172.118, 177.8602, 
    166.6158, 173.0886, 180.61, 186.5015, 180.1453, 181.6271, 185.3178, 
    187.3187,
  167.0392, 166.5454, 171.8719, 167.8862, 176.3772, 174.3398, 181.7343, 
    176.1407, 174.8461, 174.6083, 182.3814, 189.4779, 187.0962, 188.6461, 
    188.9084,
  170.1871, 166.1966, 167.8872, 167.9942, 169.7317, 170.228, 174.3819, 
    184.9376, 189.3236, 181.7934, 185.459, 191.9905, 195.149, 192.3968, 
    189.9054,
  166.9809, 168.3841, 171.9784, 176.9073, 181.7313, 183.3409, 181.9389, 
    193.6015, 192.7685, 186.6442, 191.0166, 197.0186, 191.8262, 194.0912, 
    189.1374,
  190.8308, 187.5918, 191.8385, 192.3919, 197.8343, 194.8331, 199.9394, 
    198.0772, 199.3761, 195.2043, 196.6242, 194.7293, 192.2725, 190.9979, 
    189.8168,
  200.7285, 196.9603, 196.7591, 200.2925, 200.6962, 199.346, 202.9022, 
    203.5256, 202.2992, 195.9187, 192.9168, 193.0513, 193.6865, 191.9198, 
    185.6594,
  191.2745, 191.0385, 189.2875, 183.1393, 182.3921, 186.3139, 190.5548, 
    191.2983, 190.2853, 183.6925, 187.2854, 183.0737, 182.78, 179.1937, 
    179.6217,
  198.6954, 198.9019, 193.6618, 188.0897, 180.5537, 177.6429, 174.0471, 
    173.7123, 175.9299, 175.1497, 171.751, 169.5542, 169.9831, 172.7162, 
    172.1098,
  191.3736, 195.0507, 190.6013, 191.5699, 189.7399, 191.0518, 195.992, 
    194.9349, 190.6955, 191.4325, 191.2973, 188.5169, 185.9338, 180.9052, 
    179.009,
  196.9728, 197.9207, 196.3939, 192.9644, 188.0449, 193.9179, 198.1392, 
    192.3967, 191.8536, 188.9495, 192.8283, 189.5754, 184.6782, 178.8152, 
    181.68,
  182.9255, 198.5889, 198.7511, 197.8758, 191.3747, 190.2848, 205.0328, 
    193.5398, 192.8436, 190.0915, 191.6345, 190.1419, 189.0019, 184.0932, 
    186.4572,
  173.399, 174.3815, 182.5743, 189.3062, 196.3173, 192.4206, 188.4939, 
    206.3878, 199.546, 191.3821, 193.0001, 196.9856, 190.8637, 189.7408, 
    193.3532,
  173.2329, 173.0533, 173.6056, 181.0025, 185.6984, 196.5918, 191.2878, 
    194.3407, 199.8802, 199.5283, 196.4122, 194.704, 192.8439, 195.7807, 
    196.1954,
  206.8889, 200.122, 188.4038, 178.3052, 177.2521, 174.9745, 179.2434, 
    198.0718, 202.068, 191.0545, 196.9013, 197.8477, 196.156, 197.1338, 
    196.1947,
  216.6859, 217.5269, 210.1161, 207.4043, 206.6415, 205.144, 198.3163, 
    200.0006, 202.5024, 195.9793, 192.6263, 195.3279, 197.7153, 197.6788, 
    198.3524,
  209.526, 214.8769, 216.0057, 214.6892, 218.6358, 211.9373, 211.9629, 
    209.0345, 204.6608, 195.5496, 190.0709, 191.355, 190.2866, 188.0936, 
    186.0567,
  211.443, 213.815, 211.9946, 208.5591, 216.6936, 217.5327, 213.9811, 
    205.8303, 200.2417, 195.4962, 195.7987, 192.3038, 191.249, 188.5243, 
    182.4504,
  206.595, 213.6675, 211.847, 211.6419, 213.2375, 212.6455, 205.7096, 
    196.1222, 194.8399, 191.7971, 189.1377, 183.5325, 185.7356, 182.438, 
    178.5729,
  180.0439, 180.5445, 180.3074, 184.7195, 180.0104, 184.2719, 189.6471, 
    187.8432, 190.8158, 191.9866, 192.2198, 192.7216, 191.7106, 190.9876, 
    188.7547,
  193.471, 192.1008, 187.5037, 185.5649, 184.567, 191.2122, 189.9866, 
    188.0821, 191.8379, 191.7738, 192.8606, 192.9734, 193.377, 189.303, 
    187.3243,
  204.4913, 200.3465, 194.2158, 190.5903, 188.3594, 187.2592, 192.3814, 
    188.1735, 189.788, 190.2133, 190.3686, 192.1752, 188.1215, 188.2339, 
    186.2939,
  206.8165, 204.6275, 199.0605, 193.2615, 187.0893, 188.9789, 186.418, 
    193.1604, 194.4234, 189.9918, 187.6513, 189.5129, 186.4167, 187.2093, 
    183.9772,
  202.8523, 206.4774, 204.1592, 197.497, 194.8391, 184.1793, 186.8071, 
    189.9691, 194.8651, 184.6659, 184.889, 188.1406, 183.5092, 184.2552, 
    185.4344,
  202.5473, 208.3004, 214.7621, 212.1723, 203.5574, 193.148, 182.4755, 
    187.5728, 190.7053, 183.8016, 184.6027, 184.4091, 182.5167, 184.4076, 
    184.1376,
  205.4354, 211.0607, 210.4166, 213.0109, 214.5069, 212.521, 206.6057, 
    195.5356, 196.715, 197.3407, 194.2361, 189.9701, 189.4438, 187.1324, 
    188.9443,
  205.7802, 199.2917, 204.6766, 211.1331, 208.801, 210.6762, 207.0723, 
    206.191, 205.3701, 196.9095, 197.3457, 196.3582, 197.7568, 199.5831, 
    198.7907,
  204.8037, 206.6963, 203.3938, 192.8141, 200.2944, 193.9765, 200.2788, 
    193.8431, 192.0547, 192.0992, 199.5014, 195.6145, 195.9186, 196.0623, 
    198.797,
  195.4574, 194.3308, 185.8765, 195.4966, 193.4245, 192.6344, 192.9656, 
    188.5645, 189.9329, 184.2695, 191.2838, 188.42, 189.3435, 189.9725, 
    192.8107,
  194.3575, 194.9478, 190.4254, 189.1392, 182.0735, 181.0458, 179.088, 
    170.1591, 168.9705, 166.0673, 164.2255, 167.4073, 167.7351, 174.0048, 
    174.2676,
  202.3378, 197.1005, 193.7604, 188.5478, 182.9544, 185.2925, 180.5147, 
    178.3773, 175.4833, 172.6473, 165.6229, 168.7782, 170.4633, 171.395, 
    170.4494,
  190.0944, 192.9684, 188.4733, 190.3919, 187.8796, 188.4827, 187.0135, 
    172.5683, 176.9828, 176.397, 175.2886, 172.3458, 172.8163, 173.1509, 
    172.4482,
  182.6933, 183.515, 187.7257, 186.1363, 183.6788, 185.5775, 183.3129, 
    180.6714, 181.6911, 180.947, 183.2011, 181.0525, 176.9923, 175.2939, 
    174.7851,
  187.4331, 183.9528, 188.8189, 188.3152, 187.8625, 178.4524, 181.5308, 
    184.962, 190.7359, 188.6494, 185.921, 189.336, 186.7755, 181.8557, 
    177.9449,
  193.3789, 190.3285, 187.2268, 183.6884, 186.6902, 186.4588, 177.888, 
    182.8923, 184.4246, 180.8839, 189.0917, 190.6247, 189.9738, 187.9718, 
    183.4842,
  199.8055, 202.2712, 198.5254, 197.2434, 190.1997, 187.1487, 186.9246, 
    180.897, 182.9483, 181.7626, 181.9302, 181.2603, 186.4107, 184.9473, 
    183.3737,
  200.9528, 206.1272, 204.6245, 202.6836, 201.8865, 201.7699, 196.4392, 
    201.7543, 189.7981, 182.5363, 179.5485, 181.2569, 182.8735, 184.1633, 
    183.6538,
  209.9834, 209.192, 205.5868, 209.6667, 204.9581, 205.8777, 193.7304, 
    203.0969, 195.9376, 191.137, 195.5746, 181.9213, 179.3828, 179.2018, 
    179.5053,
  210.1353, 209.8971, 206.467, 210.0753, 208.1539, 201.2595, 193.6904, 
    189.6973, 190.9131, 185.5063, 187.9221, 181.465, 180.1774, 179.0254, 
    177.3906,
  193.5452, 194.5109, 194.4209, 194.8378, 189.3527, 188.5192, 185.0185, 
    177.2049, 170.2388, 165.0171, 163.4391, 159.7028, 157.4546, 157.9586, 
    156.0098,
  196.5618, 196.2551, 190.4772, 189.7025, 190.193, 191.6678, 191.5045, 
    188.5996, 179.9248, 177.2753, 174.7106, 168.4868, 164.5108, 159.7905, 
    159.7547,
  194.638, 196.2798, 189.2915, 184.0682, 180.6282, 185.6796, 192.4268, 
    190.882, 188.1469, 183.5108, 183.5476, 180.738, 176.2931, 171.5517, 
    167.0896,
  197.8166, 205.0684, 196.7597, 187.741, 179.4731, 178.6634, 181.7225, 
    188.6986, 191.8822, 191.0407, 188.1704, 186.6345, 182.4889, 175.5088, 
    174.0602,
  198.2188, 203.754, 207.8797, 199.0466, 187.4065, 178.0133, 173.5364, 
    185.1189, 193.6276, 189.2953, 186.4847, 188.0704, 185.9702, 184.8845, 
    180.5852,
  190.6474, 200.7119, 203.4954, 200.5741, 197.2249, 187.7793, 179.3575, 
    177.1801, 178.2027, 177.7739, 187.6695, 192.446, 188.3352, 188.1834, 
    186.3195,
  190.991, 191.8747, 197.2957, 198.2598, 202.4013, 203.6498, 194.6668, 
    184.0837, 181.5137, 181.6653, 185.4124, 188.1271, 188.4719, 190.5362, 
    189.3023,
  182.9642, 183.6981, 192.553, 192.0436, 197.5926, 209.5319, 211.4371, 
    204.1457, 192.6557, 181.7688, 178.3195, 179.3293, 184.0813, 187.4676, 
    189.1676,
  181.8637, 181.5878, 186.6069, 189.5163, 191.5157, 192.807, 204.5025, 
    199.0683, 191.7021, 187.6637, 185.1637, 176.9807, 178.3127, 181.2648, 
    184.2678,
  166.4474, 170.7079, 176.6206, 181.0146, 183.141, 184.1381, 184.3907, 
    184.3234, 183.9118, 178.2811, 180.7632, 175.1425, 175.1821, 175.292, 
    181.507,
  170.9951, 176.3864, 181.1867, 185.6512, 187.2139, 191.1738, 194.9611, 
    191.122, 187.505, 184.2131, 178.6134, 174.2045, 169.144, 166.2398, 
    163.0371,
  168.6696, 172.6027, 176.4006, 181.9088, 183.4083, 194.0686, 194.2991, 
    191.7407, 189.8429, 184.7371, 182.1753, 175.9844, 170.6271, 162.8195, 
    159.3493,
  170.0861, 167.8402, 172.4878, 180.5566, 184.1029, 191.7682, 192.6031, 
    189.0331, 189.2886, 185.713, 183.7565, 176.035, 171.1142, 167.7273, 
    161.4996,
  166.7607, 165.999, 176.0896, 190.1608, 187.3549, 186.8306, 183.4437, 
    183.5415, 185.5007, 187.5394, 184.7824, 179.5435, 172.3, 169.5328, 
    161.6663,
  170.5308, 190.5073, 207.0987, 203.9237, 199.9768, 191.0368, 181.3228, 
    183.2352, 185.1689, 176.2612, 178.5762, 182.6796, 174.7822, 170.7245, 
    163.9557,
  202.1693, 211.6776, 214.5526, 212.8448, 206.7327, 199.584, 189.4709, 
    184.4483, 180.5048, 178, 184.8602, 185.6691, 179.4287, 175.0048, 168.091,
  200.9852, 203.646, 209.6626, 204.4483, 208.6484, 202.9958, 201.3426, 
    194.245, 187.7283, 187.9081, 185.6488, 183.6006, 183.1209, 179.7031, 
    172.7433,
  160.1943, 174.6086, 183.6203, 183.6284, 184.6397, 190.2129, 200.7662, 
    211.206, 196.4279, 185.9926, 182.8776, 181.2562, 182.9316, 182.5243, 
    175.2576,
  155.6238, 165.0574, 173.861, 172.7699, 170.0208, 169.6957, 177.3113, 
    189.6948, 192.4549, 189.8443, 188.7967, 179.0156, 178.7287, 178.8162, 
    178.3978,
  163.821, 169.4422, 177.5611, 179.4589, 180.9984, 173.8019, 171.1379, 
    174.9388, 179.8671, 177.6945, 179.6306, 176.3815, 175.7674, 174.1035, 
    175.8919,
  173.9761, 170.9433, 168.9139, 172.957, 175.3272, 179.322, 183.0667, 
    189.217, 185.5069, 185.7988, 185.6699, 184.8867, 179.6684, 176.6664, 
    170.9432,
  174.564, 173.6158, 171.8421, 171.1468, 170.4611, 178.0225, 179.8922, 
    182.3411, 187.8089, 184.6557, 185.4592, 185.1967, 187.171, 181.7, 174.8967,
  183.4676, 179.2804, 176.2269, 168.7809, 171.0841, 172.8593, 172.8969, 
    175.7671, 184.9691, 189.1648, 185.0255, 185.3833, 185.0972, 184.551, 
    182.834,
  186.1531, 177.9675, 173.6805, 171.3141, 167.4457, 170.1649, 170.0259, 
    179.3563, 183.1828, 188.0283, 189.6531, 189.5164, 186.4077, 185.8473, 
    186.4215,
  178.619, 177.5958, 180.317, 187.3125, 188.1865, 183.7229, 183.1345, 
    187.4137, 190.4119, 187.9588, 189.8352, 192.7536, 189.4966, 188.4555, 
    187.3902,
  199.5958, 201.1477, 190.7292, 194.8851, 199.9876, 203.4756, 204.4056, 
    199.7377, 193.213, 186.0859, 189.7494, 191.9109, 190.5634, 190.6514, 
    188.3796,
  210.6659, 206.0981, 203.2759, 195.1476, 207.3604, 210.9804, 210.9209, 
    206.4044, 199.7215, 194.1551, 191.4779, 187.4481, 187.6948, 189.1311, 
    189.8216,
  180.3836, 184.0511, 189.2475, 195.7267, 198.7722, 200.1316, 191.5031, 
    192.2018, 193.7549, 191.7028, 186.2061, 184.3755, 182.5902, 182.9866, 
    185.2204,
  150.3053, 162.5483, 167.1646, 185.9125, 204.6383, 200.6617, 195.9242, 
    180.7821, 174.244, 179.1723, 182.3572, 180.572, 179.3466, 178.5072, 
    180.5997,
  163.1222, 172.2766, 179.1166, 201.5027, 198.384, 191.527, 186.8879, 
    176.4588, 168.822, 166.4916, 170.5522, 173.9369, 174.6774, 176.5042, 
    178.8535,
  187.468, 181.3252, 172.3279, 168.9456, 160.2596, 163.448, 167.8819, 
    173.3927, 177.1664, 183.6606, 185.9617, 185.8512, 176.9566, 171.7944, 
    168.3595,
  193.7198, 183.6902, 175.3087, 166.9447, 163.35, 162.7152, 167.5466, 
    170.8436, 175.2939, 179.5694, 185.5204, 187.096, 181.8233, 171.1909, 
    165.1284,
  196.6339, 186.1681, 181.7159, 173.2963, 168.3845, 167.7318, 165.2634, 
    169.2686, 173.7506, 176.729, 182.3, 187.5475, 179.7592, 176.4331, 166.4301,
  168.202, 168.3641, 172.8048, 177.9468, 173.3377, 169.6723, 165.2095, 
    168.5098, 174.1797, 175.0671, 181.1294, 185.349, 181.2084, 177.8092, 
    170.0101,
  163.0762, 161.8517, 167.2612, 170.3604, 172.2222, 166.6529, 171.7621, 
    172.5753, 178.0899, 172.6945, 177.1248, 183.6295, 183.9717, 180.6315, 
    173.417,
  192.039, 195.2359, 193.7854, 191.7515, 189.8394, 181.5246, 172.2704, 
    171.6801, 170.1765, 171.392, 179.4952, 184.5881, 183.3146, 180.0867, 
    177.9488,
  210.4074, 212.4534, 214.7941, 210.1601, 210.8736, 207.0144, 198.7915, 
    186.2612, 183.5438, 183.6883, 183.4155, 182.0804, 183.2549, 179.251, 
    177.5217,
  210.9323, 213.7947, 210.1346, 217.4707, 212.4225, 208.8701, 206.8582, 
    205.6968, 200.1453, 193.5967, 188.8528, 185.6625, 182.6559, 181.0528, 
    177.6094,
  210.9656, 214.3378, 215.7994, 218.0444, 215.4727, 209.5173, 207.1434, 
    201.1929, 195.6868, 194.1513, 192.9025, 187.7963, 181.4904, 180.4565, 
    177.8231,
  213.0766, 215.8465, 209.6788, 206.5231, 195.3648, 188.2145, 186.845, 
    190.1488, 187.0994, 188.0965, 189.8602, 187.2382, 180.9689, 179.5878, 
    174.4476,
  194.8555, 203.0503, 199.8906, 196.3454, 186.9354, 182.1518, 178.0423, 
    177.3517, 181.8477, 183.6989, 188.7491, 188.8363, 188.9824, 191.0364, 
    192.3882,
  196.3372, 192.9512, 194.0932, 193.8326, 185.267, 189.9087, 183.5253, 
    176.138, 178.3382, 182.9104, 185.6692, 189.8785, 190.1777, 190.4312, 
    191.1823,
  200.6285, 189.6073, 177.3503, 180.1066, 186.5087, 183.7227, 184.0933, 
    174.4476, 173.7854, 177.7881, 179.8506, 181.8683, 182.4713, 188.8798, 
    187.5495,
  194.4012, 187.5913, 178.5701, 177.685, 181.0848, 182.7728, 177.6051, 
    176.1762, 174.5686, 174.3793, 173.5903, 177.6192, 178.5571, 182.0818, 
    187.7985,
  193.539, 202.0384, 188.5733, 176.36, 170.6141, 177.7761, 176.6167, 
    176.8894, 178.9847, 172.6861, 168.541, 173.189, 177.2877, 180.2678, 
    183.2906,
  202.5933, 221.4307, 207.5448, 179.1573, 167.4173, 166.7058, 167.0955, 
    178.5692, 174.8004, 166.8243, 169.903, 172.562, 176.392, 178.9203, 
    181.3796,
  207.1799, 218.3813, 216.9678, 211.9812, 196.0112, 178.804, 169.547, 
    170.1274, 168.2135, 168.9051, 169.6283, 168.2316, 175.3535, 178.5935, 
    180.6621,
  218.7665, 217.3066, 218.3995, 220.1784, 217.9611, 203.0164, 181.0711, 
    177.4723, 175.6505, 169.9225, 166.9185, 166.3647, 172.3534, 175.1233, 
    179.606,
  214.1981, 220.6456, 217.2378, 219.9272, 213.1797, 207.0127, 195.5802, 
    184.1027, 173.0745, 169.0316, 167.5521, 167.5885, 170.2878, 175.9214, 
    180.9459,
  208.1366, 216.3656, 213.8476, 204.0291, 192.4827, 187.0121, 185.0988, 
    183.6396, 176.2014, 169.5215, 168.7293, 171.3245, 172.4548, 177.1901, 
    180.09,
  191.7419, 186.2571, 181.7882, 176.3015, 168.4169, 165.7953, 170.0126, 
    171.9245, 179.1095, 177.2927, 179.5728, 178.141, 180.0869, 174.1352, 
    174.3478,
  199.9294, 190.6165, 190.694, 179.3701, 167.4408, 170.7471, 168.4906, 
    173.9144, 177.0192, 178.1506, 176.4346, 178.4019, 177.0489, 172.8537, 
    175.1835,
  207.4193, 201.4024, 196.8356, 183.4293, 173.2626, 173.646, 173.6802, 
    170.4439, 173.5949, 174.7541, 177.3581, 173.3667, 173.6102, 169.8268, 
    171.6106,
  211.4085, 204.8984, 207.6392, 201.4775, 183.6618, 177.6876, 174.5361, 
    173.6881, 172.1139, 173.2654, 170.3277, 173.0399, 174.2377, 170.5974, 
    177.0813,
  221.1262, 203.4158, 213.1809, 206.0869, 203.1026, 183.9143, 181.4579, 
    183.6914, 180.903, 175.3434, 173.1759, 171.7834, 173.896, 176.8697, 
    185.0939,
  218.1419, 214.9327, 208.5983, 201.82, 199.5215, 195.8379, 182.5486, 
    180.3153, 177.268, 176.64, 178.7555, 174.6647, 176.0173, 176.9626, 
    183.3093,
  202.8385, 217.3463, 221.135, 203.6904, 195.6653, 194.4474, 195.0909, 
    183.9854, 178.5199, 183.659, 177.2494, 172.7683, 175.1467, 177.544, 
    188.3062,
  201.8344, 218.3994, 214.4901, 212.8411, 201.7678, 202.367, 199.2786, 
    198.752, 187.4089, 181.4128, 177.2801, 176.453, 174.5045, 177.3427, 
    185.2074,
  212.6017, 211.3826, 219.2709, 212.0651, 195.6221, 198.3009, 192.9984, 
    188.498, 186.0993, 184.5359, 182.2274, 180.7241, 176.7597, 178.5473, 
    180.3568,
  217.5199, 211.1701, 207.8267, 202.9643, 190.6611, 186.7148, 186.1938, 
    187.3647, 184.8801, 184.8463, 184.7648, 180.296, 177.424, 174.4404, 
    179.1041,
  194.5956, 174.7085, 167.3259, 165.5976, 161.5631, 157.644, 162.3848, 
    168.7565, 172.8748, 176.6428, 182.8895, 190.4568, 190.6579, 188.6509, 
    185.2728,
  206.8752, 182.0612, 166.9656, 162.2061, 159.4678, 161.727, 171.545, 
    181.6573, 181.8004, 184.8339, 185.8098, 195.2655, 195.5197, 184.9023, 
    178.8348,
  212.3283, 193.1465, 170.6207, 165.8626, 167.5186, 173.1093, 185.3353, 
    187.7108, 186.2874, 186.2487, 191.1878, 191.1426, 185.8855, 183.3801, 
    176.7938,
  215.0081, 199.1404, 183.7034, 174.5121, 173.3729, 181.0314, 180.789, 
    190.2742, 188.021, 184.6603, 189.9133, 186.4931, 181.207, 179.462, 176.014,
  213.0343, 202.5644, 189.2363, 178.8223, 178.0475, 181.2428, 188.7393, 
    184.7093, 185.1888, 182.0691, 184.7321, 184.9735, 179.5699, 178.7897, 
    175.5748,
  215.6955, 207.0263, 191.0228, 182.9282, 177.0388, 181.4142, 179.5642, 
    183.5247, 186.9886, 188.6591, 184.7519, 183.6156, 175.3759, 174.2714, 
    175.8428,
  219.7469, 207.0625, 192.2356, 184.7761, 178.5896, 177.292, 180.9476, 
    180.3098, 180.5456, 181.2554, 177.6621, 175.7739, 170.4616, 169.9967, 
    174.5609,
  220.4991, 210.5155, 201.5868, 188.9492, 179.8327, 173.4744, 177.0154, 
    182.2615, 184.2964, 180.5414, 180.5548, 174.874, 172.1887, 176.5495, 
    180.2452,
  221.1065, 216.2256, 205.2593, 192.8899, 186.6308, 181.1485, 181.497, 
    178.9241, 180.467, 179.4752, 177.1958, 176.2488, 177.3219, 179.9451, 
    185.6373,
  226.3563, 206.924, 206.4135, 194.6553, 185.7991, 180.0376, 179.8206, 
    184.094, 177.9917, 176.4969, 173.26, 175.334, 177.3441, 182.9352, 187.0312,
  171.197, 164.3833, 163.2176, 165.369, 168.5007, 166.8522, 166.8158, 
    180.064, 191.4901, 184.6717, 180.5326, 180.6636, 180.5561, 178.9751, 
    179.4201,
  178.4886, 171.4635, 174.3205, 182.8532, 180.7774, 173.5981, 166.8796, 
    175.5613, 185.8259, 183.2051, 184.4003, 188.4834, 187.3916, 182.808, 
    183.0976,
  180.9193, 181.1993, 184.3194, 190.5679, 189.7545, 176.2382, 172.0868, 
    176.3125, 181.4996, 183.036, 191.8704, 191.9502, 191.1071, 191.5621, 
    187.3787,
  186.2118, 187.6296, 195.0054, 197.5463, 188.1183, 185.3801, 175.9723, 
    179.6839, 180.1144, 186.1001, 192.7164, 193.7829, 193.8223, 192.091, 
    192.5299,
  187.309, 189.405, 200.2723, 201.4403, 202.7877, 189.8524, 192.3743, 
    186.8449, 185.9734, 190.5601, 192.4503, 193.3222, 192.952, 194.1419, 
    189.9418,
  190.4317, 192.2786, 195.1188, 205.4875, 211.1324, 210.3913, 202.7469, 
    203.9469, 201.7585, 200.1782, 194.9493, 194.655, 193.4579, 187.0476, 
    183.845,
  192.8028, 194.3836, 198.5182, 201.6464, 209.7506, 212.0816, 215.4922, 
    202.7339, 201.8455, 201.1452, 195.1731, 192.6686, 188.5477, 181.2259, 
    178.2781,
  202.175, 201.0174, 202.8888, 203.9556, 207.1086, 207.6344, 214.5611, 
    205.5533, 199.4555, 195.9303, 192.3593, 185.4325, 181.1214, 178.2279, 
    179.6075,
  204.1972, 201.444, 202.4429, 196.1664, 201.3338, 200.3114, 203.4073, 
    200.6906, 195.5022, 188.8413, 185.8732, 186.1036, 182.1511, 183.664, 
    182.6333,
  199.1332, 203.9206, 206.866, 201.0634, 201.1615, 199.8278, 199.6554, 
    199.6199, 194.6295, 190.5771, 188.2266, 191.1494, 189.7319, 188.2382, 
    189.9348,
  195.3734, 201.1696, 195.969, 194.183, 190.171, 186.3177, 188.173, 186.4463, 
    193.1582, 188.2651, 186.3093, 193.0541, 189.4306, 181.4644, 166.9055,
  202.832, 201.1681, 200.6843, 197.1251, 189.0069, 182.6447, 178.3502, 
    183.4562, 191.497, 192.4301, 185.638, 188.778, 191.1798, 183.2326, 172.673,
  210.5948, 203.6172, 202.6949, 196.5469, 187.104, 177.097, 181.2694, 
    190.2001, 191.0623, 184.1185, 183.8554, 182.2961, 184.8946, 186.9524, 
    178.201,
  216.2551, 214.6951, 212.6876, 200.5653, 187.4412, 195.7196, 188.1638, 
    189.1957, 186.6345, 180.2565, 179.6396, 179.353, 181.3102, 183.1789, 
    179.8736,
  223.2972, 218.3756, 218.0056, 218.8054, 204.6476, 200.2183, 206.1223, 
    181.4877, 185.3423, 183.5919, 180.0975, 178.5196, 182.405, 183.8219, 
    182.3238,
  225.869, 221.38, 222.2462, 222.1653, 218.8843, 202.9469, 197.0741, 
    203.0045, 197.5186, 194.2743, 184.9138, 181.8285, 182.9055, 182.2076, 
    182.9126,
  223.6087, 223.0316, 218.0009, 218.3619, 218.6912, 217.123, 205.1109, 
    199.2788, 197.2109, 197.152, 189.4112, 185.7605, 180.8535, 181.1551, 
    181.679,
  218.5858, 223.932, 223.6051, 214.9822, 215.3789, 212.845, 201.6196, 
    196.6245, 194.4825, 192.8337, 189.2824, 185.9077, 182.6125, 179.9205, 
    177.6567,
  207.0224, 222.0286, 226.0964, 197.0115, 198.9303, 196.7651, 196.628, 
    195.3004, 189.4705, 184.6161, 182.6182, 183.2798, 181.6389, 175.9881, 
    177.6087,
  186.314, 189.6746, 203.278, 200.6603, 199.2188, 196.2441, 194.7383, 
    194.4484, 186.5339, 180.8766, 178.8728, 181.8847, 178.3757, 177.5099, 
    178.6763,
  199.797, 201.7819, 199.4316, 200.8895, 196.1165, 192.9035, 189.4536, 
    182.3407, 177.5789, 171.15, 169.1264, 170.1316, 173.0433, 176.6358, 
    181.186,
  203.6119, 199.2973, 200.2505, 198.812, 195.7861, 195.1181, 194.6783, 
    186.3874, 184.0848, 180.6742, 177.3438, 174.9862, 178.2787, 176.0164, 
    175.9583,
  208.9002, 204.0729, 201.716, 197.0573, 193.5902, 185.952, 194.1217, 
    193.3698, 192.4736, 188.4555, 182.9837, 182.4489, 178.9464, 178.1537, 
    176.156,
  220.4574, 223.2654, 212.3555, 198.158, 198.8283, 202.355, 187.0896, 
    188.4617, 192.9265, 190.7422, 188.6771, 187.2672, 183.3596, 182.703, 
    178.0122,
  222.1016, 224.0761, 221.6834, 217.5455, 202.2222, 200.153, 201.8595, 
    189.1699, 189.8472, 191.1338, 191.1971, 189.9729, 186.6833, 187.3413, 
    183.0607,
  227.6292, 222.6831, 221.8184, 219.6743, 215.6598, 203.1287, 200.2948, 
    198.2095, 198.244, 199.3667, 193.9574, 195.0437, 191.759, 190.2812, 
    186.5719,
  224.3068, 222.0267, 221.3375, 220.1656, 222.4919, 218.7029, 203.6309, 
    199.7187, 199.4093, 197.5083, 194.3807, 196.8517, 197.3376, 194.0477, 
    189.6871,
  225.8552, 224.6564, 218.4799, 219.8759, 219.9884, 200.3281, 202.2436, 
    202.2102, 195.839, 191.5767, 190.5451, 192.4426, 194.8649, 197.3541, 
    192.9692,
  223.334, 224.3169, 208.2013, 199.5337, 200.817, 201.9631, 200.0153, 
    198.0043, 192.3457, 189.7561, 188.2343, 187.5383, 188.9801, 194.3206, 
    192.9981,
  203.1053, 203.6799, 208.9617, 200.9492, 198.719, 191.9781, 191.088, 
    192.2898, 189.2552, 187.9337, 185.1313, 186.7303, 186.0417, 188.3649, 
    188.6961,
  199.8121, 201.2456, 198.2047, 196.513, 182.3428, 173.0681, 171.733, 
    168.0191, 167.1481, 171.0089, 180.3289, 186.8919, 192.7164, 198.1297, 
    201.4737,
  208.2661, 203.9149, 202.3382, 200.6307, 197.3693, 182.6776, 172.637, 
    170.2557, 167.9324, 173.7899, 181.2374, 188.9809, 194.2839, 199.5469, 
    199.9757,
  210.1265, 212.5956, 206.024, 202.0464, 200.2056, 189.7281, 183.0624, 
    168.1035, 168.7167, 174.0857, 180.7965, 191.2182, 199.8374, 206.9182, 
    203.2074,
  229.635, 211.1904, 214.8066, 205.7059, 205.5246, 203.7896, 183.763, 
    175.4445, 172.0393, 174.9279, 181.5213, 193.0796, 199.5138, 203.4444, 
    203.0802,
  223.354, 227.434, 225.9752, 218.9784, 208.3983, 204.0699, 198.2151, 
    180.0085, 174.3687, 177.1745, 181.4429, 192.5242, 198.1215, 201.2132, 
    200.5358,
  208.81, 218.5958, 218.6597, 216.2645, 212.3411, 205.3796, 201.2736, 
    193.6904, 185.756, 183.2722, 182.8274, 189.1457, 194.7152, 195.2356, 
    196.6314,
  205.7084, 212.4816, 217.0057, 217.8616, 214.6037, 217.3271, 209.3491, 
    196.9566, 188.4582, 187.2294, 189.0522, 189.7774, 192.8277, 192.723, 
    193.8214,
  195.3238, 200.0783, 206.6588, 212.3006, 222.1564, 218.6227, 214.9471, 
    202.8846, 194.357, 191.4544, 192.7924, 192.2323, 191.6218, 190.3697, 
    189.6127,
  189.075, 194.7336, 193.115, 201.9235, 207.8447, 213.6391, 209.8791, 
    200.135, 196.0329, 191.9142, 192.7831, 195.1018, 194.3688, 190.0454, 
    189.6421,
  178.8668, 180.7314, 185.6809, 190.0342, 197.8311, 200.6312, 199.4927, 
    197.7561, 193.0638, 192.6045, 187.9501, 191.295, 190.9037, 193.7319, 
    193.6049,
  199.0569, 202.6416, 199.277, 194.7791, 185.3346, 175.0707, 171.3688, 
    171.6584, 174.5322, 177.4572, 189.0253, 193.4778, 190.882, 193.0443, 
    195.0684,
  206.8937, 205.077, 200.8874, 194.6149, 180.2122, 171.4185, 169.9152, 
    172.961, 177.0396, 180.0327, 189.0543, 196.7174, 197.4431, 194.0473, 
    194.4257,
  222.4707, 215.0526, 204.8285, 192.5821, 180.8043, 171.5994, 171.3153, 
    170.1019, 176.6763, 181.5168, 192.3235, 197.9685, 198.0709, 198.8382, 
    195.4235,
  226.6365, 221.5781, 215.7916, 189.6907, 177.6295, 181.5632, 172.7744, 
    174.0496, 176.5763, 184.6717, 193.5114, 199.5451, 198.4098, 198.5097, 
    195.2724,
  223.2429, 225.3949, 208.2448, 189.2372, 186.0022, 190.324, 187.9747, 
    177.2771, 185.3935, 189.4913, 194.5205, 198.5718, 198.9998, 198.6543, 
    196.3606,
  224.5451, 218.6613, 209.1096, 193.8911, 201.239, 200.9499, 191.5636, 
    193.3966, 191.1359, 197.2668, 197.2737, 198.3937, 197.9803, 198.2065, 
    196.5344,
  218.806, 219.4223, 209.5042, 203.4149, 209.3864, 209.2659, 208.8026, 
    196.7433, 195.7259, 198.5919, 199.0606, 198.4754, 199.0782, 197.8848, 
    197.6537,
  218.2696, 210.7349, 207.4343, 206.2764, 211.2095, 206.555, 211.9616, 
    206.1291, 200.2526, 199.0775, 197.8857, 197.522, 199.1892, 198.3925, 
    199.2221,
  220.0624, 206.8602, 209.8062, 214.4534, 213.5585, 209.8206, 206.3567, 
    200.4602, 199.167, 197.6586, 196.7328, 197.0872, 197.8378, 198.2511, 
    198.9724,
  212.5697, 208.12, 213.0477, 208.5536, 203.7413, 200.0699, 198.3721, 
    199.3784, 196.1056, 194.0419, 193.2001, 195.4277, 196.2104, 195.7525, 
    196.5425,
  181.2627, 178.2878, 176.9413, 179.0678, 175.5317, 175.9386, 178.195, 
    178.299, 179.172, 177.5467, 182.3519, 184.697, 183.0424, 187.611, 188.0748,
  196.9567, 194.4328, 189.652, 184.4459, 177.3373, 180.2624, 176.3796, 
    179.1051, 180.349, 177.9239, 180.5097, 185.9571, 187.0477, 186.1714, 
    189.4426,
  205.0443, 204.0752, 198.2661, 187.9885, 184.65, 180.7037, 178.1223, 
    176.4433, 181.2562, 179.7392, 188.0917, 192.3795, 192.1889, 195.7556, 
    195.5702,
  223.9456, 208.4402, 204.2251, 191.3521, 186.5237, 188.8437, 178.0118, 
    181.3486, 182.5305, 181.7208, 194.5328, 195.7482, 192.0765, 196.0988, 
    196.9969,
  211.8919, 209.3282, 202.9176, 202.0149, 193.0613, 190.1222, 187.3682, 
    179.7259, 189.4698, 191.0343, 191.281, 192.7299, 191.6322, 192.1467, 
    194.6327,
  208.5676, 206.6174, 208.3075, 207.2255, 198.3253, 194.0818, 189.652, 
    192.7358, 200.0106, 198.0837, 191.3377, 187.167, 185.2503, 186.9737, 
    187.9733,
  216.2635, 210.5245, 210.1439, 201.5357, 201.8145, 207.9079, 210.3428, 
    198.8392, 198.8951, 194.5245, 188.2225, 185.0184, 182.9709, 184.1383, 
    186.2497,
  222.84, 214.2724, 213.6237, 210.8629, 212.9106, 215.6727, 199.8415, 
    203.4465, 196.869, 192.2762, 188.9932, 186.6977, 186.403, 185.4148, 
    187.4777,
  219.905, 213.3136, 212.7732, 212.2942, 208.707, 210.271, 202.7314, 
    198.9398, 195.734, 193.5004, 192.6689, 190.953, 190.6144, 192.8928, 
    193.6334,
  210.2898, 211.1845, 206.9639, 202.0292, 200.2443, 199.0959, 197.9139, 
    198.8709, 194.9643, 192.4353, 191.7318, 192.8738, 195.6996, 193.0655, 
    196.021,
  190.5823, 179.0372, 175.1193, 170.6223, 170.2758, 173.5225, 180.9314, 
    181.4496, 179.7045, 179.82, 184.5379, 188.2639, 184.5707, 184.0839, 
    180.5591,
  205.0443, 193.041, 182.8089, 175.7015, 169.7554, 170.1872, 172.0442, 
    174.0654, 175.075, 177.4228, 185.1508, 190.6814, 192.1921, 183.2975, 
    179.2971,
  216.601, 200.7852, 193.1923, 178.6272, 175.181, 168.8753, 169.5983, 
    170.8048, 174.0173, 181.4078, 190.8843, 193.8074, 193.5394, 189.575, 
    187.7067,
  219.83, 222.5122, 205.5247, 188.306, 177.7879, 174.0697, 169.7207, 
    174.4902, 181.0359, 188.866, 194.7044, 193.2266, 190.2288, 190.6588, 
    190.4997,
  217.4789, 215.7915, 209.4003, 190.5259, 187.1957, 182.106, 190.4978, 
    182.0506, 184.2387, 187.3728, 187.8996, 186.7023, 185.689, 188.7645, 
    191.8169,
  218.8761, 217.2128, 207.9619, 199.7363, 208.9713, 205.4325, 200.7815, 
    206.5807, 198.0265, 195.7845, 181.3551, 179.0547, 180.2971, 181.6648, 
    185.2359,
  218.4905, 220.1732, 220.014, 216.0909, 215.8223, 216.1573, 212.4034, 
    200.4131, 192.9801, 183.9364, 177.0567, 174.661, 174.8334, 174.5272, 
    178.8994,
  217.5867, 222.0862, 219.9929, 218.8904, 215.1432, 213.892, 200.0455, 
    199.9202, 191.0638, 180.6071, 178.076, 177.2626, 176.0683, 176.9516, 
    176.9903,
  225.112, 218.2671, 221.8647, 207.8023, 202.6807, 199.7385, 198.1108, 
    194.9887, 189.0435, 184.1391, 182.9513, 184.3465, 182.832, 182.7359, 
    183.6455,
  224.7277, 217.4059, 204.74, 202.3323, 200.0887, 197.193, 194.6336, 
    195.6679, 188.8543, 181.8527, 181.0348, 185.6436, 186.0802, 185.8227, 
    187.2318,
  197.8028, 195.5686, 189.9723, 187.6948, 182.1245, 177.9415, 185.4049, 
    186.2199, 184.3384, 179.2358, 179.2672, 183.082, 178.6544, 178.8042, 
    176.1148,
  202.1614, 194.6644, 187.9958, 182.8189, 178.4135, 176.9373, 181.6903, 
    184.4016, 183.9948, 181.8925, 181.5004, 186.3402, 186.1068, 176.4785, 
    176.1016,
  211.9183, 202.3353, 188.3718, 181.1284, 178.2063, 174.9886, 179.9337, 
    184.5225, 180.9304, 185.1603, 187.0117, 187.1946, 180.9445, 180.3874, 
    177.3297,
  213.1831, 206.3433, 191.3357, 186.3673, 173.7928, 179.684, 175.6319, 
    179.218, 178.7881, 183.408, 187.2148, 185.4459, 180.8035, 174.3099, 
    174.8797,
  209.2901, 207.0281, 196.5032, 191.6565, 180.9893, 177.0768, 188.2785, 
    179.8835, 175.6913, 183.5629, 183.5975, 182.0508, 181.4005, 177.5293, 
    173.4691,
  205.2597, 208.6967, 205.8517, 204.2844, 199.1921, 193.8151, 193.2166, 
    202.5582, 195.2455, 191.364, 181.7968, 180.3696, 179.9172, 179.1025, 
    178.3813,
  212.7064, 213.5099, 216.0176, 216.9162, 216.1969, 216.8152, 209.4794, 
    198.4453, 190.7543, 186.0919, 183.5796, 179.0883, 178.6095, 176.9335, 
    175.9675,
  219.3443, 217.9579, 215.1366, 217.6015, 218.9309, 214.914, 210.0468, 
    199.2135, 188.4924, 182.032, 177.3127, 176.8214, 175.2201, 175.783, 
    176.9779,
  223.9405, 221.6421, 216.0594, 217.8581, 201.5609, 200.0446, 199.319, 
    191.8215, 185.1871, 179.1049, 177.4043, 176.2772, 175.8517, 175.0358, 
    176.5871,
  214.4781, 214.0224, 203.6649, 200.6969, 197.0946, 195.6637, 194.2949, 
    190.7038, 184.4178, 176.5382, 174.1634, 178.5075, 178.0492, 179.0451, 
    178.546,
  202.3568, 201.3032, 199.1195, 199.6137, 196.7598, 190.8554, 183.3017, 
    177.2131, 178.025, 177.6407, 174.7542, 176.0531, 174.9778, 179.2719, 
    176.9421,
  203.6206, 201.7196, 200.6154, 197.4436, 191.0792, 183.2524, 175.9746, 
    175.221, 176.2099, 177.7408, 175.8166, 180.8487, 186.4651, 176.7982, 
    176.2988,
  214.2226, 205.4051, 200.3831, 198.4614, 195.6671, 182.9622, 180.097, 
    173.6838, 172.8908, 176.5627, 181.9656, 186.978, 189.0941, 189.6056, 
    179.7652,
  214.3607, 208.2127, 205.2987, 203.8618, 195.7134, 190.8942, 179.423, 
    178.0158, 177.9725, 179.4106, 184.6749, 187.5381, 189.8443, 183.3077, 
    172.9237,
  220.3593, 204.2152, 205.215, 204.9453, 196.9608, 185.1863, 192.1759, 
    176.3766, 169.3092, 177.2884, 183.7947, 186.1604, 185.6435, 177.728, 
    172.5074,
  219.6887, 222.0261, 215.7732, 209.981, 206.1807, 197.5449, 186.2921, 
    197.8071, 191.4539, 188.2041, 182.1609, 182.7903, 180.3931, 176.7356, 
    171.5107,
  213.303, 213.7867, 219.4842, 217.421, 208.0836, 217.5483, 203.8165, 
    192.8837, 188.537, 186.7301, 184.4674, 182.2919, 179.6334, 176.7218, 
    173.5821,
  202.377, 210.3834, 213.5296, 214.613, 215.0053, 215.9208, 208.9186, 
    195.9329, 187.501, 184.1306, 182.5483, 181.298, 178.6775, 177.0682, 
    176.6568,
  187.2005, 193.8458, 207.3526, 207.3667, 211.3207, 203.5164, 196.9201, 
    187.4334, 183.0964, 181.2111, 180.0664, 179.2795, 178.1126, 178.2882, 
    176.6134,
  183.3078, 183.496, 188.4079, 194.6811, 195.7603, 194.6539, 191.4745, 
    186.226, 179.8941, 174.872, 173.5787, 175.6979, 174.5893, 174.4631, 
    174.4561,
  204.2265, 203.9353, 201.111, 198.7422, 192.8348, 190.0801, 191.4442, 
    188.7973, 190.5993, 186.652, 184.7131, 184.3015, 186.156, 182.2953, 
    180.6136,
  204.3822, 203.0076, 199.9568, 195.8763, 188.188, 185.6854, 186.6997, 
    186.6389, 186.5883, 189.7133, 185.9768, 189.3271, 189.514, 174.7497, 
    170.5341,
  207.6176, 205.5175, 200.5558, 196.0251, 193.9175, 179.1741, 184.2713, 
    183.7287, 183.3114, 186.5471, 186.2744, 186.7089, 188.0637, 186.6861, 
    183.1501,
  215.7973, 209.713, 206.266, 201.6098, 196.9098, 200.2535, 174.9546, 
    181.2624, 180.3372, 179.824, 183.2563, 183.7608, 186.0245, 187.0779, 
    183.3072,
  211.8937, 199.1488, 199.8114, 211.7841, 196.2314, 196.942, 199.2883, 
    172.7166, 173.515, 178.7057, 177.9771, 180.2744, 183.221, 185.2679, 
    186.7528,
  219.2129, 201.5728, 197.4408, 203.9528, 205.7403, 199.2395, 195.3326, 
    195.9047, 185.2383, 178.5098, 175.2565, 178.4603, 180.9575, 184.4456, 
    185.3201,
  216.8781, 222.4372, 220.1246, 199.5465, 208.7652, 203.6681, 199.6637, 
    190.8855, 184.9431, 182.2718, 179.3663, 176.5162, 177.6907, 179.113, 
    182.0443,
  215.674, 217.8851, 220.6354, 216.5362, 196.3068, 201.5505, 201.5777, 
    191.3987, 185.1316, 181.1344, 177.5387, 176.5011, 175.058, 175.5397, 
    177.7036,
  220.5876, 215.1028, 218.5635, 212.8132, 201.0471, 202.9637, 195.8556, 
    187.7738, 182.8208, 179.5112, 176.6315, 174.9484, 174.3412, 175.8395, 
    177.9473,
  217.0534, 209.3171, 214.9909, 199.6217, 193.5389, 189.7075, 188.0836, 
    187.2879, 181.653, 175.1739, 173.1258, 175.4195, 175.2219, 176.29, 
    175.7079,
  181.5276, 187.1077, 184.8672, 188.764, 187.318, 184.8295, 190.019, 
    189.6926, 191.3616, 182.8333, 181.0008, 184.31, 183.3081, 179.5677, 
    176.9631,
  196.6148, 198.0101, 195.3923, 192.8048, 185.6138, 181.9079, 185.553, 
    186.0545, 187.1424, 189.9879, 182.2993, 186.6708, 187.7082, 171.7494, 
    168.5622,
  208.8716, 203.6399, 199.3414, 195.1041, 192.1614, 174.9433, 180.7309, 
    182.5345, 182.6243, 185.6282, 186.7291, 186.6688, 187.6447, 186.0008, 
    177.1906,
  215.0587, 206.5278, 205.587, 200.6997, 195.8939, 198.1754, 173.1338, 
    178.755, 182.1991, 180.9707, 183.5453, 185.1673, 186.6604, 185.9279, 
    180.8138,
  224.4995, 201.5605, 200.2026, 202.191, 195.1663, 196.7291, 199.8976, 
    171.2095, 172.8728, 179.36, 180.2621, 182.2935, 184.6636, 185.1378, 
    184.4669,
  222.3416, 201.7448, 203.2927, 199.8149, 199.7574, 195.9923, 195.9765, 
    195.348, 183.953, 180.5874, 178.4831, 180.9002, 182.3045, 183.1053, 
    184.2743,
  219.4342, 219.4457, 202.3115, 200.8956, 197.8514, 197.3494, 194.0029, 
    185.0003, 179.7287, 180.2375, 179.3129, 180.1497, 180.2362, 179.5888, 
    181.9008,
  222.1038, 221.2808, 216.9879, 211.7312, 200.6143, 194.1405, 194.5982, 
    181.9982, 179.2066, 177.8836, 178.6496, 179.2902, 178.5396, 178.9212, 
    181.222,
  220.092, 221.8883, 215.5396, 197.0444, 194.7097, 190.2355, 186.7475, 
    178.5477, 176.328, 176.1364, 177.3678, 178.2763, 178.2287, 178.7737, 
    179.8362,
  219.7522, 218.337, 205.4196, 195.5247, 186.6022, 181.2369, 179.6496, 
    179.1925, 177.9537, 173.7295, 171.9262, 176.0262, 176.6542, 176.6331, 
    178.3445,
  180.7321, 180.2982, 177.2731, 176.7409, 174.4086, 174.2065, 174.4981, 
    176.175, 179.8864, 177.6496, 177.3698, 179.8712, 177.2785, 175.3249, 
    170.7048,
  183.326, 179.5008, 177.3912, 178.6249, 176.1282, 174.8792, 179.7917, 
    180.4505, 182.9612, 186.0388, 179.6237, 184.3382, 185.7749, 171.9733, 
    170.0372,
  199.4625, 191.713, 186.6339, 185.7827, 187.5058, 173.5946, 178.7959, 
    181.2462, 182.55, 184.6491, 185.0254, 185.0801, 186.7584, 186.6923, 
    178.0689,
  212.9232, 206.8423, 203.4625, 200.4789, 195.5, 196.5443, 173.6529, 
    178.4517, 180.9633, 179.3116, 181.7443, 183.9112, 186.4589, 186.7536, 
    182.1709,
  215.7653, 214.059, 204.1934, 197.3044, 194.9107, 197.6663, 199.1387, 
    172.894, 169.7666, 175.2351, 178.6077, 181.7775, 185.1346, 185.5034, 
    185.619,
  217.5457, 214.5767, 202.9972, 201.7875, 198.9015, 196.1884, 197.4584, 
    198.767, 187.5264, 181.8811, 175.6102, 179.6997, 182.5374, 183.7088, 
    184.358,
  220.1148, 218.3965, 215.0846, 212.0027, 211.8445, 203.5704, 194.859, 
    190.6834, 184.9395, 181.6562, 178.7617, 178.1369, 178.305, 179.5213, 
    181.035,
  209.9906, 203.7852, 198.08, 196.3765, 197.485, 203.3499, 198.5914, 
    188.5816, 183.8653, 179.4625, 177.1316, 176.4005, 175.4971, 177.7071, 
    181.2147,
  209.8544, 201.6188, 191.3275, 185.5189, 187.6454, 193.2167, 193.3138, 
    187.1429, 182.5408, 177.6745, 176.2299, 175.2287, 174.8148, 175.5471, 
    177.2943,
  197.9276, 195.7261, 182.787, 181.6879, 184.2368, 186.9417, 188.5193, 
    187.0046, 180.2757, 172.0553, 170.1284, 173.7448, 171.268, 170.6713, 
    171.7303,
  174.1403, 177.652, 169.7721, 166.5591, 158.1076, 161.6245, 163.6142, 
    166.1344, 168.6401, 168.1886, 167.1174, 166.4598, 168.0479, 169.8888, 
    170.1189,
  174.6875, 169.1498, 166.6902, 162.0888, 162.8303, 161.3598, 160.4452, 
    164.0219, 166.8204, 166.7691, 167.7434, 170.1992, 173.5139, 171.2355, 
    170.1209,
  189.7098, 176.4777, 169.0679, 167.0823, 164.4296, 162.8756, 160.8504, 
    165.0672, 166.8017, 169.2475, 174.8855, 177.5492, 180.0211, 182.2953, 
    177.5696,
  207.0546, 192.2872, 190.9906, 180.1647, 172.8395, 172.2541, 163.4881, 
    167.9035, 172.3878, 174.1495, 177.8393, 181.8508, 185.4793, 186.3904, 
    183.8161,
  220.7477, 205.9878, 200.8925, 208.444, 193.4014, 189.1732, 189.8909, 
    170.8614, 168.5211, 173.4047, 177.0094, 182.7612, 185.3516, 186.7373, 
    187.4113,
  223.4205, 211.1638, 208.5799, 208.2674, 202.4673, 196.65, 197.2749, 
    199.0772, 186.8986, 181.353, 176.8004, 181.0265, 182.8509, 184.2948, 
    184.7134,
  205.3863, 221.8398, 223.4176, 213.3462, 208.9752, 204.6768, 198.7218, 
    191.1293, 185.2413, 183.3642, 181.4797, 179.5028, 179.3192, 180.6995, 
    180.7307,
  182.1926, 206.1967, 208.9126, 211.0399, 217.2932, 213.361, 205.0248, 
    190.1253, 185.1965, 182.2708, 179.9452, 178.7614, 176.8527, 177.0379, 
    180.1426,
  191.6264, 191.9969, 199.5299, 201.6374, 212.102, 203.062, 193.7051, 187.31, 
    182.9162, 178.0486, 175.1608, 173.8268, 172.7789, 172.1434, 178.6772,
  205.1578, 202.2347, 197.7755, 198.3329, 191.116, 184.3563, 178.0921, 
    177.284, 172.5321, 169.0066, 169.9273, 170.0058, 171.3513, 170.116, 
    172.4123,
  191.8797, 172.4679, 165.78, 162.128, 161.4488, 168.0554, 169.4108, 173.097, 
    178.2959, 182.2269, 181.7848, 177.8884, 173.0213, 169.1976, 171.8897,
  194.7186, 171.941, 162.9502, 160.5026, 160.5179, 164.1039, 165.4049, 
    168.7602, 173.2535, 178.7719, 180.7983, 176.8419, 175.5257, 170.7876, 
    167.9316,
  208.8365, 177.9945, 163.9677, 160.404, 161.0271, 163.6497, 167.1552, 
    166.1893, 169.1266, 172.8715, 172.0888, 173.6548, 174.9678, 172.8487, 
    173.4129,
  221.286, 207.6732, 174.8444, 169.0141, 163.8445, 161.6085, 167.9532, 
    168.5948, 174.9326, 174.7695, 174.4425, 175.9934, 174.272, 171.6768, 
    168.903,
  215.6852, 222.0273, 190.5289, 181.1621, 170.9537, 174.5095, 177.8293, 
    177.7846, 175.4522, 178.3082, 180.6812, 182.4458, 180.2531, 178.4639, 
    177.3367,
  212.0103, 222.1426, 202.0755, 194.7847, 188.3327, 184.0757, 187.7715, 
    193.0453, 185.0636, 181.2436, 180.1984, 183.5699, 183.7933, 180.7124, 
    178.0194,
  194.1331, 222.1178, 211.9075, 207.2153, 202.4243, 201.5385, 196.8145, 
    191.7554, 187.4535, 186.0908, 183.0766, 182.7047, 183.4109, 184.9086, 
    182.7532,
  199.9136, 214.1159, 211.2629, 205.8051, 207.4335, 205.9065, 204.5709, 
    196.3447, 195.386, 190.2249, 184.9384, 182.2933, 180.491, 179.8389, 
    185.228,
  203.151, 207.7253, 182.7829, 187.4811, 185.6253, 196.5609, 196.4506, 
    194.1934, 192.6182, 190.8574, 187.6796, 182.9501, 178.4992, 176.2565, 
    177.8235,
  194.2058, 183.5125, 174.7105, 173.3927, 178.038, 184.2901, 187.7076, 
    188.7746, 187.6971, 184.7359, 187.0724, 181.7457, 174.6925, 170.1038, 
    169.5671,
  201.6525, 201.8776, 195.3951, 186.5685, 188.6191, 190.4816, 194.8047, 
    194.9406, 192.3328, 190.1147, 192.7289, 200.7106, 204.5211, 208.4085, 
    197.5681,
  201.6096, 201.0307, 197.2174, 186.3891, 184.9546, 184.3486, 183.5989, 
    186.6424, 184.5232, 189.3092, 189.6463, 194.2046, 198.2745, 202.8293, 
    204.3876,
  202.8183, 202.6517, 199.4008, 187.7103, 182.0743, 179.1118, 180.3832, 
    181.2365, 183.2868, 183.7384, 184.5596, 186.5099, 190.2519, 196.1053, 
    196.9893,
  204.7243, 212.0728, 205.2871, 193.9684, 179.3449, 179.0198, 174.2656, 
    178.2351, 180.0626, 180.2428, 180.8884, 178.7112, 180.9897, 185.8235, 
    190.2125,
  201.2288, 208.1985, 206.4192, 197.8872, 180.7469, 176.5979, 180.0667, 
    178.0385, 177.8094, 179.615, 185.4983, 185.9868, 182.2399, 176.5291, 
    177.9191,
  198.4319, 204.9152, 204.819, 198.2235, 179.0267, 172.8015, 180.3136, 
    187.6078, 187.7601, 188.3226, 186.6101, 191.2196, 192.4153, 185.358, 
    174.9696,
  196.3313, 207.4481, 212.594, 192.8587, 180.3057, 177.6377, 186.9452, 
    193.6792, 195.2596, 194.1264, 188.4051, 186.9734, 189.0879, 192.0139, 
    186.8131,
  205.4941, 214.2446, 219.0854, 184.8709, 178.1594, 183.7851, 194.8868, 
    196.7426, 199.3704, 197.897, 196.3916, 186.4456, 183.6415, 184.906, 
    189.3171,
  212.9934, 215.1125, 202.8448, 189.9155, 188.6364, 194.2937, 195.8987, 
    194.8225, 193.9744, 192.3344, 190.8111, 189.9198, 186.9812, 183.1738, 
    182.9016,
  208.3536, 213.4464, 190.9846, 180.6644, 185.1595, 192.678, 194.8181, 
    194.1691, 190.8195, 188.1794, 190.9153, 188.512, 184.376, 181.656, 
    179.4535,
  192.1277, 190.8304, 194.226, 199.1403, 203.5314, 196.5553, 199.3831, 
    204.1155, 208.5618, 207.1992, 204.5284, 205.5101, 202.1098, 192.3255, 
    185.5832,
  194.411, 191.5038, 189.7686, 200.1048, 202.9639, 191.009, 194.8356, 
    198.2501, 203.9086, 207.1817, 203.7286, 203.4154, 204.2614, 204.5851, 
    203.6009,
  197.9759, 191.067, 186.7546, 194.0473, 203.1536, 192.6702, 190.7614, 
    193.4689, 196.0272, 198.8466, 202.075, 205.8061, 204.0972, 206.0494, 
    206.3428,
  198.4609, 192.2543, 194.154, 197.1667, 205.8589, 205.9644, 189.6186, 
    187.0266, 192.2674, 192.0637, 195.4112, 201.3785, 204.8433, 206.3019, 
    206.0459,
  197.223, 194.2936, 188.3133, 200.1915, 198.3463, 198.2781, 202.3094, 
    185.6572, 180.6397, 180.5973, 187.2497, 193.7769, 200.201, 203.6154, 
    205.2465,
  187.8895, 179.9904, 185.0038, 196.8508, 197.2874, 195.8904, 196.7046, 
    193.2522, 184.1376, 183.5846, 184.2147, 189.0005, 193.0483, 197.8174, 
    202.0299,
  181.8339, 177.4182, 181.6439, 191.5338, 198.2796, 198.658, 192.9967, 
    185.5621, 183.4396, 189.3827, 189.8832, 186.6895, 187.4138, 189.7169, 
    195.6015,
  178.8888, 173.9389, 186.2757, 187.43, 193.2697, 196.6568, 187.0721, 
    183.9836, 185.5888, 188.9262, 193.2211, 186.0089, 183.0291, 185.0291, 
    189.8886,
  177.1645, 176.2365, 185.967, 183.1008, 191.8534, 189.7155, 183.493, 
    180.3344, 184.4435, 188.8566, 192.2835, 186.8151, 182.3428, 183.0292, 
    186.1,
  173.2892, 180.519, 181.6652, 186.0594, 185.4473, 182.1912, 181.6501, 
    182.3462, 182.6513, 188.1457, 190.6801, 188.6739, 181.3195, 180.9385, 
    182.8487,
  186.4416, 182.6546, 177.6624, 176.2234, 178.1267, 176.3343, 178.0038, 
    186.4982, 197.7954, 197.6635, 198.4101, 200.4038, 207.2717, 197.8835, 
    189.271,
  187.1, 182.8798, 178.8649, 175.6482, 177.7782, 174.5121, 177.1832, 
    182.3715, 190.1238, 198.4158, 200.4604, 198.9971, 207.0303, 202.2549, 
    199.2244,
  202.2327, 191.4902, 182.3328, 178.8737, 180.6938, 181.0517, 175.3644, 
    177.5543, 182.7474, 188.8247, 195.1125, 201.4209, 204.2873, 204.7121, 
    199.7551,
  216.7649, 199.4703, 184.3308, 178.284, 177.5201, 181.9483, 180.8586, 
    179.0506, 179.1778, 183.743, 189.3917, 194.0828, 196.9195, 198.7012, 
    198.5348,
  216.4598, 212.0903, 197.9039, 182.6912, 177.7621, 180.2496, 186.1127, 
    188.7821, 192.5664, 179.9433, 183.0609, 187.0788, 192.9522, 194.4037, 
    196.3439,
  208.8405, 210.772, 205.0301, 189.7238, 180.4364, 181.5788, 185.3478, 
    188.9689, 185.581, 184.0758, 180.0471, 184.0789, 187.8509, 190.8141, 
    194.2983,
  192.4556, 195.8193, 198.6141, 194.0206, 183.2027, 185.1877, 180.425, 
    180.1148, 186.5477, 186.2835, 182.4242, 181.1414, 184.3757, 186.8034, 
    192.6277,
  193.2009, 186.3424, 185.5117, 189.6018, 192.0114, 185.6877, 181.7076, 
    182.6563, 181.2923, 184.276, 182.2435, 184.8354, 181.7989, 184.9717, 
    191.6187,
  197.8976, 187.1821, 183.2541, 184.2041, 180.8023, 183.4249, 181.4732, 
    179.5973, 177.922, 180.7039, 179.7657, 185.5637, 180.59, 183.9715, 
    189.6538,
  201.2573, 189.7372, 182.6545, 179.3111, 177.1869, 175.3123, 174.6021, 
    181.0791, 178.284, 174.3518, 178.3907, 182.9357, 179.5763, 181.7564, 
    186.1342,
  209.422, 206.7191, 204.5699, 204.4464, 193.1169, 183.9183, 174.8185, 
    169.5212, 169.8159, 169.4341, 175.1407, 181.3226, 191.8552, 195.8062, 
    201.0238,
  209.5802, 206.1155, 205.8176, 201.3164, 188.5312, 179.5703, 172.4389, 
    166.2462, 171.6452, 170.2886, 177.4569, 179.2085, 189.9144, 191.6799, 
    197.7344,
  210.9085, 206.6048, 206.4819, 199.8777, 189.6939, 176.1031, 170.0983, 
    170.9682, 169.0779, 170.1573, 172.6125, 179.4348, 187.1723, 194.3035, 
    188.793,
  219.2169, 212.1106, 207.1633, 199.3451, 187.2048, 174.6897, 169.1881, 
    169.9559, 169.3503, 171.3316, 171.7424, 178.0132, 183.6144, 188.4992, 
    188.3344,
  223.9728, 222.1454, 213.8666, 198.1226, 182.3363, 171.0794, 167.6697, 
    168.5391, 171.6953, 168.1019, 170.8697, 176.4021, 182.1919, 186.85, 
    190.2881,
  219.9579, 221.693, 215.6719, 201.8702, 179.6665, 174.8329, 169.0797, 
    165.9514, 167.1994, 168.1119, 169.7775, 177.1544, 181.4188, 185.0549, 
    188.9249,
  223.1821, 219.5367, 220.6396, 205.0846, 175.8131, 169.084, 170.0201, 
    169.1106, 170.2573, 170.8611, 173.0435, 177.0536, 179.6823, 183.5549, 
    189.052,
  226.9763, 225.1246, 218.594, 203.1095, 176.895, 169.2182, 169.0666, 
    172.0283, 169.6297, 172.5907, 173.3745, 176.1488, 177.414, 182.8257, 
    189.3158,
  227.4112, 220.5415, 214.9541, 200.3667, 180.3908, 169.5089, 168.3082, 
    168.5568, 169.4378, 170.359, 172.3161, 174.9566, 177.7767, 182.7306, 
    187.3366,
  223.986, 214.3238, 200.2357, 201.898, 189.6801, 175.0623, 167.1596, 
    165.7115, 169.1655, 167.7475, 169.6653, 175.0422, 177.9524, 181.1494, 
    185.0252,
  177.7808, 187.2497, 187.1118, 191.1398, 192.1384, 191.0068, 198.3058, 
    195.1664, 186.5433, 177.2551, 170.7641, 166.6559, 165.8177, 170.7195, 
    175.9651,
  179.9859, 182.7905, 181.7752, 188.4994, 192.274, 188.7237, 193.4153, 
    191.9776, 185.0021, 177.4688, 167.6414, 164.9576, 163.1899, 166.2775, 
    169.1413,
  183.1883, 187.4147, 184.9257, 195.498, 196.5056, 186.8245, 189.8645, 
    186.049, 178.2227, 170.3313, 161.6859, 161.2063, 162.8366, 167.6788, 
    170.1672,
  181.8501, 188.5013, 189.8258, 193.6138, 197.4038, 201.24, 188.7817, 
    182.4833, 178.2656, 168.3593, 163.0038, 159.6824, 159.8563, 164.3938, 
    170.3569,
  183.3203, 190.7544, 195.271, 194.3314, 195.6134, 202.3792, 194.5072, 
    180.3673, 175.1871, 164.1241, 160.6236, 158.9994, 165.4525, 170.1677, 
    175.743,
  185.1218, 196.1248, 205.6074, 198.0473, 205.534, 198.6898, 191.2049, 
    176.4573, 168.2779, 165.5106, 161.9649, 161.4668, 163.4334, 169.2535, 
    179.5417,
  197.0657, 198.9782, 211.1451, 204.6885, 212.4112, 198.0465, 184.8051, 
    173.161, 168.7745, 163.9112, 162.234, 165.4418, 166.9627, 175.0854, 183.64,
  199.4532, 214.2532, 224.0986, 217.8399, 210.2823, 197.8576, 175.9353, 
    173.7687, 167.1243, 165.5179, 164.5124, 167.226, 171.6023, 177.6644, 
    185.5881,
  226.2233, 228.9855, 217.1336, 218.9796, 200.749, 184.5674, 173.0771, 
    170.5001, 167.9747, 167.3706, 168.6726, 168.5701, 173.6382, 181.1239, 
    185.5519,
  230.1905, 226.9771, 221.9065, 212.4043, 196.9157, 174.5933, 170.3761, 
    170.2577, 167.0728, 168.6066, 167.5488, 169.6739, 176.6584, 180.6081, 
    183.6328,
  175.4584, 188.2339, 194.165, 191.8641, 189.4005, 185.4291, 185.6629, 
    190.3109, 189.0249, 188.8349, 186.7469, 187.566, 185.6886, 185.4733, 
    187.384,
  192.2849, 201.02, 199.7946, 192.4526, 188.6829, 188.3526, 187.7222, 
    187.3619, 184.7169, 184.0461, 184.2112, 187.9948, 184.7512, 181.4653, 
    184.0092,
  206.571, 202.4653, 198.9588, 195.8322, 191.0052, 188.9903, 183.3024, 
    183.1047, 182.1681, 183.1865, 186.5293, 185.7953, 182.4896, 179.5032, 
    184.6703,
  209.0897, 208.2248, 200.5569, 196.785, 189.3008, 189.8422, 179.2347, 
    179.648, 179.5033, 183.806, 183.2845, 182.448, 177.4642, 175.709, 174.9501,
  214.6229, 209.321, 202.3601, 196.086, 188.4903, 187.882, 187.8197, 
    182.1058, 177.1012, 180.2513, 180.6781, 179.7039, 172.29, 169.7612, 
    167.969,
  217.5185, 209.9171, 203.8099, 198.2489, 187.6535, 189.2487, 190.4721, 
    195.6792, 187.517, 185.1481, 177.8391, 173.5447, 168.9726, 166.0794, 
    163.6357,
  214.5037, 204.2678, 210.89, 198.2039, 195.2577, 200.0091, 197.0963, 
    190.4293, 186.3372, 180.5367, 173.5459, 167.9129, 161.9869, 159.0444, 
    160.6872,
  219.9657, 217.2604, 209.9165, 209.7764, 216.5612, 208.8831, 189.0681, 
    184.5278, 177.6165, 172.2974, 166.1186, 161.5255, 158.6023, 159.0933, 
    161.6066,
  223.997, 217.6409, 221.048, 211.1664, 210.6879, 186.8392, 178.0889, 
    176.2238, 169.934, 165.7708, 163.102, 160.2863, 160.5039, 159.8845, 
    164.4415,
  218.3812, 218.3553, 215.1566, 204.6494, 192.0743, 177.0975, 173.574, 
    173.0873, 168.036, 164.2487, 163.2917, 160.8365, 161.1642, 166.3965, 
    170.1999,
  206.1765, 204.1543, 204.3807, 203.4323, 201.4415, 197.4061, 195.6129, 
    195.7228, 197.8419, 197.8883, 197.89, 196.7553, 195.676, 190.7888, 
    186.5936,
  209.8355, 208.9012, 206.7326, 202.5564, 200.614, 195.4823, 193.996, 
    192.6768, 194.7986, 193.4258, 191.9444, 191.7768, 189.8136, 182.967, 
    183.5834,
  214.6915, 209.7609, 205.426, 202.7356, 200.6813, 191.8138, 192.539, 
    189.2757, 189.6126, 190.822, 188.3038, 186.5623, 183.9077, 179.2395, 
    179.7404,
  218.7212, 220.2169, 214.6793, 201.7687, 198.9868, 199.4737, 187.6509, 
    188.101, 186.5, 185.8032, 183.6206, 181.2951, 177.0575, 173.9221, 176.1809,
  220.9061, 222.4162, 216.6557, 204.5893, 197.2962, 192.8881, 196.8743, 
    180.1994, 181.2935, 180.0954, 180.1652, 179.7982, 175.6273, 174.9317, 
    176.0736,
  223.675, 220.0511, 212.2786, 206.9741, 200.7177, 191.2416, 189.2952, 
    189.7969, 189.7028, 184.6666, 179.9044, 180.1325, 178.013, 176.1462, 
    179.3594,
  219.4816, 223.6316, 210.7162, 208.3869, 207.2451, 193.9574, 190.4064, 
    187.9931, 189.067, 190.0562, 186.1892, 181.8128, 179.4178, 178.62, 178.763,
  214.8067, 216.2103, 209.4253, 200.4069, 207.2391, 200.3663, 188.8402, 
    186.4552, 186.4579, 187.1601, 185.7038, 179.7189, 176.7205, 175.9194, 
    170.1212,
  210.0465, 208.5195, 211.261, 216.0239, 211.0324, 197.7082, 188.1933, 
    184.471, 183.261, 182.3387, 179.4912, 175.9525, 172.0383, 169.9188, 
    162.4115,
  207.614, 204.1844, 203.0097, 202.194, 194.9243, 192.6925, 188.6157, 
    186.1813, 183.3391, 179.0205, 175.343, 171.6695, 168.2728, 164.1575, 
    162.7574,
  201.2073, 202.5183, 201.5204, 198.6586, 195.8504, 188.038, 188.2944, 
    187.0298, 183.7845, 183.9623, 181.3068, 181.9502, 183.7874, 189.6862, 
    192.218,
  199.9692, 202.4924, 202.799, 199.5121, 194.6779, 187.4271, 187.0413, 
    187.8912, 187.7009, 186.1497, 181.9887, 181.7605, 186.0166, 185.1205, 
    191.6568,
  200.4354, 201.6213, 202.6483, 201.7889, 200.0364, 186.2268, 188.2144, 
    182.816, 185.0643, 186.1322, 186.8597, 185.6998, 188.8878, 193.4686, 
    194.2547,
  200.8542, 206.053, 203.5512, 205.0079, 201.7583, 199.9458, 183.8261, 
    186.1957, 186.6254, 186.2153, 185.6448, 188.6731, 190.611, 194.0893, 
    195.4149,
  191.1793, 197.434, 197.9363, 204.4181, 203.8045, 201.7204, 199.5818, 
    179.2429, 185.9633, 188.7621, 185.8773, 188.2806, 188.8226, 193.2107, 
    192.9886,
  182.2586, 190.9751, 190.9045, 205.6993, 205.6288, 201.0269, 198.7921, 
    196.4053, 193.0249, 188.8237, 187.5978, 187.2474, 188.7806, 189.9819, 
    191.0394,
  178.0202, 188.1959, 185.8291, 200.0192, 210.4141, 206.412, 198.5726, 
    193.8051, 192.5863, 193.897, 192.9697, 190.9809, 190.5922, 190.3668, 
    190.3596,
  176.6122, 173.2716, 184.3507, 194.1424, 209.4889, 210.3278, 198.0795, 
    193.6121, 191.4348, 191.4185, 191.5776, 191.1826, 189.8961, 188.5744, 
    187.314,
  172.5305, 173.5165, 175.6244, 188.4975, 203.2316, 207.0844, 198.3879, 
    193.3186, 190.3197, 188.4564, 188.3522, 188.4422, 188.0485, 187.6564, 
    186.5033,
  177.8272, 176.2357, 173.399, 182.5946, 191.591, 197.7204, 197.2228, 
    195.2343, 189.5217, 184.0423, 184.581, 187.2677, 186.6772, 187.0748, 
    187.3168,
  181.3122, 172.8061, 175.4204, 193.2381, 198.2117, 190.4581, 187.8414, 
    187.625, 184.175, 182.7755, 177.264, 177.2463, 180.3289, 185.4226, 
    185.5235,
  186.893, 176.3516, 174.2383, 191.0622, 196.1385, 189.7611, 189.1045, 
    189.0291, 192.0206, 188.6164, 183.1695, 183.4663, 183.1958, 185.5764, 
    182.7498,
  193.2647, 180.7224, 175.801, 194.7932, 202.445, 188.1396, 189.2165, 
    190.6302, 192.5042, 193.0184, 193.6705, 194.1587, 195.3777, 195.4565, 
    192.5081,
  194.7833, 184.4443, 180.6074, 193.4084, 205.2182, 202.3185, 183.8918, 
    189.8564, 193.1226, 194.3613, 195.9238, 195.6189, 195.2376, 189.8194, 
    183.7461,
  201.882, 189.436, 183.7791, 192.3323, 203.3766, 202.8162, 203.0356, 
    182.4108, 187.7006, 192.4307, 190.4942, 187.1128, 184.0701, 178.5345, 
    170.2016,
  208.1871, 196.4398, 186.9081, 190.8345, 202.4723, 202.2345, 200.6079, 
    198.5957, 192.4594, 192.8505, 190.2271, 185.3691, 180.1289, 177.9322, 
    172.6982,
  213.1001, 200.9404, 191.037, 191.8199, 204.6129, 204.3296, 199.3151, 
    194.3181, 191.3724, 191.6362, 187.8837, 184.0284, 180.4398, 178.8521, 
    172.6735,
  218.4086, 208.4498, 193.8074, 192.4225, 201.4922, 204.8501, 199.4067, 
    194.6616, 190.365, 187.8261, 184.4878, 183.1358, 178.9841, 176.2617, 
    175.5963,
  220.8072, 215.9298, 199.4257, 190.3047, 200.6512, 204.1368, 199.1878, 
    194.3309, 189.7982, 186.0827, 183.9416, 180.2155, 179.814, 176.033, 
    175.1174,
  221.0298, 217.2798, 206.2156, 195.5849, 196.2638, 200.3458, 198.8198, 
    195.8584, 191.1759, 185.5907, 182.4509, 182.831, 180.9373, 176.128, 
    171.7421,
  197.0297, 197.0882, 196.4754, 196.4634, 194.2195, 191.8851, 192.4098, 
    187.0173, 188.7753, 182.5882, 181.9909, 184.0269, 180.5782, 182.2473, 
    176.8518,
  203.4268, 200.7888, 200.6891, 197.3743, 194.2031, 190.4745, 190.1341, 
    189.3991, 189.4162, 189.354, 187.6823, 192.2753, 191.8553, 180.007, 
    178.2256,
  207.3172, 203.0769, 202.243, 200.3921, 199.9882, 186.193, 186.2694, 
    181.1395, 180.5933, 187.536, 191.898, 193.7614, 192.6531, 191.1225, 
    186.1605,
  202.6124, 207.0887, 202.7695, 202.3216, 196.6862, 192.0591, 180.0917, 
    177.7865, 175.2661, 172.8724, 174.5628, 186.5307, 190.4008, 192.744, 
    191.2878,
  200.2502, 202.9844, 203.7359, 199.4717, 194.3445, 191.5145, 188.7687, 
    179.7079, 178.6518, 169.7533, 167.1225, 166.7607, 175.2126, 182.8703, 
    187.5894,
  204.8522, 203.2451, 205.1686, 201.06, 196.5261, 190.1428, 183.562, 
    180.9042, 175.1787, 166.0287, 165.0635, 166.9887, 168.3669, 176.6479, 
    183.7668,
  210.8932, 201.219, 198.6422, 199.5891, 205.577, 192.2598, 182.3307, 
    177.0838, 173.1962, 170.7138, 169.083, 168.8454, 167.1189, 172.1119, 
    176.9921,
  213.2895, 204.9826, 199.4793, 202.0855, 205.2218, 201.1027, 185.571, 
    178.8332, 173.4778, 169.353, 167.2961, 167.2771, 170.7706, 171.6818, 
    177.0555,
  217.6589, 200.3952, 200.8691, 203.2906, 201.9847, 199.1976, 191.696, 
    182.6423, 173.7606, 171.5393, 169.3698, 167.7574, 167.1947, 171.496, 
    171.618,
  206.4963, 201.2977, 206.0458, 201.6467, 199.023, 198.4476, 196.8924, 
    192.9734, 185.5861, 175.7395, 173.5044, 170.1239, 167.4517, 166.7139, 
    169.2438,
  201.4759, 200.1817, 195.9441, 196.1738, 193.3175, 187.3806, 187.5127, 
    183.9977, 183.4039, 181.0211, 181.167, 185.8054, 184.1031, 185.4805, 
    184.5573,
  203.8995, 200.5071, 197.4914, 196.5561, 193.5471, 186.4848, 184.6363, 
    184.5228, 183.0477, 184.0768, 182.1015, 187.7302, 186.4448, 180.5885, 
    180.7119,
  204.7708, 202.5616, 200.3803, 197.3582, 196.9138, 186.485, 184.4082, 
    182.3965, 180.1953, 183.0414, 186.9198, 189.202, 187.601, 183.432, 
    183.1387,
  200.6683, 198.922, 201.869, 196.9793, 194.7055, 197.5726, 180.9105, 182.9, 
    185.2673, 183.6947, 184.9027, 190.0698, 189.6139, 186.2251, 184.8252,
  198.938, 202.1162, 198.2733, 198.4146, 194.9988, 194.2046, 195.6296, 
    181.0363, 183.072, 183.9784, 185.2983, 189.7097, 190.6532, 189.1327, 
    187.0978,
  196.7562, 193.628, 195.1482, 195.252, 192.6156, 191.7914, 190.5706, 
    189.7821, 180.5298, 179.3225, 182.6644, 189.6722, 190.7981, 189.9488, 
    188.1071,
  195.1327, 193.5524, 193.3155, 193.7772, 191.8537, 195.0052, 191.3329, 
    187.0974, 180.95, 177.0147, 180.7363, 188.1722, 189.1324, 190.276, 
    188.6513,
  197.2421, 191.7166, 188.7575, 187.6915, 189.8987, 197.9525, 193.4707, 
    191.082, 184.7734, 176.4439, 172.8731, 177.669, 186.4629, 191.8916, 
    189.4043,
  199.0786, 192.2804, 196.6199, 192.3214, 198.7101, 192.5029, 194.1369, 
    192.9801, 186.6806, 176.2668, 172.0304, 169.8515, 174.4681, 184.3171, 
    190.4321,
  200.2659, 198.6425, 195.4038, 189.2566, 185.3941, 190.8121, 192.4108, 
    196.4297, 191.2801, 178.5928, 171.8651, 169.7597, 167.4496, 170.5181, 
    185.4452,
  199.0611, 199.4225, 197.4025, 196.287, 192.6373, 188.2792, 187.701, 
    189.0852, 189.637, 185.9214, 185.967, 186.5867, 183.3076, 182.0262, 
    181.025,
  202.4155, 199.56, 196.5945, 196.183, 193.8083, 185.5081, 185.4889, 
    187.6519, 188.9164, 188.9794, 185.9666, 188.0868, 189.8028, 182.2522, 
    182.3155,
  202.6139, 200.7874, 197.884, 198.2497, 196.3915, 184.9135, 186.6555, 
    186.6784, 185.0167, 186.8266, 187.883, 187.8035, 188.7741, 190.3358, 
    188.5039,
  203.4902, 202.0183, 201.5873, 198.6306, 199.7358, 198.3315, 183.0619, 
    186.133, 185.4182, 183.9733, 187.4046, 187.998, 187.9147, 188.2047, 
    189.0284,
  207.452, 207.8549, 198.8032, 196.9692, 197.5392, 197.4165, 196.9417, 
    174.4267, 177.2317, 177.9904, 184.3974, 187.3146, 186.3503, 185.8713, 
    186.9243,
  212.359, 209.0754, 196.7191, 200.6569, 196.1291, 192.7539, 188.2559, 
    186.5867, 178.7621, 176.7676, 182.0818, 187.0157, 184.5446, 181.9718, 
    182.88,
  212.1478, 203.5444, 193.4381, 200.6783, 204.4351, 193.9405, 184.4509, 
    180.6897, 173.226, 179.1631, 183.3579, 184.2804, 182.4115, 179.3764, 
    179.2827,
  205.8821, 203.9648, 192.343, 187.6089, 198.9204, 196.6113, 182.2183, 
    177.1127, 172.6557, 176.7033, 181.1505, 181.7618, 183.0107, 179.3501, 
    175.9847,
  206.4869, 190.9883, 190.9433, 215.4908, 204.6474, 191.377, 183.2605, 
    175.6276, 170.1499, 173.4521, 179.647, 181.3096, 178.9855, 178.099, 
    177.0284,
  199.8535, 203.0448, 214.0098, 196.6858, 188.7, 187.745, 184.7324, 179.9863, 
    170.5118, 170.0246, 176.555, 178.3419, 179.6209, 177.9077, 176.6414,
  193.2948, 192.7634, 192.4054, 190.7909, 190.8712, 186.8376, 185.4915, 
    183.5173, 183.675, 181.8976, 184.769, 186.2371, 185.0234, 182.8189, 
    183.0036,
  196.8354, 195.2075, 195.8649, 193.7381, 191.2082, 181.7831, 183.3434, 
    185.2311, 186.2246, 188.952, 187.9117, 189.3583, 188.6323, 185.5763, 
    181.9354,
  209.6112, 197.2912, 195.5608, 197.7439, 196.9061, 180.6879, 183.3094, 
    183.3342, 183.961, 186.861, 190.2815, 190.3096, 188.9301, 187.8184, 
    184.1956,
  221.1894, 214.9953, 209.1069, 196.7916, 197.946, 195.4755, 175.8115, 
    183.6236, 184.9138, 186.8899, 189.506, 189.991, 189.2881, 188.2778, 
    186.6003,
  220.586, 213.2316, 210.7904, 198.0043, 196.3436, 196.7437, 191.9709, 
    170.1113, 173.9652, 173.9815, 180.9515, 185.0806, 186.4129, 189.0219, 
    189.2828,
  222.5867, 208.0061, 214.6861, 204.3337, 199.5179, 193.2449, 182.6477, 
    177.7981, 175.5038, 175.0305, 176.8729, 181.6836, 183.8709, 187.3294, 
    188.6869,
  221.401, 219.9608, 216.8485, 206.6669, 208.0113, 194.1023, 181.7194, 
    176.5427, 172.8514, 177.8433, 180.6012, 180.7043, 182.446, 184.7743, 
    186.7316,
  214.3021, 213.4672, 207.311, 200.2789, 202.4896, 194.2708, 184.7812, 
    180.4762, 177.1483, 179.5835, 182.6301, 182.6967, 182.7803, 184.4209, 
    184.9277,
  216.1685, 199.5396, 199.6585, 206.4742, 194.4012, 186.3305, 184.5944, 
    181.8437, 180.7426, 181.3744, 182.0167, 183.2885, 182.8111, 183.6137, 
    181.6826,
  201.3629, 196.8153, 200.6962, 186.4743, 181.2384, 179.3517, 178.5927, 
    189.9055, 185.1394, 178.1663, 177.4303, 181.3289, 181.7429, 180.9881, 
    179.038,
  192.879, 194.0937, 192.9948, 192.9334, 189.6584, 184.6402, 185.813, 
    186.641, 186.0597, 181.1461, 181.7133, 180.2811, 175.776, 174.5251, 
    172.0895,
  199.289, 197.4346, 196.361, 195.3602, 191.7786, 185.9512, 187.6653, 
    188.3156, 189.7696, 188.0287, 186.4957, 184.9578, 180.7032, 173.1723, 
    170.6459,
  212.4552, 199.5335, 197.6473, 199.2762, 198.6094, 186.8921, 187.6262, 
    186.0432, 186.174, 187.6471, 190.0497, 191.2819, 187.568, 184.2184, 
    179.2484,
  222.8221, 218.8947, 209.5273, 199.1495, 202.2784, 198.0194, 187.8325, 
    190.0295, 186.8657, 186.2764, 189.2319, 191.4931, 191.0041, 190.6934, 
    185.5299,
  223.361, 216.3871, 210.2399, 195.9017, 192.7051, 190.106, 185.0868, 
    176.9468, 179.8392, 181.7688, 182.0802, 187.574, 187.219, 188.8313, 
    188.953,
  216.3437, 205.4845, 201.9131, 192.4739, 184.0405, 179.2755, 171.3549, 
    171.6667, 173.1012, 173.9308, 176.3836, 176.1603, 178.063, 180.9705, 
    184.7526,
  207.2042, 193.0873, 193.0872, 183.6573, 178.8036, 166.9513, 166.9028, 
    164.0345, 168.0555, 171.8047, 173.2953, 173.2836, 173.9452, 175.5051, 
    178.7475,
  195.0806, 183.1454, 180.683, 174.577, 163.3183, 163, 165.399, 167.0688, 
    168.8226, 172.6209, 170.7822, 172.1627, 173.5109, 176.0944, 178.5801,
  187.9074, 176.8064, 174.8991, 165.569, 157.6248, 163.1845, 167.5657, 
    166.7779, 173.0708, 173.8404, 171.5603, 171.0433, 169.3999, 173.1908, 
    176.0987,
  187.9552, 175.3199, 166.391, 160.5803, 160.8388, 168.6614, 172.7126, 
    178.2058, 176.2504, 169.7468, 167.2177, 166.836, 168.4869, 170.3521, 
    176.1474,
  203.4455, 197.5849, 192.9584, 193.5665, 189.4288, 185.9384, 187.0372, 
    183.6749, 183.631, 182.8144, 184.7827, 186.9264, 183.549, 185.0564, 
    182.0269,
  206.648, 204.8944, 203.4356, 202.9545, 199.61, 199.9445, 200.0645, 
    198.4658, 196.2363, 195.2196, 194.1623, 194.0348, 193.5177, 189.5557, 
    187.7598,
  217.0681, 207.5434, 203.1175, 199.9576, 205.9986, 203.3546, 202.3241, 
    193.872, 192.9202, 193.0999, 192.4213, 192.0178, 191.3522, 190.071, 
    188.8286,
  223.676, 203.6582, 189.0004, 186.2558, 192.787, 203.757, 196.8429, 
    193.9371, 185.1943, 180.9124, 182.9126, 185.4368, 183.5237, 183.1749, 
    183.6492,
  208.4018, 179.9112, 171.2866, 175.8804, 177.2888, 182.4454, 189.4646, 
    186.6656, 185.8121, 184.3467, 184.5131, 184.1693, 180.5591, 181.001, 
    179.9336,
  183.0184, 169.1715, 173.4755, 173.3092, 179.8583, 180.4233, 178.3434, 
    180.6593, 184.3298, 184.8082, 187.5794, 188.2508, 184.8733, 183.6202, 
    179.8014,
  170.274, 171.7675, 175.7733, 170.6997, 177.0344, 181.2912, 185.6857, 
    187.7958, 187.5947, 185.3861, 184.7367, 185.5756, 186.4284, 184.7189, 
    181.5467,
  173.6319, 176.1769, 177.1855, 175.9179, 182.8811, 186.0348, 189.2124, 
    187.3512, 185.5414, 183.9594, 183.4015, 183.2119, 183.8963, 184.6433, 
    182.2189,
  177.7234, 175.4656, 177.1894, 181.647, 181.8687, 187.4649, 188.056, 
    187.192, 187.1673, 186.7398, 183.1809, 181.1837, 181.2084, 180.6428, 
    179.245,
  178.9196, 178.324, 180.9008, 180.6722, 184.2582, 187.9392, 185.4897, 
    191.869, 189.8582, 182.1712, 181.8752, 179.8845, 177.0288, 177.6187, 
    176.0389,
  203.698, 204.7941, 204.752, 203.2768, 206.3322, 206.9298, 207.7653, 
    204.0455, 201.6803, 195.7861, 195.3962, 193.8073, 188.1258, 186.4405, 
    177.3138,
  203.4373, 205.192, 204.5062, 203.2435, 205.7351, 201.7262, 205.4418, 
    201.8218, 200.7231, 198.5527, 196.4328, 196.3096, 196.5216, 194.3336, 
    193.431,
  218.5046, 210.4923, 205.9746, 204.2568, 206.6875, 202.0924, 204.0591, 
    198.25, 197.4817, 195.1077, 194.2413, 194.9966, 195.0462, 194.0471, 
    192.7638,
  227.6316, 220.5382, 202.3081, 193.9413, 193.3715, 200.5331, 192.475, 
    195.8553, 192.2943, 188.7582, 190.9691, 192.7808, 192.1539, 191.5059, 
    191.9608,
  220.9264, 202.1477, 186.1066, 184.0643, 183.4674, 191.7728, 197.6772, 
    186.1227, 186.8082, 190.0055, 190.7211, 190.3591, 189.3017, 190.0123, 
    189.8422,
  204.0083, 186.8368, 181.3364, 181.3769, 188.9064, 192.007, 193.4688, 
    189.7762, 187.376, 183.7859, 186.2677, 188.3793, 188.3247, 188.5132, 
    187.8925,
  179.8406, 178.8681, 181.5255, 188.7315, 201.4154, 194.9526, 188.5332, 
    185.9574, 184.3379, 182.9764, 182.681, 183.332, 183.9682, 184.1818, 
    184.7243,
  178.0218, 182.391, 189.9794, 200.5109, 207.6874, 194.062, 187.4719, 
    185.5172, 184.6647, 183.5055, 182.519, 182.5199, 182.3783, 182.0706, 
    182.6985,
  180.7932, 177.6302, 193.5374, 209.7236, 198.4612, 190.4696, 187.313, 
    187.254, 187.6267, 187.8567, 182.6129, 180.6252, 182.4954, 183.6318, 
    182.2022,
  174.6005, 189.5168, 197.4576, 195.4514, 190.3929, 188.4501, 186.9479, 
    192.3763, 191.6478, 182.5442, 182.0813, 180.523, 181.57, 183.5173, 
    180.1484,
  165.8037, 166.9411, 172.921, 184.2728, 192.664, 197.0789, 203.9912, 
    202.3659, 198.9507, 194.142, 193.5679, 191.6068, 189.2819, 189.4507, 
    187.5408,
  164.7304, 166.2028, 174.0295, 181.1014, 189.4603, 193.2471, 196.6232, 
    197.481, 193.2639, 190.6624, 188.2358, 189.0836, 189.5046, 187.2245, 
    187.7218,
  167.5193, 169.6432, 176.576, 186.6681, 190.7526, 194.0839, 192.1912, 
    185.8013, 188.6205, 189.7124, 189.2587, 188.6663, 188.381, 187.8029, 
    187.3188,
  178.6872, 184.299, 181.2594, 185.6818, 186.1418, 193.5122, 188.2378, 
    187.9797, 188.1214, 188.0338, 189.615, 188.6808, 187.303, 186.3755, 
    185.4943,
  183.3752, 187.004, 185.2288, 187.5147, 183.1965, 185.1993, 194.6394, 
    186.5739, 182.7247, 189.1091, 191.2632, 188.0388, 185.9443, 185.4091, 
    184.9043,
  197.0555, 191.1945, 184.7901, 187.6426, 187.9609, 193.3773, 194.0258, 
    191.4704, 186.824, 182.5341, 182.657, 185.1642, 185.0478, 184.6479, 
    183.6626,
  199.4241, 191.8275, 186.3942, 188.2659, 195.5728, 195.9071, 191.7956, 
    187.5401, 185.3858, 184.2403, 184.9552, 184.5701, 184.4661, 183.3748, 
    182.6577,
  187.2778, 181.7834, 192.2384, 195.9761, 203.1218, 193.6956, 189.1349, 
    186.5941, 187.1024, 186.1955, 185.3904, 183.8513, 182.2661, 181.1439, 
    182.0542,
  173.9458, 177.8582, 185.6353, 198.838, 195.1174, 190.134, 187.631, 
    188.6525, 190.2169, 189.4721, 183.1472, 180.1629, 180.1477, 180.8486, 
    179.4622,
  172.8392, 170.4421, 183.7975, 186.4865, 184.4824, 185.8975, 186.0195, 
    192.2196, 193.24, 182.9839, 180.2023, 176.2758, 176.527, 176.636, 174.2554,
  175.9724, 170.1823, 169.0076, 172.0991, 172.5313, 177.8594, 172.755, 
    176.9474, 181.1617, 182.3493, 182.3746, 187.3828, 186.8717, 185.4085, 
    186.4053,
  170.935, 175.1809, 171.5361, 174.6407, 169.4853, 171.1913, 172.5718, 
    174.3307, 176.6905, 178.5474, 181.2594, 184.1145, 182.533, 185.2641, 
    183.9534,
  172.2829, 170.6905, 176.0199, 171.0109, 173.5424, 171.7806, 169.7609, 
    166.1398, 173.3748, 179.324, 178.5391, 180.6191, 180.0367, 180.9823, 
    184.8625,
  178.4072, 173.7473, 173.1023, 177.9476, 170.7591, 171.1565, 169.3613, 
    171.5146, 172.7391, 177.1159, 177.903, 180.8407, 179.1794, 177.7621, 
    180.4059,
  188.6908, 179.7524, 170.0943, 166.9552, 167.8453, 167.9778, 167.7243, 
    170.2038, 174.8921, 172.3541, 175.1221, 179.6303, 180.4308, 177.9227, 
    179.1429,
  203.6853, 187.6783, 177.6452, 166.02, 168.9252, 171.3779, 172.0182, 
    171.3037, 176.3115, 176.9317, 177.3873, 179.0479, 177.6431, 179.4252, 
    179.272,
  206.6603, 202.5974, 187.1301, 176.4722, 171.3234, 168.0705, 168.117, 
    166.9624, 171.0743, 173.3039, 173.2609, 174.7323, 178.2703, 182.5717, 
    181.2728,
  194.3049, 193.6693, 190.8722, 176.3098, 169.5545, 170.7807, 172.5495, 
    172.2711, 172.5486, 175.4115, 177.7385, 180.4432, 182.7721, 181.438, 
    179.7469,
  195.3456, 190.9581, 181.1118, 181.37, 175.5643, 176.3934, 172.2247, 
    172.7838, 178.1026, 182.2856, 182.4391, 182.4893, 180.5638, 178.9189, 
    175.2539,
  179.2244, 175.1221, 171.8582, 175.7705, 173.2271, 177.939, 178.6609, 
    183.9888, 187.2278, 182.9587, 178.052, 177.2991, 176.3703, 173.7308, 
    169.6646,
  195.0473, 193.8904, 192.1766, 195.2281, 197.0502, 201.212, 203.3583, 
    204.8846, 201.4613, 191.9978, 184.7503, 182.6694, 178.1173, 174.2206, 
    173.7825,
  197.6055, 194.53, 188.3891, 188.2334, 186.9963, 194.246, 195.8322, 
    196.5314, 197.2489, 190.3758, 186.8757, 181.9993, 180.8324, 177.702, 
    174.7088,
  203.899, 195.601, 188.1731, 177.2586, 180.033, 180.5697, 188.3338, 
    189.6632, 190.5788, 189.5828, 188.7641, 183.0281, 175.9838, 178.8563, 
    175.1958,
  204.931, 202.1861, 172.4725, 169.0663, 170.0751, 170.3818, 171.7466, 
    181.5319, 185.3092, 188.1175, 186.0085, 181.4956, 176.9446, 178.6691, 
    170.5425,
  205.7077, 210.0772, 175.1592, 164.5215, 165.8003, 169.2233, 172.9726, 
    180.127, 184.6207, 180.6509, 182.3663, 179.3003, 177.9847, 180.2404, 
    173.3096,
  202.1619, 198.7329, 177.0881, 165.7779, 167.589, 166.1295, 170.5104, 
    173.75, 174.0217, 174.2319, 177.6499, 176.285, 181.1286, 176.2346, 
    175.4601,
  196.8982, 205.5072, 183.2338, 161.1537, 165.2906, 164.9489, 171.1175, 
    173.1415, 175.664, 178.4346, 177.3499, 179.1379, 180.8688, 178.4733, 
    177.9778,
  185.8076, 192.8932, 185.6583, 173.1818, 164.8153, 167.8316, 173.1913, 
    174.9047, 181.3646, 180.6768, 181.1641, 180.7062, 181.7431, 180.1363, 
    178.8606,
  182.7444, 180.8779, 181.2178, 174.9573, 167.2835, 167.732, 170.8304, 
    174.3061, 179.7703, 181.7611, 184.0684, 183.6026, 183.0338, 181.2152, 
    178.9916,
  195.2567, 189.8289, 187.3477, 179.4894, 178.1899, 180.4626, 185.5876, 
    192.9387, 191.5158, 183.0182, 177.9607, 177.6675, 176.4342, 176.405, 
    176.7906,
  211.1582, 201.2314, 192.21, 190.9015, 190.7246, 195.9061, 197.4973, 
    196.9973, 198.211, 195.2218, 191.8974, 188.8972, 181.4788, 180.6371, 
    173.5666,
  198.0408, 191.1052, 190.4038, 193.3737, 193.0758, 192.2793, 192.0026, 
    193.9542, 198.0124, 198.1255, 192.3994, 187.5974, 182.4949, 176.4474, 
    173.2506,
  191.7298, 188.0948, 187.7289, 187.2083, 186.9821, 187.0859, 189.2558, 
    190.1509, 196.141, 199.2657, 197.7272, 188.8804, 184.8727, 177.7821, 
    174.9608,
  192.8403, 189.1593, 188.0968, 182.1205, 181.8763, 186.9468, 184.3866, 
    187.8653, 194.5699, 198.6384, 200.0407, 194.8546, 186.449, 173.0294, 
    169.8802,
  192.7774, 190.848, 191.0492, 183.7603, 182.1624, 181.5578, 184.0132, 
    183.2904, 187.4171, 192.2341, 197.8826, 200.081, 190.4089, 182.2698, 
    170.0603,
  195.0422, 193.0343, 190.6078, 184.5845, 184.4958, 181.9583, 182.3214, 
    178.4117, 174.267, 176.6995, 187.4745, 190.5031, 189.2083, 184.1991, 
    174.0286,
  205.9436, 199.1663, 196.2679, 189.6174, 192.937, 188.2265, 186.0726, 
    181.3143, 176.6483, 174.5353, 173.8455, 179.2177, 182.9965, 181.4037, 
    175.9942,
  201.4093, 203.7824, 195.9498, 198.0084, 197.8262, 188.6454, 188.149, 
    187.7664, 181.6098, 179.3689, 175.9437, 174.156, 175.9268, 176.9624, 
    177.2788,
  202.0795, 196.5435, 196.9605, 208.9071, 196.7721, 191.6227, 191.5574, 
    190.5792, 187.6101, 184.4386, 181.3407, 182.9269, 182.976, 181.9198, 
    180.9646,
  190.207, 194.8529, 202.2791, 195.3906, 191.4731, 189.7639, 189.9741, 
    194.6783, 188.0473, 180.4166, 178.407, 179.7249, 179.5831, 179.8807, 
    179.3984,
  213.2501, 209.2171, 207.3422, 204.8987, 201.1767, 199.6264, 201.6566, 
    201.6128, 198.4798, 196.039, 196.3783, 194.7146, 192.0163, 191.0388, 
    191.632,
  212.4831, 209.8946, 206.8614, 205.2307, 200.3608, 201.0571, 200.091, 
    201.6436, 200.8164, 197.2898, 196.2481, 193.3149, 189.8572, 188.8, 
    190.9027,
  220.4382, 213.8515, 208.3307, 203.4736, 201.0902, 195.8116, 200.8262, 
    198.6904, 196.861, 194.3918, 192.2133, 187.423, 189.311, 190.1357, 
    191.2712,
  215.7072, 216.0476, 210.8148, 199.8289, 196.4942, 198.5416, 190.1566, 
    194.1673, 187.1902, 186.3387, 189.4488, 190.3893, 188.9978, 191.9963, 
    191.295,
  204.0372, 198.5404, 196.0299, 190.2188, 193.0098, 194.7516, 196.4725, 
    181.9566, 181.3638, 186.5569, 185.9071, 188.9048, 190.6958, 191.6147, 
    192.4659,
  189.6338, 182.453, 184.1494, 185.0027, 187.6817, 192.8857, 191.0249, 
    186.7435, 182.6324, 181.2301, 182.4555, 185.2003, 185.3336, 185.1837, 
    182.3287,
  174.3138, 172.8847, 174.3706, 180.3568, 191.3509, 191.3983, 188.4997, 
    179.2331, 176.9433, 176.9189, 178.8563, 178.4296, 179.5502, 180.5643, 
    177.008,
  167.7712, 168.0853, 167.0448, 180.0647, 197.9975, 190.9579, 187.7836, 
    182.5043, 178.7821, 175.712, 176.0041, 179.3674, 179.3137, 177.8877, 
    176.733,
  171.9935, 167.8152, 169.0724, 189.3402, 197.3664, 190.4265, 186.2913, 
    181.5532, 177.9054, 174.27, 175.7898, 178.6743, 180.1462, 180.1505, 
    178.7406,
  178.0375, 180.1216, 182.7555, 187.6555, 192.6759, 188.1304, 185.5641, 
    185.3185, 179.1481, 173.5217, 173.4362, 176.764, 178.4381, 179.685, 
    180.6543,
  199.0387, 193.6236, 187.2969, 188.8604, 183.2292, 185.7798, 187.3188, 
    186.5186, 186.0714, 187.3301, 189.0245, 189.2046, 190.3439, 191.1498, 
    188.9473,
  203.1738, 204.786, 201.801, 196.7251, 193.7576, 196.8145, 196.7695, 
    196.9174, 193.2587, 187.7165, 191.8048, 192.2285, 189.329, 187.0855, 
    184.8053,
  206.5806, 203.6965, 205.1178, 202.3385, 198.8382, 198.6575, 198.1588, 
    194.3238, 188.3757, 193.2907, 192.3797, 188.1315, 184.0288, 181.297, 
    180.5675,
  189.3358, 190.7166, 199.4414, 199.6082, 193.7332, 195.5061, 191.271, 
    187.7237, 181.4388, 177.9048, 182.224, 183.6301, 182.8295, 180.8739, 
    180.5563,
  181.7194, 186.1921, 183.5311, 186.195, 185.1217, 184.1566, 180.3755, 
    174.9898, 176.4294, 178.8802, 178.8124, 180.978, 180.6255, 181.9902, 
    181.5706,
  188.8921, 186.7325, 184.5991, 188.3756, 184.19, 180.6051, 178.6224, 
    179.8964, 177.0512, 176.3884, 176.4528, 179.3245, 178.4441, 179.8074, 
    180.2309,
  195.1518, 191.1468, 195.3132, 192.5768, 190.4631, 186.0378, 183.324, 
    182.418, 181.4535, 180.8266, 179.5871, 177.0391, 177.9108, 178.2299, 
    179.0569,
  209.7012, 205.5916, 207.4209, 211.0058, 202.3643, 192.0643, 188.1506, 
    184.7942, 182.9542, 179.8536, 177.5604, 176.5299, 174.3839, 175.8665, 
    179.634,
  219.2544, 216.2653, 216.8841, 218.4255, 197.5431, 190.3763, 186.3409, 
    184.1428, 181.094, 178.059, 173.5414, 172.3276, 171.6897, 172.5961, 
    176.4926,
  219.2993, 215.562, 214.0694, 195.5348, 188.4339, 186.0586, 183.8237, 
    183.9874, 179.2988, 169.9298, 165.9466, 165.1299, 167.7944, 171.2398, 
    174.7382,
  178.2182, 166.8297, 160.7027, 153.4674, 155.4322, 163.9291, 160.2536, 
    158.9073, 166.2605, 160.9301, 167.7852, 165.0563, 161.882, 161.5674, 
    162.9144,
  180.5569, 171.5549, 163.803, 154.5045, 155.2379, 156.2884, 159.9213, 
    156.7358, 162.505, 161.7787, 163.2202, 159.3796, 166.1694, 163.5486, 
    164.3645,
  199.4822, 184.5964, 172.292, 164.352, 160.7784, 161.4958, 161.4015, 
    161.4873, 165.908, 171.6105, 170.5737, 172.1636, 175.1994, 176.7654, 
    174.5726,
  212.6278, 208.4844, 191.7402, 181.4222, 174.3748, 173.6277, 170.3663, 
    173.4536, 175.6678, 174.8177, 181.8926, 179.2737, 183.4687, 182.8028, 
    182.9862,
  224.0311, 218.3398, 211.1674, 197.2795, 190.4216, 183.5983, 179.8698, 
    177.3942, 175.7668, 174.2644, 176.401, 177.8056, 178.73, 179.8649, 
    182.8785,
  215.3927, 214.7924, 210.6829, 203.9511, 199.3966, 191.459, 189.2414, 
    186.4735, 183.0037, 176.0839, 174.5914, 179.0778, 178.8637, 181.4592, 
    180.5697,
  218.5253, 217.3448, 220.3326, 211.6675, 206.1669, 196.804, 191.7075, 
    186.4072, 181.2953, 179.4017, 180.9735, 179.2766, 181.4333, 182.9627, 
    180.7952,
  216.6057, 209.3589, 209.6937, 222.6092, 213.247, 194.9563, 189.6891, 
    185.6875, 186.4211, 185.4215, 184.958, 184.1588, 182.851, 178.7808, 
    177.597,
  208.4901, 209.4663, 216.1952, 213.335, 202.6828, 196.3709, 193.6952, 
    192.3205, 191.3439, 189.5575, 185.9758, 183.6506, 181.0845, 178.0495, 
    177.1297,
  199.6364, 202.9423, 206.0319, 201.9546, 198.4615, 196.686, 194.6076, 
    195.6183, 194.6519, 193.1623, 191.2477, 185.9193, 184.4211, 179.6944, 
    177.2936,
  194.1591, 181.1367, 172.0923, 171.2469, 176.552, 181.076, 190.97, 197.5056, 
    199.8702, 202.6452, 209.2944, 210.9494, 213.7527, 213.4485, 210.293,
  202.6046, 185.9823, 173.2072, 164.1327, 172.0783, 178.7055, 189.2227, 
    195.5649, 201.2464, 203.4709, 208.127, 208.8851, 211.5907, 208.1851, 
    199.5859,
  215.7741, 201.5038, 177.4872, 166.6345, 166.3657, 177.482, 188.2132, 
    189.1484, 193.8727, 196.5973, 202.4505, 205.4812, 201.9792, 201.2437, 
    197.7358,
  214.0339, 222.7983, 192.7218, 169.0288, 165.5599, 170.4888, 180.7157, 
    187.5244, 190.2094, 191.2971, 196.5643, 199.4426, 198.7287, 193.9961, 
    191.5769,
  212.9358, 224.3389, 224.3921, 179.2794, 169.2904, 162.7445, 173.8094, 
    182.0568, 183.7382, 188.3349, 188.0842, 190.6845, 191.5944, 190.3799, 
    185.0768,
  222.8227, 228.6058, 228.2855, 197.2769, 171.8252, 165.8776, 164.6752, 
    168.4758, 175.9382, 176.6911, 181.5204, 184.7754, 181.6889, 176.8545, 
    171.6719,
  225.7822, 229.8679, 229.37, 210.2406, 188.5528, 172.3337, 165.6993, 
    163.673, 163.594, 168.105, 169.7374, 171.7867, 169.9828, 168.8968, 
    169.2812,
  231.55, 224.1433, 228.3086, 225.289, 211.9072, 182.879, 170.4435, 165.898, 
    168.2, 164.9935, 164.2826, 166.2699, 164.8733, 164.6624, 166.7689,
  199.6974, 200.5402, 210.5565, 216.504, 208.8414, 199.7448, 184.1326, 
    174.1857, 170.9055, 166.1182, 165.9052, 162.68, 164.232, 166.9447, 
    168.8839,
  174.8295, 180.1929, 186.8212, 196.5608, 201.8821, 203.8685, 197.4621, 
    189.3109, 183.1442, 176.8697, 172.9537, 171.3421, 173.1797, 170.6044, 
    174.7805,
  213.3943, 211.0188, 209.8106, 205.2542, 199.4637, 196.1244, 200.7488, 
    200.5236, 205.5908, 209.164, 206.2279, 208.6277, 208.9902, 208.087, 
    205.3328,
  211.3348, 212.9407, 212.2777, 201.3883, 199.6506, 195.8494, 197.2435, 
    199.3678, 206.3926, 205.3555, 206.4072, 208.8449, 210.2839, 204.9085, 
    200.4804,
  207.816, 214.2308, 214.1386, 196.0677, 193.6502, 196.9324, 196.4996, 
    198.7192, 195.8265, 198.4888, 206.9731, 206.5296, 201.096, 197.5857, 
    202.907,
  201.4476, 209.6789, 210.1581, 198.3493, 189.64, 200.0914, 201.4257, 
    199.0836, 204.6582, 199.3187, 202.41, 199.5095, 199.1516, 203.2815, 
    200.6543,
  197.4025, 210.9788, 219.9155, 201.7307, 188.0165, 188.7502, 197.9314, 
    199.4219, 199.4178, 199.8132, 198.3626, 197.0723, 198.3462, 200.0072, 
    193.5888,
  205.236, 206.3557, 216.4872, 208.7458, 186.1536, 185.3303, 200.2878, 
    209.1946, 212.3397, 205.2155, 197.3193, 193.4359, 194.7285, 195.0403, 
    194.5187,
  207.4823, 203.1948, 212.0434, 212.313, 194.3793, 178.4417, 199.9605, 
    205.3541, 209.1207, 200.5322, 194.6513, 191.1769, 189.3453, 190.7569, 
    198.1822,
  199.7153, 200.5174, 204.9835, 216.6579, 210.4037, 180.7445, 186.6101, 
    205.9223, 207.3468, 198.8806, 191.2061, 189.2209, 190.6059, 188.9207, 
    191.0266,
  208.7983, 204.5156, 198.4743, 203.494, 208.0443, 185.3911, 181.9422, 
    196.1265, 199.9092, 194.1629, 187.8185, 188.605, 189.4031, 184.6687, 
    182.8044,
  219.1218, 212.632, 197.1897, 193.1008, 196.8854, 194.7796, 182.118, 
    189.0598, 194.4812, 194.6082, 185.5191, 185.2569, 183.6892, 180.1673, 
    181.5941,
  208.0718, 204.7877, 204.566, 204.7116, 208.1326, 208.3996, 211.7725, 
    209.8576, 209.6265, 206.0723, 207.0475, 209.7203, 207.9582, 206.7722, 
    204.9932,
  209.619, 205.6825, 201.7329, 202.693, 205.8292, 205.6016, 208.8195, 
    209.0456, 210.2549, 210.0824, 211.1898, 213.0058, 211.6291, 208.5515, 
    208.0545,
  217.0508, 209.9206, 206.1893, 200.9323, 200.8872, 203.2345, 206.0262, 
    206.8214, 202.9014, 204.3939, 202.6637, 202.7618, 206.4901, 212.252, 
    211.4451,
  224.3672, 217.2793, 208.4423, 200.3952, 201.7179, 205.6062, 206.1904, 
    207.2212, 210.8163, 200.0648, 208.2181, 208.0514, 209.3984, 207.3916, 
    207.3069,
  227.8171, 223.2836, 209.2769, 201.2048, 200.6972, 203.1085, 208.5849, 
    203.4252, 201.1201, 205.0045, 204.3685, 204.193, 204.4774, 203.9477, 
    199.6736,
  223.7507, 224.9317, 215.4871, 202.7008, 199.3673, 204.8596, 206.9597, 
    208.5152, 204.7622, 206.267, 207.129, 204.944, 203.2952, 200.8884, 
    197.5327,
  231.1694, 228.6056, 211.6748, 205.5956, 201.4745, 202.3161, 206.261, 
    205.6197, 204.3797, 208.3152, 206.6046, 204.35, 201.4628, 197.5344, 
    199.1696,
  228.0051, 228.6351, 210.4856, 206.2624, 197.1462, 203.1544, 206.3222, 
    209.7564, 203.9024, 205.3805, 204.2566, 197.9907, 196.9738, 197.8127, 
    196.8216,
  226.6243, 225.1416, 207.4115, 201.0277, 198.3049, 200.2801, 203.538, 
    204.6427, 202.0021, 201.5407, 194.0531, 192.0628, 196.921, 196.0727, 
    194.7483,
  216.1275, 211.541, 209.4997, 202.1971, 195.3384, 196.6133, 201.7483, 
    203.2782, 197.5041, 194.5968, 187.0965, 189.8234, 194.9762, 194.237, 
    194.5707,
  212.7554, 209.0363, 206.345, 207.4999, 201.0371, 189.9817, 195.7953, 
    200.3869, 198.304, 196.6361, 193.1138, 190.9524, 188.1336, 188.8806, 
    188.85,
  214.1119, 210.6345, 208.0863, 208.3615, 201.6016, 189.4483, 195.7154, 
    201.4955, 204.9862, 205.9053, 201.8902, 198.7772, 188.3844, 186.1884, 
    186.0048,
  221.3354, 219.1853, 212.0005, 208.3478, 205.2083, 193.5032, 198.4981, 
    203.8123, 204.369, 205.1214, 203.1876, 197.5854, 195.2955, 191.4626, 
    191.3875,
  220.2373, 224.3329, 221.1955, 212.6879, 206.8779, 202.8046, 199.9542, 
    203.3572, 208.5649, 204.6279, 205.3135, 203.4949, 200.0305, 198.4209, 
    194.7919,
  228.5087, 224.9749, 217.0715, 210.2816, 209.6624, 206.8966, 204.6468, 
    200.539, 196.7863, 202.5739, 203.8413, 202.3376, 199.584, 198.0157, 
    196.784,
  226.2711, 225.8771, 220.3606, 207.7498, 206.7045, 208.2719, 207.0613, 
    207.0934, 203.4849, 199.7535, 198.9431, 195.0328, 191.9884, 191.4076, 
    195.1285,
  217.5674, 216.8417, 210.7618, 205.361, 205.6926, 206.7772, 206.3204, 
    206.0931, 203.9896, 201.6948, 194.6477, 189.2499, 190.877, 194.6115, 
    195.5564,
  211.8767, 209.4527, 205.4894, 205.9373, 204.5796, 208.1367, 205.0865, 
    207.7794, 205.9657, 200.2176, 198.1266, 198.1746, 196.1672, 195.9578, 
    194.8609,
  214.0403, 210.9443, 206.8999, 208.0107, 210.6353, 206.8158, 205.063, 
    205.4282, 200.7779, 199.8127, 199.8721, 199.1441, 195.9562, 194.7191, 
    194.3744,
  228.8564, 222.3906, 212.4321, 206.0623, 207.434, 208.177, 206.4892, 
    206.9784, 199.6552, 199.5403, 198.7971, 196.2323, 194.5379, 193.8303, 
    194.848,
  215.5471, 209.1499, 208.8112, 208.716, 209.4644, 203.847, 202.9343, 
    200.0628, 199.9035, 197.5098, 187.1325, 189.9441, 185.3422, 185.5056, 
    190.1249,
  216.3416, 212.653, 210.5705, 210.3302, 210.916, 203.7504, 201.937, 
    201.4099, 203.2399, 199.3893, 194.0335, 194.8913, 189.7563, 187.4277, 
    185.4675,
  216.7312, 218.0803, 211.0146, 208.5181, 210.7986, 202.9909, 201.1182, 
    199.3856, 198.2915, 197.9816, 199.6577, 199.0695, 194.0194, 190.7962, 
    186.0697,
  218.2061, 220.204, 211.6117, 207.5296, 210.941, 209.7895, 198.0226, 
    196.1036, 198.0318, 197.2924, 197.3533, 198.9275, 200.1714, 196.9312, 
    190.1135,
  221.62, 211.0335, 211.4201, 208.8135, 209.6074, 209.6652, 210.1613, 
    196.1643, 193.8476, 194.565, 194.0393, 196.4375, 199.7336, 201.6197, 
    202.4667,
  221.4311, 216.1398, 210.6107, 204.3162, 208.0443, 209.2128, 207.6523, 
    208.7579, 199.1653, 193.0665, 188.9138, 191.6176, 196.2669, 198.7704, 
    201.7332,
  218.0732, 212.062, 208.6717, 202.1997, 203.511, 203.6211, 203.9602, 
    202.2152, 198.4588, 195.3171, 192.1894, 191.6119, 194.2548, 195.3038, 
    197.1856,
  221.1987, 215.5108, 203.4625, 198.0841, 197.4235, 199.6421, 198.4493, 
    197.5248, 195.7643, 193.7066, 191.3095, 191.6795, 194.2629, 194.8562, 
    194.6285,
  225.3464, 213.949, 198.8759, 192.9439, 189.8621, 193.7694, 195.528, 
    193.7759, 192.0289, 189.4976, 189.8908, 191.951, 192.3676, 193.2744, 
    194.0403,
  223.6054, 211.1112, 192.9374, 181.4897, 183.2927, 187.1367, 189.5041, 
    190.2737, 188.5473, 186.015, 187.2753, 188.2077, 189.6561, 190.7012, 
    193.9523,
  212.2133, 205.2256, 192.7721, 187.8679, 186.8231, 180.5524, 184.3181, 
    184.1715, 190.3115, 191.7207, 195.059, 196.9108, 193.5824, 190.1254, 
    185.3641,
  211.533, 200.1018, 190.0509, 186.1538, 182.4719, 178.5062, 176.1806, 
    181.5015, 183.2261, 190.9818, 193.7166, 196.6217, 199.8784, 194.141, 
    185.2676,
  214.5797, 200.7091, 186.47, 182.3882, 176.5902, 173.7014, 178.0034, 
    176.1788, 179.1993, 187.003, 191.3743, 195.7583, 201.0661, 205.3885, 
    196.4309,
  209.1545, 199.7101, 185.8767, 178.1866, 176.2668, 175.4481, 173.8166, 
    183.5345, 185.1948, 185.921, 189.7041, 191.4144, 196.9365, 201.7066, 
    204.629,
  208.2821, 198.4249, 185.515, 173.5555, 173.5856, 170.5376, 179.9713, 
    180.1263, 186.7032, 191.8896, 188.6237, 189.9659, 192.6326, 197.8952, 
    205.1207,
  200.5361, 188.6194, 182.4129, 175.7142, 174.1931, 174.4957, 182.4632, 
    186.4731, 189.5742, 188.8387, 188.3812, 187.0171, 186.431, 192.9768, 
    199.426,
  199.0151, 190.6845, 176.3589, 180.4333, 181.4479, 181.6985, 186.616, 
    187.87, 187.1064, 186.8554, 188.2296, 183.6629, 186.2708, 188.4037, 
    194.0096,
  198.1408, 191.2324, 183.7275, 186.1592, 190.3747, 190.3676, 192.1319, 
    188.353, 187.6899, 186.853, 181.1378, 181.8391, 185.2498, 186.5178, 
    188.7643,
  192.5396, 192.2507, 189.0368, 195.3477, 196.0856, 196.9217, 195.667, 
    191.262, 188.3313, 185.9518, 183.1693, 179.8451, 178.7339, 182.1161, 
    184.972,
  194.848, 190.7295, 198.6147, 197.2165, 200.8614, 202.3081, 200.6524, 
    196.3179, 191.5833, 187.2022, 183.582, 182.166, 178.1148, 176.9188, 
    181.6923,
  197.2846, 194.5761, 191.2558, 190.2468, 193.7702, 189.1576, 186.0648, 
    190.0979, 191.0205, 192.0688, 188.3593, 186.5598, 180.7483, 183.524, 
    175.7054,
  202.4304, 195.2897, 197.4298, 194.9698, 197.2673, 197.9768, 195.2673, 
    194.2302, 199.0659, 201.1964, 195.5134, 191.9749, 188.952, 181.519, 
    177.6234,
  203.7732, 199.7955, 200.1309, 199.1025, 201.9404, 198.0688, 205.3073, 
    195.0487, 199.3402, 203.2325, 200.7648, 198.0732, 190.2898, 186.0965, 
    179.4433,
  203.6285, 202.5577, 208.4182, 204.8752, 204.9686, 203.6425, 199.9263, 
    207.2116, 206.2802, 203.4082, 201.5924, 198.7379, 191.1424, 184.6605, 
    178.8192,
  206.5583, 207.3851, 206.0751, 207.4439, 205.2591, 202.7963, 200.0316, 
    195.0543, 195.886, 202.9286, 202.8312, 200.434, 190.8804, 179.5663, 
    176.4159,
  214.5717, 215.0639, 216.3566, 211.8743, 210.2412, 203.7949, 197.9631, 
    196.3113, 198.2539, 201.2343, 201.1795, 199.0699, 188.6667, 179.0393, 
    176.5224,
  213.5163, 216.7895, 214.3586, 216.7823, 209.0786, 205.0817, 201.3463, 
    198.7269, 200.3741, 203.1837, 202.3811, 200.1532, 192.4277, 179.6873, 
    187.0616,
  212.8973, 221.2099, 216.8221, 210.9735, 207.4065, 202.8363, 201.8147, 
    200.8392, 199.8789, 199.6657, 203.323, 200.8409, 191.2058, 183.4829, 
    188.3327,
  214.1534, 220.0982, 222.1563, 206.7186, 199.6475, 198.843, 198.6032, 
    199.7347, 199.8641, 200.5332, 198.9181, 198.8029, 190.7596, 183.473, 
    184.945,
  213.8044, 211.3777, 210.5211, 200.9383, 198.9007, 194.9827, 196.4594, 
    199.0672, 198.5957, 197.1857, 196.9198, 195.7628, 189.5258, 183.7056, 
    184.1879,
  206.1548, 203.582, 199.237, 199.7803, 200.0005, 197.1013, 196.2447, 
    197.5419, 197.3537, 197.3311, 200.9644, 199.8562, 196.8916, 197.0014, 
    196.8763,
  207.329, 203.9157, 202.7543, 199.3862, 201.2317, 194.4949, 194.4689, 
    195.1013, 194.5415, 196.9037, 198.9519, 199.9515, 202.2198, 197.5529, 
    193.6774,
  209.5594, 203.1128, 203.6109, 199.4383, 196.6102, 193.6378, 194.8535, 
    190.7597, 189.9143, 195.0948, 196.5919, 198.6909, 202.6289, 202.5037, 
    199.1684,
  214.5667, 204.7808, 202.3993, 197.306, 192.4298, 192.6382, 190.6357, 
    193.1039, 191.9202, 191.9717, 193.2602, 195.3747, 199.1501, 199.6533, 
    195.604,
  211.7811, 205.6503, 201.8193, 197.1502, 189.3844, 190.0387, 186.3022, 
    188.032, 189.8829, 189.1175, 188.2929, 190.8253, 195.5651, 197.698, 
    196.788,
  214.4216, 210.0131, 204.4001, 196.6186, 196.1474, 186.0689, 183.1988, 
    184.4669, 182.9789, 181.4974, 182.6479, 185.3961, 188.5101, 194.8584, 
    197.0494,
  213.9065, 208.7681, 205.6155, 195.6528, 193.3751, 189.314, 181.7205, 
    178.0359, 177.1046, 177.5144, 176.1882, 180.2158, 184.5107, 190.2193, 
    194.222,
  220.9957, 208.9547, 204.901, 199.4306, 195.5174, 188.0972, 183.0656, 
    177.5367, 176.2255, 172.434, 170.1585, 176.7494, 180.4561, 186.3611, 
    191.2219,
  218.1633, 208.6102, 207.6151, 198.7008, 193.8356, 187.373, 185.6059, 
    177.224, 174.4514, 170.1162, 169.9896, 172.8855, 177.3304, 183.2366, 
    190.4272,
  223.7778, 215.2543, 210.106, 204.6001, 200.4198, 196.3541, 189.1289, 
    177.7031, 170.9538, 166.4481, 165.3904, 169.0736, 176.3688, 187.3162, 
    189.5292,
  218.457, 213.6357, 204.8449, 197.8309, 187.9187, 184.757, 181.3617, 
    180.0778, 178.0043, 177.048, 184.5824, 181.501, 184.2949, 187.4601, 
    188.5303,
  221.8527, 217.5675, 208.4344, 197.6563, 193.1593, 185.9685, 183.618, 
    186.394, 183.0071, 176.4501, 177.4987, 180.8488, 181.3767, 183.8595, 
    184.1022,
  222.6816, 217.3574, 211.2475, 203.3899, 195.9711, 190.9698, 193.1258, 
    184.6821, 187.5643, 185.573, 181.5459, 175.9687, 175.3812, 176.9337, 
    179.067,
  222.6954, 218.1121, 214.8636, 206.7818, 199.7225, 199.1097, 192.8848, 
    195.7511, 182.9754, 181.2417, 184.7332, 175.0971, 173.7797, 172.9616, 
    175.1645,
  220.0379, 217.1126, 212.4258, 208.8176, 203.5215, 198.6531, 200.9077, 
    195.0869, 188.4066, 183.4005, 183.4851, 179.3611, 174.385, 170.916, 
    169.6342,
  215.8626, 213.8746, 211.3451, 210.4604, 206.8215, 202.785, 199.4277, 
    197.4801, 199.1716, 191.0664, 186.2673, 179.0843, 175.2523, 170.8303, 
    170.1946,
  217.0978, 214.6438, 209.3944, 210.8036, 208.012, 207.9573, 202.9001, 
    199.1569, 197.6122, 196.7782, 187.0616, 175.055, 172.7682, 168.4105, 
    169.0089,
  215.847, 212.1951, 210.1476, 208.3704, 211.417, 212.6128, 206.8757, 
    204.1805, 201.7312, 194.7747, 192.1855, 183.5382, 173.1461, 174.1658, 
    173.1244,
  219.3597, 215.0205, 213.2372, 208.3396, 210.0701, 211.1068, 209.0224, 
    207.8183, 201.0276, 194.139, 191.9995, 188.158, 184.2609, 178.3119, 
    186.7909,
  213.0065, 211.8813, 209.9911, 205.2364, 207.9617, 209.1562, 210.8573, 
    207.7156, 203.461, 197.8076, 195.2593, 191.7159, 189.3639, 194.1521, 
    196.6223,
  196.4029, 195.1645, 196.5609, 198.2817, 196.3573, 198.8232, 202.3237, 
    209.0046, 208.3223, 208.0555, 205.2662, 195.8904, 188.8705, 181.8445, 
    180.0645,
  197.7905, 196.844, 198.9886, 200.1402, 198.619, 202.0556, 203.4714, 
    208.9283, 212.741, 212.0211, 208.5831, 203.1958, 196.05, 188.4479, 
    178.1522,
  200.058, 204.2479, 200.8297, 196.7487, 195.8763, 201.3071, 200.2836, 
    203.2697, 209.072, 209.5098, 211.2498, 208.1571, 199.8144, 188.9184, 
    183.9104,
  199.6066, 203.6787, 200.6364, 200.4637, 194.6313, 199.5814, 201.3082, 
    207.0554, 211.793, 211.8344, 210.1496, 209.3009, 205.6172, 197.8709, 
    189.4307,
  203.2103, 206.9221, 205.8912, 202.2619, 197.3421, 196.1415, 200.9888, 
    202.9394, 206.6921, 211.2986, 211.9455, 210.0143, 206.571, 200.8557, 
    192.1951,
  209.8967, 207.474, 210.5569, 203.1209, 198.826, 194.0652, 194.9598, 
    202.1948, 206.0505, 207.6728, 211.3174, 212.6407, 211.3831, 204.9645, 
    193.6006,
  213.136, 211.2374, 209.0121, 204.0502, 200.6502, 193.1952, 193.0672, 
    196.4949, 201.2057, 203.3779, 207.7755, 211.5303, 212.587, 204.5272, 
    194.8259,
  215.4139, 216.2408, 211.9557, 205.1126, 198.8703, 197.3013, 194.1188, 
    195.7111, 199.1849, 201.2169, 202.2784, 204.0732, 207.4157, 205.3326, 
    200.4943,
  218.2118, 216.9352, 212.1138, 209.0378, 204.1055, 202.266, 202.6251, 
    193.4316, 195.2101, 196.8082, 194.3491, 199.0003, 200.0642, 201.2089, 
    201.573,
  221.7897, 219.8519, 217.0011, 216.5829, 211.4818, 206.892, 206.0479, 
    198.5188, 193.4124, 189.3858, 187.3519, 187.599, 189.4624, 193.5367, 
    195.3238,
  216.7926, 213.8332, 205.2184, 206.7472, 210.8124, 210.318, 208.3993, 
    208.4629, 210.6305, 208.6828, 204.4284, 205.4417, 206.3105, 206.4479, 
    204.9552,
  220.4058, 214.1216, 210.7044, 208.5252, 210.8151, 209.6501, 207.5516, 
    210.1651, 209.8459, 211.1986, 207.233, 205.1331, 206.9386, 209.3401, 
    209.8332,
  220.3985, 213.9716, 211.7566, 210.1564, 213.2037, 209.4326, 210.3644, 
    208.0206, 210.3341, 211.2057, 209.1116, 207.8623, 209.248, 208.2736, 
    207.9359,
  223.7091, 214.9805, 213.003, 211.2856, 212.8218, 212.8381, 210.6554, 
    210.745, 205.1854, 206.5562, 208.221, 208.2988, 211.0334, 209.8315, 
    207.8105,
  226.3378, 217.177, 209.2332, 213.1065, 216.2366, 215.2259, 216.3056, 
    210.6502, 204.3788, 206.647, 206.0729, 205.8401, 204.856, 206.7969, 
    209.866,
  226.4798, 220.0009, 213.989, 211.2061, 216.858, 215.1722, 213.601, 
    214.5273, 207.8196, 203.6124, 198.9297, 201.9949, 200.4452, 204.582, 
    206.2886,
  225.9594, 223.0263, 215.6621, 212.5823, 215.4574, 215.038, 213.4344, 
    209.7626, 204.2532, 202.2407, 195.868, 195.7097, 196.7017, 199.3414, 
    201.2333,
  225.505, 224.0929, 216.7371, 212.9614, 211.8612, 213.5429, 215.2106, 
    211.4165, 205.5958, 201.0989, 197.4512, 194.7704, 190.8714, 190.6754, 
    192.4685,
  225.9865, 223.2644, 219.2199, 214.3232, 213.3814, 213.0958, 210.0631, 
    212.1428, 205.5016, 198.2262, 200.0027, 196.3768, 194.1566, 187.2321, 
    185.2702,
  227.0634, 224.8689, 220.4396, 214.0284, 211.9955, 209.8365, 208.8968, 
    207.4934, 204.0319, 198.9921, 200.5617, 196.0731, 198.2206, 189.906, 
    186.2291,
  220.071, 219.4794, 220.3395, 220.1436, 218.2979, 213.2864, 209.6923, 
    203.8107, 198.9263, 199.6108, 200.2121, 203.8176, 200.0444, 202.7606, 
    205.4812,
  217.7406, 220.7316, 220.9887, 218.8545, 220.8669, 217.0248, 210.2102, 
    207.0806, 199.7111, 196.6764, 194.913, 197.4435, 200.3299, 199.4066, 
    202.0519,
  218.4594, 221.3238, 220.4727, 217.17, 218.8226, 214.1373, 211.3918, 
    207.2835, 198.1527, 198.9811, 190.7534, 191.4247, 190.7962, 199.8952, 
    199.98,
  218.9471, 220.8519, 219.1813, 216.9957, 214.5393, 215.0333, 210.3262, 
    210.4115, 200.6343, 189.3902, 187.154, 185.6843, 186.9435, 187.3808, 
    192.602,
  219.7728, 219.7081, 220.3507, 216.7067, 214.6262, 212.6523, 206.4096, 
    208.2865, 200.4361, 195.8122, 189.5606, 187.9827, 186.2368, 184.8418, 
    185.1542,
  220.9247, 218.7669, 219.3816, 217.315, 216.1405, 212.6808, 206.8356, 
    204.31, 201.7494, 197.0856, 194.6395, 189.8983, 186.3753, 183.669, 
    188.3913,
  221.7177, 217.9392, 218.3888, 218.5031, 215.8748, 210.4025, 208.2803, 
    205.3403, 201.9966, 200.415, 197.6091, 194.2491, 190.7686, 180.5002, 
    183.7312,
  217.3123, 217.1853, 218.8083, 220.6097, 218.0075, 210.0174, 206.8745, 
    204.2085, 201.1959, 200.2345, 197.3829, 197.2351, 194.2593, 189.0504, 
    184.3907,
  215.2104, 216.1831, 220.1309, 217.4695, 211.8417, 208.0337, 206.196, 
    204.4031, 202.0262, 200.5525, 198.0999, 197.4347, 195.2428, 190.2263, 
    191.4353,
  213.2355, 216.3051, 219.0122, 214.4634, 209.1772, 207.0375, 205.3099, 
    204.9041, 203.467, 198.1636, 196.114, 195.9322, 194.4076, 195.8883, 
    190.4465,
  215.2335, 208.3645, 201.3266, 198.6925, 199.0072, 199.6011, 201.4969, 
    204.8097, 204.6427, 197.5349, 195.6283, 186.9837, 186.9985, 186.0259, 
    180.4599,
  217.3603, 213.493, 202.5242, 200.6092, 200.0308, 200.434, 202.825, 
    204.4924, 204.4557, 200.2719, 198.3348, 191.4603, 186.6669, 181.5771, 
    179.8816,
  215.821, 214.8678, 211.306, 200.3921, 200.2895, 199.2348, 202.964, 
    201.7283, 201.8376, 202.443, 201.3091, 196.7617, 192.7219, 182.3438, 
    177.6754,
  218.3663, 208.7902, 211.1221, 206.0158, 199.9848, 200.429, 197.2842, 
    200.3962, 201.229, 201.5334, 200.8326, 201.5893, 195.1049, 188.5195, 
    179.7115,
  219.976, 212.0107, 208.3357, 206.2702, 204.2569, 199.7269, 199.093, 
    191.6789, 194.2277, 202.5747, 200.9102, 199.5272, 200.9065, 195.5229, 
    181.6685,
  217.0789, 209.3474, 209.9499, 210.0464, 211.3492, 200.1397, 195.3924, 
    196.3568, 195.3001, 193.7145, 193.1521, 196.1303, 198.6066, 197.3197, 
    186.5513,
  222.3401, 210.6646, 211.0123, 214.5823, 212.6977, 201.504, 196.4702, 
    194.362, 192.1089, 193.5618, 193.122, 194.2182, 197.285, 198.5886, 
    192.1245,
  223.358, 216.3478, 215.3778, 214.5775, 207.8474, 200.7023, 193.9998, 
    190.9617, 190.4101, 192.0275, 192.8527, 192.891, 194.5462, 196.7044, 
    195.8192,
  220.6798, 214.4574, 214.2575, 209.7445, 204.9503, 196.8745, 192.6568, 
    188.0518, 188.4822, 190.3315, 192.4523, 191.36, 192.1415, 195.1897, 
    198.216,
  224.1641, 217.0551, 211.9125, 206.8682, 205.6498, 198.3155, 193.6344, 
    190.6457, 186.8003, 186.0973, 189.306, 190.2986, 190.166, 193.1424, 
    196.672,
  217.0179, 210.2047, 204.6968, 201.1018, 197.1081, 192.1364, 194.7336, 
    195.5782, 195.3281, 193.6947, 193.4236, 196.7224, 195.4247, 189.9183, 
    180.1431,
  222.2933, 214.7289, 208.3921, 203.5285, 200.5639, 194.3168, 194.9601, 
    197.3974, 196.5188, 196.1645, 192.574, 195.7799, 197.8837, 194.3323, 
    183.8526,
  227.1446, 217.814, 209.9544, 204.6149, 200.0501, 194.5536, 196.13, 
    194.7704, 197.8677, 196.2254, 195.8864, 195.8721, 198.207, 198.3283, 
    189.1069,
  223.7091, 219.0545, 214.2392, 202.5371, 197.7754, 193.8679, 193.9023, 
    194.9404, 197.6578, 198.1724, 197.1432, 195.9009, 197.1202, 197.9625, 
    193.365,
  226.0545, 218.8793, 217.6709, 205.829, 202.0873, 189.7698, 193.7044, 
    191.8797, 195.2371, 199.7893, 198.8742, 195.9623, 195.0056, 197.1653, 
    197.1971,
  219.3335, 217.2442, 214.152, 207.5696, 203.6239, 191.6731, 184.0571, 
    187.1451, 193.6397, 192.3374, 194.7076, 195.3143, 193.6033, 195.3231, 
    198.6337,
  225.6765, 220.5412, 216.2274, 210.4449, 201.4507, 191.4541, 183.9822, 
    183.4693, 188.5721, 195.2594, 196.4034, 195.161, 194.2971, 193.7922, 
    197.8662,
  225.9279, 225.9148, 219.3999, 209.0611, 199.9612, 190.7173, 186.7796, 
    184.014, 185.7819, 190.7825, 195.3424, 194.914, 193.8841, 192.8434, 
    198.1723,
  227.7605, 227.3548, 219.407, 205.6269, 197.1561, 192.8824, 188.3547, 
    185.1122, 185.8449, 191.1102, 194.63, 193.9539, 192.1663, 192.8227, 
    197.7348,
  223.9086, 219.3437, 213.3834, 204.3581, 199.7119, 195.7428, 191.4281, 
    188.9454, 188.273, 188.8949, 193.4888, 193.0312, 190.8104, 191.6044, 
    195.5551,
  214.292, 210.5614, 206.3547, 204.9767, 203.2164, 202.5379, 198.7492, 
    193.8636, 193.7821, 197.1653, 196.256, 195.2692, 190.7118, 194.0483, 
    203.7074,
  218.5629, 217.1502, 205.9849, 202.2066, 199.7419, 196.9294, 187.0257, 
    183.4448, 189.5481, 193.5505, 195.3689, 195.6459, 195.3059, 195.8556, 
    201.212,
  222.4904, 216.0758, 211.0878, 200.5714, 189.2806, 185.3851, 177.8482, 
    174.6591, 185.2332, 192.7563, 197.0313, 196.7845, 194.4326, 191.5277, 
    198.8253,
  221.6661, 223.4129, 213.7645, 202.3492, 187.0446, 187.0911, 172.8561, 
    172.5467, 186.0879, 193.8457, 197.395, 196.3681, 193.2689, 190.5678, 
    197.1632,
  224.7344, 220.9304, 217.5364, 206.4323, 201.9144, 191.5505, 177.8058, 
    173.6808, 190.2628, 195.8011, 198.4633, 194.8384, 189.3319, 191.9705, 
    195.8727,
  228.0436, 221.0902, 217.8596, 209.9271, 211.9952, 199.7446, 179.0413, 
    173.1769, 185.9013, 195.797, 195.1772, 192.3714, 191.0043, 191.783, 
    197.5726,
  228.9958, 220.3911, 219.4967, 209.5213, 209.7151, 199.8394, 183.9307, 
    176.221, 181.7747, 196.5654, 194.8925, 191.3582, 190.6233, 192.2916, 
    197.1513,
  229.2479, 225.0169, 215.1072, 207.709, 200.0168, 193.2786, 189.5224, 
    190.3429, 194.1252, 194.5737, 194.282, 190.7103, 189.692, 194.212, 
    193.2007,
  228.9202, 226.9181, 215.9567, 206.64, 200.4834, 194.7494, 194.6315, 
    197.8137, 194.8112, 193.9961, 192.1856, 191.5606, 192.0083, 195.031, 
    196.0285,
  226.6973, 217.003, 212.6904, 205.3562, 203.6986, 202.7961, 200.8331, 
    200.1687, 196.7096, 192.1779, 191.3356, 190.9895, 193.5187, 194.1897, 
    196.2016,
  214.4465, 210.868, 207.3008, 203.289, 196.4825, 196.7529, 202.7814, 
    203.6153, 190.0631, 178.7191, 183.2891, 192.7206, 195.4894, 200.36, 
    202.6763,
  221.0699, 217.2081, 209.8939, 203.5816, 194.7547, 194.8265, 200.7621, 
    201.1562, 188.5182, 178.7509, 183.1828, 193.2783, 197.1636, 202.8053, 
    202.8679,
  223.8147, 223.4434, 218.5622, 205.239, 192.5612, 186.6533, 196.3008, 
    191.7575, 181.098, 174.6514, 185.8315, 195.1749, 200.5794, 207.0082, 
    206.6506,
  227.5158, 221.8702, 224.3876, 208.8663, 193.2434, 186.8744, 181.9066, 
    182.1765, 175.5237, 175.7475, 194.5734, 200.9908, 202.4412, 207.9859, 
    207.4635,
  225.743, 225.2352, 224.7828, 208.3005, 201.323, 180.6731, 180.5594, 
    182.9059, 182.4098, 190.1138, 198.7113, 201.4998, 205.4601, 207.8024, 
    208.4174,
  229.9282, 225.3691, 219.9906, 209.0173, 208.2468, 191.4774, 182.7218, 
    181.295, 188.974, 195.9832, 196.102, 200.7775, 204.7285, 205.7864, 
    208.9106,
  228.3596, 227.3452, 217.6125, 212.2793, 209.3554, 201.1358, 197.6017, 
    194.0447, 196.3031, 196.1842, 197.2021, 199.5365, 201.7598, 205.4232, 
    210.0318,
  231.0935, 226.5106, 217.6205, 207.4949, 203.9574, 202.255, 199.6285, 
    197.6875, 197.1139, 197.8357, 198.6627, 195.1006, 198.1611, 207.193, 
    207.9164,
  229.8016, 227.2988, 209.5396, 203.4928, 203.0205, 200.1549, 199.809, 
    197.6196, 196.1108, 193.6917, 189.5925, 189.5226, 197.3262, 204.7766, 
    204.533,
  228.563, 218.1, 208.9439, 203.4815, 202.0921, 198.4459, 195.4902, 194.399, 
    186.9175, 183.306, 184.6788, 187.753, 194.9435, 201.2827, 199.2237,
  203.5143, 206.0446, 205.0388, 201.17, 197.4945, 184.3704, 178.625, 
    178.6781, 190.3707, 192.1323, 185.9184, 180.8754, 184.0455, 185.7675, 
    193.6918,
  212.1207, 214.7705, 208.2149, 200.9571, 193.2948, 184.173, 173.6497, 
    169.7446, 178.8963, 180.2898, 180.548, 174.3962, 180.8952, 184.1782, 
    193.7964,
  215.9855, 225.0704, 221.9261, 201.3685, 191.8453, 178.681, 174.1921, 
    167.8884, 168.8806, 170.5006, 179.7452, 180.2897, 181.5222, 180.6459, 
    197.9247,
  222.9097, 228.1147, 222.5803, 207.8345, 192.7634, 181.3592, 173.9854, 
    175.5132, 174.0674, 173.805, 177.741, 185.4231, 189.9476, 195.8418, 
    203.8002,
  225.5943, 221.2764, 223.3723, 208.8014, 202.6061, 186.5293, 182.6719, 
    178.2532, 177.4826, 179.5142, 187.1105, 198.7933, 205.4676, 207.7679, 
    209.2511,
  223.7612, 224.1199, 216.5503, 213.8796, 210.0168, 203.0823, 189.5998, 
    189.448, 191.946, 201.5305, 204.7614, 207.8954, 209.0983, 207.9067, 
    210.1088,
  228.4962, 223.3897, 223.515, 211.0448, 208.7319, 206.2571, 206.7189, 
    205.0444, 205.1569, 205.2114, 206.5767, 208.2175, 210.0591, 209.7116, 
    211.4817,
  224.8844, 224.6911, 206.3974, 209.1878, 207.584, 206.2937, 208.2723, 
    209.2684, 208.6205, 207.9858, 207.8969, 208.0649, 208.8209, 210.2464, 
    211.4027,
  228.4929, 216.8124, 215.4933, 203.6931, 202.7292, 205.279, 207.6046, 
    207.7059, 207.5824, 207.4138, 206.4287, 210.3536, 210.6447, 210.6786, 
    211.3041,
  231.2315, 220.948, 210.5079, 203.1783, 193.5072, 189.8618, 193.7226, 
    199.4582, 205.1021, 195.2464, 203.6221, 209.0799, 211.7205, 212.3867, 
    210.2487,
  216.3712, 208.7606, 199.0186, 192.7905, 192.7878, 191.9724, 192.2158, 
    196.3782, 191.4882, 190.1826, 186.4914, 197.3437, 202.5925, 205.3976, 
    203.0442,
  220.9943, 215.0756, 204.1584, 200.1178, 198.8915, 198.8669, 195.8189, 
    197.142, 195.3243, 189.7857, 182.8786, 186.2141, 202.976, 203.4158, 
    203.2004,
  220.0597, 222.1709, 209.5518, 204.0131, 203.1259, 198.984, 203.9165, 
    199.5844, 197.178, 195.9853, 184.252, 179.2029, 192.3636, 208.1459, 
    206.6915,
  215.1646, 220.6772, 209.5912, 206.5675, 202.7871, 203.9288, 202.8759, 
    207.3942, 206.4289, 200.7083, 192.9867, 182.9892, 183.1239, 196.4857, 
    203.4201,
  211.0051, 212.8074, 211.238, 210.3204, 207.0822, 202.0351, 206.7099, 
    200.9591, 202.1749, 208.0996, 201.9302, 194.5068, 188.6933, 194.909, 
    198.5913,
  210.6426, 199.0356, 204.4802, 208.197, 208.2408, 204.0422, 204.5269, 
    204.1973, 203.9479, 207.9035, 207.0968, 204.2134, 200.3213, 198.8611, 
    199.0072,
  209.5985, 199.3, 198.323, 206.0618, 207.0761, 202.3503, 204.3851, 201.378, 
    202.3553, 210.2022, 209.5144, 207.6566, 205.0944, 205.8004, 202.7188,
  209.1674, 196.3837, 199.9214, 201.9204, 205.7046, 203.6747, 203.0758, 
    202.1399, 197.9777, 211.4191, 211.2928, 210.3399, 208.262, 206.9839, 
    207.7005,
  208.3096, 197.9008, 193.8215, 198.8365, 202.9001, 201.3854, 200.375, 
    202.027, 197.3017, 211.053, 213.1228, 212.1379, 209.7272, 207.6004, 
    204.5805,
  206.2921, 194.7946, 192.1901, 196.9189, 204.5526, 201.9482, 200.3255, 
    204.798, 201.3727, 202.1422, 213.4546, 213.1113, 212.0052, 208.9344, 
    204.2773,
  215.1974, 201.9777, 192.6148, 195.6463, 199.0271, 194.1724, 193.3956, 
    203.857, 204.7444, 198.8199, 194.3218, 200.1299, 203.097, 203.1749, 
    191.2893,
  211.004, 204.7484, 199.6612, 196.2993, 199.4656, 192.1448, 194.2133, 
    208.4339, 203.665, 198.9014, 196.5788, 199.9329, 205.6552, 205.5763, 
    200.1202,
  209.465, 211.3991, 203.1317, 196.3242, 197.5287, 194.198, 201.1141, 
    204.6759, 200.0593, 200.1413, 200.1439, 201.6451, 205.5539, 207.3452, 
    208.1321,
  209.9187, 216.1615, 203.6693, 193.9247, 189.7509, 196.6147, 202.1641, 
    211.7708, 205.6832, 203.818, 200.6839, 202.5205, 201.6587, 200.8994, 
    205.3062,
  216.5579, 217.4366, 206.6708, 190.8752, 194.1979, 203.8737, 210.1583, 
    203.8496, 200.9125, 209.1698, 202.301, 201.4781, 197.5489, 196.3912, 
    195.4422,
  220.8468, 220.6706, 207.3007, 191.2999, 195.524, 207.8983, 207.4733, 
    209.6886, 206.787, 207.2988, 204.8059, 202.6547, 198.706, 196.316, 
    188.6089,
  218.5962, 226.3965, 200.4832, 191.6486, 203.4263, 211.4864, 207.4823, 
    211.3971, 207.8043, 207.65, 206.3488, 202.8849, 199.4843, 194.7917, 
    186.4184,
  221.4837, 218.2825, 197.3994, 194.771, 209.372, 211.3618, 208.7185, 
    211.9778, 210.8335, 208.9263, 204.148, 201.6562, 198.4669, 197.5729, 
    192.0519,
  218.9021, 219.6359, 202.3946, 199.9332, 211.2493, 209.2988, 208.1123, 
    211.9172, 210.0431, 208.4859, 206.2944, 202.2018, 198.3376, 196.9529, 
    196.0341,
  221.5526, 219.6376, 208.7655, 202.492, 212.5191, 207.6433, 207.5515, 
    212.5087, 211.6134, 214.4697, 209.2271, 208.8763, 200.637, 198.9351, 
    194.6666,
  221.4283, 218.7423, 217.2774, 215.8379, 210.4825, 205.6954, 206.5482, 
    206.4134, 207.6723, 209.3322, 208.3925, 203.8851, 199.3304, 201.8508, 
    207.3199,
  220.773, 219.502, 219.5323, 216.2967, 211.2583, 212.3029, 209.7869, 
    211.1734, 209.9158, 211.3909, 207.5015, 204.1617, 200.1847, 201.8656, 
    207.2556,
  222.7271, 222.9871, 220.7523, 215.0454, 214.5021, 213.3181, 212.3441, 
    210.0819, 211.2244, 210.3093, 209.3244, 203.5728, 198.3035, 198.9598, 
    206.1947,
  220.4566, 217.2072, 223.2321, 213.1534, 212.0257, 216.3581, 210.9713, 
    212.5255, 208.8476, 210.0089, 210.5379, 202.154, 196.3617, 198.1373, 
    203.4454,
  217.8723, 215.5782, 220.1119, 215.3938, 213.9859, 212.0663, 212.4025, 
    204.7497, 202.7957, 211.1828, 205.5242, 201.6341, 197.9792, 201.586, 
    202.1794,
  217.088, 215.9673, 211.3587, 219.6226, 212.4005, 211.3394, 207.3227, 
    208.8697, 209.288, 209.7077, 205.5529, 207.8404, 203.7451, 203.2457, 
    202.7007,
  213.8765, 214.6574, 208.8948, 212.6384, 209.4198, 212.008, 208.3386, 
    208.1523, 209.527, 208.1764, 207.1993, 210.005, 203.0856, 206.3874, 
    204.387,
  213.8052, 213.6329, 208.4123, 206.5268, 206.1087, 212.1136, 208.7852, 
    209.3515, 210.592, 207.8976, 208.3396, 210.0488, 207.9467, 205.4444, 
    204.9995,
  218.3973, 214.2665, 209.9097, 206.2223, 205.5788, 211.3121, 209.461, 
    209.0024, 211.8518, 207.8734, 208.4369, 208.5387, 208.8782, 206.4368, 
    206.9441,
  218.5958, 215.6901, 213.453, 208.0023, 205.9565, 211.4395, 209.0589, 
    209.5195, 209.1039, 207.7284, 206.9098, 206.3792, 209.0707, 210.1084, 
    212.4212,
  226.4495, 219.2022, 214.9901, 210.2153, 208.8119, 211.0417, 211.1232, 
    211.0418, 210.5122, 208.759, 209.1054, 208.3499, 206.9655, 205.784, 
    204.7571,
  223.4687, 220.7908, 212.2733, 210.1633, 206.3081, 206.8846, 211.0251, 
    210.5379, 211.3802, 209.9831, 208.2757, 206.2497, 206.2565, 204.245, 
    205.5463,
  219.5023, 216.5967, 211.1857, 209.6049, 205.9632, 206.2887, 210.1828, 
    208.9412, 207.6988, 207.4097, 208.271, 204.9046, 204.74, 204.2362, 
    204.9128,
  219.8314, 214.4139, 206.5877, 207.2273, 204.7843, 208.6506, 208.0974, 
    209.4508, 208.1179, 204.382, 204.7932, 205.086, 204.6656, 204.978, 
    205.1877,
  221.9895, 208.7922, 207.6423, 209.0228, 205.3049, 207.034, 210.8808, 
    206.3621, 204.0633, 204.2222, 205.9109, 206.103, 205.9177, 206.5012, 
    206.5013,
  221.1709, 209.7562, 209.7597, 208.9544, 207.9645, 210.6564, 209.9202, 
    204.9323, 203.5371, 203.8288, 206.8529, 208.6059, 208.2194, 209.3815, 
    210.2743,
  217.1559, 207.9696, 212.3182, 209.4426, 212.1483, 213.348, 210.3474, 
    201.6214, 202.2011, 206.1369, 208.8936, 208.4622, 211.0721, 208.9952, 
    212.7004,
  215.0783, 210.062, 215.8625, 210.1991, 211.5893, 213.6479, 207.6161, 
    203.5205, 206.1047, 205.9129, 208.9799, 208.3484, 207.2304, 208.088, 
    212.3489,
  213.1326, 208.7755, 214.1783, 209.2379, 212.4655, 215.0759, 208.6838, 
    205.457, 206.9546, 208.1858, 204.6175, 203.9207, 205.5847, 206.3062, 
    208.0286,
  207.6298, 211.0819, 213.55, 208.0321, 212.9721, 214.332, 208.846, 208.598, 
    209.4141, 206.7314, 201.8384, 203.1115, 199.7613, 202.2676, 203.9997,
  208.4208, 208.5713, 209.8384, 203.8512, 211.6441, 210.5623, 209.8762, 
    210.1002, 210.7566, 206.2904, 205.4528, 204.3831, 203.2318, 204.8571, 
    204.3227,
  209.4193, 211.0552, 209.2162, 210.1295, 216.2807, 214.4006, 212.8272, 
    211.2071, 211.1767, 207.3837, 207.8058, 202.6086, 200.2924, 199.5676, 
    202.4519,
  210.426, 215.0532, 208.6301, 211.2331, 216.5959, 214.4506, 214.0595, 
    207.9801, 209.9122, 207.2102, 204.9422, 199.4211, 202.118, 204.2839, 
    203.1168,
  208.7014, 216.3897, 209.0013, 209.589, 216.7141, 216.2175, 210.3734, 
    211.6032, 210.6251, 206.7251, 204.1132, 201.6385, 203.072, 204.902, 
    202.9083,
  215.6525, 208.3419, 208.988, 211.9646, 218.9573, 215.696, 214.5499, 
    205.7938, 206.4829, 205.0626, 200.6222, 201.9324, 203.2851, 205.2307, 
    207.6505,
  213.0276, 209.424, 210.6168, 211.2956, 217.8905, 215.7085, 212.1251, 
    208.4742, 203.8643, 200.0789, 200.9479, 194.3124, 199.1577, 206.8313, 
    206.7145,
  211.8381, 209.4611, 210.9905, 212.4401, 216.6739, 216.027, 213.7851, 
    209.1621, 205.1008, 202.5514, 200.2539, 198.1667, 198.9594, 205.0041, 
    211.3379,
  214.8389, 209.902, 226.6417, 214.2281, 216.5925, 217.4871, 215.5411, 
    211.4599, 205.605, 203.4724, 199.6502, 195.0461, 198.6174, 199.6171, 
    208.2754,
  213.5019, 210.4243, 221.7369, 215.2259, 214.8892, 217.4313, 214.8994, 
    212.8468, 208.9116, 204.754, 201.9232, 201.3048, 196.587, 202.445, 
    202.5006,
  212.2641, 211.8798, 216.006, 214.5944, 214.363, 215.9081, 215.0664, 
    219.2161, 212.3759, 207.4195, 204.3024, 196.1763, 192.8184, 196.9203, 
    197.6914,
  221.7586, 218.8247, 217.5538, 214.5744, 210.752, 208.8207, 206.8058, 
    207.2036, 207.4143, 208.892, 207.7984, 207.8372, 207.7112, 205.6353, 
    204.8306,
  223.1312, 221.6472, 218.476, 215.1204, 213.065, 208.7809, 206.4227, 
    206.7616, 206.2264, 207.0051, 204.2823, 205.5485, 207.2723, 207.516, 
    205.3655,
  215.324, 217.017, 219.8907, 217.5352, 213.2409, 208.7311, 207.7394, 
    204.6867, 204.7593, 206.5169, 205.3637, 207.0712, 205.9716, 202.0217, 
    203.3842,
  213.0617, 207.9957, 209.6396, 216.326, 212.713, 209.4567, 206.4468, 
    206.3654, 206.2483, 206.1616, 206.243, 206.7465, 205.1051, 201.9633, 
    199.475,
  211.6616, 205.0328, 210.4075, 214.2746, 213.0138, 206.1067, 206.063, 
    202.6609, 206.2066, 206.0136, 205.9281, 207.6724, 206.5927, 198.7765, 
    198.8179,
  206.4091, 205.1558, 210.5676, 213.0896, 211.4082, 205.7688, 203.1889, 
    204.8793, 202.5792, 200.3276, 200.061, 206.5493, 205.9452, 202.8603, 
    196.8742,
  206.2662, 208.2098, 212.291, 215.1614, 211.8208, 208.9693, 205.067, 
    199.9598, 196.333, 198.3006, 203.56, 206.1389, 205.9676, 200.3827, 196.864,
  206.0578, 211.2836, 219.2206, 211.1092, 208.9361, 206.4354, 204.6296, 
    201.5084, 198.976, 201.3671, 202.2117, 206.75, 206.4825, 200.9277, 
    200.9365,
  209.9196, 215.0152, 213.904, 207.5204, 206.5232, 203.1787, 200.9126, 
    199.1331, 199.1673, 199.7862, 203.7617, 203.4296, 206.5686, 202.7925, 
    197.0316,
  213.8462, 222.4572, 209.9452, 205.5997, 204.1547, 202.6167, 201.601, 
    202.8934, 201.7207, 201.2527, 202.972, 203.6548, 204.052, 201.5012, 
    199.414,
  205.2905, 208.7325, 206.5909, 208.3873, 210.0842, 212.6839, 211.011, 
    210.8793, 211.4076, 210.923, 210.9535, 208.7597, 209.6779, 207.4663, 
    206.1119,
  204.7318, 208.0542, 208.5127, 210.5737, 214.396, 217.941, 214.3382, 
    212.2319, 210.615, 206.7784, 209.0819, 208.5729, 211.194, 207.9205, 
    206.3437,
  206.7175, 212.1747, 216.4656, 215.1968, 218.4201, 217.3128, 212.7713, 
    206.9238, 203.7081, 206.4485, 208.678, 208.1841, 210.7327, 211.5107, 
    209.4193,
  215.182, 219.1766, 220.5238, 217.0623, 218.6312, 215.774, 212.6488, 
    211.0016, 202.8768, 200.556, 205.4508, 206.715, 207.2419, 209.0432, 
    210.0433,
  216.8705, 224.3958, 219.0889, 220.3201, 218.7354, 212.0188, 207.8379, 
    209.0858, 204.3936, 203.2365, 200.0278, 199.7766, 197.4083, 198.2064, 
    199.4951,
  220.9385, 221.9126, 221.2772, 224.9893, 220.361, 207.8941, 203.9642, 
    201.7003, 204.6842, 200.7231, 198.2237, 196.9195, 195.4253, 195.3369, 
    194.0008,
  221.293, 220.5235, 218.3087, 223.0343, 215.442, 206.291, 201.8578, 
    198.3215, 195.7126, 199.1197, 200.3383, 201.0779, 198.0554, 198.8461, 
    194.6202,
  218.1588, 217.8283, 220.8838, 217.8776, 209.2564, 204.0114, 200.6469, 
    200.2542, 203.8262, 205.0877, 204.2076, 203.1349, 201.2232, 198.3282, 
    198.7099,
  217.4681, 219.6633, 224.1386, 212.0292, 207.7375, 205.6066, 206.5114, 
    209.7107, 207.2742, 207.5754, 206.9857, 206.0105, 203.6563, 201.6535, 
    200.8546,
  221.8506, 229.0494, 215.6104, 211.2146, 211.4289, 211.9212, 212.242, 
    212.4491, 209.4376, 208.8131, 209.2789, 208.8392, 206.3357, 203.6508, 
    203.2204,
  208.7178, 200.2657, 197.8855, 196.0196, 198.8531, 212.2521, 221.1295, 
    218.4628, 216.8068, 217.4326, 211.4062, 203.9892, 203.7425, 207.0433, 
    207.0475,
  209.2728, 204.4526, 201.4837, 198.1444, 208.1522, 219.4404, 217.4665, 
    215.5898, 211.4719, 205.2618, 203.3016, 199.9845, 201.1053, 201.3394, 
    204.4057,
  213.6707, 201.9014, 203.1478, 205.5165, 222.4809, 218.8649, 217.9644, 
    212.2103, 210.6914, 202.9394, 200.2245, 195.7047, 194.1911, 198.4397, 
    200.4184,
  211.6335, 207.1632, 207.854, 210.6236, 216.8429, 219.2897, 215.5632, 
    217.2023, 210.5288, 196.8445, 195.8993, 193.674, 190.7869, 193.4489, 
    197.4683,
  211.3414, 206.7121, 214.1833, 218.8034, 215.9249, 213.3207, 212.8326, 
    207.587, 202.9718, 199.1195, 198.503, 200.7573, 199.1279, 203.8644, 
    202.5115,
  211.1175, 211.9548, 222.5787, 221.8089, 217.7428, 213.1049, 210.9174, 
    207.155, 204.0002, 203.3202, 205.1363, 207.0685, 209.2155, 210.0291, 
    209.961,
  214.9498, 220.9496, 224.9108, 219.8656, 216.2037, 214.0844, 212.0972, 
    209.3781, 208.1941, 210.0482, 208.8505, 208.7946, 208.6661, 210.472, 
    211.6743,
  219.5278, 221.5724, 228.6902, 218.2201, 215.1701, 214.9181, 214.2955, 
    212.3184, 208.1051, 206.4038, 205.1864, 205.4891, 204.396, 203.6744, 
    206.5391,
  220.8152, 223.0073, 223.9911, 215.9202, 213.8755, 214.1054, 211.8464, 
    209.3041, 207.5873, 205.8804, 204.2406, 205.9324, 203.4602, 202.8522, 
    202.7489,
  221.0089, 222.4189, 222.3887, 211.65, 213.2933, 212.7563, 210.2966, 
    212.7098, 206.9288, 203.7329, 201.764, 205.2366, 206.6268, 205.0517, 
    205.4792,
  225.6842, 225.1984, 221.9202, 219.1975, 218.5366, 214.1122, 214.1526, 
    212.8243, 213.1184, 208.2603, 205.4632, 201.476, 197.1813, 195.895, 
    187.8942,
  223.4327, 221.6118, 221.9239, 218.5773, 217.1453, 215.4261, 214.424, 
    214.5197, 214.6329, 211.0028, 208.1447, 204.0284, 199.2045, 194.1094, 
    195.0205,
  222.3654, 221.3958, 218.9507, 216.5856, 216.0728, 210.8785, 213.9826, 
    212.2828, 209.9, 212.6102, 212.3651, 209.8047, 206.091, 199.9581, 196.5499,
  220.2886, 220.4129, 220.6428, 212.5916, 212.6932, 212.6005, 208.3446, 
    210.9148, 212.4102, 210.027, 210.8367, 210.7277, 210.4364, 203.375, 
    201.3276,
  220.4326, 217.9833, 219.2173, 213.0257, 211.312, 208.8499, 209.821, 
    204.7531, 203.6665, 207.9755, 209.2261, 207.8924, 208.6635, 209.1296, 
    208.0005,
  218.8983, 216.9592, 216.7886, 214.2413, 211.3727, 210.2749, 206.9124, 
    203.169, 201.2727, 204.481, 208.0195, 206.7687, 206.608, 208.2566, 
    207.1581,
  218.7353, 218.034, 215.5282, 211.707, 209.3167, 208.1299, 205.04, 204.1204, 
    205.3701, 204.3087, 208.6947, 208.1308, 204.8403, 206.2804, 207.5595,
  217.1646, 217.0435, 216.9771, 214.1133, 208.2392, 206.4717, 204.1308, 
    204.2102, 206.5083, 207.3125, 204.2044, 205.6999, 205.7177, 205.6043, 
    204.4301,
  213.6388, 217.5098, 217.3119, 212.8048, 207.5031, 206.1256, 204.1553, 
    202.5688, 204.3644, 205.3341, 204.0077, 202.9769, 208.1369, 210.3567, 
    208.8008,
  211.2041, 215.1341, 215.1602, 210.8642, 203.7152, 201.9358, 202.3982, 
    205.8856, 205.7832, 204.0014, 203.8074, 202.8329, 210.6222, 210.7317, 
    211.5882,
  194.9016, 199.5718, 199.8492, 206.891, 206.8501, 203.9887, 194.4277, 
    197.4158, 200.1229, 205.7645, 209.8279, 207.9146, 211.1421, 205.5823, 
    201.7758,
  194.3294, 195.7458, 196.462, 205.6994, 204.937, 201.366, 193.5338, 190.705, 
    196.9553, 201.0169, 204.8093, 206.7794, 208.4851, 208.7656, 206.7908,
  191.8129, 192.1177, 195.6976, 199.0034, 202.2685, 202.5372, 196.8471, 
    187.1874, 189.5236, 198.5979, 203.4029, 206.7779, 208.55, 211.1342, 
    210.0406,
  191.0989, 188.7255, 193.7277, 197.5811, 196.2113, 197.086, 191.1027, 
    188.5621, 189.2259, 195.3754, 199.4944, 204.2478, 207.8284, 210.679, 
    210.7503,
  186.8399, 190.8367, 190.6777, 197.544, 196.2773, 187.8594, 185.5719, 
    186.0413, 191.5577, 193.422, 199.8663, 201.3698, 205.6294, 210.2421, 
    209.9334,
  193.8723, 188.8303, 190.5712, 197.0023, 201.4165, 189.2908, 180.6966, 
    182.1271, 188.2828, 190.67, 195.6526, 202.4165, 205.9784, 209.2787, 
    207.8446,
  193.3075, 190.9227, 192.8076, 199.0365, 201.8724, 193.7164, 184.9014, 
    186.0846, 189.4639, 197.1359, 195.073, 200.9711, 205.8263, 208.3045, 
    208.6347,
  191.8577, 185.8233, 194.3833, 203.3614, 201.3979, 190.6669, 194.0496, 
    191.9996, 191.9265, 198.2413, 197.8728, 203.3017, 205.2839, 208.4495, 
    209.4296,
  193.6522, 186.0549, 197.8122, 206.4707, 197.3633, 197.0831, 196.2448, 
    194.4493, 196.0529, 196.7994, 199.7858, 203.9715, 204.9, 208.8522, 
    208.9747,
  190.1815, 191.8447, 205.503, 204.6746, 198.915, 203.6635, 200.915, 
    197.9397, 201.887, 200.5729, 202.2691, 204.3232, 205.3697, 207.5764, 
    205.793,
  198.7191, 190.9124, 184.351, 186.5214, 183.2448, 180.4183, 180.4471, 
    183.6386, 183.8327, 186.9158, 188.0655, 193.8343, 205.4789, 212.1704, 
    210.5441,
  198.5887, 197.1272, 195.863, 194.8089, 190.8893, 183.6766, 183.697, 
    188.2243, 190.1003, 193.5676, 194.5255, 193.4834, 201.2501, 209.2324, 
    208.9426,
  207.7044, 205.9643, 204.4274, 199.2424, 193.6254, 190.7629, 197.8586, 
    192.8564, 197.1591, 204.7641, 206.3521, 197.3524, 199.0137, 207.1042, 
    210.0941,
  207.9875, 207.345, 206.1398, 198.4783, 196.8001, 202.6471, 210.3714, 
    209.8868, 207.212, 207.9579, 206.2549, 197.7302, 198.5438, 202.0257, 
    206.7055,
  211.4952, 209.8596, 206.6298, 204.9468, 204.9001, 212.4918, 215.955, 
    213.4783, 208.9282, 211.1626, 202.1527, 195.3865, 193.9271, 198.9678, 
    204.003,
  211.7323, 210.0087, 204.8898, 207.7013, 209.582, 209.4287, 211.0666, 
    214.9365, 214.6613, 210.8009, 204.0862, 195.9405, 190.7563, 193.0249, 
    203.5128,
  215.0042, 206.2391, 208.0084, 214.3159, 215.3561, 214.8432, 215.5105, 
    213.8969, 211.7485, 212.3133, 208.2225, 194.2216, 189.8416, 191.4868, 
    201.3814,
  213.3038, 207.8023, 213.8714, 215.6552, 214.1278, 216.1755, 214.7642, 
    211.7996, 211.6018, 211.446, 206.9653, 201.1332, 192.4281, 195.4709, 
    202.2236,
  207.7593, 202.3087, 210.151, 213.2635, 215.3003, 214.9986, 211.5515, 
    211.4656, 210.3745, 210.3356, 208.3152, 205.4394, 203.9198, 207.1201, 
    208.0226,
  205.2333, 203.6874, 213.76, 214.8438, 215.7258, 214.3247, 213.1901, 
    212.1838, 211.1499, 208.6147, 204.4382, 204.3745, 202.8694, 204.8223, 
    206.4987,
  220.7596, 214.5732, 215.263, 219.7837, 217.706, 216.6887, 216.4428, 
    213.0911, 209.6466, 205.5109, 200.7671, 193.273, 189.1486, 192.0054, 
    198.6525,
  213.6536, 214.862, 217.7604, 216.5249, 220.7441, 215.6041, 213.9485, 
    213.4974, 212.9386, 208.1093, 207.2748, 196.4571, 190.1374, 192.7561, 
    194.7002,
  211.1512, 209.0226, 215.8225, 215.7814, 219.2932, 213.7524, 213.7763, 
    211.8174, 210.8691, 210.67, 214.9053, 210.9226, 191.8097, 189.9304, 
    191.5599,
  210.6299, 207.2696, 212.2875, 214.5802, 216.8806, 215.5794, 208.7538, 
    211.4712, 213.3525, 212.4876, 210.3054, 201.5616, 191.236, 186.0054, 
    190.9271,
  209.5842, 205.0472, 216.2489, 213.4336, 211.7889, 209.7646, 210.8057, 
    205.3203, 202.8699, 209.4677, 203.6555, 198.7172, 191.5714, 188.5697, 
    193.2853,
  216.4931, 205.7927, 210.6579, 212.4288, 210.0544, 208.8206, 206.5964, 
    206.9087, 206.6299, 208.1916, 202.6481, 199.1518, 192.8197, 189.2853, 
    195.7274,
  215.5202, 207.6236, 212.9353, 210.927, 208.3485, 205.2645, 206.1444, 
    205.4946, 205.6832, 208.1703, 202.7826, 192.3991, 193.4556, 193.3426, 
    195.3221,
  213.4, 209.476, 211.8046, 208.0486, 206.1078, 204.1001, 204.0722, 205.7434, 
    205.9095, 209.0577, 207.5007, 199.9039, 189.7436, 192.0814, 197.0455,
  213.5242, 211.3511, 210.6333, 206.3134, 202.5938, 200.996, 201.1556, 
    202.2371, 204.2847, 207.1736, 208.3132, 207.7329, 201.4919, 201.108, 
    204.7219,
  218.8281, 214.151, 208.4927, 203.7653, 200.1267, 198.6495, 198.3658, 
    201.7615, 205.3648, 206.3779, 206.8307, 205.3196, 206.7888, 207.0044, 
    209.459,
  215.8522, 207.3129, 206.2015, 203.0809, 203.2925, 204.8971, 206.7092, 
    206.6793, 207.7493, 208.0136, 208.3296, 209.4715, 213.7303, 213.1624, 
    211.7468,
  210.6851, 211.5652, 206.4701, 201.7822, 206.3891, 205.4568, 205.2224, 
    208.1605, 208.375, 207.944, 209.4372, 209.7869, 210.1781, 213.9753, 
    216.1503,
  211.025, 203.7319, 204.6398, 202.9073, 203.9174, 206.3856, 206.7607, 
    203.8645, 206.6049, 204.7777, 204.9022, 207.0675, 214.7743, 215.0037, 
    211.6801,
  209.1158, 209.716, 205.6328, 202.6223, 202.9918, 203.9452, 205.0354, 
    205.848, 207.7362, 197.4042, 194.6075, 195.0537, 198.5791, 205.6908, 
    202.3943,
  216.3023, 209.9089, 201.1706, 200.0401, 201.5113, 203.6552, 204.7838, 
    204.3591, 204.5481, 196.0882, 188.2726, 190.3833, 192.566, 195.3401, 
    194.2039,
  219.2076, 208.0967, 202.3906, 199.7662, 206.7408, 202.1307, 201.582, 
    207.1471, 205.5693, 194.1148, 185.4245, 185.6745, 186.7332, 189.0249, 
    190.7696,
  219.3987, 208.6119, 203.8756, 200.3358, 205.2919, 203.3964, 204.4867, 
    203.8973, 207.1463, 198.7481, 190.0588, 182.5637, 182.924, 186.2499, 
    189.3397,
  218.0446, 208.7365, 204.5284, 200.0976, 204.9812, 204.3533, 206.3356, 
    206.5802, 209.5686, 202.645, 194.3592, 188.2745, 181.2591, 180.3932, 
    185.2811,
  219.7886, 206.9057, 202.2033, 201.5911, 205.8828, 210.3155, 208.214, 
    208.0145, 209.2691, 207.9871, 199.7842, 191.6134, 190.5717, 188.9513, 
    197.7932,
  217.9955, 210.5536, 210.7611, 206.2036, 208.1569, 210.1306, 210.495, 
    209.135, 209.5898, 209.8201, 207.0321, 201.5923, 198.4763, 202.1124, 
    208.3136,
  209.0685, 208.7702, 215.2573, 213.0664, 212.9187, 208.4389, 206.4749, 
    203.9941, 206.0834, 207.2601, 209.1436, 205.7506, 199.7213, 195.1, 
    198.9284,
  205.7925, 213.3794, 217.1063, 214.1449, 213.1394, 209.5518, 205.5283, 
    203.1317, 206.0806, 207.8746, 210.8396, 207.5723, 208.4881, 204.3869, 
    203.4977,
  206.5654, 214.7948, 215.6559, 216.748, 213.8801, 206.9406, 204.2122, 
    192.9025, 190.5713, 206.3913, 210.7835, 207.8469, 210.0323, 210.6151, 
    208.4829,
  201.9855, 214.1902, 213.5734, 213.103, 212.8657, 210.2094, 199.7311, 
    188.3126, 186.7932, 193.4458, 208.6563, 210.9627, 210.6477, 215.65, 
    212.9475,
  206.088, 216.5516, 213.0279, 212.707, 211.9621, 208.5408, 206.1383, 
    191.0094, 186.1782, 183.207, 192.2671, 211.1273, 212.7745, 209.5003, 
    210.2996,
  203.6873, 218.8093, 215.045, 214.3293, 211.5242, 208.5411, 206.9306, 
    192.0626, 181.1075, 180.3371, 180.7973, 194.5895, 211.3045, 215.2907, 
    212.4467,
  204.5414, 218.7706, 217.3787, 211.1368, 210.6695, 209.4642, 207.4475, 
    199.5916, 183.6523, 177.5881, 172.9659, 182.6044, 196.5864, 213.7842, 
    217.156,
  206.9694, 215.6164, 215.4555, 212.2632, 210.8021, 210.1013, 210.4053, 
    207.568, 194.7158, 181.836, 177.6588, 178.5336, 185.7358, 201.9395, 
    214.2867,
  208.7805, 217.3818, 214.4534, 211.3812, 210.6935, 210.1123, 210.956, 
    209.2254, 205.0367, 189.1124, 180.535, 179.981, 182.271, 187.722, 203.5424,
  204.9276, 218.1244, 221.5201, 210.608, 210.08, 209.7476, 210.1441, 
    210.5074, 210.5765, 203.3786, 188.1952, 186.8497, 189.7676, 188.5345, 
    194.9258,
  197.0694, 198.2854, 205.3055, 214.9963, 212.5647, 210.902, 198.2332, 
    193.6427, 202.3385, 214.0764, 209.8361, 210.0238, 210.4125, 198.689, 
    196.139,
  195.2742, 201.206, 212.9952, 215.7723, 216.0399, 209.2414, 194.5064, 
    195.2895, 201.9547, 211.906, 213.6413, 210.6011, 214.9853, 202.1425, 
    199.9842,
  211.1423, 212.5664, 220.5835, 217.7019, 215.3212, 207.0127, 192.1306, 
    182.4206, 186.6092, 209.0929, 216.4063, 214.9421, 216.1402, 209.8509, 
    203.488,
  213.4397, 218.2731, 216.3437, 213.5824, 211.2128, 208.2319, 187.456, 
    177.4434, 180.9954, 198.2218, 217.9521, 216.5478, 217.1163, 216.4013, 
    209.375,
  215.4642, 214.1613, 213.1483, 212.4865, 209.235, 202.0688, 192.0331, 
    189.1853, 187.3302, 191.1449, 208.5233, 218.2323, 219.3495, 216.782, 
    214.3096,
  214.6111, 214.8374, 212.3195, 213.2235, 208.3005, 202.831, 192.3311, 
    187.0314, 182.9807, 186.547, 202.8702, 216.3342, 218.4983, 219.6666, 
    218.1938,
  216.137, 214.7159, 215.0295, 211.6078, 209.2274, 206.5789, 198.2464, 
    185.461, 183.4485, 188.131, 196.4595, 211.3002, 217.7232, 219.8739, 
    219.765,
  215.05, 214.4536, 214.8123, 210.9172, 209.3953, 208.0072, 205.143, 198.696, 
    193.7811, 189.7205, 192.4577, 205.55, 214.5454, 218.2478, 220.7663,
  216.0124, 217.6954, 218.8454, 211.2732, 209.1041, 212.4701, 212.9417, 
    208.6495, 195.1837, 194.1368, 194.5557, 201.8722, 212.2404, 217.7622, 
    217.7386,
  213.348, 215.9518, 223.1994, 212.8454, 211.6763, 217.0276, 214.1067, 
    213.0676, 208.6017, 201.4146, 197.4155, 202.2979, 207.1913, 208.2644, 
    215.78,
  196.2157, 199.4205, 210.2528, 214.4509, 213.8672, 209.9307, 211.9506, 
    211.5479, 201.0999, 213.8189, 213.9071, 214.2216, 211.2111, 196.3478, 
    188.2366,
  207.565, 209.2685, 218.754, 216.3595, 212.6576, 209.5142, 208.9899, 
    210.3822, 204.4332, 214.4599, 216.1358, 215.1712, 210.3808, 198.6733, 
    191.7217,
  218.5835, 215.4869, 217.4083, 210.886, 208.2714, 208.1452, 196.336, 
    187.2205, 195.6702, 213.9909, 216.2431, 215.3386, 214.2347, 205.6734, 
    190.7057,
  213.5159, 212.6613, 211.2553, 208.9409, 201.2016, 202.2299, 192.0778, 
    186.2434, 198.5907, 208.5878, 215.1411, 215.9507, 214.2709, 210.9501, 
    194.3628,
  212.6126, 211.5296, 210.2832, 208.3455, 202.2261, 199.9406, 200.1153, 
    203.8943, 206.4836, 209.361, 214.5524, 215.8726, 215.1664, 210.8083, 
    200.7159,
  219.7163, 215.0858, 211.4338, 209.4595, 205.7737, 203.1041, 203.3578, 
    203.7728, 201.0675, 205.6675, 213.4613, 214.5643, 216.3401, 210.4604, 
    204.5605,
  215.9014, 217.478, 212.4037, 212.0927, 211.0559, 208.6414, 207.9874, 
    206.6909, 203.6892, 204.458, 211.2326, 212.4583, 218.0647, 213.0264, 
    207.3051,
  215.1698, 220.5681, 223.4768, 216.167, 214.4625, 211.7286, 212.5063, 
    214.4386, 211.8092, 211.5629, 211.1154, 212.7946, 215.6575, 217.4991, 
    215.4267,
  210.9881, 216.758, 223.4097, 217.1986, 217.4516, 213.827, 213.2585, 
    211.9419, 212.0102, 212.3085, 213.7569, 212.6953, 211.8102, 219.0141, 
    219.1197,
  209.3247, 212.1507, 222.1614, 217.2276, 219.6219, 214.5995, 213.3206, 
    213.2823, 212.6062, 213.5008, 216.4608, 214.3952, 211.3873, 212.4298, 
    219.662,
  224.2022, 217.0697, 215.0303, 212.7811, 207.0125, 206.6946, 212.1039, 
    211.4654, 205.6642, 205.9758, 208.1892, 206.796, 208.4263, 209.2131, 
    206.4742,
  226.045, 219.8316, 215.8264, 208.2673, 207.357, 208.6471, 211.9363, 
    212.9409, 211.9349, 207.2056, 205.0787, 206.7276, 208.7455, 207.0184, 
    208.5802,
  214.7582, 212.362, 217.4061, 208.9323, 209.9493, 209.6177, 212.5828, 
    210.2796, 205.4619, 205.1398, 205.9806, 208.5667, 212.7528, 211.7029, 
    208.5358,
  213.9889, 212.7199, 215.6697, 213.2693, 212.1447, 213.8544, 212.6249, 
    212.9329, 210.9354, 204.6485, 205.3298, 209.491, 212.8763, 202.014, 
    200.7272,
  214.1872, 214.5111, 215.1732, 212.7019, 213.0164, 211.3512, 212.4316, 
    209.3743, 205.4886, 205.8624, 205.4847, 208.7379, 214.7069, 202.4986, 
    204.9829,
  212.4975, 213.1349, 215.9144, 213.615, 213.361, 210.7276, 210.0814, 
    211.5853, 210.0984, 206.7216, 205.6568, 207.3988, 209.4267, 203.0713, 
    209.3409,
  212.4052, 214.0043, 222.974, 219.5972, 213.6907, 211.41, 210.2505, 
    210.3854, 209.6939, 206.2025, 206.8994, 206.7585, 209.1839, 204.8557, 
    206.2234,
  211.5714, 213.0585, 230.6784, 218.3671, 213.9584, 211.7385, 209.8097, 
    210.447, 211.049, 211.0251, 205.994, 207.5888, 207.8156, 210.7612, 
    205.6174,
  215.9717, 228.7899, 225.9904, 217.2465, 215.217, 212.4594, 209.8193, 
    210.4095, 210.6, 213.1781, 208.3553, 206.3269, 208.4872, 208.9657, 
    205.3592,
  209.731, 224.2605, 224.3417, 218.0008, 214.3626, 213.1091, 212.751, 
    211.5953, 210.204, 213.5947, 212.5692, 206.9617, 206.6153, 206.7006, 
    208.502,
  223.037, 215.0178, 212.9115, 212.9526, 212.0383, 210.683, 213.1017, 
    213.5104, 214.1809, 207.822, 204.3129, 201.2019, 201.0188, 202.7301, 
    203.3392,
  218.5608, 213.1118, 214.3375, 212.845, 212.6364, 211.9973, 211.5217, 
    216.0548, 215.637, 210.5426, 203.8122, 203.3766, 205.5602, 205.8322, 
    203.3199,
  216.8422, 213.751, 217.0665, 212.169, 212.7775, 208.2226, 215.2076, 
    213.7611, 212.0429, 205.3562, 204.5035, 206.3031, 206.5546, 206.9769, 
    198.8756,
  214.2136, 222.5459, 213.414, 212.969, 211.3132, 212.1591, 209.1992, 
    214.9226, 215.2081, 209.0711, 207.3758, 204.5133, 206.7396, 206.4425, 
    203.4805,
  218.3648, 224.0584, 219.1056, 212.4417, 207.91, 206.5287, 209.0662, 
    208.3097, 207.1057, 211.7787, 207.1835, 207.3237, 206.1763, 214.3905, 
    209.9904,
  215.4926, 224.3323, 222.1235, 212.7329, 207.6615, 205.088, 207.7784, 
    209.8315, 210.7372, 210.7844, 207.9032, 204.338, 204.8314, 212.1427, 
    205.9135,
  211.2994, 220.4236, 224.5214, 212.5994, 204.0244, 203.8468, 207.3807, 
    209.3063, 210.0309, 210.2181, 209.009, 204.6421, 204.3287, 205.6712, 
    215.4712,
  211.2616, 215.0354, 224.2634, 211.5516, 204.5845, 202.6595, 207.6593, 
    209.9332, 211.8508, 210.6221, 210.9691, 206.1843, 204.6785, 217.632, 
    220.8721,
  221.7443, 217.6488, 221.3371, 211.651, 204.3263, 205.1318, 209.9684, 
    209.4133, 211.9019, 213.0734, 211.1704, 209.8037, 206.0469, 219.7171, 
    224.1393,
  218.1155, 221.9149, 210.4233, 209.1394, 205.6104, 205.0342, 207.083, 
    210.2985, 212.1243, 213.7125, 211.8126, 211.6749, 212.2554, 219.6775, 
    221.7265,
  219.7935, 216.4931, 213.7242, 211.06, 209.3122, 207.5599, 206.6559, 
    211.5535, 214.1663, 209.5216, 207.563, 206.9501, 205.573, 205.1104, 
    205.9405,
  220.5802, 214.6479, 213.2159, 209.3116, 208.587, 209.1109, 205.576, 
    210.3263, 211.751, 211.0307, 208.4582, 208.1669, 207.5431, 202.2921, 
    212.3297,
  217.8313, 215.0996, 211.5544, 207.3627, 209.2477, 205.7445, 208.2616, 
    206.6222, 208.1767, 206.7077, 209.098, 206.8116, 204.4963, 203.0217, 
    211.8988,
  222.7907, 215.1099, 208.825, 202.1018, 199.8162, 203.8226, 204.776, 
    206.2338, 203.518, 207.435, 206.4073, 205.6098, 204.6634, 208.2945, 
    212.8286,
  211.5952, 210.9055, 208.3046, 202.1078, 196.962, 198.5471, 201.4013, 
    203.8329, 204.7012, 203.8992, 202.4842, 206.2953, 205.0527, 210.6782, 
    214.0897,
  203.9326, 200.9796, 204.103, 194.4538, 199.1216, 199.3431, 193.9128, 
    198.7809, 201.0845, 196.4387, 200.5128, 204.2256, 205.3964, 217.646, 
    216.1028,
  202.6852, 201.47, 200.595, 202.5873, 201.8895, 200.4232, 197.4003, 
    195.2316, 195.1262, 199.9526, 205.6207, 208.2247, 205.0337, 218.9202, 
    217.0728,
  200.8461, 196.103, 202.2093, 206.0337, 204.0217, 201.6631, 198.5119, 
    198.6699, 198.669, 201.1568, 206.2016, 208.7227, 205.7131, 217.2402, 
    218.0671,
  204.2456, 202.4755, 204.8738, 210.2456, 204.5755, 201.8001, 201.7126, 
    195.7019, 199.3084, 207.8857, 212.133, 211.4362, 215.2668, 218.4953, 
    218.7119,
  206.1239, 207.9067, 211.1269, 209.2946, 206.9813, 205.6031, 200.4088, 
    200.9664, 207.106, 213.7715, 213.9285, 211.813, 218.731, 217.5963, 
    215.7759,
  207.316, 209.7947, 204.4276, 199.3297, 193.6793, 190.7424, 193.6785, 
    195.5197, 191.5431, 196.0655, 202.7892, 206.3157, 207.6167, 208.4638, 
    207.237,
  211.6786, 207.0979, 202.9177, 198.4126, 196.8125, 193.0588, 191.2307, 
    192.0744, 193.9429, 187.0909, 200.1791, 206.6896, 208.6027, 209.5209, 
    210.4777,
  207.8229, 201.156, 200.5137, 197.8471, 194.8683, 195.2773, 192.9464, 
    187.5574, 189.6376, 195.0438, 195.4272, 202.5664, 208.0457, 209.324, 
    211.005,
  209.4027, 204.0332, 201.0862, 197.9585, 199.8032, 200.6465, 197.6366, 
    200.6728, 198.6177, 194.5804, 195.8869, 201.6506, 210.0516, 208.7363, 
    210.8163,
  213.5228, 213.0552, 207.2742, 204.6888, 207.368, 206.1131, 204.9176, 
    204.4799, 208.3794, 208.263, 201.3228, 199.2566, 205.1654, 210.0856, 
    210.7788,
  220.6868, 219.4373, 209.2748, 210.5272, 210.8587, 208.6406, 206.4704, 
    206.3734, 213.5801, 209.387, 212.4053, 206.2499, 207.0409, 210.7639, 
    211.5691,
  221.5443, 219.9509, 215.4996, 211.2072, 212.6826, 211.9238, 214.5089, 
    211.2385, 210.5826, 219.0371, 214.0726, 211.4408, 210.8284, 215.4806, 
    213.1611,
  221.3711, 215.4007, 212.9946, 208.9791, 211.2205, 210.592, 213.6313, 
    214.2648, 214.5532, 218.549, 216.4275, 214.2784, 213.5445, 212.9572, 
    212.0838,
  221.1497, 219.1812, 212.8386, 210.188, 208.3785, 209.4292, 209.1241, 
    213.4736, 215.0046, 219.6732, 213.1584, 217.0598, 215.5152, 211.4998, 
    213.6344,
  224.3634, 213.6673, 214.7446, 213.976, 209.3692, 208.6041, 209.2414, 
    210.5347, 209.1082, 212.2898, 215.3201, 215.8908, 213.3771, 209.9439, 
    214.21,
  228.163, 223.7619, 219.8671, 218.1709, 215.3826, 215.4223, 213.7385, 
    207.213, 204.2332, 201.2055, 194.4662, 189.7794, 196.3265, 202.3045, 
    207.237,
  216.969, 222.2623, 218.0078, 216.1627, 215.7844, 214.5651, 208.8049, 
    210.9438, 207.8828, 198.9349, 194.364, 187.8676, 194.6696, 201.0748, 
    208.1144,
  221.289, 221.868, 218.4788, 213.5304, 214.6245, 207.2484, 207.4129, 
    207.9564, 210.7764, 207.2489, 196.8536, 190.3426, 193.0768, 202.2883, 
    209.5919,
  221.2017, 219.8799, 219.5337, 208.4226, 203.3825, 200.3031, 201.0706, 
    201.0883, 210.5381, 211.8722, 206.4988, 193.4164, 190.7484, 202.4572, 
    210.907,
  220.1007, 222.615, 219.7715, 208.2486, 203.3638, 197.1732, 199.6615, 
    201.7377, 206.5829, 214.1169, 209.0822, 201.1149, 192.7731, 202.1336, 
    211.5928,
  219.2858, 222.776, 211.4922, 202.4949, 202.6719, 200.2001, 197.3168, 
    200.6131, 203.9207, 209.5309, 213.3633, 206.7827, 200.6213, 212.3189, 
    213.6341,
  224.3351, 228.96, 216.7956, 203.3293, 208.3043, 206.4184, 204.9052, 
    200.841, 202.5047, 210.3928, 215.8454, 211.3881, 210.1291, 214.8932, 
    212.6279,
  224.8806, 223.8548, 216.0774, 207.818, 211.3395, 208.5604, 210.9872, 
    210.7014, 206.8775, 207.6837, 215.9495, 215.3462, 215.0561, 217.3015, 
    210.1821,
  229.1772, 222.578, 214.3955, 214.5207, 212.3458, 213.0423, 215.8699, 
    212.8839, 206.6462, 212.1745, 217.5705, 218.3142, 217.0089, 215.8069, 
    208.1368,
  220.6609, 222.7039, 220.387, 217.3416, 215.7116, 216.0781, 217.464, 
    214.6658, 215.1888, 212.5834, 218.0074, 218.1038, 218.015, 215.5262, 
    210.503,
  211.2481, 207.1433, 211.5451, 209.5107, 205.9095, 211.1144, 210.1912, 
    205.0762, 204.2335, 203.7222, 211.2577, 218.3, 212.156, 204.0822, 199.3422,
  218.8948, 216.8476, 211.1788, 207.3802, 204.4419, 210.4356, 206.6609, 
    204.4505, 201.233, 199.7563, 204.3996, 216.8824, 215.1242, 207.9992, 
    201.6625,
  226.4949, 227.7256, 222.2908, 208.4865, 206.2431, 208.7765, 209.3674, 
    200.2409, 201.3909, 199.1088, 203.788, 212.2643, 213.6926, 205.9067, 
    204.8532,
  235.7563, 228.6491, 228.3249, 222.0111, 212.0638, 212.767, 205.7515, 
    206.0341, 204.6784, 202.3847, 207.7566, 214.4346, 213.1252, 208.8429, 
    206.7551,
  233.9359, 232.2256, 221.5985, 221.8222, 215.2261, 213.75, 215.1533, 
    208.3967, 209.2542, 202.2829, 202.7164, 214.716, 214.0012, 207.8091, 
    208.5286,
  235.8354, 232.9117, 231.6117, 209.1195, 214.6173, 216.761, 215.4538, 
    208.5442, 205.3228, 196.8642, 201.2636, 212.8902, 212.11, 209.6544, 
    209.4944,
  234, 233.1147, 228.3883, 214.7649, 214.4272, 217.7071, 216.5067, 207.6446, 
    201.4438, 203.1513, 206.2836, 214.4158, 214.6634, 214.5166, 208.6644,
  229.8629, 230.032, 219.123, 209.0902, 211.1698, 219.008, 214.3171, 
    211.2468, 208.9812, 203.7362, 207.0816, 214.9002, 216.3704, 215.5912, 
    207.5905,
  234.1893, 226.8762, 217.8045, 213.5324, 199.6167, 218.0968, 211.4614, 
    202.5513, 199.8104, 204.581, 214.8756, 216.2709, 214.8952, 209.2616, 
    211.5804,
  232.558, 228.4198, 223.2227, 216.6477, 209.1044, 214.6432, 210.9713, 
    205.1799, 207.8359, 212.1572, 216.5564, 215.3609, 214.1419, 211.4969, 
    208.2373,
  212.5695, 219.7421, 225.518, 229.7187, 223.7138, 219.4532, 212.4679, 
    210.1175, 214.1785, 215.004, 220.9123, 220.2618, 215.5354, 199.4207, 
    190.5981,
  217.7509, 228.1948, 229.2737, 228.6412, 221.2758, 212.2244, 204.0992, 
    209.6618, 211.7582, 213.9164, 215.2931, 220.7169, 211.6562, 200.9314, 
    189.8644,
  238.162, 237.4924, 234.508, 224.1973, 217.1513, 208.9452, 197.3958, 
    206.1822, 212.3657, 209.39, 211.0719, 217.1942, 210.6842, 199.8513, 
    190.7231,
  235.404, 237.3886, 231.4595, 226.279, 215.694, 213.7038, 196.1227, 
    207.2105, 211.5748, 205.7327, 207.8337, 210.1533, 212.4816, 200.7851, 
    197.9568,
  238.2542, 234.6064, 233.1114, 227.7737, 221.2942, 213.5035, 205.4901, 
    197.8547, 208.9217, 205.9143, 206.6445, 211.6341, 208.8594, 205.9336, 
    203.6784,
  234.8663, 233.2114, 230.4946, 217.8773, 214.0678, 214.6123, 210.2767, 
    198.7276, 204.9754, 210.8624, 210.5428, 209.5601, 206.896, 207.8838, 
    207.2945,
  235.574, 235.9308, 230.8619, 215.4472, 214.2468, 211.2916, 218.1086, 
    199.3482, 205.9832, 213.3548, 205.9422, 210.6038, 208.5642, 208.7299, 
    205.3992,
  235.2131, 228.0023, 213.0514, 211.623, 217.1305, 211.5848, 215.1444, 
    204.5953, 211.8817, 216.3346, 208.8786, 208.8521, 212.9266, 210.4088, 
    205.4365,
  229.9277, 225.7198, 223.8508, 210.9392, 214.3094, 210.0029, 205.8545, 
    201.5981, 208.1699, 215.1829, 208.4784, 210.2333, 215.2056, 212.1291, 
    205.1501,
  226.6371, 221.9119, 218.5688, 215.1913, 214.0703, 208.329, 205.6582, 
    206.1157, 213.5944, 215.1478, 209.5141, 210.3571, 214.6356, 210.3859, 
    208.2981,
  225.0866, 216.9262, 218.09, 227.7016, 226.046, 223.9503, 221.9786, 
    213.3997, 208.6301, 204.4868, 216.1064, 224.8701, 223.7198, 217.4907, 
    209.2862,
  225.8957, 231.3658, 229.6155, 230.1043, 223.7142, 221.131, 216.8322, 
    215.7252, 209.2518, 208.7516, 209.9297, 218.4304, 220.7165, 206.5349, 
    201.0858,
  237.8144, 236.4557, 233.9809, 228.0373, 217.5861, 224.4266, 219.4643, 
    211.5553, 211.6299, 220.6462, 218.7814, 221.5289, 211.8167, 197.8187, 
    193.6013,
  238.6414, 236.3002, 229.5206, 223.661, 216.9468, 218.5693, 214.0423, 
    216.1359, 221.6223, 217.5429, 218.0194, 215.8521, 201.7453, 190.3776, 
    192.4788,
  235.0188, 234.038, 224.5334, 225.913, 216.8543, 210.689, 216.8932, 
    211.0024, 216.6587, 211.1721, 213.04, 205.3427, 189.4746, 188.6588, 
    187.1657,
  233.7581, 232.5193, 232.2119, 225.8887, 215.5888, 215.7229, 214.5012, 
    212.8205, 205.3274, 206.2325, 205.2136, 191.8444, 184.0354, 189.7784, 
    190.4256,
  234.9272, 233.345, 228.7811, 218.9635, 215.8298, 215.5962, 210.0077, 
    209.1453, 201.6459, 202.1578, 192.2809, 188.1146, 182.9648, 186.2234, 
    193.2228,
  231.7224, 230.4512, 209.3414, 219.3763, 214.4621, 211.2073, 207.3579, 
    198.9965, 201.2423, 195.1769, 186.7571, 185.3038, 182.9054, 186.2818, 
    192.6018,
  226.5239, 226.2916, 219.5172, 214.118, 214.1541, 213.081, 200.4678, 
    196.2159, 197.7272, 194.7894, 186.628, 182.8728, 188.307, 188.1506, 
    203.1618,
  225.6515, 225.2392, 221.694, 218.4246, 211.7294, 197.5392, 193.5388, 
    193.9182, 197.667, 191.9845, 189.1278, 188.575, 188.1601, 194.3304, 
    205.1772,
  198.5818, 199.4535, 199.4445, 204.6595, 204.9679, 205.7401, 210.1337, 
    213.4252, 213.7738, 217.3971, 220.2371, 217.9346, 217.3262, 218.6717, 
    217.6244,
  203.2925, 205.692, 206.9702, 213.149, 218.8866, 219.2503, 213.2168, 
    215.6978, 217.8894, 215.7687, 218.3138, 211.58, 209.5369, 217.5184, 
    220.2473,
  214.9951, 226.5777, 234.8065, 230.4368, 222.8588, 218.9368, 222.1124, 
    212.4531, 218.753, 220.2439, 217.9069, 212.8602, 219.1443, 221.6384, 
    222.1774,
  241.3406, 236.0667, 236.1747, 231.4216, 224.4767, 223.4677, 216.9579, 
    219.7161, 221.3241, 220.6831, 220.9982, 218.3048, 222.038, 222.5777, 
    219.8766,
  240.2574, 237.8281, 234.0608, 231.0699, 222.6828, 214.1662, 216.4684, 
    214.0467, 215.2635, 222.6529, 223.2338, 223.909, 223.3152, 220.2619, 
    213.487,
  238.752, 234.2122, 230.8713, 227.5982, 218.7595, 215.3232, 212.8648, 
    219.135, 218.9083, 222.2204, 223.0905, 222.3448, 217.0364, 213.6635, 
    204.4164,
  238.7999, 237.6502, 213.3151, 220.3807, 218.5928, 214.8025, 216.1408, 
    221.9441, 220.4107, 220.2265, 218.4393, 212.0207, 208.1512, 205.9273, 
    200.3329,
  238.2474, 234.1961, 214.3372, 219.3093, 216.394, 218.3885, 218.7665, 
    218.511, 216.7672, 209.7567, 207.9309, 203.9929, 201.8003, 204.2004, 
    207.3892,
  232.6276, 228.1061, 222.9386, 211.7939, 204.4367, 204.0617, 205.9434, 
    207.3038, 205.1047, 203.3992, 198.8888, 200.9865, 200.6856, 209.2849, 
    217.4491,
  227.8426, 228.0059, 214.9859, 200.5283, 198.1785, 196.6019, 196.8553, 
    200.7732, 196.6228, 197.2652, 193.1384, 199.4666, 207.209, 215.3352, 
    221.3738,
  211.0041, 215.1125, 214.723, 212.4152, 213.6503, 218.8347, 218.6894, 
    214.232, 211.7363, 214.1539, 210.5261, 209.816, 207.7708, 204.81, 205.1295,
  205.2113, 209.3939, 207.8157, 208.267, 208.8583, 213.579, 213.6861, 
    211.4963, 211.734, 212.1633, 212.3531, 212.9538, 214.6157, 209.7497, 
    211.6445,
  197.8654, 198.8638, 199.4585, 205.1395, 210.808, 213.047, 215.9223, 
    212.8237, 216.1918, 213.3446, 214.5115, 209.6569, 211.2321, 215.167, 
    217.9414,
  190.272, 189.0147, 198.0498, 207.1691, 209.9631, 213.8486, 211.8955, 
    218.4715, 220.7319, 218.0138, 208.8933, 212.0329, 209.3621, 217.9489, 
    215.0079,
  197.188, 205.4528, 213.717, 220.1078, 217.6106, 213.1118, 216.5845, 
    211.5357, 210.8194, 214.9223, 214.4998, 215.4389, 214.0985, 217.7203, 
    219.8879,
  210.9476, 223.7094, 229.3097, 228.3599, 223.7901, 215.6615, 210.6606, 
    214.3161, 215.8788, 213.816, 217.0736, 215.9182, 217.2719, 218.6898, 
    215.8359,
  225.9382, 236.558, 236.4209, 224.0655, 219.1909, 212.1131, 211.7257, 
    209.9121, 213.0345, 221.1064, 215.7789, 212.5575, 213.7672, 219.7795, 
    217.6836,
  238.6289, 239.8914, 232.2345, 223.2561, 214.7477, 214.0352, 219.861, 
    224.1332, 222.7376, 220.8682, 220.0655, 216.6005, 213.4707, 216.6702, 
    215.8206,
  229.3635, 234.0035, 227.7668, 217.8601, 214.4596, 222.8991, 225.8064, 
    225.1497, 222.7309, 220.3339, 220.1337, 218.8023, 214.5488, 213.5363, 
    211.9077,
  222.1114, 230.6321, 220.9616, 215.9385, 221.7896, 227.6839, 227.4009, 
    225.8825, 221.2826, 216.0051, 220.1157, 213.146, 210.2724, 211.1239, 
    210.2942,
  222.0731, 223.0637, 222.1822, 226.7214, 220.7724, 223.4543, 211.3113, 
    199.147, 190.1516, 189.3971, 189.0133, 193.7132, 199.8348, 206.8716, 
    214.0725,
  214.3421, 216.9222, 223.443, 223.1955, 220.7172, 214.5028, 205.3333, 
    198.4571, 191.7567, 194.0879, 193.6264, 197.9292, 207.724, 209.1894, 
    212.4088,
  216.2565, 218.1571, 216.4139, 212.2841, 206.4727, 199.2342, 198.42, 
    191.6404, 193.9168, 196.3484, 198.7849, 206.7669, 209.1385, 215.316, 
    210.5942,
  212.9706, 213.8121, 206.0988, 203.2252, 194.2648, 193.6432, 189.3434, 
    194.3247, 194.2243, 202.072, 208.8757, 213.2673, 211.8521, 214.3781, 
    215.5434,
  225.4324, 209.4492, 205.1291, 193.838, 188.5306, 187.8535, 197.5581, 
    200.0213, 205.0357, 214.8129, 221.4729, 216.0879, 217.7319, 218.966, 
    220.2243,
  205.015, 196.9086, 191.1211, 190.2399, 191.939, 197.8336, 208.5761, 
    221.4567, 224.4263, 223.7997, 223.9862, 223.3705, 218.266, 218.5153, 
    216.9231,
  188.3185, 186.0518, 190.7013, 193.4623, 205.5201, 221.4278, 227.8981, 
    227.6125, 224.7054, 220.3469, 213.7431, 216.6776, 218.3475, 216.436, 
    217.4565,
  186.3064, 194.3729, 198.9139, 211.0256, 226.2996, 223.2341, 227.2909, 
    225.5352, 224.2663, 221.32, 220.4718, 219.3693, 219.762, 219.35, 213.2854,
  189.8851, 196.3016, 215.2556, 222.5934, 222.3289, 226.4389, 224.3979, 
    221.2502, 220.1165, 215.9955, 217.1388, 209.6625, 209.8579, 213.1699, 
    214.4704,
  196.9375, 210.6537, 217.9607, 225.025, 226.5114, 223.4388, 220.9536, 
    219.5308, 218.5926, 218.9305, 218.9712, 211.8275, 212.2799, 216.3695, 
    211.9323,
  239.583, 240.9814, 232.1663, 226.6982, 220.7078, 218.321, 220.7472, 
    221.4798, 218.5379, 219.7009, 217.3344, 215.1808, 214.6494, 212.4756, 
    208.9075,
  238.0891, 231.7826, 218.2886, 211.7831, 210.1019, 204.4226, 203.8256, 
    204.4866, 208.8999, 210.7814, 215.8965, 214.0794, 215.6675, 210.9485, 
    209.5656,
  232.9347, 220.9759, 211.067, 206.4774, 204.5729, 201.2241, 202.3795, 
    203.2028, 204.9898, 207.2632, 209.0526, 208.8824, 211.815, 210.1067, 
    208.4245,
  229.4143, 219.207, 204.8191, 204.7791, 204.0461, 206.4382, 201.4924, 
    203.0791, 199.122, 202.6645, 214.2892, 219.8453, 212.388, 202.0043, 
    201.5336,
  221.6393, 209.2194, 201.7382, 205.2874, 205.2954, 208.5147, 209.6004, 
    205.6748, 212.853, 213.7621, 208.961, 209.1488, 205.0914, 205.582, 
    205.4238,
  212.5311, 195.7263, 202.2771, 205.4727, 208.1357, 206.6543, 211.8932, 
    216.135, 220.7355, 217.2187, 214.8682, 209.3407, 208.4235, 207.8171, 
    207.0221,
  197.2172, 194.4457, 199.9277, 203.9722, 213.9184, 221.7914, 227.024, 
    228.941, 227.7281, 218.3741, 213.9945, 208.6626, 208.01, 207.032, 207.8856,
  189.2079, 196.887, 204.4931, 215.9218, 224.1335, 227.7044, 228.5807, 
    228.5827, 227.8039, 226.2011, 222.7621, 215.8385, 214.2863, 212.9105, 
    212.7821,
  193.8278, 204.0937, 213.0159, 216.4493, 217.8655, 217.7227, 223.1002, 
    223.9275, 223.7586, 222.8101, 221.2495, 219.7973, 217.4764, 218.7453, 
    213.934,
  200.4527, 213.5346, 218.738, 217.37, 216.7138, 215.1113, 216.0496, 
    224.0653, 222.4626, 221.8518, 219.8675, 213.7913, 214.7935, 215.4741, 
    213.2564,
  192.2632, 199.6097, 204.2118, 206.9935, 212.3779, 212.6634, 218.2812, 
    223.449, 222.8922, 219.5968, 217.1295, 216.958, 215.7059, 214.4248, 
    219.3409,
  207.4669, 213.0331, 215.6661, 215.8018, 222.2014, 218.088, 220.8842, 
    221.3464, 219.4068, 216.7935, 215.5365, 211.9586, 209.7153, 208.968, 
    205.4491,
  215.1318, 218.0888, 216.0267, 216.9159, 222.1776, 216.2337, 220.798, 
    224.4591, 222.8175, 223.0934, 220.1383, 216.5042, 210.222, 208.1324, 
    202.8758,
  222.4617, 219.5805, 218.6223, 219.1794, 218.2465, 224.4974, 217.2017, 
    226.789, 226.8401, 223.5374, 224.8038, 220.1367, 213.3015, 209.1939, 
    200.1295,
  212.884, 208.2157, 214.1752, 216.5359, 218.056, 222.2466, 220.9613, 
    219.6197, 217.1853, 224.9368, 224.2143, 223.3469, 212.4997, 211.4682, 
    203.2456,
  205.7159, 202.7924, 208.5292, 221.5565, 222.3524, 223.6889, 219.6283, 
    223.862, 225.2324, 226.7644, 225.2128, 214.4657, 206.1467, 203.106, 
    200.455,
  207.3617, 206.4875, 211.136, 214.6031, 221.6796, 220.9933, 222.2104, 
    222.7068, 224.549, 225.8874, 226.2092, 201.1325, 200.7298, 198.1329, 
    199.7361,
  216.6571, 215.1249, 215.5536, 212.8004, 212.9808, 212.6979, 221.1189, 
    223.2072, 224.9032, 225.3307, 221.8698, 199.6447, 198.0999, 196.6084, 
    199.9774,
  227.4684, 215.0289, 213.3013, 211.3328, 209.39, 210.822, 219.2466, 
    223.1906, 223.9727, 224.0284, 220.2872, 199.9114, 195.6517, 196.1228, 
    198.5151,
  212.0807, 217.0078, 210.9057, 209.4094, 210.6501, 212.7656, 214.45, 
    223.2598, 223.8696, 223.4114, 217.6195, 200.9137, 199.6899, 203.6006, 
    209.3575,
  240.4457, 235.9328, 233.8991, 226.7637, 219.2782, 213.5451, 212.8415, 
    210.7612, 204.2511, 201.4448, 208.9937, 212.2206, 219.4067, 219.0872, 
    223.6749,
  235.4531, 232.9631, 232.1729, 226.5804, 218.7306, 215.6202, 215.1177, 
    207.4467, 200.0753, 196.8956, 205.4597, 212.6769, 219.8919, 221.92, 
    222.8052,
  229.662, 229.2913, 225.9825, 220.359, 217.1777, 210.1755, 207.843, 
    197.8113, 192.1469, 195.1385, 208.134, 217.0483, 224.8977, 223.9298, 
    221.9556,
  224.674, 218.7701, 217.5324, 216.064, 206.9325, 200.5931, 193.8322, 
    193.322, 193.6083, 201.8421, 208.6144, 219.7953, 226.2486, 224.5429, 
    214.2851,
  219.2643, 213.8822, 211.8801, 204.4863, 204.946, 194.5538, 195.4158, 
    196.1398, 195.8335, 209.0358, 216.2815, 223.7648, 226.5791, 215.652, 
    205.1192,
  219.9347, 212.345, 209.4993, 207.8048, 208.6965, 204.8164, 198.17, 201.541, 
    205.7977, 210.1325, 218.7294, 227.8684, 218.0564, 205.1866, 205.4604,
  224.7894, 216.5288, 209.2365, 213.7065, 210.1904, 206.14, 207.3984, 
    207.4622, 209.852, 217.5434, 226.3554, 222.2331, 215.0557, 201.52, 
    204.8674,
  229.8076, 216.3709, 214.5057, 213.2731, 213.0191, 213.7628, 216.4154, 
    221.3781, 221.4958, 226.0279, 227.2896, 218.9399, 207.5572, 198.5019, 
    204.7739,
  236.6472, 223.1279, 214.2779, 210.9723, 211.295, 211.6384, 214.4206, 
    222.2864, 223.841, 226.1396, 215.7845, 209.8311, 198.0552, 196.3316, 
    207.7278,
  230.2661, 219.1377, 211.3073, 214.3971, 214.6891, 220.4655, 221.5174, 
    223.5888, 225.2531, 222.049, 212.5276, 207.8285, 208.9349, 213.9078, 
    216.1398,
  226.455, 223.7621, 224.1277, 224.5548, 226.8165, 220.4225, 210.6919, 
    210.424, 208.9924, 214.383, 216.0986, 204.6591, 192.9572, 189.2671, 
    188.367,
  216.7503, 220.3624, 224.2834, 226.5397, 226.0937, 221.6906, 207.5337, 
    207.3108, 208.4995, 204.3306, 196.409, 189.6473, 190.8267, 188.4646, 
    202.261,
  219.7033, 221.0541, 223.0823, 227.7842, 223.8831, 217.3424, 206.3095, 
    194.4423, 193.4865, 194.3182, 190.2369, 190.8112, 197.8022, 212.0722, 
    229.2041,
  222.1355, 223.5345, 229.5964, 226.3389, 220.5065, 224.066, 197.6353, 
    190.1848, 189.2164, 187.4866, 189.4878, 199.156, 218.5795, 228.459, 
    225.9783,
  230.7126, 226.4826, 235.6084, 222.4415, 219.2988, 214.781, 200.6021, 
    184.8239, 182.0161, 187.1562, 192.1244, 208.223, 224.1435, 225.6683, 
    218.2727,
  241.0979, 224.2644, 222.6034, 218.1281, 216.1895, 215.8382, 207.4493, 
    187.6015, 180.0185, 185.6359, 190.1472, 216.1411, 224.7434, 225.8251, 
    223.7148,
  238.9707, 223.2717, 216.1366, 212.5675, 214.3426, 215.5111, 216.4364, 
    191.5936, 183.7115, 190.814, 202.5434, 220.6899, 224.5458, 222.0512, 
    220.8077,
  240.8967, 221.4279, 214.4814, 210.3796, 210.2324, 212.6087, 216.1009, 
    216.9514, 200.8337, 202.7896, 214.1307, 216.1945, 213.8785, 212.2603, 
    209.5013,
  235.1634, 224.4166, 217.2398, 210.9602, 210.261, 212.0721, 215.1708, 
    224.4232, 217.4882, 212.6871, 218.6636, 213.0975, 213.894, 213.3175, 
    212.6868,
  228.1866, 225.7275, 215.7336, 214.2132, 210.3295, 216.2896, 219.0868, 
    224.9969, 219.8671, 219.1545, 210.8512, 214.4246, 216.2128, 216.4776, 
    219.6658,
  205.3354, 204.8205, 209.4098, 222.996, 228.9578, 229.4076, 225.6271, 
    220.9524, 211.9654, 211.2488, 217.0205, 217.229, 219.5693, 217.5023, 
    204.7886,
  205.4658, 211.5223, 221.1691, 227.8409, 232.4546, 229.3594, 224.6545, 
    221.0524, 213.3839, 209.5108, 215.2376, 216.0513, 220.3429, 219.4498, 
    220.0364,
  211.1997, 221.0112, 229.5426, 232.7094, 230.5896, 228.6913, 224.675, 
    214.9996, 208.0366, 200.6371, 208.5707, 212.0871, 215.4471, 216.8276, 
    217.1167,
  218.1727, 232.3627, 234.3568, 229.8445, 227.4299, 229.9739, 219.9677, 
    216.9938, 206.9393, 199.5299, 207.2362, 209.5184, 212.007, 214.7498, 
    216.5658,
  233.7107, 240.9121, 231.6652, 226.817, 223.6925, 215.5186, 217.57, 
    214.5094, 201.2138, 200.9044, 207.158, 206.6002, 207.3752, 211.5674, 
    214.4332,
  244.3594, 235.7626, 231.6442, 219.3754, 206.5949, 207.6926, 210.348, 
    215.8182, 203.3574, 200.5443, 210.6718, 206.5556, 205.1105, 205.3737, 
    211.5316,
  230.6675, 225.8064, 220.9777, 212.1679, 206.9401, 201.2314, 208.8027, 
    213.6882, 206.6165, 207.2459, 212.4193, 205.6018, 204.056, 203.1955, 
    204.8997,
  244.3157, 239.0143, 230.3249, 224.0439, 215.0963, 213.1403, 212.6331, 
    215.8842, 204.2386, 210.3732, 210.5877, 205.8736, 207.1466, 209.2217, 
    205.2655,
  238.4354, 231.5023, 230.2888, 228.5063, 218.8556, 216.9601, 212.9727, 
    217.7413, 202.3941, 212.8118, 207.2892, 207.844, 206.9593, 207.2349, 
    208.5753,
  234.2861, 228.6725, 228.2104, 227.6684, 227.8868, 219.8043, 215.7671, 
    215.7143, 205.9769, 213.0565, 207.8581, 209.3532, 206.9574, 209.0771, 
    208.6772,
  189.0663, 187.7963, 190.6548, 207.8731, 223.952, 230.1846, 227.865, 
    226.8217, 226.8935, 217.0555, 206.6003, 207.6149, 216.7972, 216.7038, 
    218.3084,
  185.8498, 191.2254, 204.2708, 224.7363, 231.9134, 231.3018, 227.1691, 
    226.1952, 224.5117, 219.4964, 207.065, 209.4756, 218.0284, 217.6447, 
    220.438,
  188.8398, 204.5898, 228.0796, 234.1432, 234.1981, 231.3235, 228.3302, 
    222.4405, 223.0219, 217.7483, 210.1935, 207.5295, 216.0989, 218.971, 
    220.48,
  200.392, 226.514, 238.2897, 238.8881, 232.1096, 232.6681, 220.7524, 
    226.2133, 222.749, 214.3093, 210.0949, 206.1535, 210.8516, 217.0957, 
    217.7695,
  216.5974, 222.1222, 226.6511, 229.0008, 231.7587, 218.0866, 216.3886, 
    216.8223, 214.6785, 217.663, 212.2597, 208.8247, 207.3918, 212.553, 
    213.9301,
  220.6331, 236.6494, 237.1842, 222.7778, 221.4142, 214.7813, 218.7778, 
    219.9398, 219.178, 214.8897, 212.9588, 211.4683, 208.3341, 210.0147, 
    209.0125,
  226.9085, 232.2406, 231.7686, 229.2781, 225.7495, 220.9447, 217.7051, 
    219.7355, 219.8006, 217.8076, 215.1718, 211.7102, 208.1539, 208.4334, 
    209.7989,
  233.0779, 230.4257, 228.1345, 224.9982, 220.6733, 220.9524, 220.3749, 
    222.3723, 216.8952, 215.6545, 210.0126, 208.4455, 208.0343, 208.034, 
    208.9177,
  230.7591, 229.7335, 224.8817, 222.6496, 220.3637, 219.3743, 222.2731, 
    220.6942, 216.6858, 212.2426, 208.6194, 205.8773, 203.7523, 210.3128, 
    206.6286,
  228.0977, 226.3445, 225.2802, 221.568, 220.4291, 220.9762, 218.6628, 
    218.5581, 216.7603, 213.0732, 207.8752, 200.8416, 202.149, 209.0389, 
    210.5874,
  236.2702, 231.6741, 228.8562, 229.3549, 229.6035, 230.8561, 227.9542, 
    225.2523, 222.5036, 219.241, 217.4719, 215.6816, 209.9411, 203.5383, 
    203.474,
  231.0381, 228.3839, 229.5871, 228.881, 231.1015, 228.3773, 225.2018, 
    224.0764, 223.3584, 218.3154, 215.9084, 208.4789, 206.5434, 206.4031, 
    207.0399,
  221.9149, 225.7595, 228.572, 228.558, 230.547, 223.941, 224.8536, 220.9946, 
    217.6937, 216.3658, 210.5712, 202.7602, 202.3805, 207.1345, 206.7608,
  218.1989, 224.7915, 226.5567, 229.4388, 225.0952, 223.9693, 220.0705, 
    224.2037, 218.53, 214.458, 212.2202, 201.3894, 207.8869, 209.289, 205.6318,
  215.375, 221.0231, 224.9027, 230.4999, 225.0543, 221.0771, 220.12, 
    218.1842, 216.9114, 216.2475, 210.7615, 205.6417, 203.1191, 206.5906, 
    205.7374,
  216.1411, 224.7542, 227.1121, 226.0898, 222.3361, 219.7684, 217.6167, 
    217.9378, 218.1969, 213.9035, 210.1515, 205.9918, 205.7131, 211.2835, 
    203.739,
  226.9671, 228.1846, 225.9206, 223.0214, 219.8855, 219.0339, 215.9575, 
    216.1938, 216.9563, 214.7961, 208.9658, 207.1667, 208.9569, 208.8921, 
    206.744,
  228.9657, 227.2202, 225.4281, 222.1926, 218.3553, 216.5654, 215.1459, 
    218.8732, 217.4189, 216.0653, 210.3478, 209.6624, 213.2852, 213.1415, 
    208.7056,
  227.6605, 225.1839, 226.4165, 221.2732, 217.0484, 215.5524, 218.4494, 
    219.3187, 218.7952, 216.3326, 213.6326, 210.9542, 210.0257, 212.3222, 
    213.337,
  225.9254, 228.3143, 225.1857, 220.7538, 217.2746, 216.6169, 216.0199, 
    217.8725, 219.3579, 219.3956, 215.4208, 214.8285, 213.8919, 210.0605, 
    208.0416,
  231.5619, 225.778, 229.9298, 229.8941, 227.81, 225.7989, 223.0863, 
    220.3149, 216.144, 213.9912, 211.4413, 211.0699, 211.0294, 205.5719, 
    204.2776,
  227.9218, 227.351, 229.5474, 227.321, 226.4352, 224.8017, 220.1498, 
    220.3858, 215.6277, 213.5964, 211.9162, 213.0313, 209.3006, 205.9993, 
    206.3805,
  226.8252, 227.9652, 228.3152, 226.5557, 226.9439, 220.381, 220.7993, 
    212.7015, 215.1843, 213.7492, 212.6675, 211.5967, 209.5078, 206.1443, 
    206.4711,
  227.6431, 228.4005, 228.4767, 227.0081, 222.9065, 221.1246, 217.0004, 
    214.2162, 216.9812, 213.5777, 212.0457, 212.3191, 208.3949, 205.3803, 
    204.0422,
  230.9759, 230.0893, 229.0965, 223.8952, 219.7087, 216.1886, 217.0014, 
    216.6974, 216.3035, 215.7579, 208.6967, 209.8423, 209.667, 203.9085, 
    201.6755,
  229.5706, 227.2094, 225.9878, 223.0608, 218.4228, 214.7005, 211.6472, 
    217.0275, 219.272, 216.004, 212.2504, 208.9051, 210.0362, 203.9743, 
    201.7547,
  229.3161, 228.1484, 225.0571, 222.2077, 216.744, 214.5759, 215.061, 
    216.9416, 217.5192, 216.2056, 213.1663, 209.1218, 212.4824, 208.5713, 
    202.0022,
  228.1623, 225.8416, 224.2074, 220.8289, 217.7254, 218.0962, 217.2531, 
    218.2584, 218.4733, 216.5394, 211.0525, 208.5189, 206.1047, 207.1704, 
    210.9856,
  227.5606, 227.3609, 223.5947, 221.0637, 217.3825, 218.5515, 216.9239, 
    214.7637, 214.441, 212.662, 209.3824, 204.4213, 201.2425, 206.281, 
    212.3536,
  230.741, 226.2505, 223.7791, 222.286, 220.4854, 217.4796, 215.1461, 
    213.4611, 210.8371, 208.8579, 208.8563, 205.7603, 203.1136, 208.8192, 
    213.4778,
  240.6207, 231.3828, 231.9231, 228.2804, 226.0684, 222.0991, 218.1428, 
    218.7553, 213.9417, 210.9549, 209.9278, 208.3599, 214.6451, 211.231, 
    205.2709,
  230.89, 235.0695, 230.2151, 227.1026, 223.4028, 220.2887, 213.1876, 
    217.3276, 218.6752, 210.353, 209.3312, 214.478, 215.865, 216.0209, 
    210.5401,
  234.6486, 231.0927, 229.9498, 225.5289, 222.1904, 219.9542, 217.7373, 
    205.9829, 210.0182, 209.8395, 214.5538, 216.8163, 216.0058, 212.3523, 
    208.5404,
  230.8552, 232.0472, 228.4763, 224.6836, 220.9627, 221.6546, 215.999, 
    213.9941, 213.2914, 209.7421, 212.7971, 215.1627, 215.7881, 211.646, 
    208.9312,
  231.6435, 229.8443, 227.3658, 223.8007, 220.9352, 216.7605, 215.1271, 
    213.2371, 213.8739, 212.3447, 212.0123, 213.6851, 211.2207, 209.3148, 
    205.0513,
  237.7118, 229.2269, 226.4643, 223.3558, 221.7098, 216.5831, 210.8529, 
    209.9205, 212.5195, 210.9345, 211.6777, 214.321, 209.7697, 207.9968, 
    206.2176,
  233.6429, 229.4317, 225.621, 225.4959, 223.2296, 215.809, 210.362, 
    211.5758, 207.6388, 209.4863, 213.6897, 211.7564, 207.0936, 206.6877, 
    205.0313,
  232.8828, 229.5423, 226.8939, 225.711, 222.7349, 213.376, 213.1708, 
    211.5718, 210.8878, 207.8383, 210.2057, 209.0491, 208.0143, 209.451, 
    208.8755,
  233.1717, 229.1425, 227.1885, 224.8238, 221.9138, 215.1091, 213.8085, 
    213.4072, 209.7042, 209.5774, 212.0697, 209.5892, 216.331, 216.1381, 
    213.9857,
  233.4263, 231.265, 227.4861, 226.0911, 220.6244, 217.2237, 215.7048, 
    214.8031, 212.5541, 211.1702, 212.2349, 211.0477, 217.364, 213.6738, 
    215.4846,
  241.7833, 236.3028, 232.8217, 227.2216, 225.0049, 221.9755, 217.3262, 
    214.3236, 208.1986, 210.4294, 205.3348, 206.8421, 211.7626, 219.0785, 
    213.7913,
  237.3904, 232.1352, 228.8211, 225.3851, 223.6473, 221.8121, 214.9915, 
    214.3369, 211.9464, 209.6305, 206.6121, 205.2426, 211.6398, 209.0863, 
    217.8465,
  232.869, 231.9451, 227.1778, 223.9242, 222.8797, 218.693, 214.7677, 
    206.6136, 207.0297, 207.7282, 205.7065, 207.8087, 212.3728, 210.0044, 
    211.8726,
  236.009, 230.5449, 226.9095, 223.5545, 221.3558, 214.737, 215.5629, 
    212.1537, 201.8686, 201.5063, 203.4132, 210.3447, 215.0143, 210.1309, 
    211.105,
  232.5709, 229.0312, 225.9835, 223.491, 218.346, 207.3271, 208.7516, 
    211.4218, 203.8304, 203.6785, 204.0104, 206.7275, 214.4888, 211.4755, 
    210.8797,
  234.2854, 228.6971, 225.4477, 222.4491, 216.0997, 205.1227, 200.7823, 
    201.6965, 203.966, 204.2055, 205.315, 206.084, 212.8597, 215.0583, 
    212.3061,
  234.4076, 230.1508, 228.6169, 221.1871, 213.8953, 205.7246, 202.0245, 
    199.5946, 205.5811, 207.6221, 205.3208, 217.4214, 215.6406, 215.8367, 
    215.4494,
  233.4043, 229.6886, 227.2356, 222.6302, 216.4616, 210.6923, 204.0163, 
    201.3356, 204.6434, 208.1654, 208.3552, 218.1385, 212.4942, 217.5944, 
    217.5707,
  233.3437, 229.7491, 227.3567, 222.9921, 217.9675, 211.8129, 206.5038, 
    203.0378, 206.7502, 211.025, 211.6236, 212.0072, 223.4954, 219.9234, 
    219.0208,
  238.3315, 233.5512, 228.52, 227.2717, 220.5416, 215.2054, 208.6886, 
    206.2468, 206.9517, 213.0675, 213.4357, 206.0041, 221.1102, 223.8839, 
    219.812,
  247.1855, 237.1736, 230.9689, 227.1533, 224.8666, 219.8089, 215.7499, 
    212.9151, 208.8975, 205.7041, 215.3627, 222.1007, 217.5473, 220.1398, 
    219.8653,
  235.6483, 231.6397, 229.1231, 228.3934, 223.4273, 215.3681, 209.1436, 
    211.3083, 211.3688, 205.6775, 213.2171, 222.3047, 218.4301, 218.4143, 
    219.1898,
  233.812, 229.1741, 226.475, 221.8522, 218.2374, 213.6617, 206.881, 
    203.3322, 209.6413, 207.4526, 206.0325, 215.7719, 218.3555, 216.1276, 
    216.8572,
  232.4849, 227.6508, 226.742, 222.2089, 215.1147, 211.2968, 202.7569, 
    203.08, 212.5444, 208.4311, 202.3134, 213.8051, 220.9808, 214.5603, 
    218.7986,
  231.6362, 227.5661, 227.5726, 223.7049, 214.5713, 210.5175, 202.4571, 
    199.6688, 204.8576, 209.7724, 203.7443, 208.8172, 213.2381, 215.3402, 
    218.1244,
  231.4345, 227.5716, 229.4234, 224.7126, 219.2972, 210.2629, 202.863, 
    207.341, 208.4641, 204.4191, 200.7039, 206.0158, 210.6038, 214.0351, 
    215.9397,
  230.8819, 230.6953, 228.053, 227.4306, 220.3772, 210.8624, 209.2308, 
    216.6171, 212.9527, 212.0469, 202.6585, 207.6008, 208.8391, 211.0112, 
    217.2872,
  230.3817, 228.9207, 228.2374, 228.009, 223.6791, 211.7218, 211.3244, 
    222.5364, 219.7982, 218.8433, 204.5232, 209.9474, 208.258, 211.4971, 
    215.7463,
  230.1292, 228.4999, 227.9261, 225.9666, 222.622, 212.2015, 209.1969, 
    219.2978, 221.4592, 215.1059, 204.8417, 207.7111, 208.4628, 211.2395, 
    215.1122,
  230.4373, 228.3165, 227.6166, 225.2956, 220.5806, 214.9546, 208.0713, 
    204.9778, 203.126, 203.4341, 205.444, 208.7615, 210.6445, 211.4039, 
    215.369,
  210.9859, 209.0942, 215.7616, 221.839, 225.4461, 221.6109, 213.7504, 
    213.1562, 210.2716, 211.3104, 215.4229, 223.193, 227.9371, 232.5877, 
    218.2008,
  204.3748, 211.7374, 221.0268, 226.7803, 222.7231, 213.6038, 210.9854, 
    211.3954, 211.3795, 209.6823, 212.3467, 222.1862, 226.2722, 220.8046, 
    211.4448,
  201.7142, 214.6877, 226.0302, 227.1544, 218.5021, 210.653, 202.6136, 
    206.9725, 209.252, 202.4084, 213.5247, 219.0382, 224.6202, 215.9122, 
    203.7632,
  207.7872, 222.8659, 227.8482, 227.7992, 215.6775, 207.3998, 211.9518, 
    208.8286, 208.945, 207.904, 212.6114, 218.9083, 220.3216, 210.8955, 
    209.8369,
  220.0807, 226.0784, 228.1912, 228.0181, 208.9211, 206.9981, 205.0788, 
    196.1023, 212.8332, 217.0136, 215.0443, 217.7093, 213.2256, 207.5999, 
    215.3236,
  225.1764, 227.6687, 227.9024, 226.8801, 210.1837, 206.905, 214.8772, 
    220.791, 217.8894, 216.1524, 216.9949, 213.5658, 210.7888, 208.9549, 
    216.0846,
  229.3409, 228.062, 227.4339, 225.4407, 212.2672, 219.778, 228.371, 
    218.1447, 213.2197, 212.4569, 211.7268, 203.5897, 204.1302, 206.3992, 
    211.0612,
  228.611, 228.6537, 226.0733, 210.3668, 205.6517, 209.5777, 216.1083, 
    211.9928, 211.8177, 210.0946, 206.8, 204.4452, 200.0713, 210.4742, 
    209.1929,
  228.6066, 225.1695, 212.284, 206.1761, 205.4841, 206.0928, 207.8786, 
    211.1905, 203.0598, 204.756, 201.8857, 204.4486, 200.4737, 204.0758, 
    208.3694,
  229.8139, 219.2335, 208.8163, 206.493, 205.5705, 209.6048, 207.0402, 
    206.312, 203.1693, 202.7235, 201.1614, 205.4839, 203.565, 204.919, 208.197,
  213.2373, 214.132, 211.1348, 213.0421, 217.0403, 219.8755, 220.4068, 
    219.5668, 222.845, 228.1831, 221.1464, 223.962, 229.0872, 235.4131, 
    214.5815,
  209.6616, 209.7065, 209.4664, 213.674, 218.4324, 218.162, 220.5663, 
    222.0298, 218.8931, 216.4696, 219.311, 226.1541, 232.5364, 231.2745, 
    211.4991,
  202.5523, 200.8199, 208.2617, 214.0445, 222.989, 222.4247, 216.9622, 
    215.0042, 213.0946, 226.7107, 227.969, 223.6619, 232.0784, 227.4648, 
    206.5574,
  193.5884, 200.2625, 211.8401, 220.6575, 228.8938, 223.4897, 227.433, 
    228.5904, 211.4458, 220.7359, 223.7514, 224.4166, 232.48, 221.5208, 
    208.9325,
  198.7116, 215.7977, 224.1859, 226.7412, 225.5772, 208.0179, 213.9202, 
    207.129, 224.5865, 228.5891, 226.0777, 226.6771, 229.7599, 213.6526, 
    210.6634,
  223.2496, 226.8834, 227.1697, 227.4057, 215.1972, 206.7851, 211.2007, 
    222.9944, 218.0025, 227.6266, 231.5293, 231.4414, 220.3948, 210.429, 
    216.294,
  228.0991, 228.0924, 227.0806, 224.3987, 213.5464, 214.7932, 213.3513, 
    219.7507, 220.407, 231.749, 230.814, 223.3108, 213.3141, 212.3636, 
    215.1471,
  230.6999, 230.6018, 226.8853, 219.133, 210.8235, 216.3231, 212.1337, 
    216.1209, 225.3626, 228.4352, 221.1592, 211.4538, 210.6834, 216.0412, 
    222.873,
  236.5971, 221.7711, 207.5591, 206.5909, 208.6271, 213.31, 207.2582, 
    214.9127, 221.2161, 213.2378, 204.4866, 204.2484, 214.4635, 220.8382, 
    224.5087,
  236.6501, 208.3403, 207.0698, 212.2627, 211.558, 208.6376, 214.2631, 
    216.4745, 204.6175, 201.5473, 200.226, 209.9937, 218.6824, 219.4424, 
    225.2406,
  203.7457, 218.2937, 225.2027, 230.4531, 230.2181, 232.4099, 229.1558, 
    224.6168, 223.981, 225.0929, 232.0989, 231.1916, 239.3402, 235.386, 
    228.335,
  192.426, 205.3578, 220.337, 220.2266, 223.4544, 223.1678, 220.4244, 
    223.125, 227.8533, 231.8934, 234.9728, 231.5438, 237.2495, 230.7636, 
    212.8038,
  188.9259, 195.7003, 204.4789, 213.1307, 215.7975, 223.0928, 220.0547, 
    223.3659, 229.2992, 231.909, 233.0383, 231.3192, 236.6853, 221.9878, 
    200.0142,
  189.629, 193.9517, 201.5426, 208.1432, 211.1957, 220.5137, 226.0398, 
    229.4085, 233.5707, 233.3581, 231.2729, 232.1257, 228.1195, 208.9495, 
    202.864,
  196.7724, 199.776, 205.6162, 209.5213, 216.4095, 220.2458, 232.2705, 
    223.5724, 228.3141, 237.0014, 233.2941, 228.5083, 218.7133, 212.2117, 
    213.78,
  207.6611, 213.9254, 220.7713, 221.5681, 226.883, 225.3976, 221.9807, 
    228.8108, 237.0869, 237.1185, 234.0771, 225.6946, 218.118, 219.7881, 
    217.7732,
  224.2646, 224.6653, 225.6839, 228.1309, 225.422, 221.2342, 219.808, 
    224.6714, 236.0761, 236.395, 229.0268, 221.7818, 224.1183, 217.6338, 
    217.8774,
  225.3976, 224.6386, 231.3557, 231.3295, 217.7152, 216.3774, 222.7852, 
    230.9123, 235.5681, 232.2047, 224.6013, 222.739, 220.3784, 215.8074, 
    214.0729,
  240.2464, 226.3723, 224.8843, 214.1663, 222.9687, 221.3297, 230.7922, 
    225.8794, 232.2522, 226.3319, 222.6556, 223.5463, 214.9113, 214.5702, 
    219.2216,
  236.8118, 213.2847, 211.1399, 216.979, 229.2968, 225.4006, 235.6525, 
    233.1236, 228.1358, 223.5305, 214.6175, 214.4284, 212.6275, 220.4531, 
    230.2983,
  243.8565, 239.6293, 232.1072, 218.9565, 209.0144, 220.683, 233.697, 
    240.3847, 233.993, 227.6685, 229.4752, 233.0442, 235.6497, 236.3769, 
    237.3465,
  235.4369, 236.4509, 227.1471, 210.4055, 205.8542, 220.3476, 235.1062, 
    238.6224, 233.5772, 228.9285, 230.1977, 234.057, 234.1379, 234.6812, 
    236.0764,
  234.5907, 229.2842, 222.9052, 208.1306, 206.306, 212.8472, 232.6854, 
    231.5639, 226.2087, 227.6943, 229.3104, 233.9506, 234.542, 234.0641, 
    231.7209,
  225.8043, 227.0661, 213.0736, 198.4529, 198.3759, 210.79, 228.6937, 
    229.7277, 226.5499, 227.8387, 235.0162, 234.8113, 232.7793, 227.6284, 
    231.5097,
  214.0889, 212.9894, 198.9506, 192.1756, 190.366, 195.8284, 211.6333, 
    223.2829, 226.1703, 233.2069, 239.0389, 234.8678, 231.8471, 223.0377, 
    227.7194,
  206.2849, 200.531, 190.801, 182.8051, 188.2599, 195.8225, 202.3677, 
    216.2245, 231.3909, 236.4613, 237.1996, 234.7519, 228.6054, 225.3837, 
    225.0052,
  197.7662, 191.7133, 188.1444, 186.8778, 192.1479, 201.0168, 216.0167, 
    228.4412, 233.9177, 236.7765, 235.2067, 231.354, 227.709, 221.9393, 
    218.3743,
  204.8162, 195.0569, 191.2337, 192.5318, 199.4497, 211.0134, 225.2795, 
    233.4577, 236.1897, 238.9095, 232.4519, 222.0752, 222.3085, 221.4833, 
    220.4265,
  210.6569, 204.6845, 201.0439, 199.9511, 201.645, 214.0589, 226.5197, 
    233.1428, 236.6125, 238.8814, 227.1549, 221.2546, 215.9098, 224.7996, 
    217.9013,
  220.3179, 212.9401, 204.6247, 203.2823, 210.6, 216.9172, 228.2869, 
    240.0453, 240.3805, 236.2143, 221.3556, 220.5387, 220.2273, 225.5343, 
    219.7292,
  181.6585, 198.7924, 216.6106, 222.4678, 218.046, 219.1959, 225.8738, 
    227.6202, 231.5118, 236.4701, 238.6718, 238.3856, 237.4927, 236.6201, 
    237.9839,
  188.2446, 205.4455, 215.3682, 217.9694, 220.1207, 224.435, 227.7275, 
    228.3293, 231.7931, 235.4464, 234.5268, 234.9687, 236.0778, 236.3439, 
    238.7724,
  198.8521, 204.4157, 214.0029, 218.1913, 221.15, 222.9254, 226.7144, 226.93, 
    230.4918, 232.1548, 232.3569, 233.7015, 234.7015, 233.5441, 234.667,
  194.9765, 197.9308, 213.2778, 224.5797, 221.2814, 224.1316, 225.6956, 
    231.7914, 230.6328, 231.42, 233.1374, 233.3122, 233.5928, 227.67, 230.3058,
  189.7827, 199.5837, 215.1391, 228.4765, 224.5775, 216.3709, 220.4955, 
    232.1545, 229.8187, 231.1699, 229.9832, 234.0361, 230.781, 224.8273, 
    223.9925,
  197.5249, 205.7188, 223.0957, 234.3923, 230.7823, 224.9241, 215.018, 
    221.5037, 223.7299, 228.6252, 229.4902, 226.4045, 224.0559, 225.2333, 
    229.668,
  198.5078, 211.0683, 229.3648, 232.2987, 228.1233, 220.9048, 214.1421, 
    219.4823, 223.6599, 226.6963, 231.1955, 224.7373, 225.1243, 222.5994, 
    221.018,
  205.4304, 217.4451, 224.2894, 223.8149, 220.2087, 216.0871, 220.3826, 
    230.738, 236.7273, 235.0435, 226.3578, 222.1478, 225.1112, 224.7474, 
    220.0456,
  203.8147, 215.546, 216.1377, 218.8693, 208.2229, 208.515, 225.8739, 
    236.4676, 237.3652, 227.1704, 219.2214, 216.5932, 216.403, 218.8982, 
    208.6275,
  203.2436, 211.5282, 210.0394, 207.4465, 198.8574, 203.9712, 233.7192, 
    239.9274, 238.7912, 227.2927, 220.9588, 214.678, 214.394, 209.4044, 
    205.0641,
  232.6882, 231.6779, 207.9024, 208.4314, 222.6413, 241.0419, 243.1321, 
    228.8328, 213.2241, 199.4952, 199.3206, 210.6748, 218.8727, 224.8541, 
    235.328,
  216.0068, 223.2119, 213.7029, 217.4036, 232.0557, 244.0977, 244.8031, 
    234.5465, 222.1455, 203.9635, 205.8971, 210.7868, 220.1478, 228.6341, 
    234.7158,
  216.7341, 228.5647, 221.8786, 224.8969, 236.3547, 244.0577, 244.7737, 
    237.0307, 218.8777, 208.3644, 205.8453, 206.9796, 216.4315, 226.7567, 
    231.7699,
  233.8152, 239.5957, 236.6224, 228.976, 239.4872, 243.8667, 239.1826, 
    238.1304, 233.6772, 218.6236, 208.8794, 207.1736, 216.1684, 222.2904, 
    228.3012,
  233.2215, 239.4437, 240.1246, 237.0925, 237.654, 232.756, 230.771, 
    231.3792, 233.6584, 224.7523, 213.2345, 210.6846, 209.9749, 219.2415, 
    215.7571,
  230.1068, 234.294, 237.6518, 237.1971, 236.3952, 230.3783, 222.1225, 
    214.3992, 215.3617, 214.4906, 212.7492, 204.661, 205.1736, 208.5784, 
    215.9089,
  230.1441, 234.8084, 235.6456, 234.4875, 227.4478, 223.257, 220.6962, 
    207.3174, 203.985, 202.3411, 205.1601, 201.5242, 201.8647, 205.9759, 
    215.9808,
  232.3178, 232.5294, 229.4765, 228.4574, 227.7039, 218.1687, 212.1769, 
    210.6068, 211.4833, 215.1991, 212.2529, 210.9911, 220.3148, 226.5552, 
    230.8425,
  234.9531, 231.1423, 228.5243, 223.8066, 225.5167, 224.1611, 232.7816, 
    237.1454, 233.3905, 235.4746, 232.1374, 230.0834, 226.6476, 235.3255, 
    233.7436,
  234.7067, 233.17, 232.0251, 230.8983, 236.3518, 241.7473, 245.9798, 
    245.3116, 237.6274, 225.1715, 222.5594, 220.5778, 229.2917, 232.425, 
    226.1683,
  235.3768, 230.7709, 226.4242, 205.5764, 217.5042, 235.5336, 244.2941, 
    238.4805, 230.3049, 231.4028, 232.5287, 242.6408, 243.1389, 242.303, 
    244.0432,
  230.4418, 216.2142, 199.4302, 193.7354, 205.7857, 233.8514, 239.9915, 
    236.4759, 230.8804, 228.3936, 231.8593, 234.4775, 230.6993, 233.1772, 
    233.9303,
  217.223, 203.5081, 188.1159, 187.9206, 209.1137, 223.5652, 236.6246, 
    228.0824, 221.022, 220.9148, 230.2078, 226.8585, 224.4971, 219.5806, 
    221.6399,
  212.8843, 198.2873, 185.7823, 189.3016, 205.5667, 221.6279, 227.3811, 
    229.6401, 219.3839, 215.5343, 220.1805, 226.2611, 220.312, 216.6954, 
    214.107,
  213.4118, 202.6976, 196.102, 198.1109, 208.107, 225.1616, 232.8544, 
    230.2668, 228.1338, 209.1571, 211.6297, 218.138, 214.6366, 212.708, 
    211.2048,
  231.0715, 231.1264, 223.1455, 218.0734, 222.4079, 231.1216, 238.1221, 
    228.5978, 226.5942, 210.4799, 202.1704, 206.0567, 206.6034, 208.3334, 
    205.6177,
  239.4909, 240.4994, 242.6088, 242.9386, 236.5618, 236.6102, 240.5291, 
    227.38, 225.7691, 215.0191, 203.7264, 198.3769, 200.7869, 197.7175, 
    196.074,
  238.6757, 238.9025, 241.4197, 244.0607, 242.0416, 239.1582, 235.7117, 
    224.8533, 226.0376, 217.9694, 207.2216, 197.4068, 192.9967, 191.8, 
    194.0344,
  226.0499, 226.4744, 225.9908, 226.8324, 228.6597, 230.8997, 228.4283, 
    220.7207, 221.1406, 220.8143, 215.1481, 208.3085, 206.5002, 202.2472, 
    204.6929,
  232.2514, 234.3431, 236.093, 235.898, 234.262, 234.7285, 235.5591, 
    231.4371, 231.0216, 230.5433, 226.02, 220.3843, 219.1606, 215.5879, 
    212.8973,
  221.5739, 223.8502, 223.5961, 224.5466, 216.2454, 216.323, 218.0318, 
    220.0919, 230.8981, 230.5748, 235.7254, 235.2439, 242.2378, 245.1086, 
    248.3774,
  223.0389, 221.011, 217.5643, 220.8911, 222.5843, 230.2139, 225.6295, 
    222.4255, 227.5144, 233.7041, 234.949, 237.8145, 244.5146, 245.8629, 
    248.6919,
  223.9041, 219.8085, 215.0285, 211.8677, 221.0408, 228.2117, 234.5687, 
    223.0089, 227.8452, 235.0489, 235.9532, 239.9815, 245.6449, 246.5942, 
    247.8618,
  228.1338, 221.2574, 206.0034, 209.1508, 208.6004, 230.1185, 230.2399, 
    228.5702, 232.4587, 235.4718, 237.3383, 241.6789, 245.8481, 247.1883, 
    245.8032,
  231.4676, 223.118, 207.0641, 209.6001, 212.9177, 218.7517, 234.0111, 
    230.0776, 233.6869, 240.6306, 238.1806, 244.8391, 246.359, 247.7328, 
    247.8042,
  227.9824, 223.3125, 217.8141, 221.1389, 223.8408, 224.917, 234.5037, 
    238.1592, 237.8811, 237.1283, 240.1087, 244.9962, 247.2524, 247.7467, 
    249.341,
  220.1097, 219.0649, 222.4987, 228.2735, 223.1319, 227.4462, 235.4273, 
    237.3566, 236.4668, 240.371, 243.3092, 245.843, 247.8274, 247.4059, 
    250.6546,
  218.6466, 221.3064, 219.796, 215.99, 220.1438, 222.6598, 236.1132, 
    237.1056, 237.6961, 238.6021, 237.0403, 244.5181, 246.4834, 246.4419, 
    246.4512,
  220.934, 215.3126, 212.957, 213.397, 212.4086, 220.4607, 232.8462, 
    230.1016, 234.3944, 235.5793, 234.7357, 236.3515, 236.6957, 240.5027, 
    239.3039,
  222.404, 218.0735, 215.5591, 212.5752, 216.9552, 221.0264, 226.9513, 
    222.5891, 225.1836, 227.146, 227.0051, 229.8296, 231.6939, 232.8139, 
    229.0707,
  223.2181, 224.2133, 226.9783, 226.7123, 221.8453, 228.3086, 230.5004, 
    225.3742, 227.3695, 224.2677, 226.2319, 222.5804, 212.5746, 216.5136, 
    218.2606,
  225.9468, 229.2014, 228.8574, 228.5586, 225.5347, 224.2658, 224.0867, 
    227.0924, 230.9926, 223.6819, 219.3603, 220.7286, 208.3767, 210.7963, 
    216.4337,
  232.0686, 229.8251, 227.9168, 224.7868, 222.0747, 223.9088, 226.5683, 
    224.6039, 228.3086, 226.5158, 216.5729, 209.1851, 202.9803, 208.3301, 
    215.1453,
  222.7982, 219.4231, 224.6075, 225.8673, 222.646, 224.9226, 223.9399, 
    229.015, 234.6982, 232.8201, 217.5291, 206.6542, 205.7697, 210.319, 
    219.6607,
  215.6062, 220.5843, 225.4134, 223.7922, 224.0085, 219.2366, 221.3192, 
    222.3221, 227.0601, 234.6251, 214.4813, 206.7717, 208.5051, 216.4138, 
    223.8925,
  215.6519, 219.0511, 222.9734, 228.1626, 229.4593, 219.6146, 220.517, 
    222.5368, 235.4279, 231.3696, 211.5207, 211.8406, 217.5041, 223.0186, 
    229.0593,
  215.8557, 217.0025, 215.648, 222.1234, 227.5866, 220.9964, 220.9262, 
    215.5895, 227.9319, 227.3615, 211.9706, 217.301, 223.7324, 227.9672, 
    230.6437,
  216.6077, 209.3486, 207.5897, 227.2168, 224.8757, 217.6021, 219.3861, 
    221.0217, 236.8921, 223.324, 210.5954, 219.2059, 227.3544, 225.7801, 
    229.8036,
  217.0446, 214.73, 205.631, 217.1795, 221.4513, 212.6097, 219.7914, 
    212.8539, 233.4362, 214.4941, 215.5487, 221.7427, 225.6229, 225.277, 
    227.0822,
  216.8705, 214.2807, 208.8815, 209.0054, 211.2098, 213.2782, 212.5953, 
    216.2986, 229.3186, 216.6679, 219.945, 223.2298, 222.3412, 225.5265, 
    229.4496,
  225.1909, 221.3838, 222.9129, 223.0831, 227.1875, 228.0489, 227.2734, 
    226.3473, 229.5252, 231.6224, 233.6955, 232.6559, 233.6245, 238.478, 
    240.302,
  225.0883, 229.3286, 233.5889, 233.5118, 233.5164, 233.9919, 229.3384, 
    228.4121, 232.7984, 229.0032, 227.7078, 235.1154, 234.9569, 236.4529, 
    240.9556,
  236.8054, 237.4704, 232.7117, 229.2994, 228.6291, 225.8955, 228.6353, 
    221.0786, 223.7588, 226.9113, 227.1632, 225.6374, 227.396, 235.8628, 
    238.6774,
  238.4193, 233.4429, 228.1577, 223.1236, 222.4739, 225.8878, 221.7803, 
    225.3293, 224.7804, 224.3093, 225.5303, 222.6926, 230.7321, 234.6483, 
    231.2621,
  229.4424, 221.2874, 213.4487, 214.6297, 216.9206, 217.7792, 222.2825, 
    220.8435, 224.6894, 226.9344, 223.259, 217.8026, 221.6058, 228.951, 
    227.9351,
  215.6023, 209.2676, 208.7603, 209.6087, 210.8537, 216.0055, 220.733, 
    226.219, 227.3817, 230.2271, 223.2472, 216.8539, 221.0178, 228.1045, 
    225.7706,
  209.4623, 208.8334, 203.6755, 203.7921, 209.8112, 222.2481, 222.2976, 
    226.0651, 228.9291, 231.1373, 216.0096, 214.6409, 219.5412, 226.629, 
    227.062,
  206.6279, 206.5443, 212.3997, 211.045, 217.5102, 225.6575, 227.9031, 
    232.598, 231.4825, 219.2182, 210.8541, 212.9316, 222.9839, 230.0175, 
    229.4623,
  205.9138, 210.8678, 213.0966, 214.2885, 222.1289, 221.0086, 229.5746, 
    230.7321, 220.0236, 207.6678, 206.5667, 215.9605, 228.6801, 233.7299, 
    236.2652,
  205.6689, 212.2731, 212.7956, 212.6393, 219.9415, 228.8289, 226.85, 
    221.9415, 206.1372, 203.679, 212.3797, 222.0747, 232.0253, 237.1483, 
    242.9528,
  193.3564, 196.8316, 195.8792, 200.6293, 208.6065, 212.4978, 216.5932, 
    217.701, 221.7605, 224.9422, 242.5103, 240.3171, 238.4062, 239.7228, 
    214.5438,
  189.7324, 194.8593, 204.5413, 206.6967, 216.0488, 220.6978, 224.063, 
    234.4513, 239.0372, 240.1349, 240.5141, 238.7945, 239.0695, 233.9555, 
    205.3163,
  194.8558, 201.3677, 212.8478, 215.4864, 219.7663, 224.127, 228.7536, 
    234.2572, 238.6221, 238.2172, 237.5964, 239.2402, 240.5966, 226.554, 
    194.635,
  210.0652, 215.8045, 222.8542, 230.3336, 229.1755, 234.2607, 233.2152, 
    237.4382, 239.2656, 239.3295, 239.701, 240.0927, 239.2566, 212.8487, 
    189.8219,
  217.5285, 219.9324, 221.4244, 225.4549, 227.0314, 225.5079, 226.9327, 
    226.6002, 234.0328, 235.3242, 235.7077, 237.2438, 232.596, 204.4186, 
    195.0267,
  222.7057, 222.4834, 222.3174, 223.2077, 223.8933, 221.8819, 221.3874, 
    224.4793, 225.4889, 230.9568, 238.7609, 238.6518, 233.8787, 203.149, 
    205.0109,
  230.4989, 226.8032, 227.4189, 226.3541, 221.9274, 216.1709, 214.2803, 
    212.1544, 214.7234, 231.5499, 234.9977, 235.8978, 229.1782, 203.3726, 
    208.2927,
  224.4973, 223.4862, 225.0271, 219.2815, 212.7663, 209.3705, 209.4845, 
    212.7907, 222.6502, 233.857, 234.1572, 235.2937, 227.2332, 206.3295, 
    222.4584,
  224.9667, 222.2244, 217.2674, 214.0194, 209.6598, 205.4804, 207.5286, 
    211.2193, 220.6198, 231.718, 233.9541, 234.3656, 226.3956, 217.7827, 
    229.5496,
  227.8926, 221.1884, 212.1341, 212.2734, 215.6869, 215.159, 214.3885, 
    217.226, 226.3337, 233.0889, 235.3635, 232.6285, 223.4861, 229.3408, 
    230.0187,
  233.8932, 233.5543, 212.5764, 196.9617, 194.0328, 203.2165, 190.5847, 
    189.3407, 183.1716, 199.7603, 209.0072, 227.7322, 242.101, 243.9348, 
    238.3363,
  210.8469, 232.035, 218.9996, 202.1289, 194.4668, 195.1902, 189.7603, 
    190.1082, 192.6819, 205.5416, 215.781, 229.3499, 241.6837, 239.8033, 
    239.4375,
  197.7114, 216.5677, 215.8087, 202.026, 193.6364, 193.8997, 190.0691, 
    187.0832, 198.9636, 205.8053, 217.6404, 235.5489, 240.4572, 240.2, 
    241.9553,
  193.4859, 195.799, 199.4008, 198.7806, 200.122, 198.773, 194.7867, 195.836, 
    199.0319, 210.1746, 221.4202, 236.807, 240.8923, 238.5478, 240.1793,
  191.3618, 186.7668, 188.3304, 192.6219, 198.1673, 193.9007, 204.3202, 
    208.4523, 209.1641, 211.7021, 225.9111, 240.7391, 238.6359, 232.6477, 
    233.809,
  198.1893, 182.8519, 190.7107, 194.0692, 203.8918, 200.378, 200.0233, 
    203.6486, 211.6266, 223.3981, 235.6851, 238.3597, 235.4066, 227.378, 
    224.4807,
  223.4992, 190.825, 190.4183, 199.8686, 203.1287, 205.7682, 210.8393, 
    210.1149, 219.8129, 233.2719, 238.4247, 236.2508, 229.5435, 219.6691, 
    220.1576,
  240.366, 206.6431, 197.3357, 201.8294, 211.9553, 212.6469, 220.4941, 
    234.1641, 238.1142, 237.6395, 236.3813, 234.3936, 225.4068, 211.9786, 
    213.6153,
  233.1075, 227.6909, 206.8587, 204.2009, 211.2674, 216.5997, 223.7946, 
    235.1184, 237.0517, 235.6847, 235.4966, 230.2488, 212.1358, 204.8037, 
    216.4476,
  235.1809, 235.0178, 221.9885, 214.8771, 214.0978, 216.8968, 222.0681, 
    229.7017, 233.6784, 234.4278, 231.6351, 225.3495, 199.6632, 205.8323, 
    225.9479,
  232.9039, 228.8556, 217.0599, 225.2899, 245.4102, 247.7832, 236.7652, 
    212.1138, 197.6374, 197.6371, 192.6161, 190.8188, 194.8118, 200.5932, 
    210.9334,
  223.149, 227.2727, 216.3191, 220.1467, 234.4907, 230.1478, 207.3616, 
    200.0831, 194.2999, 184.8822, 188.4537, 191.5076, 194.8569, 208.6119, 
    230.6464,
  223.0424, 223.1498, 218.3394, 212.3233, 221.8886, 211.9737, 199.9219, 
    192.9056, 194.2996, 186.6134, 185.5662, 191.4894, 205.3145, 226.3326, 
    238.3873,
  220.0286, 222.7027, 224.96, 211.8488, 206.6029, 208.3571, 195.7967, 
    202.0191, 200.598, 194.9612, 189.3714, 197.2842, 223.102, 237.3159, 
    239.3859,
  219.3465, 220.0656, 222.9111, 225.2313, 215.2902, 204.1475, 213.9293, 
    224.812, 206.7223, 191.4599, 195.1757, 212.4457, 234.4577, 236.4772, 
    236.4666,
  223.282, 223.4724, 223.1059, 232.0927, 225.9159, 224.8214, 218.1661, 
    201.7288, 195.9034, 196.6427, 205.0454, 232.6213, 234.5188, 234.0659, 
    234.5161,
  232.0304, 235.6432, 221.3838, 230.8432, 222.7591, 218.3004, 218.7741, 
    203.1881, 199.1821, 210.3647, 233.0433, 234.3983, 233.2983, 233.9695, 
    230.3272,
  229.3644, 231.4822, 216.643, 220.4748, 220.5832, 210.2544, 205.7312, 
    198.8206, 208.3987, 226.6499, 234.3235, 231.9195, 230.3727, 226.7814, 
    226.1358,
  235.267, 236.0991, 214.3447, 210.8741, 207.7775, 200.2338, 197.6147, 
    197.1145, 211.5181, 231.0116, 231.594, 230.5963, 228.2086, 224.3212, 
    228.6074,
  233.6772, 232.319, 212.0986, 200.9548, 199.7484, 197.8598, 190.7153, 
    200.612, 224.5048, 231.2141, 231.2008, 229.2861, 222.7788, 228.445, 
    228.8339,
  227.4355, 211.1537, 204.0038, 214.2346, 225.917, 226.3843, 231.8068, 
    243.3823, 240.6288, 233.0563, 221.1526, 203.2467, 193.7964, 193.4632, 
    204.0321,
  225.5057, 210.7784, 203.8175, 209.8734, 223.4875, 224.5155, 229.1316, 
    238.8689, 240.6045, 239.32, 232.4732, 224.7131, 222.2451, 214.7966, 
    220.8366,
  218.9558, 203.0539, 201.017, 203.5303, 217.5161, 225.0908, 228.6156, 
    227.8936, 238.0003, 237.3331, 224.7188, 218.4689, 215.1792, 224.7515, 
    239.5529,
  227.7529, 218.5411, 207.4715, 207.3308, 209.1351, 216.7082, 225.2754, 
    228.7339, 227.8477, 223.04, 212.5369, 210.2301, 218.6508, 235.3069, 
    239.8385,
  233.8766, 224.6097, 217.5175, 211.513, 214.6207, 213.887, 222.606, 231.147, 
    218.6843, 208.2868, 205.5371, 205.8881, 223.031, 234.584, 237.6301,
  230.1591, 220.5527, 215.9938, 215.6423, 218.6672, 216.5128, 220.8888, 
    215.1958, 213.6073, 214.6389, 210.567, 222.0966, 227.2177, 233.5182, 
    233.1284,
  231.1844, 224.9036, 220.5518, 217.2502, 213.7192, 215.6339, 213.6213, 
    208.732, 209.1436, 209.9981, 215.7522, 221.5368, 232.4788, 233.7131, 
    229.7643,
  220.9905, 214.6154, 212.0433, 214.3004, 208.303, 205.4033, 206.282, 
    204.2368, 207.8163, 208.1599, 219.5637, 230.2452, 230.4217, 229.0341, 
    226.0291,
  205.9721, 197.4445, 198.267, 200.856, 201.9835, 200.6082, 203.2457, 
    204.9884, 206.4667, 212.4509, 226.9346, 230.9226, 229.3438, 222.868, 
    219.3669,
  201.8398, 195.5645, 191.9274, 195.291, 197.5567, 197.7311, 206.5251, 
    210.5964, 210.7793, 225.2542, 230.6246, 230.2162, 226.4344, 218.9104, 
    215.5273,
  212.1373, 211.4645, 209.3459, 214.7063, 217.4784, 216.5102, 216.9803, 
    221.489, 220.2251, 225.4379, 225.2335, 227.3814, 226.0611, 225.0934, 
    224.6414,
  201.6047, 203.7884, 204.1212, 209.1316, 215.6748, 217.6799, 212.4996, 
    219.509, 220.4533, 221.6731, 217.828, 219.6246, 219.8911, 217.3004, 
    218.4618,
  205.1149, 210.1594, 211.3011, 212.7013, 213.9224, 217.6292, 216.8686, 
    216.1225, 215.263, 218.9864, 217.4727, 213.2886, 214.0169, 212.2008, 
    218.0916,
  214.2582, 221.095, 223.552, 229.944, 233.8579, 236.381, 231.1816, 227.1534, 
    219.1246, 208.5629, 210.7301, 207.9856, 210.051, 200.9675, 208.3322,
  228.2875, 231.5012, 236.0602, 239.1767, 240.9201, 240.86, 238.4907, 
    231.2074, 223.8734, 217.7775, 209.8907, 209.8148, 203.0442, 203.7946, 
    208.0577,
  235.7225, 239.1222, 243.4181, 243.437, 245.1461, 246.1259, 241.2783, 
    234.7967, 225.6002, 219.3944, 212.2898, 208.332, 206.5272, 208.9653, 
    216.1288,
  246.4062, 246.4787, 245.0202, 245.3422, 246.1201, 246.0664, 242.6093, 
    234.9075, 222.7189, 219.5014, 217.2791, 211.7906, 208.2614, 212.7231, 
    221.8955,
  249.377, 247.1793, 244.0599, 243.6416, 242.7796, 240.6259, 237.6258, 
    228.871, 226.5476, 221.0791, 212.6879, 215.2787, 214.1404, 217.5267, 
    224.0862,
  245.3155, 242.8262, 236.5745, 232.3473, 232.843, 233.3112, 230.7989, 
    225.3329, 220.7073, 215.342, 215.0272, 216.5005, 215.8082, 222.028, 
    230.0125,
  242.9129, 237.8369, 207.6736, 207.3154, 222.7248, 227.814, 226.2933, 
    219.8578, 217.0526, 213.825, 213.3226, 216.2479, 224.2063, 230.8844, 
    229.5596,
  233.0447, 231.1306, 226.4648, 214.2286, 203.9998, 197.0162, 189.933, 
    184.6035, 191.8851, 196.6282, 198.8411, 198.1552, 201.2751, 202.6329, 
    202.7668,
  213.8008, 212.5733, 207.2597, 201.6803, 201.6925, 194.5819, 192.6786, 
    194.4365, 199.134, 201.5652, 204.327, 203.3835, 206.5298, 209.0508, 
    208.6186,
  203.3674, 198.8929, 198.8288, 197.8212, 204.3573, 197.8343, 196.6916, 
    194.6496, 202.3402, 208.2335, 207.3523, 208.7152, 211.3526, 210.0558, 
    211.0121,
  196.3768, 190.4572, 192.1681, 197.8602, 200.4344, 206.7331, 210.4715, 
    211.8435, 212.7457, 211.1578, 216.3104, 218.5476, 215.6786, 214.3209, 
    215.177,
  199.2659, 199.1958, 200.4466, 212.4091, 214.4592, 220.9709, 225.5859, 
    231.8728, 232.9188, 236.1295, 234.6285, 237.6068, 235.2934, 228.8314, 
    227.9191,
  210.5469, 216.3977, 220.9871, 226.9428, 230.7907, 235.3595, 235.7024, 
    236.8624, 236.1792, 236.087, 236.8812, 238.2792, 236.8324, 232.109, 
    225.3367,
  226.6348, 228.1179, 230.5205, 234.3251, 237.1691, 236.9095, 234.882, 
    233.8998, 234.4252, 232.342, 232.7245, 235.7742, 235.2339, 230.131, 
    222.6708,
  229.9903, 233.9103, 235.5396, 236.4801, 235.6122, 230.4663, 226.0536, 
    221.398, 215.7087, 215.7013, 214.3844, 219.6937, 225.0996, 217.2457, 
    216.9047,
  233.445, 235.6252, 236.3595, 233.6953, 232.3244, 227.8374, 225.0693, 
    220.0182, 216.3441, 213.4326, 215.9727, 221.6668, 220.2735, 214.9733, 
    211.2678,
  239.2115, 237.9176, 230.9167, 235.0964, 237.2668, 233.5022, 235.0778, 
    225.7983, 217.5711, 218.8798, 220.2471, 217.627, 216.0914, 209.4648, 
    207.5628,
  249.9071, 248.5664, 251.6884, 252.6509, 252.7127, 247.6509, 247.998, 
    246.2189, 239.4387, 237.144, 229.4282, 227.8615, 222.9231, 216.3741, 
    206.7218,
  246.9531, 251.9555, 255.6944, 255.9936, 251.4956, 250.9415, 247.0278, 
    240.6621, 232.2897, 225.9182, 219.6294, 218.4546, 215.2915, 214.3331, 
    209.1046,
  239.3121, 247.367, 250.9401, 248.5905, 247.6339, 241.0838, 236.7479, 
    228.838, 226.9431, 218.3115, 219.224, 215.4239, 212.4803, 210.7891, 
    207.5015,
  216.6924, 221.3248, 225.0834, 232.3468, 230.9314, 232.0199, 224.8499, 
    223.1994, 222.3846, 220.06, 216.5169, 213.924, 213.8326, 213.5739, 
    214.2624,
  212.0005, 208.3409, 206.4538, 202.5038, 210.1599, 215.3987, 217.9498, 
    219.7, 220.5663, 220.4049, 217.204, 220.3161, 219.8436, 219.3761, 214.8541,
  211.2268, 199.5826, 192.3951, 192.7706, 191.2525, 194.2412, 200.6974, 
    213.9684, 221.1691, 226.3429, 224.4585, 224.8073, 225.0465, 224.5197, 
    224.7996,
  217.1706, 208.2424, 199.9779, 195.7665, 203.817, 204.2147, 211.3773, 
    212.2904, 216.0026, 215.9601, 220.2485, 224.0361, 225.2097, 232.5794, 
    233.9255,
  220.4095, 222.3795, 224.4276, 221.7343, 228.4421, 231.2455, 233.5798, 
    235.5984, 234.4582, 231.22, 228.4677, 226.853, 228.9155, 234.9863, 
    228.3379,
  225.4346, 228.5003, 230.6781, 229.4978, 232.3746, 234.8038, 235.5926, 
    235.5114, 235.2802, 232.0349, 224.0921, 223.8697, 223.3235, 232.489, 
    224.4708,
  232.1382, 228.3563, 229.984, 230.4785, 231.0706, 234.5507, 237.3251, 
    237.8217, 235.0884, 227.6994, 219.8825, 214.29, 221.0827, 219.9729, 
    221.9068,
  191.5568, 198.1664, 208.1706, 220.466, 229.3293, 235.6639, 240.4408, 
    244.0519, 245.968, 248.9027, 250.7735, 250.9243, 252.3778, 254.0195, 
    254.7836,
  190.2015, 197.9411, 205.0031, 212.7832, 222.1759, 234.9513, 243.0036, 
    244.5457, 246.2313, 248.2635, 251.3577, 250.0071, 250.5658, 249.7991, 
    251.2179,
  198.703, 204.5285, 210.721, 213.9781, 223.0762, 231.6847, 239.7445, 
    242.2293, 244.5381, 245.8599, 248.166, 248.8096, 250.1616, 248.972, 
    247.1322,
  213.9625, 215.4253, 218.5232, 220.869, 224.877, 228.1958, 231.3519, 
    239.991, 241.8349, 244.9668, 246.7101, 248.4741, 249.6021, 248.2326, 
    246.4597,
  226.2503, 226.0314, 226.0698, 226.4966, 227.268, 225.083, 230.0127, 
    233.0823, 232.1731, 239.3133, 241.7297, 245.1665, 247.591, 246.785, 
    242.712,
  233.733, 230.2814, 231.1816, 230.5959, 228.7379, 224.632, 220.6618, 
    226.9778, 224.7347, 229.248, 229.8925, 229.1026, 234.8927, 235.1512, 
    230.4906,
  228.481, 229.3543, 227.4965, 225.3319, 222.9301, 219.5928, 221.0327, 
    223.1704, 225.6817, 223.9911, 218.1671, 213.107, 217.2886, 217.192, 
    209.6563,
  223.8699, 223.6278, 219.8349, 218.908, 219.1218, 220.57, 222.6755, 
    228.6416, 228.5079, 230.0027, 227.4343, 216.287, 209.7374, 206.3083, 
    196.384,
  223.6017, 216.5697, 217.7259, 220.2826, 222.2631, 224.8403, 226.2442, 
    229.4518, 231.7917, 232.5396, 228.1682, 226.3103, 221.8369, 207.5623, 
    196.7935,
  221.1726, 219.7241, 222.3589, 223.7826, 227.2769, 225.9272, 225.7003, 
    224.5132, 230.5492, 221.6938, 228.0397, 229.8901, 226.5563, 218.9919, 
    211.1911,
  236.111, 221.4462, 218.3574, 218.6555, 220.3793, 232.7458, 237.0042, 
    231.4822, 231.4081, 235.8167, 236.1674, 230.2048, 233.3646, 238.6544, 
    242.2753,
  235.6611, 234.8472, 223.4671, 212.4765, 224.0438, 222.1543, 233.8484, 
    231.9486, 236.1199, 232.654, 234.021, 231.1452, 236.5265, 240.2395, 
    241.6925,
  230.4277, 228.9053, 221.8634, 215.9494, 213.6113, 210.8388, 220.6318, 
    221.2444, 225.8657, 229.6191, 230.486, 228.9338, 234.5698, 240.4058, 
    237.404,
  217.855, 217.9902, 213.6703, 210.9823, 207.3353, 204.3744, 204.5234, 
    208.1198, 214.0022, 215.7372, 219.0817, 224.8902, 229.9007, 233.8059, 
    232.4263,
  208.7146, 208.1461, 209.7354, 206.6202, 204.3766, 195.6787, 199.9402, 
    205.8268, 213.1966, 207.6865, 213.6049, 223.0483, 226.4054, 229.1562, 
    228.0958,
  217.3688, 208.5357, 208.8861, 206.4097, 205.7955, 204.1987, 204.8147, 
    204.9479, 211.204, 213.1217, 223.8112, 225.7636, 230.0257, 223.78, 
    224.5456,
  229.901, 222.6174, 215.5976, 212.7705, 212.1714, 213.3423, 213.4075, 
    211.0054, 210.7116, 217.34, 225.3033, 231.8219, 229.6997, 221.6116, 
    211.7631,
  234.629, 232.1327, 222.3859, 220.167, 217.5545, 218.0997, 221.3236, 
    222.6927, 220.2399, 224.8599, 227.7986, 230.9718, 224.098, 213.9267, 
    203.6355,
  229.9635, 226.3661, 225.3363, 224.6664, 222.7647, 224.3887, 228.1673, 
    227.6064, 226.2289, 230.2105, 231.2535, 227.2929, 221.9945, 209.4379, 
    195.3387,
  223.2346, 220.3094, 219.9553, 223.4225, 225.9072, 223.1489, 231.4004, 
    229.3681, 230.0403, 235.416, 234.4647, 223.8793, 215.3262, 199.0314, 
    194.2726,
  234.5627, 233.784, 220.1011, 226.3414, 235.238, 250.7794, 256.2926, 
    259.5032, 261.3705, 267.117, 260.7005, 252.8294, 247.7337, 239.1315, 
    234.6898,
  238.9826, 240.9124, 231.0428, 227.2079, 234.9389, 251.1798, 255.4991, 
    256.2188, 257.7749, 261.2321, 261.7845, 254.1542, 246.3024, 237.5173, 
    233.2184,
  239.3361, 244.0801, 242.8588, 236.8583, 234.0979, 238.8165, 251.7926, 
    251.9655, 256.0924, 256.6736, 256.7635, 250.2411, 241.3942, 232.2763, 
    227.5277,
  236.2406, 243.0542, 247.8731, 242.3559, 240.2651, 236.0866, 233.8911, 
    247.6239, 250.9033, 252.2001, 248.4915, 240.0048, 233.5392, 229.4776, 
    220.2931,
  232.3475, 238.8062, 244.7953, 245.5055, 244.9845, 236.3391, 233.8716, 
    239.4512, 239.0827, 241.1247, 236.1748, 233.8404, 231.6753, 219.5702, 
    206.0323,
  230.8199, 233.2981, 239.7125, 243.5641, 246.5573, 240.6917, 226.6324, 
    227.4739, 226.3906, 221.5511, 222.1232, 217.8808, 208.3131, 200.6836, 
    197.6695,
  231.054, 232.0509, 232.4479, 237.0314, 242.8802, 236.1645, 231.0806, 
    215.1233, 210.0235, 210.5607, 216.6667, 203.6598, 204.6252, 193.285, 
    197.6263,
  234.3469, 232.1318, 231.9555, 228.8881, 234.8873, 240.119, 231.0613, 
    224.5971, 215.6579, 208.6192, 204.4021, 201.7581, 198.7572, 199.2143, 
    205.2776,
  228.0531, 234.0722, 229.9683, 227.7948, 226.0086, 230.1396, 228.8205, 
    220.0034, 218.578, 206.0552, 202.7228, 201.9255, 198.572, 206.432, 
    214.3148,
  218.6391, 222.033, 229.6054, 228.4372, 223.6263, 222.3635, 220.2063, 
    219.9726, 214.424, 206.3552, 203.0524, 200.1641, 208.5983, 215.2362, 
    218.3646,
  199.4574, 196.2631, 205.8965, 224.5815, 231.6651, 237.8209, 241.0139, 
    249.6678, 258.5923, 267.5862, 260.2731, 258.7933, 258.4945, 250.506, 
    242.7901,
  206.2025, 196.2026, 202.1923, 211.999, 227.7428, 233.7495, 236.4157, 
    246.5838, 255.9561, 258.7852, 261.5283, 249.5561, 251.4442, 253.4894, 
    244.0687,
  215.5177, 204.4455, 202.6072, 203.1171, 214.1984, 230.2126, 231.9119, 
    238.8033, 251.7061, 256.9734, 260.0964, 251.3588, 252.7532, 247.7598, 
    245.8393,
  230.4947, 221.1936, 208.4865, 206.698, 206.695, 220.9369, 229.4225, 
    233.3229, 240.7299, 250.9642, 256.3381, 258.2939, 255.2235, 249.6363, 
    245.5338,
  233.5878, 232.5072, 225.9369, 218.762, 208.4444, 214.3677, 228.6588, 
    239.3191, 240.7887, 238.8799, 244.7499, 255.0328, 256.5784, 247.378, 
    234.9985,
  235.191, 235.2614, 233.9913, 233.7472, 226.7883, 218.6109, 224.0387, 
    232.1074, 232.4911, 232.3521, 235.0929, 244.7783, 245.0095, 241.3215, 
    232.5254,
  237.2952, 235.9469, 235.4522, 234.0896, 238.4949, 231.3897, 232.2364, 
    228.1475, 229.4622, 233.5252, 230.7104, 231.5676, 233.2157, 228.211, 
    219.4315,
  236.3364, 238.4751, 236.0143, 236.4175, 240.037, 241.9161, 241.7447, 
    238.6165, 235.192, 233.5356, 226.6246, 229.0442, 227.0808, 217.2172, 
    206.5611,
  218.689, 236.3264, 235.59, 235.2948, 239.971, 241.1875, 245.9939, 245.8584, 
    241.0977, 236.0215, 229.6567, 223.81, 216.1125, 210.8925, 200.01,
  214.5515, 224.4139, 229.4468, 235.4197, 238.2397, 239.723, 243.6559, 
    246.079, 245.4543, 238.2042, 230.0175, 220.2011, 208.1238, 203.2844, 
    195.227,
  180.5534, 206.145, 217.0072, 236.3246, 240.2831, 241.8218, 239.9564, 
    240.456, 248.3438, 264.117, 271.6079, 268.5232, 264.1258, 266.8839, 
    263.7141,
  176.4645, 191.6134, 209.7929, 230.2965, 231.1637, 235.812, 236.4314, 
    239.9538, 250.5803, 264.1349, 269.5805, 267.4523, 267.0102, 266.2644, 
    264.7225,
  177.8796, 180.3837, 200.2013, 217.6124, 231.7065, 232.2059, 231.7889, 
    232.875, 242.0522, 257.3746, 259.4128, 264.0154, 266.0686, 264.2179, 
    260.7179,
  184.5273, 179.2676, 189.5608, 208.3917, 222.5415, 229.6392, 228.1015, 
    230.1653, 233.1365, 249.3527, 247.1602, 257.3311, 262.7585, 265.7847, 
    264.9785,
  198.9484, 186.8194, 184.3707, 194.4436, 212.0589, 222.4718, 227.1492, 
    235.8223, 239.4034, 240.842, 240.189, 248.1551, 254.6402, 259.6753, 
    259.3092,
  213.0233, 200.2903, 193.5917, 194.5337, 198.1615, 210.9357, 220.2358, 
    225.3418, 221.5576, 229.5344, 238.7223, 238.9492, 245.6209, 246.1876, 
    248.195,
  226.2997, 216.5899, 207.0754, 198.6653, 200.4409, 205.248, 212.2786, 
    216.8391, 220.3189, 232.2978, 235.0058, 237.7464, 239.1866, 237.1599, 
    238.9479,
  242.8565, 226.9958, 223.2535, 212.2184, 209.418, 207.8299, 211.9664, 
    216.9185, 222.3967, 230.5937, 229.4084, 233.5357, 233.2316, 234.0868, 
    225.9381,
  247.1685, 237.6983, 233.5363, 225.0871, 218.6576, 213.1272, 215.954, 
    220.2624, 221.093, 223.232, 225.6859, 229.8079, 228.3624, 225.0717, 
    220.0718,
  235.0833, 231.0002, 230.5333, 234.0062, 228.4597, 223.2594, 222.0407, 
    224.703, 226.5773, 228.2859, 231.3071, 232.7978, 226.1349, 221.107, 
    215.2145,
  236.6359, 248.2789, 250.5479, 242.136, 249.3474, 247.4157, 229.5436, 
    222.0291, 238.5788, 270.042, 274.7439, 271.9362, 273.7631, 273.1014, 
    275.0076,
  225.7246, 242.9617, 249.8186, 248.0169, 253.5615, 249.5029, 230.4604, 
    218.1282, 229.1107, 261.9495, 274.9818, 272.3704, 264.2052, 272.052, 
    273.7268,
  218.2738, 231.9518, 246.3734, 246.4992, 252.0228, 244.1496, 229.0929, 
    215.3479, 216.1566, 245.6367, 269.1483, 263.6473, 257.9081, 262.4837, 
    264.7911,
  208.7031, 222.7514, 234.868, 240.2073, 244.6761, 241.9828, 223.3072, 
    217.3318, 215.6174, 235.9465, 252.4947, 262.6743, 262.5494, 261.6198, 
    268.0125,
  196.1335, 206.2195, 223.8137, 233.8872, 237.706, 231.2299, 228.0385, 
    219.2542, 223.8217, 228.8947, 246.8255, 254.7131, 260.5304, 263.2678, 
    262.601,
  190.92, 199.058, 212.7715, 226.1349, 229.9642, 228.1145, 218.9417, 
    213.4656, 214.7299, 225.6483, 237.5632, 239.7039, 246.0636, 254.9085, 
    259.9293,
  201.8233, 196.5874, 205.2793, 218.4914, 222.309, 221.7664, 221.439, 
    213.8795, 213.0959, 220.0217, 226.3548, 228.8249, 232.69, 242.2185, 
    244.6257,
  207.87, 199.3625, 202.9152, 211.03, 218.3318, 216.6996, 223.1269, 216.4991, 
    216.0521, 218.9584, 217.6285, 222.9943, 223.1917, 226.0767, 231.6519,
  228.1712, 212.9107, 204.2232, 206.5377, 212.6403, 216.1958, 216.9594, 
    214.8454, 214.985, 216.1362, 216.9462, 222.6511, 222.3151, 221.1282, 
    228.2869,
  244.8583, 234.3861, 216.1891, 211.1723, 213.8547, 212.0585, 209.6662, 
    210.8457, 212.0568, 212.0336, 220.498, 216.7249, 224.8115, 218.9094, 
    224.8608,
  220.5218, 234.2147, 238.0629, 240.9611, 249.3366, 229.2299, 209.1154, 
    202.0933, 226.3521, 264.2501, 278.97, 274.9008, 276.8175, 275.1948, 
    275.2541,
  213.9538, 237.5028, 242.0008, 235.5128, 249.105, 230.1906, 213.1585, 
    202.7149, 226.6689, 263.1315, 277.7831, 270.7949, 268.3537, 275.0404, 
    275.4844,
  209.0927, 239.1858, 236.7117, 236.0597, 248.0198, 224.0719, 218.3327, 
    202.8442, 229.896, 257.9935, 266.0493, 267.5958, 261.3578, 267.0197, 
    266.7899,
  207.3985, 236.1906, 234.4105, 236.4064, 242.3868, 226.8712, 223.0081, 
    212.7579, 232.9366, 250.4554, 260.1165, 261.3156, 261.8705, 263.3888, 
    264.009,
  205.1525, 231.6814, 233.6273, 235.5393, 242.1454, 221.8463, 226.8334, 
    221.7347, 235.961, 248.2565, 260.9196, 261.5734, 261.2706, 264.0983, 
    264.6234,
  207.6431, 217.5871, 234.5968, 235.1007, 240.499, 225.0429, 223.1901, 
    219.075, 228.7648, 239.8624, 261.5081, 261.2874, 263.2581, 259.1862, 
    259.3053,
  215.031, 209.7635, 228.2228, 236.9808, 234.588, 228.5337, 230.1569, 
    217.3597, 221.6606, 236.4857, 253.7704, 259.5526, 261.2688, 259.3016, 
    253.7011,
  208.1229, 203.419, 216.7387, 224.725, 227.5204, 231.6075, 232.8396, 
    228.3263, 232.2803, 234.4052, 243.0382, 254.4297, 260.6484, 261.1338, 
    253.4228,
  217.596, 222.3463, 212.1731, 221.7749, 225.049, 227.9713, 234.1797, 
    232.3124, 229.856, 233.4745, 237.459, 249.9227, 258.759, 257.1741, 
    250.3958,
  234.5631, 222.1236, 222.445, 223.3408, 221.6558, 223.957, 238.2709, 
    241.2001, 239.476, 231.3938, 236.3692, 236.8792, 243.6516, 246.1664, 
    247.5103,
  231.8349, 234.5791, 237.318, 239.4944, 241.7964, 246.7532, 242.7123, 
    226.749, 222.9822, 250.8469, 272.0692, 273.4205, 268.3123, 246.4048, 
    220.1726,
  228.7959, 233.6604, 237.0271, 238.2746, 242.7077, 246.11, 243.7751, 
    227.7037, 229.7536, 249.9338, 271.118, 268.5411, 259.8788, 227.378, 
    227.593,
  229.7797, 233.5297, 235.6644, 236.9028, 239.8439, 238.8383, 242.6461, 
    226.6886, 228.3225, 249.6333, 261.951, 262.8384, 247.5019, 226.7992, 
    245.1722,
  225.0059, 233.2863, 234.4145, 236.1016, 235.7523, 240.9745, 231.8621, 
    229.8366, 236.3062, 251.9511, 258.4194, 252.214, 238.944, 231.6497, 
    258.1149,
  224.2922, 230.9673, 233.4681, 233.5255, 234.2545, 230.6581, 230.3495, 
    227.8952, 236.8182, 252.2173, 259.8015, 250.4752, 238.1498, 250.778, 
    260.472,
  221.5782, 229.5214, 232.8731, 232.5379, 233.0382, 228.0345, 219.965, 
    222.495, 239.4569, 256.165, 260.3333, 248.584, 242.8983, 255.8011, 255.423,
  221.7128, 225.5606, 231.6822, 234.6011, 232.093, 226.1994, 215.505, 
    215.5064, 238.8571, 260.5901, 257.4875, 250.1138, 249.4276, 251.376, 
    251.1192,
  216.9063, 221.5029, 225.6393, 234.1361, 232.362, 220.0513, 214.1118, 
    220.7338, 242.8821, 260.5422, 256.7117, 249.489, 253.1091, 246.7889, 
    246.824,
  218.0034, 216.1636, 223.9857, 229.7669, 228.6614, 218.6678, 212.7885, 
    217.6864, 242.2143, 260.0143, 259.1034, 254.8306, 251.7899, 251.8527, 
    242.3656,
  224.3624, 220.6311, 217.7755, 224.4346, 223.5302, 213.9463, 214.185, 
    219.0167, 239.4806, 258.6704, 256.6684, 255.0825, 251.3847, 245.5486, 
    246.7536,
  252.9655, 245.5742, 240.2141, 239.973, 239.041, 239.1818, 238.8331, 
    237.2494, 239.8116, 246.0832, 251.8342, 256.5992, 253.1906, 251.9265, 
    267.1861,
  240.86, 241.6926, 239.7943, 241.6694, 240.4916, 240.4405, 239.9438, 
    240.7859, 239.3145, 243.8773, 249.942, 255.1837, 253.7054, 254.2996, 
    264.7396,
  236.008, 235.1404, 237.6151, 240.0407, 242.3601, 239.7492, 242.1114, 
    242.2669, 240.9411, 242.2352, 248.5983, 254.797, 252.4426, 251.0022, 
    260.546,
  233.4656, 231.4221, 236.4257, 237.3183, 239.6095, 242.8121, 239.7907, 
    247.706, 245.7859, 241.9763, 249.0771, 252.8597, 250.6115, 252.0663, 
    257.4886,
  234.4327, 231.6933, 234.1728, 235.553, 237.0779, 240.6003, 243.5789, 
    240.7199, 244.1689, 239.2489, 243.8742, 249.3222, 249.7109, 253.69, 
    254.5539,
  228.241, 230.3715, 231.7026, 232.9852, 236.389, 238.1664, 241.7514, 
    245.3586, 246.1267, 236.246, 238.4616, 242.7088, 251.9364, 254.0342, 
    254.0432,
  223.9172, 224.5577, 223.7686, 226.2202, 231.0787, 236.5314, 241.0754, 
    244.8923, 246.0559, 241.7884, 229.6226, 234.3433, 250.956, 256.4683, 
    253.9469,
  223.8476, 216.9578, 219.9807, 226.7954, 230.8822, 235.9021, 238.6861, 
    246.2643, 248.0165, 242.9058, 227.0118, 236.7857, 254.2268, 257.4297, 
    253.6717,
  217.7197, 215.5569, 217.3441, 217.8736, 225.2115, 234.9481, 239.7014, 
    244.3854, 249.6075, 244.9194, 229.1452, 234.5172, 253.8214, 258.1422, 
    253.8985,
  218.8631, 216.9656, 216.6229, 216.5639, 229.1513, 236.6265, 241.7434, 
    247.6663, 250.7118, 244.0954, 225.8888, 228.758, 252.5748, 254.8409, 
    251.7384,
  234.205, 232.8179, 240.9131, 239.9978, 240.1906, 239.6878, 237.7355, 
    236.4928, 239.2634, 242.7151, 241.9993, 245.3641, 238.2394, 230.4248, 
    238.2418,
  238.8893, 238.8347, 239.4315, 238.2801, 240.3382, 241.5369, 241.0527, 
    238.6052, 239.7303, 238.9651, 245.6306, 243.4711, 234.9494, 231.5994, 
    240.4377,
  233.4594, 240.0672, 241.8719, 238.738, 239.1457, 238.597, 244.5452, 
    239.1143, 241.7387, 240.8024, 245.1597, 245.9566, 231.5506, 225.7306, 
    231.7396,
  228.3762, 229.2777, 238.2759, 241.572, 238.5106, 238.9854, 238.0906, 
    244.2261, 246.6004, 241.0512, 241.3476, 242.1944, 229.9107, 226.8819, 
    234.3665,
  244.1967, 243.028, 237.0155, 238.8395, 238.6758, 237.3685, 238.4566, 
    239.3843, 238.8495, 239.5332, 239.6086, 245.3059, 237.7821, 227.5367, 
    229.9864,
  239.2871, 235.579, 231.3354, 230.2606, 234.6837, 239.8602, 240.842, 
    239.9614, 239.8961, 240.1958, 235.1825, 243.7505, 240.6444, 228.5412, 
    221.5841,
  227.8252, 228.5731, 228.2935, 230.5475, 229.2736, 230.1884, 234.2422, 
    238.0889, 241.9276, 240.8187, 238.543, 240.1321, 248.8992, 236.0924, 
    219.6272,
  229.0299, 229.8016, 229.0027, 230.1527, 229.742, 230.0505, 232.9888, 
    240.861, 241.4668, 241.3854, 239.6404, 238.6757, 247.742, 245.184, 227.952,
  233.36, 231.7883, 230.3364, 229.8862, 226.8472, 225.2549, 230.4318, 
    236.3889, 241.3778, 243.5217, 241.1802, 237.9205, 243.5052, 250.3836, 
    238.6144,
  235.6463, 228.9053, 228.3373, 229.5976, 226.6281, 227.1329, 229.5943, 
    235.0193, 238.9756, 242.1906, 242.0661, 236.5254, 242.9973, 250.2889, 
    244.1418 ;

 scalar_axis = 0 ;

 sftlf =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.141347, 0.07456003, 0.2762221, 0, 0.2154952, 0.5089986, 0.007178012, 0, 
    0.1467785, 25.31165, 20.60715, 2.120196, 15.979, 48.81725, 63.64272,
  0.001503375, 0, 0, 0, 0.8848332, 11.68672, 0, 0, 0, 0.4694104, 0.9680001, 
    0.09868675, 1.334438, 150.908, 101.0153,
  0, 0, 0, 0, 8.803595, 280.9762, 7.478715, 0, 0, 0, 0.0046135, 0, 
    0.00845787, 0.9458157, 6.678408,
  0, 0, 0, 0, 0, 12.95772, 307.1121, 15.76765, 0, 0, 0, 0, 0.001950179, 
    0.08926713, 2.882818,
  0, 0, 0, 0, 0, 0, 9.245329, 485.3841, 540.1508, 15.00115, 0.01623012, 0, 0, 
    0.06344586, 0.01027276,
  0, 0, 0, 0, 0, 0, 0, 1.278773, 12.13823, 0.8518202, 0.2699268, 0, 0, 
    0.01012854, 0.01599434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05785002, 0, 0, 0, 0, 0.2725836,
  0, 0, 0, 0, 0, 0, 0, 0.3482242, 1.154397, 3.605569, 0.8750445, 0, 0.158783, 
    0.02233585, 0.6264485 ;
}
