netcdf atmos.1980-1981.aliq {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 11:53:49 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.nc reduced/atmos.1980-1981.aliq.nc\n",
			"Mon Aug 25 14:39:17 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -6.136523e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.254924e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.112337e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.07579e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 2.890782e-05, 0, -1.363373e-06, 0, 0, 0, -9.73065e-08, 0, 0, 
    2.526224e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.1657e-06, 0, 0, 0, 0,
  0, 0, 0, -3.880526e-07, 0, -2.098912e-07, -1.469291e-06, 0, 0, 
    -2.442881e-07, -9.019695e-07, 0, 4.371262e-05, 0, 5.485918e-06, 
    -6.187642e-11, 0, 0, 0, 0, 0, 0, 0, 0, -1.352705e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -4.484093e-07, 2.405397e-06, 0, -3.350173e-07, 
    -5.324855e-07, 0, -3.569248e-07, 0, 0, 0, 0, 0, 0, 0, 0, -2.064459e-07, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 3.438136e-05, 5.870911e-05, 1.494414e-05, 0, 
    -2.481991e-06, 0, 0, 0, 0, 0, 0, -2.141107e-07, -1.236259e-06, 0, 0, 
    2.564439e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -2.738298e-06, 6.504583e-05, -1.99626e-07, -8.337548e-08, 
    8.119186e-06, 8.997665e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 7.503704e-07, 0.0002950877, 6.573232e-06, 3.551227e-05, 0, 
    -1.248489e-06, -6.020026e-07, -2.398529e-06, -8.059528e-07, 5.642353e-06, 
    7.741545e-05, 1.833506e-05, 2.857688e-05, -2.373882e-07, 0, 5.874296e-07, 
    0, 0, 0, 0, 0, 0, -4.055553e-06, 0, 0, 0, 0,
  0, 0, 3.678203e-06, -4.108795e-06, -3.023277e-06, 3.262934e-05, 
    -4.407873e-06, 2.347701e-06, 1.303532e-05, -2.977098e-06, 2.202641e-05, 
    1.095381e-05, 9.218875e-05, -5.838169e-06, 0.000134762, -2.232185e-06, 0, 
    -1.240803e-07, 0, 0, 0, 0, 0, -1.42364e-06, -5.332435e-06, 1.055829e-05, 
    0, 0, 0,
  0, 5.776115e-06, -1.435026e-06, 0, 1.091255e-06, 1.103804e-06, 0, 
    -3.38519e-07, -1.19904e-06, 8.18146e-05, -2.455446e-06, -2.345127e-06, 
    5.312474e-05, 2.562815e-07, 5.184525e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -8.718501e-07, 7.889109e-09, 0, 0, -2.656939e-07, 0,
  0, 0, 0, 0, 0, 0, 0, 5.164693e-05, -2.219964e-06, 6.709639e-05, 
    0.0002452189, 3.316299e-05, 0.000122059, 8.421825e-05, -1.138004e-06, 0, 
    -1.163189e-06, -1.115705e-06, 0, -1.733143e-07, 4.259954e-05, 
    3.730318e-05, 5.406658e-05, 1.038775e-06, 5.325181e-05, 0, -3.750349e-07, 
    0, 0,
  0, 0, 0, 0, 0, 0, 1.017189e-05, 8.394452e-05, -1.232763e-06, 1.155462e-05, 
    0.0003449228, 0.0002504748, -1.494427e-06, 0, 0, 0, 0, 0, 0, 0, 
    -6.196097e-07, 0, -1.352211e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.707784e-06, 6.659714e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 8.577484e-05, 0, 0, 0, 0, 9.370727e-05, 0, 0, 0, 0, 0, 0, 
    -5.228511e-07, 0, 0, 0, 0, 0, 0, 0, 0, -1.07831e-07, 0, 0, 0,
  0, -9.184159e-07, 3.317356e-06, 0.0004956687, 1.5732e-05, 0.0001924253, 0, 
    0.0001390938, 6.078876e-05, 1.160524e-05, -6.348633e-07, 9.894445e-05, 
    0.0001589483, 0.0001425175, 0.0001107694, -5.496449e-06, 0, 1.23889e-05, 
    0, 0, 0, 0, 0, -7.489882e-09, 7.272392e-05, 3.026143e-05, 0, 0, 0,
  0, 0, 0.0001426013, -4.690183e-06, 7.206705e-05, 0.0001439939, 
    -1.815477e-05, 0.0001994687, 0.0001650703, 8.869915e-06, 0.0001329719, 
    6.860141e-05, 0.0002286307, 1.881084e-05, 0.0003995104, 0.0003442488, 
    2.192732e-06, -1.461065e-06, -7.200829e-07, 0, 0, 0, 0, 5.137535e-06, 
    9.174056e-05, 8.494688e-05, 0, 0, 0,
  -5.342646e-07, 0.0001581547, 8.494599e-06, 0, 3.271409e-06, 0.0003439685, 
    8.917954e-06, -1.068209e-06, -1.253525e-06, 0.0002782514, 2.08821e-05, 
    -5.529619e-06, 0.0003094958, 0.0001107501, 9.700518e-05, -1.846361e-08, 
    -5.735412e-07, 0, 0, 0, 0, 0, 0, 2.67135e-05, 3.162188e-05, 9.250919e-05, 
    1.748167e-05, -6.372564e-07, 0,
  -1.668654e-07, -3.371535e-07, 0, 0, 0, 0, -7.020166e-07, 0.0002652147, 
    6.491068e-06, 0.0002681242, 0.0009567462, 0.0001146483, 0.0005508801, 
    0.000357464, 5.427959e-05, 0.000142649, 0.0002197675, 6.065584e-05, 
    1.008535e-05, -8.096215e-06, 0.00039081, 0.0004243999, 0.0002340823, 
    3.825703e-06, 0.0001484415, -4.144323e-07, 5.297301e-05, 1.722141e-05, 
    -9.241738e-07,
  0, 0, 0, 0, 0, 0, 0.0005294149, 0.0001667399, -3.657828e-06, 8.476552e-05, 
    0.0009956262, 0.0005427265, -1.305608e-05, 1.260862e-05, 0, 0, 0, 0, 0, 
    0, -7.684181e-06, 4.057306e-05, -4.254083e-06, 2.675333e-05, 
    -2.69497e-07, -2.004228e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.091068e-05, 0.0001675732, 1.189526e-05, 
    -1.791452e-06, 2.316095e-07, 1.316746e-05, 0, 0, 0, 0, 0, 0, 0, 
    -2.609174e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.020382e-07, 1.807498e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 1.724251e-05, 0, -8.329946e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.736471e-06, 0, 0, 0, 0,
  0, 0, 0, -2.963954e-07, 0.0003171631, -3.041313e-06, -2.827647e-06, 0, 0, 
    0.0002107495, 0, -1.360409e-09, 2.666623e-05, -5.499271e-07, 0, 
    -2.337353e-06, -7.063715e-06, 0, -1.315572e-07, -5.295728e-07, 0, 0, 0, 
    0, -2.08179e-06, -6.365056e-06, -2.941194e-06, 0, 0,
  0, -3.926499e-06, 2.941714e-05, 0.0008299379, 0.0001793485, 0.0003494378, 
    6.67296e-06, 0.0003154779, 0.0002723942, 0.0002038245, 9.246691e-05, 
    0.0001890401, 0.0003310167, 0.0003392776, 0.0002137039, 1.762804e-05, 
    -1.72545e-05, 2.270096e-05, 0, 0, 0, 0, 0, -2.246964e-08, 0.0002602255, 
    0.0002733522, -6.678434e-06, 0, 0,
  0, 5.01867e-05, 0.0002565707, 2.598505e-05, 0.0002237189, 0.0005915824, 
    0.0002790524, 0.000493695, 0.0004585033, 7.953632e-05, 0.0002514192, 
    0.0001431833, 0.0008781581, 0.0003580261, 0.0009799293, 0.0009516105, 
    9.482446e-05, 1.83813e-05, 3.599413e-05, 0, 0, -8.872264e-07, 0, 
    0.0001174445, 0.0003682391, 0.0002885363, 0, 0, 0,
  4.297304e-05, 0.0004943172, 0.0001009272, 0, -6.8501e-06, 0.0007786419, 
    0.0002435575, 0.0001698735, 2.65178e-06, 0.001060063, 0.0002783139, 
    -5.016048e-06, 0.0008929409, 0.0004842205, 0.0004093527, 2.822535e-06, 
    -3.827251e-06, -4.092311e-06, 0, 0, 0, 1.323655e-06, 0, 0.0001381651, 
    0.0001917006, 0.0002370895, 0.0001215593, 1.011294e-06, -7.27245e-07,
  -2.967214e-06, 4.602592e-06, 8.899287e-06, -1.122827e-06, 0, -1.569241e-06, 
    -9.274698e-06, 0.001025568, 0.0001702495, 0.0007295532, 0.001782796, 
    0.0006837462, 0.002069508, 0.001282519, 0.0001392881, 0.0003349575, 
    0.0009254793, 0.0004559935, 0.0001659405, 0.0002157636, 0.001288342, 
    0.001380655, 0.0005713395, 1.392867e-05, 0.0003481515, 1.469701e-05, 
    0.0002505122, 0.0002894198, 0.0003256046,
  0, 0, 0, 0, 0, -5.691844e-07, 0.001419445, 0.0004255939, 3.196565e-05, 
    0.0002402475, 0.002074744, 0.001408782, 4.564977e-05, 0.0004235335, 0, 0, 
    0, 0, 0, -7.255049e-08, 1.372259e-05, 3.905788e-05, 6.08562e-06, 
    0.0004891404, 7.164566e-06, 3.048695e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 1.656879e-05, 3.409945e-05, 0.0003654582, 8.700965e-05, 
    2.875435e-05, 9.240842e-06, 4.05727e-05, 0.0001080675, -9.248015e-07, 0, 
    0, 0, 0, 0, -4.591958e-06, 0, 5.658536e-06, 3.039131e-05, 0, 
    -3.003171e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.306507e-09, -3.596205e-10, 1.748223e-06, 
    7.2137e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.409656e-08, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0.0001704271, -1.327984e-07, 2.966957e-05, 0, 0, 0, 0, 0, 0, 0, 
    -1.540976e-09, -3.107326e-07, 0, 6.312802e-06, 8.065216e-06, 0, 0, 0, 0, 
    0, 0, 9.277543e-05, -3.611995e-07, 6.740362e-05, 0, 0,
  0, 0, -2.522866e-07, -4.132077e-06, 0.0006778809, 2.107059e-05, 
    2.47566e-05, 0, 0, 0.0003254187, 0, -2.720818e-09, 6.648435e-05, 
    7.721877e-06, 5.728129e-06, 1.348536e-05, 6.775105e-05, 0.0001246088, 
    0.0001620586, -8.619948e-07, 0, 0, 0, 0, 3.828285e-05, -8.539814e-06, 
    4.27217e-05, 0, 0,
  0, 9.177459e-06, 0.0001972107, 0.00105605, 0.0006732337, 0.0007931656, 
    0.0003963389, 0.0005681839, 0.0003516976, 0.0005117054, 0.0002014638, 
    0.0002589175, 0.0008298442, 0.0006588857, 0.000590889, 0.0001453266, 
    9.885717e-05, 5.943449e-05, -3.421782e-07, 0, 0, 0, 0, -2.48834e-07, 
    0.0008345377, 0.0007289079, 2.980853e-05, 0, 0,
  0, 0.0003661683, 0.0008327896, 0.0002805041, 0.0006336261, 0.001390886, 
    0.0009207246, 0.001221467, 0.001253643, 0.0001480883, 0.0009876954, 
    0.0004518909, 0.002597143, 0.001321092, 0.002119505, 0.001773714, 
    0.0003539632, 0.0001686148, 0.0002056107, 0, 0, -2.939039e-06, 0, 
    0.0005478273, 0.001091852, 0.00058451, 8.76635e-06, 0, 0,
  6.535755e-05, 0.001107685, 0.000426668, 0, 0.000242057, 0.001554085, 
    0.0005218964, 0.0003304349, 7.232199e-05, 0.002452794, 0.0008237893, 
    7.481519e-05, 0.00264707, 0.002011803, 0.001939775, 9.567744e-06, 
    -6.809771e-06, -5.876599e-06, -1.868844e-06, 0, 0, 3.68767e-06, 
    4.216752e-05, 0.000624178, 0.0005596134, 0.0007230112, 0.0005377269, 
    3.548472e-07, -1.617175e-06,
  1.311839e-05, 2.656939e-05, 0.0001605735, -4.317396e-06, 7.703851e-06, 
    -4.804549e-06, 5.416795e-05, 0.001659907, 0.0006312084, 0.001716063, 
    0.002877794, 0.002108308, 0.0056289, 0.003371631, 0.0005593617, 
    0.00132357, 0.001914201, 0.001469685, 0.0008632492, 0.00147183, 
    0.004068576, 0.00320254, 0.0013181, 1.801831e-05, 0.0006002401, 
    8.894017e-05, 0.0007290103, 0.0008542162, 0.0007148745,
  0, 0, 0, -6.089145e-08, 9.967441e-06, 3.80504e-05, 0.00337791, 
    0.0008950551, 0.0005120909, 0.000964029, 0.004371686, 0.004463729, 
    0.0008216465, 0.001556018, -4.261071e-08, -1.454921e-06, 0, 
    -1.451668e-06, 3.654974e-05, -1.765992e-07, 5.921669e-05, 0.0001544945, 
    0.0001212044, 0.0008409012, 6.246007e-05, 0.0001292096, 0, 0, 0,
  0, 0, 0, 0, -1.006919e-06, 0, 0.0001233787, 9.779523e-05, 0.0009005829, 
    0.0003913871, 0.0005751671, 8.463401e-05, 0.0003584907, 0.0001959734, 
    2.540953e-05, -7.023448e-07, 0, 0, 0, 0, 1.006232e-05, 0, 5.354299e-05, 
    0.0002726744, 0, -3.661831e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 3.401807e-07, -2.723744e-08, 0.0001182114, 
    8.932687e-05, 0.0008991349, -2.043546e-06, 1.832464e-05, 0, 0, 0, 0, 0, 
    -1.548096e-06, 8.351838e-06, -9.885126e-07, 1.239656e-05, -7.395398e-07, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.046645e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.197431e-06, -9.167797e-07, 0, 2.942649e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.74035e-06, 0, 0, 0, 0, 0, 0, 
    -5.568836e-10, 0, 0, 0, 0, 0, -3.657907e-07, 0, 0, -2.355826e-08,
  0, 0, 0, 0.0005530587, 3.539032e-05, 0.0002187589, 1.107263e-06, 0, 0, 0, 
    2.400212e-05, -2.185013e-06, 1.912973e-05, 1.899109e-05, 4.001885e-05, 
    -6.18129e-07, 0.000107031, 4.521423e-05, 3.066501e-05, 5.741805e-06, 
    5.20765e-06, 1.038787e-05, 0, 0, 0.0002946829, 0.0001619768, 
    0.0001998958, 1.329103e-05, 0,
  0, 0, 1.294148e-06, 0.0001158753, 0.001592743, 0.0003305777, 0.0006634129, 
    0, 0, 0.0004540946, 0, -7.541312e-07, 9.335846e-05, 0.0002604975, 
    0.0005030183, 0.0001312878, 0.0005168456, 0.000609217, 0.0008830542, 
    2.564115e-05, 1.382155e-05, 0, 0, 0, 0.00012606, 0.00049513, 
    0.0004056936, 0, 0,
  0, 0.0001248539, 0.0003746988, 0.001646712, 0.002023178, 0.001727514, 
    0.0008175949, 0.001173379, 0.000531538, 0.0008974034, 0.0006200154, 
    0.0005798484, 0.00180675, 0.001339346, 0.001279764, 0.0008402365, 
    0.001018904, 0.0004657679, 4.50349e-05, -2.754692e-06, 0, 0, 0, 
    -1.117124e-06, 0.001501711, 0.00129261, 0.0001560761, 0, 0,
  0, 0.0006195923, 0.001470074, 0.0005995597, 0.001548421, 0.002753104, 
    0.002495732, 0.002669916, 0.00222946, 0.000340058, 0.001976425, 
    0.001281783, 0.004419104, 0.003436895, 0.00440711, 0.00374231, 
    0.001086673, 0.0004471324, 0.0006400002, 0, 0, -1.02136e-05, 0, 
    0.00127175, 0.002108463, 0.0009090472, 0.000163852, 0, 0,
  0.00023151, 0.002359767, 0.001399086, -7.823898e-07, 0.0009516035, 
    0.003123498, 0.001143803, 0.0009686664, 0.0008143578, 0.005030042, 
    0.002003646, 0.0002906602, 0.005593397, 0.00379673, 0.002926609, 
    0.0001383556, 3.456523e-05, -3.976455e-06, 2.079982e-06, 5.046678e-07, 
    -8.567859e-07, 1.707217e-05, 0.0002885859, 0.001472146, 0.001147707, 
    0.002072469, 0.001431425, 4.495174e-05, 1.72054e-05,
  0.0001047764, 0.0001447779, 0.0002225342, -7.393027e-06, 7.497873e-05, 
    -1.284955e-05, 0.0002146155, 0.002464583, 0.001635972, 0.00369725, 
    0.005101148, 0.004536056, 0.01131762, 0.007706775, 0.001521966, 
    0.002895426, 0.003585331, 0.004033749, 0.00254454, 0.003600027, 
    0.009125054, 0.006672204, 0.00266514, 0.0003060048, 0.0008523478, 
    0.0002187399, 0.001420468, 0.002071482, 0.001480836,
  0, 0, 0, 9.604516e-06, 1.437223e-05, 0.0001352738, 0.00643475, 0.001610239, 
    0.001165828, 0.002488324, 0.008722627, 0.008468685, 0.002394188, 
    0.003263271, -2.257011e-07, -3.606863e-06, -2.731078e-07, -1.030152e-06, 
    0.0002148007, -8.82941e-07, 0.0003722622, 0.0006037496, 0.0004809232, 
    0.00119117, 0.0002450455, 0.0002857512, -7.16314e-07, 0, 0,
  0, 0, -1.055742e-07, -6.313507e-07, 5.194396e-06, -3.673462e-07, 
    0.0002559491, 0.0005119753, 0.002083299, 0.001382562, 0.002266347, 
    0.0005385517, 0.001069244, 0.0005319701, 9.065601e-05, -4.885811e-06, 
    -4.685378e-07, 1.519798e-05, 0, 0, 3.417875e-05, -9.116515e-06, 
    0.0002147972, 0.0004543419, 8.114241e-06, 0.000100424, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.417464e-06, 9.222049e-06, 0.0002784311, 
    0.0005921028, 0.0005967675, 0.002275918, 0.0002701228, 1.995869e-05, 
    3.693151e-05, 0.000100257, 0, 0, 0, 1.981394e-05, 0.0004095865, 
    -8.435877e-06, 0.0003264569, -6.713735e-06, 1.203623e-06, -1.294568e-07, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.719081e-06, 9.543392e-06, -7.314091e-07, 
    2.745764e-05, -7.519798e-07, 3.508489e-06, -1.477844e-06, 0, 0, 0, 0, 
    5.379316e-05, 7.357423e-05, 2.722508e-05, 8.28949e-05, -2.520851e-09, 
    1.063453e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.08014e-07, 0, -1.761243e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -8.020239e-08, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -6.523547e-07, 0, 0, 0, 0.0001106319, 0, -1.555618e-06, -5.145332e-06, 0, 
    0, 0, 1.985493e-06, 0.0001534767, -6.560345e-06, 3.324759e-05, 
    -6.594778e-09, 0, -1.373221e-06, 0, 5.867633e-07, 0, 0, 0, 0, 
    -4.090195e-07, -3.131351e-06, 1.344226e-05, 3.186315e-06, -7.067477e-08,
  -4.228522e-07, 0, 4.616621e-06, 0.001117109, 0.0006449802, 0.0008436373, 
    5.090532e-05, 0.0001852774, 0, 1.716944e-06, 9.499039e-05, 0.000118913, 
    0.0003337985, 0.0002367513, 0.0001428823, 6.002776e-05, 0.0003699639, 
    0.0008372444, 0.0004560695, 0.0001844314, 0.0002921715, 0.0002858021, 0, 
    0, 0.001197765, 0.001299998, 0.00114457, 0.0002972772, 0.0001406412,
  0, 0, 1.78276e-05, 0.0008374591, 0.003614143, 0.0009770035, 0.001828333, 0, 
    3.696328e-06, 0.0005338635, 3.679092e-05, 3.729444e-05, 0.0002089859, 
    0.0008390543, 0.001605367, 0.001019725, 0.001597882, 0.001332913, 
    0.001699351, 0.0006278917, 0.0001481953, -2.124993e-06, 0, 0, 
    0.0003927651, 0.002118153, 0.001748796, 4.908239e-05, 1.322301e-06,
  0, 0.0003746499, 0.0006781602, 0.00265722, 0.004752352, 0.003198935, 
    0.001912846, 0.001906082, 0.0009032017, 0.001651079, 0.0017092, 
    0.001280139, 0.003580673, 0.00222881, 0.00305713, 0.002771851, 
    0.002480837, 0.001319176, 0.0002975092, 4.418721e-05, 1.605956e-05, 0, 0, 
    -2.948845e-06, 0.002620221, 0.002584231, 0.0006019713, 0, -3.075131e-07,
  0, 0.001232438, 0.003075391, 0.001111935, 0.003066073, 0.004706974, 
    0.005393348, 0.006685759, 0.004475224, 0.0009914779, 0.003553786, 
    0.00231307, 0.00763555, 0.007419823, 0.00857169, 0.007473091, 
    0.002323869, 0.0007883844, 0.0009909426, 0, 0, 3.801477e-05, 0, 
    0.002351121, 0.003937921, 0.001402893, 0.0005337365, -2.047753e-07, 0,
  0.0006172475, 0.004573764, 0.002287549, 7.162255e-06, 0.001656964, 
    0.00627498, 0.002594777, 0.001875343, 0.002050057, 0.009282975, 
    0.0034794, 0.00131217, 0.01013539, 0.006653044, 0.005227296, 
    0.0006259062, 0.0002516474, 0.0001559167, 5.101951e-05, -8.170302e-07, 
    -8.060282e-07, 0.0002067844, 0.000584429, 0.003249074, 0.001960211, 
    0.003726829, 0.002656471, 8.82052e-05, 1.520847e-05,
  0.0003991086, 0.000607371, 0.0005806431, 0.0001215649, 0.0002364207, 
    9.250287e-05, 0.00077715, 0.00370325, 0.003695496, 0.007005259, 
    0.008635097, 0.009724697, 0.02039116, 0.01565365, 0.00389326, 
    0.006306727, 0.006860932, 0.00829106, 0.005972059, 0.007155154, 
    0.01678163, 0.01279954, 0.004563196, 0.0008534543, 0.001208812, 
    0.0008586552, 0.002463125, 0.00477772, 0.002854249,
  0, 0, 0, 9.450155e-05, 0.0001899637, 0.0006569762, 0.01247457, 0.003071135, 
    0.002556681, 0.005892169, 0.01637397, 0.01366411, 0.005714779, 
    0.005860002, 1.478171e-06, 2.634746e-05, -4.558051e-06, -2.368073e-06, 
    0.0006209114, -4.784982e-06, 0.0008893405, 0.001818957, 0.001114783, 
    0.001467368, 0.0008746001, 0.0007862495, 2.207742e-05, 0, 0,
  0, 0, 4.908174e-05, 2.582028e-05, 0.0001013146, 3.192154e-07, 0.0008478248, 
    0.001027507, 0.003978914, 0.003415901, 0.005777127, 0.002360191, 
    0.00313358, 0.00157114, 0.0005599211, 0.0001954659, 1.045506e-06, 
    0.0002824935, 4.825155e-05, 0, 0.0001305078, 7.659331e-05, 0.0006076663, 
    0.000936334, 0.0004296901, 0.0005120976, 9.059861e-05, 0, 0,
  8.822825e-06, 1.331907e-07, -5.104713e-08, 0, 1.666483e-05, 8.31736e-08, 
    -3.157996e-09, 0, 0.0001102654, 0.0003388412, 0.001705338, 0.003179912, 
    0.002198888, 0.004916097, 0.00151892, 0.0002149221, 0.000228399, 
    0.000376428, 0, 0, -1.367039e-07, 0.0002869709, 0.00163978, 0.000341356, 
    0.0008624825, 0.000929617, 0.0001605023, -3.138602e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.141574e-06, 6.882639e-06, -6.873171e-06, 
    0.000259788, 0.0001275415, 0.0001895357, 0.0002616679, 0.0002936381, 
    6.625299e-05, 1.931045e-07, 0, 0, 1.684173e-05, 0.0006213785, 
    0.0006171403, 0.001054159, 0.0003666456, 0.0003586794, 0.0001312712, 
    -2.133212e-06, 5.190518e-05,
  0, -2.768659e-06, -1.815782e-07, 0, 0, -8.59041e-07, 0, 0, 0, 
    -9.785707e-07, -2.628446e-07, 3.678967e-06, -4.148885e-07, 2.889638e-05, 
    -6.350252e-07, 8.402989e-06, 0, 0, 0, 0, -7.011287e-08, 0, 7.702161e-05, 
    -6.73963e-07, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2.463607e-06, 0, -3.676579e-07, 0, 0, 0, 6.744734e-07, 
    1.678001e-05, 0, -3.563049e-07, 0, 0, -2.345404e-06, 0, 0, 0, 
    1.372117e-06, 0, 0, 0, 0, 1.954465e-05,
  4.143469e-05, -3.480857e-07, 0, 3.517111e-05, 0.0007867372, 0.0002476617, 
    0.0001178488, 0.0003328889, 9.719568e-05, 0, 0, 7.977791e-05, 
    0.0006871722, 0.0003378867, 0.0002644071, 7.830388e-05, 2.258352e-05, 
    2.320132e-05, 7.090635e-05, 0.0003778881, 0.0001439769, 8.253221e-05, 
    0.0001098171, -7.343725e-07, -2.270129e-06, 0.0001770613, 0.0004344134, 
    0.0001941798, 3.549596e-05,
  -9.874597e-06, -3.447319e-06, 0.0001514136, 0.002333167, 0.002980775, 
    0.002433853, 0.0005981472, 0.0005806139, 0, 0.0001481829, 0.0004184357, 
    0.0009633349, 0.0009934161, 0.001496171, 0.0007674173, 0.0005039895, 
    0.002024844, 0.002209419, 0.002398085, 0.001018634, 0.001767344, 
    0.0007844559, 0.0001910598, 1.236491e-05, 0.003394892, 0.005229586, 
    0.003332033, 0.001116935, 0.000459313,
  0, -1.871113e-06, 0.0001306984, 0.002988101, 0.006907009, 0.002870082, 
    0.004347946, -4.88401e-06, 0.0001150436, 0.0006725478, 0.0004996513, 
    0.0005864348, 0.001043131, 0.00308318, 0.003364223, 0.004892586, 
    0.005237624, 0.003839108, 0.00458512, 0.001749674, 0.000712719, 
    -1.296282e-05, 0, 0, 0.002002365, 0.00772831, 0.005419146, 0.0002140737, 
    0.0001476207,
  0, 0.001031073, 0.001724576, 0.004198727, 0.01147402, 0.005356066, 
    0.003975668, 0.003184127, 0.001812141, 0.003440628, 0.003071745, 
    0.003059224, 0.006313806, 0.004163367, 0.006690084, 0.008516629, 
    0.006574722, 0.003710947, 0.0009337988, 8.143124e-05, 9.451068e-05, 0, 
    3.834121e-05, 0.000140997, 0.005852815, 0.004588706, 0.001770505, 0, 
    -3.26879e-07,
  0, 0.002609456, 0.006076861, 0.0025617, 0.008214037, 0.01055138, 
    0.01192866, 0.01349795, 0.00832222, 0.002096369, 0.006831108, 
    0.005157196, 0.01437181, 0.01759814, 0.01681903, 0.01335938, 0.005759994, 
    0.002103921, 0.001563072, -1.05309e-06, 0, 4.581339e-05, 0, 0.005175256, 
    0.008219271, 0.003424153, 0.00115317, -2.856992e-06, 0,
  0.001166489, 0.00788073, 0.003771036, 8.351752e-05, 0.003084504, 
    0.01102419, 0.006693865, 0.004513303, 0.004710669, 0.01566467, 
    0.006393429, 0.004753506, 0.0183473, 0.0146262, 0.01090944, 0.0014, 
    0.001053783, 0.0009506898, 0.0002579331, 3.823715e-05, 3.787539e-05, 
    0.0005446282, 0.001145332, 0.007667518, 0.004046369, 0.006696343, 
    0.004765177, 0.0003896506, 0.0004896134,
  0.001127878, 0.001211007, 0.001072179, 0.0006926605, 0.0003963627, 
    0.0003758955, 0.00167783, 0.006157731, 0.006257073, 0.01303682, 
    0.01583043, 0.02097237, 0.03497081, 0.0276664, 0.01018005, 0.01254976, 
    0.01333821, 0.01539428, 0.01198693, 0.01379655, 0.03131696, 0.02391619, 
    0.009490472, 0.002207221, 0.002053139, 0.003117478, 0.004071303, 
    0.01198901, 0.004634425,
  0, -8.766746e-11, -2.698084e-12, 0.0005419492, 0.0004459201, 0.001931812, 
    0.02031045, 0.007060154, 0.006931343, 0.01071053, 0.02706255, 0.0234556, 
    0.01259702, 0.01002304, 6.787185e-05, 7.361617e-05, 0.0001661586, 
    0.001124225, 0.00131329, 0.0002075796, 0.00250686, 0.004187691, 
    0.002651291, 0.002897572, 0.001901072, 0.001530713, 0.0003344943, 
    -3.256412e-07, 0,
  0, -2.37596e-06, 0.0001402759, 0.0001639003, 0.0002952855, 8.123909e-05, 
    0.002930449, 0.001973071, 0.007315648, 0.007189418, 0.01106071, 
    0.007442639, 0.008198305, 0.003678919, 0.0020943, 0.001054274, 
    0.0002977118, 0.001380105, 0.0003407518, 4.250385e-05, 0.0002991616, 
    0.0006663459, 0.002089112, 0.002415933, 0.001312442, 0.001381941, 
    0.0005187849, 0, 0,
  0.0001198648, 8.884456e-05, 6.22383e-05, -6.62701e-09, 0.0001594535, 
    0.0001520294, 3.651422e-05, -1.043332e-08, 0.0005301666, 0.00119506, 
    0.004487136, 0.007576888, 0.007350487, 0.009361882, 0.004979472, 
    0.00186339, 0.00096875, 0.0006320179, -5.847705e-07, -2.638969e-06, 
    -1.200735e-06, 0.001750628, 0.004382414, 0.002062509, 0.003097323, 
    0.003483057, 0.0005522863, 5.690746e-05, -1.092326e-06,
  2.909038e-05, -8.052545e-07, 5.074234e-06, 1.064616e-05, 4.891867e-05, 
    1.077845e-05, 0, -3.169532e-06, 1.162546e-05, 0.0006882294, 0.0008480473, 
    0.001587595, 0.001346159, 0.001701098, 0.0009349753, 0.0009158014, 
    0.0003673836, 0.0002199015, -4.331777e-06, 0, 0.0003121342, 0.001312666, 
    0.002309358, 0.002358711, 0.001902765, 0.001318104, 0.0008496931, 
    0.0001874508, 0.0001778232,
  9.262481e-06, -5.150888e-06, 0.0001252263, -1.375048e-07, -9.66586e-08, 
    -1.243396e-05, 9.507313e-05, -1.716827e-06, 1.178867e-05, 6.521585e-05, 
    3.378963e-05, 0.0007761291, 0.0002819993, 0.0001327509, -2.090797e-06, 
    0.0002573837, -6.566916e-06, 0, 0, 0, -8.384764e-06, 7.138918e-06, 
    0.0001703355, 3.964709e-06, 9.838216e-05, -8.058289e-06, 9.348241e-09, 
    -1.83941e-11, 5.012776e-06,
  0, 0, 0, -1.46977e-06, 0, 0, 0, 0, 0, 0, -2.068584e-06, 1.221568e-09, 0, 
    3.993203e-10, 0, 0, 0, 0, 0, 0, -1.496259e-07, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.910303e-11, 5.154954e-09, 
    1.7268e-08, -1.735501e-11, 0, 0, 0, 0, 0, 0, -6.662993e-12, 
    -4.784483e-11, 2.146498e-10, -5.640593e-11, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.336138e-11, 0, 0, 0, 
    0, 0, 0, -5.598166e-07, 0, 0, 0, 0,
  0, 0, -4.194577e-08, -4.505735e-07, 0, 3.765821e-06, -6.561997e-06, 
    1.713604e-05, 5.443056e-07, 6.160628e-06, -3.130133e-11, -2.226209e-08, 
    -5.124627e-06, 0.0003185146, 0.0001317245, 3.181229e-07, 0.0002508239, 
    -9.937221e-06, 0.0001511773, 1.939759e-05, 2.338804e-07, 0, -9.05828e-07, 
    6.059174e-05, 0, 0, -8.538655e-07, 7.461706e-05, 5.249638e-05,
  0.0004810396, 2.90778e-05, 2.444376e-06, 0.0002855638, 0.002519726, 
    0.001078235, 0.0008106229, 0.000899985, 0.0005220821, 2.399237e-06, 
    1.830278e-05, 0.0001421016, 0.001577139, 0.001771621, 0.0004655088, 
    0.001534925, 0.0005134364, 0.0004922317, 0.0004744242, 0.001175188, 
    0.0008862155, 0.0005187679, 0.0006175198, 9.862866e-05, 2.171203e-05, 
    0.001357652, 0.001976992, 0.001021127, 0.0008211384,
  0.0002830519, 3.999905e-05, 0.0003851561, 0.004745455, 0.006841906, 
    0.005967798, 0.002482861, 0.001643151, -2.250897e-07, 0.0006386507, 
    0.001728354, 0.003383891, 0.002349034, 0.004693422, 0.002150556, 
    0.002825881, 0.00565252, 0.005380918, 0.009050894, 0.005401212, 
    0.005320231, 0.003172781, 0.0009079747, 0.000302623, 0.006414688, 
    0.01259744, 0.009140843, 0.002961506, 0.001222521,
  -1.712479e-06, -4.968612e-06, 0.0009866687, 0.007390792, 0.01109124, 
    0.008669855, 0.008701344, 0.0001022416, 0.001192365, 0.001255022, 
    0.001384575, 0.00190443, 0.002638076, 0.006612192, 0.009553171, 
    0.01446732, 0.01312786, 0.01213203, 0.01546036, 0.004554791, 0.002491549, 
    -1.595509e-05, 0, 2.11172e-08, 0.005197042, 0.0170961, 0.01291987, 
    0.001177622, 0.0004550829,
  1.611188e-07, 0.002718335, 0.003892577, 0.007048812, 0.02034036, 
    0.01016618, 0.007713697, 0.004564157, 0.003265836, 0.005792395, 
    0.007458895, 0.008341402, 0.01139554, 0.008994672, 0.01458385, 
    0.01978967, 0.01581546, 0.009218534, 0.002745861, 0.0005175711, 
    0.0004015267, -1.805105e-07, 1.941109e-05, 0.0009484013, 0.01566131, 
    0.0093979, 0.005127899, 1.502774e-05, -8.561476e-07,
  -7.996103e-08, 0.005711363, 0.01271695, 0.007184647, 0.0176191, 0.02120428, 
    0.02586236, 0.02545404, 0.01775448, 0.005541295, 0.01287401, 0.01464051, 
    0.02663683, 0.04221684, 0.03713237, 0.02492351, 0.0124206, 0.004014446, 
    0.002193769, -3.454068e-07, -4.963899e-06, 0.000160428, -3.852005e-07, 
    0.02122482, 0.02702814, 0.008258192, 0.001766102, 8.540233e-06, 
    1.179298e-07,
  0.003220916, 0.01560937, 0.009839154, 0.0004041374, 0.00746042, 0.02142066, 
    0.01670036, 0.01105798, 0.01803919, 0.03301645, 0.0137326, 0.01458057, 
    0.03946031, 0.0356239, 0.02074502, 0.003058471, 0.002455615, 0.002315826, 
    0.0007448627, 0.0003383829, 0.0006655358, 0.001304303, 0.002574033, 
    0.02867183, 0.01061462, 0.01186602, 0.007831465, 0.001439896, 0.002461855,
  0.004210462, 0.002415967, 0.002322918, 0.002089876, 0.0009075204, 
    0.001172885, 0.005597401, 0.01560898, 0.01371022, 0.02586111, 0.02922418, 
    0.04459711, 0.06920499, 0.05101082, 0.02362701, 0.02597041, 0.02583492, 
    0.02772891, 0.02167743, 0.02486393, 0.05155712, 0.04275416, 0.0274843, 
    0.007778961, 0.004529664, 0.00746284, 0.007655129, 0.02082288, 0.009258986,
  -5.502971e-08, -1.069105e-07, 2.586875e-05, 0.001538589, 0.002012898, 
    0.01147754, 0.03110808, 0.03045611, 0.01923501, 0.02402855, 0.04277398, 
    0.03705501, 0.02635598, 0.01610051, 0.0008662364, 0.000655996, 
    0.001636506, 0.006403603, 0.004359624, 0.002262613, 0.006806847, 
    0.01162572, 0.004838623, 0.005288533, 0.003124569, 0.003049142, 
    0.001123682, 0.0001843816, 6.677862e-05,
  0, -8.968398e-06, 0.0003427592, 0.0005334612, 0.0009300514, 0.0002705785, 
    0.01764163, 0.003998469, 0.01285215, 0.02130333, 0.02178951, 0.01610921, 
    0.0199168, 0.008861132, 0.005740428, 0.003580711, 0.00150715, 0.00408193, 
    0.001437183, 0.0005021475, 0.0008789908, 0.003669041, 0.008300247, 
    0.006169883, 0.003878488, 0.003716531, 0.00106537, -2.598071e-06, 
    -5.428863e-06,
  0.0002056409, 0.0005235658, 0.0002420349, 7.048732e-05, 0.0005929436, 
    0.0003445979, 0.0003094085, 3.455102e-05, 0.001805994, 0.003310767, 
    0.0104806, 0.0162927, 0.01671723, 0.0185645, 0.01123529, 0.005813825, 
    0.003207758, 0.001908659, 0.0004545175, 6.762482e-05, 5.148334e-05, 
    0.003772408, 0.008900097, 0.006128426, 0.008826664, 0.008851464, 
    0.002340508, 0.0006583053, 0.0002199576,
  0.0002463952, 0.0003114458, 0.0004253326, 0.0002228339, 0.0002117439, 
    5.052751e-05, -1.253885e-06, 4.500562e-05, 0.0007921829, 0.002374857, 
    0.002892792, 0.004815456, 0.005427947, 0.005650831, 0.002253159, 
    0.001572339, 0.002174319, 0.001471925, 0.000540139, -5.412221e-06, 
    0.001150717, 0.002791423, 0.004746463, 0.004808043, 0.006131148, 
    0.00447034, 0.004077903, 0.001476994, 0.0006497749,
  0.0002276017, 0.0004430191, 0.0004142973, -3.488125e-06, 0.0005041274, 
    9.07366e-05, 0.0001986054, 0.0001093198, 0.0001864626, 0.0006959864, 
    0.0003441922, 0.002974623, 0.001505428, 0.0008378188, 0.0004379985, 
    0.0007439813, 0.0003760235, -2.605765e-07, 4.058261e-05, -1.07494e-06, 
    0.000227322, 0.0001690217, 0.0006165692, 0.0005769192, 0.0008897783, 
    0.0005702345, 0.0002305832, -1.120376e-05, 0.0001245816,
  0, -1.434625e-09, -1.784611e-08, -5.504507e-06, -3.302611e-06, 
    -3.717086e-06, 8.979304e-05, 0.0001518177, 0.000110725, 3.01505e-05, 
    -2.054915e-06, -4.60993e-06, -4.860215e-06, -4.6615e-06, -9.823689e-07, 
    0, 0, 0, 0, -3.609449e-06, 3.167688e-05, -7.202232e-07, -8.893576e-07, 
    -1.112473e-10, 8.079535e-05, -3.167056e-07, 0, 0, -1.874589e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.599162e-12, -6.899097e-11, 
    9.91641e-09, 1.066449e-08, 0, 0, 1.022264e-10, -5.997156e-12, 0, 0, 
    2.146159e-11, 2.08709e-09, -2.977834e-10, 1.196863e-09, -1.70156e-12, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.67427e-06, 0, 0, 0, 
    -1.322752e-06, 0, 0, 7.095442e-05, 0, -3.100918e-07, -4.794864e-06, 0, 0, 
    0, 0,
  9.874618e-05, -1.041716e-06, -6.973242e-07, 4.526132e-06, 7.82014e-05, 
    0.0002839167, 0.0002221856, 0.0002101681, 0.0002214424, 0.0001718235, 
    2.134511e-06, 3.325097e-05, 3.711723e-05, 0.0007320507, 0.0009529897, 
    1.928533e-05, 0.0006390027, 0.0005219335, 0.0004481793, 0.0001162993, 
    0.0001252173, 2.960603e-06, 1.547991e-05, 0.0002455923, 4.094406e-07, 
    -5.962141e-07, 0.0001190124, 0.000111654, 0.0001169605,
  0.002171885, 0.001541471, 0.000340108, 0.001507969, 0.006565722, 
    0.004380269, 0.003055806, 0.002892683, 0.001539624, 0.0006415854, 
    0.0001498095, 0.0006253769, 0.002874739, 0.004921651, 0.002065663, 
    0.003017615, 0.001637719, 0.001971314, 0.001855266, 0.003263064, 
    0.003194753, 0.002678621, 0.002436103, 0.0007528234, 0.0003003387, 
    0.003883419, 0.005486508, 0.004159363, 0.003432257,
  0.002573659, 0.001134328, 0.0008586479, 0.0104687, 0.01533753, 0.01321368, 
    0.006483898, 0.003709086, 0.0003023122, 0.001436323, 0.004175204, 
    0.00731858, 0.005055268, 0.01037099, 0.007000614, 0.01116656, 0.01100531, 
    0.01317787, 0.02079283, 0.01949919, 0.01328591, 0.007486518, 0.002988044, 
    0.001298232, 0.01116313, 0.02291088, 0.02114483, 0.00929335, 0.005452447,
  9.381653e-05, 0.0003143811, 0.003731901, 0.01737562, 0.02044194, 
    0.01901425, 0.01656067, 0.001091673, 0.004903501, 0.003839662, 
    0.005645206, 0.006002584, 0.004851977, 0.01362552, 0.02351727, 
    0.03342176, 0.03069561, 0.03165267, 0.03847897, 0.012213, 0.007602446, 
    0.0008155772, 0.0003634771, 0.0006162578, 0.0126751, 0.03281082, 
    0.02702694, 0.003003128, 0.001206503,
  5.005053e-05, 0.01106616, 0.01578759, 0.02364481, 0.04328537, 0.02901541, 
    0.01764212, 0.008229728, 0.009340366, 0.01499098, 0.03417956, 0.03059406, 
    0.03499246, 0.03070381, 0.05062833, 0.0553577, 0.04455576, 0.02792151, 
    0.007380448, 0.001938292, 0.0009637089, 7.946522e-05, 0.0001517803, 
    0.01917823, 0.07708925, 0.0175353, 0.01015385, 0.0001022057, 1.935265e-05,
  4.633685e-05, 0.02849422, 0.03508749, 0.01920459, 0.04075919, 0.05337564, 
    0.05636874, 0.06884212, 0.06108934, 0.04521764, 0.03813611, 0.08804182, 
    0.1018046, 0.1554452, 0.1358926, 0.08430523, 0.03902297, 0.01207714, 
    0.005009852, 0.0002855962, 0.0001342567, 0.000801962, 0.002378488, 
    0.08795626, 0.1215075, 0.02725829, 0.005626099, 0.0002834921, 0.0001072105,
  0.01947033, 0.03597961, 0.03711713, 0.001333602, 0.01499909, 0.03877638, 
    0.04442638, 0.05499807, 0.07549809, 0.09112228, 0.08833785, 0.1107986, 
    0.1582847, 0.1278766, 0.08704292, 0.02658859, 0.0109721, 0.008149676, 
    0.002734094, 0.003491065, 0.003069517, 0.005864337, 0.01118811, 
    0.1114859, 0.0637693, 0.02723846, 0.01734859, 0.007937508, 0.0119643,
  0.02200934, 0.009457314, 0.007888312, 0.004025691, 0.003029399, 0.01615446, 
    0.06742686, 0.1909274, 0.1635218, 0.1546581, 0.1619445, 0.1763268, 
    0.2172071, 0.1518842, 0.1132241, 0.08672122, 0.05799107, 0.0520794, 
    0.04208402, 0.05304778, 0.1033185, 0.1133257, 0.06689318, 0.04232989, 
    0.01667816, 0.01704695, 0.0153908, 0.04140248, 0.02481277,
  0.0003479463, 1.870974e-05, 0.001178096, 0.008894043, 0.02287371, 
    0.04287836, 0.09098148, 0.08198497, 0.1078412, 0.07707785, 0.1053708, 
    0.09741886, 0.1004945, 0.04237259, 0.00973435, 0.003772531, 0.006480494, 
    0.01710343, 0.01567343, 0.01021737, 0.03736431, 0.04792911, 0.02155974, 
    0.02168017, 0.006021362, 0.005678236, 0.002903818, 0.001307063, 
    0.0003248022,
  7.429087e-05, 0.0002043104, 0.0008085587, 0.00139468, 0.002546717, 
    0.001999782, 0.01950751, 0.007409996, 0.02222431, 0.0574096, 0.06360663, 
    0.06276793, 0.06824704, 0.03710617, 0.02039718, 0.00997424, 0.0066027, 
    0.01057525, 0.004776005, 0.001989923, 0.003445315, 0.02289646, 
    0.03956071, 0.01800729, 0.009782541, 0.009430634, 0.002831729, 
    0.0001036135, 0.0001117715,
  0.00100977, 0.002162627, 0.0006878283, 0.0004205293, 0.001440973, 
    0.001011382, 0.0007365444, 0.001506422, 0.009727016, 0.010918, 
    0.03174091, 0.04674301, 0.05073709, 0.0440827, 0.0287916, 0.01955401, 
    0.01044189, 0.007871796, 0.002007907, 0.000435016, 0.000160255, 
    0.007119123, 0.01726467, 0.01857777, 0.02156751, 0.01857367, 0.008462051, 
    0.002342462, 0.0004529054,
  0.001362497, 0.001587666, 0.002688025, 0.001269277, 0.0004678736, 
    0.0005201807, 3.703713e-05, 0.0005953939, 0.002676095, 0.005634265, 
    0.00771643, 0.01155893, 0.01445184, 0.01377977, 0.00878601, 0.004308808, 
    0.006976799, 0.005381433, 0.002205329, 8.79821e-05, 0.002665834, 
    0.005668201, 0.008369147, 0.008421877, 0.01170162, 0.01250585, 
    0.01342419, 0.006268308, 0.002867309,
  0.001165243, 0.0009721118, 0.001470635, 0.000189742, 0.001506956, 
    0.0008485719, 0.0005732565, 0.0008217851, 0.0005131707, 0.002187943, 
    0.001746728, 0.00511011, 0.00324442, 0.002166714, 0.00132687, 0.0014251, 
    0.00107052, 0.0002961482, 0.0002023691, 0.0004992905, 0.0007916164, 
    0.0005193193, 0.002328051, 0.001241896, 0.003580747, 0.002755147, 
    0.001607735, 0.0003336544, 0.001890263,
  0, -1.293418e-06, 1.793378e-05, 8.74875e-05, 2.148802e-05, 0.0001094029, 
    0.0003538756, 0.0004460246, 0.0002746666, 0.0002541183, 0.0001627619, 
    7.897963e-06, 2.089876e-05, 3.377886e-05, 9.162027e-05, -7.056379e-08, 
    -2.060807e-07, -9.8882e-07, -6.857553e-07, 3.481746e-06, 0.0006463618, 
    2.721361e-05, 1.966043e-05, -1.992636e-06, 0.0002763441, -1.376278e-06, 
    -1.319471e-07, 9.791792e-05, 0.000114523,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 6.036712e-06, -8.673499e-08, -4.438897e-11, 
    1.855446e-09, 1.5128e-05, -1.470608e-05, -7.959151e-10, 0, 0, 0, 0, 0, 0, 
    0, -8.065917e-11, -4.241045e-09, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.202541e-06, -1.91132e-06, 1.408826e-05, 0, 0, 0, 0,
  -9.99515e-06, 0, 0, -1.511612e-07, 0, 0, -4.426236e-07, -1.846349e-06, 
    -1.636011e-12, 0, 0, 0, -5.458616e-06, -4.662136e-06, 0.0001676659, 
    1.37364e-09, -2.236668e-11, 0.0001136595, 1.333516e-06, 8.986511e-06, 0, 
    0.0002316921, -4.682393e-07, 4.319131e-06, 2.296209e-06, 0, 0, 
    7.680275e-05, 0.00015911,
  0.0003994303, 7.522265e-05, 2.600429e-05, 0.0001380672, 0.0005692818, 
    0.001301001, 0.001662902, 0.001407609, 0.0009135971, 0.0002936068, 
    6.551377e-05, 0.0002482726, 0.0004116664, 0.001247591, 0.002816202, 
    0.0007970939, 0.001878885, 0.001583408, 0.001282873, 0.0004881998, 
    0.0006134156, 7.688961e-05, 0.001026258, 0.0007075936, 0.0004453096, 
    0.0001069754, 0.0004602202, 0.0004136978, 0.000233025,
  0.007277032, 0.005049112, 0.001882734, 0.004195153, 0.01462315, 0.01227634, 
    0.008207466, 0.00802369, 0.004192907, 0.002330296, 0.0008338802, 
    0.00188737, 0.005786501, 0.01033418, 0.007071896, 0.00592237, 
    0.005927646, 0.005715122, 0.007576076, 0.007924535, 0.00847088, 
    0.007335726, 0.007758634, 0.003496695, 0.001719207, 0.00821069, 
    0.01177254, 0.01116833, 0.008504128,
  0.01107568, 0.004684628, 0.003210562, 0.02122341, 0.03313477, 0.03503617, 
    0.02048142, 0.0105499, 0.003207968, 0.004747761, 0.01026675, 0.0149771, 
    0.01214056, 0.02092703, 0.01873362, 0.02642061, 0.02685634, 0.03206063, 
    0.04505742, 0.04557805, 0.03500894, 0.0186589, 0.00650826, 0.004160082, 
    0.01880551, 0.03821113, 0.04571827, 0.03181493, 0.01856285,
  0.002416648, 0.002043482, 0.02132724, 0.04737281, 0.0523108, 0.05619872, 
    0.04967938, 0.02023927, 0.02399443, 0.01886705, 0.02219822, 0.02385312, 
    0.01331479, 0.03458906, 0.05657909, 0.0782887, 0.08358478, 0.09839262, 
    0.1203528, 0.04599742, 0.01868901, 0.01101482, 0.002750669, 0.005729794, 
    0.03790033, 0.08971908, 0.08792423, 0.02925521, 0.01048324,
  0.001491253, 0.04035131, 0.08147129, 0.03804974, 0.065446, 0.05656357, 
    0.04003971, 0.01991281, 0.01898325, 0.02445106, 0.0501519, 0.04123725, 
    0.04040774, 0.04680081, 0.08190723, 0.1050487, 0.1162537, 0.1273133, 
    0.08613334, 0.02946983, 0.007357708, 0.004551654, 0.005779858, 
    0.03899139, 0.1073338, 0.09356166, 0.06499231, 0.02602668, 0.006258065,
  0.001831316, 0.06570164, 0.1930535, 0.08467282, 0.07718398, 0.09121349, 
    0.09932335, 0.1039856, 0.07251969, 0.04740888, 0.04669333, 0.08230665, 
    0.09391349, 0.1457562, 0.1358758, 0.09993177, 0.06500324, 0.02719643, 
    0.02018542, 0.007498342, 0.004642254, 0.004224181, 0.01397737, 0.2430185, 
    0.2156655, 0.1333802, 0.0617912, 0.02656485, 0.001981039,
  0.04825455, 0.2228079, 0.2748346, 0.02643049, 0.04514833, 0.1040851, 
    0.1375007, 0.1649089, 0.2837998, 0.3047686, 0.122373, 0.1264329, 
    0.1562653, 0.117028, 0.07473179, 0.02127087, 0.01172112, 0.01174353, 
    0.005934307, 0.01318282, 0.01832367, 0.02315364, 0.0535582, 0.2980507, 
    0.1835147, 0.07712278, 0.07090621, 0.0396429, 0.02564996,
  0.1172637, 0.1016625, 0.08436049, 0.007734298, 0.01869701, 0.03735558, 
    0.1014375, 0.1776847, 0.1448657, 0.1376026, 0.1383051, 0.1507728, 
    0.1879579, 0.1345106, 0.1166749, 0.1215881, 0.09441966, 0.09615029, 
    0.08601528, 0.1115977, 0.1738651, 0.1484708, 0.1673666, 0.1115678, 
    0.05685109, 0.06832036, 0.0746353, 0.1244688, 0.1404249,
  0.02021248, 0.005175686, 0.004233647, 0.0152915, 0.02839908, 0.04674017, 
    0.09672508, 0.07141458, 0.1134575, 0.06462329, 0.09698393, 0.08418573, 
    0.0944878, 0.06688179, 0.05588425, 0.04772523, 0.04261997, 0.06278237, 
    0.07133801, 0.0548569, 0.1016198, 0.08437407, 0.05759993, 0.08272077, 
    0.07004485, 0.03648344, 0.02058816, 0.04482024, 0.02351472,
  0.002115989, 0.002567287, 0.001845831, 0.003080324, 0.004877937, 
    0.003615227, 0.01609696, 0.01394806, 0.04093023, 0.07903636, 0.08668647, 
    0.08915565, 0.09844608, 0.07902803, 0.07431704, 0.04648222, 0.04256241, 
    0.03608693, 0.01318651, 0.009895437, 0.02122765, 0.06407113, 0.09052949, 
    0.08794115, 0.07672488, 0.04880229, 0.01385568, 0.005624107, 0.0009239387,
  0.004671707, 0.00628533, 0.001803998, 0.001325209, 0.003767043, 
    0.002843125, 0.002342479, 0.009498038, 0.02377156, 0.0292867, 0.05928404, 
    0.08022718, 0.09579722, 0.1038698, 0.08198807, 0.07578281, 0.04476317, 
    0.0345087, 0.01421544, 0.001898473, 0.0007870522, 0.02471743, 0.04713021, 
    0.05611348, 0.07550945, 0.05488493, 0.03202182, 0.01133547, 0.003640873,
  0.004697137, 0.004456494, 0.005630808, 0.00280806, 0.00250178, 0.003416396, 
    0.0009609551, 0.001133402, 0.00487647, 0.01139133, 0.02157487, 
    0.03412902, 0.03613912, 0.04356409, 0.03139998, 0.02595679, 0.02477721, 
    0.02294108, 0.01194444, 0.001234622, 0.005005225, 0.01069881, 0.01572284, 
    0.01754745, 0.02486124, 0.03308789, 0.03610301, 0.01946168, 0.01130277,
  0.00349763, 0.001976816, 0.002958252, 0.001236268, 0.002553698, 
    0.002040226, 0.002176189, 0.00381247, 0.00175259, 0.004826873, 
    0.006059204, 0.009679306, 0.01004714, 0.009786025, 0.008684059, 
    0.00629895, 0.0024393, 0.00260984, 0.0008705633, 0.001346662, 
    0.002455869, 0.002035004, 0.004811159, 0.002644462, 0.009197724, 
    0.01068421, 0.007936982, 0.004232693, 0.004262301,
  -8.270718e-06, 0.0002784441, 0.0003425182, 0.0004574405, 0.0003964649, 
    0.0005661705, 0.0007475929, 0.001021614, 0.0006321018, 0.0009278799, 
    0.0004895974, 0.0001687218, 0.0003386085, 0.001201299, 0.001210946, 
    0.0001891683, 0.0001713627, 3.063745e-05, 1.741797e-06, 0.0001125955, 
    0.001728584, 0.0004718991, 0.0004819891, 0.0002235919, 0.0007119805, 
    0.0001122677, 2.424012e-05, 0.0007507784, 0.000539429,
  0, -2.609875e-08, 1.407751e-10, -1.42834e-05, -9.797009e-07, 0, 0, 
    -5.746724e-06, -2.531843e-05, 0.0002022608, -5.787267e-06, -1.689191e-06, 
    5.513838e-05, 5.132195e-05, 0.000160743, -6.03107e-07, -1.395636e-07, 
    -1.034398e-06, 2.806698e-06, -1.570257e-07, 0.0001912734, -3.266836e-06, 
    0, -9.412636e-07, -2.878816e-09, 0, 0, -5.777748e-15, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.95239e-07, -4.351936e-08, 
    -5.377989e-09, 2.487017e-05, 2.20178e-05, 1.141306e-06, -2.920485e-08, 0, 
    0, 9.694416e-06, 1.33825e-05, 1.408826e-05, -1.881389e-06, 0, 0, 0,
  0.0003692244, 4.566551e-05, -2.184962e-06, 1.168566e-06, -1.055401e-10, 
    -9.792692e-07, 0.0002696184, -1.121669e-05, -1.276712e-06, 0, 0, 0, 
    5.893693e-05, 3.088068e-05, 0.0006499857, 0.0004069229, 0.0003071325, 
    0.0002432628, 0.0007773575, 0.001214587, 0.0001808549, 0.0006266406, 
    0.0003915864, 3.458528e-05, 0.0002059462, 0, 1.781855e-05, 0.0002554194, 
    0.0002386259,
  0.001666738, 0.001175628, 0.0002769322, 0.0007489499, 0.001775894, 
    0.002897596, 0.003754803, 0.002400877, 0.002725363, 0.001375799, 
    0.0004490542, 0.001258299, 0.00142898, 0.003417509, 0.008812311, 
    0.007438728, 0.007244855, 0.005887468, 0.004153842, 0.002198999, 
    0.002625843, 0.001776888, 0.002838578, 0.003270231, 0.0020379, 
    0.0009397765, 0.001789392, 0.002036431, 0.001291071,
  0.02433475, 0.01864372, 0.01155353, 0.01568222, 0.03381698, 0.0323492, 
    0.02707541, 0.02273511, 0.01791157, 0.01232191, 0.008407873, 0.009492137, 
    0.01352291, 0.02406676, 0.0242861, 0.02287469, 0.02601784, 0.02050026, 
    0.01880813, 0.02378883, 0.02800208, 0.0273323, 0.02533991, 0.0116249, 
    0.007960722, 0.01947213, 0.02481347, 0.03146345, 0.02929291,
  0.04485215, 0.02594024, 0.02377409, 0.05000681, 0.06481788, 0.07063948, 
    0.05138727, 0.03629659, 0.0271544, 0.02682288, 0.03624288, 0.04152576, 
    0.0319965, 0.04433242, 0.04160905, 0.05772436, 0.05708244, 0.06656607, 
    0.08469099, 0.1112589, 0.09564451, 0.06204423, 0.02922077, 0.01385088, 
    0.04035044, 0.07402673, 0.08643565, 0.0817318, 0.05917022,
  0.02047556, 0.01473877, 0.0384201, 0.06038909, 0.07012708, 0.07765389, 
    0.07128882, 0.03884568, 0.04055645, 0.03995313, 0.05597003, 0.04761897, 
    0.03332963, 0.05900764, 0.08160079, 0.1125171, 0.1238987, 0.1468144, 
    0.2076098, 0.1431828, 0.09228463, 0.04112998, 0.0172772, 0.01924099, 
    0.0519106, 0.107971, 0.12754, 0.07308263, 0.03862603,
  0.0004332738, 0.03178573, 0.08438483, 0.0344899, 0.05979825, 0.04654346, 
    0.03351329, 0.01783676, 0.01915302, 0.02166808, 0.04685127, 0.03409575, 
    0.03424412, 0.04309122, 0.07822173, 0.09857418, 0.1058314, 0.1158016, 
    0.07795107, 0.03262907, 0.01867682, 0.003386798, 0.002081467, 0.0311668, 
    0.08604682, 0.1043078, 0.05807911, 0.02861191, 0.006400016,
  0.0004726518, 0.04855732, 0.1705846, 0.06808664, 0.0592178, 0.06494121, 
    0.07579817, 0.08198703, 0.05916443, 0.03713738, 0.03693642, 0.0638426, 
    0.07420312, 0.1170829, 0.1088458, 0.0768922, 0.04716449, 0.01978419, 
    0.01432049, 0.00451198, 0.002686261, 0.00205015, 0.007297414, 0.2083103, 
    0.1794457, 0.1135076, 0.0487572, 0.01580437, 0.0008533255,
  0.0299829, 0.1829631, 0.1926618, 0.01898378, 0.0295416, 0.074138, 
    0.09464185, 0.1173981, 0.2223934, 0.2508735, 0.08511136, 0.09693044, 
    0.1219002, 0.09352998, 0.0579289, 0.01458731, 0.008818333, 0.008895601, 
    0.004358488, 0.0040229, 0.005578616, 0.0117281, 0.03539708, 0.2336187, 
    0.138068, 0.06080421, 0.05095434, 0.02351246, 0.01404276,
  0.09517543, 0.08286964, 0.06679387, 0.04349329, 0.01367991, 0.02357276, 
    0.06358032, 0.1267055, 0.1156264, 0.09556171, 0.1031613, 0.1191786, 
    0.1588706, 0.1138603, 0.08868434, 0.09585015, 0.07736306, 0.07731052, 
    0.06238826, 0.08158788, 0.138935, 0.1197235, 0.1365972, 0.08083385, 
    0.03879836, 0.04847619, 0.05565311, 0.1047215, 0.1309564,
  0.07701819, 0.0160534, 0.006130317, 0.01518545, 0.0356866, 0.04355858, 
    0.09333567, 0.06007696, 0.1015472, 0.05520406, 0.08844019, 0.07340968, 
    0.07990996, 0.05139988, 0.04415262, 0.03849267, 0.04201475, 0.06293097, 
    0.07788016, 0.05797177, 0.08463476, 0.07148091, 0.04406901, 0.06601358, 
    0.05591927, 0.04197708, 0.03639806, 0.06586504, 0.08435201,
  0.02648148, 0.02219989, 0.01446294, 0.01067291, 0.01326297, 0.01347851, 
    0.02896748, 0.03378744, 0.06686612, 0.08558387, 0.09770244, 0.1010633, 
    0.1055967, 0.0854515, 0.09165371, 0.08543476, 0.08743005, 0.06825907, 
    0.05416355, 0.034402, 0.038507, 0.1013339, 0.1224209, 0.115724, 
    0.1210076, 0.1025716, 0.05490193, 0.02035466, 0.01691164,
  0.02847991, 0.02098884, 0.00724111, 0.004565698, 0.01349475, 0.01399508, 
    0.004936929, 0.02670557, 0.04696266, 0.04444202, 0.07502344, 0.08875312, 
    0.1160506, 0.1303083, 0.1155019, 0.1341336, 0.1047696, 0.09958182, 
    0.04450221, 0.00848657, 0.01123389, 0.04126855, 0.0637646, 0.08415995, 
    0.1163835, 0.1100828, 0.08502473, 0.04359371, 0.02340522,
  0.03151259, 0.0143785, 0.01667119, 0.009713665, 0.01410505, 0.01639582, 
    0.009427223, 0.003192818, 0.008891374, 0.02949985, 0.04064308, 
    0.05018249, 0.05044736, 0.06050307, 0.05806695, 0.05331986, 0.05950896, 
    0.07124462, 0.05443512, 0.006886368, 0.01808262, 0.03420457, 0.03208486, 
    0.03650557, 0.05145429, 0.07312673, 0.08338362, 0.06656535, 0.0499772,
  0.02031559, 0.006491961, 0.01054663, 0.005860924, 0.008338723, 0.01185761, 
    0.01170077, 0.01019214, 0.008007612, 0.01613648, 0.02458015, 0.02508235, 
    0.01842067, 0.02218003, 0.02187842, 0.018207, 0.01258751, 0.01578332, 
    0.003657555, 0.006424379, 0.008127208, 0.01216878, 0.01297527, 
    0.00938149, 0.01985458, 0.021979, 0.02127724, 0.01907634, 0.01950226,
  0.001626761, 0.002161591, 0.002748398, 0.004199574, 0.00230727, 0.00164604, 
    0.002884996, 0.003921815, 0.004240874, 0.005530067, 0.005337401, 
    0.004415329, 0.004845524, 0.007714522, 0.003794924, 0.002778041, 
    0.002378698, 0.003728706, 0.004171525, 0.00401214, 0.005766835, 
    0.002077827, 0.001818178, 0.001116014, 0.001955999, 0.0003020223, 
    0.0002058363, 0.00373001, 0.003724775,
  1.54337e-05, -4.129195e-06, 5.434338e-05, 6.07982e-05, -1.283916e-05, 
    0.0001029414, 2.874413e-05, 0.0002355669, 1.022264e-05, 0.0002644448, 
    0.0001106805, -7.337316e-06, 7.728166e-05, 0.0003772147, 0.0005766149, 
    0.0001667602, 0.0001293405, 5.678922e-05, 0.0001648499, -1.982624e-06, 
    0.0003130818, 0.0001376218, 3.195804e-05, -1.203323e-06, -1.041254e-05, 
    7.535477e-07, -1.319975e-11, -2.146227e-06, 5.140118e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.085346e-05, -1.160376e-05, 
    -2.205898e-05, 0.0001059588, 7.42676e-05, 2.42625e-06, -6.420087e-07, 0, 
    0, 5.618183e-05, 2.460812e-05, 1.644592e-05, -9.673499e-06, 
    -1.281071e-06, 0, 0,
  0.001024881, 0.0009230383, 0.0005832639, 0.0001601274, -5.06711e-07, 
    4.212452e-05, 0.0005871829, 8.148809e-05, -1.877833e-05, -2.780183e-06, 
    -9.7855e-07, -3.936027e-06, 0.0003069739, 0.0009714838, 0.002554771, 
    0.002522123, 0.003199304, 0.003020574, 0.003435065, 0.004815018, 
    0.003329393, 0.002689295, 0.001192126, 0.001133041, 0.001301149, 
    1.357921e-05, 3.557392e-05, 0.0004051768, 0.0004421523,
  0.005682683, 0.007524446, 0.005836536, 0.00316293, 0.008043365, 0.01019764, 
    0.01373011, 0.01204703, 0.01167235, 0.008913966, 0.006365373, 
    0.005447316, 0.008379017, 0.01431007, 0.0234032, 0.02335135, 0.02330616, 
    0.01916942, 0.01745064, 0.01242078, 0.01142904, 0.007325706, 0.00930136, 
    0.01098097, 0.01158348, 0.009848769, 0.009310478, 0.009364658, 0.006570823,
  0.06399422, 0.05800762, 0.05015082, 0.0623435, 0.08587021, 0.08356272, 
    0.06821688, 0.06965478, 0.06094683, 0.04829907, 0.04298663, 0.04734347, 
    0.0500214, 0.06252771, 0.05532036, 0.05420412, 0.05676328, 0.05536835, 
    0.05819977, 0.05869441, 0.07353915, 0.0747727, 0.08249433, 0.03627519, 
    0.04169317, 0.06399359, 0.06556934, 0.06881261, 0.06946304,
  0.0804058, 0.06249766, 0.05630348, 0.08713246, 0.1028068, 0.09839583, 
    0.08022383, 0.07686118, 0.05881695, 0.05424664, 0.06841566, 0.07067815, 
    0.05515795, 0.07381596, 0.07189945, 0.09457821, 0.09961577, 0.09717739, 
    0.1191991, 0.1478183, 0.1437393, 0.1211815, 0.07838069, 0.04000093, 
    0.08959624, 0.1133367, 0.1244346, 0.1231983, 0.1051918,
  0.02344118, 0.01351019, 0.05987515, 0.05876252, 0.07052914, 0.07642234, 
    0.06985519, 0.03883649, 0.03976133, 0.04094235, 0.06187875, 0.05067891, 
    0.04208466, 0.06251071, 0.08738786, 0.1123839, 0.1300273, 0.1501362, 
    0.2097398, 0.1453975, 0.08823464, 0.04452797, 0.01896495, 0.02100064, 
    0.04842303, 0.1032189, 0.124041, 0.07208668, 0.0405826,
  0.0002537064, 0.02572007, 0.07370892, 0.03112742, 0.05475878, 0.04191867, 
    0.03022988, 0.01599568, 0.01943136, 0.01832772, 0.04547419, 0.02976559, 
    0.02947108, 0.04512966, 0.0764764, 0.09091774, 0.09695747, 0.09840243, 
    0.05804291, 0.02163427, 0.01334126, 0.00155968, 0.0007141102, 0.0256727, 
    0.07129539, 0.09581129, 0.0462261, 0.01871006, 0.002988747,
  0.0001587111, 0.04142156, 0.1466929, 0.06284907, 0.05192656, 0.05348399, 
    0.06619858, 0.07374629, 0.05607161, 0.03402257, 0.03423956, 0.05478648, 
    0.06593801, 0.102336, 0.09869469, 0.0695496, 0.04302296, 0.01742266, 
    0.01024393, 0.001913605, 0.00146315, 0.000592032, 0.003317342, 0.1854377, 
    0.1630616, 0.1012259, 0.03443988, 0.01046227, 0.000154332,
  0.01935447, 0.1585778, 0.141994, 0.01055319, 0.02283063, 0.06266055, 
    0.0770533, 0.08963058, 0.1825255, 0.2171441, 0.06777162, 0.07986864, 
    0.1117346, 0.08729199, 0.05340068, 0.01272489, 0.007460531, 0.007875249, 
    0.003167005, 0.001834039, 0.00319393, 0.00595653, 0.02856778, 0.1902722, 
    0.1136959, 0.0582537, 0.04299949, 0.01702138, 0.008268598,
  0.08428802, 0.07770345, 0.05961073, 0.03361244, 0.01231389, 0.01585853, 
    0.04878287, 0.08277984, 0.100273, 0.07663074, 0.08379015, 0.1044589, 
    0.1409651, 0.104709, 0.07632955, 0.08324596, 0.07172067, 0.07167009, 
    0.05371372, 0.07153488, 0.1219472, 0.1065797, 0.1165361, 0.06916519, 
    0.03228462, 0.04074199, 0.04715509, 0.09040877, 0.1193608,
  0.06752352, 0.0169368, 0.004546297, 0.01436466, 0.03297007, 0.04095327, 
    0.09155429, 0.0510793, 0.09331453, 0.04806592, 0.07795516, 0.06690152, 
    0.07010362, 0.04570012, 0.03743248, 0.02948211, 0.0364191, 0.05173418, 
    0.06993027, 0.04726768, 0.06742299, 0.05835862, 0.0383206, 0.05639422, 
    0.04438723, 0.03715242, 0.03522821, 0.05919814, 0.08557115,
  0.04677945, 0.03850898, 0.02627843, 0.02773179, 0.02425467, 0.02761971, 
    0.04486831, 0.04498483, 0.08422284, 0.09813941, 0.1048986, 0.1009024, 
    0.1087755, 0.08940092, 0.09735842, 0.09491356, 0.08906636, 0.08746695, 
    0.07711703, 0.04680161, 0.06309699, 0.1009772, 0.1198893, 0.112131, 
    0.113543, 0.1012237, 0.07418908, 0.03684707, 0.03864209,
  0.06784932, 0.04977625, 0.02849561, 0.01640287, 0.03507218, 0.03583716, 
    0.009504217, 0.0551526, 0.07464409, 0.06554679, 0.08840799, 0.1019869, 
    0.1278782, 0.1476915, 0.1393299, 0.1707178, 0.1529051, 0.1633729, 
    0.08493046, 0.03090634, 0.02579288, 0.05691087, 0.09301947, 0.1221216, 
    0.1495276, 0.1522727, 0.1306105, 0.08324843, 0.05734665,
  0.07194155, 0.05210445, 0.05153643, 0.04857057, 0.04279115, 0.04936435, 
    0.02817465, 0.0109231, 0.02694136, 0.04623988, 0.0485408, 0.06274755, 
    0.0600878, 0.06894117, 0.07489643, 0.08002251, 0.09465811, 0.1241894, 
    0.1127419, 0.02538445, 0.03892933, 0.05352207, 0.04708692, 0.0557757, 
    0.0795596, 0.1102003, 0.12532, 0.110371, 0.09527206,
  0.06064236, 0.03719851, 0.03067903, 0.02638504, 0.02680386, 0.03097995, 
    0.03544275, 0.02904596, 0.02576252, 0.03109868, 0.03797079, 0.04180938, 
    0.03290979, 0.0456665, 0.03574036, 0.03677126, 0.02902718, 0.04907716, 
    0.02276668, 0.03288762, 0.03729142, 0.04452625, 0.03286671, 0.027201, 
    0.04720669, 0.04684215, 0.05353324, 0.05034031, 0.05872914,
  0.01869392, 0.02057477, 0.01489, 0.01730957, 0.01363561, 0.01185314, 
    0.01317686, 0.01642222, 0.01714092, 0.02580242, 0.02163327, 0.01734822, 
    0.02615844, 0.02668661, 0.02613236, 0.01983156, 0.018502, 0.01527745, 
    0.01528195, 0.02385492, 0.02253568, 0.01640018, 0.00941144, 0.004192234, 
    0.0152475, 0.0005642799, 0.000664487, 0.0256351, 0.02174008,
  0.002894879, 0.003931042, 0.006606709, 0.004867501, 0.002578166, 
    0.004193543, 0.002317076, 0.003107313, 0.002674604, 0.004476844, 
    0.005344527, 0.006098742, 0.004322062, 0.005341751, 0.003693787, 
    0.005232378, 0.005431039, 0.005905773, 0.006087409, 0.005526002, 
    0.006698978, 0.006849091, 0.00307048, -6.132152e-05, 0.0001133637, 
    1.691433e-05, -0.0001090261, 0.0004518092, 0.004043923,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.783305e-09, 0.0007897037, 
    -3.555289e-05, 0.0005060769, 0.0008737987, 0.0008372249, 0.0006889898, 
    0.0002084224, -1.979878e-05, -3.539687e-06, 0.0001772446, 0.0003894677, 
    0.0005278328, -6.40527e-05, 9.899814e-05, -3.331779e-06, 0,
  0.003845043, 0.00365426, 0.0029545, 0.00106951, -2.345483e-05, 
    9.217153e-05, 0.004250078, 0.0004110568, 2.740853e-05, -8.586352e-05, 
    -4.53093e-06, 1.22058e-05, 0.001034033, 0.006929608, 0.01102785, 
    0.01117242, 0.01084414, 0.01054543, 0.01410823, 0.01222321, 0.01072279, 
    0.006425907, 0.005204251, 0.005468658, 0.008245979, 0.003652572, 
    0.002244204, 0.002335588, 0.004264127,
  0.03206569, 0.0290234, 0.02126731, 0.02529497, 0.02637607, 0.02982277, 
    0.03508913, 0.03314792, 0.03401258, 0.0308757, 0.02790773, 0.02986348, 
    0.04144548, 0.05310782, 0.06123052, 0.06179715, 0.06131479, 0.0537774, 
    0.05152534, 0.04242904, 0.04018873, 0.03788886, 0.0409627, 0.04346975, 
    0.04331305, 0.04369788, 0.03464179, 0.03389728, 0.0292265,
  0.1159739, 0.1094439, 0.1145912, 0.1274133, 0.1386565, 0.1347894, 
    0.1125563, 0.1179671, 0.1103578, 0.1014834, 0.09955997, 0.1060343, 
    0.1037754, 0.1055681, 0.09916887, 0.09817653, 0.1067215, 0.106447, 
    0.1024058, 0.104298, 0.1188222, 0.1225656, 0.1341351, 0.07342757, 
    0.08826392, 0.1220654, 0.1139651, 0.1169877, 0.1189572,
  0.1132694, 0.08292192, 0.0727322, 0.1044377, 0.1088648, 0.1034943, 
    0.09325997, 0.0898921, 0.07413352, 0.07243279, 0.08437014, 0.08610611, 
    0.0731618, 0.09414428, 0.09173454, 0.1072659, 0.1158911, 0.1174384, 
    0.1340349, 0.1601117, 0.1534854, 0.1353415, 0.1007795, 0.06794202, 
    0.1142709, 0.1266491, 0.1418943, 0.1389255, 0.130536,
  0.0200459, 0.009610539, 0.0551013, 0.05181681, 0.06477658, 0.06891081, 
    0.06357308, 0.03162219, 0.03664241, 0.03627938, 0.0632366, 0.04993176, 
    0.04282621, 0.05827296, 0.08244885, 0.1041048, 0.1199109, 0.1388725, 
    0.1931855, 0.1315847, 0.07305446, 0.03591427, 0.01692447, 0.01382741, 
    0.04293678, 0.09449679, 0.1136161, 0.06060028, 0.03672604,
  0.0001028113, 0.02146481, 0.0630441, 0.02592563, 0.04921823, 0.03791893, 
    0.02759473, 0.01693626, 0.02015666, 0.01546255, 0.04134369, 0.02457294, 
    0.02863752, 0.04723139, 0.0789929, 0.08494274, 0.08648767, 0.08462, 
    0.04672706, 0.01637927, 0.007379017, 0.00271492, 0.001777711, 0.02174721, 
    0.0572226, 0.09237738, 0.04016974, 0.01285984, 0.002902562,
  0.0001524575, 0.03763396, 0.125719, 0.05366813, 0.04617978, 0.04406004, 
    0.05957528, 0.06622569, 0.05045529, 0.03018958, 0.03228131, 0.04885041, 
    0.06232794, 0.08846577, 0.08794846, 0.06091612, 0.0380117, 0.01422531, 
    0.008080124, 0.000965468, 0.0005514619, 1.970741e-05, 0.001853304, 
    0.1477075, 0.142565, 0.08445619, 0.02463584, 0.005497958, 1.223026e-05,
  0.01426552, 0.1310907, 0.1010859, 0.008132638, 0.01963871, 0.05272583, 
    0.06323041, 0.06504742, 0.1358677, 0.1760619, 0.05219873, 0.06637477, 
    0.09740707, 0.07694346, 0.04915988, 0.01233297, 0.007290273, 0.00609158, 
    0.002920929, 0.001549444, 0.003621517, 0.003030664, 0.02304544, 0.147884, 
    0.08982792, 0.06383204, 0.03745253, 0.01190949, 0.006545592,
  0.07032982, 0.06818301, 0.04853229, 0.028262, 0.01133238, 0.01076209, 
    0.03913402, 0.0537113, 0.08711622, 0.06328676, 0.07231065, 0.08919667, 
    0.1228287, 0.09609459, 0.06515729, 0.07222682, 0.06869093, 0.06833509, 
    0.04924912, 0.06563892, 0.1084431, 0.0919165, 0.09075605, 0.05100337, 
    0.02755001, 0.03753598, 0.04231552, 0.07999092, 0.1003955,
  0.05388316, 0.01179837, 0.003538673, 0.01369004, 0.02835022, 0.03698675, 
    0.08649425, 0.04284132, 0.0874913, 0.04345287, 0.07218835, 0.06005373, 
    0.05790954, 0.04001693, 0.02928929, 0.02379199, 0.0283516, 0.03908318, 
    0.0548306, 0.03958157, 0.05744787, 0.04918119, 0.03052706, 0.04762124, 
    0.03297579, 0.03251713, 0.02919117, 0.05192367, 0.07402851,
  0.04839177, 0.04151285, 0.02822778, 0.03106022, 0.02715214, 0.03131477, 
    0.0432508, 0.04457232, 0.09950729, 0.104754, 0.1016804, 0.1001535, 
    0.10463, 0.08892418, 0.09360963, 0.08802154, 0.07807141, 0.07827597, 
    0.06349058, 0.03505376, 0.06545576, 0.08444472, 0.09751065, 0.09722269, 
    0.09515283, 0.0846249, 0.05994697, 0.03364991, 0.04577834,
  0.09826127, 0.07114244, 0.05014849, 0.03651, 0.05343983, 0.05285057, 
    0.02174267, 0.08169737, 0.09024806, 0.07790658, 0.09813541, 0.1147508, 
    0.140112, 0.1615089, 0.1540416, 0.1801596, 0.1714433, 0.1784409, 
    0.09950113, 0.06295961, 0.04137084, 0.07733262, 0.1186161, 0.136149, 
    0.1566593, 0.1650355, 0.1408292, 0.09322902, 0.08548802,
  0.1221044, 0.09566373, 0.07704511, 0.07191416, 0.08179183, 0.07214083, 
    0.0450516, 0.02503337, 0.04514835, 0.05832161, 0.05872234, 0.07212869, 
    0.07585921, 0.08177917, 0.0963835, 0.1078835, 0.1321194, 0.1616231, 
    0.1539809, 0.05384946, 0.06202113, 0.07492115, 0.06758236, 0.08060177, 
    0.1063567, 0.1411441, 0.1594511, 0.1442201, 0.1368784,
  0.1068093, 0.06675798, 0.06552374, 0.05698881, 0.05349901, 0.05314577, 
    0.07116309, 0.05779817, 0.04394101, 0.0447837, 0.05118465, 0.05464667, 
    0.04556185, 0.0644266, 0.05121208, 0.07385902, 0.0578256, 0.09945545, 
    0.06861461, 0.06206263, 0.05783333, 0.06567746, 0.05217484, 0.05236964, 
    0.08819535, 0.09534824, 0.09428633, 0.1010958, 0.1115928,
  0.05508713, 0.05815896, 0.04783062, 0.04709297, 0.05060549, 0.04821404, 
    0.04236557, 0.04424868, 0.03953901, 0.03795815, 0.03559072, 0.03378572, 
    0.04182287, 0.03906534, 0.04545928, 0.0431235, 0.04623627, 0.05486349, 
    0.05946703, 0.07041781, 0.05407522, 0.03851315, 0.03065296, 0.01589698, 
    0.05093844, 0.003197182, 0.001755713, 0.06686226, 0.06001326,
  0.02251051, 0.02823885, 0.03132833, 0.02667128, 0.02555766, 0.02205708, 
    0.0211793, 0.02421475, 0.02282652, 0.02407446, 0.02909544, 0.02728393, 
    0.02417711, 0.02027544, 0.0195222, 0.02407165, 0.03140434, 0.03308626, 
    0.03394981, 0.03006138, 0.02271285, 0.02601788, 0.0155653, 0.007963674, 
    0.008591882, 0.001027801, 3.407403e-05, 0.008566044, 0.02164566,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.130374e-05, 0.001360853, 0.001488549, 
    0.002961621, 0.00333017, 0.002770245, 0.00205845, 0.0007741603, 
    5.805073e-06, -3.850354e-06, 0.001041016, 0.008543018, 0.006860781, 
    0.004295836, 0.004994595, 8.434042e-06, 0,
  0.01264228, 0.01209611, 0.009934346, 0.005924158, -6.147451e-05, 
    0.001231622, 0.01748039, 0.001003169, 0.0008036708, 0.0005034084, 
    0.0003281112, 0.0002905978, 0.001922798, 0.03063903, 0.03793217, 
    0.03561648, 0.03694525, 0.03676856, 0.03464692, 0.03454299, 0.03643796, 
    0.03635988, 0.02818665, 0.02206831, 0.03317, 0.02445317, 0.01999857, 
    0.01707556, 0.01381622,
  0.07254883, 0.07018412, 0.0672833, 0.07760751, 0.07560056, 0.06877053, 
    0.07994672, 0.07404038, 0.07424013, 0.06958773, 0.07291089, 0.08591372, 
    0.111467, 0.124856, 0.1184273, 0.1210011, 0.1139044, 0.1074077, 
    0.1058837, 0.09720968, 0.09240495, 0.09136806, 0.101619, 0.1104955, 
    0.110062, 0.09697545, 0.09154245, 0.08278616, 0.07594331,
  0.1504757, 0.1543972, 0.1654149, 0.1772495, 0.1776876, 0.1697677, 
    0.1431214, 0.1503217, 0.1459571, 0.1447004, 0.147957, 0.150151, 
    0.1469972, 0.1403752, 0.1407901, 0.1374235, 0.1323225, 0.1338347, 
    0.1336342, 0.1340188, 0.1517577, 0.1496169, 0.1681845, 0.1157038, 
    0.1215491, 0.1685486, 0.1569808, 0.1500929, 0.1504147,
  0.1140026, 0.08079366, 0.0713552, 0.1008866, 0.09873784, 0.09541102, 
    0.09225135, 0.08830757, 0.07324789, 0.07350679, 0.08361737, 0.09459346, 
    0.08239589, 0.1077101, 0.1013229, 0.1182876, 0.1202328, 0.1189203, 
    0.1299685, 0.1581201, 0.1470618, 0.1353642, 0.1049119, 0.08482107, 
    0.105318, 0.1162429, 0.1347485, 0.1362978, 0.1287331,
  0.01604326, 0.006018375, 0.04809014, 0.04507704, 0.05923091, 0.06181396, 
    0.05750511, 0.02698325, 0.03088102, 0.03101954, 0.05856769, 0.04686856, 
    0.04070746, 0.05373422, 0.07695205, 0.09635922, 0.1102312, 0.1283588, 
    0.1810809, 0.1183612, 0.06512208, 0.02677174, 0.0110883, 0.009722464, 
    0.03910311, 0.08682685, 0.09989747, 0.05165996, 0.03182334,
  0.0001627347, 0.01892741, 0.05293613, 0.02192748, 0.04550097, 0.03281715, 
    0.02553947, 0.01648824, 0.01740481, 0.01371622, 0.03393594, 0.02030339, 
    0.02779195, 0.04835396, 0.0746907, 0.08212896, 0.07546928, 0.07192925, 
    0.03786223, 0.012341, 0.003893705, 0.001722923, 0.001745795, 0.01828626, 
    0.04564057, 0.08569959, 0.0351232, 0.009349083, 0.002111254,
  0.0003086571, 0.0331663, 0.1044589, 0.04609192, 0.03970859, 0.03656529, 
    0.05317449, 0.0586024, 0.04326409, 0.0249046, 0.03216509, 0.04103827, 
    0.05798836, 0.07236405, 0.0739779, 0.05545958, 0.03155001, 0.01159896, 
    0.006004632, 0.0006988775, 0.0004750644, -3.77166e-05, 0.0009484703, 
    0.1097762, 0.1229822, 0.06774937, 0.01960073, 0.001656876, 1.157133e-05,
  0.01226903, 0.1126364, 0.07765614, 0.007469947, 0.01821485, 0.04400982, 
    0.05018778, 0.04628256, 0.09563877, 0.1457885, 0.04117171, 0.05028951, 
    0.08057895, 0.06127756, 0.0408241, 0.01109486, 0.006886959, 0.005099565, 
    0.001805301, 0.001878813, 0.002502995, 0.001801575, 0.02137142, 
    0.1135423, 0.07114089, 0.06957714, 0.03484562, 0.009189364, 0.006276069,
  0.05563959, 0.0557139, 0.04326067, 0.02971106, 0.01127096, 0.008029997, 
    0.03037908, 0.03629364, 0.06955543, 0.05247325, 0.05927354, 0.07427102, 
    0.104254, 0.08691623, 0.05741522, 0.06021309, 0.06747171, 0.06333726, 
    0.05209075, 0.06610635, 0.09522755, 0.07883997, 0.07274829, 0.03624167, 
    0.02449984, 0.03520612, 0.03831522, 0.07417405, 0.08668226,
  0.04081728, 0.007370356, 0.002859663, 0.01269278, 0.02895017, 0.03628889, 
    0.08019793, 0.03626655, 0.07877728, 0.03983865, 0.06916175, 0.05386507, 
    0.04625583, 0.03549386, 0.02035568, 0.01877112, 0.02171315, 0.03121645, 
    0.04319377, 0.03132046, 0.04967507, 0.04386326, 0.02245089, 0.03890936, 
    0.02674662, 0.02893811, 0.02454038, 0.04265685, 0.05728811,
  0.04150658, 0.037096, 0.02534313, 0.02611852, 0.02701287, 0.0288644, 
    0.03771858, 0.04554266, 0.1126185, 0.1027236, 0.09836503, 0.09631661, 
    0.101883, 0.08269387, 0.08564729, 0.0806028, 0.06839907, 0.06361946, 
    0.0481335, 0.02606453, 0.05528153, 0.06776395, 0.07844622, 0.07936435, 
    0.07730015, 0.07103624, 0.04721321, 0.02693484, 0.03935005,
  0.1015985, 0.08061555, 0.06553771, 0.05968152, 0.07091956, 0.0707956, 
    0.04082399, 0.1067114, 0.09785885, 0.08107461, 0.106881, 0.1248262, 
    0.1445315, 0.1667295, 0.170297, 0.1791738, 0.1711841, 0.1685684, 
    0.09512664, 0.08390911, 0.05848364, 0.08924779, 0.1226419, 0.1305734, 
    0.1514843, 0.157558, 0.1316703, 0.08376659, 0.08184563,
  0.1446937, 0.1329219, 0.1171464, 0.1113059, 0.1151035, 0.1058037, 
    0.06792799, 0.04225073, 0.05749383, 0.07318068, 0.07466294, 0.08107515, 
    0.09359712, 0.09867511, 0.1220672, 0.1330623, 0.1516937, 0.1766825, 
    0.1763697, 0.0905695, 0.08595403, 0.09615441, 0.101506, 0.1051044, 
    0.1280531, 0.1528313, 0.1716124, 0.1536016, 0.148264,
  0.1609838, 0.1160331, 0.09940968, 0.1029755, 0.09948882, 0.08906879, 
    0.1058777, 0.09025734, 0.06503846, 0.06303134, 0.06307957, 0.06385086, 
    0.05575602, 0.07800873, 0.08061302, 0.1110993, 0.1068745, 0.1423921, 
    0.1173733, 0.08518399, 0.08248472, 0.08526466, 0.07632405, 0.07824774, 
    0.1221377, 0.1258098, 0.1274762, 0.1473709, 0.1555221,
  0.1030561, 0.09639909, 0.07961246, 0.0690533, 0.08053152, 0.08082438, 
    0.06224874, 0.06063516, 0.05173582, 0.04907376, 0.04868523, 0.04186591, 
    0.05095923, 0.05672659, 0.0740312, 0.07746379, 0.09021145, 0.09013104, 
    0.08456734, 0.09743366, 0.0747109, 0.06290098, 0.06466229, 0.0439681, 
    0.07953911, 0.01670301, 0.004246802, 0.1128108, 0.1040418,
  0.05016585, 0.05510022, 0.0532664, 0.04546226, 0.04899993, 0.05566373, 
    0.0591029, 0.05510172, 0.05058114, 0.04744136, 0.05110396, 0.04714867, 
    0.04336938, 0.03914402, 0.04187404, 0.05249808, 0.06069253, 0.06292354, 
    0.06740603, 0.0605924, 0.04954633, 0.05210305, 0.03498022, 0.01869363, 
    0.03026826, 0.008640277, 0.009212804, 0.02015544, 0.04831699,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.10124e-06, 0.0002142576, 0.0002695889, 
    0.00298499, 0.007547922, 0.01729297, 0.025589, 0.01830797, 0.007613771, 
    0.003170957, 0.001093157, 0.0001727745, 0.006198118, 0.03382958, 
    0.02680432, 0.01382439, 0.01581103, 0.002953606, 1.589121e-05,
  0.04777897, 0.05342361, 0.0554363, 0.03857526, 0.0002919543, 0.005382907, 
    0.03750373, 0.00353313, 0.002770533, 0.002899107, 0.002014182, 
    0.0008914306, 0.01136679, 0.07906379, 0.08373148, 0.07721862, 0.07748714, 
    0.08136157, 0.07750794, 0.08351453, 0.07943518, 0.09199964, 0.09607504, 
    0.08298788, 0.1000287, 0.07779513, 0.07385497, 0.06129234, 0.05716662,
  0.1312008, 0.1247397, 0.1288968, 0.1415512, 0.1350322, 0.1248622, 
    0.1295036, 0.1282621, 0.1290134, 0.1256514, 0.1357161, 0.1651368, 
    0.1882338, 0.1921108, 0.1803273, 0.1790681, 0.1771759, 0.1670138, 
    0.1575301, 0.1543047, 0.1512978, 0.1493324, 0.1636185, 0.1701514, 
    0.1781419, 0.1625403, 0.1442566, 0.1399246, 0.1350504,
  0.1686348, 0.1732418, 0.1827494, 0.1946421, 0.1846138, 0.1747151, 
    0.1534473, 0.1627406, 0.165082, 0.1655752, 0.1764765, 0.1728882, 
    0.1723237, 0.1681292, 0.1543718, 0.140922, 0.144716, 0.1473505, 
    0.1493016, 0.1551176, 0.1756884, 0.1723365, 0.1884134, 0.1463984, 
    0.1370895, 0.1794545, 0.1740825, 0.1640563, 0.1690671,
  0.1077208, 0.07399372, 0.06434996, 0.09381443, 0.08804082, 0.08775819, 
    0.08933765, 0.08261815, 0.06820226, 0.06866938, 0.07837438, 0.09425837, 
    0.08362687, 0.1079151, 0.1070849, 0.1168662, 0.1134963, 0.1160812, 
    0.1220251, 0.15124, 0.1447261, 0.1317569, 0.1077859, 0.08824951, 
    0.09117822, 0.1056678, 0.1246447, 0.1285906, 0.1227785,
  0.01284411, 0.00417411, 0.04336659, 0.04338095, 0.05315789, 0.05964058, 
    0.04688046, 0.02349264, 0.02538912, 0.02440758, 0.05215445, 0.04728071, 
    0.03875691, 0.04960756, 0.07005786, 0.08926191, 0.1026413, 0.1213585, 
    0.1686322, 0.1036316, 0.05546621, 0.0186795, 0.007485419, 0.008336983, 
    0.03693961, 0.07935023, 0.08625892, 0.04670923, 0.02831187,
  0.0002087502, 0.01726259, 0.04364121, 0.01826822, 0.04365951, 0.02995371, 
    0.02336679, 0.01557454, 0.01336185, 0.01228992, 0.02615218, 0.01764438, 
    0.02740967, 0.04649864, 0.06900335, 0.07852392, 0.06781309, 0.06064987, 
    0.03076173, 0.01100365, 0.001642691, 0.0002561049, 0.001034988, 
    0.01635969, 0.03901718, 0.0793668, 0.03118139, 0.006572453, 0.0006780794,
  0.0005434601, 0.03283106, 0.08599556, 0.03888062, 0.03988295, 0.03347282, 
    0.05021879, 0.05558568, 0.0386262, 0.02152198, 0.03061514, 0.03790278, 
    0.06079756, 0.06565227, 0.06755425, 0.05044, 0.02824443, 0.01046715, 
    0.005116533, 0.0007427197, 0.0001813826, -7.827803e-06, 0.001109133, 
    0.08573146, 0.1090323, 0.05538727, 0.01551907, 0.0003672384, 1.194362e-05,
  0.01568487, 0.09714787, 0.06340793, 0.008555353, 0.01722176, 0.04121437, 
    0.04418674, 0.03792149, 0.06962456, 0.1320235, 0.03628167, 0.04145487, 
    0.07013221, 0.05317871, 0.03513563, 0.01069168, 0.00820626, 0.004990671, 
    0.002430488, 0.002426196, 0.002716571, 0.002340152, 0.02405749, 
    0.09162547, 0.06389222, 0.07508783, 0.03527652, 0.009931466, 0.006822817,
  0.04497157, 0.04570425, 0.03915859, 0.03063787, 0.009220295, 0.007375041, 
    0.02513937, 0.03026574, 0.05790309, 0.04706562, 0.05451686, 0.0659536, 
    0.09176329, 0.0815532, 0.05421773, 0.05630039, 0.06611349, 0.06196031, 
    0.05618123, 0.07024888, 0.09325718, 0.07028699, 0.06135202, 0.02787994, 
    0.02473455, 0.03537238, 0.03324758, 0.06471666, 0.07556907,
  0.0280869, 0.004414679, 0.003036772, 0.01358684, 0.02611846, 0.03372994, 
    0.07180837, 0.03154857, 0.06902076, 0.03898522, 0.06843976, 0.05141845, 
    0.03964508, 0.03228614, 0.01438233, 0.01626923, 0.01739259, 0.02665024, 
    0.0305186, 0.0279131, 0.04197923, 0.04204677, 0.01625891, 0.03374352, 
    0.02112854, 0.0211441, 0.01810342, 0.03318658, 0.04349185,
  0.03248408, 0.03285909, 0.02389424, 0.0240311, 0.02524456, 0.02660625, 
    0.03495914, 0.05236311, 0.1298868, 0.1040944, 0.0938261, 0.0897564, 
    0.09704244, 0.07927456, 0.07647388, 0.07127956, 0.05725286, 0.05188035, 
    0.03680455, 0.01922686, 0.04522553, 0.05458169, 0.06448067, 0.06444732, 
    0.0639269, 0.0567821, 0.03819001, 0.0214185, 0.03575228,
  0.09394285, 0.07956311, 0.06844366, 0.07648648, 0.08221085, 0.08261599, 
    0.06611869, 0.1169586, 0.1019372, 0.08210331, 0.1128433, 0.1281274, 
    0.1496885, 0.1690453, 0.1691788, 0.1758487, 0.1728531, 0.1598745, 
    0.08726945, 0.08714966, 0.08153185, 0.09217227, 0.1145024, 0.1244106, 
    0.145068, 0.1475029, 0.1206688, 0.0756868, 0.07402363,
  0.1492203, 0.148341, 0.1354476, 0.1361833, 0.1455341, 0.1415377, 0.1039545, 
    0.055099, 0.07436849, 0.0897723, 0.09485345, 0.09309123, 0.1161314, 
    0.1182353, 0.1433526, 0.1515934, 0.1689247, 0.1860783, 0.1774025, 
    0.1141186, 0.09680244, 0.1126929, 0.1268166, 0.1326233, 0.1431004, 
    0.1549115, 0.1732062, 0.1544245, 0.1518982,
  0.1811894, 0.1505519, 0.1301388, 0.1395339, 0.1375007, 0.1344408, 
    0.1524481, 0.1358865, 0.1023511, 0.08375365, 0.06786083, 0.06795385, 
    0.06949252, 0.1091493, 0.1177461, 0.1510386, 0.1407661, 0.1830432, 
    0.155809, 0.1172169, 0.1028664, 0.1156211, 0.09844651, 0.1072891, 
    0.151999, 0.1562071, 0.1485381, 0.1794741, 0.1783442,
  0.141846, 0.1300508, 0.1116725, 0.1118396, 0.1183375, 0.1096829, 
    0.09481618, 0.08794507, 0.06400594, 0.06752084, 0.06232492, 0.07022727, 
    0.0724442, 0.08863185, 0.1094889, 0.1143658, 0.1263553, 0.121364, 
    0.1134658, 0.1196246, 0.09878427, 0.07656387, 0.07906505, 0.06891106, 
    0.1062921, 0.05002949, 0.01710146, 0.1462096, 0.1423703,
  0.07421429, 0.0813783, 0.07748724, 0.07453278, 0.07561658, 0.07768248, 
    0.08079261, 0.08007865, 0.06841971, 0.06804315, 0.07092825, 0.07244614, 
    0.07666489, 0.08001921, 0.08927751, 0.09898004, 0.09458675, 0.0893385, 
    0.09186446, 0.08388146, 0.07043108, 0.07445568, 0.05781107, 0.03252554, 
    0.04973772, 0.0225189, 0.02287961, 0.03268643, 0.07654507,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -1.890131e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003680586, 0.0004497501, 
    0.0006023283, 0.009180469, 0.02443177, 0.04452658, 0.06406297, 
    0.05489253, 0.02996953, 0.00797982, 0.005966169, 0.002080285, 0.02136994, 
    0.07438561, 0.06698094, 0.04009981, 0.05078088, 0.0112157, 0.0005254779,
  0.1094019, 0.1247852, 0.1203456, 0.09480736, 0.003212357, 0.0145887, 
    0.06667379, 0.00950564, 0.008635211, 0.006593939, 0.005390494, 
    0.003816091, 0.04335658, 0.1569039, 0.1599714, 0.1469335, 0.1441511, 
    0.147634, 0.1362671, 0.1441026, 0.1479108, 0.1604076, 0.1834498, 
    0.1623656, 0.1963781, 0.1456034, 0.1386932, 0.1223182, 0.1177729,
  0.1731981, 0.1704497, 0.187071, 0.1964016, 0.1844789, 0.1722884, 0.1685314, 
    0.1695175, 0.1750385, 0.1806366, 0.1902376, 0.2237885, 0.2413615, 
    0.2319876, 0.2142758, 0.2034138, 0.1995812, 0.1957582, 0.1918316, 
    0.197898, 0.2049059, 0.2088761, 0.2192264, 0.2180397, 0.2331106, 
    0.2042052, 0.1880867, 0.176236, 0.1883234,
  0.1724589, 0.1792302, 0.1820475, 0.1917435, 0.1801502, 0.1744155, 
    0.1547651, 0.1662374, 0.1719269, 0.1771304, 0.1884554, 0.1797339, 
    0.1725242, 0.1624086, 0.1490227, 0.1341496, 0.1446336, 0.1472502, 
    0.1483442, 0.1613677, 0.181572, 0.1756323, 0.1955603, 0.1587285, 
    0.1380212, 0.1768101, 0.1741184, 0.1686072, 0.1746701,
  0.1009381, 0.06833658, 0.0574616, 0.08892679, 0.08254281, 0.08113279, 
    0.08881386, 0.08050038, 0.06678502, 0.05837915, 0.07200904, 0.08661908, 
    0.07794072, 0.09975245, 0.1016673, 0.1141323, 0.106951, 0.1094264, 
    0.1170185, 0.1398198, 0.1366176, 0.1295995, 0.1059978, 0.08901071, 
    0.08166766, 0.09647573, 0.1154326, 0.1198875, 0.1138267,
  0.01117266, 0.005117807, 0.04035083, 0.04195195, 0.05025576, 0.05637662, 
    0.03916574, 0.01795464, 0.02062799, 0.02077981, 0.05042288, 0.04776723, 
    0.03737815, 0.04953681, 0.06593407, 0.08253333, 0.09606415, 0.1170637, 
    0.159064, 0.08663538, 0.0520627, 0.01532252, 0.005538125, 0.007513975, 
    0.03587285, 0.07528292, 0.07805807, 0.04203542, 0.02731261,
  0.0002888275, 0.01516034, 0.03619125, 0.01583274, 0.04248105, 0.02711665, 
    0.02440013, 0.01574799, 0.01078766, 0.01122472, 0.02406287, 0.01502821, 
    0.02795564, 0.04591844, 0.06359194, 0.07513334, 0.06199024, 0.05527735, 
    0.02740175, 0.01024865, 0.0003779742, 5.239829e-05, 0.0001227478, 
    0.01207066, 0.03447247, 0.07516168, 0.02709841, 0.006781295, 0.0008131789,
  0.001048998, 0.03391756, 0.07453075, 0.0359171, 0.03754983, 0.03441735, 
    0.04949703, 0.05240281, 0.03489801, 0.0196947, 0.03328886, 0.03684689, 
    0.06434927, 0.06418595, 0.06675666, 0.04603324, 0.02646622, 0.0114442, 
    0.005208763, 0.0009633247, 2.246868e-05, -1.441351e-05, 0.000876456, 
    0.07077678, 0.1042181, 0.04862181, 0.01215643, 0.0001991733, 1.01897e-05,
  0.02229495, 0.09181074, 0.05856966, 0.01017985, 0.01977993, 0.04236511, 
    0.0412954, 0.03556794, 0.05554585, 0.1267566, 0.03630201, 0.03627153, 
    0.06464726, 0.04679201, 0.03383722, 0.009966171, 0.006577797, 
    0.004083244, 0.00379396, 0.002680918, 0.003717028, 0.002893446, 
    0.03021236, 0.08216213, 0.06710903, 0.08049932, 0.04029646, 0.01241359, 
    0.008139848,
  0.03939965, 0.04144998, 0.03975558, 0.03679559, 0.0107316, 0.007846661, 
    0.0238381, 0.02679862, 0.0526995, 0.0458238, 0.05269773, 0.06192917, 
    0.08421656, 0.07668862, 0.05480079, 0.05733978, 0.06572944, 0.06141418, 
    0.06435081, 0.07754377, 0.09363181, 0.06623749, 0.0543847, 0.0238144, 
    0.02516122, 0.03497745, 0.03288893, 0.05960274, 0.06844047,
  0.02503966, 0.003860285, 0.003985215, 0.0126652, 0.02491351, 0.03274382, 
    0.06916524, 0.03011126, 0.06638009, 0.03893362, 0.06807888, 0.0538906, 
    0.03638541, 0.02732776, 0.0106402, 0.01375064, 0.01626395, 0.02091201, 
    0.02521351, 0.02473835, 0.03335765, 0.04160049, 0.01266849, 0.03098148, 
    0.01647129, 0.0182905, 0.01718131, 0.0263638, 0.03379589,
  0.02907318, 0.03171885, 0.02179867, 0.02349414, 0.02459736, 0.02525588, 
    0.03525714, 0.06581233, 0.1487633, 0.1079816, 0.09336641, 0.08501934, 
    0.09671692, 0.07737447, 0.07049138, 0.06134646, 0.04836852, 0.04874589, 
    0.03143989, 0.01548389, 0.03617754, 0.04418433, 0.05851825, 0.05383583, 
    0.05537964, 0.05156467, 0.02956614, 0.01908404, 0.03269807,
  0.08269799, 0.07741256, 0.06794188, 0.0905441, 0.07920388, 0.07638876, 
    0.08495779, 0.1147026, 0.09929743, 0.09088185, 0.1127889, 0.122546, 
    0.1471684, 0.1643228, 0.165231, 0.1733116, 0.1677871, 0.1483141, 
    0.08037788, 0.08754633, 0.09301715, 0.09278778, 0.1091388, 0.1222979, 
    0.1389814, 0.1368311, 0.1094058, 0.06911398, 0.0713158,
  0.147026, 0.1534644, 0.1384515, 0.1399512, 0.1431567, 0.1445171, 0.1296545, 
    0.07530015, 0.0899231, 0.1103867, 0.1164759, 0.113102, 0.1379687, 
    0.1453625, 0.1657743, 0.1665615, 0.1746741, 0.1878956, 0.1772018, 
    0.1210041, 0.1081798, 0.1295144, 0.148424, 0.1541583, 0.1582975, 
    0.1602935, 0.1725473, 0.1540651, 0.1528642,
  0.1946135, 0.1678416, 0.1498419, 0.1733887, 0.1687387, 0.1681406, 
    0.1823823, 0.1756261, 0.1513866, 0.1209785, 0.08387843, 0.07776531, 
    0.09626044, 0.1470112, 0.1541667, 0.1771525, 0.167097, 0.2194809, 
    0.1833308, 0.1369781, 0.1281858, 0.1411228, 0.1218653, 0.1372918, 
    0.1774049, 0.1875384, 0.1717091, 0.1993843, 0.1951708,
  0.1675191, 0.1576543, 0.1500039, 0.1483036, 0.1557538, 0.1455833, 
    0.1323474, 0.12747, 0.08892874, 0.1062121, 0.08309418, 0.1005901, 
    0.1043347, 0.1198536, 0.1382693, 0.1278847, 0.1441264, 0.1456271, 
    0.1387755, 0.1477836, 0.1251794, 0.09475905, 0.1029355, 0.08798764, 
    0.1235186, 0.08395299, 0.0426653, 0.1675412, 0.1678463,
  0.1131617, 0.1158465, 0.1086858, 0.110287, 0.1095058, 0.1063069, 0.0972301, 
    0.09597021, 0.08024701, 0.08384431, 0.0910044, 0.1006048, 0.1088752, 
    0.1136434, 0.1223426, 0.1227406, 0.1106802, 0.1090112, 0.1121747, 
    0.1062143, 0.09322288, 0.09845824, 0.08128012, 0.05112708, 0.07115899, 
    0.03647462, 0.036027, 0.05477737, 0.1146747,
  0.00016626, 9.834013e-05, 3.042031e-05, -3.749953e-05, -0.0001054194, 
    -0.0001733392, -0.000241259, -1.049732e-05, -4.730774e-06, 1.035769e-06, 
    6.802311e-06, 1.256885e-05, 1.83354e-05, 2.410194e-05, 0.0001396364, 
    0.0001405711, 0.0001415058, 0.0001424405, 0.0001433752, 0.0001443099, 
    0.0001452447, -0.0003016227, -0.0002404041, -0.0001791855, -0.0001179669, 
    -5.674834e-05, 4.470241e-06, 6.568883e-05, 0.0002205958,
  0.0001816021, 0.0003363212, 0.000198141, -4.157478e-06, 0, -3.550298e-05, 
    0, 0, 0, 0.0002787744, 0.0005484839, 0.0007133326, 0.0005743934, 
    0.03778711, 0.06495676, 0.09314507, 0.1139913, 0.111309, 0.06336021, 
    0.03067113, 0.01988921, 0.01139847, 0.05435544, 0.1544539, 0.1441167, 
    0.09336518, 0.1073351, 0.04162775, 0.006023417,
  0.1565764, 0.1879865, 0.184911, 0.1459061, 0.02013875, 0.03750545, 
    0.1024688, 0.02310352, 0.01756942, 0.02032524, 0.01499949, 0.01496443, 
    0.09521011, 0.2034761, 0.2058409, 0.1903464, 0.1860413, 0.1959466, 
    0.1931447, 0.1962628, 0.2056944, 0.223242, 0.2569125, 0.2480918, 
    0.2651124, 0.1943025, 0.1918827, 0.1750914, 0.1862573,
  0.1987744, 0.203301, 0.2272068, 0.2318407, 0.2210364, 0.2053166, 0.1943433, 
    0.203049, 0.2069295, 0.2228502, 0.2370698, 0.2634301, 0.2629937, 
    0.2490585, 0.2254836, 0.2129505, 0.2033008, 0.2026126, 0.2091888, 
    0.2204483, 0.2326909, 0.2390061, 0.2445822, 0.2404788, 0.2497215, 
    0.2246585, 0.2133263, 0.1996463, 0.217798,
  0.174598, 0.1811502, 0.1836445, 0.1887856, 0.1741744, 0.1704478, 0.1544511, 
    0.1692667, 0.1770242, 0.1864388, 0.1921412, 0.1799009, 0.1703113, 
    0.1553706, 0.1440067, 0.1259992, 0.1377207, 0.1413126, 0.1441799, 
    0.1597264, 0.1752795, 0.1779779, 0.1916716, 0.1617077, 0.1311153, 
    0.1725561, 0.1715584, 0.1696166, 0.1759801,
  0.0979421, 0.06427895, 0.05204358, 0.08565449, 0.08072907, 0.07729642, 
    0.08642956, 0.07567437, 0.06215543, 0.05442676, 0.06982832, 0.08186498, 
    0.07369479, 0.09518816, 0.09816863, 0.1076649, 0.1010573, 0.1024658, 
    0.1115028, 0.1298243, 0.1314031, 0.124814, 0.1034427, 0.08681232, 
    0.07293808, 0.09392645, 0.1056125, 0.1161866, 0.1094148,
  0.009614315, 0.007487838, 0.04111693, 0.04078113, 0.04593476, 0.05335191, 
    0.03212992, 0.01507251, 0.01723348, 0.01822033, 0.0523376, 0.05010207, 
    0.03790409, 0.04905329, 0.06103254, 0.07564037, 0.09053314, 0.1103847, 
    0.1476828, 0.07767744, 0.04674342, 0.01549857, 0.004551748, 0.007966325, 
    0.03567328, 0.07215334, 0.07480558, 0.03989124, 0.02723549,
  0.0005049731, 0.01703073, 0.03315504, 0.01709175, 0.04300087, 0.02570147, 
    0.0253793, 0.01722419, 0.01098054, 0.00834797, 0.02449398, 0.01453464, 
    0.02656431, 0.04630698, 0.05984315, 0.06869809, 0.05830944, 0.05192114, 
    0.02572598, 0.0101552, 0.0001062962, 9.945819e-05, 3.310433e-06, 
    0.00831008, 0.03395158, 0.07250568, 0.0249031, 0.005060044, 0.0005922676,
  0.0005369326, 0.03951772, 0.07282276, 0.03707925, 0.03799549, 0.03616832, 
    0.05077044, 0.04907954, 0.03392044, 0.02056502, 0.03483021, 0.03588673, 
    0.06864285, 0.06189553, 0.06490939, 0.04489802, 0.02516519, 0.01226061, 
    0.004763325, 0.001257626, 0.0001351407, -2.143507e-05, 0.0009633565, 
    0.05993406, 0.1015004, 0.04657304, 0.009128076, 0.0001824221, 0.000397246,
  0.03995064, 0.09255725, 0.05876468, 0.01324932, 0.02123508, 0.04036928, 
    0.03983215, 0.03341774, 0.05100131, 0.1238398, 0.0359694, 0.03257141, 
    0.05999391, 0.04352244, 0.03187364, 0.01054856, 0.007468168, 0.003622657, 
    0.005765065, 0.004231308, 0.004497123, 0.004678434, 0.03888255, 
    0.08068652, 0.06619712, 0.08075552, 0.04016363, 0.01422973, 0.0126649,
  0.03750667, 0.03891783, 0.0409209, 0.04415753, 0.01549848, 0.008799641, 
    0.02192767, 0.02521149, 0.04765378, 0.04591744, 0.05305524, 0.0589228, 
    0.08119396, 0.07612148, 0.05269649, 0.05992043, 0.06481539, 0.06346589, 
    0.07109003, 0.08952257, 0.09414449, 0.0644919, 0.05302588, 0.02224257, 
    0.02492083, 0.03141084, 0.0324805, 0.05713907, 0.06643002,
  0.0254087, 0.004988133, 0.004187043, 0.01092349, 0.02120803, 0.02667762, 
    0.06935458, 0.03261719, 0.06796753, 0.03874435, 0.0723479, 0.05701647, 
    0.03583386, 0.02546373, 0.008760083, 0.01197786, 0.01582403, 0.01553304, 
    0.02179774, 0.02031981, 0.02607436, 0.0423398, 0.01121194, 0.02886621, 
    0.01302661, 0.01860731, 0.01502005, 0.02148251, 0.02725496,
  0.0263756, 0.02725148, 0.01885952, 0.02458384, 0.02578939, 0.02382401, 
    0.03457168, 0.07637754, 0.1684961, 0.1132433, 0.09377823, 0.082651, 
    0.0935391, 0.0738572, 0.0634109, 0.05385735, 0.04332601, 0.04394969, 
    0.02601333, 0.01395893, 0.03083291, 0.0414486, 0.05353783, 0.04771066, 
    0.04901719, 0.04521573, 0.02426172, 0.01754404, 0.02926394,
  0.07491416, 0.0723726, 0.06861661, 0.09745371, 0.07379283, 0.06650464, 
    0.1115786, 0.1005556, 0.09054828, 0.09090855, 0.1071136, 0.1145771, 
    0.1412969, 0.1623386, 0.1596666, 0.1682541, 0.1620527, 0.1382568, 
    0.07336897, 0.08713361, 0.1037671, 0.09344544, 0.1098361, 0.1209327, 
    0.1378429, 0.1291802, 0.09721234, 0.06219613, 0.06414588,
  0.1383569, 0.1525823, 0.1342952, 0.1396197, 0.1352264, 0.1396068, 
    0.1345673, 0.1025847, 0.1152134, 0.1338684, 0.1358154, 0.1326427, 
    0.1540189, 0.1663517, 0.1725309, 0.1771929, 0.1824837, 0.1872029, 
    0.1716441, 0.1301975, 0.1147341, 0.1370966, 0.1603049, 0.1708069, 
    0.1687962, 0.1651056, 0.1687706, 0.1560497, 0.1505716,
  0.205456, 0.1827623, 0.1632513, 0.1962775, 0.1903162, 0.1877031, 0.2066461, 
    0.2001084, 0.1892854, 0.157729, 0.1105313, 0.1019634, 0.1202227, 
    0.1746465, 0.1787846, 0.1930611, 0.1918966, 0.2514314, 0.213204, 
    0.1524221, 0.1445527, 0.1657237, 0.1466563, 0.171624, 0.1994586, 
    0.2207349, 0.1831074, 0.2144285, 0.2076888,
  0.1905963, 0.1867836, 0.1921541, 0.1838089, 0.1913048, 0.1808549, 
    0.1751549, 0.1754692, 0.1268697, 0.137981, 0.105442, 0.1437241, 0.136825, 
    0.154332, 0.1622697, 0.1420257, 0.1607931, 0.1698439, 0.1679941, 
    0.1721367, 0.1488404, 0.1139768, 0.134295, 0.1114388, 0.1431147, 
    0.1130723, 0.0655527, 0.1915184, 0.1882752,
  0.1435439, 0.1498126, 0.1399979, 0.1429149, 0.1279811, 0.1247551, 
    0.1212945, 0.1191922, 0.1065743, 0.109108, 0.1155169, 0.1246139, 
    0.1357762, 0.1478385, 0.1569061, 0.1579735, 0.1430849, 0.1352934, 
    0.1321942, 0.1247433, 0.1096441, 0.1174275, 0.1004391, 0.06263558, 
    0.08879069, 0.05310698, 0.05662367, 0.07493658, 0.1496041,
  0.003762479, 0.003652136, 0.003541793, 0.00343145, 0.003321107, 
    0.003210763, 0.003100421, 0.003494198, 0.003384356, 0.003274515, 
    0.003164674, 0.003054833, 0.002944991, 0.00283515, 0.001976876, 
    0.002206491, 0.002436107, 0.002665723, 0.002895338, 0.003124954, 
    0.00335457, 0.004145918, 0.004136486, 0.004127054, 0.004117623, 
    0.004108191, 0.00409876, 0.004089329, 0.003850753,
  0.008397367, 0.0007188815, 0.0005710291, 0.0001830681, 7.88352e-05, 
    0.0001310354, -5.044847e-05, -1.625474e-05, 2.298983e-05, 0.0007650605, 
    0.0006566088, 0.0008869024, 0.002014976, 0.08867482, 0.09791227, 
    0.1270544, 0.1593074, 0.1617246, 0.1087244, 0.06693347, 0.04545304, 
    0.0339783, 0.09790436, 0.2038656, 0.1922429, 0.1661575, 0.1756233, 
    0.08383818, 0.02444876,
  0.1949392, 0.2341766, 0.2237546, 0.2049746, 0.06718218, 0.06930462, 
    0.1375781, 0.04859918, 0.03912144, 0.05152923, 0.0404537, 0.03881094, 
    0.1481372, 0.2363906, 0.23958, 0.2221357, 0.2095992, 0.2331271, 
    0.2351173, 0.2367435, 0.2432826, 0.259846, 0.2894079, 0.3034626, 
    0.2960139, 0.2119812, 0.2123691, 0.1992234, 0.2230949,
  0.2105558, 0.2248619, 0.2492595, 0.2481283, 0.2442327, 0.2282843, 
    0.2172502, 0.2247117, 0.2360661, 0.2534941, 0.2647129, 0.2786716, 
    0.2661345, 0.2536279, 0.2290968, 0.2126964, 0.2072636, 0.2051406, 
    0.2127785, 0.2313235, 0.2418262, 0.2521298, 0.2588285, 0.2470456, 
    0.2499034, 0.229791, 0.2126923, 0.2078625, 0.2230331,
  0.1767825, 0.1806248, 0.1806195, 0.182745, 0.168868, 0.1678001, 0.1575716, 
    0.1734643, 0.18273, 0.1948383, 0.193939, 0.1776647, 0.1645137, 0.154771, 
    0.1444117, 0.1137372, 0.1298543, 0.1353831, 0.140185, 0.1539643, 
    0.1718906, 0.1725224, 0.1835196, 0.1538349, 0.1224362, 0.1671644, 
    0.1693291, 0.1670355, 0.1710259,
  0.09276105, 0.06473099, 0.04697023, 0.08625469, 0.07843497, 0.07239372, 
    0.08352, 0.0752356, 0.06035011, 0.04802502, 0.06760293, 0.077753, 
    0.07268056, 0.09373414, 0.09618025, 0.1036443, 0.09847694, 0.101402, 
    0.1066521, 0.1242614, 0.1222678, 0.1140842, 0.09815668, 0.08582975, 
    0.06779265, 0.08724938, 0.0995158, 0.1092375, 0.1061708,
  0.01083819, 0.01004447, 0.0460275, 0.04013501, 0.04427861, 0.05163255, 
    0.0270666, 0.01225395, 0.01445762, 0.0160717, 0.05346178, 0.05097998, 
    0.03996731, 0.0473128, 0.05730978, 0.07060794, 0.08628064, 0.1020478, 
    0.1359474, 0.07370157, 0.04385147, 0.01638953, 0.004976005, 0.008610032, 
    0.03798855, 0.07197479, 0.07473784, 0.03867488, 0.02884384,
  0.0005365951, 0.02000744, 0.03515081, 0.01813283, 0.04764612, 0.02710079, 
    0.02557168, 0.01850462, 0.01020379, 0.009252715, 0.0331997, 0.01542563, 
    0.02669113, 0.0499857, 0.06307241, 0.0692312, 0.0565685, 0.0517649, 
    0.02469272, 0.009784007, 0.0001964594, 0.0004678625, 2.796502e-06, 
    0.00680766, 0.03890625, 0.07398547, 0.02625844, 0.003768292, 0.0009569085,
  0.002178801, 0.04617408, 0.07509382, 0.04253298, 0.04081933, 0.03911937, 
    0.05503133, 0.05101112, 0.03398309, 0.02307667, 0.04006001, 0.03763157, 
    0.07781712, 0.06334102, 0.06748429, 0.04599001, 0.02746666, 0.0135503, 
    0.004777818, 0.001299943, 0.0001724189, 9.581313e-05, 0.00288096, 
    0.06071909, 0.1097621, 0.04723229, 0.009070025, 0.0001869124, 0.001125421,
  0.0771988, 0.09723968, 0.07285704, 0.01661922, 0.01937504, 0.03829701, 
    0.04096576, 0.03440711, 0.05374736, 0.1276141, 0.03705801, 0.03439632, 
    0.062163, 0.04560107, 0.03127537, 0.01092777, 0.007774895, 0.004284378, 
    0.007418736, 0.006142164, 0.009366875, 0.006417163, 0.05118828, 
    0.08664089, 0.07407168, 0.07778236, 0.0429573, 0.01802733, 0.02531534,
  0.03819723, 0.03773632, 0.04051504, 0.06283118, 0.0206129, 0.009937743, 
    0.02480907, 0.02621338, 0.05098223, 0.05320428, 0.0599281, 0.05965424, 
    0.0851398, 0.08270732, 0.05672547, 0.06876295, 0.07023044, 0.07098705, 
    0.08049975, 0.0992502, 0.1014375, 0.06390214, 0.05713368, 0.02406717, 
    0.02599235, 0.0311032, 0.03550064, 0.0563221, 0.06673644,
  0.0208188, 0.005436759, 0.003894157, 0.01053128, 0.01797086, 0.025966, 
    0.07809577, 0.0406406, 0.07673914, 0.04468583, 0.08078911, 0.06251456, 
    0.03973303, 0.02365334, 0.008473362, 0.01039603, 0.01497701, 0.01308411, 
    0.0186439, 0.01765956, 0.02430605, 0.04499006, 0.01208828, 0.0303937, 
    0.01175977, 0.01947153, 0.01318126, 0.01490337, 0.02406328,
  0.01821487, 0.02166955, 0.01486463, 0.02187276, 0.03043636, 0.0220165, 
    0.03770873, 0.08809128, 0.186722, 0.1193704, 0.09610298, 0.08724272, 
    0.09389116, 0.07325616, 0.06165728, 0.04949766, 0.03773124, 0.03988781, 
    0.02194496, 0.009769928, 0.02906605, 0.0387478, 0.05171576, 0.04372384, 
    0.04420562, 0.04057867, 0.02346842, 0.0154381, 0.02608284,
  0.06756523, 0.06808317, 0.06978179, 0.1007316, 0.06868736, 0.05763675, 
    0.1317503, 0.08317458, 0.07681349, 0.08711101, 0.1032006, 0.1086405, 
    0.1360295, 0.1589399, 0.1554407, 0.1644635, 0.1512306, 0.1284976, 
    0.06673028, 0.08429314, 0.1134885, 0.09039454, 0.1096613, 0.118771, 
    0.1337518, 0.1205841, 0.09030075, 0.05704322, 0.06012784,
  0.1310413, 0.1477171, 0.1320487, 0.136455, 0.1327884, 0.1382758, 0.1373857, 
    0.1329226, 0.1372024, 0.1424413, 0.1399722, 0.1458087, 0.1596995, 
    0.169551, 0.1770608, 0.1756784, 0.1811178, 0.1826754, 0.1677708, 
    0.1379828, 0.1200535, 0.1395691, 0.1684908, 0.1836471, 0.171469, 
    0.1647209, 0.1665275, 0.1491811, 0.1402639,
  0.1969768, 0.1875455, 0.1621545, 0.2041115, 0.2001373, 0.20288, 0.2155449, 
    0.2224881, 0.2108311, 0.189707, 0.1367833, 0.1249742, 0.1505601, 
    0.1920443, 0.1832254, 0.1987625, 0.2006679, 0.2690257, 0.2385793, 
    0.1672629, 0.1507773, 0.1782971, 0.1687741, 0.2045732, 0.2151584, 
    0.2449894, 0.1930598, 0.2179828, 0.2037814,
  0.2061206, 0.2009137, 0.2189036, 0.2044071, 0.2055629, 0.1977284, 
    0.2017846, 0.2117254, 0.1705034, 0.1741254, 0.1380288, 0.169068, 
    0.1645581, 0.1707233, 0.1836848, 0.1530526, 0.1770982, 0.1834595, 
    0.183166, 0.1801426, 0.1644524, 0.1257749, 0.1519806, 0.1356376, 
    0.1567979, 0.143325, 0.1036779, 0.2073877, 0.1937304,
  0.1601369, 0.1815825, 0.1671515, 0.1606026, 0.1486502, 0.1509933, 
    0.1475613, 0.1525166, 0.1453279, 0.1424928, 0.143907, 0.14583, 0.162112, 
    0.1793138, 0.1975631, 0.1940083, 0.1763132, 0.1573045, 0.1538396, 
    0.1517175, 0.1409123, 0.1481024, 0.1187245, 0.07298551, 0.1080677, 
    0.0698768, 0.07468978, 0.09805001, 0.1797225,
  0.007422621, 0.007148488, 0.006874355, 0.006600223, 0.00632609, 
    0.006051957, 0.005777824, 0.005908438, 0.005946374, 0.005984309, 
    0.006022244, 0.00606018, 0.006098115, 0.00613605, 0.005890391, 
    0.006173217, 0.006456044, 0.006738869, 0.007021695, 0.007304522, 
    0.007587348, 0.008179569, 0.00813294, 0.008086312, 0.008039683, 
    0.007993056, 0.007946426, 0.007899798, 0.007641927,
  0.02534367, 0.006702114, 0.001696978, 0.002233988, 0.002571383, 
    0.0009707591, 0.001137512, 0.001618928, 0.002200192, 0.00188823, 
    0.001732207, 0.004244455, 0.008555661, 0.1273396, 0.1256059, 0.1540394, 
    0.1871123, 0.2008377, 0.1527365, 0.1097778, 0.08791804, 0.07874002, 
    0.1534141, 0.2289787, 0.2070553, 0.1832155, 0.1977947, 0.1422815, 
    0.04857497,
  0.2115792, 0.2511179, 0.2370361, 0.244605, 0.1131037, 0.1045822, 0.1633856, 
    0.08917772, 0.07483654, 0.09298119, 0.09041721, 0.08636843, 0.1917316, 
    0.249325, 0.252007, 0.2364754, 0.2265848, 0.2462554, 0.2527341, 
    0.2514472, 0.2609571, 0.2808797, 0.3069225, 0.3283108, 0.30643, 
    0.2108778, 0.2155453, 0.2058181, 0.2368024,
  0.2203587, 0.238518, 0.2618552, 0.2619391, 0.2572669, 0.2454154, 0.2384244, 
    0.2412485, 0.2559933, 0.2651854, 0.2699933, 0.2808248, 0.2696922, 
    0.252963, 0.2307253, 0.2114595, 0.2145924, 0.2093963, 0.2229132, 
    0.2373811, 0.2443587, 0.2543772, 0.2524886, 0.2447212, 0.2459534, 
    0.2266448, 0.2116204, 0.2129954, 0.2283627,
  0.1790732, 0.1768561, 0.1817219, 0.1814146, 0.1665314, 0.167191, 0.1614859, 
    0.1742479, 0.1801844, 0.1935639, 0.1914026, 0.1793917, 0.1617761, 
    0.1513117, 0.142411, 0.1153624, 0.1286653, 0.1336741, 0.1446457, 
    0.1562195, 0.1678101, 0.1688482, 0.1771295, 0.1445419, 0.1173687, 
    0.1640052, 0.1645998, 0.1685787, 0.1721836,
  0.0902741, 0.06551985, 0.04722138, 0.08700632, 0.07787138, 0.07422905, 
    0.08265954, 0.07475064, 0.06259625, 0.0472271, 0.06763273, 0.07434329, 
    0.07366899, 0.0941428, 0.09489753, 0.1005547, 0.09204856, 0.09951898, 
    0.1060786, 0.1175779, 0.1157989, 0.1095764, 0.09519716, 0.08664254, 
    0.06715846, 0.08489207, 0.09581257, 0.1063886, 0.1061358,
  0.009068675, 0.007172556, 0.05482453, 0.04200176, 0.04458923, 0.05284205, 
    0.02395515, 0.01262641, 0.0144321, 0.01644595, 0.049693, 0.04911311, 
    0.04422856, 0.04726814, 0.05828068, 0.06856257, 0.0860956, 0.09857357, 
    0.1280918, 0.07264362, 0.04613004, 0.01887826, 0.005795782, 0.0081046, 
    0.04454057, 0.07590405, 0.07666389, 0.04000753, 0.0299661,
  0.00108596, 0.02665101, 0.04468128, 0.02056697, 0.05696798, 0.0322838, 
    0.0285287, 0.02024474, 0.01174343, 0.01267443, 0.04707265, 0.02469691, 
    0.02874683, 0.05294197, 0.06789352, 0.0735355, 0.05994006, 0.05813102, 
    0.02636703, 0.01070788, 0.0002090632, 0.0008765445, 7.080131e-06, 
    0.005229016, 0.04943157, 0.08048562, 0.02759547, 0.002480116, 0.00115735,
  0.003509799, 0.05975186, 0.09029039, 0.05371441, 0.04673508, 0.04901636, 
    0.06549032, 0.058766, 0.03986378, 0.02965474, 0.04763729, 0.04601106, 
    0.09508272, 0.07679048, 0.08092115, 0.05121797, 0.03270031, 0.01583583, 
    0.005275145, 0.001664274, 0.0002267232, 0.0009866136, 0.002768604, 
    0.07400404, 0.1308077, 0.05680446, 0.01019973, 0.0003128487, 0.002166609,
  0.1046884, 0.1186353, 0.1008433, 0.01807606, 0.01892766, 0.04083135, 
    0.04473038, 0.04131599, 0.06894096, 0.144552, 0.0482545, 0.04296637, 
    0.07338797, 0.0530955, 0.0336233, 0.01225399, 0.009275354, 0.005175137, 
    0.007301388, 0.005199992, 0.01014651, 0.01340545, 0.06122793, 0.1066796, 
    0.08401549, 0.08214294, 0.04781925, 0.01827398, 0.03956863,
  0.04171163, 0.04521495, 0.04547415, 0.1006631, 0.0234182, 0.01178179, 
    0.03159696, 0.03318077, 0.06610785, 0.0681238, 0.07752449, 0.07244221, 
    0.1006049, 0.09655121, 0.0687599, 0.08098315, 0.07788118, 0.08109698, 
    0.0929032, 0.1126124, 0.11392, 0.07441691, 0.06847479, 0.03149239, 
    0.03042031, 0.03749523, 0.04285011, 0.06734078, 0.07957826,
  0.0154945, 0.003435777, 0.003147638, 0.00955754, 0.01844067, 0.02572541, 
    0.09254231, 0.05321578, 0.09367272, 0.0570376, 0.09319232, 0.07217367, 
    0.04766472, 0.02593175, 0.01122451, 0.0117612, 0.01518578, 0.01421484, 
    0.0138086, 0.01812014, 0.0290522, 0.05280009, 0.01680795, 0.03536144, 
    0.01344326, 0.02329358, 0.01420524, 0.01423567, 0.02195047,
  0.01115731, 0.01836392, 0.01054145, 0.01534814, 0.03322303, 0.02165565, 
    0.04142767, 0.1010056, 0.2046346, 0.1250696, 0.1013437, 0.09587873, 
    0.09986614, 0.07448471, 0.06316616, 0.05103333, 0.03667038, 0.04048333, 
    0.01767577, 0.008057208, 0.03225887, 0.03954023, 0.05516816, 0.04515402, 
    0.04466695, 0.03917768, 0.02459372, 0.01351926, 0.02417888,
  0.05860378, 0.06109839, 0.06862577, 0.1026901, 0.06326588, 0.05038814, 
    0.1456062, 0.06712641, 0.06390502, 0.08390649, 0.1008405, 0.1030358, 
    0.130225, 0.1553346, 0.1529405, 0.1630237, 0.1489679, 0.1213212, 
    0.06395063, 0.08015204, 0.1104601, 0.08687006, 0.1077873, 0.1190931, 
    0.1308798, 0.117896, 0.08535763, 0.0552047, 0.0571879,
  0.1233127, 0.1455288, 0.1336099, 0.1382493, 0.1281042, 0.1361106, 0.132188, 
    0.1488757, 0.153944, 0.1429226, 0.1408131, 0.1506748, 0.1646786, 
    0.1740371, 0.1784294, 0.1750199, 0.1749977, 0.1774203, 0.1620014, 
    0.1458472, 0.1258123, 0.1356723, 0.1696982, 0.1967191, 0.1796551, 
    0.1652202, 0.1616371, 0.1456753, 0.1380903,
  0.1943552, 0.1919188, 0.1617893, 0.2040531, 0.2082175, 0.2092282, 
    0.2167988, 0.2289016, 0.22942, 0.2112539, 0.1580608, 0.1455369, 
    0.1802686, 0.2024294, 0.1865547, 0.1975813, 0.2053417, 0.278027, 
    0.2525435, 0.1721633, 0.1525956, 0.1809524, 0.1847146, 0.227514, 
    0.2282507, 0.2624572, 0.1872742, 0.2158802, 0.2032795,
  0.2040617, 0.1951134, 0.23411, 0.2122668, 0.2157027, 0.2108497, 0.2207782, 
    0.2380391, 0.1970944, 0.1944168, 0.1604635, 0.1875486, 0.1762725, 
    0.1870321, 0.1884182, 0.1632043, 0.189325, 0.188012, 0.1900994, 
    0.1869986, 0.1746948, 0.1482639, 0.170469, 0.1539315, 0.176082, 0.175192, 
    0.1363289, 0.2098215, 0.1902698,
  0.1565621, 0.1850236, 0.1759783, 0.1711969, 0.1617596, 0.1621216, 
    0.1670528, 0.1771619, 0.1723423, 0.1725935, 0.1622618, 0.1701828, 
    0.1862836, 0.1970178, 0.2166635, 0.2069457, 0.1952601, 0.1810436, 
    0.1731256, 0.1712961, 0.159151, 0.1718682, 0.1459301, 0.08843762, 
    0.1287199, 0.08400529, 0.09809693, 0.1266748, 0.1806637,
  0.01756209, 0.01687397, 0.01618586, 0.01549774, 0.01480962, 0.01412151, 
    0.01343339, 0.0162074, 0.01654152, 0.01687564, 0.01720976, 0.01754387, 
    0.01787799, 0.01821211, 0.01482039, 0.01574801, 0.01667562, 0.01760323, 
    0.01853084, 0.01945845, 0.02038606, 0.02274762, 0.02217401, 0.0216004, 
    0.02102678, 0.02045317, 0.01987956, 0.01930595, 0.01811258,
  0.04826006, 0.02261262, 0.006581211, 0.00490777, 0.003915946, 0.002846458, 
    0.003697555, 0.003982069, 0.003527407, 0.003945148, 0.006390993, 
    0.01448322, 0.03027052, 0.1553456, 0.1323955, 0.1617892, 0.2017801, 
    0.223304, 0.1865774, 0.1639522, 0.1417627, 0.1436327, 0.2076533, 
    0.2312918, 0.2105405, 0.1889666, 0.2095964, 0.1773098, 0.07287292,
  0.2201645, 0.263398, 0.2456619, 0.2642938, 0.1529751, 0.1353295, 0.183714, 
    0.1335103, 0.1142038, 0.1511529, 0.1471316, 0.1389088, 0.2143564, 
    0.2521565, 0.2570021, 0.2412636, 0.2346036, 0.2560986, 0.2734327, 
    0.2649296, 0.2754443, 0.2936639, 0.3089631, 0.3459659, 0.3092973, 
    0.2130724, 0.2175902, 0.2089079, 0.2446986,
  0.228825, 0.2454094, 0.2687935, 0.2747681, 0.2683025, 0.2518712, 0.2444603, 
    0.2520776, 0.2627591, 0.279809, 0.2755463, 0.2843324, 0.2671428, 
    0.2499044, 0.2292875, 0.2113715, 0.2163564, 0.2154972, 0.2317551, 
    0.2435867, 0.2559065, 0.2435339, 0.2573499, 0.2498725, 0.2468521, 
    0.2268587, 0.2126023, 0.2100016, 0.2299472,
  0.1842051, 0.1763914, 0.1823958, 0.1810513, 0.1690594, 0.1683002, 
    0.1582529, 0.1762044, 0.1824213, 0.1948307, 0.1970332, 0.1826064, 
    0.1653224, 0.1564724, 0.1394802, 0.1178363, 0.1269543, 0.133305, 
    0.1388249, 0.1572106, 0.1697837, 0.1691867, 0.1752451, 0.1394053, 
    0.1164774, 0.1589944, 0.1606648, 0.1648274, 0.1709131,
  0.08802799, 0.06898338, 0.0492741, 0.08872716, 0.08045436, 0.07691658, 
    0.08534561, 0.07845351, 0.06513552, 0.05368691, 0.06835929, 0.07498382, 
    0.07664598, 0.09420988, 0.09939541, 0.09671782, 0.09095449, 0.09516281, 
    0.1075794, 0.1155295, 0.1154668, 0.105054, 0.08899631, 0.08908813, 
    0.06673743, 0.08554889, 0.09731698, 0.1057801, 0.1075982,
  0.009821498, 0.005869183, 0.0634885, 0.04593202, 0.04879292, 0.05850254, 
    0.02481421, 0.01495932, 0.01575778, 0.01818813, 0.04928083, 0.04446537, 
    0.04992283, 0.04976469, 0.06201623, 0.07047619, 0.0854509, 0.09899592, 
    0.127054, 0.07872801, 0.05477814, 0.02166338, 0.008061595, 0.007243865, 
    0.05451326, 0.08226001, 0.08241385, 0.04191593, 0.02836642,
  0.0008039656, 0.03474992, 0.05702279, 0.02237349, 0.06670776, 0.03877874, 
    0.0337477, 0.02109742, 0.01260827, 0.01523023, 0.05219074, 0.02909862, 
    0.02976533, 0.05392888, 0.07144183, 0.08038469, 0.06577066, 0.06831785, 
    0.03319342, 0.01284903, 0.0009657708, 0.0005551318, 6.960446e-06, 
    0.003000912, 0.06470038, 0.09123552, 0.02891023, 0.002296569, 0.0009812356,
  0.004005471, 0.06429042, 0.1235706, 0.06747355, 0.05259541, 0.05719901, 
    0.07480391, 0.06551962, 0.04663342, 0.03475803, 0.05254593, 0.05425696, 
    0.109683, 0.08832257, 0.09004659, 0.05860305, 0.03589891, 0.01827728, 
    0.006126883, 0.001628728, 0.0001910126, 0.002116061, 0.004555415, 
    0.09408663, 0.1548672, 0.08220341, 0.01143258, 0.0003408639, 0.001059186,
  0.1108129, 0.1493295, 0.1349574, 0.02039864, 0.01857509, 0.04302119, 
    0.04992072, 0.04953813, 0.09207074, 0.1766745, 0.05658458, 0.05030837, 
    0.08221279, 0.05974108, 0.03659189, 0.01361175, 0.009322271, 0.006322744, 
    0.008680991, 0.007047118, 0.01149194, 0.01642951, 0.07849266, 0.1395393, 
    0.1042996, 0.08236647, 0.05030107, 0.01929221, 0.03690055,
  0.05210212, 0.05457017, 0.05198278, 0.1396786, 0.02398582, 0.01404831, 
    0.03856259, 0.04151028, 0.07755984, 0.0734556, 0.09372776, 0.08162843, 
    0.1126696, 0.1036645, 0.07973924, 0.0873493, 0.08432577, 0.09092755, 
    0.1002905, 0.126404, 0.1270871, 0.08257824, 0.08289642, 0.04134156, 
    0.03470881, 0.04295624, 0.04833503, 0.07785101, 0.09546477,
  0.01012743, 0.002645848, 0.003606984, 0.007861521, 0.01770275, 0.02064744, 
    0.1105155, 0.05487113, 0.1163619, 0.06413679, 0.09835643, 0.07674334, 
    0.05108735, 0.02965962, 0.01375445, 0.01371687, 0.01816364, 0.01435837, 
    0.01216203, 0.01917381, 0.03539129, 0.06187076, 0.01935791, 0.04315297, 
    0.01557805, 0.02617813, 0.01404986, 0.01242321, 0.01574441,
  0.004736083, 0.01358462, 0.008624622, 0.0114065, 0.03530217, 0.02155355, 
    0.03606546, 0.1107265, 0.2141751, 0.1302343, 0.1037762, 0.09762383, 
    0.1072085, 0.0801406, 0.06888262, 0.05355155, 0.03819608, 0.04011725, 
    0.01672585, 0.007113572, 0.03636874, 0.0425549, 0.05715384, 0.04945235, 
    0.05124722, 0.04241163, 0.02438927, 0.01256556, 0.02036886,
  0.05282471, 0.05454555, 0.06831034, 0.1063835, 0.06239506, 0.04355555, 
    0.1474205, 0.05176542, 0.04951718, 0.08086246, 0.1005182, 0.09837694, 
    0.1298461, 0.156414, 0.1580376, 0.1635547, 0.1472316, 0.1185264, 
    0.06399214, 0.07823041, 0.1023874, 0.08769617, 0.1069336, 0.1226722, 
    0.1335776, 0.1186234, 0.09013933, 0.05423924, 0.05854662,
  0.1251124, 0.148378, 0.1340408, 0.1388781, 0.1265395, 0.1339251, 0.1319666, 
    0.1566759, 0.1535438, 0.1384305, 0.1388646, 0.1519459, 0.1612452, 
    0.178403, 0.1848112, 0.1744949, 0.177696, 0.1777908, 0.1639918, 
    0.1500425, 0.1254116, 0.1329095, 0.173727, 0.2067339, 0.1871134, 
    0.1672418, 0.164983, 0.147824, 0.137856,
  0.1909328, 0.1924043, 0.1639257, 0.2120339, 0.211417, 0.2125121, 0.2165183, 
    0.2329732, 0.2332801, 0.2223408, 0.1730318, 0.1558388, 0.1953607, 
    0.2082931, 0.1900901, 0.2057595, 0.2079546, 0.2883898, 0.2569694, 
    0.1756404, 0.1548976, 0.1826693, 0.1965119, 0.2467655, 0.2407809, 
    0.2714291, 0.1903015, 0.2158039, 0.2044064,
  0.2058859, 0.1931008, 0.2332031, 0.216776, 0.2283751, 0.2239674, 0.2230067, 
    0.2607396, 0.2170021, 0.206975, 0.176194, 0.1967795, 0.1887887, 0.185518, 
    0.1920472, 0.1593007, 0.1915372, 0.1906601, 0.193508, 0.1911264, 
    0.183877, 0.1566464, 0.1726137, 0.1757301, 0.1750923, 0.2149514, 
    0.1661966, 0.2080906, 0.1891309,
  0.1536288, 0.1891449, 0.179051, 0.1761023, 0.1795803, 0.177439, 0.1773094, 
    0.1886157, 0.1838712, 0.1880568, 0.1797068, 0.1892571, 0.1945692, 
    0.2116169, 0.2237637, 0.2125008, 0.2112289, 0.1968283, 0.183862, 
    0.1905254, 0.1772956, 0.1955898, 0.1735129, 0.1024197, 0.1388349, 
    0.1005748, 0.1206911, 0.1312128, 0.1819614,
  0.03771275, 0.03617186, 0.03463098, 0.0330901, 0.03154921, 0.03000833, 
    0.02846744, 0.03101798, 0.03229271, 0.03356743, 0.03484215, 0.03611687, 
    0.0373916, 0.03866632, 0.03630328, 0.03789236, 0.03948143, 0.04107051, 
    0.04265959, 0.04424866, 0.04583774, 0.04952262, 0.0481997, 0.04687679, 
    0.04555387, 0.04423096, 0.04290804, 0.04158513, 0.03894546,
  0.06625129, 0.04184896, 0.02502471, 0.0119102, 0.01032039, 0.007673877, 
    0.00700963, 0.006884492, 0.00721173, 0.01191936, 0.01570923, 0.0378049, 
    0.06217385, 0.1681136, 0.1357275, 0.1696111, 0.208427, 0.2394383, 
    0.2060132, 0.2023216, 0.206453, 0.219477, 0.234778, 0.231329, 0.2092435, 
    0.1899293, 0.209975, 0.1934554, 0.1117949,
  0.2336045, 0.277128, 0.2575918, 0.2784199, 0.1956915, 0.1573725, 0.2024365, 
    0.1738344, 0.1584074, 0.1978851, 0.1929239, 0.178268, 0.2267245, 
    0.2610413, 0.2689953, 0.2483005, 0.259158, 0.2741028, 0.2792764, 
    0.2797318, 0.2867342, 0.3031455, 0.307409, 0.3543823, 0.311756, 
    0.2085983, 0.211472, 0.2180771, 0.2441964,
  0.2498214, 0.2647416, 0.2865925, 0.2957919, 0.2912722, 0.2689672, 
    0.2693313, 0.2747593, 0.2800973, 0.2852068, 0.2777813, 0.2858875, 
    0.2699352, 0.2536242, 0.2329228, 0.2143224, 0.217156, 0.2200348, 
    0.2338219, 0.2497526, 0.2584954, 0.2493044, 0.2626164, 0.2473247, 
    0.2411982, 0.230423, 0.2185725, 0.2212216, 0.2449276,
  0.1925626, 0.1805296, 0.1881725, 0.1835693, 0.1754532, 0.1722577, 
    0.1631305, 0.1888794, 0.1900987, 0.1959547, 0.2079566, 0.192121, 
    0.1676366, 0.153303, 0.1324696, 0.11834, 0.1276789, 0.1374565, 0.1453464, 
    0.1599739, 0.1698727, 0.1732599, 0.1703035, 0.1393122, 0.1185308, 
    0.1519392, 0.1578313, 0.1643762, 0.1738453,
  0.09407051, 0.07384305, 0.05253049, 0.08895739, 0.08469224, 0.08033465, 
    0.08633253, 0.08344982, 0.07114266, 0.05645365, 0.06815728, 0.07631499, 
    0.07855573, 0.09725914, 0.1045018, 0.09812, 0.0956068, 0.09841511, 
    0.1083001, 0.1168856, 0.116477, 0.1051652, 0.09090292, 0.09183424, 
    0.06829081, 0.08630253, 0.1005735, 0.1089782, 0.1134555,
  0.01156762, 0.005460331, 0.06972218, 0.04817171, 0.05151823, 0.0638376, 
    0.02838927, 0.01706651, 0.0173937, 0.01686399, 0.04185669, 0.03456, 
    0.0598921, 0.05540905, 0.06660045, 0.07537586, 0.0898528, 0.1015798, 
    0.1289585, 0.08681747, 0.06412076, 0.02568258, 0.00995873, 0.005228465, 
    0.06245402, 0.09046029, 0.08753652, 0.04581584, 0.03122982,
  0.0003321955, 0.03853837, 0.06641412, 0.02217774, 0.06529088, 0.0369569, 
    0.0361252, 0.02147827, 0.01152478, 0.01216367, 0.0463423, 0.03009683, 
    0.02904659, 0.05168009, 0.06620118, 0.0763637, 0.06594744, 0.06834443, 
    0.0395062, 0.01475978, 0.002626959, 0.000714294, 2.777138e-06, 
    0.0007864711, 0.06192946, 0.1076991, 0.02973076, 0.002544144, 0.0001157123,
  0.002061879, 0.04677938, 0.1562539, 0.07286182, 0.05052081, 0.05681917, 
    0.07041115, 0.06328476, 0.04158138, 0.02842994, 0.05060377, 0.04110302, 
    0.1017531, 0.07337114, 0.07745177, 0.05594182, 0.03607804, 0.0201698, 
    0.006239517, 0.001431203, 0.000362815, 0.002850781, 0.002444522, 
    0.09936209, 0.150947, 0.1155559, 0.01208116, 0.0003705427, 0.0005030496,
  0.08418878, 0.1744018, 0.1489659, 0.02455025, 0.01760865, 0.04050793, 
    0.04945447, 0.04550563, 0.1021896, 0.197084, 0.05261476, 0.0372333, 
    0.06698601, 0.0496968, 0.03225757, 0.01312601, 0.008844109, 0.006137733, 
    0.009361298, 0.00573546, 0.00951426, 0.01654025, 0.08270752, 0.1561024, 
    0.1180596, 0.07704449, 0.0495882, 0.01807356, 0.02730206,
  0.04766656, 0.05500847, 0.05132781, 0.1655799, 0.01944602, 0.01314005, 
    0.0403972, 0.03475886, 0.05535627, 0.05944141, 0.08332347, 0.06490962, 
    0.08801449, 0.0874692, 0.07116771, 0.08087278, 0.08295289, 0.09308451, 
    0.102018, 0.1261454, 0.1220871, 0.0728531, 0.08993304, 0.04468165, 
    0.03196057, 0.04446087, 0.0443991, 0.06599475, 0.1035453,
  0.003377738, 0.00147415, 0.00189133, 0.005972756, 0.01059077, 0.0132905, 
    0.09402727, 0.04683832, 0.1295063, 0.05792759, 0.08984658, 0.06622984, 
    0.04065428, 0.02610013, 0.01409552, 0.01473221, 0.02132485, 0.01410852, 
    0.01219732, 0.02066359, 0.02916029, 0.06585734, 0.01892837, 0.04133172, 
    0.01776093, 0.02904155, 0.01283013, 0.01189577, 0.009194355,
  0.002163046, 0.009463666, 0.007433772, 0.01157159, 0.03739349, 0.02114662, 
    0.02977524, 0.1235161, 0.2284458, 0.130163, 0.1015672, 0.09173415, 
    0.1028704, 0.07735186, 0.0738002, 0.05653208, 0.04103236, 0.0408811, 
    0.01664959, 0.007331521, 0.03858173, 0.04264878, 0.05518796, 0.0515006, 
    0.05678469, 0.04594596, 0.0266883, 0.01217113, 0.01549431,
  0.04958984, 0.04693864, 0.07213498, 0.1124536, 0.06203427, 0.037953, 
    0.1452331, 0.0383538, 0.03632897, 0.07766164, 0.1023675, 0.09375542, 
    0.1292094, 0.1580064, 0.163871, 0.1708286, 0.1495459, 0.1217324, 
    0.06408697, 0.0800334, 0.09904209, 0.08252735, 0.1095503, 0.1246176, 
    0.1367097, 0.120064, 0.09600458, 0.05672308, 0.06133316,
  0.122543, 0.1450876, 0.1402373, 0.1432164, 0.1212916, 0.1305554, 0.1304768, 
    0.1632178, 0.1463319, 0.1342312, 0.1408458, 0.1538175, 0.1633764, 
    0.181572, 0.1967515, 0.1835799, 0.1819783, 0.182597, 0.1649178, 
    0.1529281, 0.1278113, 0.1333866, 0.186125, 0.2115906, 0.1962374, 
    0.1712429, 0.1691822, 0.1507521, 0.1405381,
  0.1917513, 0.2010349, 0.1775739, 0.2176452, 0.2189263, 0.2163532, 
    0.2185565, 0.2393054, 0.2371356, 0.2319681, 0.1870613, 0.1634099, 
    0.2075216, 0.2199922, 0.1907946, 0.2117994, 0.2102271, 0.3118379, 
    0.2588087, 0.1756828, 0.160233, 0.1976755, 0.207542, 0.2568465, 
    0.2367531, 0.2734598, 0.1982268, 0.2236892, 0.2120266,
  0.2138517, 0.1963115, 0.2445655, 0.2302436, 0.230366, 0.2277985, 0.2289491, 
    0.2713437, 0.2238183, 0.2165266, 0.1875954, 0.2067016, 0.1999752, 
    0.1880407, 0.1999096, 0.1658569, 0.1945955, 0.1978537, 0.1897619, 
    0.2004152, 0.1870156, 0.1640158, 0.1798235, 0.1871025, 0.1789667, 
    0.2505927, 0.1974861, 0.2092463, 0.1919248,
  0.1548668, 0.1842711, 0.1809694, 0.17631, 0.1798757, 0.1764231, 0.1800101, 
    0.1963397, 0.1971461, 0.2008248, 0.1937204, 0.202864, 0.2001184, 
    0.2127944, 0.2227845, 0.2179116, 0.2060953, 0.198417, 0.1907424, 
    0.2007883, 0.1938364, 0.2159242, 0.1904802, 0.1143385, 0.1412098, 
    0.1132816, 0.1335687, 0.1427082, 0.1864925,
  0.06248819, 0.06117525, 0.0598623, 0.05854936, 0.05723641, 0.05592347, 
    0.05461052, 0.05558119, 0.05747441, 0.05936763, 0.06126085, 0.06315406, 
    0.06504729, 0.06694051, 0.06909335, 0.07053878, 0.07198421, 0.07342964, 
    0.07487506, 0.07632049, 0.07776592, 0.077092, 0.0750663, 0.0730406, 
    0.0710149, 0.06898919, 0.06696349, 0.06493779, 0.06353855,
  0.09972171, 0.05361447, 0.04589437, 0.02862191, 0.0224047, 0.02302107, 
    0.01943078, 0.0159275, 0.02201193, 0.02905031, 0.03991574, 0.05861851, 
    0.09311652, 0.1759042, 0.1373644, 0.1883542, 0.2134421, 0.2493093, 
    0.2120859, 0.2239629, 0.2556442, 0.2985866, 0.2511481, 0.2381259, 
    0.2141496, 0.1913963, 0.2121765, 0.1980904, 0.1417432,
  0.2470183, 0.2871639, 0.2717116, 0.2939829, 0.23209, 0.1732569, 0.220635, 
    0.2176729, 0.1978393, 0.2359666, 0.2261956, 0.2045, 0.231825, 0.276183, 
    0.2863812, 0.2700339, 0.2708738, 0.3030518, 0.3073747, 0.3079051, 
    0.3136193, 0.3289235, 0.3285919, 0.3772796, 0.311575, 0.2154856, 
    0.2323955, 0.2465415, 0.2629292,
  0.2717269, 0.286299, 0.3037178, 0.3142141, 0.2965898, 0.2843614, 0.2811011, 
    0.2936485, 0.3033002, 0.3083467, 0.3006425, 0.2947327, 0.2755526, 
    0.2525787, 0.2402701, 0.2172596, 0.2235728, 0.2278599, 0.2500004, 
    0.2598787, 0.2691372, 0.2593302, 0.2672852, 0.2460022, 0.2398368, 
    0.2342142, 0.2309932, 0.2330094, 0.2636481,
  0.2029096, 0.1890793, 0.1951804, 0.192471, 0.1795984, 0.1806124, 0.1726629, 
    0.1985477, 0.2009693, 0.2076741, 0.2152784, 0.1952671, 0.170279, 
    0.1566159, 0.1359896, 0.1249882, 0.1324916, 0.145172, 0.1545098, 
    0.1658248, 0.1755946, 0.1746667, 0.1713488, 0.1435734, 0.1172731, 
    0.1525428, 0.1608631, 0.1656089, 0.177062,
  0.1043875, 0.08451491, 0.05859369, 0.08972212, 0.09419613, 0.09012246, 
    0.09328934, 0.08793461, 0.07871348, 0.06456904, 0.06934004, 0.07546654, 
    0.08178591, 0.1050137, 0.1133734, 0.1048554, 0.1039043, 0.1038413, 
    0.1118499, 0.1171279, 0.1211537, 0.1078286, 0.09366461, 0.09632701, 
    0.0660854, 0.09065822, 0.1066681, 0.1169131, 0.1211022,
  0.01427313, 0.005863723, 0.07316518, 0.046428, 0.05489869, 0.06555878, 
    0.03355631, 0.01876937, 0.01842725, 0.01672791, 0.02903722, 0.0238807, 
    0.06603723, 0.05984174, 0.06990135, 0.08069483, 0.09136869, 0.1022638, 
    0.130463, 0.09312157, 0.07378553, 0.03239635, 0.01307776, 0.004132629, 
    0.06102088, 0.08689255, 0.09006228, 0.05302449, 0.0336314,
  0.0002152855, 0.03345763, 0.06336938, 0.0219683, 0.06196026, 0.03616617, 
    0.03767033, 0.02085277, 0.01062066, 0.008480151, 0.03409719, 0.02617427, 
    0.0302433, 0.05135109, 0.06413097, 0.0692864, 0.0635092, 0.06184686, 
    0.04495233, 0.02212941, 0.005283247, 0.0009107823, 9.253504e-07, 
    0.0002134513, 0.05721034, 0.1168083, 0.02916058, 0.003497737, 0.0002377049,
  0.0007583351, 0.02773356, 0.1594068, 0.06501777, 0.04832049, 0.05345972, 
    0.06283461, 0.06043269, 0.03773471, 0.02378243, 0.04607693, 0.03445238, 
    0.09962532, 0.06434402, 0.06876759, 0.05327983, 0.0375714, 0.02184366, 
    0.007443334, 0.001465049, 0.0007505909, 0.00141928, 0.001340493, 
    0.07116834, 0.1103808, 0.08933791, 0.01461687, 0.0005358225, 5.204256e-05,
  0.05435039, 0.1408775, 0.1046855, 0.02981816, 0.01615379, 0.03738218, 
    0.0464172, 0.03965524, 0.08986565, 0.1730268, 0.0493408, 0.02856272, 
    0.05632148, 0.04322187, 0.02888097, 0.01328587, 0.009306072, 0.005397687, 
    0.008178738, 0.005556967, 0.009902939, 0.01347215, 0.07814438, 0.1332145, 
    0.125049, 0.06959839, 0.05076089, 0.01739288, 0.01875872,
  0.02760099, 0.03379815, 0.03106176, 0.2101593, 0.0201856, 0.01270706, 
    0.04269899, 0.03048518, 0.04470924, 0.050124, 0.07983535, 0.05511988, 
    0.07205174, 0.07493933, 0.06532604, 0.07460198, 0.077092, 0.08976854, 
    0.09994499, 0.1243464, 0.1139385, 0.06639198, 0.08683498, 0.0420712, 
    0.02952783, 0.03806372, 0.03923727, 0.05028272, 0.07385956,
  0.0009717622, 0.0005018669, 0.00172639, 0.005305208, 0.007588834, 
    0.008807587, 0.08143981, 0.04605162, 0.1148769, 0.05425129, 0.08908689, 
    0.05626121, 0.03540946, 0.02301473, 0.01535379, 0.01625132, 0.02149758, 
    0.0154544, 0.0124612, 0.01687939, 0.02026668, 0.07047766, 0.01772971, 
    0.03524571, 0.01970911, 0.03043957, 0.008641594, 0.007096334, 0.003637397,
  0.001560042, 0.007885139, 0.0074807, 0.01219049, 0.03932328, 0.01972284, 
    0.0253748, 0.13483, 0.2462751, 0.1289627, 0.09431675, 0.0893626, 
    0.1001857, 0.07392016, 0.07538939, 0.06066783, 0.0464872, 0.04450276, 
    0.01991993, 0.008571599, 0.03604229, 0.0425871, 0.05293014, 0.04902544, 
    0.05747569, 0.04861353, 0.02826135, 0.01198397, 0.01161754,
  0.04778287, 0.04391662, 0.07450632, 0.1231748, 0.0609391, 0.03245802, 
    0.14166, 0.03038426, 0.02685378, 0.0740606, 0.1012325, 0.09233991, 
    0.1312213, 0.1598144, 0.1585798, 0.1735674, 0.1533967, 0.1280501, 
    0.06824152, 0.08387569, 0.09992357, 0.0791922, 0.1125594, 0.1214727, 
    0.1386383, 0.1256041, 0.1006299, 0.06251521, 0.06547098,
  0.1249944, 0.154755, 0.1439288, 0.1545988, 0.1230343, 0.1285605, 0.1300516, 
    0.172004, 0.1402159, 0.1309326, 0.143416, 0.1571082, 0.1627708, 
    0.1918926, 0.2101446, 0.1960876, 0.1870312, 0.1889899, 0.1696599, 
    0.161154, 0.1370065, 0.1321121, 0.1891468, 0.2299008, 0.1986921, 
    0.1730564, 0.1765801, 0.1624431, 0.144758,
  0.2008184, 0.2071722, 0.1850925, 0.2271444, 0.2378316, 0.2275995, 
    0.2357478, 0.2541883, 0.2456689, 0.2476025, 0.2027183, 0.176622, 
    0.220532, 0.2338742, 0.2049075, 0.2204668, 0.221466, 0.3326774, 
    0.2692848, 0.1797501, 0.1693784, 0.2035162, 0.218031, 0.2623322, 
    0.2414947, 0.2757565, 0.2066837, 0.2245956, 0.2163941,
  0.2243326, 0.2058957, 0.2554854, 0.2406893, 0.2516364, 0.2510925, 
    0.2405775, 0.2803384, 0.2345601, 0.2266645, 0.1992686, 0.2072844, 
    0.1991023, 0.1972531, 0.2071442, 0.1715771, 0.2071116, 0.2082052, 
    0.1878179, 0.2076273, 0.19631, 0.1779822, 0.202395, 0.2011352, 0.1701208, 
    0.2855695, 0.2308803, 0.2206706, 0.206161,
  0.1700366, 0.2028525, 0.2024681, 0.1894334, 0.1850802, 0.1819192, 
    0.1909689, 0.2139295, 0.2065345, 0.2050672, 0.1962009, 0.2082506, 
    0.2159449, 0.2228383, 0.2442311, 0.2319909, 0.2167285, 0.2015826, 
    0.2070294, 0.2087603, 0.1998646, 0.2222813, 0.2063152, 0.1297778, 
    0.144584, 0.1207412, 0.1438167, 0.1439582, 0.1986989,
  0.0887723, 0.08673253, 0.08469276, 0.082653, 0.08061323, 0.07857347, 
    0.0765337, 0.08157372, 0.08402761, 0.0864815, 0.0889354, 0.09138929, 
    0.09384318, 0.09629708, 0.0925364, 0.09549689, 0.09845739, 0.1014179, 
    0.1043784, 0.1073389, 0.1102994, 0.1091528, 0.1057782, 0.1024036, 
    0.09902894, 0.09565432, 0.09227969, 0.08890507, 0.09040411,
  0.1337874, 0.07650184, 0.05829519, 0.05173636, 0.04006158, 0.04691411, 
    0.03928802, 0.03612028, 0.03182587, 0.04510874, 0.05471575, 0.08193554, 
    0.1197092, 0.17246, 0.12701, 0.1701477, 0.2060861, 0.2418414, 0.2172634, 
    0.226634, 0.2834637, 0.3440051, 0.2588681, 0.2387912, 0.2111145, 
    0.1891304, 0.2128551, 0.202655, 0.1611433,
  0.2598282, 0.2993932, 0.2800763, 0.309696, 0.2595056, 0.1886495, 0.2311267, 
    0.2495252, 0.23202, 0.2613905, 0.2591676, 0.2198443, 0.2367686, 
    0.2874609, 0.2956126, 0.2928974, 0.2844384, 0.2923539, 0.3237986, 
    0.3222379, 0.3286092, 0.3317793, 0.3423442, 0.4056809, 0.3116997, 
    0.2174477, 0.2340066, 0.259419, 0.2728394,
  0.292349, 0.3159141, 0.3341655, 0.335557, 0.3235181, 0.3092568, 0.3054551, 
    0.3200962, 0.3311612, 0.3294865, 0.3222361, 0.3068288, 0.2933802, 
    0.272696, 0.2658744, 0.2414981, 0.2454746, 0.2507512, 0.274963, 
    0.2913807, 0.2951179, 0.2692911, 0.2722578, 0.2668699, 0.2537916, 
    0.2480335, 0.2424442, 0.2404481, 0.2805095,
  0.2205735, 0.2059181, 0.213133, 0.2062561, 0.1894955, 0.1876372, 0.1847294, 
    0.210824, 0.2087542, 0.2216042, 0.2285276, 0.2039158, 0.1800805, 
    0.1661306, 0.1389285, 0.1393862, 0.1469559, 0.1648533, 0.1722541, 
    0.1785938, 0.1952301, 0.1844574, 0.1850831, 0.153582, 0.1212588, 
    0.1558377, 0.1707403, 0.1782092, 0.1918757,
  0.1204225, 0.09727446, 0.07024211, 0.09656464, 0.1067531, 0.1007301, 
    0.1092229, 0.1046097, 0.090652, 0.07928413, 0.07911848, 0.07880057, 
    0.08752459, 0.1139337, 0.1289159, 0.1160539, 0.1175213, 0.1114156, 
    0.1191406, 0.1226377, 0.1288679, 0.1206837, 0.1040852, 0.102442, 
    0.06579927, 0.0982381, 0.1161689, 0.1261563, 0.1305358,
  0.02008877, 0.007183479, 0.07491576, 0.04187147, 0.05290506, 0.06605349, 
    0.03927877, 0.02516218, 0.02175512, 0.0165196, 0.01814302, 0.01606726, 
    0.07164229, 0.06166971, 0.07605848, 0.08821889, 0.09887533, 0.1044384, 
    0.1258231, 0.09696534, 0.08129454, 0.04303405, 0.01809376, 0.003286687, 
    0.05608121, 0.08914217, 0.08902703, 0.0569353, 0.04221153,
  0.0002508654, 0.02490235, 0.05655398, 0.024037, 0.06686912, 0.03945385, 
    0.04056542, 0.0264082, 0.01279284, 0.009130514, 0.02496472, 0.02411925, 
    0.03399635, 0.05015972, 0.06447805, 0.06572494, 0.06200338, 0.06089724, 
    0.05431969, 0.03883107, 0.01220933, 0.001586517, -7.705486e-06, 
    8.578836e-05, 0.06018038, 0.1065864, 0.03533145, 0.008128121, 0.0014382,
  0.0006521873, 0.02115894, 0.116572, 0.07824649, 0.04875316, 0.0535157, 
    0.05983029, 0.06049089, 0.03670038, 0.02154877, 0.04573707, 0.03258738, 
    0.1023074, 0.06095769, 0.06443753, 0.054719, 0.04355804, 0.02693619, 
    0.01120181, 0.003487856, 0.0007188951, 0.0007287961, 0.0005048173, 
    0.06776385, 0.09387804, 0.07027677, 0.02303933, 0.0008912117, 7.490622e-05,
  0.03946236, 0.1152969, 0.07627885, 0.04193258, 0.01663015, 0.03604113, 
    0.04423604, 0.03760557, 0.09003096, 0.1651277, 0.04701511, 0.0232681, 
    0.05018566, 0.04008717, 0.03024721, 0.0180588, 0.01117932, 0.005633619, 
    0.008602486, 0.004872303, 0.008298685, 0.01281779, 0.07017392, 0.1281957, 
    0.1356023, 0.06327967, 0.05388794, 0.01731568, 0.01599387,
  0.02124017, 0.022907, 0.02246611, 0.2217151, 0.02048189, 0.01378222, 
    0.04602388, 0.03106726, 0.04263301, 0.04798321, 0.08027991, 0.05321111, 
    0.0654982, 0.06966468, 0.06448918, 0.07073972, 0.07614511, 0.09112717, 
    0.1012391, 0.123606, 0.1077391, 0.06373676, 0.09049552, 0.04281245, 
    0.03036617, 0.03377562, 0.03681011, 0.04455283, 0.05976207,
  0.0001411642, 4.671567e-05, 0.001256344, 0.005459404, 0.007853359, 
    0.00663871, 0.07212865, 0.04888124, 0.116957, 0.05737676, 0.08824077, 
    0.05437648, 0.03498302, 0.02484758, 0.02060715, 0.02105582, 0.02412186, 
    0.01837463, 0.01134644, 0.01646594, 0.01594687, 0.07996222, 0.01885279, 
    0.03832275, 0.0238635, 0.03367044, 0.008959052, 0.002841681, 0.002201169,
  0.00203314, 0.006730544, 0.01241438, 0.01351264, 0.04090226, 0.01890088, 
    0.02135725, 0.141589, 0.2472172, 0.1289178, 0.09326678, 0.09229849, 
    0.09626498, 0.07353251, 0.07756255, 0.06847797, 0.05521936, 0.05160225, 
    0.026667, 0.01153954, 0.03356775, 0.04775734, 0.05570826, 0.04925627, 
    0.05916401, 0.05042854, 0.03024027, 0.01456105, 0.009930646,
  0.04536484, 0.04413006, 0.07864397, 0.133995, 0.06024592, 0.02883457, 
    0.136535, 0.02383497, 0.01921245, 0.07123387, 0.101681, 0.09557169, 
    0.1376724, 0.1634381, 0.156623, 0.1742528, 0.1569342, 0.1353305, 
    0.07591823, 0.08942734, 0.1013574, 0.07143234, 0.1192448, 0.1233693, 
    0.1397376, 0.1307415, 0.1062447, 0.07613946, 0.0722395,
  0.1404824, 0.1643518, 0.1567843, 0.1628967, 0.1330765, 0.1393649, 0.13763, 
    0.1805124, 0.1356499, 0.1260684, 0.1402304, 0.1628514, 0.1755743, 
    0.210501, 0.2220656, 0.205879, 0.1996913, 0.2028475, 0.1755704, 0.171226, 
    0.1333507, 0.1257008, 0.1981954, 0.2435707, 0.2085769, 0.1828787, 
    0.1858462, 0.1723144, 0.1548772,
  0.2065565, 0.2197656, 0.2117077, 0.2494059, 0.2656389, 0.2492151, 
    0.2562726, 0.2650818, 0.2536044, 0.2610315, 0.2306623, 0.1852645, 
    0.23832, 0.2486196, 0.2177665, 0.2481599, 0.2462188, 0.3572541, 
    0.2848935, 0.1886813, 0.1704331, 0.2094851, 0.2294579, 0.2713889, 
    0.2490733, 0.281161, 0.2224736, 0.2385526, 0.2266558,
  0.256648, 0.2222259, 0.2806761, 0.2638312, 0.2734321, 0.2639072, 0.2649092, 
    0.3086093, 0.2571507, 0.2409661, 0.2149979, 0.2267486, 0.1998461, 
    0.1990672, 0.228383, 0.1846106, 0.219237, 0.2186577, 0.1891999, 
    0.2197299, 0.2050283, 0.1910431, 0.1996304, 0.198863, 0.1718023, 
    0.3157147, 0.2474039, 0.2268001, 0.2321252,
  0.1808893, 0.2236923, 0.2199062, 0.2094608, 0.2008102, 0.1994333, 0.205965, 
    0.2315964, 0.2176808, 0.2186684, 0.217445, 0.2294847, 0.2409203, 
    0.2413833, 0.253284, 0.2506361, 0.2320934, 0.2116259, 0.2171102, 
    0.2215067, 0.2153356, 0.2393967, 0.2117029, 0.1341172, 0.1497067, 
    0.1345675, 0.1558402, 0.1516102, 0.2156023,
  0.1229036, 0.1203569, 0.1178102, 0.1152635, 0.1127167, 0.11017, 0.1076233, 
    0.1184467, 0.1221792, 0.1259118, 0.1296443, 0.1333768, 0.1371093, 
    0.1408419, 0.140065, 0.144, 0.147935, 0.1518701, 0.1558051, 0.1597401, 
    0.1636751, 0.1585609, 0.15344, 0.1483192, 0.1431984, 0.1380776, 
    0.1329568, 0.127836, 0.124941,
  0.1582586, 0.1100379, 0.07182302, 0.06729865, 0.05827625, 0.06658445, 
    0.05814843, 0.05022167, 0.04899843, 0.06560257, 0.07404587, 0.1047925, 
    0.1479252, 0.1664312, 0.123963, 0.1547715, 0.1837751, 0.2217437, 
    0.2151267, 0.220606, 0.2990754, 0.3674439, 0.270547, 0.2350483, 
    0.2026598, 0.1829491, 0.2086808, 0.2045084, 0.1760838,
  0.2488482, 0.2786006, 0.2691969, 0.2922246, 0.2754223, 0.1989215, 
    0.2384098, 0.2741258, 0.2625286, 0.2800731, 0.2732103, 0.2239791, 
    0.2308771, 0.2742602, 0.2814054, 0.2852932, 0.2656244, 0.2849773, 
    0.3040928, 0.2829838, 0.2939428, 0.3046869, 0.319254, 0.4017979, 
    0.2902928, 0.203298, 0.215852, 0.2494339, 0.2705217,
  0.2800656, 0.3028908, 0.3237209, 0.3308704, 0.3325057, 0.3149028, 
    0.3048288, 0.3048463, 0.3320388, 0.3240405, 0.3222195, 0.3181916, 
    0.2970293, 0.2834347, 0.2767439, 0.2574618, 0.2610778, 0.2736213, 
    0.2913657, 0.3016502, 0.2967295, 0.2778911, 0.2825505, 0.2745467, 
    0.2619778, 0.2453064, 0.2460721, 0.2505175, 0.2695822,
  0.2331698, 0.2234746, 0.2284266, 0.2141531, 0.2023303, 0.2016162, 
    0.1973746, 0.2292547, 0.2225127, 0.2369574, 0.2461718, 0.2185743, 
    0.1962218, 0.177258, 0.1533734, 0.1538613, 0.1708275, 0.1842054, 
    0.1982469, 0.1966842, 0.2095701, 0.2037211, 0.2009399, 0.1665937, 
    0.1156977, 0.1579365, 0.178655, 0.1924129, 0.202466,
  0.1328596, 0.1136158, 0.08548224, 0.1108077, 0.117538, 0.1146398, 
    0.1227003, 0.1229995, 0.1117335, 0.09464478, 0.09146106, 0.08811673, 
    0.09079714, 0.1206899, 0.1470753, 0.1303183, 0.1326746, 0.1225647, 
    0.1278251, 0.1287567, 0.1414178, 0.1320153, 0.119445, 0.1113551, 
    0.06327996, 0.1075727, 0.1252588, 0.1348783, 0.1450692,
  0.02659864, 0.008990904, 0.06574003, 0.04023324, 0.05299778, 0.06955478, 
    0.0434143, 0.02895437, 0.02760881, 0.01858291, 0.01133136, 0.009525893, 
    0.07023254, 0.06144917, 0.08390854, 0.09350978, 0.1027847, 0.1089793, 
    0.1249774, 0.1004801, 0.08691345, 0.05706917, 0.02181456, 0.00322006, 
    0.05075818, 0.08904057, 0.0913216, 0.06245854, 0.0523945,
  0.0009285967, 0.0162324, 0.05931606, 0.02721148, 0.07273962, 0.04540769, 
    0.04584433, 0.03364466, 0.01736351, 0.008273247, 0.01828478, 0.0243051, 
    0.03723186, 0.05321064, 0.06975298, 0.06408879, 0.05939147, 0.06283163, 
    0.06134352, 0.05453102, 0.03339672, 0.005996049, 0.000407058, 
    0.0001001172, 0.06079918, 0.09599628, 0.05045745, 0.02267919, 0.003891088,
  0.000426303, 0.01797472, 0.09618659, 0.09435973, 0.05029162, 0.05416571, 
    0.05933898, 0.06364741, 0.0379871, 0.02232432, 0.04964003, 0.03379329, 
    0.1085024, 0.05958521, 0.05983945, 0.05292206, 0.04662313, 0.03245448, 
    0.01740051, 0.006577918, 0.001172281, 0.0005849635, 0.0003780128, 
    0.06628446, 0.07975031, 0.06915715, 0.03670375, 0.001513178, 0.0001599448,
  0.03140831, 0.1031124, 0.06171973, 0.05722434, 0.0185111, 0.03577555, 
    0.04333689, 0.03592922, 0.09792562, 0.164803, 0.04488209, 0.02131842, 
    0.04634557, 0.03727972, 0.03078349, 0.02254787, 0.01389891, 0.008039184, 
    0.01022568, 0.00675621, 0.009647164, 0.01368951, 0.05795629, 0.1241353, 
    0.126476, 0.0564981, 0.05569679, 0.02227568, 0.01700441,
  0.01708107, 0.01760954, 0.01592794, 0.1718898, 0.01906782, 0.0159409, 
    0.04833882, 0.03084209, 0.04267095, 0.04722555, 0.08506958, 0.05341151, 
    0.06268936, 0.06774023, 0.06303627, 0.0693884, 0.07488149, 0.09322327, 
    0.1082399, 0.1231892, 0.1052378, 0.06483477, 0.1012209, 0.04704358, 
    0.03308723, 0.03224951, 0.03601305, 0.04179274, 0.05201688,
  1.609348e-05, 2.481788e-05, 0.001482665, 0.006062025, 0.003869057, 
    0.005132406, 0.06681605, 0.05235545, 0.1205919, 0.06146776, 0.08587855, 
    0.05717251, 0.03942446, 0.03021083, 0.0268904, 0.02609414, 0.02837859, 
    0.02032567, 0.01112737, 0.01854418, 0.01388587, 0.09396613, 0.02128343, 
    0.03915114, 0.02772621, 0.038945, 0.01414134, 0.001361785, 0.001437142,
  0.002022571, 0.005428543, 0.01951085, 0.01623483, 0.04001793, 0.01746081, 
    0.0138811, 0.1368073, 0.2311913, 0.1276561, 0.09526057, 0.09754746, 
    0.09812132, 0.07647593, 0.08179227, 0.07380461, 0.06199409, 0.0583927, 
    0.03118788, 0.01308185, 0.03056284, 0.04992597, 0.06045769, 0.05246115, 
    0.06160663, 0.05380734, 0.03621585, 0.01815462, 0.008952046,
  0.03830831, 0.04520927, 0.08149758, 0.1440967, 0.05360642, 0.02600043, 
    0.1296599, 0.01810396, 0.01296346, 0.05979297, 0.1020751, 0.1043873, 
    0.1483956, 0.1706937, 0.1622483, 0.1789, 0.1656666, 0.1425511, 
    0.08663955, 0.0960707, 0.09483957, 0.06383649, 0.1227219, 0.1237156, 
    0.1491108, 0.1384701, 0.1134413, 0.08459885, 0.08177552,
  0.1471798, 0.1787992, 0.1647467, 0.1648447, 0.1239071, 0.132652, 0.1315859, 
    0.1858356, 0.1329045, 0.1163683, 0.1350428, 0.1708772, 0.1880253, 
    0.2317333, 0.2339778, 0.2218718, 0.2147675, 0.2143699, 0.1817745, 
    0.1809423, 0.1238426, 0.1158795, 0.1972683, 0.2516908, 0.2115082, 
    0.1979473, 0.1994272, 0.1882965, 0.1599584,
  0.2188027, 0.2282628, 0.216894, 0.2616698, 0.280361, 0.2556334, 0.2586872, 
    0.276606, 0.2545267, 0.2680667, 0.2478284, 0.1949, 0.2426431, 0.2543302, 
    0.2261064, 0.2576156, 0.26637, 0.3675556, 0.2849322, 0.1866327, 
    0.1664515, 0.2020611, 0.2169814, 0.2758865, 0.2414398, 0.2882091, 
    0.2434171, 0.2595045, 0.2494182,
  0.2722999, 0.2408611, 0.2794205, 0.2690529, 0.2839483, 0.2665442, 
    0.2682147, 0.3200208, 0.2657068, 0.2534826, 0.2311293, 0.2371378, 
    0.2000578, 0.2113489, 0.2279838, 0.1874178, 0.2225773, 0.223154, 
    0.1854708, 0.2123846, 0.2049929, 0.1837561, 0.1999008, 0.1885552, 
    0.1728361, 0.3437832, 0.2475068, 0.2336387, 0.2496734,
  0.2002698, 0.2374796, 0.2300314, 0.2149026, 0.2062345, 0.2063146, 
    0.2059507, 0.2357028, 0.2249966, 0.2221844, 0.2231881, 0.2259005, 
    0.236637, 0.2421684, 0.2442977, 0.2436595, 0.2239113, 0.1931777, 
    0.2034015, 0.2221834, 0.2148429, 0.2474316, 0.2170049, 0.1457863, 
    0.1454923, 0.134906, 0.1485363, 0.1560644, 0.2231897,
  0.1592884, 0.15696, 0.1546317, 0.1523034, 0.149975, 0.1476467, 0.1453184, 
    0.1634193, 0.1684697, 0.17352, 0.1785704, 0.1836207, 0.1886711, 
    0.1937214, 0.1906431, 0.1942183, 0.1977934, 0.2013685, 0.2049437, 
    0.2085188, 0.2120939, 0.1996512, 0.193354, 0.1870568, 0.1807597, 
    0.1744625, 0.1681654, 0.1618682, 0.1611511,
  0.1745473, 0.1436609, 0.09600423, 0.07791159, 0.06698003, 0.0784501, 
    0.07517356, 0.07154155, 0.06791876, 0.08245033, 0.09778358, 0.122076, 
    0.1721526, 0.1471344, 0.1262668, 0.1385894, 0.1764195, 0.2003065, 
    0.1985547, 0.2178937, 0.3234025, 0.3835748, 0.2859625, 0.2325438, 
    0.2090085, 0.1872971, 0.2177128, 0.2075171, 0.1864478,
  0.2422268, 0.2636343, 0.2618711, 0.2818075, 0.2830867, 0.2084673, 
    0.2468454, 0.2924793, 0.2838243, 0.2899745, 0.2799742, 0.2260672, 
    0.227115, 0.2715965, 0.2786466, 0.2696564, 0.2583908, 0.2658246, 
    0.2821592, 0.2769542, 0.2766837, 0.288043, 0.2976997, 0.3825823, 
    0.269535, 0.193221, 0.2246723, 0.2562407, 0.2662549,
  0.26857, 0.293292, 0.320765, 0.3218392, 0.3230783, 0.3047361, 0.297282, 
    0.3012243, 0.3202139, 0.3230361, 0.3148643, 0.3049205, 0.2868689, 
    0.2814407, 0.2761144, 0.2570753, 0.260191, 0.2640762, 0.2900568, 
    0.3021799, 0.2969405, 0.2813453, 0.287745, 0.2694307, 0.2536916, 
    0.2291568, 0.236619, 0.2482184, 0.2654656,
  0.2368853, 0.2343863, 0.2355024, 0.2268984, 0.2172538, 0.2096426, 
    0.2105536, 0.2461041, 0.2406291, 0.2529136, 0.2670352, 0.2321381, 
    0.2177495, 0.1911425, 0.1665786, 0.1702499, 0.1863168, 0.2037234, 
    0.2210774, 0.2151628, 0.2253912, 0.2198908, 0.2151364, 0.1745668, 
    0.1085447, 0.1583281, 0.1819763, 0.1965353, 0.2145735,
  0.1487563, 0.1339154, 0.103626, 0.130862, 0.1300705, 0.1291334, 0.1326235, 
    0.1398441, 0.1321685, 0.1118672, 0.1028643, 0.1025179, 0.09412349, 
    0.1292602, 0.1620187, 0.1434229, 0.1446102, 0.1373459, 0.1397843, 
    0.1390528, 0.1541909, 0.1463518, 0.1369195, 0.1223551, 0.05874466, 
    0.117924, 0.1393365, 0.1486886, 0.1584539,
  0.03715778, 0.01295312, 0.0556332, 0.04265743, 0.05847349, 0.07379539, 
    0.05578081, 0.0413694, 0.03857481, 0.02693425, 0.01092544, 0.006335053, 
    0.05421429, 0.07004837, 0.08654325, 0.0970725, 0.1092677, 0.1155225, 
    0.1266228, 0.1036676, 0.09201273, 0.07280247, 0.02854305, 0.003169733, 
    0.04581827, 0.08708299, 0.09681931, 0.07039811, 0.06636871,
  0.001948291, 0.0104917, 0.0559356, 0.0290707, 0.06912952, 0.05031382, 
    0.05177576, 0.04078051, 0.02058085, 0.009695636, 0.01499462, 0.01590472, 
    0.04002313, 0.054868, 0.07172967, 0.06147818, 0.05852255, 0.06238724, 
    0.05886967, 0.05829635, 0.06291153, 0.02674568, 0.0008307098, 
    0.0001559114, 0.06074081, 0.09617712, 0.0547476, 0.04697319, 0.01593896,
  0.0001848602, 0.01477993, 0.08595498, 0.09555639, 0.04936868, 0.05486763, 
    0.05847314, 0.06680325, 0.04009436, 0.02506505, 0.05499641, 0.03775105, 
    0.1113935, 0.05428952, 0.05130286, 0.04519298, 0.04199549, 0.03076858, 
    0.02109868, 0.01390973, 0.002660798, 0.001128596, 0.0006054329, 
    0.06307188, 0.0686569, 0.04708667, 0.04506785, 0.003924785, 0.00117722,
  0.02759217, 0.09786764, 0.05402869, 0.06034761, 0.02308363, 0.03613608, 
    0.0402784, 0.0328214, 0.1029292, 0.1685997, 0.04322766, 0.01932875, 
    0.04007156, 0.03294513, 0.02899368, 0.02327909, 0.0178675, 0.0124567, 
    0.01216928, 0.00922469, 0.01239596, 0.01538593, 0.04588007, 0.1198227, 
    0.1125473, 0.04883669, 0.05314027, 0.02732384, 0.01816684,
  0.01586413, 0.01527594, 0.01300602, 0.1202615, 0.0200892, 0.01890578, 
    0.04891066, 0.02906526, 0.03962095, 0.04568087, 0.08353162, 0.04935601, 
    0.05691976, 0.06145722, 0.05954306, 0.06620312, 0.07312713, 0.09346948, 
    0.1133478, 0.1201052, 0.1016217, 0.06219678, 0.111923, 0.05350745, 
    0.03196977, 0.03223855, 0.03607241, 0.0398108, 0.04540555,
  4.440001e-06, 5.76297e-06, 0.00069695, 0.009053178, 0.001670725, 
    0.004677597, 0.06407192, 0.05265846, 0.1210032, 0.07024235, 0.08232757, 
    0.06319582, 0.04164891, 0.0337431, 0.03466336, 0.03125212, 0.03771298, 
    0.0281682, 0.01434162, 0.02255103, 0.01200692, 0.1092477, 0.02378372, 
    0.0383641, 0.03036925, 0.04186576, 0.01905288, 0.001238107, 0.0007122387,
  0.002165876, 0.009853628, 0.02386152, 0.01460708, 0.03675466, 0.01629598, 
    0.008130182, 0.1146376, 0.2146453, 0.1216128, 0.0998895, 0.1135627, 
    0.1021335, 0.07978708, 0.08666687, 0.08293247, 0.0751886, 0.06579095, 
    0.03481141, 0.01447691, 0.02575135, 0.05166695, 0.05951265, 0.05913785, 
    0.06511477, 0.05894051, 0.04636342, 0.0244452, 0.007878994,
  0.03188505, 0.04673334, 0.08005107, 0.1534182, 0.04856027, 0.02377322, 
    0.1218442, 0.01410573, 0.009839623, 0.05667285, 0.1031482, 0.1232591, 
    0.1650617, 0.1880386, 0.1762126, 0.1914925, 0.1788824, 0.1525068, 
    0.09904122, 0.09770525, 0.08998312, 0.06195775, 0.1242221, 0.1232625, 
    0.1651825, 0.143799, 0.1208321, 0.09502733, 0.08628788,
  0.1492888, 0.1892625, 0.166184, 0.1616809, 0.1046715, 0.1197743, 0.1179495, 
    0.1847355, 0.1263656, 0.1034532, 0.1299415, 0.177883, 0.1967991, 
    0.2532591, 0.2462901, 0.2334015, 0.2225054, 0.2227838, 0.1861217, 
    0.1904246, 0.1196429, 0.1132086, 0.1889132, 0.2657448, 0.2165365, 
    0.2151178, 0.2187984, 0.203383, 0.1684108,
  0.2275323, 0.2272634, 0.2182924, 0.2642955, 0.2730335, 0.2502625, 
    0.2526115, 0.2636983, 0.2523582, 0.2748085, 0.2450067, 0.1944447, 
    0.2469747, 0.2628118, 0.2378537, 0.2474411, 0.2740773, 0.3731481, 
    0.2860736, 0.1802716, 0.1651305, 0.1901881, 0.2141676, 0.2725241, 
    0.2433413, 0.2851465, 0.2614346, 0.2722648, 0.2600818,
  0.2757644, 0.2540613, 0.2879443, 0.2705487, 0.2625317, 0.2610846, 
    0.2602953, 0.322439, 0.2645041, 0.268753, 0.2387688, 0.2277144, 
    0.1954503, 0.2150728, 0.2238013, 0.1719025, 0.207996, 0.2224855, 
    0.1754406, 0.20986, 0.2092621, 0.1870685, 0.2132992, 0.1833016, 
    0.1634972, 0.3643067, 0.2532715, 0.2332083, 0.2541582,
  0.1969577, 0.2139338, 0.2271808, 0.1994081, 0.1966573, 0.200038, 0.2078122, 
    0.2276121, 0.214179, 0.2156238, 0.2112346, 0.2110537, 0.2216849, 
    0.232371, 0.2252338, 0.2326576, 0.2157479, 0.1863118, 0.2036379, 
    0.2285255, 0.216226, 0.2443585, 0.219269, 0.1467572, 0.1398885, 
    0.1392227, 0.1510603, 0.1720609, 0.2320334,
  0.1881205, 0.1859854, 0.1838503, 0.1817152, 0.1795801, 0.177445, 0.1753099, 
    0.1936975, 0.1997289, 0.2057603, 0.2117916, 0.217823, 0.2238544, 
    0.2298858, 0.2306628, 0.2339374, 0.2372121, 0.2404867, 0.2437614, 
    0.2470361, 0.2503107, 0.2387824, 0.2316115, 0.2244406, 0.2172697, 
    0.2100987, 0.2029278, 0.1957569, 0.1898286,
  0.1838825, 0.1716024, 0.1265236, 0.09691143, 0.07912271, 0.09483447, 
    0.09970126, 0.08526592, 0.07972412, 0.09564076, 0.1218032, 0.132286, 
    0.1989971, 0.1278105, 0.130514, 0.1480156, 0.1778155, 0.1877248, 
    0.1883334, 0.208834, 0.3540004, 0.3947461, 0.305628, 0.2361854, 
    0.2212815, 0.1925408, 0.2199064, 0.1979923, 0.1999457,
  0.2537659, 0.2645548, 0.2664459, 0.2585717, 0.2797404, 0.213202, 0.2387745, 
    0.3027802, 0.2947802, 0.2971399, 0.2814426, 0.218187, 0.2206774, 
    0.2801857, 0.3059235, 0.2856842, 0.2767129, 0.2916503, 0.314999, 
    0.3018318, 0.3112095, 0.2990144, 0.3058463, 0.3887413, 0.2653519, 
    0.2226937, 0.2335538, 0.2795268, 0.2824134,
  0.3090092, 0.3134557, 0.3429536, 0.3480793, 0.3367524, 0.3193002, 
    0.3363032, 0.3332425, 0.3539613, 0.3632403, 0.3399687, 0.3225711, 
    0.3113604, 0.3162516, 0.3002351, 0.284799, 0.2872034, 0.2888151, 
    0.323958, 0.3389589, 0.3205378, 0.3130786, 0.316337, 0.2965339, 
    0.2691478, 0.2507848, 0.2585664, 0.2751315, 0.3042178,
  0.267313, 0.2638142, 0.2682553, 0.257659, 0.2478939, 0.2365727, 0.2367151, 
    0.2849376, 0.2652441, 0.2793354, 0.293668, 0.2615402, 0.2409522, 
    0.2187181, 0.1817101, 0.197717, 0.2201402, 0.2477968, 0.2638869, 
    0.2588226, 0.2508173, 0.2419682, 0.2460582, 0.1850538, 0.109766, 
    0.1716613, 0.2101899, 0.2325634, 0.2470832,
  0.1818009, 0.1673415, 0.1392718, 0.1660492, 0.1600222, 0.1650316, 
    0.1554189, 0.1693662, 0.1663738, 0.1430758, 0.1293331, 0.1209109, 
    0.1019912, 0.1448618, 0.1816212, 0.1573895, 0.1678945, 0.1629089, 
    0.1710915, 0.1674923, 0.18016, 0.1753782, 0.1669546, 0.1355018, 
    0.06267755, 0.1416175, 0.1661281, 0.1736347, 0.179399,
  0.06649666, 0.02642644, 0.04923868, 0.06160453, 0.06907295, 0.08790883, 
    0.073702, 0.07129758, 0.05867217, 0.04357582, 0.00920266, 0.005109601, 
    0.04233889, 0.08922759, 0.09767707, 0.1094069, 0.120344, 0.1351608, 
    0.1370908, 0.1098953, 0.1045826, 0.09585851, 0.05119698, 0.003382333, 
    0.04227649, 0.0969074, 0.1071245, 0.08317545, 0.09007732,
  0.01290328, 0.00773846, 0.04451823, 0.03099079, 0.06605631, 0.05403209, 
    0.06431966, 0.06201149, 0.04888769, 0.01729972, 0.01239968, 0.01282537, 
    0.04662691, 0.0575923, 0.07559409, 0.06330448, 0.06239522, 0.06111688, 
    0.05467391, 0.05511965, 0.08093572, 0.07571069, 0.009339226, 
    0.0002779556, 0.06487305, 0.09682193, 0.05277182, 0.07631117, 0.05134542,
  0.001285341, 0.01146631, 0.07602268, 0.08725462, 0.04535788, 0.05250327, 
    0.05715956, 0.0655765, 0.04052162, 0.02790339, 0.05797319, 0.04073672, 
    0.1151721, 0.04872054, 0.04319211, 0.03845807, 0.03614881, 0.02729032, 
    0.02203844, 0.02334454, 0.009042282, 0.003310406, 0.002870104, 
    0.05904385, 0.05948521, 0.0336681, 0.05025291, 0.01364872, 0.00511829,
  0.02652583, 0.09634478, 0.04885753, 0.05433548, 0.0262975, 0.03622216, 
    0.0356965, 0.0297799, 0.1028597, 0.1764725, 0.03977573, 0.01775539, 
    0.03530261, 0.02847444, 0.02730386, 0.02181171, 0.01956915, 0.01547817, 
    0.01668156, 0.0126956, 0.01448275, 0.01655797, 0.03442563, 0.1129928, 
    0.1018573, 0.04128558, 0.04826054, 0.02803457, 0.01775698,
  0.01653511, 0.01413011, 0.0113522, 0.08713458, 0.02852839, 0.02217203, 
    0.04762055, 0.02761376, 0.03844561, 0.04278712, 0.08219103, 0.04292782, 
    0.04913487, 0.05381502, 0.05396374, 0.05970322, 0.07160925, 0.09362547, 
    0.1139979, 0.1112474, 0.09287024, 0.05652424, 0.1172002, 0.05891304, 
    0.03110736, 0.03423256, 0.03774009, 0.03720793, 0.04031193,
  1.136587e-06, 1.052003e-06, 0.0001256689, 0.01466457, 0.0009828481, 
    0.01358077, 0.06307722, 0.04871394, 0.1247676, 0.08943971, 0.08708397, 
    0.06926891, 0.04333102, 0.03853961, 0.04198505, 0.03983192, 0.04606298, 
    0.04922183, 0.02319184, 0.02670979, 0.0117034, 0.1268455, 0.02821138, 
    0.03711597, 0.03392096, 0.04479243, 0.03105222, 0.001654116, 0.0001948628,
  0.0009863345, 0.01258191, 0.0295474, 0.01493203, 0.03431943, 0.01373506, 
    0.005975058, 0.09320126, 0.2075884, 0.1159277, 0.1236409, 0.1466136, 
    0.121268, 0.09988081, 0.1022202, 0.1051761, 0.09476874, 0.08517378, 
    0.05270506, 0.0213015, 0.02619669, 0.06045972, 0.06046829, 0.07549502, 
    0.07334653, 0.06761542, 0.06182095, 0.04183237, 0.00676897,
  0.02785254, 0.04785734, 0.07506504, 0.1643769, 0.04681953, 0.0225021, 
    0.1121011, 0.01053286, 0.008311058, 0.05451279, 0.1077342, 0.1501336, 
    0.1952094, 0.2064756, 0.2054477, 0.2182993, 0.2095959, 0.184356, 
    0.1281424, 0.1043831, 0.08758619, 0.06404855, 0.1339908, 0.1340497, 
    0.1967224, 0.1605067, 0.1464431, 0.1219943, 0.09364163,
  0.1605079, 0.2042768, 0.1880895, 0.1695454, 0.09855362, 0.120082, 
    0.1092903, 0.1925868, 0.1150267, 0.09109132, 0.1281085, 0.1815646, 
    0.2177404, 0.2823857, 0.2768633, 0.2611328, 0.2532612, 0.2569209, 
    0.2123479, 0.2009752, 0.1208124, 0.1239103, 0.1994236, 0.2759545, 
    0.2275039, 0.2462403, 0.2476177, 0.2238, 0.1846574,
  0.2372737, 0.2362831, 0.2284641, 0.2663179, 0.2802297, 0.2357702, 
    0.2541676, 0.2779418, 0.2636883, 0.2890922, 0.2584473, 0.2022658, 
    0.2524158, 0.2808021, 0.2771206, 0.262869, 0.2924405, 0.38103, 0.2964049, 
    0.1771835, 0.1697622, 0.1971881, 0.2233077, 0.2804958, 0.2776171, 
    0.2712727, 0.2943039, 0.2997178, 0.2778717,
  0.3077717, 0.2695436, 0.3045132, 0.2968912, 0.2920953, 0.2695382, 
    0.2732229, 0.3337372, 0.2648501, 0.2850474, 0.2525203, 0.2403607, 
    0.209296, 0.2330638, 0.2405676, 0.1704576, 0.2241922, 0.2266634, 
    0.1734805, 0.2200917, 0.2270264, 0.2045076, 0.2286593, 0.1857988, 
    0.164025, 0.3720753, 0.2574317, 0.2319408, 0.2961431,
  0.2098707, 0.2162113, 0.2364138, 0.2098288, 0.1942254, 0.2199127, 
    0.2262178, 0.2436831, 0.2406892, 0.2327835, 0.2314364, 0.2344507, 
    0.2382286, 0.2453814, 0.2333496, 0.2390999, 0.2332576, 0.2119382, 
    0.2227852, 0.24168, 0.2234941, 0.2489884, 0.2200079, 0.1563578, 
    0.1409526, 0.1511403, 0.157794, 0.1837321, 0.2642746,
  0.2188936, 0.2175433, 0.216193, 0.2148427, 0.2134924, 0.2121422, 0.2107919, 
    0.2230685, 0.2294238, 0.2357791, 0.2421344, 0.2484897, 0.254845, 
    0.2612003, 0.2675368, 0.2698729, 0.2722091, 0.2745453, 0.2768814, 
    0.2792176, 0.2815537, 0.2653515, 0.2580103, 0.2506691, 0.2433279, 
    0.2359868, 0.2286456, 0.2213044, 0.2199738,
  0.1915635, 0.1893245, 0.1619689, 0.1135452, 0.09417121, 0.1159292, 
    0.1238541, 0.1068073, 0.09592978, 0.1158331, 0.1427984, 0.1545729, 
    0.215711, 0.1050515, 0.1353241, 0.1563943, 0.1840485, 0.1911214, 
    0.1905321, 0.2015769, 0.3775863, 0.4135138, 0.3323168, 0.240044, 
    0.2240107, 0.1977589, 0.222226, 0.1915096, 0.2086902,
  0.2800094, 0.2660715, 0.2666487, 0.2331904, 0.2668291, 0.2214857, 
    0.2204683, 0.3159483, 0.3006049, 0.300226, 0.2805867, 0.2093209, 
    0.2190901, 0.2741168, 0.3463112, 0.3182633, 0.3220978, 0.3455936, 
    0.3565062, 0.3466024, 0.3287581, 0.3259227, 0.3202609, 0.4060246, 
    0.2697577, 0.2605179, 0.2730023, 0.3297802, 0.3194512,
  0.3628578, 0.3501007, 0.3862736, 0.3885513, 0.3837804, 0.3733988, 
    0.3826219, 0.38487, 0.412619, 0.4015409, 0.3667434, 0.3613047, 0.3672498, 
    0.3637509, 0.3401467, 0.3286227, 0.3376459, 0.3428486, 0.3700536, 
    0.3715253, 0.3391585, 0.3303317, 0.3522679, 0.3446124, 0.3264713, 
    0.3123179, 0.3054227, 0.3247686, 0.3580553,
  0.3158571, 0.3026802, 0.3086109, 0.2935328, 0.2776393, 0.2649038, 0.270571, 
    0.3141524, 0.2845718, 0.30313, 0.3168547, 0.2982376, 0.2731043, 
    0.2573106, 0.2095484, 0.2405405, 0.2612921, 0.2846669, 0.2974181, 
    0.3032829, 0.2896868, 0.2746935, 0.2823886, 0.1934427, 0.1165582, 
    0.2006305, 0.2598001, 0.2783392, 0.2933656,
  0.227829, 0.2067137, 0.1806279, 0.2006597, 0.2062715, 0.1977371, 0.198698, 
    0.2142336, 0.2044122, 0.1752447, 0.1588797, 0.1372468, 0.1086293, 
    0.167002, 0.2061614, 0.1807156, 0.2025749, 0.210453, 0.2132422, 
    0.2107935, 0.2250207, 0.2134089, 0.2058048, 0.153621, 0.0720195, 
    0.1641544, 0.1893334, 0.1982355, 0.2149467,
  0.1156684, 0.04398577, 0.0427138, 0.0891367, 0.09594212, 0.1182456, 
    0.1097704, 0.1321861, 0.1198151, 0.06890615, 0.006475648, 0.00277589, 
    0.03256915, 0.1058148, 0.1181814, 0.1272001, 0.1372361, 0.1509601, 
    0.1478005, 0.1318685, 0.1271162, 0.1290775, 0.1128697, 0.00423715, 
    0.04634776, 0.1172995, 0.1291608, 0.1086627, 0.1264239,
  0.0708026, 0.005742757, 0.03403034, 0.04356853, 0.0673676, 0.0588048, 
    0.08343662, 0.1023412, 0.09575056, 0.01680234, 0.01078505, 0.009603467, 
    0.07114541, 0.07997893, 0.07939361, 0.06720674, 0.07096977, 0.06173428, 
    0.0561504, 0.05979392, 0.1157248, 0.1707995, 0.05796188, 0.0001741014, 
    0.0682647, 0.1013653, 0.05763216, 0.1081314, 0.1505084,
  0.005485652, 0.01178694, 0.06726623, 0.07672725, 0.0434238, 0.04951784, 
    0.0561043, 0.06148998, 0.04365927, 0.03298879, 0.05911151, 0.04407409, 
    0.1149554, 0.04540051, 0.03929001, 0.03777574, 0.03510899, 0.02849367, 
    0.02532426, 0.0306032, 0.03784108, 0.01795199, 0.008439058, 0.05617142, 
    0.05296219, 0.02707647, 0.06166494, 0.03832796, 0.0231421,
  0.03108671, 0.1008068, 0.04218202, 0.04680493, 0.02999387, 0.03597062, 
    0.03455736, 0.02940256, 0.1014132, 0.1807262, 0.03809743, 0.01877744, 
    0.03288881, 0.02838254, 0.02806682, 0.02224434, 0.01859212, 0.0158088, 
    0.01996268, 0.01931981, 0.019505, 0.01435917, 0.02613396, 0.10715, 
    0.0951019, 0.0369513, 0.04490715, 0.03225933, 0.02314886,
  0.01757115, 0.01345133, 0.008917614, 0.06500382, 0.04068861, 0.02974996, 
    0.04391892, 0.03563625, 0.0434038, 0.04520676, 0.0750434, 0.04081702, 
    0.04320426, 0.04920847, 0.05074031, 0.05530511, 0.06702137, 0.09257637, 
    0.1130921, 0.1023209, 0.08386257, 0.0514852, 0.1218826, 0.06158002, 
    0.03399729, 0.04045279, 0.04234739, 0.03467515, 0.03689307,
  4.800123e-07, 2.443918e-07, 4.773116e-05, 0.01329816, 0.000595048, 
    0.02422707, 0.05731033, 0.05027588, 0.1216328, 0.1155135, 0.107656, 
    0.08580609, 0.05543749, 0.05336368, 0.05901048, 0.0543585, 0.06867653, 
    0.07426994, 0.05213647, 0.04597718, 0.01288041, 0.1455583, 0.04514855, 
    0.04004048, 0.04453188, 0.05919574, 0.06274384, 0.00639211, 7.477948e-05,
  0.001491121, 0.016596, 0.03870323, 0.01686091, 0.03347893, 0.01116985, 
    0.003584184, 0.07958435, 0.207017, 0.1122515, 0.172966, 0.1640675, 
    0.1297746, 0.1135032, 0.1279424, 0.1329415, 0.1261066, 0.1258076, 
    0.09850225, 0.03427938, 0.02739013, 0.07337679, 0.069194, 0.1095281, 
    0.08920906, 0.08783362, 0.08570617, 0.07193667, 0.008225283,
  0.02695712, 0.04225438, 0.07291958, 0.1785243, 0.05133443, 0.02413675, 
    0.1011799, 0.006790806, 0.006997066, 0.04699542, 0.1162471, 0.1785245, 
    0.2304761, 0.2253113, 0.2287519, 0.2457383, 0.2551973, 0.233821, 
    0.1699029, 0.1119956, 0.08307438, 0.06790711, 0.1473583, 0.143994, 
    0.2324366, 0.1883879, 0.1721438, 0.152765, 0.1053943,
  0.1666224, 0.2262431, 0.190863, 0.173051, 0.1050204, 0.1293588, 0.1125897, 
    0.1978438, 0.1082128, 0.08728414, 0.116522, 0.1881059, 0.2508862, 
    0.3011081, 0.3034205, 0.2952599, 0.2933112, 0.2925298, 0.2391942, 
    0.2044276, 0.1135458, 0.1233692, 0.2062395, 0.2898264, 0.2424532, 
    0.2798406, 0.281378, 0.2449259, 0.2021814,
  0.2606002, 0.2380337, 0.2312646, 0.2760836, 0.2920638, 0.2407102, 
    0.2675679, 0.2899021, 0.2700323, 0.2981468, 0.2805047, 0.2174489, 
    0.2540176, 0.3063838, 0.3557208, 0.3004282, 0.3127299, 0.3854032, 
    0.3017534, 0.171199, 0.1760702, 0.2077423, 0.2419818, 0.3022189, 
    0.3364637, 0.2583484, 0.3222353, 0.3279112, 0.2916556,
  0.3463311, 0.2865469, 0.3281752, 0.3352978, 0.3252033, 0.2971807, 
    0.3099402, 0.3387535, 0.2746586, 0.3089044, 0.2777713, 0.2603361, 
    0.226927, 0.2525212, 0.2631432, 0.1857029, 0.2491203, 0.2404451, 
    0.1815627, 0.2444418, 0.2551458, 0.2394796, 0.2567205, 0.2017224, 
    0.1712406, 0.3754661, 0.2619497, 0.2364732, 0.356888,
  0.2454293, 0.2589807, 0.2580653, 0.2212167, 0.2164283, 0.2500065, 
    0.2614703, 0.2661112, 0.2745436, 0.2651874, 0.2678615, 0.2642642, 
    0.2698558, 0.2748055, 0.2741616, 0.2704825, 0.2678153, 0.2521466, 
    0.2515222, 0.2784374, 0.246619, 0.2646583, 0.2275067, 0.1668181, 
    0.1461224, 0.1563091, 0.1573626, 0.2053411, 0.2874013,
  0.245364, 0.2448738, 0.2443836, 0.2438934, 0.2434033, 0.2429131, 0.2424229, 
    0.2515553, 0.2578467, 0.2641381, 0.2704296, 0.276721, 0.2830124, 
    0.2893038, 0.2996378, 0.3009256, 0.3022134, 0.3035012, 0.3047889, 
    0.3060767, 0.3073645, 0.2835552, 0.2764661, 0.2693771, 0.2622881, 
    0.2551991, 0.24811, 0.241021, 0.2457561,
  0.2044701, 0.2034926, 0.1848519, 0.1368512, 0.111652, 0.138272, 0.141056, 
    0.1273739, 0.1049649, 0.1287106, 0.1589695, 0.1756801, 0.2317559, 
    0.08036853, 0.1391366, 0.1522873, 0.1780479, 0.1866828, 0.1884227, 
    0.2077259, 0.404646, 0.4265227, 0.3457986, 0.2355437, 0.2368492, 
    0.2234636, 0.210171, 0.1861045, 0.216824,
  0.2918561, 0.2597938, 0.2652232, 0.2030073, 0.2536041, 0.2376701, 
    0.1845161, 0.3201139, 0.3047346, 0.3072362, 0.2827637, 0.2088554, 
    0.2106044, 0.2626746, 0.3424039, 0.3503323, 0.3501841, 0.3835382, 
    0.3956007, 0.3771201, 0.3656431, 0.3692547, 0.3445458, 0.4265842, 
    0.2752043, 0.2924965, 0.3465265, 0.3620254, 0.3449066,
  0.403802, 0.387748, 0.4150301, 0.41582, 0.4164873, 0.4218709, 0.4089456, 
    0.4326242, 0.4388502, 0.4038593, 0.3835263, 0.3876301, 0.4077933, 
    0.3985287, 0.35499, 0.3584462, 0.3791193, 0.3987383, 0.3976052, 
    0.3582595, 0.3440718, 0.329077, 0.3568423, 0.3612548, 0.3828778, 
    0.3722526, 0.3674151, 0.3860317, 0.3999226,
  0.349718, 0.3378264, 0.3424656, 0.3122138, 0.3112952, 0.2988383, 0.3003012, 
    0.3224318, 0.3064946, 0.3146442, 0.3156992, 0.302512, 0.2760149, 
    0.2740636, 0.2423525, 0.2669128, 0.296649, 0.311464, 0.3160146, 
    0.3242308, 0.3064084, 0.2977165, 0.3031815, 0.2064169, 0.1148613, 
    0.2306037, 0.319397, 0.3286418, 0.3318003,
  0.2558498, 0.2391146, 0.1813777, 0.2226531, 0.2376046, 0.2346752, 0.238322, 
    0.2642745, 0.2636399, 0.2132082, 0.1762783, 0.1403216, 0.1015873, 
    0.1850075, 0.2405828, 0.2151781, 0.2352823, 0.2520224, 0.2416273, 
    0.2322862, 0.2434825, 0.2387272, 0.2233531, 0.1823134, 0.06688823, 
    0.1660228, 0.2029067, 0.2129263, 0.2500321,
  0.1881638, 0.06002465, 0.03844154, 0.1124054, 0.1136688, 0.1393745, 
    0.1637623, 0.1852752, 0.2059004, 0.06447542, 0.006003705, 0.001870334, 
    0.02440495, 0.1026606, 0.1282125, 0.1359835, 0.1504162, 0.1606284, 
    0.1602365, 0.1368719, 0.1365145, 0.159309, 0.1882094, 0.005011967, 
    0.05045364, 0.1308446, 0.136463, 0.1229699, 0.1577433,
  0.2058729, 0.005272284, 0.02675204, 0.04976493, 0.07789325, 0.06650861, 
    0.09205911, 0.1290354, 0.1489047, 0.01730117, 0.00870613, 0.007038618, 
    0.08092742, 0.1046623, 0.09431166, 0.08393732, 0.08574024, 0.07390426, 
    0.06608608, 0.0798298, 0.1244015, 0.2577398, 0.2398489, 0.0005688959, 
    0.06522664, 0.1002079, 0.07024004, 0.1241945, 0.2277829,
  0.030106, 0.0162225, 0.05054431, 0.07126751, 0.04918716, 0.05650723, 
    0.06244759, 0.07092385, 0.06133663, 0.05046561, 0.06189096, 0.05641117, 
    0.1145726, 0.04924449, 0.0462115, 0.04904426, 0.04797899, 0.04818927, 
    0.04862381, 0.06186476, 0.1004278, 0.09943144, 0.0228813, 0.05261043, 
    0.04372223, 0.01893148, 0.08807524, 0.08422047, 0.09759617,
  0.05165604, 0.1004716, 0.0321001, 0.0410438, 0.04078687, 0.05082658, 
    0.04714592, 0.03658663, 0.09710911, 0.1697531, 0.04470069, 0.02406049, 
    0.03881693, 0.0377447, 0.04515311, 0.03831468, 0.02321559, 0.01715947, 
    0.02290959, 0.02699707, 0.03081321, 0.02130496, 0.0190529, 0.09353019, 
    0.07893673, 0.03848969, 0.05134862, 0.04122366, 0.0356331,
  0.01729705, 0.01273416, 0.006194833, 0.0514957, 0.04404004, 0.07561646, 
    0.03682866, 0.06012094, 0.05326174, 0.05616478, 0.07202908, 0.04683682, 
    0.04600494, 0.05402064, 0.05646979, 0.0608627, 0.07014871, 0.097469, 
    0.113404, 0.0965122, 0.08104703, 0.0592837, 0.1261545, 0.06092436, 
    0.04900114, 0.07600742, 0.08872341, 0.03536864, 0.03244154,
  2.884711e-07, -3.161878e-07, 1.445333e-05, 0.008283503, 0.0004267851, 
    0.03254879, 0.04391545, 0.05020975, 0.1136554, 0.1456795, 0.1185552, 
    0.1049322, 0.07248648, 0.06994533, 0.07398739, 0.07546587, 0.0998914, 
    0.1057896, 0.1367404, 0.09388266, 0.01516162, 0.1608628, 0.05923003, 
    0.04353945, 0.06126105, 0.07516089, 0.09805172, 0.01691081, 4.252064e-05,
  0.0008315475, 0.02546669, 0.02924566, 0.0216977, 0.03323052, 0.01076185, 
    0.001336448, 0.07582276, 0.2000652, 0.1064299, 0.1825304, 0.1459149, 
    0.1301657, 0.1114601, 0.1486786, 0.1534688, 0.1585419, 0.1596558, 
    0.1809264, 0.04695435, 0.02775806, 0.08937743, 0.07775792, 0.1138198, 
    0.09573192, 0.09906808, 0.111151, 0.1153968, 0.00835858,
  0.02933272, 0.0406926, 0.07165211, 0.1897217, 0.04742103, 0.02221009, 
    0.09390727, 0.004147215, 0.006538972, 0.04044373, 0.1273065, 0.1575273, 
    0.223405, 0.2183528, 0.2327593, 0.2584502, 0.2872097, 0.278115, 
    0.2199451, 0.1171222, 0.08004177, 0.07736829, 0.1610626, 0.1498602, 
    0.227715, 0.2060905, 0.1950046, 0.2007207, 0.1275811,
  0.1777014, 0.2347095, 0.1928282, 0.1743824, 0.1286232, 0.1351083, 
    0.1211623, 0.1998204, 0.09772256, 0.08760868, 0.1093104, 0.1936648, 
    0.2650001, 0.2954664, 0.3083534, 0.3292949, 0.3326205, 0.3114997, 
    0.2634973, 0.2088575, 0.1076233, 0.1312394, 0.2136203, 0.3033217, 
    0.2513911, 0.3054727, 0.2888751, 0.2560974, 0.2184319,
  0.248393, 0.2227006, 0.2433408, 0.2829799, 0.3078629, 0.2518418, 0.2784393, 
    0.2895996, 0.2710281, 0.3062732, 0.2844304, 0.2220854, 0.2468968, 
    0.3073037, 0.4233936, 0.3267457, 0.3322142, 0.3825008, 0.3095947, 
    0.1600896, 0.1840668, 0.22148, 0.2467424, 0.317333, 0.3984306, 0.221736, 
    0.3197489, 0.329007, 0.2827495,
  0.3567706, 0.2836403, 0.3391548, 0.3427161, 0.355463, 0.3205698, 0.3243914, 
    0.3604879, 0.2909054, 0.3299942, 0.2976534, 0.2830306, 0.2595587, 
    0.2831558, 0.2939424, 0.2271177, 0.2735038, 0.263707, 0.2082551, 0.27827, 
    0.2829268, 0.2697473, 0.2762506, 0.2164926, 0.178477, 0.3777393, 
    0.2635424, 0.2339505, 0.4133464,
  0.2697908, 0.2974986, 0.290304, 0.2585185, 0.2740192, 0.2975229, 0.3214169, 
    0.3148312, 0.3180436, 0.3216175, 0.3215943, 0.3064457, 0.3193218, 
    0.3314969, 0.3202676, 0.3235151, 0.3097085, 0.2844797, 0.2963103, 
    0.314862, 0.282748, 0.2795587, 0.2405212, 0.1947616, 0.1595675, 
    0.1705594, 0.1603929, 0.230965, 0.3078717,
  0.2707674, 0.2704709, 0.2701744, 0.2698779, 0.2695813, 0.2692848, 
    0.2689883, 0.2774458, 0.283434, 0.2894223, 0.2954105, 0.3013988, 
    0.307387, 0.3133753, 0.3260612, 0.3264925, 0.3269238, 0.3273551, 
    0.3277864, 0.3282177, 0.328649, 0.3061133, 0.2999903, 0.2938672, 
    0.2877442, 0.2816212, 0.2754982, 0.2693751, 0.2710046,
  0.2223164, 0.2236928, 0.2063513, 0.1588133, 0.1299264, 0.155223, 0.1579166, 
    0.141381, 0.1182218, 0.145013, 0.1813046, 0.2025587, 0.2452893, 
    0.05634099, 0.1297162, 0.1531553, 0.1723967, 0.1976444, 0.1873246, 
    0.2102793, 0.435769, 0.4492405, 0.3516583, 0.2250276, 0.2361779, 
    0.253368, 0.1978985, 0.1711096, 0.2283431,
  0.2795274, 0.2436963, 0.2629256, 0.1623153, 0.2276707, 0.2424682, 
    0.1402343, 0.3166524, 0.3062871, 0.3088282, 0.2810643, 0.20595, 
    0.1955402, 0.2465711, 0.3375787, 0.383013, 0.3747548, 0.4033352, 
    0.4048931, 0.3825415, 0.3948922, 0.3822406, 0.3675674, 0.4414912, 
    0.274072, 0.3081149, 0.3666669, 0.3701116, 0.3324625,
  0.4124339, 0.3931672, 0.4175847, 0.4031977, 0.4146337, 0.4342283, 
    0.4162854, 0.4360647, 0.4256327, 0.3672325, 0.362038, 0.3892503, 
    0.4344202, 0.4079202, 0.3566448, 0.3757211, 0.4159839, 0.4348046, 
    0.4138826, 0.335831, 0.3264572, 0.3172216, 0.3478335, 0.3653189, 
    0.3972874, 0.4094974, 0.4173501, 0.4209377, 0.4273185,
  0.3705893, 0.3593784, 0.3605696, 0.33658, 0.3364836, 0.3343966, 0.3302411, 
    0.31288, 0.3088364, 0.317808, 0.301714, 0.3066252, 0.2685657, 0.2617625, 
    0.2460103, 0.2708446, 0.3119684, 0.3392054, 0.3169549, 0.3193776, 
    0.2998842, 0.3050566, 0.2936793, 0.2152551, 0.1090675, 0.2355753, 
    0.3383239, 0.3542339, 0.3494191,
  0.2674769, 0.2295108, 0.1473529, 0.2115375, 0.2266741, 0.2140848, 
    0.2373129, 0.2644525, 0.2749413, 0.22393, 0.2006108, 0.1242436, 
    0.07382467, 0.1810497, 0.2710253, 0.2214981, 0.2396161, 0.2633717, 
    0.2326235, 0.2306836, 0.2263735, 0.2309745, 0.2225844, 0.20878, 
    0.05242098, 0.1567658, 0.2056275, 0.2229193, 0.2525842,
  0.2146367, 0.09481819, 0.0331703, 0.1066286, 0.1208163, 0.1417689, 
    0.1570714, 0.1890431, 0.2173649, 0.04292215, 0.009096904, 0.001143878, 
    0.01823946, 0.08588034, 0.1216103, 0.1297643, 0.1362345, 0.161679, 
    0.1515683, 0.1293699, 0.143108, 0.1485659, 0.2419257, 0.008241557, 
    0.04968886, 0.1242197, 0.1249111, 0.1183257, 0.1578578,
  0.3501035, 0.007952333, 0.02080587, 0.06956165, 0.08192464, 0.06320622, 
    0.07631283, 0.09956474, 0.1654633, 0.02446528, 0.006913127, 0.004574486, 
    0.06679215, 0.1147704, 0.1083108, 0.1007093, 0.09525862, 0.08650497, 
    0.0736184, 0.0641688, 0.08677929, 0.1935144, 0.4462873, 0.002031066, 
    0.05863485, 0.09607644, 0.07523672, 0.09263334, 0.1972312,
  0.2062188, 0.03951798, 0.03477023, 0.06115526, 0.0638943, 0.07270693, 
    0.08082188, 0.08341107, 0.090414, 0.07898606, 0.05415297, 0.06777181, 
    0.1193186, 0.07563899, 0.06291668, 0.06743511, 0.06095888, 0.06553211, 
    0.06094301, 0.06957907, 0.14483, 0.3097571, 0.1173656, 0.03648679, 
    0.0289332, 0.01225298, 0.09389312, 0.1239504, 0.2663605,
  0.0978849, 0.08685829, 0.02024479, 0.0411622, 0.09289514, 0.1152266, 
    0.1189102, 0.0861031, 0.07971103, 0.1367078, 0.07365953, 0.08150596, 
    0.08221644, 0.07201441, 0.07238061, 0.06589103, 0.04339621, 0.0351677, 
    0.04465859, 0.04518612, 0.06643637, 0.0497228, 0.02510959, 0.06576844, 
    0.05018518, 0.0634123, 0.06860816, 0.08115665, 0.07356627,
  0.01598224, 0.0107752, 0.003864299, 0.04290915, 0.05474725, 0.1109718, 
    0.04156993, 0.08597091, 0.05343809, 0.09198807, 0.07209592, 0.07745588, 
    0.05412305, 0.05886162, 0.06146505, 0.07031717, 0.08214653, 0.1187904, 
    0.128274, 0.1186738, 0.1041116, 0.07505566, 0.1629216, 0.06670485, 
    0.05692364, 0.08705531, 0.1433136, 0.04811574, 0.02607507,
  2.083186e-07, -1.002595e-06, 8.31681e-05, 0.004363502, 0.0001287345, 
    0.02342588, 0.03407915, 0.0476565, 0.09274521, 0.1563688, 0.1053907, 
    0.09367315, 0.07325361, 0.07205505, 0.06639307, 0.06280743, 0.08793544, 
    0.1112076, 0.216599, 0.1730007, 0.02865531, 0.1715174, 0.0662954, 
    0.03646395, 0.05423852, 0.07649656, 0.1292637, 0.03303836, 1.76275e-05,
  0.0001736089, 0.02249464, 0.01909729, 0.02037747, 0.03140027, 0.009975674, 
    0.0005934297, 0.07852852, 0.1934585, 0.1006233, 0.1585337, 0.1283554, 
    0.1317216, 0.1177872, 0.1472386, 0.1502859, 0.1516728, 0.1737126, 
    0.2557136, 0.07031594, 0.02988685, 0.1014064, 0.07648157, 0.1120199, 
    0.1011083, 0.1247248, 0.1238554, 0.1814255, 0.009175034,
  0.0285743, 0.03910074, 0.06814417, 0.2049205, 0.03426438, 0.02240635, 
    0.09133729, 0.003401189, 0.005123292, 0.0366438, 0.1351239, 0.1142557, 
    0.2062507, 0.2251788, 0.2409984, 0.2712635, 0.30363, 0.2937702, 
    0.2680012, 0.1229864, 0.07624331, 0.08358026, 0.1659181, 0.1481958, 
    0.2053766, 0.2179256, 0.2127725, 0.2386473, 0.1366842,
  0.1923434, 0.2377097, 0.1916371, 0.1901164, 0.1527458, 0.1391578, 
    0.1215275, 0.1985137, 0.08803581, 0.09108399, 0.1005183, 0.1953527, 
    0.2522904, 0.2835552, 0.310365, 0.3418477, 0.3493453, 0.3354745, 
    0.2823567, 0.2184187, 0.1083183, 0.1353806, 0.2092525, 0.3176429, 
    0.2570423, 0.3068644, 0.2953331, 0.2556233, 0.2357081,
  0.2235453, 0.2133185, 0.2621007, 0.3003656, 0.3261697, 0.2465778, 
    0.2958142, 0.2954184, 0.2798916, 0.3068366, 0.2848421, 0.2332908, 
    0.2424985, 0.2891736, 0.4339972, 0.355175, 0.3435951, 0.3749684, 
    0.3139989, 0.1543487, 0.1985462, 0.2289961, 0.2519355, 0.3081414, 
    0.419087, 0.1849298, 0.3036175, 0.3076636, 0.2737481,
  0.3401797, 0.2494226, 0.3250783, 0.3216605, 0.3630641, 0.3403946, 
    0.3385331, 0.3760236, 0.28707, 0.3358157, 0.3178751, 0.3000484, 
    0.2832529, 0.3183974, 0.3287316, 0.2921765, 0.3088883, 0.2828364, 
    0.2331545, 0.3111309, 0.3072382, 0.3105131, 0.2839085, 0.2474138, 
    0.1975272, 0.3763708, 0.269075, 0.2229748, 0.4161159,
  0.3109336, 0.3394124, 0.330062, 0.3063888, 0.3361224, 0.3538779, 0.3759783, 
    0.3825185, 0.374361, 0.3847753, 0.3604482, 0.353148, 0.3627796, 
    0.3883447, 0.372058, 0.3643682, 0.3551804, 0.3375347, 0.3552963, 
    0.3667754, 0.3476071, 0.3001137, 0.2551613, 0.2240529, 0.178043, 
    0.181301, 0.1716077, 0.2569885, 0.3397559,
  0.2942314, 0.2949615, 0.2956915, 0.2964215, 0.2971515, 0.2978816, 
    0.2986116, 0.3002399, 0.3054448, 0.3106498, 0.3158546, 0.3210596, 
    0.3262645, 0.3314694, 0.3457715, 0.345066, 0.3443605, 0.3436549, 
    0.3429494, 0.3422439, 0.3415384, 0.320287, 0.3150576, 0.3098282, 
    0.3045987, 0.2993693, 0.2941399, 0.2889104, 0.2936474,
  0.2380839, 0.2434604, 0.2219701, 0.1796226, 0.1513886, 0.1595509, 
    0.1678693, 0.1532301, 0.1312757, 0.1543815, 0.1965212, 0.2241131, 
    0.2684456, 0.03857536, 0.1297744, 0.1708403, 0.1883305, 0.2003733, 
    0.1829006, 0.2032347, 0.4429813, 0.4579712, 0.3458411, 0.2164816, 
    0.2217719, 0.2581453, 0.1853774, 0.1574376, 0.2312563,
  0.263995, 0.1994852, 0.2449337, 0.1224924, 0.1877949, 0.2273611, 
    0.09707339, 0.2932911, 0.2917323, 0.2927118, 0.2654532, 0.1947303, 
    0.1689357, 0.2130891, 0.3328272, 0.3884322, 0.3797382, 0.4011552, 
    0.4082714, 0.3911363, 0.4059583, 0.3960278, 0.3808543, 0.4487314, 
    0.2721791, 0.3155916, 0.3573599, 0.3634302, 0.3284678,
  0.4151936, 0.3842868, 0.3859163, 0.372671, 0.3849108, 0.4150546, 0.4031827, 
    0.4071231, 0.3899786, 0.3202672, 0.3327554, 0.3657312, 0.4255186, 
    0.4004333, 0.3543691, 0.3854793, 0.4254658, 0.4494741, 0.4036691, 
    0.3098181, 0.2982309, 0.2975637, 0.326563, 0.3434542, 0.3863819, 
    0.4207619, 0.4432368, 0.4324234, 0.4316642,
  0.361729, 0.3547562, 0.3685679, 0.3360476, 0.3397605, 0.3409182, 0.3344263, 
    0.3064124, 0.3047067, 0.3037527, 0.276945, 0.2793886, 0.2371017, 
    0.2361582, 0.2198387, 0.2599029, 0.293652, 0.3275036, 0.3183493, 
    0.3000554, 0.274656, 0.2903392, 0.2787601, 0.2116885, 0.09287674, 
    0.2314335, 0.3467758, 0.3481119, 0.3609836,
  0.2393297, 0.1793612, 0.1070443, 0.1807824, 0.1954822, 0.191105, 0.2228336, 
    0.2296411, 0.2488136, 0.1773746, 0.148868, 0.07796352, 0.05088449, 
    0.145462, 0.2872734, 0.1896353, 0.1963937, 0.2139013, 0.2101319, 
    0.1948519, 0.2110457, 0.2176877, 0.184908, 0.2285187, 0.04329531, 
    0.1463117, 0.1859147, 0.211785, 0.2349801,
  0.1287868, 0.09209992, 0.02748321, 0.07837468, 0.1053182, 0.1086356, 
    0.09268148, 0.1050348, 0.1392423, 0.02326561, 0.009127825, 0.0009408526, 
    0.01515881, 0.05897335, 0.09564183, 0.09445649, 0.1071618, 0.1382692, 
    0.1380624, 0.1016231, 0.1094201, 0.07546216, 0.148121, 0.01441561, 
    0.04573352, 0.1050867, 0.09679582, 0.07108169, 0.09270576,
  0.215511, 0.01460909, 0.01546499, 0.06144324, 0.04233412, 0.03668767, 
    0.03721103, 0.04838596, 0.1010758, 0.02673913, 0.005655364, 0.002949678, 
    0.05185458, 0.06722911, 0.08010432, 0.07849913, 0.07869639, 0.06914563, 
    0.03606103, 0.02356761, 0.02637632, 0.06880761, 0.265937, 0.07166316, 
    0.05224214, 0.08864859, 0.03034595, 0.03292712, 0.09674625,
  0.4022066, 0.1062955, 0.02483856, 0.06002453, 0.05123963, 0.05142712, 
    0.04498426, 0.04721567, 0.04539567, 0.06694099, 0.0367028, 0.03568578, 
    0.09285776, 0.05097784, 0.0340778, 0.02508886, 0.0218272, 0.0214367, 
    0.01647771, 0.01784156, 0.04420213, 0.1682236, 0.3391879, 0.02065319, 
    0.01958733, 0.007851431, 0.02745713, 0.04568174, 0.1807732,
  0.1618856, 0.06225492, 0.01245659, 0.04160012, 0.07896338, 0.05823787, 
    0.06117405, 0.05861048, 0.06123539, 0.0982398, 0.05406937, 0.103531, 
    0.03393661, 0.02721017, 0.02876705, 0.03830779, 0.04583938, 0.04052834, 
    0.04304294, 0.05821206, 0.1329545, 0.228139, 0.0723885, 0.04088625, 
    0.02725269, 0.04392262, 0.04484043, 0.07273306, 0.1599698,
  0.01019608, 0.0088079, 0.002479321, 0.03886272, 0.05307608, 0.03660992, 
    0.03563448, 0.03154058, 0.02097042, 0.04523847, 0.05573225, 0.05775419, 
    0.03743024, 0.04283772, 0.03443082, 0.04290372, 0.05345099, 0.08173769, 
    0.1006544, 0.1113145, 0.083396, 0.06445964, 0.2433129, 0.07697296, 
    0.02389096, 0.03707178, 0.09458381, 0.08943059, 0.01917541,
  1.725809e-07, -3.208807e-06, 0.0002669983, 0.001541129, 0.0002116881, 
    0.0406841, 0.0327768, 0.03356211, 0.07365429, 0.146106, 0.09084372, 
    0.06099915, 0.035143, 0.03401255, 0.02919518, 0.02590538, 0.03639821, 
    0.0622235, 0.19282, 0.2164819, 0.0392584, 0.1573626, 0.01737769, 
    0.01471995, 0.02572202, 0.03378515, 0.09185392, 0.0578335, 7.788482e-06,
  7.965501e-05, 0.01598968, 0.009031425, 0.0150849, 0.02936277, 0.008089115, 
    -0.0003873942, 0.08210867, 0.1846358, 0.09774049, 0.1380437, 0.1187009, 
    0.1322007, 0.1099578, 0.1345479, 0.1348003, 0.1227156, 0.1239906, 
    0.2252863, 0.09982935, 0.02984068, 0.1057126, 0.06539647, 0.1005467, 
    0.09252907, 0.09194121, 0.08261674, 0.125409, 0.009767445,
  0.02568311, 0.02561358, 0.05315025, 0.2185159, 0.02199219, 0.02270633, 
    0.08845297, 0.002783611, 0.00402212, 0.03455038, 0.1397161, 0.09918212, 
    0.2088489, 0.230914, 0.2461986, 0.2712177, 0.3034855, 0.2971522, 
    0.2704735, 0.1276411, 0.07022418, 0.08442396, 0.1554241, 0.1369532, 
    0.1925598, 0.2038984, 0.1931031, 0.2114773, 0.1423252,
  0.1851275, 0.2318313, 0.184479, 0.1999567, 0.1547095, 0.1421825, 0.1117421, 
    0.1919157, 0.08007918, 0.09154071, 0.09235997, 0.1942245, 0.24551, 
    0.2811973, 0.3088813, 0.3451889, 0.3578765, 0.3387501, 0.2833304, 
    0.2274881, 0.1085212, 0.1255607, 0.1873852, 0.3205383, 0.2478904, 
    0.291064, 0.2722845, 0.258862, 0.2355134,
  0.2006851, 0.2221209, 0.2643104, 0.3218713, 0.3431271, 0.2441145, 
    0.3087662, 0.2959254, 0.2776997, 0.2967723, 0.2889452, 0.2512228, 
    0.2407062, 0.2656103, 0.3848317, 0.3645077, 0.3488871, 0.3553165, 
    0.3088358, 0.1564454, 0.2150113, 0.2229519, 0.2364841, 0.2947725, 
    0.4000309, 0.1621263, 0.2759516, 0.26891, 0.2447214,
  0.3017377, 0.2133874, 0.3032091, 0.2779296, 0.3548015, 0.3535513, 
    0.3678391, 0.3739925, 0.2663167, 0.3262224, 0.3346196, 0.3025705, 
    0.2982582, 0.3374023, 0.361181, 0.3378508, 0.3369706, 0.2804755, 
    0.2531708, 0.3269732, 0.3304874, 0.3542159, 0.284085, 0.2705081, 
    0.1946422, 0.371103, 0.2730487, 0.2073261, 0.3962574,
  0.3605247, 0.3610489, 0.3754035, 0.3621134, 0.4160116, 0.4394716, 
    0.4442664, 0.440547, 0.4267348, 0.4431995, 0.4302936, 0.4243951, 
    0.4294646, 0.4554654, 0.4359479, 0.4269703, 0.4131212, 0.3923084, 
    0.4093213, 0.4373228, 0.3958599, 0.3222443, 0.2551487, 0.2643484, 
    0.1950941, 0.1750294, 0.1703591, 0.2720441, 0.3866813,
  0.3005395, 0.300936, 0.3013326, 0.3017291, 0.3021257, 0.3025222, 0.3029188, 
    0.2939391, 0.2990462, 0.3041534, 0.3092605, 0.3143677, 0.3194749, 
    0.324582, 0.3455819, 0.3444043, 0.3432267, 0.342049, 0.3408714, 
    0.3396938, 0.3385161, 0.3276685, 0.3233424, 0.3190163, 0.3146902, 
    0.3103641, 0.306038, 0.3017119, 0.3002222,
  0.2468371, 0.2602445, 0.2221327, 0.1885006, 0.1568855, 0.1519095, 
    0.1664779, 0.1638993, 0.1289627, 0.1526368, 0.1809134, 0.2058068, 
    0.2856954, 0.02319526, 0.1398391, 0.2003705, 0.216911, 0.2051368, 
    0.1693806, 0.1986922, 0.4295063, 0.4569397, 0.3232891, 0.2016396, 
    0.2129914, 0.2522105, 0.1741392, 0.1433273, 0.2343097,
  0.230159, 0.1588135, 0.2152602, 0.08841438, 0.1419966, 0.2015171, 
    0.06630243, 0.2585066, 0.2669862, 0.2648614, 0.2374122, 0.1826963, 
    0.1377537, 0.1817476, 0.319835, 0.382345, 0.3831807, 0.3879775, 
    0.3911307, 0.3889884, 0.4017448, 0.401193, 0.392682, 0.4489603, 
    0.2719389, 0.3334039, 0.3602496, 0.3496027, 0.3198991,
  0.402341, 0.3714807, 0.3421945, 0.3292076, 0.3460633, 0.372577, 0.3795287, 
    0.3612415, 0.3494403, 0.2755102, 0.2935396, 0.3342396, 0.4052649, 
    0.3804495, 0.3420786, 0.3726524, 0.4143156, 0.4391088, 0.3748993, 
    0.2823579, 0.2672003, 0.2670768, 0.294819, 0.3072001, 0.356027, 
    0.4269369, 0.4469877, 0.4300434, 0.4245319,
  0.3403115, 0.3400998, 0.3514009, 0.3205883, 0.3331054, 0.3302339, 0.321233, 
    0.2776321, 0.287818, 0.2812039, 0.2346098, 0.239781, 0.199419, 0.2156707, 
    0.1948567, 0.2417471, 0.2667791, 0.2948209, 0.2861008, 0.2730348, 
    0.2414711, 0.2615436, 0.2483873, 0.19063, 0.08139043, 0.2258577, 
    0.3413791, 0.3318468, 0.3467572,
  0.2055101, 0.1244438, 0.07488813, 0.1499832, 0.1721314, 0.1658994, 
    0.1814054, 0.1919888, 0.1910176, 0.1239708, 0.08975859, 0.04722653, 
    0.03051043, 0.1199216, 0.2758446, 0.1506737, 0.1571971, 0.1632235, 
    0.1734216, 0.1709881, 0.1900515, 0.1858111, 0.1408968, 0.2353806, 
    0.03999723, 0.1263922, 0.1763671, 0.1861689, 0.2114772,
  0.06233081, 0.05821744, 0.02236382, 0.05299294, 0.07952017, 0.06851452, 
    0.05277513, 0.04609026, 0.06800982, 0.01184712, 0.006687758, 
    0.0004962508, 0.01342293, 0.03829556, 0.0702836, 0.07058071, 0.0866401, 
    0.118132, 0.1170717, 0.07604948, 0.06062474, 0.03545083, 0.06297553, 
    0.0286283, 0.03996645, 0.08140701, 0.07293386, 0.03492496, 0.0452718,
  0.09515121, 0.0279947, 0.0121402, 0.01961428, 0.01319633, 0.01418234, 
    0.01498867, 0.02057584, 0.04291463, 0.01819336, 0.004422074, 0.002077143, 
    0.02020649, 0.03672878, 0.04314573, 0.04436227, 0.03444114, 0.02881112, 
    0.01367259, 0.007050545, 0.006558498, 0.02090525, 0.09800657, 0.09731316, 
    0.040879, 0.087396, 0.01097815, 0.008742363, 0.03584071,
  0.2010042, 0.124047, 0.0199171, 0.07007218, 0.01368507, 0.01569127, 
    0.01712251, 0.01724705, 0.01266945, 0.01301065, 0.02092732, 0.01020634, 
    0.06341377, 0.01790088, 0.01316812, 0.008533663, 0.004890147, 
    0.004612389, 0.002717945, 0.003176556, 0.01080203, 0.0523193, 0.2111005, 
    0.01353607, 0.01552738, 0.00627736, 0.003116554, 0.01061527, 0.06312765,
  0.08442768, 0.04847656, 0.009217623, 0.03655489, 0.0307472, 0.01572434, 
    0.01619473, 0.01490776, 0.05353873, 0.06642133, 0.01786038, 0.01913681, 
    0.01605287, 0.009120557, 0.008992374, 0.007163655, 0.01461811, 
    0.01734173, 0.01962601, 0.04050971, 0.08133505, 0.2921064, 0.303637, 
    0.02882217, 0.01697828, 0.01891834, 0.0191324, 0.01912408, 0.07957575,
  0.006443122, 0.008048376, 0.001884524, 0.03816888, 0.0398081, 0.008546873, 
    0.02804647, 0.007509239, 0.006106935, 0.01607047, 0.0305422, 0.01681338, 
    0.01674547, 0.01589206, 0.01307226, 0.02114081, 0.02697272, 0.04429037, 
    0.05610238, 0.06160586, 0.03978493, 0.03254123, 0.2776129, 0.06973354, 
    0.005456034, 0.01312343, 0.03765798, 0.06655359, 0.01577274,
  1.574445e-07, -3.544126e-06, 0.0001643822, 0.0007336029, 0.0002119146, 
    0.04143999, 0.02917461, 0.01888403, 0.06677615, 0.1263006, 0.04671568, 
    0.02655373, 0.01008155, 0.009810955, 0.008231836, 0.005704848, 
    0.01461875, 0.02612529, 0.09477034, 0.187651, 0.05453572, 0.1288421, 
    0.003910964, 0.003737303, 0.006177871, 0.01267987, 0.03756311, 
    0.04522949, 1.719439e-06,
  0.0001760396, 0.01070231, 0.005420534, 0.009675563, 0.02685018, 
    0.006764484, -0.0009036785, 0.08181137, 0.1735183, 0.09015303, 0.116959, 
    0.1082982, 0.1127988, 0.08905812, 0.1012922, 0.1035191, 0.08456254, 
    0.07238144, 0.1275776, 0.1241326, 0.02773835, 0.09981308, 0.05616232, 
    0.06694558, 0.05115185, 0.04418787, 0.03594762, 0.05476939, 0.0115458,
  0.01816797, 0.01574428, 0.03622867, 0.2256292, 0.01455695, 0.02428944, 
    0.0832845, 0.002149113, 0.002957757, 0.03181481, 0.1411363, 0.08859298, 
    0.2101074, 0.2306546, 0.2377371, 0.2555822, 0.2969453, 0.2609144, 
    0.2428472, 0.1268066, 0.06258619, 0.07870089, 0.1378962, 0.1365342, 
    0.1666781, 0.1771742, 0.1524644, 0.1554703, 0.1323482,
  0.1624485, 0.2132493, 0.180492, 0.1991367, 0.1469336, 0.1409925, 
    0.09116878, 0.1799261, 0.06974711, 0.08458452, 0.0852269, 0.1962501, 
    0.2539993, 0.282644, 0.3136308, 0.3385507, 0.3496585, 0.3244115, 
    0.2556058, 0.2354494, 0.099412, 0.1130965, 0.1723218, 0.3214012, 
    0.2250095, 0.2709104, 0.2456134, 0.2362963, 0.216373,
  0.1828327, 0.234538, 0.2530961, 0.3406207, 0.3547032, 0.2418813, 0.3071162, 
    0.2889967, 0.2734231, 0.2903204, 0.2926141, 0.2791951, 0.2404767, 
    0.2424156, 0.334611, 0.3606228, 0.3547271, 0.3307674, 0.3030796, 
    0.1654603, 0.2403543, 0.2061987, 0.226623, 0.2693626, 0.3759679, 
    0.141149, 0.2397129, 0.2271401, 0.2114683,
  0.2688099, 0.1769733, 0.282844, 0.2323739, 0.3331857, 0.3494336, 0.3959624, 
    0.3589561, 0.2437195, 0.3084733, 0.3512783, 0.30524, 0.2974361, 
    0.3518693, 0.3651718, 0.3427974, 0.3498571, 0.2728676, 0.2675134, 
    0.3298571, 0.3357969, 0.3792737, 0.2930551, 0.2887254, 0.2118638, 
    0.3554645, 0.269823, 0.1843742, 0.3570621,
  0.3945556, 0.3733885, 0.3850529, 0.3896149, 0.4403673, 0.4779342, 
    0.4793506, 0.4669224, 0.4576146, 0.4856269, 0.4745748, 0.4725165, 
    0.4771252, 0.494507, 0.4828077, 0.4828792, 0.458036, 0.4459782, 
    0.4631395, 0.4881979, 0.4364668, 0.326145, 0.2647879, 0.3021259, 
    0.2023577, 0.1761683, 0.166664, 0.2908095, 0.4226764,
  0.2486719, 0.2486272, 0.2485824, 0.2485377, 0.248493, 0.2484483, 0.2484035, 
    0.2384836, 0.2452942, 0.2521048, 0.2589154, 0.265726, 0.2725366, 
    0.2793472, 0.3062149, 0.3047838, 0.3033528, 0.3019217, 0.3004906, 
    0.2990595, 0.2976285, 0.3008419, 0.2955071, 0.2901723, 0.2848375, 
    0.2795027, 0.2741679, 0.2688331, 0.2487077,
  0.2436712, 0.2491352, 0.1979369, 0.1737797, 0.1503701, 0.1299326, 
    0.1480257, 0.1607638, 0.118162, 0.1188555, 0.1301076, 0.1616783, 
    0.2773692, 0.01321188, 0.1538164, 0.2235274, 0.2636228, 0.2179618, 
    0.1592782, 0.1994513, 0.415317, 0.4535168, 0.2862838, 0.1755915, 
    0.2055138, 0.2524708, 0.1671568, 0.126762, 0.2194638,
  0.1981211, 0.1220119, 0.1735428, 0.05982576, 0.1021433, 0.1746128, 
    0.04560418, 0.2147232, 0.2369607, 0.2297467, 0.2047907, 0.1747606, 
    0.1100118, 0.1509898, 0.3070597, 0.3724971, 0.3739641, 0.3665571, 
    0.3574128, 0.3730259, 0.3790403, 0.3887465, 0.3802135, 0.4362061, 
    0.264904, 0.3568336, 0.3716955, 0.3385746, 0.297798,
  0.3721831, 0.3369347, 0.2896109, 0.2718996, 0.2918294, 0.3161913, 
    0.3431748, 0.3090298, 0.2973291, 0.2342786, 0.2503842, 0.2946799, 
    0.375637, 0.3471636, 0.3016036, 0.3456824, 0.3821296, 0.4103521, 
    0.3343411, 0.2421155, 0.2314722, 0.2295014, 0.2509436, 0.2620242, 
    0.3222263, 0.4202612, 0.4317138, 0.4040268, 0.4000657,
  0.3011231, 0.3054527, 0.3117851, 0.2901265, 0.3155341, 0.3067831, 
    0.2933948, 0.2361788, 0.2511772, 0.2430295, 0.1881793, 0.1933466, 
    0.1583104, 0.1819633, 0.1755496, 0.2120676, 0.2196947, 0.2465395, 
    0.2393557, 0.2337412, 0.2049727, 0.2220595, 0.2057521, 0.1594402, 
    0.07281882, 0.2089295, 0.3160063, 0.3064165, 0.3233097,
  0.1617957, 0.07981318, 0.04915956, 0.1197736, 0.1416045, 0.1322634, 
    0.1381293, 0.1514019, 0.1391973, 0.08083518, 0.05501059, 0.02668589, 
    0.02145642, 0.09464241, 0.2471647, 0.1155698, 0.1235851, 0.1326627, 
    0.1389784, 0.1473076, 0.1576117, 0.1460655, 0.1016794, 0.2318918, 
    0.03463022, 0.1004042, 0.1512796, 0.1525553, 0.1704136,
  0.02673628, 0.02631572, 0.01875849, 0.03348783, 0.04995793, 0.04180618, 
    0.03048096, 0.02211514, 0.03405679, 0.008837383, 0.004250765, 
    0.0002751109, 0.01255576, 0.02416011, 0.04939025, 0.04739508, 0.06618125, 
    0.08957149, 0.09042692, 0.04918943, 0.03154776, 0.01696816, 0.02693263, 
    0.02902652, 0.03351728, 0.055308, 0.04775573, 0.01796616, 0.02323355,
  0.04008934, 0.03569429, 0.008043364, 0.006049315, 0.00267951, 0.004721831, 
    0.005195417, 0.01025063, 0.01879434, 0.009721047, 0.003401896, 
    0.001708869, 0.007715276, 0.01861843, 0.0208263, 0.01971433, 0.01265947, 
    0.01034431, 0.00591038, 0.003677028, 0.002461295, 0.007918956, 
    0.03889248, 0.05008002, 0.03023397, 0.08531011, 0.004651838, 0.003151297, 
    0.0139241,
  0.08538222, 0.06427954, 0.01757376, 0.07091887, 0.004430392, 0.004471034, 
    0.005908977, 0.006410017, 0.003515167, 0.002350239, 0.01228278, 
    0.003308119, 0.03676786, 0.004778015, 0.004860546, 0.00362035, 
    0.001559129, 0.001684941, 0.0009925709, 0.001186477, 0.004074672, 
    0.01958782, 0.0870617, 0.01185669, 0.01402172, 0.005583697, 0.0004827388, 
    0.003848051, 0.02355551,
  0.02627361, 0.04520824, 0.00831717, 0.02944974, 0.008015078, 0.006341706, 
    0.007811703, 0.005324274, 0.0486584, 0.05230755, 0.004816683, 
    0.005085999, 0.008254075, 0.004284928, 0.004181132, 0.001756305, 
    0.002874963, 0.002825153, 0.003743648, 0.007071364, 0.02100584, 
    0.1104811, 0.1717184, 0.02509201, 0.01326384, 0.01026901, 0.009403284, 
    0.003771009, 0.02061217,
  0.004259884, 0.007705347, 0.001220895, 0.03928975, 0.02647717, 0.002759182, 
    0.02202583, 0.002569061, 0.002183027, 0.005248037, 0.01347628, 
    0.005563135, 0.006550478, 0.005894183, 0.004281331, 0.00856403, 
    0.01227224, 0.02099225, 0.02736629, 0.02505909, 0.01862656, 0.01169063, 
    0.2471116, 0.05609281, 0.001716312, 0.004695119, 0.01298394, 0.02450847, 
    0.01442147,
  1.495912e-07, -2.667658e-06, 4.293413e-05, 0.0004710454, 0.0001448136, 
    0.02072718, 0.02117254, 0.006799829, 0.06341566, 0.0725498, 0.0190852, 
    0.01071221, 0.002964396, 0.003419073, 0.002237361, 0.001765896, 
    0.006988853, 0.01050502, 0.0423512, 0.1058085, 0.02118219, 0.1001723, 
    0.001333841, 0.0001879769, 0.001997181, 0.004923497, 0.01482867, 
    0.02301467, -7.620112e-07,
  7.911985e-05, 0.007010645, 0.003383916, 0.006611331, 0.02380071, 
    0.005137995, -0.0009813261, 0.07756401, 0.1617294, 0.07881498, 
    0.09908194, 0.08444732, 0.08877659, 0.05974041, 0.06622873, 0.07312677, 
    0.05101583, 0.04086449, 0.06418675, 0.1148516, 0.02418316, 0.08715656, 
    0.04698814, 0.04370649, 0.03046553, 0.02492577, 0.01407935, 0.02298506, 
    0.01236779,
  0.01337012, 0.01011075, 0.02366003, 0.2228775, 0.007703516, 0.02068053, 
    0.07642103, 0.001566565, 0.002835826, 0.0257586, 0.1402125, 0.08100155, 
    0.1968536, 0.2175495, 0.2182568, 0.2178479, 0.2523689, 0.2025672, 
    0.1721726, 0.1198556, 0.05513956, 0.07053072, 0.1195042, 0.1301169, 
    0.1219322, 0.1373362, 0.1075456, 0.1006149, 0.1076874,
  0.1288127, 0.1925315, 0.1636714, 0.1855257, 0.1383936, 0.1270216, 
    0.06773768, 0.1604409, 0.06034032, 0.07562859, 0.07771219, 0.1956868, 
    0.2691547, 0.2733111, 0.2967416, 0.3071204, 0.3173273, 0.2879786, 
    0.219973, 0.2333868, 0.08471803, 0.0932563, 0.1515851, 0.3131694, 
    0.1949068, 0.2506366, 0.2161773, 0.1967845, 0.1856456,
  0.1508235, 0.238134, 0.2413478, 0.3348954, 0.3474835, 0.233084, 0.289777, 
    0.2712711, 0.2670004, 0.2763168, 0.2817424, 0.2973929, 0.2312977, 
    0.2210014, 0.2997089, 0.3555389, 0.3516803, 0.2992591, 0.2836244, 
    0.1658438, 0.2548587, 0.185339, 0.2199852, 0.25029, 0.3409892, 0.1237032, 
    0.2025875, 0.1865557, 0.1822545,
  0.2442777, 0.1457565, 0.261995, 0.1847807, 0.3064307, 0.3394521, 0.403926, 
    0.3257158, 0.2254096, 0.3009872, 0.3564973, 0.3065599, 0.3135535, 
    0.3607259, 0.3640731, 0.3439927, 0.3513938, 0.2710225, 0.275335, 
    0.3142297, 0.3355791, 0.4010433, 0.3005241, 0.3076023, 0.2287719, 
    0.3179076, 0.2638074, 0.1575074, 0.3235175,
  0.4282869, 0.3503946, 0.3965591, 0.4023604, 0.4241801, 0.4905741, 
    0.5056569, 0.4951308, 0.4839295, 0.5166374, 0.5033448, 0.5045097, 
    0.516424, 0.5168148, 0.5121821, 0.5179527, 0.4959263, 0.4929237, 
    0.5056118, 0.5052397, 0.4592603, 0.3076037, 0.2717094, 0.3287369, 
    0.1918607, 0.1725745, 0.1516399, 0.3045987, 0.45051,
  0.1996761, 0.2001206, 0.2005652, 0.2010097, 0.2014543, 0.2018988, 
    0.2023433, 0.1843715, 0.1909343, 0.1974972, 0.2040601, 0.210623, 
    0.2171858, 0.2237487, 0.2596587, 0.2582262, 0.2567936, 0.2553611, 
    0.2539285, 0.2524959, 0.2510634, 0.2473005, 0.2417257, 0.2361508, 
    0.2305759, 0.2250011, 0.2194262, 0.2138514, 0.1993205,
  0.2275716, 0.2113436, 0.1511225, 0.1431862, 0.1358351, 0.1012134, 0.117069, 
    0.1426727, 0.08707375, 0.07980116, 0.07889647, 0.1273232, 0.2413951, 
    0.00757651, 0.1867785, 0.2801638, 0.3083942, 0.2352346, 0.1409948, 
    0.2073843, 0.4005377, 0.4564448, 0.2355257, 0.1423387, 0.2053297, 
    0.279386, 0.1635607, 0.1077631, 0.1971358,
  0.1758677, 0.09493413, 0.1357162, 0.04058374, 0.07467327, 0.1479883, 
    0.03401015, 0.1665573, 0.2036327, 0.1880387, 0.1708031, 0.1645633, 
    0.08622648, 0.1219815, 0.29332, 0.3427148, 0.3357378, 0.3260207, 
    0.3085922, 0.3327307, 0.3405496, 0.3597035, 0.3580177, 0.4035849, 
    0.2439571, 0.3591576, 0.3587435, 0.3158763, 0.2706598,
  0.3205734, 0.2840433, 0.2308852, 0.2108152, 0.2281095, 0.2475609, 
    0.2883168, 0.2474728, 0.237973, 0.1892453, 0.205475, 0.2470236, 
    0.3248949, 0.2939285, 0.2451606, 0.2906621, 0.3271528, 0.3549708, 
    0.2818685, 0.1982475, 0.1905238, 0.1815973, 0.1981701, 0.2051516, 
    0.2847638, 0.3858056, 0.3896205, 0.3527846, 0.3427598,
  0.2522746, 0.2488243, 0.2537265, 0.2432895, 0.2702327, 0.2569858, 
    0.2473436, 0.187849, 0.2011269, 0.1894878, 0.1384666, 0.1393768, 
    0.1135031, 0.1365935, 0.1522373, 0.1709075, 0.1686182, 0.1896158, 
    0.1828008, 0.1815592, 0.1579303, 0.1712904, 0.1563071, 0.1294258, 
    0.06328995, 0.1791994, 0.2703949, 0.2626015, 0.2795872,
  0.1187713, 0.04916594, 0.03271341, 0.09123158, 0.1042013, 0.09412066, 
    0.09848671, 0.1126589, 0.09781751, 0.05228617, 0.03515706, 0.01514292, 
    0.01512113, 0.06917138, 0.209643, 0.08509856, 0.09395304, 0.1069695, 
    0.1114572, 0.118017, 0.1219618, 0.1075779, 0.06826823, 0.2175053, 
    0.02966193, 0.07628527, 0.1136832, 0.1122598, 0.1295612,
  0.01419805, 0.01347165, 0.01500856, 0.01889622, 0.02612836, 0.02461388, 
    0.01706915, 0.0130882, 0.01932573, 0.005622793, 0.00231705, 0.000124933, 
    0.01009916, 0.01337457, 0.0319497, 0.03027228, 0.04518194, 0.06476423, 
    0.06335389, 0.02812077, 0.01660296, 0.008783105, 0.01398452, 0.01964678, 
    0.02729132, 0.03235463, 0.02978579, 0.009371711, 0.01297566,
  0.02121463, 0.03176809, 0.004694397, 0.002817693, -0.000275962, 
    0.001838524, 0.001715709, 0.004655689, 0.009500006, 0.004163655, 
    0.002341821, 0.001046636, 0.003483383, 0.008157838, 0.009361505, 
    0.007980642, 0.00487633, 0.004238117, 0.00285231, 0.001944336, 
    0.001132053, 0.004083183, 0.019935, 0.02819221, 0.02260036, 0.07807405, 
    0.002102069, 0.001498309, 0.006724451,
  0.04440907, 0.03075678, 0.01701222, 0.05745476, 0.00182688, 0.00163601, 
    0.002349881, 0.002355424, 0.001453374, 0.000701769, 0.007472588, 
    0.001559297, 0.01821936, 0.001548093, 0.002422831, 0.001723628, 
    0.0006646506, 0.0008236066, 0.0004713862, 0.0006496481, 0.002188402, 
    0.01002377, 0.04630824, 0.01149912, 0.01439898, 0.005264014, 
    1.285612e-05, 0.00200275, 0.01184186,
  0.01195684, 0.04593255, 0.009634841, 0.02288495, 0.003163347, 0.003178311, 
    0.004195188, 0.002633776, 0.04158065, 0.05230004, 0.002118528, 
    0.002470007, 0.004551178, 0.002389651, 0.002705169, 0.0007166376, 
    0.001143404, 0.000862777, 0.001472617, 0.002271326, 0.006250774, 
    0.04437028, 0.08107192, 0.02537045, 0.01299315, 0.005265361, 0.005356983, 
    0.001622325, 0.009259533,
  0.00327145, 0.00679844, 0.0005643658, 0.03877281, 0.01652126, 0.001427798, 
    0.01413849, 0.001308119, 0.0008481464, 0.002074405, 0.005671861, 
    0.002337891, 0.002617231, 0.002365062, 0.001504538, 0.003992485, 
    0.005471353, 0.01134355, 0.01316035, 0.0106847, 0.00872509, 0.004862723, 
    0.1909495, 0.04653423, 0.0007142246, 0.002157606, 0.005993432, 
    0.01140548, 0.0118757,
  1.431012e-07, -1.160204e-06, 1.583121e-05, 0.0002728143, 0.0001238634, 
    0.01022645, 0.01176634, 0.001904889, 0.05722306, 0.03534762, 0.008389299, 
    0.004820507, 0.001301687, 0.001452752, 0.0008943718, 0.0008293558, 
    0.003446379, 0.004587685, 0.02206371, 0.05979472, 0.01263785, 0.07738214, 
    0.0006748162, -0.0005628631, 0.0009736198, 0.00235379, 0.007370179, 
    0.01254218, -7.216061e-07,
  2.6966e-05, 0.005245565, 0.002304755, 0.004347233, 0.02035673, 0.004315396, 
    -0.0008483586, 0.0713772, 0.1475499, 0.05940879, 0.08224243, 0.05924921, 
    0.06005245, 0.03580144, 0.0406114, 0.0438812, 0.03127376, 0.02380423, 
    0.03559924, 0.08264321, 0.0203324, 0.07383273, 0.03802947, 0.0243839, 
    0.01924706, 0.01310355, 0.007246247, 0.01160657, 0.01080719,
  0.009553264, 0.006127711, 0.01569421, 0.2109208, 0.006252736, 0.01591693, 
    0.0682793, 0.001193593, 0.002073712, 0.02127289, 0.132231, 0.08291657, 
    0.1765506, 0.1856639, 0.1816428, 0.1739995, 0.19239, 0.1519161, 
    0.1180011, 0.1107756, 0.04755814, 0.06006572, 0.09813199, 0.1140373, 
    0.0827447, 0.09120324, 0.06725194, 0.0610305, 0.08225688,
  0.09711766, 0.1673791, 0.1334827, 0.1628484, 0.1175833, 0.101366, 
    0.05043951, 0.1384102, 0.05253575, 0.06946236, 0.07023051, 0.188134, 
    0.2637905, 0.2437787, 0.2574048, 0.2625241, 0.2700949, 0.2382409, 
    0.1790016, 0.2221261, 0.06912284, 0.06834929, 0.1258208, 0.2938666, 
    0.1659549, 0.2379753, 0.1814829, 0.1550942, 0.1462991,
  0.118731, 0.2313662, 0.2129373, 0.3063881, 0.320591, 0.2120446, 0.255679, 
    0.2402155, 0.2475868, 0.25, 0.2651536, 0.2975973, 0.2209884, 0.2027946, 
    0.2678288, 0.3241187, 0.3456595, 0.260826, 0.244566, 0.1629012, 
    0.2544791, 0.165182, 0.2049589, 0.2337983, 0.3037367, 0.1062281, 
    0.1691395, 0.1481305, 0.1470454,
  0.2164697, 0.118547, 0.243004, 0.1472273, 0.2743219, 0.3191158, 0.3845164, 
    0.2902131, 0.2076596, 0.2936802, 0.3718169, 0.2966312, 0.3579263, 
    0.3444693, 0.3461119, 0.3415918, 0.3188256, 0.2565705, 0.2722978, 
    0.2815852, 0.3291954, 0.4259869, 0.3099601, 0.3219768, 0.2396459, 
    0.272131, 0.262933, 0.1366195, 0.290656,
  0.4505492, 0.3238301, 0.4049685, 0.4129943, 0.4239761, 0.4963765, 
    0.5255043, 0.5052173, 0.4974551, 0.5290481, 0.5147371, 0.5137172, 
    0.5180787, 0.5237542, 0.5128982, 0.5260882, 0.5123641, 0.5108131, 
    0.4988136, 0.4987404, 0.4738215, 0.2772067, 0.2686201, 0.3488634, 
    0.1664879, 0.1591474, 0.1343011, 0.2833777, 0.4460146,
  0.1482668, 0.1485025, 0.1487381, 0.1489738, 0.1492095, 0.1494451, 
    0.1496808, 0.1258224, 0.1316411, 0.1374599, 0.1432786, 0.1490974, 
    0.1549162, 0.1607349, 0.2071489, 0.2062897, 0.2054305, 0.2045713, 
    0.2037122, 0.202853, 0.2019938, 0.1901522, 0.1849569, 0.1797617, 
    0.1745664, 0.1693711, 0.1641759, 0.1589806, 0.1480782,
  0.2140481, 0.168981, 0.1070603, 0.1099649, 0.110914, 0.0742327, 0.08724525, 
    0.09814319, 0.06715301, 0.06016264, 0.05464011, 0.08679695, 0.1747395, 
    0.004566222, 0.2212127, 0.3142534, 0.3042207, 0.2357479, 0.1220571, 
    0.2172807, 0.3905941, 0.4651545, 0.1947279, 0.1113111, 0.2041004, 
    0.3117866, 0.1608135, 0.09092642, 0.1821561,
  0.1516932, 0.07458551, 0.1076321, 0.02930572, 0.05692617, 0.1244653, 
    0.02742876, 0.1210945, 0.1660099, 0.1504716, 0.1439588, 0.15089, 
    0.06762179, 0.1005585, 0.2683601, 0.2976174, 0.2852747, 0.2691678, 
    0.2532178, 0.2801858, 0.2851573, 0.3128525, 0.3181577, 0.3579055, 
    0.2241841, 0.3345388, 0.3183245, 0.2708036, 0.2352226,
  0.2531022, 0.2198714, 0.1743874, 0.1561422, 0.1689694, 0.1853732, 
    0.2277196, 0.1925212, 0.1844215, 0.1433661, 0.1575316, 0.1930538, 
    0.2602907, 0.2299567, 0.1823201, 0.2228807, 0.2595322, 0.2889903, 
    0.2262853, 0.1543889, 0.1452084, 0.1290908, 0.1425579, 0.1466226, 
    0.2327087, 0.3260583, 0.3248729, 0.2877933, 0.2716697,
  0.2000725, 0.1928613, 0.196896, 0.1926346, 0.2190201, 0.2052175, 0.1974123, 
    0.1412435, 0.150052, 0.1364882, 0.09247972, 0.08974367, 0.07363392, 
    0.09178862, 0.1201725, 0.1230566, 0.1182379, 0.1322135, 0.1280774, 
    0.1281221, 0.1106881, 0.1193972, 0.1072586, 0.1061844, 0.04917886, 
    0.1399478, 0.2160436, 0.2101362, 0.2282439,
  0.08067314, 0.02948632, 0.02222136, 0.06190272, 0.0676725, 0.06022428, 
    0.06501383, 0.07740864, 0.06278574, 0.03178964, 0.0216525, 0.009069319, 
    0.01046787, 0.04624842, 0.1745027, 0.05494476, 0.06228475, 0.07778689, 
    0.08096463, 0.08346613, 0.08532882, 0.07274824, 0.04055416, 0.1992732, 
    0.02399332, 0.05286532, 0.07761879, 0.07279383, 0.08817832,
  0.008924232, 0.008071755, 0.0110396, 0.00921235, 0.01323399, 0.01291896, 
    0.00970142, 0.008409021, 0.01201581, 0.003864448, 0.001470087, 
    0.0001057939, 0.008124731, 0.006966269, 0.0189089, 0.01813109, 
    0.02667358, 0.0423659, 0.03720641, 0.01535303, 0.008081258, 0.004860141, 
    0.008811681, 0.01286986, 0.02167306, 0.01656509, 0.01678059, 0.004553743, 
    0.007154691,
  0.0135759, 0.02398271, 0.002391333, 0.001684397, -0.001042068, 
    0.0008024295, 0.0007760496, 0.002141953, 0.005472868, 0.00228858, 
    0.001474201, 0.0004882454, 0.001809644, 0.003895039, 0.004004832, 
    0.003264562, 0.00220721, 0.001887089, 0.001281539, 0.0009889191, 
    0.000663376, 0.002572893, 0.01264151, 0.01927911, 0.01621902, 0.06590477, 
    0.001022722, 0.0009120646, 0.004064183,
  0.02810115, 0.01593314, 0.01564154, 0.04374097, 0.0008914773, 0.0007359043, 
    0.001025197, 0.0009555263, 0.0007692224, 0.0005278336, 0.004312572, 
    0.0007341144, 0.007963718, 0.0005998609, 0.001106202, 0.0007794473, 
    0.0003110302, 0.0004365424, 0.0002821638, 0.0004283559, 0.001416113, 
    0.006334787, 0.02966252, 0.01009205, 0.01378049, 0.00446227, 
    4.494741e-06, 0.001275098, 0.007421277,
  0.006889558, 0.04102528, 0.008476936, 0.01738128, 0.001649008, 0.001634242, 
    0.002182747, 0.001362438, 0.03462653, 0.05370984, 0.001075521, 
    0.001455772, 0.002091941, 0.001167452, 0.001496396, 0.0004099616, 
    0.0005839647, 0.0004958012, 0.0008034937, 0.001267681, 0.003193697, 
    0.02446016, 0.04806699, 0.02346029, 0.01279172, 0.002474506, 0.002589384, 
    0.0009028561, 0.005183616,
  0.002037402, 0.004629675, 0.0002189811, 0.03518024, 0.009416116, 
    0.0009379372, 0.007543096, 0.0007797895, 0.0003974485, 0.0009771284, 
    0.002403264, 0.001136995, 0.001078265, 0.00104042, 0.0005747068, 
    0.001855823, 0.002421355, 0.005468251, 0.006023953, 0.00472714, 
    0.003903148, 0.002174302, 0.1503155, 0.03987028, 0.0003222166, 
    0.001113683, 0.003349919, 0.006100469, 0.008553299,
  1.386489e-07, -6.247046e-07, 9.482309e-06, 0.0001614137, 4.659837e-05, 
    0.005551241, 0.005132209, 0.0007901588, 0.04544385, 0.01726828, 
    0.003673549, 0.002236845, 0.0007467275, 0.0007680596, 0.0005159344, 
    0.0005240398, 0.001747886, 0.002232555, 0.01327826, 0.0359856, 
    0.007547427, 0.06073478, 0.0004328906, -0.0008190293, 0.0005773001, 
    0.001332778, 0.004570191, 0.007143068, -4.521299e-07,
  1.492068e-05, 0.003683703, 0.001531764, 0.002864806, 0.01680943, 
    0.003620575, -0.0005941327, 0.06628136, 0.1324662, 0.03958658, 
    0.06196363, 0.03676056, 0.03379262, 0.01971747, 0.02486716, 0.02636816, 
    0.01893907, 0.01455922, 0.02113272, 0.06163315, 0.01641759, 0.05975704, 
    0.02981534, 0.01339649, 0.01102859, 0.007084705, 0.004383638, 
    0.006988744, 0.008768908,
  0.00675064, 0.004290993, 0.0109416, 0.1939306, 0.004900216, 0.01223136, 
    0.0595542, 0.001060579, 0.001371195, 0.0175602, 0.1170618, 0.0773099, 
    0.1475672, 0.1513615, 0.1390166, 0.1283829, 0.1355959, 0.1068199, 
    0.07896983, 0.09990542, 0.04050552, 0.0486523, 0.07926573, 0.09804273, 
    0.05354019, 0.05368141, 0.0384062, 0.03428518, 0.05877679,
  0.07000513, 0.1401567, 0.1068318, 0.1360774, 0.09451854, 0.08268697, 
    0.03853188, 0.1213149, 0.04995925, 0.06385026, 0.06115667, 0.174352, 
    0.2335265, 0.2070467, 0.211346, 0.2106247, 0.2084703, 0.1764064, 
    0.1294239, 0.2071453, 0.05443889, 0.05000031, 0.09971158, 0.2633709, 
    0.1425522, 0.2144367, 0.1381091, 0.1098353, 0.1023334,
  0.08986107, 0.2189946, 0.1827927, 0.2668687, 0.28584, 0.1817055, 0.2194996, 
    0.2008122, 0.2154393, 0.2144707, 0.2331368, 0.2960595, 0.2184728, 
    0.1806544, 0.2312155, 0.272515, 0.3335475, 0.2253224, 0.2049448, 
    0.1530778, 0.243754, 0.1557565, 0.1774199, 0.2259534, 0.2680984, 
    0.08946219, 0.1246109, 0.1044107, 0.1079619,
  0.1746357, 0.09043361, 0.2283189, 0.116524, 0.2423009, 0.288835, 0.3552582, 
    0.2652686, 0.2074988, 0.2945686, 0.3618793, 0.2632573, 0.373555, 
    0.2943223, 0.3004293, 0.3090069, 0.2803321, 0.2219821, 0.263888, 
    0.2432229, 0.2927364, 0.4251347, 0.3061008, 0.3400313, 0.2239634, 
    0.2258478, 0.2733704, 0.1192774, 0.248288,
  0.4439245, 0.3036563, 0.3860673, 0.3929171, 0.4046144, 0.4602989, 
    0.4787011, 0.4597066, 0.4594316, 0.4705936, 0.4731014, 0.4607356, 
    0.4648682, 0.4655381, 0.4492551, 0.4631442, 0.4491397, 0.4516248, 
    0.4401252, 0.4449584, 0.434029, 0.2461146, 0.2590368, 0.3712737, 
    0.1444886, 0.1360709, 0.1197377, 0.2637493, 0.4088367,
  0.1061729, 0.1068213, 0.1074696, 0.108118, 0.1087663, 0.1094147, 0.110063, 
    0.09293592, 0.09673602, 0.1005361, 0.1043362, 0.1081363, 0.1119364, 
    0.1157365, 0.149237, 0.1487735, 0.14831, 0.1478464, 0.1473829, 0.1469194, 
    0.1464559, 0.1350376, 0.1310526, 0.1270677, 0.1230828, 0.1190978, 
    0.1151129, 0.111128, 0.1056543,
  0.190404, 0.1284906, 0.07559129, 0.07686892, 0.08472022, 0.05915213, 
    0.05971489, 0.06375529, 0.04533656, 0.04272433, 0.03858577, 0.06577154, 
    0.1310299, 0.003069258, 0.2517863, 0.2973473, 0.282537, 0.2336004, 
    0.1038047, 0.246944, 0.3832193, 0.4687526, 0.170629, 0.09428695, 
    0.2001731, 0.3216048, 0.1632578, 0.07726327, 0.1636422,
  0.1335589, 0.06139776, 0.08978777, 0.02345763, 0.04516557, 0.1054932, 
    0.02303977, 0.09834164, 0.1400277, 0.1265882, 0.1303441, 0.1435608, 
    0.05706754, 0.08554869, 0.2432711, 0.2585859, 0.2422606, 0.2286624, 
    0.2121032, 0.2369329, 0.2426013, 0.2671976, 0.2798328, 0.3188164, 
    0.2008806, 0.2957288, 0.2731737, 0.2245983, 0.2019602,
  0.2067792, 0.1757665, 0.1392641, 0.1246786, 0.1326181, 0.1492176, 
    0.1881524, 0.1567889, 0.1476947, 0.114984, 0.1258097, 0.1549028, 
    0.2105613, 0.1848797, 0.1398532, 0.1754434, 0.2116727, 0.2410011, 
    0.1852457, 0.1226952, 0.1124415, 0.0959277, 0.1068538, 0.1085079, 
    0.1886612, 0.2707402, 0.2717336, 0.2405135, 0.2238606,
  0.163925, 0.1564334, 0.159429, 0.158658, 0.1827699, 0.1721723, 0.1642972, 
    0.1105499, 0.1168375, 0.1026188, 0.06551263, 0.0616085, 0.04951178, 
    0.06347576, 0.09123223, 0.08761544, 0.08310705, 0.0917025, 0.09167363, 
    0.09257892, 0.07947873, 0.08660007, 0.07741427, 0.09535911, 0.03638536, 
    0.1077334, 0.1737903, 0.1702136, 0.1902089,
  0.05450317, 0.01868534, 0.01518289, 0.04041083, 0.04350709, 0.03853207, 
    0.04297788, 0.05319168, 0.04057811, 0.02047461, 0.01377972, 0.006177352, 
    0.007492334, 0.03021804, 0.1483727, 0.03534338, 0.04010858, 0.05359944, 
    0.05524307, 0.05684726, 0.05710233, 0.04872309, 0.02544576, 0.1823537, 
    0.01937451, 0.03603005, 0.05095507, 0.04829022, 0.05960816,
  0.006339298, 0.005625754, 0.008672649, 0.005270774, 0.007649852, 
    0.007180531, 0.006112327, 0.005608023, 0.008678652, 0.002915969, 
    0.0008985348, 0.000191359, 0.007139857, 0.003884721, 0.01120416, 
    0.01025606, 0.01549731, 0.02594185, 0.02184487, 0.008971285, 0.004396898, 
    0.003054829, 0.006487388, 0.009808507, 0.0174081, 0.009312003, 
    0.00906989, 0.002753821, 0.004487582,
  0.009991338, 0.01780625, 0.001288802, 0.001193398, -0.000945587, 
    0.0004524385, 0.0004919594, 0.001248943, 0.003840717, 0.001563327, 
    0.0008037965, 0.0002472346, 0.001158273, 0.002208445, 0.002172861, 
    0.001744057, 0.001280735, 0.001076061, 0.0006865753, 0.0005413705, 
    0.0004668276, 0.001866777, 0.009223084, 0.01493055, 0.01239141, 
    0.0557169, 0.0005765115, 0.0006543027, 0.002893248,
  0.02047492, 0.009665374, 0.01481282, 0.03824505, 0.0005238692, 0.000433386, 
    0.0005357471, 0.0004694356, 0.0005079355, 0.0004909615, 0.002808291, 
    0.0004084657, 0.003895989, 0.0003210017, 0.0005417273, 0.0004109887, 
    0.0001820491, 0.0002703817, 0.0002066047, 0.0003192629, 0.001045387, 
    0.004611037, 0.02177737, 0.01007608, 0.01077133, 0.003768968, 
    4.887387e-06, 0.0009308763, 0.005373,
  0.004690881, 0.0370631, 0.006012633, 0.01431957, 0.001011526, 0.0009268499, 
    0.001233167, 0.0007858764, 0.03143744, 0.05849371, 0.0005940183, 
    0.0009624242, 0.001046252, 0.0006039204, 0.000778647, 0.0002817915, 
    0.0003749051, 0.000346075, 0.0005403742, 0.0008664216, 0.002099593, 
    0.01669153, 0.03389728, 0.01805619, 0.01128665, 0.001222796, 0.001214268, 
    0.0005980625, 0.003448957,
  0.001577734, 0.00282236, 9.759539e-05, 0.03013927, 0.006175822, 
    0.0006998834, 0.004108732, 0.0005374471, 0.000210496, 0.0005735327, 
    0.001199686, 0.0006608821, 0.0005229277, 0.0005414338, 0.000303244, 
    0.000908747, 0.001138796, 0.002607525, 0.002856789, 0.00232402, 
    0.001880286, 0.001077234, 0.1199433, 0.03418938, 0.0001732377, 
    0.0006660205, 0.002183948, 0.003820686, 0.005875009,
  1.349498e-07, -3.448899e-07, 6.963425e-06, 0.0001053707, 2.284691e-05, 
    0.003727647, 0.003454688, 0.0004739241, 0.03566806, 0.01040246, 
    0.002059952, 0.001231834, 0.000490714, 0.0004973788, 0.0003707508, 
    0.0003883623, 0.0009989801, 0.001409217, 0.009008166, 0.02469709, 
    0.005130142, 0.05022812, 0.0003260249, -0.0009177474, 0.0003899542, 
    0.0008651611, 0.003292728, 0.004669751, -8.787202e-07,
  1.02186e-05, 0.002758037, 0.001020787, 0.002152499, 0.01441802, 
    0.002925089, -0.0001462434, 0.0665143, 0.1227133, 0.02804506, 0.04503413, 
    0.0221029, 0.02014759, 0.01185991, 0.01583228, 0.01610493, 0.01213794, 
    0.009058608, 0.01394561, 0.04881943, 0.01402394, 0.05065568, 0.02566888, 
    0.007580475, 0.006275687, 0.004303327, 0.003101742, 0.004982506, 
    0.006971853,
  0.005290062, 0.003495242, 0.008287036, 0.1797443, 0.003981825, 0.009944871, 
    0.05349898, 0.001094004, 0.0009034296, 0.01587181, 0.1046454, 0.06433615, 
    0.1180321, 0.122595, 0.105248, 0.0942124, 0.09483419, 0.07235821, 
    0.05383651, 0.09053266, 0.03689485, 0.04169626, 0.06660604, 0.08115555, 
    0.03633756, 0.03214136, 0.02214486, 0.02098542, 0.04349105,
  0.05383373, 0.1228396, 0.0923049, 0.1190079, 0.0813354, 0.07314107, 
    0.0322353, 0.1161476, 0.06124386, 0.0583362, 0.05572086, 0.1634333, 
    0.197212, 0.1710787, 0.1699228, 0.1602687, 0.1577931, 0.1293967, 
    0.09167042, 0.1965989, 0.04577905, 0.04021933, 0.08475645, 0.2356351, 
    0.1271345, 0.1865427, 0.1022205, 0.07630954, 0.06961136,
  0.06777395, 0.2131294, 0.1644593, 0.2390015, 0.2595299, 0.1592703, 
    0.1910389, 0.1722016, 0.1875439, 0.1836764, 0.2052668, 0.3111998, 
    0.2295514, 0.1700893, 0.1952862, 0.2217054, 0.3175851, 0.2060316, 
    0.1911165, 0.1457043, 0.2228158, 0.1561924, 0.1443472, 0.2173071, 
    0.2367785, 0.07678635, 0.09140168, 0.07281598, 0.07942481,
  0.1324579, 0.06919754, 0.2262751, 0.09496024, 0.2177773, 0.2550706, 
    0.3335961, 0.2559783, 0.2271984, 0.2917474, 0.3531725, 0.2418877, 
    0.3473105, 0.2395788, 0.2523866, 0.2651357, 0.2591653, 0.1930442, 
    0.2416471, 0.204798, 0.2527862, 0.379479, 0.2759193, 0.3401682, 
    0.2068173, 0.1882063, 0.3054264, 0.1061118, 0.2033974,
  0.4186822, 0.2875506, 0.3468316, 0.3351718, 0.342614, 0.3781308, 0.3764443, 
    0.353056, 0.3644704, 0.3571201, 0.3502035, 0.3416845, 0.3422742, 
    0.3415573, 0.3335353, 0.3468263, 0.3401979, 0.3436601, 0.3233635, 
    0.3307891, 0.3345158, 0.2209394, 0.2519443, 0.4013867, 0.1363991, 
    0.1099993, 0.114069, 0.24808, 0.3489218,
  0.07781415, 0.07808875, 0.07836334, 0.07863792, 0.07891251, 0.0791871, 
    0.07946169, 0.06739618, 0.07076774, 0.07413929, 0.07751085, 0.08088241, 
    0.08425396, 0.08762552, 0.1129076, 0.1128496, 0.1127917, 0.1127337, 
    0.1126757, 0.1126178, 0.1125598, 0.107113, 0.1035249, 0.09993669, 
    0.09634852, 0.09276035, 0.08917217, 0.085584, 0.07759449,
  0.1565333, 0.09634557, 0.05568308, 0.06098904, 0.06662235, 0.05061504, 
    0.04828269, 0.05339696, 0.03936224, 0.03590476, 0.03048497, 0.05721033, 
    0.1153735, 0.003071262, 0.2826219, 0.2603983, 0.255891, 0.2478797, 
    0.1063286, 0.2666916, 0.3720236, 0.4670913, 0.1638463, 0.09155796, 
    0.1856752, 0.3137435, 0.1663452, 0.07732617, 0.1402474,
  0.1286774, 0.06009919, 0.08432642, 0.0216364, 0.04144895, 0.09542956, 
    0.02160467, 0.09097686, 0.1316558, 0.1191328, 0.1232945, 0.1410844, 
    0.05371585, 0.07981884, 0.2274813, 0.236505, 0.2203997, 0.2069264, 
    0.187395, 0.2136591, 0.218545, 0.2433181, 0.2546427, 0.2920966, 
    0.1867763, 0.2673677, 0.2440919, 0.1986285, 0.1817661,
  0.1823839, 0.1545518, 0.121058, 0.1084337, 0.1141008, 0.1301099, 0.1668184, 
    0.1385042, 0.1280122, 0.09762742, 0.1067372, 0.1313736, 0.1793649, 
    0.1554185, 0.1154573, 0.1479579, 0.1810942, 0.2076784, 0.157938, 
    0.1032956, 0.09361651, 0.07859033, 0.08735628, 0.08863006, 0.1582891, 
    0.2355952, 0.2430746, 0.2131567, 0.1985036,
  0.1389153, 0.1324478, 0.1340312, 0.1318211, 0.1548736, 0.1455549, 
    0.1390467, 0.09261928, 0.09816059, 0.08547846, 0.05198846, 0.04783512, 
    0.03772956, 0.04829848, 0.07101516, 0.0676044, 0.06298637, 0.06897104, 
    0.07017223, 0.07162423, 0.06215072, 0.06748319, 0.06122945, 0.1098284, 
    0.02892515, 0.08600739, 0.1435344, 0.1438053, 0.16177,
  0.0405577, 0.0135814, 0.01085125, 0.02866891, 0.03087831, 0.02691892, 
    0.03063507, 0.03859571, 0.02852544, 0.0150448, 0.009829603, 0.004813833, 
    0.00542044, 0.02153507, 0.146685, 0.02437139, 0.02744386, 0.03840372, 
    0.03958052, 0.04079387, 0.04120843, 0.03468727, 0.01807296, 0.1819225, 
    0.0154145, 0.02592552, 0.03672411, 0.03530253, 0.04354554,
  0.004983461, 0.00452235, 0.011255, 0.003708491, 0.004933278, 0.004765176, 
    0.004282269, 0.004200036, 0.006820509, 0.002448536, 0.0006230119, 
    0.000451792, 0.0110094, 0.00262645, 0.006860797, 0.006230305, 
    0.009537755, 0.01632882, 0.01412591, 0.005658807, 0.002936817, 
    0.002320895, 0.005379266, 0.008232372, 0.0235619, 0.006053329, 
    0.005443814, 0.001969134, 0.003385082,
  0.008261831, 0.01426928, 0.001997243, 0.0009666129, -0.001004599, 
    0.0003290032, 0.0003823795, 0.0009459003, 0.003108562, 0.001237309, 
    0.0007540418, 0.0002746799, 0.0008833139, 0.0014955, 0.00140585, 
    0.001207795, 0.0009417183, 0.000788386, 0.0004648519, 0.0003792829, 
    0.0003786186, 0.001539373, 0.007624513, 0.01256112, 0.02104632, 
    0.07821541, 0.000422639, 0.0005357583, 0.002349988,
  0.01674197, 0.006996633, 0.02881872, 0.06779411, 0.0003754044, 0.000321661, 
    0.0003727585, 0.0003221766, 0.0004001678, 0.0002787234, 0.002158432, 
    0.0002920181, 0.002530328, 0.0002386071, 0.0003616177, 0.0002816904, 
    0.0001367528, 0.0002081157, 0.0001711868, 0.0002669471, 0.0008715685, 
    0.003804503, 0.01788475, 0.05199997, 0.02565769, 0.01333644, 
    -6.100679e-06, 0.0007683743, 0.0044048,
  0.003727725, 0.06552418, 0.008288094, 0.01482376, 0.0007451493, 
    0.0006724227, 0.0008681536, 0.0005755849, 0.04771128, 0.08976738, 
    0.0004295734, 0.0007416051, 0.0006983199, 0.0004047671, 0.000512176, 
    0.0002271692, 0.000291354, 0.0002778232, 0.0004252207, 0.0006809832, 
    0.001619112, 0.01308507, 0.02710365, 0.04514832, 0.037676, 0.000794159, 
    0.0007314634, 0.0004712367, 0.002695156,
  0.01194498, 0.003250527, 0.0001098644, 0.03070533, 0.004643384, 
    0.000584485, 0.00604035, 0.0004233015, -0.0007601702, 0.0004290951, 
    0.0007819053, 0.0004842766, 0.0003520739, 0.0003777661, 0.0002211356, 
    0.000572925, 0.0007090537, 0.001609439, 0.001766869, 0.001545087, 
    0.001212713, 0.000708058, 0.1611309, 0.03728749, 0.0001254757, 
    0.0005056842, 0.001706782, 0.002894412, 0.01612127,
  1.337212e-07, -1.997797e-07, 5.383104e-06, 8.030561e-05, 1.434335e-05, 
    0.002856708, 0.003655246, 0.0003332748, 0.05740475, 0.006831106, 
    0.001446541, 0.0008561384, 0.0003815699, 0.0003891608, 0.000307394, 
    0.0003256546, 0.0007191995, 0.001090777, 0.00696549, 0.01919012, 
    0.003922973, 0.04586766, 0.000275202, -0.001386071, 0.0003094568, 
    0.000677984, 0.002693363, 0.003627159, -5.524289e-07,
  7.803445e-06, 0.002274597, 0.0008557306, 0.001977149, 0.01377049, 
    0.002632699, 0.000837922, 0.08184307, 0.1303765, 0.02536125, 0.03201563, 
    0.01402529, 0.01327787, 0.00800073, 0.0109023, 0.01066881, 0.008182499, 
    0.006162437, 0.01057628, 0.04153075, 0.01245653, 0.06242096, 0.04052068, 
    0.005145658, 0.003996746, 0.003103473, 0.002459092, 0.004034871, 
    0.005875072,
  0.005394003, 0.002937131, 0.00704497, 0.1788108, 0.003434506, 0.008627504, 
    0.05237505, 0.001300797, 0.0007516273, 0.01571387, 0.1112186, 0.05022641, 
    0.09287222, 0.09268157, 0.07911246, 0.0705684, 0.07121255, 0.05219309, 
    0.03890412, 0.0879076, 0.03736332, 0.04056641, 0.06859598, 0.06721907, 
    0.02775194, 0.02167247, 0.01469472, 0.01449631, 0.03621585,
  0.04489202, 0.12434, 0.09330691, 0.1171943, 0.07558893, 0.06937321, 
    0.0303218, 0.1479461, 0.09748019, 0.06467092, 0.07681773, 0.1828327, 
    0.1665679, 0.1425036, 0.1376292, 0.1267739, 0.1232174, 0.09974075, 
    0.06884591, 0.2050433, 0.04474035, 0.0397696, 0.09477796, 0.2471984, 
    0.1228635, 0.157921, 0.0797577, 0.05738651, 0.05144328,
  0.05453246, 0.2480256, 0.1683238, 0.2365031, 0.2700579, 0.1768003, 
    0.1969375, 0.1860476, 0.210489, 0.1982705, 0.2110114, 0.3567905, 
    0.2692175, 0.182674, 0.1700493, 0.1916282, 0.3370385, 0.2032335, 
    0.2187306, 0.1659578, 0.2222048, 0.1769047, 0.1233532, 0.2355272, 
    0.214805, 0.06848948, 0.07320996, 0.05654976, 0.06335582,
  0.1062014, 0.05614967, 0.2540846, 0.07833936, 0.2012275, 0.2380518, 
    0.324703, 0.2678935, 0.2679998, 0.2973441, 0.3711534, 0.2785921, 
    0.318621, 0.216809, 0.2312089, 0.2339382, 0.2690991, 0.1926734, 
    0.2282941, 0.1857854, 0.2275272, 0.3452947, 0.2616279, 0.3467202, 
    0.1898732, 0.170351, 0.3484495, 0.09808543, 0.1684205,
  0.3999889, 0.2715926, 0.314945, 0.2846454, 0.2879981, 0.3213643, 0.3113503, 
    0.28813, 0.3005413, 0.2830135, 0.274259, 0.2636993, 0.2661233, 0.2686609, 
    0.2619899, 0.2753419, 0.2707057, 0.2733123, 0.2594999, 0.2682944, 
    0.2724241, 0.2059829, 0.2617159, 0.4171001, 0.132534, 0.09806781, 
    0.1171735, 0.2488771, 0.3062815 ;

 average_DT = 720 ;

 average_T1 = 350.5 ;

 average_T2 = 1080.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 715.5 ;

 time_bnds =
  350.5, 1080.5 ;
}
