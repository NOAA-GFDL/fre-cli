netcdf atmos_month.198001-198012.alb_sfc {
dimensions:
	time = UNLIMITED ; // (12 currently)
	lat = 2 ;
	lon = 2 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_methods = "time: mean" ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:10 2025" ;
		:hostname = "pp033" ;
		:history = "Tue Sep 23 14:27:36 2025: ncks -d lon,0,1 atmos_month.198001-198012.alb_sfc.nc_lat01 atmos_month.198001-198012.alb_sfc.nc_lat01_lon01\n",
			"Tue Sep 23 14:26:17 2025: ncks -d lat,0,1 atmos_month.198001-198012.alb_sfc.nc atmos_month.198001-198012.alb_sfc.nc_lat01\n",
			"Mon Aug 11 16:13:43 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198001-198012.alb_sfc.nc reduced/atmos_month.198001-198012.alb_sfc.nc\n",
			"Mon Aug 11 20:02:14 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.3.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.21249, 76.21249,
  76.5369, 76.35718,
  76.45917, 76.45917,
  73.2886, 73.07695,
  47.00509, 47.00509,
  43.41802, 43.26198,
  0, 0,
  10.06781, 10.30963,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  2.493829, 2.492429,
  20.90129, 20.90129,
  33.09964, 33.03193,
  76.34792, 76.34792,
  64.8836, 64.57207,
  76.27164, 76.27164,
  76.35242, 76.16932,
  76.13555, 76.13555,
  76.35452, 76.19527 ;

 lat = -89.5, -79.5 ;

 lat_bnds =
  -90, -89,
  -80, -79 ;

 lon = 0.625, 13.125 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75 ;

 time = 380.5, 410.5, 440.5, 471, 501.5, 532, 562.5, 593.5, 624, 654.5, 685, 
    715.5 ;

 time_bnds =
  365, 396,
  396, 425,
  425, 456,
  456, 486,
  486, 517,
  517, 547,
  547, 578,
  578, 609,
  609, 639,
  639, 670,
  670, 700,
  700, 731 ;
}
