netcdf \20030101.atmos_static_cmip.tile5 {
dimensions:
	grid_xt = 96 ;
	grid_yt = 96 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:associated_files = "area: 20030101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 time = 0 ;

 orog =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01534718, 
    0.004565009, 0.008999515, 0.009599131, 0.0008479413, 0, 0, 0.0007195598, 
    0.004574103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7068716, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003399682, 
    0.0147934, 0.002706561, 0, 0, 0, 0.004826599, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004755895, 
    0.00314351, 0.002793752, 0, 0, 0, 0.006179405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006290677, 
    0.007201957, 0, 0.01463142, 0.003162183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008779748, 0, 0, 0, 
    0.00300725, 0.002690252, 0.005241457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.506357, 3.305288, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.007343553, 0, 0.009825814, 0.01535672, 0.006712195, 0, 0, 0.005644962, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19.68891, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008339305, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00178691, 18.51452, 0.01244308, 0, 0, 0, 
    0, 0.009080717, 0, 0, 0, 0, 0.006611669, 0.003060021, 0.008406991, 0, 
    0.005074322, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01017599, 
    0, 0, 0, 0.004030156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003469607, 0, 0, 0, 0, 0, 0.002995649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004560474, 0, 0, 0.01124365, 0.003597797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01154227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2431989, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.001374771, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.06463672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1425494, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  33.14798, 0, 34.79201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0004971988, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  668.3605, 750.8135, 625.5392, 386.1679, 158.3386, 2.453814, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1070.732, 1178.2, 1004.681, 772.6516, 403.6846, 150.0447, 26.30301, 
    1.64736, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1507.715, 1421.274, 1144.302, 833.4024, 441.414, 72.99273, 109.9673, 
    184.5779, 220.3756, 0.00647221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1551.811, 1623.509, 1564.146, 1482.56, 1154.821, 803.4989, 487.0388, 
    202.9149, 268.4435, 226.8269, 46.07853, 0.3954178, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1557.897, 1671.874, 1696.626, 1635.232, 1700.021, 1734.235, 1559.076, 
    995.3284, 449.7531, 276.2559, 565.8065, 21.12218, 0.8193069, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1468.874, 1600.571, 1614.583, 1414.91, 1396.924, 1757.31, 2173.984, 
    2018.616, 1396.95, 1025.211, 762.0422, 232.5291, 8.014444, 1.140886, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1326.019, 1541.283, 1555.617, 1480.098, 1514.677, 1689.735, 1982.568, 
    2007.651, 1670.599, 1186.88, 1048.513, 684.1181, 117.3529, 0.1669138, 0, 
    0, 0, 14.15248, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1146.4, 1447.466, 1700.664, 1654.412, 1747.869, 2042.93, 1975.362, 
    1731.381, 1260.238, 1003.032, 874.1664, 965.1847, 711.4643, 390.3766, 
    173.5833, 3.412067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1373.781, 1329.12, 1740.19, 1867.481, 1919.821, 2046.155, 2020.59, 
    1730.883, 1388.832, 990.3948, 863.0721, 733.3089, 488.1863, 444.3896, 
    642.3708, 630.8365, 208.2363, 11.2473, 0.03753853, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1914.861, 1386.722, 1730.161, 1876.041, 1894.845, 2047.599, 1965.026, 
    1787.49, 1283.865, 1007.386, 831.1433, 589.1078, 291.1984, 130.3001, 
    245.2175, 308.7728, 423.5323, 287.8249, 17.96172, 32.98395, 0.1041703, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1970985, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  2061.196, 1476.068, 1648.332, 1574.314, 1569.191, 1744.371, 1828.933, 
    1790.968, 1558.644, 1149.688, 1213.996, 906.5831, 504.1509, 233.0578, 
    183.2224, 38.9668, 0.0118664, 233.6236, 272.1967, 144.2618, 56.46022, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1840.156, 1504.441, 1582.167, 1490.926, 1402.836, 1518.827, 1694.572, 
    2058.519, 1824.339, 1671.718, 1643.01, 1482.167, 815.0604, 396.3656, 
    379.8361, 318.8223, 100.745, 65.86816, 107.3457, 244.7698, 250.1199, 
    15.35586, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1837.63, 1728.632, 1902.097, 1719.298, 1875.763, 1918.201, 2012.239, 
    2196.799, 2065.854, 1799.648, 1839.158, 1689.026, 1220.946, 556.4898, 
    653.7017, 762.9083, 615.2339, 393.6399, 83.12075, 4.564439, 169.0518, 
    231.0936, 86.59752, 8.810427, 0, 0, 0, 0, 0.004199471, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2287.553, 2375.422, 2227.182, 2205.671, 2448.729, 2173.713, 2069.91, 
    1804.564, 1718.86, 1645.912, 1760.087, 1774.775, 1588.443, 1158.239, 
    1042.855, 1238.964, 1055.679, 720.4163, 300.8953, 74.61289, 2.083953, 
    10.21264, 134.772, 93.68505, 9.525565, 0, 0, 0, 0.06281511, 3.428892, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2614.957, 2546.323, 2390.928, 2148.965, 2257.577, 2052.22, 1766.787, 
    1770.134, 1673.074, 1765.732, 1825.648, 1895.919, 1992.829, 1695.072, 
    1362.996, 1422.211, 1302.389, 1040.16, 627.5578, 400.1667, 51.56722, 
    2.257818, 0.1849899, 56.72547, 250.1037, 1.460486, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.967957, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1897.78, 2076.201, 2129.073, 2115.72, 2166.538, 1872.045, 2072.919, 
    1904.649, 2256.727, 1803.393, 1983.677, 2108.663, 2195.764, 2050.119, 
    1605.954, 1432.204, 1511.048, 1487.268, 1426.227, 1196.583, 721.2061, 
    185.3391, 24.12744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004704067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2958491, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1716.921, 1748.802, 1939.11, 2058.646, 2214.479, 2215.264, 2299.508, 
    2683.908, 2679.552, 2308.606, 2102.935, 2086.155, 2177.915, 2051.186, 
    1598.307, 1383.17, 1438.509, 1773.132, 2076.03, 2118.625, 1700.985, 
    1170.254, 459.9845, 48.66238, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1594.9, 1717.709, 1846.341, 2183, 2416.479, 2646.638, 2920.714, 2901.701, 
    3107.744, 2624.682, 2306.014, 2028.034, 1806.9, 1723.413, 1505.019, 
    1253.708, 1291.276, 1617.983, 1898.304, 2037.906, 2075.454, 2108.36, 
    1570.701, 841.1761, 129.8114, 0.2389687, 3.660637, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1414.581, 1499.586, 1735.549, 1988.982, 2430.141, 2544.231, 2714.589, 
    2826.258, 2566.761, 2620.082, 2419.738, 2052.477, 1891.764, 1767.929, 
    1617.863, 1432.407, 1338.126, 1367.179, 1424.379, 1473.549, 1661.907, 
    2049.929, 2230.574, 1919.274, 1373.336, 316.5095, 39.45748, 94.61289, 
    39.49365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.207365e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1235.553, 1437.662, 1381.895, 1611.005, 1679.951, 1728.312, 1922.424, 
    1964.016, 1953.016, 2112.162, 2098.977, 1710.801, 1526.079, 1414.803, 
    1368.911, 1237.472, 1292.035, 1341.555, 1204.039, 1329.621, 1429.259, 
    1572.953, 1800.086, 2189.089, 2119.821, 1455.417, 1083.626, 1022.557, 
    862.4561, 51.87525, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1174.93, 1228.427, 1291.553, 1290.888, 1424, 1351.69, 1468.16, 1589.555, 
    1427.788, 1689.11, 1630.9, 1414.054, 1334.024, 1248.547, 1122.594, 
    1033.518, 1091.201, 1192.766, 1168.232, 1309.946, 1314.83, 1245.706, 
    1400.043, 1858.552, 2194.833, 2118.342, 1668, 1707.535, 1364.425, 
    595.4224, 15.76594, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  823.5144, 966.8268, 1033.309, 1192.71, 1210.489, 1193.993, 1280.92, 
    1308.805, 1209.215, 1289.174, 1294.622, 1176.932, 1193.732, 1146.91, 
    1025.355, 875.7115, 882.8735, 978.463, 1033.714, 1232.486, 1255.239, 
    1216.565, 1342.363, 1716.272, 2074.805, 2120.552, 2071.005, 1786.363, 
    1785.419, 844.6271, 169.2518, 0.001837272, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  661.3832, 741.7489, 952.168, 1073.759, 1053.268, 1013.894, 1031.548, 
    1062.557, 1014.31, 1013.214, 1007.304, 1006.718, 987.2679, 929.3942, 
    846.1819, 807.7843, 729.1191, 717.0919, 644.5469, 733.0809, 815.4983, 
    1055.672, 1469.535, 1941.911, 2045.901, 2101.024, 2062.683, 2086.129, 
    1883.878, 989.241, 529.9884, 1.092551, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  574.1776, 618.1168, 795.5441, 907.0357, 894.5935, 851.0385, 820.7712, 
    843.4498, 837.6264, 813.8089, 821.1804, 790.303, 694.8225, 637.4512, 
    626.2227, 661.035, 688.275, 597.9715, 427.0944, 299.6628, 342.4961, 
    676.9834, 1214.729, 1706.491, 1881.969, 1649.495, 1733.168, 2044.59, 
    2105.82, 1415.646, 915.3256, 166.6185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  503.9159, 538.9011, 631.793, 737.8944, 750.1324, 703.1216, 655.9878, 
    654.8143, 672.593, 642.7423, 621.7355, 602.098, 473.79, 425.5311, 
    461.755, 530.6566, 568.3069, 558.3639, 330.7892, 179.9599, 143.326, 
    168.8803, 392.449, 875.6781, 1042.997, 940.2807, 1005.778, 1682.482, 
    2467.645, 1832.106, 1341.977, 441.4869, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  453.9662, 441.7195, 504.0019, 592.8539, 608.1069, 578.1291, 526.2635, 
    513.4938, 532.1535, 479.4901, 447.4254, 444.3315, 379.7191, 325.8571, 
    347.1577, 396.39, 397.7914, 382.2119, 225.9507, 114.7197, 95.74188, 
    70.67721, 57.3841, 157.933, 314.682, 123.271, 156.6136, 1009.174, 
    2106.859, 2219.086, 1513.035, 924.8544, 29.27477, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  503.6515, 465.5753, 433.9768, 478.4191, 482.0991, 473.893, 436.3061, 
    425.1155, 431.4804, 382.6123, 325.8517, 340.3661, 314.822, 260.5178, 
    239.2539, 233.0164, 209.3085, 185.2675, 99.46118, 35.69082, 15.04999, 
    5.81494, 7.321244, 7.285094, 10.49513, 6.034019, 12.30279, 178.9217, 
    1494.86, 1747.576, 1843.446, 1614.362, 380.1558, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  438.2668, 471.7402, 408.1164, 400.8929, 380.3304, 374.7529, 382.5601, 
    372.2382, 382.916, 320.6809, 264.4974, 252.2818, 258.8326, 194.5873, 
    162.8055, 141.8769, 114.3217, 85.31949, 39.80796, 4.830305, 0, 0, 0, 0, 
    0, 0, 0, 0.02132653, 176.2921, 430.069, 932.7458, 1392.24, 747.5593, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  375.052, 414.3507, 415.5859, 381.3595, 361.0887, 329.3397, 313.1617, 
    313.8601, 298.01, 280.3281, 250.9803, 220.6591, 244.4896, 157.4741, 
    126.7682, 118.9209, 91.80339, 46.5208, 11.15798, 0.09899135, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50.89595, 153.9082, 606.8809, 122.0387, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  304.4448, 364.8189, 357.5074, 352.7218, 337.0601, 318.3467, 277.0119, 
    265.5412, 282.2703, 328.1339, 341.168, 288.7758, 254.3146, 138.1611, 
    97.54157, 97.74657, 73.76514, 23.01658, 0.5496842, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.476873, 75.94135, 449.1298, 34.83492, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  306.857, 361.5244, 342.5269, 300.4066, 292.6741, 274.3279, 251.7741, 
    245.3346, 294.167, 380.9618, 372.6419, 271.2439, 204.3829, 99.51021, 
    69.604, 73.45421, 50.67704, 12.05578, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.512501, 149.8454, 851.515, 526.5105, 5.040119, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  319.7339, 346.4661, 325.2934, 268.1579, 235.2851, 243.1511, 224.0061, 
    242.3429, 319.4263, 334.612, 274.955, 164.2817, 109.9028, 55.26638, 
    47.65622, 41.80495, 35.97699, 2.775469, 0.03288275, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6.357764, 280.3884, 1031.42, 1222.137, 606.0325, 0.7514994, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07952388, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  294.8905, 319.0948, 294.4915, 238.6062, 212.2333, 193.6535, 202.8654, 
    221.7048, 288.9077, 248.9493, 137.382, 84.58096, 51.21586, 40.6296, 
    44.39739, 63.04242, 40.62316, 8.783824, 0.268134, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.7404718, 15.12963, 65.80754, 738.6376, 1257.209, 1292.93, 64.7064, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13.92286, 118.2891, 0.07517834, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  313.3622, 298.425, 277.4745, 233.6075, 198.1856, 187.4898, 173.2009, 
    175.6373, 200.6465, 144.9214, 80.57291, 77.81576, 66.51388, 73.39558, 
    92.76784, 95.03912, 61.3536, 3.831983, 0.1158118, 0, 0, 0, 0, 0, 0, 0, 
    0.6463583, 18.92656, 71.69862, 132.442, 95.90388, 289.954, 763.129, 
    1148.201, 229.1096, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.065996, 
    17.50426, 2.459143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  289.323, 276.3043, 265.5132, 220.7219, 216.1242, 195.0884, 181.3391, 
    143.4675, 147.2648, 111.0426, 110.6656, 125.9561, 122.3719, 105.6208, 
    113.7486, 98.84241, 43.68995, 0.9661562, 0.02680171, 0, 0, 0, 0, 0, 0, 0, 
    3.878528, 38.69389, 97.16181, 132.8956, 207.0652, 216.3446, 424.0393, 
    918.3037, 351.0448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.011113, 
    0.1137814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  230.5823, 241.4872, 225.9881, 214.9098, 207.3458, 206.6044, 173.4783, 
    138.0395, 130.4559, 142.9235, 167.6159, 175.7432, 143.494, 103.3232, 
    73.60364, 63.91725, 27.10206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.20466, 
    20.16096, 25.27402, 21.63544, 14.64767, 43.60937, 331.3476, 893.1275, 
    454.1429, 1.288543, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  191.6571, 178.5321, 189.9285, 201.3738, 214.7888, 215.5745, 179.5497, 
    147.2228, 153.1658, 179.6961, 230.3224, 239.8835, 194.1318, 137.8888, 
    87.66043, 69.8594, 27.32165, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.084438, 
    6.930506, 0.584422, 0.003764597, 0.003457344, 0.4655042, 543.0778, 
    932.6347, 615.3885, 85.28525, 0.2777186, 0, 0, 0, 0, 0, 0.422377, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  231.2289, 207.4846, 224.9596, 237.2916, 248.9516, 252.8323, 212.7034, 
    195.5234, 197.4957, 263.0653, 303.2209, 280.5213, 264.7434, 194.2222, 
    116.7919, 78.11273, 25.05218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.827813, 526.7432, 777.7427, 639.5916, 362.6419, 79.72997, 29.67748, 
    0.912546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  278.9553, 267.2621, 269.6895, 261.4806, 287.7636, 281.252, 243.8186, 
    240.3938, 298.7545, 342.4502, 399.08, 363.9893, 266.6101, 221.5975, 
    126.7727, 76.75681, 26.75876, 0.9402217, 0, 0, 0, 0, 0, 0, 0, 0.3805751, 
    0, 0, 0, 0, 0, 3.231741, 309.7996, 351.9758, 387.7886, 218.6437, 153.275, 
    263.9878, 54.07672, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  241.8856, 246.4237, 245.6055, 259.1919, 286.3187, 285.9484, 254.3894, 
    280.3928, 369.3888, 439.415, 618.7897, 387.4653, 291.7344, 174.3447, 
    113.5729, 67.22175, 24.12755, 0, 0, 0, 0, 0, 0, 0, 20.0383, 16.96434, 0, 
    0, 0, 0, 0.003687347, 0.00572379, 52.21835, 70.8857, 55.61906, 70.92522, 
    123.4313, 420.684, 636.3296, 6.528507, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  202.4083, 219.8558, 207.086, 261.2129, 295.0167, 264.0109, 249.5903, 
    352.6951, 497.0891, 679.3617, 595.9517, 404.6982, 150.7021, 114.5868, 
    78.8996, 54.99938, 26.96955, 5.426031, 1.965392, 0.1738949, 0, 0, 0, 0, 
    39.73782, 6.958992, 0, 0, 0, 0, 0, 0.0001729098, 1.584328, 6.905681, 
    0.7596173, 0.490705, 0, 84.19572, 863.5649, 289.1957, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  210.9862, 176.5489, 218.8383, 299.7639, 293.6812, 247.376, 300.3907, 
    490.8528, 720.3207, 577.838, 503.2361, 148.1991, 107.7899, 63.81637, 
    42.55847, 31.07135, 27.5754, 28.17957, 28.8343, 16.63614, 2.660592, 0, 
    0.01031376, 0.9608897, 33.86351, 0.509288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05132846, 0, 0, 160.5816, 333.4066, 8.909275, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  247.1366, 214.9977, 272.471, 323.8452, 298.5703, 362.521, 537.7053, 
    668.5198, 624.8367, 453.5524, 165.6625, 102.4959, 57.48196, 21.7608, 
    4.573749, 1.787246, 5.738702, 13.79587, 21.61514, 15.3555, 7.805641, 
    1.753023, 0.05135195, 1.186182, 39.27137, 0.8040789, 0, 0.01927231, 
    0.09756799, 0, 0, 0, 0, 0, 0.1619276, 0, 0, 0, 9.406398, 314.6326, 
    92.01137, 0, 0, 0.001729056, 0, 0, 0, 0, 0.6381596, 31.72947, 4.45034, 
    6.862898, 161.6274, 35.41436, 10.87154, 0.005455857, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.744836, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  229.433, 306.0153, 351.427, 376.3137, 463.0498, 627.9566, 686.7066, 
    565.6674, 405.129, 181.5926, 102.0433, 47.04384, 16.67009, 1.10613, 0, 0, 
    0, 0.09115441, 1.67472, 5.002741, 3.653378, 0.914476, 0.0004763628, 
    1.392298, 81.95518, 36.95679, 0, 0.102858, 0, 0, 0, 0, 0, 7.409501e-05, 
    0, 0, 0, 0, 55.38284, 97.32481, 47.17434, 0, 0, 0, 0, 0, 0.03468706, 
    60.15501, 130.7003, 244.7536, 135.677, 424.9022, 731.8262, 553.5016, 
    151.7469, 15.67891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1039039, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.4516, 455.0074, 496.0555, 490.0974, 549.4736, 625.2988, 487.0647, 
    277.1122, 157.1025, 104.1153, 47.97492, 9.955524, 1.711641, 0, 0, 0, 0, 
    0, 0, 0.08672119, 0.02051163, 0.0005947647, 0, 0.02029713, 58.99087, 
    18.83587, 0.0248516, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 110.5765, 3.497101, 
    0, 0, 0, 0, 0, 0.05597858, 47.99405, 655.0215, 1362.752, 1510.303, 
    1890.99, 1900.117, 1904.355, 1649.458, 1608.771, 1245.189, 378.5316, 
    4.13827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.282194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  430.407, 573.2601, 458.0574, 384.715, 322.2038, 270.0156, 169.9159, 
    89.97162, 81.54353, 47.91539, 13.97083, 0.9449826, 0, 0, 0, 0, 0, 0, 
    0.0004252571, 0.3309443, 0.03876647, 1.728635, 0.4185002, 0, 15.5728, 
    39.27885, 1.380751, 0.007368555, 55.84319, 1.191139, 0, 0, 0, 0, 0, 0, 0, 
    0, 115.976, 114.2675, 74.08803, 0, 0, 0, 0.3069585, 74.61648, 1023.105, 
    1976.442, 2391.624, 2180.577, 1604.411, 1326.77, 901.5997, 1351.656, 
    2254.224, 2631.384, 2637.751, 1822.456, 620.1605, 20.8799, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  430.7066, 471.0601, 333.3573, 224.1613, 108.1152, 65.5984, 26.94351, 
    37.64307, 24.10448, 10.83371, 1.795868, 0, 0, 0, 0, 0, 0, 0, 0, 0.421066, 
    0.211959, 0.211567, 0.4754283, 0, 1.457668, 49.35142, 77.70663, 0.225208, 
    177.6199, 27.2492, 0, 0, 0, 0, 0, 0, 0, 0, 16.10499, 144.5139, 247.1739, 
    155.9424, 68.87181, 112.7537, 548.5216, 1326.625, 1537.927, 1522.117, 
    1053.582, 538.7177, 494.4248, 237.3714, 225.9437, 723.8336, 1495.832, 
    2103.182, 2873.699, 3292.384, 3380.365, 2269.825, 515.0248, 4.337821, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  431.9473, 396.6402, 222.4012, 114.462, 25.37888, 7.691118, 6.677791, 
    7.348661, 3.157577, 0.984972, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3024256, 
    0.2389092, 0.1394803, 0.00746349, 0, 70.57438, 149.7564, 0, 80.11617, 
    0.0417327, 0, 0, 0, 0, 0, 0, 0, 0.01057512, 27.73273, 266.8832, 915.6628, 
    1100.12, 1117.166, 1315.549, 1758.784, 2041.483, 1431.61, 474.8531, 
    232.1502, 208.0247, 196.3371, 166.9769, 139.262, 189.603, 539.9, 
    636.6401, 1134.973, 2116.188, 3255.661, 3725.555, 3525.62, 2041.445, 
    414.1652, 93.96832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  441.435, 319.8361, 136.8747, 29.58521, 4.141918, 2.825089, 0.08903898, 
    0.08046266, 0.2208437, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3990609, 
    0.3265876, 0.0633444, 0.05431467, 84.71734, 149.596, 0, 0.04963135, 0, 0, 
    0, 0, 0, 0, 0, 27.05583, 59.55542, 2.632703, 383.2401, 1071.188, 
    1466.155, 1676.46, 1735.292, 1635.764, 1205.279, 587.2426, 204.6946, 
    192.8305, 201.6285, 192.1485, 173.3057, 135.0386, 115.5985, 154.6932, 
    207.6518, 252.7319, 408.4037, 1234.129, 2512.059, 3625.666, 3840.744, 
    2953.312, 1398.119, 200.1961, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  298.2758, 155.1034, 25.55248, 4.920603, 0.003125044, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1279996, 0.02609903, 0.3170911, 0, 23.67887, 
    68.64729, 35.86671, 72.66331, 0, 0, 0, 0, 0, 0, 27.26858, 361.5938, 
    62.6906, 207.8889, 270.3431, 466.9674, 991.8314, 1723.766, 1665.32, 
    1134.25, 697.3764, 239.1669, 204.7155, 192.0341, 177.9332, 167.6514, 
    147.1711, 124.0248, 116.1455, 138.7632, 205.803, 202.1669, 218.9659, 
    445.2673, 918.5952, 2052.283, 3110.208, 3814.63, 3245.299, 1978.916, 
    128.154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.621783, 0, 0, 1.331606, 2.106077,
  156.3812, 18.64756, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.02620244, 0.1723592, 0.6139864, 0.7052164, 39.91206, 73.66648, 
    34.73109, 0, 0, 0, 0, 0, 0, 103.6746, 970.1916, 637.6611, 308.0594, 
    768.11, 1294.207, 1777.075, 1670.896, 1144.713, 449.2721, 228.4367, 
    250.4818, 226.3325, 198.0396, 169.848, 146.4091, 131.5473, 124.774, 
    133.6427, 162.3437, 232.3307, 229.8633, 231.2848, 277.8121, 478.211, 
    827.6024, 1960.805, 3358.45, 4059.359, 3432.779, 1310.91, 0.5703501, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.00629, 
    172.8352, 183.9977, 46.27448, 129.1229, 178.4515, 97.62695,
  36.70903, 1.210476, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.226078, 0.04288947, 3.178066, 257.9394, 343.0803, 13.00084, 0, 
    0, 0, 0, 0, 2.137605, 96.99342, 646.0239, 147.4564, 527.7556, 1280.455, 
    1827.782, 1949.41, 1110.227, 192.4001, 183.5117, 228.3509, 244.9112, 
    227.8943, 192.5254, 159.7048, 137.4386, 124.2721, 122.957, 142.0076, 
    164.3923, 198.738, 229.3472, 259.537, 313.7084, 313.5366, 602.6287, 
    1546.649, 3188.223, 4339.325, 4235.496, 2657.681, 348.9787, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.4312, 110.2107, 
    133.0185, 292.7062, 324.6068, 298.3218, 359.0092, 476.8519, 554.6548,
  1.995229, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4212663, 0.04588909, 11.18899, 517.642, 542.4244, 51.31382, 0, 0, 0, 0, 
    0, 43.47145, 14.86237, 90.16446, 49.90094, 852.6797, 695.9244, 698.5693, 
    469.248, 149.1092, 136.4317, 196.3584, 211.3587, 231.4343, 214.1757, 
    171.0396, 141.9184, 127.4874, 119.4414, 115.9838, 130.7626, 159.6196, 
    192.4039, 226.2965, 268.5108, 312.2362, 358.5796, 389.9218, 1083.607, 
    2472.518, 4258.277, 4571.348, 3741.117, 2121.892, 269.5249, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.388186, 133.4869, 148.3846, 211.8387, 382.2953, 
    257.1787, 180.7228, 149.7092, 212.2956, 459.678, 761.8045, 1055.912, 
    1120.853, 1110.582, 1166.25, 1085.751, 1108.78,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001913318, 33.17125, 520.3718, 399.8852, 0, 0, 0, 0, 0, 0, 0.8113799, 
    95.28371, 460.3841, 937.3494, 915.1066, 445.8253, 106.3576, 103.3282, 
    112.4795, 164.6748, 183.3819, 200.0266, 220.7052, 195.8168, 166.651, 
    121.4309, 123.9416, 113.4673, 102.3118, 125.9921, 156.5412, 179.7962, 
    206.3467, 238.4389, 260.7508, 315.1216, 328.1903, 360.6142, 1509.248, 
    3565.005, 4402.538, 4396.66, 3602.803, 2091.149, 261.0787, 82.22005, 
    0.2868135, 0, 0.5076911, 60.36261, 183.4623, 519.5708, 450.9728, 
    353.2507, 488.7053, 617.8168, 1421.896, 2045.6, 2299.798, 2328.442, 
    2164.863, 1835.325, 1553.868, 1649.168, 1826.316, 1985.27, 1961.338, 
    1556.79, 1371.403, 1288.084, 1040.601, 1072.717,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.771062, 165.8212, 28.28846, 0, 0, 0, 0, 0, 0.1610673, 17.69787, 
    260.4066, 714.0234, 586.6948, 462.326, 79.98116, 88.8905, 101.472, 
    127.5234, 151.2906, 172.9191, 187.4914, 183.702, 173.0886, 139.7318, 
    124.8896, 118.3931, 105.5773, 109.4129, 131.1672, 156.9932, 163.0083, 
    184.8383, 204.416, 225.2426, 266.9706, 316.145, 224.5979, 381.9278, 
    2492.509, 3806.261, 4259.841, 4400.584, 3759.828, 2950.103, 2123.126, 
    1457.011, 1071.604, 1158.814, 1261.4, 1360.847, 1651.959, 2091.039, 
    2134.101, 2298.518, 2832.512, 3516.553, 3862.269, 3539.123, 3228.904, 
    3070.49, 3133.28, 3088.744, 2907.435, 2507.032, 2134.26, 1858.328, 
    1274.926, 962.0797, 842.9384, 710.9687, 939.0226,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 51.69876, 6.425387, 0, 0, 0, 0, 0, 0, 2.873953, 169.8395, 449.1624, 
    300.1902, 62.32654, 69.31486, 78.20786, 85.0916, 97.69564, 127.4337, 
    145.2199, 162.7987, 148.36, 126.3364, 126.9805, 112.7666, 113.0274, 
    97.65716, 107.4775, 138.243, 148.1546, 151.6598, 170.6716, 190.0256, 
    201.0505, 226.6755, 261.319, 232.2254, 219.3973, 932.7808, 2511.412, 
    3070.967, 3937.193, 4288.645, 4117.858, 3970.56, 3654.04, 3348.081, 
    3098.408, 2970.42, 2560.729, 2923.75, 3655.134, 3966.941, 4254.809, 
    4391.425, 4123.873, 3285.485, 2428.365, 1895.18, 1763.043, 1610.22, 
    1446.99, 1407.953, 1387.499, 1476.249, 1487.882, 1047.58, 652.7329, 
    528.4442, 542.4118, 917.0056,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.3669669, 0.3634669, 0, 0, 0, 0, 0, 0, 0.6933007, 13.2217, 484.2191, 
    144.2932, 49.07107, 47.2271, 55.1874, 111.1454, 210.9041, 104.5796, 
    116.9778, 131.3689, 115.879, 101.3334, 98.76527, 97.77927, 91.92683, 
    82.82296, 102.0775, 115.0132, 128.6879, 136.6141, 155.6852, 166.7384, 
    172.6179, 192.5376, 207.4939, 206.3573, 175.2231, 245.1321, 792.022, 
    1577.401, 2693.881, 3723.349, 4046.354, 3911.702, 3846.095, 3873.51, 
    4067.074, 4060.027, 3885.769, 3648.284, 4000.79, 4255.121, 4298.765, 
    3941.536, 2986.297, 2167.081, 1555.988, 1086.933, 981.1671, 671.5908, 
    517.9108, 560.5896, 604.6505, 737.5284, 838.4316, 663.5747, 487.8661, 
    405.7701, 432.4994, 598.6184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 87.07624, 9.664433, 0, 0, 0, 0, 0, 0, 0.1396964, 165.1147, 498.7843, 
    209.5764, 50.07817, 49.66368, 196.0763, 442.8151, 358.6526, 227.8948, 
    104.9866, 105.646, 125.2638, 109.2299, 82.44156, 78.38992, 73.12806, 
    72.46248, 85.68304, 100.9489, 111.212, 121.0391, 131.6541, 139.9958, 
    153.3166, 166.8747, 176.9339, 177.9256, 166.0943, 164.8257, 217.7268, 
    390.218, 1575.724, 3050.704, 3828.212, 3839.21, 3919.247, 3790.678, 
    3970.27, 4419.288, 4398.239, 4177.742, 4184.263, 4184.499, 4041.16, 
    3409.468, 2121.299, 1508.151, 989.2469, 766.4855, 749.4873, 491.5999, 
    500.2154, 587.9318, 432.9168, 407.4583, 403.593, 373.3047, 314.6314, 
    310.2964, 287.6699, 288.7629,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 137.5109, 1.268968, 0, 0, 0, 0, 0, 0, 0.1147682, 82.57735, 311.5683, 
    151.4449, 78.04676, 128.0494, 376.5229, 522.9591, 427.1115, 256.4601, 
    112.6585, 142.7851, 266.511, 196.9078, 88.25249, 66.20465, 58.85111, 
    66.82548, 83.11908, 91.31876, 101.4318, 105.2445, 110.9949, 121.9766, 
    145.8439, 152.8409, 158.7673, 160.5151, 158.0549, 151.2477, 147.5351, 
    168.9152, 567.9518, 1848.487, 3247.352, 3623.287, 3933.537, 4026.396, 
    3815.863, 3989.005, 4117.667, 4075.111, 3740.598, 3347.181, 3151.984, 
    2783.441, 1733.658, 1189.891, 689.3563, 352.485, 479.9682, 518.3051, 
    654.5156, 843.5643, 637.5115, 436.4144, 356.3743, 315.6976, 287.2369, 
    264.154, 245.379, 203.1721,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0005155665, 0.00535053, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5.954806, 0.008552877, 0, 0, 0, 0, 0, 0, 0, 
    1.392343, 147.5822, 117.1248, 79.08617, 161.021, 478.1805, 672.9123, 
    747.8989, 659.3046, 435.462, 300.6021, 411.5335, 261.7856, 93.77441, 
    56.53286, 59.12653, 61.15051, 76.3445, 85.60712, 87.65303, 86.02962, 
    90.52665, 104.9385, 125.5316, 141.8028, 161.3927, 151.9469, 148.933, 
    141.536, 144.3197, 149.6154, 172.0073, 623.9898, 1684.723, 2641.521, 
    3090.655, 3319.659, 3217.01, 3316.014, 3452.869, 3067.782, 2450.786, 
    1764.937, 1428.371, 1315.265, 759.3845, 608.1971, 375.0185, 229.107, 
    391.8174, 639.2117, 819.7453, 915.3849, 607.8117, 379.9553, 305.7845, 
    306.8441, 298.1168, 286.4967, 240.3828, 184.6151,
  0, 0, 0, 0, 0, 0, 0, 0, 0.121945, 0.03938331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.3118506, 3.291815, 0.01598853, 0, 0, 0, 0, 0, 0.1340173, 
    4.044582, 143.5697, 233.638, 191.9344, 118.6989, 147.4646, 285.2692, 
    535.5562, 720.2246, 908.1365, 672.2578, 505.0814, 365.3874, 130.3261, 
    44.65852, 61.89712, 58.099, 59.19082, 61.83461, 73.12101, 69.1452, 
    71.91867, 79.77286, 88.05507, 108.2875, 147.0296, 195.7139, 207.4643, 
    157.7728, 145.7407, 144.7948, 163.3843, 160.5329, 192.4493, 810.9302, 
    1566.056, 2149.559, 2256.098, 2102.709, 1810.442, 1541.477, 1113.111, 
    754.5137, 622.1283, 649.4427, 513.0068, 210.115, 259.1717, 228.6151, 
    216.1971, 473.4304, 783.3362, 789.3256, 686.4561, 419.5589, 249.4682, 
    205.099, 202.2573, 216.5917, 217.1671, 199.7617, 132.155,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.005494107, 0.4346767, 0, 0, 0, 0, 0, 0, 0, 9.391527, 298.571, 237.2993, 
    140.6926, 155.2257, 256.6727, 406.4414, 433.8806, 600.3461, 683.2579, 
    620.795, 483.5708, 265.2493, 69.42221, 44.01501, 51.81279, 60.87005, 
    53.39784, 52.44471, 56.40654, 59.58292, 67.88076, 74.34882, 81.33792, 
    95.65347, 148.0806, 236.6955, 255.9585, 205.559, 151.0034, 159.6844, 
    176.646, 199.4624, 204.3659, 270.1312, 848.1915, 1003.153, 1148.617, 
    1003.102, 887.6286, 594.8246, 321.8112, 230.0089, 347.2778, 260.032, 
    255.0762, 190.1423, 159.5509, 136.5862, 182.9312, 271.9562, 310.1284, 
    283.9276, 277.2419, 213.3407, 155.9381, 136.6259, 129.9663, 124.8657, 
    144.5141, 150.6962, 106.1049,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2010026, 5.480222, 1.905644, 0, 0, 0, 0, 0, 0, 10.41574, 79.70645, 
    33.17719, 101.7773, 211.8761, 328.2486, 519.1068, 687.5656, 568.6201, 
    426.9638, 407.4171, 258.6449, 133.8155, 46.44923, 40.82528, 43.58858, 
    52.29549, 51.97647, 43.10914, 47.15418, 57.30152, 61.27217, 67.14295, 
    78.3484, 97.84009, 141.1024, 209.3585, 245.7221, 223.8985, 178.6274, 
    164.8928, 205.0671, 272.722, 329.3512, 281.3043, 329.6042, 396.7708, 
    453.139, 536.9029, 418.7523, 345.6891, 235.4872, 214.9491, 197.1605, 
    217.0889, 210.202, 187.8262, 155.8819, 114.6811, 108.0696, 103.5813, 
    75.537, 103.2833, 131.8954, 130.8562, 121.067, 118.0025, 105.5169, 
    96.54052, 119.8245, 176.6302, 195.5793,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.086443, 9.708963, 25.8066, 0, 0, 0, 0.6762983, 7.368328, 15.26273, 
    7.240432, 15.79535, 109.3353, 221.0537, 269.0515, 704.3265, 939.6818, 
    701.0948, 330.6563, 190.7539, 178.3714, 105.7215, 59.61247, 39.14966, 
    45.20544, 46.21466, 48.67001, 35.86091, 46.08049, 52.98456, 62.92745, 
    69.35141, 85.43824, 110.8834, 142.6441, 180.2906, 238.7265, 252.6595, 
    239.7324, 184.5832, 228.8213, 276.7168, 392.7193, 388.6469, 296.1601, 
    280.3641, 341.4388, 353.615, 317.2159, 244.4351, 223.8407, 201.6992, 
    183.6967, 176.9333, 172.614, 165.7017, 145.3332, 110.9088, 80.85966, 
    70.93066, 76.48385, 91.80798, 97.15785, 91.67457, 100.7875, 107.6938, 
    96.9532, 86.08794, 101.3551, 185.22, 281.0552,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.485921, 26.4163, 34.1476, 13.50462, 14.0831, 0.4166287, 2.192102, 
    29.53002, 14.33252, 3.286679, 52.2133, 156.3645, 257.6373, 649.4648, 
    1054.655, 614.7567, 162.2067, 99.85813, 116.9508, 77.15819, 48.32669, 
    64.66377, 56.2935, 65.67332, 46.97363, 33.90272, 37.93755, 51.28942, 
    58.10233, 78.93856, 106.3503, 116.9305, 149.4504, 180.898, 213.7403, 
    292.1611, 291.1207, 281.1519, 252.0287, 285.7556, 316.2794, 374.6313, 
    325.8148, 322.2468, 325.9581, 276.3282, 228.0858, 195.2241, 187.3171, 
    175.7014, 163.5601, 151.0618, 141.3108, 129.977, 114.84, 86.42167, 
    68.05943, 63.20282, 64.60545, 60.11647, 42.99261, 50.01132, 55.99592, 
    74.10268, 81.50942, 73.58952, 83.45282, 127.7083, 226.8334,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.984597, 0.01858864, 0, 0.0009470581, 16.01784, 
    87.35822, 173.5935, 488.2748, 759.5725, 523.7241, 141.7197, 113.1382, 
    159.5228, 147.7596, 115.4366, 107.1132, 102.7932, 85.72213, 66.42902, 
    30.98574, 37.11678, 45.43555, 64.23547, 99.53561, 129.9766, 138.2153, 
    142.8759, 176.7178, 267.0287, 349.3065, 417.0574, 373.9982, 391.8378, 
    306.8354, 254.5319, 312.5648, 296.5179, 377.6109, 330.0472, 242.8435, 
    164.2536, 149.3302, 147.9863, 144.5899, 139.069, 133.0572, 122.3601, 
    110.4266, 95.19322, 77.43336, 63.58871, 58.07784, 51.05425, 36.38617, 
    36.80247, 46.6338, 42.84441, 35.56261, 47.46378, 56.36189, 58.939, 
    105.9327, 189.9787,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.923116, 0, 0, 0, 0, 0, 6.078897, 54.77836, 77.55535, 
    204.2334, 410.9161, 330.8391, 185.1925, 194.0988, 249.267, 253.3829, 
    177.0466, 158.8476, 113.1643, 101.53, 68.00449, 31.76886, 36.63785, 
    58.77195, 90.80497, 133.0862, 161.9473, 164.7115, 165.2141, 201.0824, 
    279.0718, 359.1356, 398.5262, 459.7346, 501.9608, 511.8822, 352.2849, 
    246.1968, 246.5588, 279.2735, 323.1726, 191.8587, 143.4464, 112.1324, 
    117.9595, 116.5617, 114.9787, 113.5484, 107.3903, 97.09441, 84.3097, 
    70.09772, 57.50354, 51.82816, 43.33216, 40.77794, 45.42603, 66.79871, 
    45.82823, 21.87241, 20.00079, 29.68418, 34.1625, 55.23173, 131.1202,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007114115, 12.30466, 48.17017, 
    51.3419, 136.4395, 140.1926, 152.5834, 214.4402, 290.774, 334.6097, 
    242.1319, 179.8538, 138.1877, 94.74007, 53.06939, 31.48326, 46.89961, 
    89.87615, 131.2574, 140.4565, 168.6543, 171.5402, 207.168, 234.0502, 
    297.8369, 300.6861, 321.7401, 399.447, 557.8159, 602.8211, 392.1693, 
    231.2913, 117.9363, 190.2211, 228.4644, 181.8213, 100.4968, 90.92713, 
    91.9957, 95.57886, 98.97549, 93.66434, 91.03915, 82.98544, 72.89633, 
    60.49364, 58.69539, 60.83919, 60.2387, 64.67129, 64.97378, 60.37475, 
    50.22374, 26.93556, 10.59541, 21.63067, 16.65605, 21.7373, 41.34349,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.366938, 28.12142, 64.29294, 
    128.7759, 176.1391, 224.7735, 297.6988, 326.8529, 254.3473, 185.0925, 
    128.5998, 87.42819, 38.13975, 29.44325, 68.62458, 118.0892, 143.8512, 
    173.974, 164.9058, 204.4256, 210.1949, 267.1867, 300.9321, 309.5306, 
    297.9662, 355.8887, 461.3635, 509.2478, 310.7938, 206.6006, 123.8932, 
    125.1484, 178.9654, 129.2888, 94.40868, 92.13621, 118.3059, 139.3436, 
    102.2285, 87.8205, 78.24416, 72.41794, 72.99378, 69.93626, 64.41702, 
    66.0837, 67.51834, 70.63937, 64.17177, 65.43086, 61.57732, 57.59845, 
    48.39719, 66.22498, 19.65588, 7.979198, 7.954746,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1979136, 16.10868, 94.42965, 
    187.4814, 245.3877, 271.5805, 257.391, 297.2609, 210.7862, 164.771, 
    95.62947, 56.90887, 40.72773, 52.8884, 92.41105, 126.1473, 166.0383, 
    207.8445, 272.0114, 271.0105, 294.9529, 248.3746, 307.0643, 316.8501, 
    327.4612, 325.9547, 386.9184, 403.7983, 311.1118, 240.8184, 164.2083, 
    103.1077, 117.4106, 99.13666, 106.3574, 154.6648, 260.3508, 285.6964, 
    234.8461, 154.5512, 112.9279, 100.7134, 123.8555, 127.3378, 90.11683, 
    76.42348, 68.03311, 66.51344, 75.3875, 112.4858, 142.2936, 124.5137, 
    93.33791, 99.31126, 54.70262, 4.06266, 0.262289,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04155033, 10.73219, 79.11258, 
    190.445, 274.9487, 342.6148, 355.8712, 312.3603, 292.6754, 221.7762, 
    115.474, 47.77611, 50.80471, 84.23752, 95.56871, 148.4016, 177.4802, 
    241.8285, 273.5516, 339.5761, 337.356, 326.2194, 277.1494, 336.4698, 
    352.6033, 363.4337, 382.938, 416.9631, 325.3823, 303.8384, 203.988, 
    116.0254, 110.5155, 121.6094, 106.5421, 137.3756, 210.812, 317.8851, 
    344.7708, 323.2015, 252.112, 193.5985, 213.3652, 191.4196, 156.1301, 
    106.2765, 104.4049, 72.89532, 100.3581, 157.0007, 215.9135, 191.733, 
    119.1055, 115.4301, 99.49779, 31.93542, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.542466, 22.26523, 77.77408, 
    140.4331, 240.0608, 343.6068, 376.1221, 378.217, 372.9897, 356.2578, 
    217.9453, 48.16224, 56.58264, 94.03797, 155.6086, 206.1189, 244.8234, 
    262.5258, 267.4071, 294.3894, 384.4132, 383.2951, 330.3748, 318.6039, 
    351.7903, 366.8914, 400.56, 447.5571, 438.7595, 508.2295, 383.2372, 
    246.7716, 200.7712, 148.0255, 184.6252, 228.8072, 293.0768, 384.8521, 
    451.6723, 470.1341, 383.5, 297.7384, 261.2184, 257.7826, 233.8021, 
    230.1151, 168.3038, 140.5308, 159.7929, 141.3796, 184.5563, 169.6956, 
    127.2488, 153.812, 157.5335, 129.1637, 8.482048 ;
}
