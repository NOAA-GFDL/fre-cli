netcdf \00010101.atmos_daily.tile3.pv350K {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;


 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  2.017718e-08, 1.976381e-08, 1.961709e-08, 1.986073e-08, 2.047343e-08, 
    2.118852e-08, 2.208785e-08, 2.274241e-08, 2.334492e-08, 2.370841e-08, 
    2.389475e-08, 2.402058e-08, 2.377232e-08, 2.368855e-08, 2.355447e-08,
  2.190678e-08, 2.139531e-08, 2.09069e-08, 2.059836e-08, 2.078039e-08, 
    2.189722e-08, 2.27305e-08, 2.347991e-08, 2.374091e-08, 2.397768e-08, 
    2.402963e-08, 2.406372e-08, 2.403866e-08, 2.372944e-08, 2.331324e-08,
  2.329143e-08, 2.251149e-08, 2.131385e-08, 2.068825e-08, 2.123963e-08, 
    2.275906e-08, 2.409936e-08, 2.450796e-08, 2.439861e-08, 2.420946e-08, 
    2.398099e-08, 2.382929e-08, 2.370662e-08, 2.359628e-08, 2.340611e-08,
  2.394707e-08, 2.312124e-08, 2.177468e-08, 2.116737e-08, 2.172701e-08, 
    2.366735e-08, 2.489848e-08, 2.431501e-08, 2.403957e-08, 2.387475e-08, 
    2.358344e-08, 2.347759e-08, 2.339066e-08, 2.32351e-08, 2.337963e-08,
  2.418862e-08, 2.364578e-08, 2.251291e-08, 2.188292e-08, 2.225765e-08, 
    2.372152e-08, 2.429897e-08, 2.440821e-08, 2.369208e-08, 2.190219e-08, 
    2.174546e-08, 2.265097e-08, 2.287587e-08, 2.296371e-08, 2.300941e-08,
  2.35327e-08, 2.394826e-08, 2.326776e-08, 2.257785e-08, 2.251337e-08, 
    2.327823e-08, 2.320986e-08, 2.246457e-08, 2.153551e-08, 2.072541e-08, 
    2.117874e-08, 2.199677e-08, 2.239311e-08, 2.269771e-08, 2.290329e-08,
  2.262755e-08, 2.352544e-08, 2.380145e-08, 2.336093e-08, 2.318407e-08, 
    2.304087e-08, 2.244303e-08, 2.184942e-08, 2.115291e-08, 2.083576e-08, 
    2.109996e-08, 2.18049e-08, 2.221965e-08, 2.258342e-08, 2.249154e-08,
  2.160614e-08, 2.287316e-08, 2.378406e-08, 2.379613e-08, 2.368718e-08, 
    2.362781e-08, 2.288075e-08, 2.153551e-08, 2.109016e-08, 2.101563e-08, 
    2.12975e-08, 2.185383e-08, 2.233667e-08, 2.218719e-08, 2.200407e-08,
  2.075658e-08, 2.202219e-08, 2.338382e-08, 2.391924e-08, 2.402308e-08, 
    2.414219e-08, 2.39554e-08, 2.273239e-08, 2.134076e-08, 2.104014e-08, 
    2.172136e-08, 2.173235e-08, 2.200942e-08, 2.167903e-08, 2.129734e-08,
  2.117451e-08, 2.169673e-08, 2.262507e-08, 2.371684e-08, 2.401337e-08, 
    2.419306e-08, 2.482425e-08, 2.472738e-08, 2.39908e-08, 2.346141e-08, 
    2.275862e-08, 2.199752e-08, 2.180575e-08, 2.136235e-08, 2.148007e-08,
  2.403501e-08, 2.337882e-08, 2.266398e-08, 2.127729e-08, 1.951859e-08, 
    2.036092e-08, 2.306692e-08, 2.361765e-08, 2.377142e-08, 2.35035e-08, 
    2.366152e-08, 2.375429e-08, 2.425484e-08, 2.384802e-08, 2.380567e-08,
  2.384711e-08, 2.333777e-08, 2.276363e-08, 2.243803e-08, 2.090667e-08, 
    2.033364e-08, 2.145131e-08, 2.28213e-08, 2.322077e-08, 2.311993e-08, 
    2.328802e-08, 2.333665e-08, 2.356926e-08, 2.345454e-08, 2.355723e-08,
  2.419242e-08, 2.357465e-08, 2.326587e-08, 2.242611e-08, 2.165548e-08, 
    2.070542e-08, 2.117653e-08, 2.209061e-08, 2.260989e-08, 2.265834e-08, 
    2.302478e-08, 2.311866e-08, 2.32128e-08, 2.339601e-08, 2.371418e-08,
  2.438417e-08, 2.401683e-08, 2.39114e-08, 2.334487e-08, 2.264205e-08, 
    2.193884e-08, 2.162726e-08, 2.218293e-08, 2.321621e-08, 2.321116e-08, 
    2.335677e-08, 2.340308e-08, 2.355227e-08, 2.367302e-08, 2.444887e-08,
  2.459692e-08, 2.428617e-08, 2.434583e-08, 2.393395e-08, 2.373014e-08, 
    2.305892e-08, 2.270703e-08, 2.259691e-08, 2.325375e-08, 2.300309e-08, 
    2.358136e-08, 2.369919e-08, 2.387315e-08, 2.374584e-08, 2.423142e-08,
  2.444149e-08, 2.422463e-08, 2.422239e-08, 2.369573e-08, 2.315899e-08, 
    2.272403e-08, 2.23625e-08, 2.216222e-08, 2.285307e-08, 2.305049e-08, 
    2.328946e-08, 2.339169e-08, 2.377731e-08, 2.371738e-08, 2.410993e-08,
  2.437455e-08, 2.412435e-08, 2.394439e-08, 2.332123e-08, 2.246552e-08, 
    2.182723e-08, 2.179253e-08, 2.197686e-08, 2.226782e-08, 2.244078e-08, 
    2.275749e-08, 2.304007e-08, 2.348464e-08, 2.361435e-08, 2.398894e-08,
  2.401193e-08, 2.411686e-08, 2.380542e-08, 2.323109e-08, 2.22097e-08, 
    2.147238e-08, 2.117551e-08, 2.167377e-08, 2.202874e-08, 2.224935e-08, 
    2.253875e-08, 2.270845e-08, 2.301436e-08, 2.335512e-08, 2.377731e-08,
  2.382161e-08, 2.396762e-08, 2.385737e-08, 2.356454e-08, 2.282571e-08, 
    2.200727e-08, 2.13954e-08, 2.142302e-08, 2.170582e-08, 2.192785e-08, 
    2.237131e-08, 2.264211e-08, 2.291727e-08, 2.314198e-08, 2.338239e-08,
  2.371851e-08, 2.391914e-08, 2.375707e-08, 2.339014e-08, 2.298749e-08, 
    2.246359e-08, 2.202242e-08, 2.167566e-08, 2.167909e-08, 2.207242e-08, 
    2.24127e-08, 2.262316e-08, 2.274083e-08, 2.291827e-08, 2.317872e-08,
  2.464277e-08, 2.456013e-08, 2.343494e-08, 2.3289e-08, 2.120369e-08, 
    2.073402e-08, 2.283465e-08, 2.372655e-08, 2.374169e-08, 2.370829e-08, 
    2.330046e-08, 2.313745e-08, 2.292166e-08, 2.170394e-08, 2.152543e-08,
  2.457843e-08, 2.460217e-08, 2.381676e-08, 2.295156e-08, 2.066516e-08, 
    2.086715e-08, 2.32789e-08, 2.393812e-08, 2.381476e-08, 2.354573e-08, 
    2.332725e-08, 2.329241e-08, 2.221556e-08, 2.057118e-08, 2.319158e-08,
  2.419801e-08, 2.427405e-08, 2.385238e-08, 2.232604e-08, 2.100653e-08, 
    2.135724e-08, 2.392965e-08, 2.396387e-08, 2.370434e-08, 2.353405e-08, 
    2.305944e-08, 2.261782e-08, 2.11423e-08, 2.19321e-08, 2.408206e-08,
  2.365366e-08, 2.375765e-08, 2.349691e-08, 2.225969e-08, 2.118682e-08, 
    2.18011e-08, 2.389753e-08, 2.430848e-08, 2.365599e-08, 2.33174e-08, 
    2.310525e-08, 2.261861e-08, 2.211235e-08, 2.26709e-08, 2.447075e-08,
  2.282039e-08, 2.304541e-08, 2.321925e-08, 2.236626e-08, 2.168948e-08, 
    2.224434e-08, 2.357432e-08, 2.402338e-08, 2.375861e-08, 2.350148e-08, 
    2.298851e-08, 2.288642e-08, 2.2921e-08, 2.44913e-08, 2.506973e-08,
  2.229867e-08, 2.223508e-08, 2.25287e-08, 2.226308e-08, 2.21247e-08, 
    2.285208e-08, 2.362244e-08, 2.365081e-08, 2.320325e-08, 2.326869e-08, 
    2.30874e-08, 2.332149e-08, 2.371222e-08, 2.38324e-08, 2.392177e-08,
  2.20876e-08, 2.203843e-08, 2.205344e-08, 2.214171e-08, 2.254606e-08, 
    2.317647e-08, 2.336018e-08, 2.343914e-08, 2.318103e-08, 2.314478e-08, 
    2.275098e-08, 2.26097e-08, 2.319702e-08, 2.330828e-08, 2.4485e-08,
  2.211049e-08, 2.203887e-08, 2.197497e-08, 2.22096e-08, 2.276494e-08, 
    2.322855e-08, 2.330005e-08, 2.316272e-08, 2.286553e-08, 2.303445e-08, 
    2.284684e-08, 2.257292e-08, 2.251021e-08, 2.340474e-08, 2.452223e-08,
  2.232416e-08, 2.206122e-08, 2.212531e-08, 2.225496e-08, 2.26516e-08, 
    2.305115e-08, 2.321536e-08, 2.313656e-08, 2.291448e-08, 2.269719e-08, 
    2.184748e-08, 2.180379e-08, 2.262302e-08, 2.362868e-08, 2.367004e-08,
  2.228698e-08, 2.22388e-08, 2.200685e-08, 2.217627e-08, 2.243457e-08, 
    2.280544e-08, 2.311099e-08, 2.302383e-08, 2.296766e-08, 2.286314e-08, 
    2.252872e-08, 2.239044e-08, 2.298069e-08, 2.330167e-08, 2.322462e-08,
  2.309548e-08, 2.426678e-08, 2.389979e-08, 2.399121e-08, 2.340163e-08, 
    2.252829e-08, 2.223612e-08, 2.21916e-08, 2.214398e-08, 2.233669e-08, 
    2.286416e-08, 2.355194e-08, 2.35802e-08, 2.317278e-08, 2.391998e-08,
  2.333153e-08, 2.429645e-08, 2.384469e-08, 2.316277e-08, 2.191234e-08, 
    2.167254e-08, 2.207215e-08, 2.253594e-08, 2.262557e-08, 2.279396e-08, 
    2.353036e-08, 2.357849e-08, 2.282489e-08, 2.321014e-08, 2.561947e-08,
  2.376228e-08, 2.390348e-08, 2.291384e-08, 2.168622e-08, 2.145776e-08, 
    2.212733e-08, 2.2866e-08, 2.28046e-08, 2.290791e-08, 2.341657e-08, 
    2.349635e-08, 2.269409e-08, 2.296634e-08, 2.484544e-08, 2.594786e-08,
  2.372229e-08, 2.297984e-08, 2.18297e-08, 2.14225e-08, 2.176547e-08, 
    2.262018e-08, 2.314271e-08, 2.348566e-08, 2.341645e-08, 2.324324e-08, 
    2.28935e-08, 2.277675e-08, 2.425853e-08, 2.586016e-08, 2.507865e-08,
  2.326481e-08, 2.220471e-08, 2.156697e-08, 2.163325e-08, 2.274632e-08, 
    2.350211e-08, 2.344883e-08, 2.319312e-08, 2.289919e-08, 2.274053e-08, 
    2.295643e-08, 2.378175e-08, 2.576742e-08, 2.542277e-08, 2.390215e-08,
  2.265797e-08, 2.187628e-08, 2.163026e-08, 2.240899e-08, 2.340832e-08, 
    2.361187e-08, 2.28308e-08, 2.190974e-08, 2.237187e-08, 2.406978e-08, 
    2.407709e-08, 2.536832e-08, 2.573769e-08, 2.413863e-08, 2.314038e-08,
  2.238059e-08, 2.189088e-08, 2.214161e-08, 2.318383e-08, 2.378846e-08, 
    2.373754e-08, 2.303679e-08, 2.275699e-08, 2.32485e-08, 2.407651e-08, 
    2.487254e-08, 2.569925e-08, 2.449842e-08, 2.338548e-08, 2.319493e-08,
  2.224953e-08, 2.212169e-08, 2.2814e-08, 2.373076e-08, 2.376121e-08, 
    2.354854e-08, 2.262805e-08, 2.257564e-08, 2.312466e-08, 2.433778e-08, 
    2.527714e-08, 2.477034e-08, 2.381838e-08, 2.356355e-08, 2.334968e-08,
  2.238007e-08, 2.271885e-08, 2.350736e-08, 2.401384e-08, 2.3698e-08, 
    2.326265e-08, 2.268108e-08, 2.317574e-08, 2.372065e-08, 2.459902e-08, 
    2.464427e-08, 2.395344e-08, 2.381023e-08, 2.333573e-08, 2.274043e-08,
  2.278156e-08, 2.332094e-08, 2.383139e-08, 2.387423e-08, 2.308351e-08, 
    2.27374e-08, 2.288771e-08, 2.372944e-08, 2.391034e-08, 2.462064e-08, 
    2.385161e-08, 2.362795e-08, 2.351588e-08, 2.29181e-08, 2.310598e-08,
  2.36226e-08, 2.358721e-08, 2.375519e-08, 2.439376e-08, 2.423621e-08, 
    2.351133e-08, 2.284033e-08, 2.215243e-08, 2.120684e-08, 2.174007e-08, 
    2.252502e-08, 2.2904e-08, 2.361845e-08, 2.440523e-08, 2.415187e-08,
  2.326723e-08, 2.340951e-08, 2.394855e-08, 2.439306e-08, 2.376222e-08, 
    2.304406e-08, 2.253362e-08, 2.187308e-08, 2.16449e-08, 2.191564e-08, 
    2.273758e-08, 2.339289e-08, 2.38047e-08, 2.392024e-08, 2.405213e-08,
  2.318077e-08, 2.364307e-08, 2.399595e-08, 2.381557e-08, 2.321044e-08, 
    2.282313e-08, 2.221747e-08, 2.136933e-08, 2.124265e-08, 2.211746e-08, 
    2.342626e-08, 2.376327e-08, 2.397623e-08, 2.398294e-08, 2.410878e-08,
  2.329283e-08, 2.362956e-08, 2.349237e-08, 2.313907e-08, 2.262001e-08, 
    2.232494e-08, 2.198508e-08, 2.165974e-08, 2.219079e-08, 2.284931e-08, 
    2.384413e-08, 2.403652e-08, 2.411955e-08, 2.427261e-08, 2.399191e-08,
  2.329048e-08, 2.330922e-08, 2.291384e-08, 2.249723e-08, 2.249852e-08, 
    2.22262e-08, 2.180906e-08, 2.192214e-08, 2.211409e-08, 2.134437e-08, 
    2.406793e-08, 2.415063e-08, 2.440137e-08, 2.430525e-08, 2.397586e-08,
  2.329095e-08, 2.263031e-08, 2.231767e-08, 2.24837e-08, 2.237139e-08, 
    2.186341e-08, 2.028837e-08, 1.730256e-08, 1.837613e-08, 2.565464e-08, 
    2.77516e-08, 2.458084e-08, 2.459695e-08, 2.4393e-08, 2.400909e-08,
  2.259444e-08, 2.224841e-08, 2.223805e-08, 2.240864e-08, 2.209938e-08, 
    2.091965e-08, 1.848722e-08, 1.823328e-08, 2.425497e-08, 3.008197e-08, 
    2.651142e-08, 2.452563e-08, 2.466397e-08, 2.449682e-08, 2.404029e-08,
  2.247932e-08, 2.203074e-08, 2.231087e-08, 2.251304e-08, 2.172853e-08, 
    1.946789e-08, 1.855914e-08, 2.232642e-08, 2.846934e-08, 2.886962e-08, 
    2.505063e-08, 2.447735e-08, 2.468282e-08, 2.458844e-08, 2.424169e-08,
  2.196066e-08, 2.208689e-08, 2.267295e-08, 2.22127e-08, 2.038004e-08, 
    1.895518e-08, 2.108476e-08, 2.681895e-08, 2.914657e-08, 2.66493e-08, 
    2.437729e-08, 2.434729e-08, 2.457882e-08, 2.475537e-08, 2.435665e-08,
  2.234045e-08, 2.282919e-08, 2.285152e-08, 2.139554e-08, 1.988607e-08, 
    2.026006e-08, 2.514812e-08, 2.830386e-08, 2.801807e-08, 2.534394e-08, 
    2.403122e-08, 2.430795e-08, 2.473801e-08, 2.481985e-08, 2.451333e-08,
  2.425702e-08, 2.425064e-08, 2.416034e-08, 2.376818e-08, 2.395241e-08, 
    2.387802e-08, 2.269847e-08, 2.234339e-08, 2.375291e-08, 2.518552e-08, 
    2.675398e-08, 2.773689e-08, 2.847016e-08, 2.837047e-08, 2.798258e-08,
  2.459205e-08, 2.451783e-08, 2.415606e-08, 2.377793e-08, 2.401522e-08, 
    2.382638e-08, 2.21913e-08, 2.231331e-08, 2.35994e-08, 2.543032e-08, 
    2.667183e-08, 2.71148e-08, 2.685792e-08, 2.742279e-08, 2.787467e-08,
  2.440675e-08, 2.463968e-08, 2.422137e-08, 2.40399e-08, 2.404427e-08, 
    2.335539e-08, 2.221386e-08, 2.219107e-08, 2.412225e-08, 2.574791e-08, 
    2.627258e-08, 2.622895e-08, 2.700956e-08, 2.783975e-08, 2.784809e-08,
  2.418622e-08, 2.436204e-08, 2.414785e-08, 2.405703e-08, 2.395163e-08, 
    2.307333e-08, 2.185769e-08, 2.257556e-08, 2.441924e-08, 2.542313e-08, 
    2.565032e-08, 2.605005e-08, 2.70809e-08, 2.686045e-08, 2.66887e-08,
  2.397179e-08, 2.416057e-08, 2.424173e-08, 2.413279e-08, 2.386418e-08, 
    2.291074e-08, 2.150299e-08, 2.213248e-08, 2.440682e-08, 2.542517e-08, 
    2.553915e-08, 2.586767e-08, 2.598142e-08, 2.520324e-08, 2.501446e-08,
  2.42124e-08, 2.410087e-08, 2.407124e-08, 2.396402e-08, 2.371035e-08, 
    2.280596e-08, 2.170933e-08, 2.234673e-08, 2.444091e-08, 2.572622e-08, 
    2.554749e-08, 2.519328e-08, 2.494375e-08, 2.348208e-08, 2.316243e-08,
  2.427954e-08, 2.412056e-08, 2.406951e-08, 2.382257e-08, 2.354675e-08, 
    2.275907e-08, 2.201489e-08, 2.248301e-08, 2.273442e-08, 2.504838e-08, 
    2.510756e-08, 2.457527e-08, 2.381023e-08, 2.176941e-08, 2.098853e-08,
  2.414205e-08, 2.394234e-08, 2.377907e-08, 2.35927e-08, 2.341185e-08, 
    2.253693e-08, 2.191097e-08, 2.237348e-08, 2.372995e-08, 2.594394e-08, 
    2.504584e-08, 2.410917e-08, 2.307843e-08, 2.083067e-08, 2.037639e-08,
  2.370009e-08, 2.371539e-08, 2.355882e-08, 2.343254e-08, 2.30819e-08, 
    2.241079e-08, 2.158259e-08, 2.216813e-08, 2.365632e-08, 2.573546e-08, 
    2.455837e-08, 2.379706e-08, 2.275165e-08, 2.081747e-08, 2.040189e-08,
  2.339308e-08, 2.336765e-08, 2.340023e-08, 2.316687e-08, 2.28656e-08, 
    2.181044e-08, 2.116902e-08, 2.209445e-08, 2.378006e-08, 2.570015e-08, 
    2.404662e-08, 2.355157e-08, 2.273418e-08, 2.124347e-08, 2.075102e-08,
  2.260301e-08, 2.307946e-08, 2.39176e-08, 2.415913e-08, 2.3241e-08, 
    2.398275e-08, 2.548509e-08, 2.811771e-08, 2.880423e-08, 2.854159e-08, 
    2.698248e-08, 2.504573e-08, 2.307609e-08, 2.175472e-08, 2.062212e-08,
  2.34113e-08, 2.345747e-08, 2.398489e-08, 2.372322e-08, 2.27172e-08, 
    2.446876e-08, 2.573755e-08, 2.83688e-08, 2.88135e-08, 2.820921e-08, 
    2.59962e-08, 2.411367e-08, 2.261396e-08, 2.180655e-08, 2.101694e-08,
  2.292568e-08, 2.310914e-08, 2.395532e-08, 2.356631e-08, 2.291123e-08, 
    2.472571e-08, 2.604743e-08, 2.846701e-08, 2.901208e-08, 2.733464e-08, 
    2.493955e-08, 2.370862e-08, 2.299252e-08, 2.230163e-08, 2.161509e-08,
  2.274881e-08, 2.289711e-08, 2.373651e-08, 2.375661e-08, 2.402079e-08, 
    2.441562e-08, 2.558759e-08, 2.888077e-08, 2.867427e-08, 2.645646e-08, 
    2.495445e-08, 2.436581e-08, 2.372011e-08, 2.284764e-08, 2.247376e-08,
  2.285477e-08, 2.263768e-08, 2.378127e-08, 2.388317e-08, 2.404866e-08, 
    2.404347e-08, 2.521948e-08, 2.871911e-08, 2.887659e-08, 2.64375e-08, 
    2.538799e-08, 2.485216e-08, 2.437599e-08, 2.369455e-08, 2.380584e-08,
  2.424057e-08, 2.3131e-08, 2.340941e-08, 2.418034e-08, 2.437931e-08, 
    2.412728e-08, 2.474391e-08, 2.798802e-08, 2.831231e-08, 2.700692e-08, 
    2.606619e-08, 2.55739e-08, 2.515172e-08, 2.506053e-08, 2.49679e-08,
  2.400106e-08, 2.418497e-08, 2.371708e-08, 2.396243e-08, 2.42271e-08, 
    2.380847e-08, 2.456275e-08, 2.765547e-08, 2.803201e-08, 2.717433e-08, 
    2.672105e-08, 2.593251e-08, 2.538584e-08, 2.468079e-08, 2.502799e-08,
  2.320075e-08, 2.404337e-08, 2.401865e-08, 2.431332e-08, 2.448409e-08, 
    2.391828e-08, 2.405002e-08, 2.723308e-08, 2.814216e-08, 2.750853e-08, 
    2.709802e-08, 2.601946e-08, 2.502719e-08, 2.41935e-08, 2.459052e-08,
  2.228428e-08, 2.409987e-08, 2.416748e-08, 2.411837e-08, 2.427266e-08, 
    2.374389e-08, 2.353377e-08, 2.666106e-08, 2.805507e-08, 2.756715e-08, 
    2.733545e-08, 2.590493e-08, 2.425398e-08, 2.387493e-08, 2.465395e-08,
  2.222077e-08, 2.39155e-08, 2.435554e-08, 2.455067e-08, 2.461366e-08, 
    2.402683e-08, 2.326276e-08, 2.581493e-08, 2.803666e-08, 2.779688e-08, 
    2.736308e-08, 2.566762e-08, 2.400413e-08, 2.368408e-08, 2.463997e-08,
  2.398232e-08, 2.410108e-08, 2.350012e-08, 2.388435e-08, 2.510369e-08, 
    2.662423e-08, 2.527126e-08, 2.275715e-08, 2.134395e-08, 2.056249e-08, 
    2.035781e-08, 2.044764e-08, 2.09124e-08, 2.113395e-08, 2.130655e-08,
  2.386208e-08, 2.396808e-08, 2.380819e-08, 2.351546e-08, 2.368673e-08, 
    2.742655e-08, 2.594603e-08, 2.312305e-08, 2.126489e-08, 2.038342e-08, 
    2.010667e-08, 2.008245e-08, 2.043943e-08, 2.060275e-08, 2.0654e-08,
  2.345725e-08, 2.328526e-08, 2.337112e-08, 2.343038e-08, 2.293396e-08, 
    2.714397e-08, 2.678538e-08, 2.343498e-08, 2.099131e-08, 2.013063e-08, 
    1.981462e-08, 1.990823e-08, 2.045961e-08, 2.061105e-08, 2.064681e-08,
  2.349801e-08, 2.367871e-08, 2.311219e-08, 2.357178e-08, 2.17434e-08, 
    2.664169e-08, 2.918547e-08, 2.487687e-08, 2.134344e-08, 1.99571e-08, 
    1.96206e-08, 1.994288e-08, 2.053217e-08, 2.086838e-08, 2.116614e-08,
  2.354905e-08, 2.356088e-08, 2.309893e-08, 2.353192e-08, 2.211326e-08, 
    2.650922e-08, 2.972665e-08, 2.546655e-08, 2.101502e-08, 1.988121e-08, 
    1.945733e-08, 2.030596e-08, 2.105588e-08, 2.189222e-08, 2.21612e-08,
  2.301423e-08, 2.399356e-08, 2.346719e-08, 2.343922e-08, 2.299259e-08, 
    2.572902e-08, 2.958874e-08, 2.60097e-08, 2.115406e-08, 1.980099e-08, 
    1.946931e-08, 2.095511e-08, 2.184507e-08, 2.282367e-08, 2.26894e-08,
  2.108326e-08, 2.312635e-08, 2.373553e-08, 2.360548e-08, 2.296237e-08, 
    2.499412e-08, 2.940801e-08, 2.676639e-08, 2.167941e-08, 2.01752e-08, 
    1.995656e-08, 2.152697e-08, 2.252442e-08, 2.33796e-08, 2.336334e-08,
  2.005938e-08, 2.198284e-08, 2.372592e-08, 2.361632e-08, 2.352218e-08, 
    2.433183e-08, 2.899863e-08, 2.728801e-08, 2.206179e-08, 2.068469e-08, 
    2.053013e-08, 2.187946e-08, 2.286416e-08, 2.335557e-08, 2.33513e-08,
  1.982865e-08, 2.072412e-08, 2.315271e-08, 2.365271e-08, 2.345781e-08, 
    2.383462e-08, 2.836961e-08, 2.800519e-08, 2.278862e-08, 2.131019e-08, 
    2.113086e-08, 2.215373e-08, 2.279562e-08, 2.287758e-08, 2.303461e-08,
  2.10853e-08, 2.08454e-08, 2.235856e-08, 2.312233e-08, 2.411402e-08, 
    2.342893e-08, 2.736585e-08, 2.852991e-08, 2.363207e-08, 2.204949e-08, 
    2.16788e-08, 2.225423e-08, 2.275697e-08, 2.302074e-08, 2.317191e-08,
  2.240313e-08, 2.31823e-08, 2.391957e-08, 2.5077e-08, 2.384426e-08, 
    2.17235e-08, 2.238512e-08, 2.245258e-08, 2.266164e-08, 2.270572e-08, 
    2.2728e-08, 2.27801e-08, 2.319866e-08, 2.351638e-08, 2.343913e-08,
  2.240878e-08, 2.335675e-08, 2.376844e-08, 2.421534e-08, 2.295543e-08, 
    2.196929e-08, 2.172629e-08, 2.232651e-08, 2.243256e-08, 2.226082e-08, 
    2.262136e-08, 2.27466e-08, 2.306138e-08, 2.296338e-08, 2.273498e-08,
  2.202067e-08, 2.342598e-08, 2.334509e-08, 2.242349e-08, 2.276675e-08, 
    2.158704e-08, 2.083012e-08, 2.246692e-08, 2.197537e-08, 2.217313e-08, 
    2.238502e-08, 2.237141e-08, 2.24757e-08, 2.235171e-08, 2.226574e-08,
  2.162094e-08, 2.345739e-08, 2.36656e-08, 2.271464e-08, 2.029332e-08, 
    2.212065e-08, 2.30791e-08, 2.236883e-08, 2.166547e-08, 2.19197e-08, 
    2.220772e-08, 2.196369e-08, 2.190536e-08, 2.178846e-08, 2.178904e-08,
  2.093271e-08, 2.301527e-08, 2.338828e-08, 2.324619e-08, 2.050446e-08, 
    2.304167e-08, 2.401224e-08, 2.351237e-08, 2.194624e-08, 2.186279e-08, 
    2.192365e-08, 2.145321e-08, 2.137819e-08, 2.125151e-08, 2.137586e-08,
  2.088911e-08, 2.165203e-08, 2.351557e-08, 2.398665e-08, 2.103848e-08, 
    2.407722e-08, 2.599656e-08, 2.150615e-08, 2.078538e-08, 2.318292e-08, 
    2.199158e-08, 2.143603e-08, 2.107581e-08, 2.116002e-08, 2.143912e-08,
  2.157813e-08, 2.041372e-08, 2.307805e-08, 2.464429e-08, 2.160584e-08, 
    2.440709e-08, 2.738893e-08, 2.184691e-08, 2.063495e-08, 2.222044e-08, 
    2.14419e-08, 2.149844e-08, 2.114862e-08, 2.125453e-08, 2.144735e-08,
  2.250937e-08, 2.075689e-08, 2.188195e-08, 2.441288e-08, 2.267174e-08, 
    2.399225e-08, 2.832014e-08, 2.325288e-08, 2.050837e-08, 2.132568e-08, 
    2.104237e-08, 2.158312e-08, 2.153496e-08, 2.16284e-08, 2.197658e-08,
  2.340386e-08, 2.18269e-08, 2.108061e-08, 2.368755e-08, 2.314354e-08, 
    2.318568e-08, 2.835942e-08, 2.531659e-08, 2.084684e-08, 2.066759e-08, 
    2.065215e-08, 2.187745e-08, 2.202088e-08, 2.210245e-08, 2.216956e-08,
  2.416165e-08, 2.29421e-08, 2.170049e-08, 2.249819e-08, 2.39177e-08, 
    2.293683e-08, 2.734398e-08, 2.704267e-08, 2.201875e-08, 2.013712e-08, 
    2.036863e-08, 2.213809e-08, 2.249952e-08, 2.248363e-08, 2.228413e-08,
  2.186645e-08, 2.376549e-08, 2.472708e-08, 2.378559e-08, 2.228157e-08, 
    2.354935e-08, 2.400867e-08, 2.377704e-08, 2.438045e-08, 2.436185e-08, 
    2.424285e-08, 2.42376e-08, 2.345045e-08, 2.179996e-08, 2.143767e-08,
  2.212848e-08, 2.435803e-08, 2.414624e-08, 2.274415e-08, 2.176929e-08, 
    2.353264e-08, 2.274749e-08, 2.320766e-08, 2.354115e-08, 2.36034e-08, 
    2.386085e-08, 2.404756e-08, 2.386142e-08, 2.245269e-08, 2.191303e-08,
  2.185651e-08, 2.378785e-08, 2.278861e-08, 2.157895e-08, 2.208961e-08, 
    2.213657e-08, 2.293729e-08, 2.310888e-08, 2.292155e-08, 2.320359e-08, 
    2.331113e-08, 2.337367e-08, 2.321315e-08, 2.273575e-08, 2.248155e-08,
  2.177456e-08, 2.355409e-08, 2.300891e-08, 2.13639e-08, 2.166205e-08, 
    2.215644e-08, 2.484214e-08, 2.294593e-08, 2.265064e-08, 2.294497e-08, 
    2.30167e-08, 2.285238e-08, 2.265821e-08, 2.225873e-08, 2.240944e-08,
  2.221049e-08, 2.209574e-08, 2.362982e-08, 2.13884e-08, 2.045247e-08, 
    2.082865e-08, 2.440767e-08, 2.415735e-08, 2.281558e-08, 2.281806e-08, 
    2.262581e-08, 2.26368e-08, 2.248155e-08, 2.232979e-08, 2.218866e-08,
  2.268054e-08, 2.109856e-08, 2.381833e-08, 2.2547e-08, 2.067428e-08, 
    2.039597e-08, 2.374733e-08, 2.405189e-08, 2.281137e-08, 2.330422e-08, 
    2.262237e-08, 2.260222e-08, 2.250494e-08, 2.219381e-08, 2.160484e-08,
  2.420334e-08, 2.233191e-08, 2.274851e-08, 2.369203e-08, 2.130603e-08, 
    2.098673e-08, 2.272743e-08, 2.331008e-08, 2.289087e-08, 2.402855e-08, 
    2.273926e-08, 2.241709e-08, 2.232968e-08, 2.183578e-08, 2.10182e-08,
  2.517726e-08, 2.403038e-08, 2.204668e-08, 2.39836e-08, 2.240184e-08, 
    2.293497e-08, 2.321178e-08, 2.227297e-08, 2.272415e-08, 2.407582e-08, 
    2.246205e-08, 2.226463e-08, 2.227578e-08, 2.317307e-08, 2.436146e-08,
  2.473187e-08, 2.501574e-08, 2.348006e-08, 2.359703e-08, 2.260622e-08, 
    2.297077e-08, 2.389922e-08, 2.229791e-08, 2.236534e-08, 2.436409e-08, 
    2.218953e-08, 2.19782e-08, 2.242876e-08, 2.361772e-08, 2.62335e-08,
  2.403458e-08, 2.482404e-08, 2.508886e-08, 2.381124e-08, 2.336481e-08, 
    2.281829e-08, 2.46502e-08, 2.326688e-08, 2.156715e-08, 2.243705e-08, 
    2.225739e-08, 2.324496e-08, 2.194197e-08, 2.353394e-08, 2.607099e-08,
  2.325322e-08, 2.404679e-08, 2.274614e-08, 2.2598e-08, 2.328898e-08, 
    2.346513e-08, 2.262434e-08, 2.309733e-08, 2.338898e-08, 2.338159e-08, 
    2.335642e-08, 2.324861e-08, 2.318812e-08, 2.148062e-08, 2.111628e-08,
  2.301598e-08, 2.316047e-08, 2.225028e-08, 2.258596e-08, 2.358729e-08, 
    2.384694e-08, 2.259259e-08, 2.179054e-08, 2.257305e-08, 2.23843e-08, 
    2.258359e-08, 2.348467e-08, 2.409265e-08, 2.372041e-08, 2.237855e-08,
  2.292812e-08, 2.272003e-08, 2.194902e-08, 2.175792e-08, 2.298235e-08, 
    2.454543e-08, 2.356948e-08, 2.128801e-08, 2.218072e-08, 2.18322e-08, 
    2.175938e-08, 2.240435e-08, 2.353691e-08, 2.460994e-08, 2.428952e-08,
  2.320829e-08, 2.326765e-08, 2.254244e-08, 2.160736e-08, 2.178548e-08, 
    2.39298e-08, 2.475573e-08, 2.255887e-08, 2.110121e-08, 2.166801e-08, 
    2.14875e-08, 2.201394e-08, 2.267505e-08, 2.406897e-08, 2.450581e-08,
  2.34758e-08, 2.343305e-08, 2.372875e-08, 2.224124e-08, 2.121122e-08, 
    2.222827e-08, 2.406727e-08, 2.371549e-08, 2.196179e-08, 2.087302e-08, 
    2.028811e-08, 2.076125e-08, 2.141129e-08, 2.30155e-08, 2.374366e-08,
  2.402442e-08, 2.395257e-08, 2.412813e-08, 2.386791e-08, 2.236465e-08, 
    2.163017e-08, 2.347008e-08, 2.388815e-08, 2.385171e-08, 2.264333e-08, 
    2.076736e-08, 1.978808e-08, 1.941481e-08, 2.06966e-08, 2.297994e-08,
  2.405943e-08, 2.39669e-08, 2.45582e-08, 2.452773e-08, 2.356837e-08, 
    2.219262e-08, 2.293881e-08, 2.344468e-08, 2.380675e-08, 2.430415e-08, 
    2.287403e-08, 2.212187e-08, 2.081994e-08, 1.916536e-08, 1.925773e-08,
  2.423184e-08, 2.380429e-08, 2.442455e-08, 2.509954e-08, 2.452755e-08, 
    2.326147e-08, 2.309503e-08, 2.316841e-08, 2.304801e-08, 2.336029e-08, 
    2.341554e-08, 2.470387e-08, 2.625456e-08, 2.658981e-08, 2.404641e-08,
  2.483874e-08, 2.404405e-08, 2.394126e-08, 2.479318e-08, 2.554761e-08, 
    2.385475e-08, 2.328932e-08, 2.323476e-08, 2.30737e-08, 2.357068e-08, 
    2.33994e-08, 2.531553e-08, 2.854678e-08, 3.23476e-08, 3.446285e-08,
  2.489864e-08, 2.475631e-08, 2.384251e-08, 2.394184e-08, 2.550116e-08, 
    2.536399e-08, 2.383641e-08, 2.366579e-08, 2.288304e-08, 2.307488e-08, 
    2.383909e-08, 2.577121e-08, 2.778748e-08, 3.218101e-08, 3.391145e-08,
  2.303909e-08, 2.299379e-08, 2.297121e-08, 2.265053e-08, 2.320433e-08, 
    2.42309e-08, 2.11259e-08, 2.023684e-08, 2.194196e-08, 2.3146e-08, 
    2.470576e-08, 2.526887e-08, 2.419112e-08, 2.183767e-08, 2.195483e-08,
  2.337361e-08, 2.36926e-08, 2.34876e-08, 2.26459e-08, 2.301701e-08, 
    2.475158e-08, 2.18508e-08, 1.910304e-08, 2.09425e-08, 2.245e-08, 
    2.392703e-08, 2.464077e-08, 2.461949e-08, 2.29903e-08, 2.269451e-08,
  2.391672e-08, 2.434287e-08, 2.418022e-08, 2.310398e-08, 2.24535e-08, 
    2.420588e-08, 2.369902e-08, 1.918597e-08, 1.979467e-08, 2.161052e-08, 
    2.286243e-08, 2.380935e-08, 2.372721e-08, 2.374999e-08, 2.318877e-08,
  2.407555e-08, 2.473129e-08, 2.484761e-08, 2.408214e-08, 2.313486e-08, 
    2.405563e-08, 2.512386e-08, 2.174211e-08, 1.890126e-08, 2.018258e-08, 
    2.168271e-08, 2.312887e-08, 2.316308e-08, 2.269449e-08, 2.270508e-08,
  2.388687e-08, 2.458533e-08, 2.515061e-08, 2.469916e-08, 2.323308e-08, 
    2.340262e-08, 2.453062e-08, 2.407759e-08, 2.127859e-08, 2.017221e-08, 
    2.03697e-08, 2.193869e-08, 2.242784e-08, 2.175239e-08, 2.196814e-08,
  2.380249e-08, 2.397125e-08, 2.49384e-08, 2.565933e-08, 2.406223e-08, 
    2.340481e-08, 2.413412e-08, 2.460202e-08, 2.440633e-08, 2.256628e-08, 
    2.172567e-08, 2.10828e-08, 2.124642e-08, 2.100299e-08, 2.09022e-08,
  2.431833e-08, 2.356029e-08, 2.404274e-08, 2.556945e-08, 2.523285e-08, 
    2.363676e-08, 2.348858e-08, 2.392816e-08, 2.439991e-08, 2.483572e-08, 
    2.514991e-08, 2.540826e-08, 2.256538e-08, 2.04573e-08, 2.035858e-08,
  2.488408e-08, 2.369798e-08, 2.281786e-08, 2.471661e-08, 2.61708e-08, 
    2.448743e-08, 2.35214e-08, 2.374012e-08, 2.42288e-08, 2.490876e-08, 
    2.715109e-08, 3.048382e-08, 3.085469e-08, 2.721912e-08, 2.621618e-08,
  2.501594e-08, 2.432417e-08, 2.290574e-08, 2.301242e-08, 2.533043e-08, 
    2.599394e-08, 2.425479e-08, 2.367315e-08, 2.431928e-08, 2.564148e-08, 
    2.823786e-08, 3.197682e-08, 3.344955e-08, 3.264172e-08, 3.226906e-08,
  2.511726e-08, 2.471218e-08, 2.328017e-08, 2.27625e-08, 2.375909e-08, 
    2.518125e-08, 2.569792e-08, 2.412489e-08, 2.370757e-08, 2.437983e-08, 
    2.727002e-08, 3.046337e-08, 3.183252e-08, 3.092022e-08, 2.824107e-08,
  2.449395e-08, 2.416332e-08, 2.418804e-08, 2.45338e-08, 2.421704e-08, 
    2.417234e-08, 2.335372e-08, 2.073334e-08, 2.123483e-08, 2.23709e-08, 
    2.29923e-08, 2.239177e-08, 2.223695e-08, 2.250675e-08, 2.366815e-08,
  2.431535e-08, 2.414036e-08, 2.457272e-08, 2.490439e-08, 2.439283e-08, 
    2.379636e-08, 2.366597e-08, 2.151725e-08, 2.151401e-08, 2.223263e-08, 
    2.249715e-08, 2.167262e-08, 2.15162e-08, 2.185505e-08, 2.306239e-08,
  2.406418e-08, 2.418395e-08, 2.481465e-08, 2.495642e-08, 2.432223e-08, 
    2.387384e-08, 2.408437e-08, 2.235892e-08, 2.16306e-08, 2.242427e-08, 
    2.310412e-08, 2.235672e-08, 2.065737e-08, 2.224713e-08, 2.3038e-08,
  2.36704e-08, 2.407278e-08, 2.506199e-08, 2.51124e-08, 2.415175e-08, 
    2.465874e-08, 2.42559e-08, 2.3173e-08, 2.21861e-08, 2.318268e-08, 
    2.453582e-08, 2.441059e-08, 2.223705e-08, 2.069005e-08, 2.151326e-08,
  2.31097e-08, 2.387576e-08, 2.524454e-08, 2.546022e-08, 2.41026e-08, 
    2.407867e-08, 2.441207e-08, 2.38638e-08, 2.384004e-08, 2.513756e-08, 
    2.742125e-08, 2.776403e-08, 2.488334e-08, 2.181152e-08, 2.052946e-08,
  2.312693e-08, 2.351125e-08, 2.507957e-08, 2.572697e-08, 2.481895e-08, 
    2.440066e-08, 2.46916e-08, 2.48576e-08, 2.540746e-08, 2.686608e-08, 
    3.01371e-08, 3.118093e-08, 2.889852e-08, 2.556268e-08, 2.124808e-08,
  2.319489e-08, 2.316897e-08, 2.427585e-08, 2.538844e-08, 2.524488e-08, 
    2.456017e-08, 2.471659e-08, 2.50179e-08, 2.599394e-08, 2.798418e-08, 
    3.034048e-08, 3.19185e-08, 3.263323e-08, 3.188244e-08, 2.976024e-08,
  2.392802e-08, 2.334961e-08, 2.34286e-08, 2.470521e-08, 2.51035e-08, 
    2.486683e-08, 2.471327e-08, 2.503769e-08, 2.583148e-08, 2.703317e-08, 
    2.940736e-08, 3.062468e-08, 3.186893e-08, 3.452334e-08, 3.66234e-08,
  2.464622e-08, 2.410101e-08, 2.356832e-08, 2.325977e-08, 2.39182e-08, 
    2.463881e-08, 2.461797e-08, 2.452122e-08, 2.47841e-08, 2.555234e-08, 
    2.690904e-08, 2.817593e-08, 2.789941e-08, 2.85458e-08, 3.167515e-08,
  2.44457e-08, 2.453927e-08, 2.422619e-08, 2.34126e-08, 2.26813e-08, 
    2.273048e-08, 2.374694e-08, 2.411808e-08, 2.407803e-08, 2.425608e-08, 
    2.465494e-08, 2.605509e-08, 2.667868e-08, 2.460119e-08, 2.39437e-08,
  2.48002e-08, 2.475808e-08, 2.483242e-08, 2.456408e-08, 2.452744e-08, 
    2.461298e-08, 2.453762e-08, 2.468574e-08, 2.420281e-08, 2.369648e-08, 
    2.376406e-08, 2.692623e-08, 2.805003e-08, 2.343991e-08, 2.181865e-08,
  2.484487e-08, 2.489862e-08, 2.462112e-08, 2.445734e-08, 2.459724e-08, 
    2.459446e-08, 2.462433e-08, 2.473693e-08, 2.404406e-08, 2.389673e-08, 
    2.559326e-08, 3.00019e-08, 2.933218e-08, 2.332854e-08, 2.097832e-08,
  2.467485e-08, 2.445871e-08, 2.428684e-08, 2.423127e-08, 2.464202e-08, 
    2.467968e-08, 2.460716e-08, 2.458577e-08, 2.399922e-08, 2.487912e-08, 
    2.836177e-08, 3.183116e-08, 2.973587e-08, 2.410742e-08, 2.174846e-08,
  2.456309e-08, 2.424149e-08, 2.409909e-08, 2.446227e-08, 2.463426e-08, 
    2.494789e-08, 2.500198e-08, 2.431885e-08, 2.462311e-08, 2.686355e-08, 
    2.993188e-08, 3.234538e-08, 3.202125e-08, 2.564976e-08, 2.182294e-08,
  2.422298e-08, 2.389306e-08, 2.390187e-08, 2.442934e-08, 2.52402e-08, 
    2.485801e-08, 2.517459e-08, 2.443725e-08, 2.577142e-08, 2.803252e-08, 
    2.943927e-08, 3.22497e-08, 3.305704e-08, 2.988638e-08, 2.275199e-08,
  2.380167e-08, 2.344952e-08, 2.381297e-08, 2.466947e-08, 2.538699e-08, 
    2.533833e-08, 2.499189e-08, 2.580905e-08, 2.727557e-08, 2.674785e-08, 
    2.84867e-08, 3.116763e-08, 3.41475e-08, 3.331117e-08, 2.495336e-08,
  2.377382e-08, 2.355015e-08, 2.36462e-08, 2.454298e-08, 2.515226e-08, 
    2.514268e-08, 2.537825e-08, 2.581788e-08, 2.594278e-08, 2.61029e-08, 
    2.686598e-08, 2.830244e-08, 3.113705e-08, 3.421225e-08, 3.216958e-08,
  2.418739e-08, 2.367271e-08, 2.338231e-08, 2.394634e-08, 2.443996e-08, 
    2.470174e-08, 2.480956e-08, 2.5164e-08, 2.455672e-08, 2.493598e-08, 
    2.533075e-08, 2.603957e-08, 2.621286e-08, 3.038455e-08, 3.319075e-08,
  2.446313e-08, 2.438702e-08, 2.361791e-08, 2.326497e-08, 2.328128e-08, 
    2.340657e-08, 2.353213e-08, 2.341067e-08, 2.393931e-08, 2.399398e-08, 
    2.420579e-08, 2.47157e-08, 2.504398e-08, 2.430036e-08, 2.636564e-08,
  2.462172e-08, 2.48873e-08, 2.489762e-08, 2.387178e-08, 2.335417e-08, 
    2.29344e-08, 2.285689e-08, 2.28545e-08, 2.292149e-08, 2.320106e-08, 
    2.356963e-08, 2.41792e-08, 2.499069e-08, 2.434024e-08, 2.36618e-08,
  2.45535e-08, 2.451211e-08, 2.449843e-08, 2.483545e-08, 2.477691e-08, 
    2.461426e-08, 2.434537e-08, 2.453285e-08, 2.486088e-08, 2.567623e-08, 
    2.580109e-08, 2.925323e-08, 3.266243e-08, 2.59062e-08, 2.18395e-08,
  2.469425e-08, 2.497791e-08, 2.496853e-08, 2.493591e-08, 2.498553e-08, 
    2.457575e-08, 2.443066e-08, 2.464089e-08, 2.519745e-08, 2.583415e-08, 
    2.611949e-08, 2.955818e-08, 3.222345e-08, 2.544482e-08, 2.172644e-08,
  2.47453e-08, 2.516198e-08, 2.511887e-08, 2.510286e-08, 2.494858e-08, 
    2.440188e-08, 2.418954e-08, 2.462268e-08, 2.532204e-08, 2.585785e-08, 
    2.603144e-08, 2.943745e-08, 3.173004e-08, 2.543817e-08, 2.184234e-08,
  2.480747e-08, 2.499264e-08, 2.491321e-08, 2.497623e-08, 2.462084e-08, 
    2.432964e-08, 2.481434e-08, 2.475395e-08, 2.559629e-08, 2.590757e-08, 
    2.593847e-08, 2.891419e-08, 3.095134e-08, 2.567823e-08, 2.171327e-08,
  2.475306e-08, 2.468643e-08, 2.487934e-08, 2.476942e-08, 2.453413e-08, 
    2.41283e-08, 2.479715e-08, 2.494042e-08, 2.577245e-08, 2.54765e-08, 
    2.555004e-08, 2.732071e-08, 2.957495e-08, 2.646572e-08, 2.231357e-08,
  2.471365e-08, 2.459649e-08, 2.45643e-08, 2.442527e-08, 2.403378e-08, 
    2.420162e-08, 2.41889e-08, 2.484691e-08, 2.521797e-08, 2.505041e-08, 
    2.496468e-08, 2.583375e-08, 2.810476e-08, 2.743787e-08, 2.292391e-08,
  2.482251e-08, 2.459316e-08, 2.452188e-08, 2.420673e-08, 2.411257e-08, 
    2.410523e-08, 2.442556e-08, 2.473797e-08, 2.470128e-08, 2.482935e-08, 
    2.42009e-08, 2.494122e-08, 2.610857e-08, 2.736378e-08, 2.481314e-08,
  2.463609e-08, 2.46205e-08, 2.44232e-08, 2.414784e-08, 2.398455e-08, 
    2.401522e-08, 2.406748e-08, 2.410274e-08, 2.402783e-08, 2.381909e-08, 
    2.386717e-08, 2.445575e-08, 2.484694e-08, 2.537684e-08, 2.557576e-08,
  2.424632e-08, 2.430352e-08, 2.421831e-08, 2.404567e-08, 2.394361e-08, 
    2.367168e-08, 2.359057e-08, 2.318673e-08, 2.314999e-08, 2.327117e-08, 
    2.344393e-08, 2.371425e-08, 2.439507e-08, 2.425676e-08, 2.479444e-08,
  2.441408e-08, 2.435122e-08, 2.444549e-08, 2.433455e-08, 2.415245e-08, 
    2.392193e-08, 2.360645e-08, 2.344194e-08, 2.324873e-08, 2.306255e-08, 
    2.310974e-08, 2.329906e-08, 2.374883e-08, 2.454448e-08, 2.39603e-08,
  2.441226e-08, 2.42003e-08, 2.430896e-08, 2.493745e-08, 2.530346e-08, 
    2.506821e-08, 2.484688e-08, 2.436714e-08, 2.510461e-08, 2.544767e-08, 
    2.555987e-08, 2.636285e-08, 2.492996e-08, 2.384634e-08, 2.452436e-08,
  2.457686e-08, 2.422855e-08, 2.441919e-08, 2.511767e-08, 2.549647e-08, 
    2.476794e-08, 2.476705e-08, 2.42029e-08, 2.508631e-08, 2.533604e-08, 
    2.517935e-08, 2.59678e-08, 2.497553e-08, 2.383622e-08, 2.455685e-08,
  2.413568e-08, 2.44044e-08, 2.464218e-08, 2.523472e-08, 2.520775e-08, 
    2.484049e-08, 2.455103e-08, 2.436629e-08, 2.477879e-08, 2.495403e-08, 
    2.482247e-08, 2.591135e-08, 2.512895e-08, 2.43455e-08, 2.437497e-08,
  2.415873e-08, 2.463688e-08, 2.488144e-08, 2.495515e-08, 2.500151e-08, 
    2.500897e-08, 2.461915e-08, 2.415752e-08, 2.462819e-08, 2.469456e-08, 
    2.44167e-08, 2.543702e-08, 2.522388e-08, 2.41015e-08, 2.43529e-08,
  2.436261e-08, 2.461615e-08, 2.468745e-08, 2.46692e-08, 2.48385e-08, 
    2.467024e-08, 2.459444e-08, 2.409852e-08, 2.432724e-08, 2.417508e-08, 
    2.410841e-08, 2.476129e-08, 2.524116e-08, 2.434618e-08, 2.446466e-08,
  2.462675e-08, 2.470771e-08, 2.461326e-08, 2.474805e-08, 2.471536e-08, 
    2.472225e-08, 2.433986e-08, 2.416589e-08, 2.42029e-08, 2.394165e-08, 
    2.380182e-08, 2.410825e-08, 2.494358e-08, 2.43452e-08, 2.397444e-08,
  2.572617e-08, 2.550351e-08, 2.51558e-08, 2.491231e-08, 2.48776e-08, 
    2.467185e-08, 2.45059e-08, 2.441734e-08, 2.4159e-08, 2.385921e-08, 
    2.356087e-08, 2.361265e-08, 2.435715e-08, 2.466069e-08, 2.42679e-08,
  2.500119e-08, 2.516553e-08, 2.508884e-08, 2.492691e-08, 2.475104e-08, 
    2.452283e-08, 2.435173e-08, 2.411706e-08, 2.398437e-08, 2.390968e-08, 
    2.365969e-08, 2.354191e-08, 2.389907e-08, 2.441104e-08, 2.468306e-08,
  2.428232e-08, 2.439356e-08, 2.438691e-08, 2.434246e-08, 2.424739e-08, 
    2.430903e-08, 2.436096e-08, 2.440061e-08, 2.449837e-08, 2.453419e-08, 
    2.416124e-08, 2.353231e-08, 2.350093e-08, 2.448316e-08, 2.406952e-08,
  2.45604e-08, 2.443625e-08, 2.431191e-08, 2.432047e-08, 2.433022e-08, 
    2.450662e-08, 2.460923e-08, 2.468768e-08, 2.450869e-08, 2.454258e-08, 
    2.421613e-08, 2.38837e-08, 2.332871e-08, 2.385831e-08, 2.392247e-08,
  2.475649e-08, 2.491311e-08, 2.407392e-08, 2.514901e-08, 2.521675e-08, 
    2.469726e-08, 2.48893e-08, 2.460509e-08, 2.445389e-08, 2.436248e-08, 
    2.458165e-08, 2.491195e-08, 2.459429e-08, 2.292754e-08, 2.19484e-08,
  2.500351e-08, 2.469405e-08, 2.441546e-08, 2.56123e-08, 2.528109e-08, 
    2.4634e-08, 2.491427e-08, 2.456602e-08, 2.442154e-08, 2.436226e-08, 
    2.443052e-08, 2.471427e-08, 2.465484e-08, 2.309282e-08, 2.200412e-08,
  2.457999e-08, 2.41237e-08, 2.44531e-08, 2.495276e-08, 2.47579e-08, 
    2.465731e-08, 2.467768e-08, 2.502618e-08, 2.451245e-08, 2.435493e-08, 
    2.412679e-08, 2.445235e-08, 2.447475e-08, 2.372889e-08, 2.204934e-08,
  2.443574e-08, 2.427097e-08, 2.454681e-08, 2.490494e-08, 2.495788e-08, 
    2.526857e-08, 2.49351e-08, 2.453667e-08, 2.447491e-08, 2.46323e-08, 
    2.417396e-08, 2.41956e-08, 2.441263e-08, 2.351117e-08, 2.262794e-08,
  2.478661e-08, 2.46444e-08, 2.458732e-08, 2.480724e-08, 2.477947e-08, 
    2.480324e-08, 2.508198e-08, 2.471105e-08, 2.475114e-08, 2.463642e-08, 
    2.432609e-08, 2.399051e-08, 2.449718e-08, 2.377116e-08, 2.262258e-08,
  2.499993e-08, 2.479297e-08, 2.471151e-08, 2.514698e-08, 2.523921e-08, 
    2.516047e-08, 2.480311e-08, 2.463322e-08, 2.453331e-08, 2.476795e-08, 
    2.474487e-08, 2.398572e-08, 2.422983e-08, 2.393802e-08, 2.236096e-08,
  2.526599e-08, 2.527388e-08, 2.52191e-08, 2.525699e-08, 2.509885e-08, 
    2.473458e-08, 2.454616e-08, 2.442483e-08, 2.442172e-08, 2.477948e-08, 
    2.517929e-08, 2.458235e-08, 2.402837e-08, 2.44844e-08, 2.231415e-08,
  2.398285e-08, 2.421302e-08, 2.451235e-08, 2.46252e-08, 2.45415e-08, 
    2.434517e-08, 2.434777e-08, 2.404609e-08, 2.459852e-08, 2.499159e-08, 
    2.526506e-08, 2.494648e-08, 2.386637e-08, 2.481961e-08, 2.364952e-08,
  2.385118e-08, 2.41708e-08, 2.425317e-08, 2.439989e-08, 2.429563e-08, 
    2.436454e-08, 2.420092e-08, 2.435974e-08, 2.47883e-08, 2.470566e-08, 
    2.476388e-08, 2.504373e-08, 2.414537e-08, 2.426221e-08, 2.426742e-08,
  2.495156e-08, 2.490866e-08, 2.479163e-08, 2.464327e-08, 2.439376e-08, 
    2.432753e-08, 2.421248e-08, 2.440026e-08, 2.419486e-08, 2.42355e-08, 
    2.441752e-08, 2.459567e-08, 2.432295e-08, 2.385223e-08, 2.426934e-08,
  2.477426e-08, 2.527825e-08, 2.400562e-08, 2.454414e-08, 2.544603e-08, 
    2.520229e-08, 2.503196e-08, 2.507207e-08, 2.461941e-08, 2.479362e-08, 
    2.421257e-08, 2.326553e-08, 2.256957e-08, 2.186268e-08, 2.232155e-08,
  2.486708e-08, 2.511053e-08, 2.400477e-08, 2.455698e-08, 2.530619e-08, 
    2.496176e-08, 2.559819e-08, 2.502565e-08, 2.461995e-08, 2.490564e-08, 
    2.449237e-08, 2.327926e-08, 2.22515e-08, 2.229574e-08, 2.278298e-08,
  2.492879e-08, 2.442138e-08, 2.390927e-08, 2.460459e-08, 2.521887e-08, 
    2.498272e-08, 2.497886e-08, 2.497598e-08, 2.458047e-08, 2.487944e-08, 
    2.464367e-08, 2.325031e-08, 2.252072e-08, 2.276962e-08, 2.274542e-08,
  2.485334e-08, 2.458487e-08, 2.440785e-08, 2.484445e-08, 2.51841e-08, 
    2.5762e-08, 2.513239e-08, 2.454179e-08, 2.437408e-08, 2.478579e-08, 
    2.50216e-08, 2.354934e-08, 2.221594e-08, 2.231164e-08, 2.305588e-08,
  2.531594e-08, 2.518546e-08, 2.491614e-08, 2.493949e-08, 2.509518e-08, 
    2.487386e-08, 2.508793e-08, 2.441674e-08, 2.435717e-08, 2.451612e-08, 
    2.51542e-08, 2.393861e-08, 2.239881e-08, 2.246034e-08, 2.326227e-08,
  2.523073e-08, 2.512427e-08, 2.483472e-08, 2.474818e-08, 2.466792e-08, 
    2.464981e-08, 2.441713e-08, 2.446902e-08, 2.420663e-08, 2.437523e-08, 
    2.503499e-08, 2.459935e-08, 2.234941e-08, 2.19425e-08, 2.280753e-08,
  2.472678e-08, 2.46759e-08, 2.45017e-08, 2.437789e-08, 2.439481e-08, 
    2.435276e-08, 2.454371e-08, 2.423042e-08, 2.417812e-08, 2.466474e-08, 
    2.462867e-08, 2.506656e-08, 2.287376e-08, 2.159996e-08, 2.200036e-08,
  2.460269e-08, 2.445469e-08, 2.434385e-08, 2.442448e-08, 2.443778e-08, 
    2.462356e-08, 2.451856e-08, 2.440723e-08, 2.450349e-08, 2.440812e-08, 
    2.428871e-08, 2.49963e-08, 2.38298e-08, 2.215244e-08, 2.182293e-08,
  2.491347e-08, 2.491542e-08, 2.48374e-08, 2.486405e-08, 2.492474e-08, 
    2.478951e-08, 2.451313e-08, 2.449625e-08, 2.443353e-08, 2.42991e-08, 
    2.406182e-08, 2.468302e-08, 2.441148e-08, 2.310705e-08, 2.210964e-08,
  2.453503e-08, 2.454497e-08, 2.454023e-08, 2.484175e-08, 2.486368e-08, 
    2.468365e-08, 2.467074e-08, 2.467964e-08, 2.45414e-08, 2.426303e-08, 
    2.410152e-08, 2.416252e-08, 2.458559e-08, 2.392994e-08, 2.256911e-08,
  2.410082e-08, 2.490991e-08, 2.475826e-08, 2.45902e-08, 2.501802e-08, 
    2.507456e-08, 2.525514e-08, 2.498416e-08, 2.41019e-08, 2.428212e-08, 
    2.38508e-08, 2.275415e-08, 2.380599e-08, 2.443293e-08, 2.463991e-08,
  2.444173e-08, 2.518924e-08, 2.488772e-08, 2.472484e-08, 2.507653e-08, 
    2.486512e-08, 2.502674e-08, 2.440857e-08, 2.410961e-08, 2.446375e-08, 
    2.42036e-08, 2.304197e-08, 2.373637e-08, 2.465304e-08, 2.474074e-08,
  2.492009e-08, 2.526494e-08, 2.502278e-08, 2.49944e-08, 2.495353e-08, 
    2.460901e-08, 2.463167e-08, 2.452681e-08, 2.417652e-08, 2.428011e-08, 
    2.425041e-08, 2.318692e-08, 2.354801e-08, 2.509456e-08, 2.497349e-08,
  2.513213e-08, 2.521968e-08, 2.517513e-08, 2.491051e-08, 2.477509e-08, 
    2.53489e-08, 2.461091e-08, 2.448439e-08, 2.42957e-08, 2.444017e-08, 
    2.45183e-08, 2.342306e-08, 2.29273e-08, 2.426246e-08, 2.516358e-08,
  2.520569e-08, 2.515968e-08, 2.507914e-08, 2.484727e-08, 2.462373e-08, 
    2.445758e-08, 2.521113e-08, 2.449804e-08, 2.435206e-08, 2.455045e-08, 
    2.452773e-08, 2.371235e-08, 2.275908e-08, 2.423815e-08, 2.525118e-08,
  2.509917e-08, 2.497706e-08, 2.496243e-08, 2.469695e-08, 2.470193e-08, 
    2.497598e-08, 2.480467e-08, 2.504123e-08, 2.486507e-08, 2.464385e-08, 
    2.449071e-08, 2.413656e-08, 2.234716e-08, 2.31886e-08, 2.500754e-08,
  2.490684e-08, 2.495666e-08, 2.49138e-08, 2.479423e-08, 2.497232e-08, 
    2.507389e-08, 2.504576e-08, 2.488862e-08, 2.476685e-08, 2.490241e-08, 
    2.450981e-08, 2.461431e-08, 2.29132e-08, 2.27883e-08, 2.490875e-08,
  2.478832e-08, 2.480888e-08, 2.475757e-08, 2.48256e-08, 2.502764e-08, 
    2.506367e-08, 2.507669e-08, 2.50049e-08, 2.505799e-08, 2.513702e-08, 
    2.470061e-08, 2.47072e-08, 2.379414e-08, 2.220751e-08, 2.485952e-08,
  2.427356e-08, 2.442613e-08, 2.45145e-08, 2.478194e-08, 2.499833e-08, 
    2.51487e-08, 2.511845e-08, 2.507931e-08, 2.506636e-08, 2.542619e-08, 
    2.507984e-08, 2.457353e-08, 2.455859e-08, 2.260243e-08, 2.264758e-08,
  2.437175e-08, 2.44054e-08, 2.449319e-08, 2.472908e-08, 2.479828e-08, 
    2.479027e-08, 2.493196e-08, 2.509958e-08, 2.520697e-08, 2.501766e-08, 
    2.48695e-08, 2.443946e-08, 2.460735e-08, 2.371283e-08, 2.213226e-08,
  2.466259e-08, 2.471857e-08, 2.488665e-08, 2.483131e-08, 2.488389e-08, 
    2.469569e-08, 2.458745e-08, 2.490355e-08, 2.492298e-08, 2.481852e-08, 
    2.497346e-08, 2.476661e-08, 2.415774e-08, 2.400928e-08, 2.517464e-08,
  2.479793e-08, 2.469167e-08, 2.472193e-08, 2.46404e-08, 2.466569e-08, 
    2.449208e-08, 2.46676e-08, 2.479308e-08, 2.479333e-08, 2.501964e-08, 
    2.508939e-08, 2.486283e-08, 2.417546e-08, 2.401129e-08, 2.493681e-08,
  2.456042e-08, 2.447551e-08, 2.44378e-08, 2.440853e-08, 2.447372e-08, 
    2.434223e-08, 2.460867e-08, 2.477712e-08, 2.480678e-08, 2.520494e-08, 
    2.519373e-08, 2.501175e-08, 2.416202e-08, 2.433332e-08, 2.480019e-08,
  2.438331e-08, 2.429715e-08, 2.430163e-08, 2.430523e-08, 2.429844e-08, 
    2.473785e-08, 2.456047e-08, 2.455013e-08, 2.48143e-08, 2.541154e-08, 
    2.537886e-08, 2.501852e-08, 2.430811e-08, 2.395188e-08, 2.415013e-08,
  2.422438e-08, 2.414577e-08, 2.409613e-08, 2.413113e-08, 2.427612e-08, 
    2.432401e-08, 2.48315e-08, 2.455825e-08, 2.470731e-08, 2.551731e-08, 
    2.540415e-08, 2.49785e-08, 2.442383e-08, 2.434577e-08, 2.422088e-08,
  2.394407e-08, 2.391512e-08, 2.393672e-08, 2.410629e-08, 2.414258e-08, 
    2.447889e-08, 2.44867e-08, 2.472942e-08, 2.51286e-08, 2.561704e-08, 
    2.550146e-08, 2.482088e-08, 2.457727e-08, 2.43216e-08, 2.441727e-08,
  2.384079e-08, 2.393611e-08, 2.394751e-08, 2.406043e-08, 2.429092e-08, 
    2.434426e-08, 2.451185e-08, 2.449293e-08, 2.47923e-08, 2.562268e-08, 
    2.555977e-08, 2.456642e-08, 2.457089e-08, 2.474425e-08, 2.636578e-08,
  2.394073e-08, 2.396871e-08, 2.39052e-08, 2.413099e-08, 2.411025e-08, 
    2.417471e-08, 2.429335e-08, 2.459203e-08, 2.522221e-08, 2.596564e-08, 
    2.535197e-08, 2.418475e-08, 2.442777e-08, 2.427571e-08, 2.717353e-08,
  2.4094e-08, 2.402346e-08, 2.41323e-08, 2.429119e-08, 2.416424e-08, 
    2.416997e-08, 2.435416e-08, 2.476935e-08, 2.547719e-08, 2.594919e-08, 
    2.486423e-08, 2.388306e-08, 2.426867e-08, 2.389987e-08, 2.450866e-08,
  2.433811e-08, 2.425522e-08, 2.438165e-08, 2.441064e-08, 2.407152e-08, 
    2.413822e-08, 2.427247e-08, 2.472407e-08, 2.567891e-08, 2.571397e-08, 
    2.45982e-08, 2.394989e-08, 2.420042e-08, 2.44053e-08, 2.36693e-08,
  2.461485e-08, 2.459363e-08, 2.45329e-08, 2.449245e-08, 2.446323e-08, 
    2.437561e-08, 2.444344e-08, 2.428675e-08, 2.399754e-08, 2.437121e-08, 
    2.550075e-08, 2.570097e-08, 2.52069e-08, 2.448648e-08, 2.491704e-08,
  2.490353e-08, 2.495645e-08, 2.487971e-08, 2.471105e-08, 2.456045e-08, 
    2.4408e-08, 2.444805e-08, 2.430918e-08, 2.420515e-08, 2.480026e-08, 
    2.587043e-08, 2.586523e-08, 2.50786e-08, 2.445285e-08, 2.488872e-08,
  2.485299e-08, 2.494387e-08, 2.482642e-08, 2.472868e-08, 2.452068e-08, 
    2.442705e-08, 2.420367e-08, 2.410246e-08, 2.411746e-08, 2.508874e-08, 
    2.595175e-08, 2.583032e-08, 2.493021e-08, 2.451828e-08, 2.517231e-08,
  2.494273e-08, 2.499525e-08, 2.483739e-08, 2.461797e-08, 2.444658e-08, 
    2.436233e-08, 2.41758e-08, 2.371925e-08, 2.437763e-08, 2.535948e-08, 
    2.595227e-08, 2.588791e-08, 2.500344e-08, 2.450811e-08, 2.507275e-08,
  2.481828e-08, 2.486262e-08, 2.469687e-08, 2.45611e-08, 2.440462e-08, 
    2.419761e-08, 2.411539e-08, 2.389272e-08, 2.470969e-08, 2.51573e-08, 
    2.567794e-08, 2.612832e-08, 2.512938e-08, 2.447475e-08, 2.554519e-08,
  2.486187e-08, 2.487472e-08, 2.467713e-08, 2.437648e-08, 2.431775e-08, 
    2.419232e-08, 2.394185e-08, 2.392296e-08, 2.454449e-08, 2.454057e-08, 
    2.548233e-08, 2.642566e-08, 2.520166e-08, 2.434572e-08, 2.541775e-08,
  2.473625e-08, 2.482262e-08, 2.451267e-08, 2.399564e-08, 2.408441e-08, 
    2.408255e-08, 2.396481e-08, 2.379241e-08, 2.402481e-08, 2.445582e-08, 
    2.588734e-08, 2.681962e-08, 2.532421e-08, 2.440859e-08, 2.569069e-08,
  2.461959e-08, 2.481066e-08, 2.437837e-08, 2.37155e-08, 2.392961e-08, 
    2.405008e-08, 2.395555e-08, 2.385238e-08, 2.408479e-08, 2.469986e-08, 
    2.563973e-08, 2.678392e-08, 2.553162e-08, 2.430662e-08, 2.553686e-08,
  2.447416e-08, 2.48124e-08, 2.434382e-08, 2.328982e-08, 2.36592e-08, 
    2.391285e-08, 2.390285e-08, 2.393213e-08, 2.40516e-08, 2.403912e-08, 
    2.53184e-08, 2.715074e-08, 2.572076e-08, 2.444574e-08, 2.512611e-08,
  2.427073e-08, 2.463647e-08, 2.415667e-08, 2.295749e-08, 2.335408e-08, 
    2.378837e-08, 2.388307e-08, 2.395324e-08, 2.36058e-08, 2.339896e-08, 
    2.478691e-08, 2.702116e-08, 2.57759e-08, 2.429362e-08, 2.512916e-08,
  2.366457e-08, 2.337931e-08, 2.306964e-08, 2.329165e-08, 2.346733e-08, 
    2.363589e-08, 2.414103e-08, 2.457344e-08, 2.432033e-08, 2.35377e-08, 
    2.298107e-08, 2.5187e-08, 2.702881e-08, 2.548457e-08, 2.53257e-08,
  2.369744e-08, 2.339886e-08, 2.295246e-08, 2.318949e-08, 2.338711e-08, 
    2.347385e-08, 2.418408e-08, 2.47623e-08, 2.465275e-08, 2.352398e-08, 
    2.24664e-08, 2.487069e-08, 2.695616e-08, 2.560905e-08, 2.523427e-08,
  2.391856e-08, 2.355356e-08, 2.298516e-08, 2.305944e-08, 2.312125e-08, 
    2.294721e-08, 2.35146e-08, 2.439812e-08, 2.464364e-08, 2.330108e-08, 
    2.190207e-08, 2.441404e-08, 2.660518e-08, 2.558723e-08, 2.535022e-08,
  2.407611e-08, 2.387955e-08, 2.325983e-08, 2.31544e-08, 2.317718e-08, 
    2.363515e-08, 2.3298e-08, 2.430376e-08, 2.470477e-08, 2.30597e-08, 
    2.165071e-08, 2.392692e-08, 2.657752e-08, 2.534543e-08, 2.505415e-08,
  2.433485e-08, 2.428036e-08, 2.351978e-08, 2.328704e-08, 2.290634e-08, 
    2.27126e-08, 2.370204e-08, 2.391348e-08, 2.442176e-08, 2.261872e-08, 
    2.161578e-08, 2.372055e-08, 2.614561e-08, 2.537006e-08, 2.486309e-08,
  2.429717e-08, 2.438144e-08, 2.385582e-08, 2.371064e-08, 2.320944e-08, 
    2.288907e-08, 2.282956e-08, 2.353536e-08, 2.363513e-08, 2.237639e-08, 
    2.208603e-08, 2.345331e-08, 2.600093e-08, 2.533048e-08, 2.451664e-08,
  2.441288e-08, 2.454679e-08, 2.409712e-08, 2.393969e-08, 2.311571e-08, 
    2.260014e-08, 2.283229e-08, 2.324433e-08, 2.352826e-08, 2.303963e-08, 
    2.250942e-08, 2.329503e-08, 2.563544e-08, 2.515786e-08, 2.448837e-08,
  2.448376e-08, 2.45484e-08, 2.429453e-08, 2.423206e-08, 2.330641e-08, 
    2.277777e-08, 2.26729e-08, 2.316962e-08, 2.348493e-08, 2.352203e-08, 
    2.261011e-08, 2.314036e-08, 2.541741e-08, 2.50449e-08, 2.414207e-08,
  2.461939e-08, 2.46786e-08, 2.444086e-08, 2.414508e-08, 2.312125e-08, 
    2.267564e-08, 2.274366e-08, 2.304105e-08, 2.334265e-08, 2.33538e-08, 
    2.273806e-08, 2.294099e-08, 2.50318e-08, 2.488162e-08, 2.406592e-08,
  2.448428e-08, 2.435024e-08, 2.418904e-08, 2.389276e-08, 2.322836e-08, 
    2.296228e-08, 2.26063e-08, 2.259102e-08, 2.29572e-08, 2.318392e-08, 
    2.277721e-08, 2.294405e-08, 2.478313e-08, 2.471044e-08, 2.437399e-08,
  2.421327e-08, 2.433472e-08, 2.410716e-08, 2.417469e-08, 2.390961e-08, 
    2.343813e-08, 2.307871e-08, 2.350351e-08, 2.407376e-08, 2.301348e-08, 
    2.235514e-08, 2.293865e-08, 2.504098e-08, 2.499886e-08, 2.419537e-08,
  2.436173e-08, 2.446785e-08, 2.4015e-08, 2.424435e-08, 2.404521e-08, 
    2.352151e-08, 2.316091e-08, 2.322763e-08, 2.385865e-08, 2.294831e-08, 
    2.265135e-08, 2.297065e-08, 2.500852e-08, 2.493127e-08, 2.377852e-08,
  2.407112e-08, 2.434131e-08, 2.399955e-08, 2.396224e-08, 2.403734e-08, 
    2.357589e-08, 2.339475e-08, 2.324715e-08, 2.341114e-08, 2.300567e-08, 
    2.294715e-08, 2.297461e-08, 2.483988e-08, 2.483396e-08, 2.348326e-08,
  2.384734e-08, 2.430905e-08, 2.412092e-08, 2.399701e-08, 2.380655e-08, 
    2.383104e-08, 2.341525e-08, 2.316828e-08, 2.352586e-08, 2.268112e-08, 
    2.288828e-08, 2.288857e-08, 2.450913e-08, 2.457758e-08, 2.318071e-08,
  2.362021e-08, 2.402867e-08, 2.380398e-08, 2.347774e-08, 2.37012e-08, 
    2.322061e-08, 2.376928e-08, 2.318028e-08, 2.334131e-08, 2.259888e-08, 
    2.287535e-08, 2.302738e-08, 2.418974e-08, 2.459884e-08, 2.314938e-08,
  2.355572e-08, 2.39277e-08, 2.3944e-08, 2.383289e-08, 2.368396e-08, 
    2.393537e-08, 2.308955e-08, 2.351016e-08, 2.340607e-08, 2.2638e-08, 
    2.26821e-08, 2.288997e-08, 2.384116e-08, 2.455925e-08, 2.300834e-08,
  2.361954e-08, 2.357563e-08, 2.337488e-08, 2.29282e-08, 2.29005e-08, 
    2.265664e-08, 2.324426e-08, 2.324049e-08, 2.276394e-08, 2.224073e-08, 
    2.274743e-08, 2.295428e-08, 2.346581e-08, 2.459297e-08, 2.26032e-08,
  2.352496e-08, 2.340793e-08, 2.317004e-08, 2.292021e-08, 2.298232e-08, 
    2.306e-08, 2.339857e-08, 2.284757e-08, 2.274977e-08, 2.25307e-08, 
    2.252424e-08, 2.269277e-08, 2.318968e-08, 2.459537e-08, 2.247795e-08,
  2.357579e-08, 2.3313e-08, 2.270001e-08, 2.22328e-08, 2.230349e-08, 
    2.228478e-08, 2.271833e-08, 2.246831e-08, 2.283835e-08, 2.221091e-08, 
    2.234926e-08, 2.292362e-08, 2.299311e-08, 2.443832e-08, 2.259566e-08,
  2.325125e-08, 2.292122e-08, 2.234217e-08, 2.20821e-08, 2.215216e-08, 
    2.227428e-08, 2.271237e-08, 2.217487e-08, 2.24632e-08, 2.21826e-08, 
    2.241992e-08, 2.276112e-08, 2.292975e-08, 2.405994e-08, 2.390557e-08,
  2.308222e-08, 2.36171e-08, 2.375469e-08, 2.37864e-08, 2.309304e-08, 
    2.298309e-08, 2.363151e-08, 2.391592e-08, 2.343084e-08, 2.268621e-08, 
    2.286241e-08, 2.387029e-08, 2.410387e-08, 2.29185e-08, 2.342972e-08,
  2.326388e-08, 2.364098e-08, 2.382225e-08, 2.401851e-08, 2.336946e-08, 
    2.254563e-08, 2.344315e-08, 2.35074e-08, 2.379797e-08, 2.301009e-08, 
    2.292207e-08, 2.357389e-08, 2.394854e-08, 2.309303e-08, 2.380523e-08,
  2.339214e-08, 2.326798e-08, 2.387789e-08, 2.398623e-08, 2.383565e-08, 
    2.249007e-08, 2.296352e-08, 2.308781e-08, 2.36798e-08, 2.3163e-08, 
    2.299338e-08, 2.340986e-08, 2.39515e-08, 2.363695e-08, 2.403887e-08,
  2.324599e-08, 2.326913e-08, 2.37917e-08, 2.378821e-08, 2.386008e-08, 
    2.326244e-08, 2.257485e-08, 2.259903e-08, 2.351668e-08, 2.334763e-08, 
    2.292341e-08, 2.328543e-08, 2.357939e-08, 2.32423e-08, 2.398095e-08,
  2.340838e-08, 2.347939e-08, 2.312706e-08, 2.364603e-08, 2.341364e-08, 
    2.305892e-08, 2.312749e-08, 2.242265e-08, 2.32946e-08, 2.365479e-08, 
    2.292692e-08, 2.308573e-08, 2.356935e-08, 2.322063e-08, 2.339215e-08,
  2.352787e-08, 2.320768e-08, 2.326056e-08, 2.31246e-08, 2.278245e-08, 
    2.299144e-08, 2.262168e-08, 2.257301e-08, 2.330675e-08, 2.290075e-08, 
    2.248504e-08, 2.282855e-08, 2.321524e-08, 2.338989e-08, 2.350367e-08,
  2.363837e-08, 2.353259e-08, 2.315236e-08, 2.256926e-08, 2.291499e-08, 
    2.249675e-08, 2.234984e-08, 2.262487e-08, 2.235048e-08, 2.205484e-08, 
    2.277013e-08, 2.299701e-08, 2.311389e-08, 2.350685e-08, 2.321251e-08,
  2.36427e-08, 2.350582e-08, 2.298355e-08, 2.274155e-08, 2.21165e-08, 
    2.186358e-08, 2.247448e-08, 2.276387e-08, 2.214741e-08, 2.326047e-08, 
    2.335856e-08, 2.270743e-08, 2.279764e-08, 2.367039e-08, 2.270574e-08,
  2.339167e-08, 2.348723e-08, 2.31656e-08, 2.245045e-08, 2.225363e-08, 
    2.195526e-08, 2.21274e-08, 2.139198e-08, 2.290866e-08, 2.31945e-08, 
    2.303268e-08, 2.296888e-08, 2.301212e-08, 2.378769e-08, 2.233929e-08,
  2.285025e-08, 2.308401e-08, 2.302282e-08, 2.288283e-08, 2.25159e-08, 
    2.262209e-08, 2.256237e-08, 2.220288e-08, 2.159655e-08, 2.334781e-08, 
    2.399791e-08, 2.309458e-08, 2.252855e-08, 2.37604e-08, 2.254026e-08,
  2.344795e-08, 2.3106e-08, 2.345698e-08, 2.379235e-08, 2.32638e-08, 
    2.23825e-08, 2.274033e-08, 2.384867e-08, 2.260391e-08, 2.316206e-08, 
    2.393966e-08, 2.395386e-08, 2.383215e-08, 2.404787e-08, 2.426511e-08,
  2.399161e-08, 2.319361e-08, 2.373387e-08, 2.364513e-08, 2.310348e-08, 
    2.27555e-08, 2.301632e-08, 2.310336e-08, 2.343278e-08, 2.354958e-08, 
    2.389439e-08, 2.405192e-08, 2.410861e-08, 2.460927e-08, 2.468555e-08,
  2.355905e-08, 2.306133e-08, 2.37007e-08, 2.372667e-08, 2.312253e-08, 
    2.247915e-08, 2.265071e-08, 2.316044e-08, 2.337571e-08, 2.3514e-08, 
    2.386294e-08, 2.425634e-08, 2.454676e-08, 2.500001e-08, 2.495686e-08,
  2.363593e-08, 2.33931e-08, 2.332523e-08, 2.380828e-08, 2.309594e-08, 
    2.229393e-08, 2.253411e-08, 2.343331e-08, 2.325934e-08, 2.309628e-08, 
    2.390169e-08, 2.43583e-08, 2.478799e-08, 2.524065e-08, 2.520383e-08,
  2.418227e-08, 2.323994e-08, 2.29154e-08, 2.314452e-08, 2.307355e-08, 
    2.271942e-08, 2.287053e-08, 2.285507e-08, 2.324424e-08, 2.337213e-08, 
    2.389333e-08, 2.399204e-08, 2.441638e-08, 2.470328e-08, 2.490186e-08,
  2.402083e-08, 2.332045e-08, 2.334562e-08, 2.304974e-08, 2.296197e-08, 
    2.247768e-08, 2.11377e-08, 2.304506e-08, 2.408417e-08, 2.375955e-08, 
    2.375987e-08, 2.382502e-08, 2.431309e-08, 2.488756e-08, 2.514043e-08,
  2.348994e-08, 2.354715e-08, 2.292005e-08, 2.311685e-08, 2.272199e-08, 
    2.275803e-08, 2.269718e-08, 2.365111e-08, 2.326051e-08, 2.294179e-08, 
    2.332298e-08, 2.3762e-08, 2.426719e-08, 2.48264e-08, 2.49976e-08,
  2.179506e-08, 2.314115e-08, 2.325115e-08, 2.301101e-08, 2.247374e-08, 
    2.240848e-08, 2.246883e-08, 2.305435e-08, 2.237508e-08, 2.276914e-08, 
    2.330945e-08, 2.368725e-08, 2.40975e-08, 2.453893e-08, 2.445634e-08,
  2.027348e-08, 2.162238e-08, 2.27702e-08, 2.34378e-08, 2.343499e-08, 
    2.299526e-08, 2.269375e-08, 2.25023e-08, 2.297317e-08, 2.275943e-08, 
    2.31025e-08, 2.349372e-08, 2.387206e-08, 2.397558e-08, 2.373197e-08,
  1.986083e-08, 2.057496e-08, 2.143646e-08, 2.256026e-08, 2.356966e-08, 
    2.384808e-08, 2.358478e-08, 2.226334e-08, 2.242895e-08, 2.371172e-08, 
    2.423708e-08, 2.376095e-08, 2.337783e-08, 2.351598e-08, 2.350507e-08,
  2.398788e-08, 2.31603e-08, 2.334838e-08, 2.355245e-08, 2.237252e-08, 
    2.261422e-08, 2.329839e-08, 2.302483e-08, 2.282977e-08, 2.3433e-08, 
    2.388412e-08, 2.331606e-08, 2.378142e-08, 2.51708e-08, 2.56303e-08,
  2.414542e-08, 2.331272e-08, 2.351676e-08, 2.305528e-08, 2.233292e-08, 
    2.265372e-08, 2.256135e-08, 2.319602e-08, 2.333578e-08, 2.433947e-08, 
    2.421997e-08, 2.396124e-08, 2.4377e-08, 2.514896e-08, 2.532153e-08,
  2.347113e-08, 2.354425e-08, 2.351625e-08, 2.257216e-08, 2.181486e-08, 
    2.124387e-08, 2.172082e-08, 2.303156e-08, 2.397675e-08, 2.453732e-08, 
    2.391898e-08, 2.456118e-08, 2.48487e-08, 2.522831e-08, 2.454558e-08,
  2.371366e-08, 2.36313e-08, 2.333352e-08, 2.229265e-08, 2.098187e-08, 
    2.140193e-08, 2.22558e-08, 2.347727e-08, 2.441969e-08, 2.434565e-08, 
    2.464809e-08, 2.47567e-08, 2.489282e-08, 2.486765e-08, 2.402231e-08,
  2.382003e-08, 2.316428e-08, 2.317643e-08, 2.248293e-08, 2.164306e-08, 
    2.143295e-08, 2.405672e-08, 2.573833e-08, 2.34934e-08, 2.353407e-08, 
    2.436517e-08, 2.487138e-08, 2.500494e-08, 2.459786e-08, 2.391783e-08,
  2.375185e-08, 2.312114e-08, 2.31427e-08, 2.234606e-08, 2.119336e-08, 
    2.111119e-08, 2.305087e-08, 2.32857e-08, 2.377643e-08, 2.618015e-08, 
    2.658918e-08, 2.563023e-08, 2.490419e-08, 2.462052e-08, 2.421432e-08,
  2.370131e-08, 2.307497e-08, 2.314389e-08, 2.234708e-08, 2.172618e-08, 
    2.217448e-08, 2.415143e-08, 2.526221e-08, 2.630486e-08, 2.848004e-08, 
    2.656958e-08, 2.528152e-08, 2.500811e-08, 2.485545e-08, 2.453144e-08,
  2.324961e-08, 2.314536e-08, 2.290727e-08, 2.246073e-08, 2.241917e-08, 
    2.330969e-08, 2.455112e-08, 2.521377e-08, 2.624846e-08, 2.713407e-08, 
    2.530903e-08, 2.513686e-08, 2.512906e-08, 2.502058e-08, 2.501968e-08,
  2.222839e-08, 2.285532e-08, 2.292243e-08, 2.292622e-08, 2.307987e-08, 
    2.366505e-08, 2.471472e-08, 2.507596e-08, 2.51678e-08, 2.503605e-08, 
    2.497369e-08, 2.51602e-08, 2.520387e-08, 2.516109e-08, 2.542909e-08,
  2.160797e-08, 2.245215e-08, 2.285946e-08, 2.336201e-08, 2.339571e-08, 
    2.36046e-08, 2.347021e-08, 2.310646e-08, 2.394015e-08, 2.48211e-08, 
    2.49914e-08, 2.499509e-08, 2.500485e-08, 2.516058e-08, 2.55692e-08,
  2.32188e-08, 2.323367e-08, 2.323224e-08, 2.324374e-08, 2.364837e-08, 
    2.353243e-08, 2.397279e-08, 2.37884e-08, 2.331614e-08, 2.283517e-08, 
    2.343205e-08, 2.375582e-08, 2.458205e-08, 2.523968e-08, 2.496298e-08,
  2.294636e-08, 2.34906e-08, 2.3478e-08, 2.360254e-08, 2.29436e-08, 
    2.279116e-08, 2.252188e-08, 2.311115e-08, 2.303382e-08, 2.33147e-08, 
    2.385713e-08, 2.394601e-08, 2.496882e-08, 2.51963e-08, 2.475867e-08,
  2.29899e-08, 2.348332e-08, 2.363562e-08, 2.339185e-08, 2.240506e-08, 
    2.044752e-08, 2.212228e-08, 2.315585e-08, 2.298565e-08, 2.352336e-08, 
    2.373573e-08, 2.442809e-08, 2.544815e-08, 2.533318e-08, 2.423445e-08,
  2.302669e-08, 2.347446e-08, 2.343031e-08, 2.284919e-08, 2.100621e-08, 
    2.010574e-08, 2.226227e-08, 2.270575e-08, 2.360381e-08, 2.383347e-08, 
    2.419526e-08, 2.473695e-08, 2.510055e-08, 2.458189e-08, 2.351831e-08,
  2.342165e-08, 2.359052e-08, 2.334213e-08, 2.243929e-08, 2.093405e-08, 
    2.029187e-08, 2.188468e-08, 2.567953e-08, 2.360281e-08, 2.28009e-08, 
    2.410802e-08, 2.481433e-08, 2.477403e-08, 2.396444e-08, 2.338702e-08,
  2.34575e-08, 2.34551e-08, 2.307541e-08, 2.20579e-08, 2.076736e-08, 
    2.126523e-08, 2.42304e-08, 2.16272e-08, 2.251681e-08, 2.511598e-08, 
    2.48409e-08, 2.497999e-08, 2.422354e-08, 2.350363e-08, 2.31655e-08,
  2.354952e-08, 2.331014e-08, 2.279248e-08, 2.178558e-08, 2.091516e-08, 
    2.224648e-08, 2.495697e-08, 2.218711e-08, 2.458017e-08, 2.849898e-08, 
    2.539204e-08, 2.49614e-08, 2.38183e-08, 2.320891e-08, 2.277346e-08,
  2.367561e-08, 2.304233e-08, 2.228531e-08, 2.141161e-08, 2.148696e-08, 
    2.388157e-08, 2.463909e-08, 2.290885e-08, 2.681088e-08, 2.845739e-08, 
    2.538882e-08, 2.460216e-08, 2.37021e-08, 2.307684e-08, 2.270773e-08,
  2.336058e-08, 2.252894e-08, 2.19132e-08, 2.180127e-08, 2.319326e-08, 
    2.502754e-08, 2.577511e-08, 2.557232e-08, 2.810058e-08, 2.731191e-08, 
    2.499318e-08, 2.462639e-08, 2.375731e-08, 2.315898e-08, 2.289538e-08,
  2.277342e-08, 2.240482e-08, 2.261304e-08, 2.323796e-08, 2.445758e-08, 
    2.586349e-08, 2.623904e-08, 2.661553e-08, 2.719005e-08, 2.649671e-08, 
    2.516203e-08, 2.465267e-08, 2.403321e-08, 2.365564e-08, 2.320456e-08,
  2.256262e-08, 2.285435e-08, 2.340391e-08, 2.324484e-08, 2.34761e-08, 
    2.492368e-08, 2.509131e-08, 2.401706e-08, 2.369607e-08, 2.395043e-08, 
    2.469135e-08, 2.510759e-08, 2.488391e-08, 2.482116e-08, 2.519089e-08,
  2.221422e-08, 2.276449e-08, 2.328414e-08, 2.364543e-08, 2.39493e-08, 
    2.366443e-08, 2.310889e-08, 2.365055e-08, 2.383353e-08, 2.45711e-08, 
    2.505858e-08, 2.500618e-08, 2.461866e-08, 2.470556e-08, 2.534425e-08,
  2.211984e-08, 2.269753e-08, 2.31797e-08, 2.354281e-08, 2.395779e-08, 
    2.304185e-08, 2.231114e-08, 2.278971e-08, 2.422051e-08, 2.462431e-08, 
    2.504591e-08, 2.502861e-08, 2.491591e-08, 2.525123e-08, 2.554381e-08,
  2.18839e-08, 2.204877e-08, 2.271505e-08, 2.361731e-08, 2.355637e-08, 
    2.200147e-08, 2.33271e-08, 2.297056e-08, 2.34594e-08, 2.476042e-08, 
    2.48945e-08, 2.497224e-08, 2.528131e-08, 2.534448e-08, 2.477142e-08,
  2.19944e-08, 2.210393e-08, 2.252026e-08, 2.364238e-08, 2.338092e-08, 
    2.204325e-08, 2.331612e-08, 2.417106e-08, 2.444514e-08, 2.426208e-08, 
    2.481218e-08, 2.500691e-08, 2.517007e-08, 2.501781e-08, 2.472682e-08,
  2.218572e-08, 2.210544e-08, 2.243115e-08, 2.348639e-08, 2.345896e-08, 
    2.170742e-08, 2.268769e-08, 2.334258e-08, 2.466354e-08, 2.419433e-08, 
    2.479181e-08, 2.489967e-08, 2.489465e-08, 2.455043e-08, 2.463768e-08,
  2.25594e-08, 2.232525e-08, 2.252835e-08, 2.342367e-08, 2.318421e-08, 
    2.15374e-08, 2.176559e-08, 2.401653e-08, 2.429419e-08, 2.496305e-08, 
    2.46674e-08, 2.472555e-08, 2.441267e-08, 2.42785e-08, 2.463569e-08,
  2.258708e-08, 2.247965e-08, 2.276647e-08, 2.364135e-08, 2.320092e-08, 
    2.109145e-08, 2.167238e-08, 2.300657e-08, 2.385516e-08, 2.537188e-08, 
    2.449896e-08, 2.452783e-08, 2.415702e-08, 2.414259e-08, 2.462361e-08,
  2.29413e-08, 2.289622e-08, 2.289094e-08, 2.338917e-08, 2.284379e-08, 
    2.126629e-08, 2.221512e-08, 2.225778e-08, 2.399972e-08, 2.59735e-08, 
    2.464961e-08, 2.446663e-08, 2.404947e-08, 2.397241e-08, 2.443432e-08,
  2.316353e-08, 2.301158e-08, 2.307948e-08, 2.341999e-08, 2.274753e-08, 
    2.154294e-08, 2.26224e-08, 2.2344e-08, 2.443045e-08, 2.661864e-08, 
    2.470443e-08, 2.427599e-08, 2.37588e-08, 2.382376e-08, 2.423273e-08,
  2.229381e-08, 2.234098e-08, 2.294005e-08, 2.262723e-08, 2.263653e-08, 
    2.436106e-08, 2.406403e-08, 2.412991e-08, 2.363492e-08, 2.311421e-08, 
    2.345406e-08, 2.393746e-08, 2.469664e-08, 2.531095e-08, 2.493826e-08,
  2.263483e-08, 2.255344e-08, 2.34496e-08, 2.2951e-08, 2.309538e-08, 
    2.375826e-08, 2.456814e-08, 2.373163e-08, 2.355283e-08, 2.361116e-08, 
    2.375192e-08, 2.410259e-08, 2.456248e-08, 2.490654e-08, 2.568519e-08,
  2.238539e-08, 2.273374e-08, 2.342206e-08, 2.284875e-08, 2.327723e-08, 
    2.429528e-08, 2.243437e-08, 2.312482e-08, 2.379615e-08, 2.379087e-08, 
    2.39449e-08, 2.428339e-08, 2.461947e-08, 2.527014e-08, 2.628718e-08,
  2.194692e-08, 2.288029e-08, 2.331939e-08, 2.284201e-08, 2.303761e-08, 
    2.36179e-08, 2.357911e-08, 2.266644e-08, 2.402527e-08, 2.439208e-08, 
    2.435502e-08, 2.438113e-08, 2.46241e-08, 2.553245e-08, 2.654864e-08,
  2.163218e-08, 2.26259e-08, 2.29842e-08, 2.263357e-08, 2.306215e-08, 
    2.361781e-08, 2.354035e-08, 2.516284e-08, 2.497575e-08, 2.339166e-08, 
    2.415588e-08, 2.42755e-08, 2.449816e-08, 2.562671e-08, 2.672858e-08,
  2.132186e-08, 2.230333e-08, 2.292302e-08, 2.300021e-08, 2.335967e-08, 
    2.424021e-08, 2.498927e-08, 2.479897e-08, 2.329009e-08, 2.330727e-08, 
    2.534225e-08, 2.428523e-08, 2.465178e-08, 2.530229e-08, 2.635997e-08,
  2.129164e-08, 2.226193e-08, 2.294209e-08, 2.34621e-08, 2.409146e-08, 
    2.456393e-08, 2.472871e-08, 2.462476e-08, 2.42872e-08, 2.50768e-08, 
    2.517666e-08, 2.437328e-08, 2.470228e-08, 2.507911e-08, 2.575093e-08,
  2.128249e-08, 2.22063e-08, 2.297017e-08, 2.3445e-08, 2.403893e-08, 
    2.428306e-08, 2.446851e-08, 2.482853e-08, 2.503142e-08, 2.521387e-08, 
    2.509108e-08, 2.457756e-08, 2.500644e-08, 2.501272e-08, 2.53213e-08,
  2.153567e-08, 2.223852e-08, 2.283917e-08, 2.33985e-08, 2.405133e-08, 
    2.357372e-08, 2.379262e-08, 2.451404e-08, 2.386555e-08, 2.499987e-08, 
    2.428245e-08, 2.459695e-08, 2.507818e-08, 2.489131e-08, 2.493352e-08,
  2.193743e-08, 2.222311e-08, 2.27293e-08, 2.313007e-08, 2.343691e-08, 
    2.292493e-08, 2.329793e-08, 2.337748e-08, 2.337093e-08, 2.414862e-08, 
    2.339272e-08, 2.51953e-08, 2.527579e-08, 2.50325e-08, 2.47825e-08,
  2.167227e-08, 2.131942e-08, 2.154774e-08, 2.188927e-08, 2.184285e-08, 
    2.207016e-08, 2.271721e-08, 2.310248e-08, 2.316627e-08, 2.366402e-08, 
    2.473137e-08, 2.323644e-08, 2.131738e-08, 1.944742e-08, 2.090262e-08,
  2.156209e-08, 2.132927e-08, 2.1664e-08, 2.168408e-08, 2.170601e-08, 
    2.17715e-08, 2.228632e-08, 2.311794e-08, 2.356971e-08, 2.429696e-08, 
    2.474834e-08, 2.272914e-08, 2.082347e-08, 2.07465e-08, 2.37499e-08,
  2.17355e-08, 2.129978e-08, 2.182972e-08, 2.17977e-08, 2.158449e-08, 
    2.185875e-08, 2.2146e-08, 2.253176e-08, 2.330611e-08, 2.370247e-08, 
    2.43089e-08, 2.270586e-08, 2.208598e-08, 2.316968e-08, 2.438827e-08,
  2.166744e-08, 2.139906e-08, 2.192901e-08, 2.17063e-08, 2.102787e-08, 
    2.168412e-08, 2.34758e-08, 2.264397e-08, 2.361078e-08, 2.437355e-08, 
    2.465957e-08, 2.298336e-08, 2.273738e-08, 2.360668e-08, 2.430624e-08,
  2.158661e-08, 2.146945e-08, 2.206137e-08, 2.190735e-08, 2.150012e-08, 
    2.32078e-08, 2.32899e-08, 2.422296e-08, 2.485794e-08, 2.254463e-08, 
    2.36069e-08, 2.332836e-08, 2.322843e-08, 2.352997e-08, 2.430582e-08,
  2.152759e-08, 2.171234e-08, 2.209233e-08, 2.18596e-08, 2.154358e-08, 
    2.318115e-08, 2.344043e-08, 2.333783e-08, 2.218356e-08, 2.131028e-08, 
    2.583826e-08, 2.456046e-08, 2.380641e-08, 2.357874e-08, 2.444318e-08,
  2.157937e-08, 2.160158e-08, 2.206476e-08, 2.198474e-08, 2.195855e-08, 
    2.306422e-08, 2.336647e-08, 2.371902e-08, 2.244552e-08, 2.344187e-08, 
    2.586225e-08, 2.502334e-08, 2.39923e-08, 2.396242e-08, 2.44798e-08,
  2.153767e-08, 2.179904e-08, 2.217473e-08, 2.212675e-08, 2.19585e-08, 
    2.292133e-08, 2.305401e-08, 2.351832e-08, 2.270378e-08, 2.398915e-08, 
    2.641886e-08, 2.545861e-08, 2.478756e-08, 2.42523e-08, 2.467177e-08,
  2.144941e-08, 2.175713e-08, 2.231188e-08, 2.236785e-08, 2.236281e-08, 
    2.302098e-08, 2.329099e-08, 2.373605e-08, 2.32556e-08, 2.260155e-08, 
    2.434171e-08, 2.522097e-08, 2.449136e-08, 2.481381e-08, 2.43126e-08,
  2.121311e-08, 2.19923e-08, 2.262679e-08, 2.285059e-08, 2.264306e-08, 
    2.310745e-08, 2.334969e-08, 2.365783e-08, 2.116372e-08, 1.89533e-08, 
    2.46216e-08, 2.752873e-08, 2.574211e-08, 2.507695e-08, 2.476751e-08,
  2.491216e-08, 2.397285e-08, 2.29885e-08, 2.18551e-08, 2.206917e-08, 
    2.213096e-08, 2.338897e-08, 2.368352e-08, 2.295667e-08, 2.12222e-08, 
    1.992945e-08, 1.863476e-08, 1.994009e-08, 2.246993e-08, 2.501407e-08,
  2.481321e-08, 2.393993e-08, 2.251164e-08, 2.169516e-08, 2.199817e-08, 
    2.220638e-08, 2.310721e-08, 2.377909e-08, 2.340632e-08, 2.236234e-08, 
    2.02801e-08, 1.855789e-08, 2.169979e-08, 2.747324e-08, 2.856778e-08,
  2.49745e-08, 2.380588e-08, 2.245014e-08, 2.179438e-08, 2.189863e-08, 
    2.263596e-08, 2.289356e-08, 2.234182e-08, 2.301012e-08, 2.182995e-08, 
    1.982555e-08, 1.868373e-08, 2.290457e-08, 2.779161e-08, 2.920072e-08,
  2.506991e-08, 2.400594e-08, 2.232437e-08, 2.179006e-08, 2.168425e-08, 
    2.095958e-08, 2.230922e-08, 2.226347e-08, 2.30809e-08, 2.249317e-08, 
    2.033793e-08, 1.837657e-08, 2.188412e-08, 2.534049e-08, 2.719551e-08,
  2.506545e-08, 2.379302e-08, 2.226482e-08, 2.175575e-08, 2.171055e-08, 
    2.161417e-08, 2.23823e-08, 2.427544e-08, 2.496641e-08, 2.059988e-08, 
    1.895514e-08, 1.783164e-08, 2.092086e-08, 2.379464e-08, 2.528095e-08,
  2.485019e-08, 2.381274e-08, 2.230625e-08, 2.171255e-08, 2.125127e-08, 
    2.155e-08, 2.272036e-08, 2.285768e-08, 2.037394e-08, 1.736546e-08, 
    2.30426e-08, 1.985478e-08, 2.071753e-08, 2.2911e-08, 2.49261e-08,
  2.433087e-08, 2.34944e-08, 2.22541e-08, 2.169288e-08, 2.13063e-08, 
    2.154277e-08, 2.252326e-08, 2.364481e-08, 2.08313e-08, 2.145803e-08, 
    2.366929e-08, 2.123932e-08, 2.101989e-08, 2.249299e-08, 2.470868e-08,
  2.374592e-08, 2.327659e-08, 2.237905e-08, 2.172784e-08, 2.092689e-08, 
    2.112484e-08, 2.232245e-08, 2.316021e-08, 2.084838e-08, 2.168732e-08, 
    2.414848e-08, 2.294457e-08, 2.24908e-08, 2.31314e-08, 2.42634e-08,
  2.313607e-08, 2.280475e-08, 2.224352e-08, 2.177165e-08, 2.130419e-08, 
    2.1307e-08, 2.214498e-08, 2.346802e-08, 2.155189e-08, 2.08984e-08, 
    2.262076e-08, 2.28703e-08, 2.285852e-08, 2.322993e-08, 2.426778e-08,
  2.261113e-08, 2.248491e-08, 2.216938e-08, 2.165384e-08, 2.101506e-08, 
    2.10376e-08, 2.169277e-08, 2.278149e-08, 2.113335e-08, 1.916606e-08, 
    2.240304e-08, 2.569613e-08, 2.449149e-08, 2.404901e-08, 2.473077e-08,
  2.311208e-08, 2.404459e-08, 2.55097e-08, 2.576595e-08, 2.445639e-08, 
    2.290982e-08, 2.249461e-08, 2.171411e-08, 2.093108e-08, 2.105481e-08, 
    2.197841e-08, 2.289161e-08, 2.34282e-08, 2.362005e-08, 2.44647e-08,
  2.313003e-08, 2.395915e-08, 2.518596e-08, 2.549482e-08, 2.477796e-08, 
    2.334943e-08, 2.20826e-08, 2.232828e-08, 2.117802e-08, 2.148671e-08, 
    2.176563e-08, 2.262912e-08, 2.402263e-08, 2.391821e-08, 2.440314e-08,
  2.288895e-08, 2.375008e-08, 2.477465e-08, 2.531618e-08, 2.500934e-08, 
    2.371085e-08, 2.265478e-08, 2.181487e-08, 2.203052e-08, 2.122948e-08, 
    2.091189e-08, 2.291662e-08, 2.516862e-08, 2.535643e-08, 2.45562e-08,
  2.267513e-08, 2.366169e-08, 2.447266e-08, 2.492876e-08, 2.512321e-08, 
    2.345977e-08, 2.262919e-08, 2.232023e-08, 2.161013e-08, 2.097319e-08, 
    2.092392e-08, 2.321461e-08, 2.549049e-08, 2.579186e-08, 2.512757e-08,
  2.261949e-08, 2.324898e-08, 2.439638e-08, 2.441367e-08, 2.51911e-08, 
    2.385933e-08, 2.232092e-08, 2.297835e-08, 2.263619e-08, 2.038853e-08, 
    1.956504e-08, 2.236069e-08, 2.525076e-08, 2.548365e-08, 2.373765e-08,
  2.287522e-08, 2.339113e-08, 2.415267e-08, 2.43553e-08, 2.46035e-08, 
    2.391419e-08, 2.237305e-08, 2.230741e-08, 2.162997e-08, 1.890389e-08, 
    2.013127e-08, 2.241547e-08, 2.448855e-08, 2.586362e-08, 2.466908e-08,
  2.285721e-08, 2.342953e-08, 2.41457e-08, 2.420123e-08, 2.441594e-08, 
    2.394601e-08, 2.259301e-08, 2.22453e-08, 2.153561e-08, 1.992561e-08, 
    2.080688e-08, 2.178935e-08, 2.435719e-08, 2.60124e-08, 2.562088e-08,
  2.316045e-08, 2.383007e-08, 2.417256e-08, 2.448819e-08, 2.374743e-08, 
    2.386431e-08, 2.269982e-08, 2.234252e-08, 2.166375e-08, 2.020765e-08, 
    2.058611e-08, 2.144381e-08, 2.316322e-08, 2.548225e-08, 2.575437e-08,
  2.390324e-08, 2.417508e-08, 2.440982e-08, 2.449547e-08, 2.416457e-08, 
    2.384009e-08, 2.289409e-08, 2.249976e-08, 2.209009e-08, 2.04633e-08, 
    2.095251e-08, 2.150323e-08, 2.271256e-08, 2.448018e-08, 2.489803e-08,
  2.430573e-08, 2.49151e-08, 2.500841e-08, 2.495176e-08, 2.379594e-08, 
    2.404286e-08, 2.307753e-08, 2.256503e-08, 2.248731e-08, 2.048175e-08, 
    2.065952e-08, 2.204533e-08, 2.254329e-08, 2.33604e-08, 2.389538e-08,
  2.498395e-08, 2.446387e-08, 2.323569e-08, 2.344945e-08, 2.392646e-08, 
    2.324067e-08, 2.334693e-08, 2.247239e-08, 2.209758e-08, 2.16351e-08, 
    2.140862e-08, 2.144516e-08, 2.076206e-08, 1.915255e-08, 2.086744e-08,
  2.48277e-08, 2.429067e-08, 2.325429e-08, 2.310595e-08, 2.375809e-08, 
    2.409154e-08, 2.23428e-08, 2.274058e-08, 2.174587e-08, 2.138693e-08, 
    2.154567e-08, 2.178255e-08, 2.119773e-08, 1.984916e-08, 2.231141e-08,
  2.462134e-08, 2.402817e-08, 2.315632e-08, 2.311728e-08, 2.322156e-08, 
    2.409218e-08, 2.374355e-08, 2.220439e-08, 2.173764e-08, 2.181364e-08, 
    2.183819e-08, 2.198723e-08, 2.181302e-08, 2.078788e-08, 2.283006e-08,
  2.427524e-08, 2.368545e-08, 2.306754e-08, 2.278738e-08, 2.308837e-08, 
    2.376328e-08, 2.391818e-08, 2.325209e-08, 2.214299e-08, 2.162892e-08, 
    2.184018e-08, 2.205054e-08, 2.210892e-08, 2.150163e-08, 2.291577e-08,
  2.419048e-08, 2.362346e-08, 2.303812e-08, 2.269373e-08, 2.28235e-08, 
    2.348329e-08, 2.425437e-08, 2.395079e-08, 2.295085e-08, 2.197354e-08, 
    2.168681e-08, 2.192742e-08, 2.198247e-08, 2.172139e-08, 2.290083e-08,
  2.411504e-08, 2.351913e-08, 2.303228e-08, 2.25399e-08, 2.273339e-08, 
    2.329397e-08, 2.416682e-08, 2.394355e-08, 2.284016e-08, 2.2292e-08, 
    2.143253e-08, 2.155381e-08, 2.167366e-08, 2.153537e-08, 2.245397e-08,
  2.448067e-08, 2.382394e-08, 2.328846e-08, 2.276964e-08, 2.251796e-08, 
    2.31151e-08, 2.366659e-08, 2.400088e-08, 2.30121e-08, 2.240177e-08, 
    2.167912e-08, 2.147231e-08, 2.143612e-08, 2.111202e-08, 2.190555e-08,
  2.503574e-08, 2.445716e-08, 2.403278e-08, 2.346215e-08, 2.304109e-08, 
    2.299428e-08, 2.372338e-08, 2.410311e-08, 2.356948e-08, 2.281052e-08, 
    2.180802e-08, 2.132411e-08, 2.151655e-08, 2.120239e-08, 2.151438e-08,
  2.478364e-08, 2.454808e-08, 2.413944e-08, 2.35729e-08, 2.313938e-08, 
    2.302026e-08, 2.325457e-08, 2.380602e-08, 2.373397e-08, 2.343748e-08, 
    2.23024e-08, 2.144504e-08, 2.132386e-08, 2.16878e-08, 2.134906e-08,
  2.393551e-08, 2.390052e-08, 2.373282e-08, 2.354896e-08, 2.307847e-08, 
    2.299784e-08, 2.30452e-08, 2.346975e-08, 2.374849e-08, 2.383158e-08, 
    2.312047e-08, 2.182043e-08, 2.13286e-08, 2.182393e-08, 2.193316e-08,
  2.611537e-08, 2.620839e-08, 2.615031e-08, 2.564341e-08, 2.479694e-08, 
    2.372291e-08, 2.440451e-08, 2.432072e-08, 2.380081e-08, 2.280951e-08, 
    2.2003e-08, 2.184015e-08, 2.226449e-08, 2.237874e-08, 2.08184e-08,
  2.589372e-08, 2.590452e-08, 2.583389e-08, 2.56006e-08, 2.459496e-08, 
    2.429987e-08, 2.392601e-08, 2.389425e-08, 2.346252e-08, 2.284083e-08, 
    2.194434e-08, 2.165345e-08, 2.200991e-08, 2.210418e-08, 2.061053e-08,
  2.539682e-08, 2.550028e-08, 2.574993e-08, 2.53841e-08, 2.543696e-08, 
    2.413074e-08, 2.404358e-08, 2.393567e-08, 2.352468e-08, 2.30603e-08, 
    2.214062e-08, 2.168505e-08, 2.197534e-08, 2.223616e-08, 2.045392e-08,
  2.443918e-08, 2.482422e-08, 2.521417e-08, 2.525691e-08, 2.508294e-08, 
    2.438635e-08, 2.368151e-08, 2.37256e-08, 2.338542e-08, 2.320175e-08, 
    2.237232e-08, 2.171143e-08, 2.192847e-08, 2.238405e-08, 2.079299e-08,
  2.498277e-08, 2.519699e-08, 2.529775e-08, 2.551796e-08, 2.500147e-08, 
    2.479555e-08, 2.388912e-08, 2.355115e-08, 2.292586e-08, 2.319679e-08, 
    2.282186e-08, 2.202323e-08, 2.197201e-08, 2.240675e-08, 2.114959e-08,
  2.45693e-08, 2.530706e-08, 2.525868e-08, 2.554856e-08, 2.52273e-08, 
    2.455712e-08, 2.433819e-08, 2.368108e-08, 2.304719e-08, 2.303326e-08, 
    2.278567e-08, 2.240489e-08, 2.207484e-08, 2.25611e-08, 2.178348e-08,
  2.452085e-08, 2.541504e-08, 2.553558e-08, 2.583615e-08, 2.545218e-08, 
    2.475632e-08, 2.403458e-08, 2.387628e-08, 2.329137e-08, 2.31999e-08, 
    2.277078e-08, 2.248142e-08, 2.209913e-08, 2.225816e-08, 2.225611e-08,
  2.523652e-08, 2.584986e-08, 2.604433e-08, 2.628173e-08, 2.593701e-08, 
    2.531126e-08, 2.432455e-08, 2.371436e-08, 2.341672e-08, 2.315545e-08, 
    2.306317e-08, 2.267467e-08, 2.225429e-08, 2.213615e-08, 2.220052e-08,
  2.262495e-08, 2.458184e-08, 2.577425e-08, 2.660508e-08, 2.614321e-08, 
    2.582335e-08, 2.510317e-08, 2.420717e-08, 2.361164e-08, 2.334075e-08, 
    2.303326e-08, 2.287563e-08, 2.224493e-08, 2.202809e-08, 2.187928e-08,
  2.048123e-08, 2.209784e-08, 2.372378e-08, 2.509322e-08, 2.532724e-08, 
    2.55627e-08, 2.568753e-08, 2.527491e-08, 2.453531e-08, 2.402773e-08, 
    2.362119e-08, 2.339063e-08, 2.281724e-08, 2.219742e-08, 2.184591e-08,
  2.421208e-08, 2.40314e-08, 2.388893e-08, 2.42088e-08, 2.48467e-08, 
    2.573741e-08, 2.592181e-08, 2.501571e-08, 2.39234e-08, 2.327709e-08, 
    2.33033e-08, 2.330661e-08, 2.272102e-08, 2.2556e-08, 2.272599e-08,
  2.359083e-08, 2.339313e-08, 2.340823e-08, 2.363163e-08, 2.46163e-08, 
    2.556158e-08, 2.580154e-08, 2.492012e-08, 2.400432e-08, 2.343909e-08, 
    2.326028e-08, 2.321793e-08, 2.264489e-08, 2.202382e-08, 2.248882e-08,
  2.309291e-08, 2.302231e-08, 2.306535e-08, 2.326452e-08, 2.47087e-08, 
    2.527204e-08, 2.595942e-08, 2.52691e-08, 2.426633e-08, 2.356691e-08, 
    2.321253e-08, 2.306809e-08, 2.258667e-08, 2.207027e-08, 2.258159e-08,
  2.325778e-08, 2.3105e-08, 2.331574e-08, 2.324471e-08, 2.391201e-08, 
    2.489387e-08, 2.538293e-08, 2.534411e-08, 2.46444e-08, 2.383625e-08, 
    2.33969e-08, 2.307105e-08, 2.252063e-08, 2.201406e-08, 2.261724e-08,
  2.304934e-08, 2.33368e-08, 2.349582e-08, 2.368867e-08, 2.387722e-08, 
    2.494318e-08, 2.511365e-08, 2.52481e-08, 2.48904e-08, 2.432502e-08, 
    2.358061e-08, 2.32216e-08, 2.259338e-08, 2.20092e-08, 2.230626e-08,
  2.262273e-08, 2.292174e-08, 2.290841e-08, 2.329845e-08, 2.385049e-08, 
    2.488961e-08, 2.519388e-08, 2.405715e-08, 2.416891e-08, 2.498846e-08, 
    2.451069e-08, 2.398833e-08, 2.281764e-08, 2.207393e-08, 2.211338e-08,
  2.248819e-08, 2.226977e-08, 2.237504e-08, 2.259865e-08, 2.362482e-08, 
    2.465256e-08, 2.548583e-08, 2.531351e-08, 2.439059e-08, 2.475581e-08, 
    2.465796e-08, 2.435095e-08, 2.338718e-08, 2.222307e-08, 2.185945e-08,
  2.22079e-08, 2.173569e-08, 2.197204e-08, 2.242208e-08, 2.392694e-08, 
    2.495502e-08, 2.575573e-08, 2.571055e-08, 2.485646e-08, 2.443575e-08, 
    2.445897e-08, 2.444006e-08, 2.407984e-08, 2.302207e-08, 2.183323e-08,
  2.136341e-08, 2.097429e-08, 2.139496e-08, 2.235139e-08, 2.433807e-08, 
    2.579065e-08, 2.603423e-08, 2.614502e-08, 2.513335e-08, 2.458517e-08, 
    2.406231e-08, 2.407753e-08, 2.393386e-08, 2.373338e-08, 2.264636e-08,
  2.204663e-08, 2.141684e-08, 2.115384e-08, 2.251474e-08, 2.458493e-08, 
    2.618077e-08, 2.667228e-08, 2.59181e-08, 2.41447e-08, 2.399006e-08, 
    2.458981e-08, 2.463268e-08, 2.397729e-08, 2.374883e-08, 2.324255e-08,
  2.331066e-08, 2.341553e-08, 2.335009e-08, 2.315904e-08, 2.3073e-08, 
    2.296281e-08, 2.35974e-08, 2.535186e-08, 2.640483e-08, 2.55341e-08, 
    2.478845e-08, 2.46813e-08, 2.473479e-08, 2.432679e-08, 2.335481e-08,
  2.30909e-08, 2.328825e-08, 2.323e-08, 2.30507e-08, 2.304044e-08, 
    2.317697e-08, 2.399059e-08, 2.563835e-08, 2.617574e-08, 2.52843e-08, 
    2.443821e-08, 2.439609e-08, 2.45954e-08, 2.397838e-08, 2.316972e-08,
  2.297234e-08, 2.311376e-08, 2.295988e-08, 2.282731e-08, 2.310561e-08, 
    2.332152e-08, 2.416736e-08, 2.566686e-08, 2.637735e-08, 2.519994e-08, 
    2.433022e-08, 2.413819e-08, 2.428452e-08, 2.405696e-08, 2.322945e-08,
  2.304188e-08, 2.304026e-08, 2.27045e-08, 2.284177e-08, 2.278445e-08, 
    2.320031e-08, 2.377443e-08, 2.565116e-08, 2.603318e-08, 2.496162e-08, 
    2.403441e-08, 2.399234e-08, 2.417942e-08, 2.383219e-08, 2.317653e-08,
  2.327736e-08, 2.308719e-08, 2.260938e-08, 2.236185e-08, 2.243693e-08, 
    2.327902e-08, 2.393742e-08, 2.497672e-08, 2.549856e-08, 2.45561e-08, 
    2.421873e-08, 2.376897e-08, 2.391059e-08, 2.369466e-08, 2.315215e-08,
  2.354074e-08, 2.315655e-08, 2.254482e-08, 2.217253e-08, 2.212574e-08, 
    2.294899e-08, 2.320558e-08, 2.175186e-08, 2.294761e-08, 2.420303e-08, 
    2.440883e-08, 2.420752e-08, 2.387285e-08, 2.352261e-08, 2.305677e-08,
  2.359127e-08, 2.320845e-08, 2.260385e-08, 2.221812e-08, 2.194517e-08, 
    2.238564e-08, 2.361788e-08, 2.370015e-08, 2.390518e-08, 2.481748e-08, 
    2.503755e-08, 2.437006e-08, 2.389449e-08, 2.340934e-08, 2.305618e-08,
  2.356033e-08, 2.348726e-08, 2.287259e-08, 2.235113e-08, 2.204336e-08, 
    2.215243e-08, 2.373592e-08, 2.483263e-08, 2.462137e-08, 2.50881e-08, 
    2.536403e-08, 2.47968e-08, 2.411332e-08, 2.336124e-08, 2.303345e-08,
  2.359178e-08, 2.374708e-08, 2.333361e-08, 2.292929e-08, 2.21898e-08, 
    2.235293e-08, 2.366405e-08, 2.526363e-08, 2.513056e-08, 2.534859e-08, 
    2.562163e-08, 2.509289e-08, 2.43818e-08, 2.36087e-08, 2.30877e-08,
  2.372175e-08, 2.391075e-08, 2.368627e-08, 2.332361e-08, 2.27757e-08, 
    2.31114e-08, 2.401548e-08, 2.559536e-08, 2.516154e-08, 2.389383e-08, 
    2.486992e-08, 2.581627e-08, 2.503079e-08, 2.394492e-08, 2.330692e-08,
  2.447644e-08, 2.46033e-08, 2.464669e-08, 2.420471e-08, 2.374763e-08, 
    2.332747e-08, 2.313825e-08, 2.317104e-08, 2.405883e-08, 2.522177e-08, 
    2.587658e-08, 2.587098e-08, 2.566665e-08, 2.549126e-08, 2.531187e-08,
  2.467191e-08, 2.490051e-08, 2.486414e-08, 2.428469e-08, 2.376297e-08, 
    2.32409e-08, 2.318613e-08, 2.328172e-08, 2.423099e-08, 2.53197e-08, 
    2.5975e-08, 2.595116e-08, 2.58509e-08, 2.542297e-08, 2.497934e-08,
  2.494518e-08, 2.50679e-08, 2.492074e-08, 2.427259e-08, 2.375429e-08, 
    2.328071e-08, 2.311768e-08, 2.325073e-08, 2.428221e-08, 2.54215e-08, 
    2.610187e-08, 2.59606e-08, 2.579118e-08, 2.556216e-08, 2.509969e-08,
  2.561138e-08, 2.553517e-08, 2.502248e-08, 2.438221e-08, 2.36774e-08, 
    2.347535e-08, 2.320214e-08, 2.325525e-08, 2.430599e-08, 2.525773e-08, 
    2.565241e-08, 2.555401e-08, 2.563378e-08, 2.559042e-08, 2.513985e-08,
  2.602237e-08, 2.535187e-08, 2.475855e-08, 2.425777e-08, 2.399346e-08, 
    2.315494e-08, 2.322281e-08, 2.303579e-08, 2.340358e-08, 2.46961e-08, 
    2.530046e-08, 2.526716e-08, 2.52723e-08, 2.534269e-08, 2.511423e-08,
  2.60779e-08, 2.524838e-08, 2.471084e-08, 2.448012e-08, 2.418477e-08, 
    2.350063e-08, 2.301079e-08, 2.290923e-08, 2.258949e-08, 2.325238e-08, 
    2.446899e-08, 2.465617e-08, 2.499007e-08, 2.515682e-08, 2.497879e-08,
  2.581636e-08, 2.493788e-08, 2.458961e-08, 2.443822e-08, 2.422995e-08, 
    2.346945e-08, 2.291524e-08, 2.314905e-08, 2.338456e-08, 2.354019e-08, 
    2.418525e-08, 2.473088e-08, 2.467259e-08, 2.493591e-08, 2.482756e-08,
  2.535992e-08, 2.480669e-08, 2.478959e-08, 2.459793e-08, 2.423636e-08, 
    2.36905e-08, 2.290791e-08, 2.328515e-08, 2.406287e-08, 2.400502e-08, 
    2.428758e-08, 2.4446e-08, 2.457526e-08, 2.47229e-08, 2.463992e-08,
  2.50417e-08, 2.49234e-08, 2.508014e-08, 2.452988e-08, 2.398076e-08, 
    2.377251e-08, 2.308735e-08, 2.381318e-08, 2.459097e-08, 2.463586e-08, 
    2.46415e-08, 2.459985e-08, 2.452495e-08, 2.450489e-08, 2.445393e-08,
  2.489626e-08, 2.495898e-08, 2.498357e-08, 2.42809e-08, 2.405456e-08, 
    2.430997e-08, 2.372406e-08, 2.433973e-08, 2.479118e-08, 2.467904e-08, 
    2.505704e-08, 2.490277e-08, 2.441647e-08, 2.438252e-08, 2.42416e-08,
  2.484111e-08, 2.444142e-08, 2.409409e-08, 2.420325e-08, 2.436985e-08, 
    2.459187e-08, 2.464357e-08, 2.489385e-08, 2.478159e-08, 2.449979e-08, 
    2.426128e-08, 2.441317e-08, 2.486883e-08, 2.522899e-08, 2.558405e-08,
  2.401879e-08, 2.398705e-08, 2.399323e-08, 2.441926e-08, 2.47859e-08, 
    2.501504e-08, 2.530636e-08, 2.538612e-08, 2.488958e-08, 2.448254e-08, 
    2.425737e-08, 2.442378e-08, 2.51106e-08, 2.528157e-08, 2.559305e-08,
  2.422436e-08, 2.470103e-08, 2.506386e-08, 2.562881e-08, 2.598214e-08, 
    2.618266e-08, 2.587791e-08, 2.543846e-08, 2.489064e-08, 2.437925e-08, 
    2.413624e-08, 2.444481e-08, 2.510281e-08, 2.549112e-08, 2.568433e-08,
  2.600857e-08, 2.657586e-08, 2.699589e-08, 2.71485e-08, 2.673975e-08, 
    2.671091e-08, 2.595253e-08, 2.546328e-08, 2.484894e-08, 2.433021e-08, 
    2.408335e-08, 2.441621e-08, 2.49873e-08, 2.556553e-08, 2.57804e-08,
  2.692843e-08, 2.724171e-08, 2.72809e-08, 2.689257e-08, 2.667293e-08, 
    2.593276e-08, 2.571307e-08, 2.546637e-08, 2.474009e-08, 2.403061e-08, 
    2.383604e-08, 2.42137e-08, 2.496853e-08, 2.585855e-08, 2.582484e-08,
  2.646532e-08, 2.65162e-08, 2.601281e-08, 2.592496e-08, 2.548151e-08, 
    2.538406e-08, 2.501323e-08, 2.471327e-08, 2.426739e-08, 2.388555e-08, 
    2.345132e-08, 2.368108e-08, 2.455243e-08, 2.580295e-08, 2.592042e-08,
  2.576516e-08, 2.544274e-08, 2.516446e-08, 2.499637e-08, 2.501727e-08, 
    2.502738e-08, 2.500944e-08, 2.4657e-08, 2.428171e-08, 2.386614e-08, 
    2.356507e-08, 2.362312e-08, 2.439858e-08, 2.567365e-08, 2.592828e-08,
  2.49751e-08, 2.49608e-08, 2.470589e-08, 2.517087e-08, 2.519627e-08, 
    2.519088e-08, 2.489428e-08, 2.445763e-08, 2.402594e-08, 2.382532e-08, 
    2.367958e-08, 2.379315e-08, 2.438359e-08, 2.543761e-08, 2.584489e-08,
  2.502589e-08, 2.499975e-08, 2.508813e-08, 2.547522e-08, 2.515736e-08, 
    2.482941e-08, 2.442888e-08, 2.403991e-08, 2.387946e-08, 2.39069e-08, 
    2.389277e-08, 2.399784e-08, 2.440339e-08, 2.53078e-08, 2.562284e-08,
  2.519561e-08, 2.516955e-08, 2.542336e-08, 2.563619e-08, 2.504811e-08, 
    2.451335e-08, 2.433586e-08, 2.438854e-08, 2.429708e-08, 2.446978e-08, 
    2.450172e-08, 2.436503e-08, 2.451768e-08, 2.516351e-08, 2.546026e-08,
  2.566125e-08, 2.568881e-08, 2.570297e-08, 2.591149e-08, 2.57638e-08, 
    2.589735e-08, 2.568632e-08, 2.547632e-08, 2.523727e-08, 2.530519e-08, 
    2.525784e-08, 2.549887e-08, 2.538543e-08, 2.523418e-08, 2.499133e-08,
  2.555057e-08, 2.537035e-08, 2.567255e-08, 2.541935e-08, 2.578211e-08, 
    2.539397e-08, 2.54992e-08, 2.534975e-08, 2.536592e-08, 2.549097e-08, 
    2.570128e-08, 2.559378e-08, 2.55977e-08, 2.534886e-08, 2.521236e-08,
  2.537438e-08, 2.538843e-08, 2.566875e-08, 2.555067e-08, 2.551437e-08, 
    2.593359e-08, 2.587944e-08, 2.648954e-08, 2.65267e-08, 2.659674e-08, 
    2.628277e-08, 2.615916e-08, 2.57813e-08, 2.556746e-08, 2.527866e-08,
  2.498003e-08, 2.518172e-08, 2.521042e-08, 2.570894e-08, 2.494419e-08, 
    2.532056e-08, 2.632537e-08, 2.680349e-08, 2.731873e-08, 2.720664e-08, 
    2.687763e-08, 2.657427e-08, 2.613168e-08, 2.553801e-08, 2.520506e-08,
  2.482295e-08, 2.501506e-08, 2.514127e-08, 2.528833e-08, 2.570211e-08, 
    2.506764e-08, 2.600872e-08, 2.626527e-08, 2.663257e-08, 2.659765e-08, 
    2.672212e-08, 2.64651e-08, 2.596266e-08, 2.517882e-08, 2.493123e-08,
  2.482339e-08, 2.500297e-08, 2.503295e-08, 2.519042e-08, 2.526364e-08, 
    2.520457e-08, 2.545159e-08, 2.54267e-08, 2.535601e-08, 2.59209e-08, 
    2.602755e-08, 2.594932e-08, 2.531362e-08, 2.470223e-08, 2.473262e-08,
  2.464072e-08, 2.471863e-08, 2.496022e-08, 2.5173e-08, 2.503005e-08, 
    2.50947e-08, 2.49079e-08, 2.499936e-08, 2.504715e-08, 2.522026e-08, 
    2.529961e-08, 2.523828e-08, 2.47215e-08, 2.427015e-08, 2.463951e-08,
  2.42171e-08, 2.46548e-08, 2.511791e-08, 2.516159e-08, 2.518876e-08, 
    2.523784e-08, 2.528946e-08, 2.526291e-08, 2.511076e-08, 2.516205e-08, 
    2.511911e-08, 2.492357e-08, 2.44993e-08, 2.416326e-08, 2.471893e-08,
  2.425238e-08, 2.46217e-08, 2.483477e-08, 2.509721e-08, 2.528597e-08, 
    2.545322e-08, 2.559622e-08, 2.543478e-08, 2.525399e-08, 2.502098e-08, 
    2.471661e-08, 2.459364e-08, 2.431314e-08, 2.414956e-08, 2.487286e-08,
  2.406282e-08, 2.439094e-08, 2.473017e-08, 2.487943e-08, 2.514452e-08, 
    2.519089e-08, 2.507655e-08, 2.494818e-08, 2.489861e-08, 2.475494e-08, 
    2.445547e-08, 2.424457e-08, 2.413127e-08, 2.413174e-08, 2.510375e-08,
  2.49149e-08, 2.487014e-08, 2.48094e-08, 2.485048e-08, 2.479824e-08, 
    2.50059e-08, 2.520157e-08, 2.524173e-08, 2.540038e-08, 2.551092e-08, 
    2.542437e-08, 2.567054e-08, 2.576021e-08, 2.57709e-08, 2.572189e-08,
  2.516604e-08, 2.498472e-08, 2.477647e-08, 2.464277e-08, 2.459435e-08, 
    2.477304e-08, 2.48663e-08, 2.520613e-08, 2.521536e-08, 2.52963e-08, 
    2.539151e-08, 2.55656e-08, 2.579935e-08, 2.546027e-08, 2.550998e-08,
  2.524507e-08, 2.488687e-08, 2.447898e-08, 2.419894e-08, 2.444065e-08, 
    2.421474e-08, 2.445565e-08, 2.488271e-08, 2.517082e-08, 2.543692e-08, 
    2.583656e-08, 2.607944e-08, 2.615333e-08, 2.559908e-08, 2.577378e-08,
  2.524967e-08, 2.481183e-08, 2.433754e-08, 2.423744e-08, 2.394518e-08, 
    2.41418e-08, 2.399382e-08, 2.397194e-08, 2.449697e-08, 2.504366e-08, 
    2.561703e-08, 2.614994e-08, 2.608015e-08, 2.633839e-08, 2.649094e-08,
  2.541925e-08, 2.483521e-08, 2.435546e-08, 2.389892e-08, 2.40775e-08, 
    2.376129e-08, 2.424652e-08, 2.429927e-08, 2.444553e-08, 2.452915e-08, 
    2.499467e-08, 2.536883e-08, 2.570785e-08, 2.642879e-08, 2.681528e-08,
  2.54825e-08, 2.48258e-08, 2.403743e-08, 2.402507e-08, 2.388725e-08, 
    2.431984e-08, 2.444151e-08, 2.473762e-08, 2.414994e-08, 2.44886e-08, 
    2.500691e-08, 2.543744e-08, 2.581965e-08, 2.656355e-08, 2.668027e-08,
  2.532985e-08, 2.471581e-08, 2.424571e-08, 2.414265e-08, 2.419551e-08, 
    2.447236e-08, 2.451773e-08, 2.488872e-08, 2.511264e-08, 2.487591e-08, 
    2.490268e-08, 2.531032e-08, 2.572945e-08, 2.621072e-08, 2.645228e-08,
  2.525315e-08, 2.498061e-08, 2.435782e-08, 2.423295e-08, 2.429899e-08, 
    2.442016e-08, 2.455631e-08, 2.496143e-08, 2.514739e-08, 2.516938e-08, 
    2.510872e-08, 2.521021e-08, 2.551415e-08, 2.59113e-08, 2.622534e-08,
  2.534429e-08, 2.480431e-08, 2.449933e-08, 2.448808e-08, 2.442064e-08, 
    2.439749e-08, 2.459334e-08, 2.496614e-08, 2.523148e-08, 2.538257e-08, 
    2.526256e-08, 2.52398e-08, 2.52671e-08, 2.560271e-08, 2.590662e-08,
  2.512152e-08, 2.461511e-08, 2.482682e-08, 2.471366e-08, 2.448508e-08, 
    2.454624e-08, 2.46547e-08, 2.48638e-08, 2.521561e-08, 2.547388e-08, 
    2.536068e-08, 2.524428e-08, 2.518056e-08, 2.55144e-08, 2.563938e-08,
  2.603754e-08, 2.655864e-08, 2.69263e-08, 2.701779e-08, 2.677993e-08, 
    2.654699e-08, 2.604354e-08, 2.559851e-08, 2.517815e-08, 2.489166e-08, 
    2.459401e-08, 2.44162e-08, 2.431445e-08, 2.422329e-08, 2.447401e-08,
  2.655816e-08, 2.709233e-08, 2.751781e-08, 2.730306e-08, 2.720161e-08, 
    2.651708e-08, 2.6145e-08, 2.54155e-08, 2.493642e-08, 2.465266e-08, 
    2.45316e-08, 2.438464e-08, 2.451231e-08, 2.443898e-08, 2.419217e-08,
  2.699266e-08, 2.73549e-08, 2.740092e-08, 2.703868e-08, 2.734769e-08, 
    2.633831e-08, 2.552681e-08, 2.490995e-08, 2.448104e-08, 2.414187e-08, 
    2.411965e-08, 2.409246e-08, 2.42733e-08, 2.445197e-08, 2.452741e-08,
  2.683759e-08, 2.68961e-08, 2.680349e-08, 2.682484e-08, 2.629659e-08, 
    2.662217e-08, 2.53136e-08, 2.472636e-08, 2.415401e-08, 2.405707e-08, 
    2.390454e-08, 2.392485e-08, 2.410527e-08, 2.42574e-08, 2.47901e-08,
  2.636254e-08, 2.637119e-08, 2.640971e-08, 2.605969e-08, 2.595553e-08, 
    2.54832e-08, 2.563817e-08, 2.507966e-08, 2.421581e-08, 2.396572e-08, 
    2.36535e-08, 2.377664e-08, 2.37918e-08, 2.405899e-08, 2.423501e-08,
  2.584541e-08, 2.595204e-08, 2.570461e-08, 2.574725e-08, 2.529821e-08, 
    2.525225e-08, 2.506246e-08, 2.489559e-08, 2.469938e-08, 2.424989e-08, 
    2.378551e-08, 2.393418e-08, 2.39528e-08, 2.415418e-08, 2.429765e-08,
  2.549727e-08, 2.55921e-08, 2.555062e-08, 2.546843e-08, 2.514281e-08, 
    2.513625e-08, 2.509034e-08, 2.492309e-08, 2.466929e-08, 2.441702e-08, 
    2.41483e-08, 2.417103e-08, 2.422868e-08, 2.436416e-08, 2.455884e-08,
  2.533254e-08, 2.535245e-08, 2.525781e-08, 2.512922e-08, 2.527248e-08, 
    2.52092e-08, 2.504891e-08, 2.499107e-08, 2.468304e-08, 2.454853e-08, 
    2.44649e-08, 2.44497e-08, 2.444624e-08, 2.463568e-08, 2.456108e-08,
  2.544052e-08, 2.528385e-08, 2.500724e-08, 2.513461e-08, 2.549755e-08, 
    2.536902e-08, 2.516344e-08, 2.497483e-08, 2.473963e-08, 2.465809e-08, 
    2.466651e-08, 2.481804e-08, 2.478029e-08, 2.48649e-08, 2.47604e-08,
  2.574715e-08, 2.541869e-08, 2.519734e-08, 2.546315e-08, 2.57638e-08, 
    2.56789e-08, 2.524279e-08, 2.493583e-08, 2.479098e-08, 2.471513e-08, 
    2.484551e-08, 2.508229e-08, 2.514228e-08, 2.50215e-08, 2.499023e-08,
  2.573555e-08, 2.56019e-08, 2.578016e-08, 2.592592e-08, 2.612505e-08, 
    2.673632e-08, 2.74378e-08, 2.741702e-08, 2.744986e-08, 2.746045e-08, 
    2.743452e-08, 2.728833e-08, 2.678942e-08, 2.620953e-08, 2.552228e-08,
  2.592496e-08, 2.573319e-08, 2.587316e-08, 2.574663e-08, 2.617813e-08, 
    2.683346e-08, 2.747113e-08, 2.715015e-08, 2.666967e-08, 2.674961e-08, 
    2.701297e-08, 2.664571e-08, 2.663069e-08, 2.595311e-08, 2.532681e-08,
  2.59418e-08, 2.575618e-08, 2.560013e-08, 2.547573e-08, 2.60292e-08, 
    2.688346e-08, 2.592856e-08, 2.570414e-08, 2.575793e-08, 2.582185e-08, 
    2.608866e-08, 2.59981e-08, 2.577902e-08, 2.541267e-08, 2.514594e-08,
  2.61626e-08, 2.595532e-08, 2.579484e-08, 2.557743e-08, 2.602287e-08, 
    2.528784e-08, 2.44321e-08, 2.461559e-08, 2.468569e-08, 2.531109e-08, 
    2.560009e-08, 2.552562e-08, 2.514925e-08, 2.490545e-08, 2.485601e-08,
  2.639717e-08, 2.613012e-08, 2.568954e-08, 2.552516e-08, 2.541534e-08, 
    2.4407e-08, 2.524575e-08, 2.472297e-08, 2.542759e-08, 2.595359e-08, 
    2.594648e-08, 2.557756e-08, 2.503685e-08, 2.441119e-08, 2.444024e-08,
  2.644595e-08, 2.60937e-08, 2.554939e-08, 2.544364e-08, 2.577601e-08, 
    2.540207e-08, 2.475335e-08, 2.485667e-08, 2.531925e-08, 2.562843e-08, 
    2.522207e-08, 2.482627e-08, 2.436874e-08, 2.408056e-08, 2.383932e-08,
  2.642368e-08, 2.597598e-08, 2.564303e-08, 2.547453e-08, 2.582403e-08, 
    2.497585e-08, 2.502528e-08, 2.457326e-08, 2.486597e-08, 2.504117e-08, 
    2.51342e-08, 2.489736e-08, 2.430145e-08, 2.39769e-08, 2.375335e-08,
  2.627359e-08, 2.554521e-08, 2.530557e-08, 2.528648e-08, 2.589747e-08, 
    2.519831e-08, 2.479935e-08, 2.431691e-08, 2.46459e-08, 2.510145e-08, 
    2.538569e-08, 2.507791e-08, 2.450416e-08, 2.416431e-08, 2.348804e-08,
  2.623567e-08, 2.548464e-08, 2.54212e-08, 2.573566e-08, 2.589102e-08, 
    2.492962e-08, 2.469477e-08, 2.433453e-08, 2.441547e-08, 2.483768e-08, 
    2.50785e-08, 2.476058e-08, 2.448091e-08, 2.436162e-08, 2.37564e-08,
  2.578082e-08, 2.523616e-08, 2.475738e-08, 2.516216e-08, 2.591699e-08, 
    2.478623e-08, 2.432338e-08, 2.41186e-08, 2.430338e-08, 2.476306e-08, 
    2.489899e-08, 2.478735e-08, 2.458337e-08, 2.437355e-08, 2.399195e-08,
  2.659741e-08, 2.542111e-08, 2.519432e-08, 2.529142e-08, 2.544631e-08, 
    2.515534e-08, 2.515736e-08, 2.525877e-08, 2.452282e-08, 2.388037e-08, 
    2.430514e-08, 2.511579e-08, 2.602888e-08, 2.711183e-08, 2.771826e-08,
  2.535919e-08, 2.476449e-08, 2.459713e-08, 2.505815e-08, 2.533276e-08, 
    2.460193e-08, 2.476373e-08, 2.498122e-08, 2.42888e-08, 2.381116e-08, 
    2.445355e-08, 2.53476e-08, 2.635291e-08, 2.700444e-08, 2.737257e-08,
  2.430653e-08, 2.412532e-08, 2.460088e-08, 2.523257e-08, 2.505798e-08, 
    2.451082e-08, 2.442666e-08, 2.496445e-08, 2.477138e-08, 2.38922e-08, 
    2.448439e-08, 2.565957e-08, 2.623863e-08, 2.635438e-08, 2.707863e-08,
  2.407867e-08, 2.451761e-08, 2.484352e-08, 2.506982e-08, 2.544607e-08, 
    2.523072e-08, 2.502334e-08, 2.468937e-08, 2.472644e-08, 2.421131e-08, 
    2.456927e-08, 2.564483e-08, 2.590782e-08, 2.594369e-08, 2.62635e-08,
  2.442511e-08, 2.444909e-08, 2.441629e-08, 2.519138e-08, 2.535801e-08, 
    2.510456e-08, 2.583472e-08, 2.498843e-08, 2.523728e-08, 2.414249e-08, 
    2.425621e-08, 2.534462e-08, 2.547469e-08, 2.548524e-08, 2.593693e-08,
  2.352321e-08, 2.344929e-08, 2.401042e-08, 2.460416e-08, 2.544836e-08, 
    2.550851e-08, 2.509607e-08, 2.655523e-08, 2.64107e-08, 2.513235e-08, 
    2.455119e-08, 2.51171e-08, 2.484686e-08, 2.486877e-08, 2.525838e-08,
  2.279259e-08, 2.254729e-08, 2.313984e-08, 2.431464e-08, 2.483871e-08, 
    2.565307e-08, 2.56055e-08, 2.499067e-08, 2.500667e-08, 2.558493e-08, 
    2.534517e-08, 2.528907e-08, 2.473446e-08, 2.453314e-08, 2.467703e-08,
  2.259658e-08, 2.236036e-08, 2.258918e-08, 2.334312e-08, 2.432083e-08, 
    2.515297e-08, 2.529287e-08, 2.533797e-08, 2.563347e-08, 2.537391e-08, 
    2.53583e-08, 2.51293e-08, 2.474958e-08, 2.445405e-08, 2.413758e-08,
  2.329375e-08, 2.281442e-08, 2.297545e-08, 2.335534e-08, 2.371512e-08, 
    2.505022e-08, 2.558488e-08, 2.51508e-08, 2.507472e-08, 2.569509e-08, 
    2.561155e-08, 2.531992e-08, 2.471909e-08, 2.450022e-08, 2.361427e-08,
  2.404438e-08, 2.349026e-08, 2.322132e-08, 2.328889e-08, 2.361599e-08, 
    2.423793e-08, 2.532434e-08, 2.547633e-08, 2.515142e-08, 2.506373e-08, 
    2.54321e-08, 2.570323e-08, 2.500407e-08, 2.449554e-08, 2.359115e-08,
  2.413112e-08, 2.410194e-08, 2.447237e-08, 2.519955e-08, 2.52332e-08, 
    2.454582e-08, 2.53565e-08, 2.604388e-08, 2.520078e-08, 2.459211e-08, 
    2.479857e-08, 2.584046e-08, 2.671358e-08, 2.694819e-08, 2.74201e-08,
  2.376436e-08, 2.401793e-08, 2.426426e-08, 2.504143e-08, 2.520167e-08, 
    2.456169e-08, 2.49248e-08, 2.607264e-08, 2.551295e-08, 2.48001e-08, 
    2.454194e-08, 2.537553e-08, 2.62604e-08, 2.6874e-08, 2.731935e-08,
  2.338836e-08, 2.400704e-08, 2.449603e-08, 2.480864e-08, 2.488909e-08, 
    2.469279e-08, 2.480756e-08, 2.601888e-08, 2.583612e-08, 2.496172e-08, 
    2.480072e-08, 2.498556e-08, 2.579084e-08, 2.706455e-08, 2.741119e-08,
  2.361281e-08, 2.437342e-08, 2.48533e-08, 2.494363e-08, 2.530264e-08, 
    2.52761e-08, 2.484554e-08, 2.498274e-08, 2.544388e-08, 2.550177e-08, 
    2.475417e-08, 2.458484e-08, 2.48154e-08, 2.5385e-08, 2.631429e-08,
  2.375669e-08, 2.466178e-08, 2.5162e-08, 2.504173e-08, 2.517756e-08, 
    2.569704e-08, 2.598126e-08, 2.492043e-08, 2.488185e-08, 2.543894e-08, 
    2.564598e-08, 2.471281e-08, 2.472876e-08, 2.504737e-08, 2.523749e-08,
  2.445008e-08, 2.513744e-08, 2.523995e-08, 2.514147e-08, 2.550398e-08, 
    2.538161e-08, 2.530092e-08, 2.583564e-08, 2.559433e-08, 2.482025e-08, 
    2.565232e-08, 2.526368e-08, 2.442202e-08, 2.42621e-08, 2.472377e-08,
  2.517824e-08, 2.569751e-08, 2.553613e-08, 2.553066e-08, 2.588207e-08, 
    2.598009e-08, 2.556223e-08, 2.504135e-08, 2.56753e-08, 2.549165e-08, 
    2.511111e-08, 2.553261e-08, 2.49363e-08, 2.408857e-08, 2.367975e-08,
  2.557066e-08, 2.577604e-08, 2.542776e-08, 2.563933e-08, 2.625384e-08, 
    2.645952e-08, 2.642284e-08, 2.588669e-08, 2.627246e-08, 2.562132e-08, 
    2.486602e-08, 2.539272e-08, 2.537768e-08, 2.466928e-08, 2.333169e-08,
  2.589671e-08, 2.568582e-08, 2.550265e-08, 2.610036e-08, 2.682377e-08, 
    2.721362e-08, 2.68707e-08, 2.616865e-08, 2.653608e-08, 2.628937e-08, 
    2.493456e-08, 2.541399e-08, 2.513562e-08, 2.54791e-08, 2.396312e-08,
  2.577386e-08, 2.538079e-08, 2.528079e-08, 2.607705e-08, 2.730865e-08, 
    2.789261e-08, 2.740906e-08, 2.64373e-08, 2.687013e-08, 2.403713e-08, 
    2.434009e-08, 2.591735e-08, 2.508068e-08, 2.536897e-08, 2.510082e-08,
  2.409237e-08, 2.382034e-08, 2.494633e-08, 2.567118e-08, 2.609828e-08, 
    2.636208e-08, 2.682093e-08, 2.775404e-08, 2.729872e-08, 2.566944e-08, 
    2.450196e-08, 2.484314e-08, 2.568559e-08, 2.624271e-08, 2.645912e-08,
  2.393533e-08, 2.475454e-08, 2.575308e-08, 2.58211e-08, 2.62827e-08, 
    2.627262e-08, 2.689129e-08, 2.720631e-08, 2.733069e-08, 2.635152e-08, 
    2.48862e-08, 2.452859e-08, 2.487348e-08, 2.582128e-08, 2.591179e-08,
  2.429022e-08, 2.547486e-08, 2.599842e-08, 2.58349e-08, 2.620742e-08, 
    2.657734e-08, 2.67926e-08, 2.724503e-08, 2.755864e-08, 2.686147e-08, 
    2.528358e-08, 2.468038e-08, 2.424539e-08, 2.569019e-08, 2.580541e-08,
  2.515118e-08, 2.591567e-08, 2.599468e-08, 2.571136e-08, 2.605761e-08, 
    2.637762e-08, 2.670555e-08, 2.675101e-08, 2.733205e-08, 2.70201e-08, 
    2.563623e-08, 2.524849e-08, 2.418531e-08, 2.388498e-08, 2.504904e-08,
  2.596115e-08, 2.596494e-08, 2.56907e-08, 2.546557e-08, 2.589504e-08, 
    2.583303e-08, 2.649814e-08, 2.685375e-08, 2.731979e-08, 2.672726e-08, 
    2.527112e-08, 2.579871e-08, 2.479276e-08, 2.404357e-08, 2.430354e-08,
  2.628303e-08, 2.575582e-08, 2.526239e-08, 2.526618e-08, 2.532861e-08, 
    2.55025e-08, 2.593422e-08, 2.646337e-08, 2.716665e-08, 2.635895e-08, 
    2.463022e-08, 2.484325e-08, 2.515473e-08, 2.4357e-08, 2.394759e-08,
  2.640038e-08, 2.563674e-08, 2.511695e-08, 2.4868e-08, 2.498705e-08, 
    2.513585e-08, 2.57422e-08, 2.60722e-08, 2.627766e-08, 2.629851e-08, 
    2.464028e-08, 2.44034e-08, 2.439035e-08, 2.48591e-08, 2.421714e-08,
  2.592462e-08, 2.548587e-08, 2.487326e-08, 2.469375e-08, 2.453566e-08, 
    2.432525e-08, 2.526498e-08, 2.584943e-08, 2.608644e-08, 2.630139e-08, 
    2.458487e-08, 2.392498e-08, 2.353322e-08, 2.38764e-08, 2.495418e-08,
  2.548974e-08, 2.502474e-08, 2.484746e-08, 2.452114e-08, 2.433144e-08, 
    2.425938e-08, 2.500372e-08, 2.536024e-08, 2.574523e-08, 2.560483e-08, 
    2.419813e-08, 2.433392e-08, 2.338751e-08, 2.354354e-08, 2.384171e-08,
  2.491288e-08, 2.440755e-08, 2.43853e-08, 2.406733e-08, 2.401302e-08, 
    2.400347e-08, 2.46324e-08, 2.464155e-08, 2.486768e-08, 2.393922e-08, 
    2.383122e-08, 2.410131e-08, 2.425837e-08, 2.364529e-08, 2.344703e-08,
  2.428044e-08, 2.477629e-08, 2.493801e-08, 2.454619e-08, 2.460965e-08, 
    2.449725e-08, 2.46273e-08, 2.460324e-08, 2.483596e-08, 2.504717e-08, 
    2.499336e-08, 2.479263e-08, 2.444624e-08, 2.446186e-08, 2.504149e-08,
  2.463961e-08, 2.493332e-08, 2.495724e-08, 2.452357e-08, 2.446261e-08, 
    2.429625e-08, 2.45779e-08, 2.45847e-08, 2.48027e-08, 2.484664e-08, 
    2.482029e-08, 2.474738e-08, 2.468844e-08, 2.422571e-08, 2.450531e-08,
  2.471243e-08, 2.504455e-08, 2.524805e-08, 2.491505e-08, 2.46662e-08, 
    2.439977e-08, 2.496274e-08, 2.496651e-08, 2.479637e-08, 2.46562e-08, 
    2.457746e-08, 2.446555e-08, 2.459065e-08, 2.473879e-08, 2.448555e-08,
  2.525111e-08, 2.534762e-08, 2.549766e-08, 2.5764e-08, 2.623633e-08, 
    2.573416e-08, 2.4957e-08, 2.501655e-08, 2.475875e-08, 2.487471e-08, 
    2.444928e-08, 2.442096e-08, 2.443806e-08, 2.438344e-08, 2.452069e-08,
  2.576727e-08, 2.670714e-08, 2.726799e-08, 2.656356e-08, 2.547644e-08, 
    2.570942e-08, 2.586754e-08, 2.48781e-08, 2.4763e-08, 2.495732e-08, 
    2.461095e-08, 2.433738e-08, 2.435382e-08, 2.444014e-08, 2.458856e-08,
  2.711347e-08, 2.816093e-08, 2.605885e-08, 2.544577e-08, 2.569362e-08, 
    2.463799e-08, 2.429174e-08, 2.514619e-08, 2.508206e-08, 2.461723e-08, 
    2.470376e-08, 2.450397e-08, 2.44618e-08, 2.433185e-08, 2.444707e-08,
  2.746825e-08, 2.667635e-08, 2.458737e-08, 2.312941e-08, 2.297028e-08, 
    2.370127e-08, 2.324638e-08, 2.288584e-08, 2.313062e-08, 2.405142e-08, 
    2.435857e-08, 2.431971e-08, 2.456481e-08, 2.469653e-08, 2.45796e-08,
  2.769576e-08, 2.55223e-08, 2.459002e-08, 2.355137e-08, 2.225486e-08, 
    2.322163e-08, 2.301424e-08, 2.318514e-08, 2.298623e-08, 2.334228e-08, 
    2.383617e-08, 2.39748e-08, 2.42907e-08, 2.482951e-08, 2.482597e-08,
  2.819078e-08, 2.724935e-08, 2.579389e-08, 2.454722e-08, 2.278409e-08, 
    2.465781e-08, 2.394725e-08, 2.314527e-08, 2.265426e-08, 2.2941e-08, 
    2.325367e-08, 2.355075e-08, 2.410892e-08, 2.475504e-08, 2.503938e-08,
  2.758508e-08, 2.821961e-08, 2.871799e-08, 2.975406e-08, 2.683754e-08, 
    2.696555e-08, 2.526554e-08, 2.309226e-08, 2.206983e-08, 2.222076e-08, 
    2.278526e-08, 2.337015e-08, 2.397065e-08, 2.482636e-08, 2.545033e-08,
  2.43932e-08, 2.45351e-08, 2.538864e-08, 2.555716e-08, 2.55296e-08, 
    2.607704e-08, 2.603092e-08, 2.454989e-08, 2.351867e-08, 2.258857e-08, 
    2.244471e-08, 2.257756e-08, 2.297277e-08, 2.253431e-08, 2.241056e-08,
  2.471256e-08, 2.529802e-08, 2.584798e-08, 2.605882e-08, 2.647295e-08, 
    2.694526e-08, 2.602514e-08, 2.448515e-08, 2.351803e-08, 2.34376e-08, 
    2.484312e-08, 2.572466e-08, 2.465625e-08, 2.196212e-08, 2.223233e-08,
  2.510979e-08, 2.592142e-08, 2.593641e-08, 2.689556e-08, 2.711543e-08, 
    2.953027e-08, 2.733342e-08, 2.484662e-08, 2.364143e-08, 2.645207e-08, 
    2.860559e-08, 2.727233e-08, 2.41643e-08, 2.220718e-08, 2.401036e-08,
  2.579714e-08, 2.661509e-08, 2.69911e-08, 2.830836e-08, 2.693514e-08, 
    2.544678e-08, 2.634944e-08, 2.533675e-08, 2.568478e-08, 3.103335e-08, 
    2.892522e-08, 2.475303e-08, 2.241045e-08, 2.297025e-08, 2.58956e-08,
  2.679618e-08, 2.723648e-08, 2.713075e-08, 2.795961e-08, 2.760953e-08, 
    2.519962e-08, 2.392194e-08, 2.446058e-08, 2.831055e-08, 3.208076e-08, 
    2.626826e-08, 2.256832e-08, 2.2299e-08, 2.419639e-08, 2.558139e-08,
  2.796198e-08, 2.713269e-08, 2.634626e-08, 2.691537e-08, 2.671661e-08, 
    2.539705e-08, 2.594719e-08, 2.794414e-08, 2.987521e-08, 2.576131e-08, 
    2.250974e-08, 2.197769e-08, 2.310161e-08, 2.379289e-08, 2.379603e-08,
  2.877714e-08, 2.86937e-08, 2.497993e-08, 2.528766e-08, 2.595858e-08, 
    2.86376e-08, 3.075289e-08, 2.958565e-08, 2.838579e-08, 2.561822e-08, 
    2.508064e-08, 2.390068e-08, 2.299315e-08, 2.252429e-08, 2.337023e-08,
  2.980186e-08, 2.956861e-08, 2.893916e-08, 2.925738e-08, 3.084726e-08, 
    3.263033e-08, 3.088147e-08, 3.029264e-08, 2.946253e-08, 2.834103e-08, 
    2.56772e-08, 2.280225e-08, 2.187083e-08, 2.255443e-08, 2.325352e-08,
  3.133045e-08, 3.06249e-08, 3.108065e-08, 3.108305e-08, 3.191757e-08, 
    3.134891e-08, 3.021781e-08, 2.929493e-08, 2.768169e-08, 2.574189e-08, 
    2.30863e-08, 2.182854e-08, 2.24558e-08, 2.316986e-08, 2.395693e-08,
  2.938164e-08, 2.931969e-08, 2.948216e-08, 2.987452e-08, 2.92247e-08, 
    3.003608e-08, 2.90275e-08, 2.792187e-08, 2.538538e-08, 2.399208e-08, 
    2.253226e-08, 2.27689e-08, 2.427034e-08, 2.428858e-08, 2.480125e-08,
  2.347579e-08, 2.361826e-08, 2.410589e-08, 2.413477e-08, 2.419467e-08, 
    2.483776e-08, 2.533187e-08, 2.553347e-08, 2.5806e-08, 2.593387e-08, 
    2.793382e-08, 3.038123e-08, 2.929326e-08, 2.774138e-08, 2.618938e-08,
  2.359153e-08, 2.3753e-08, 2.392113e-08, 2.374311e-08, 2.351172e-08, 
    2.445048e-08, 2.641211e-08, 2.717688e-08, 2.771442e-08, 2.828495e-08, 
    2.930892e-08, 2.978084e-08, 2.784021e-08, 2.593323e-08, 2.457107e-08,
  2.26137e-08, 2.297375e-08, 2.296897e-08, 2.341126e-08, 2.234188e-08, 
    2.550514e-08, 3.026904e-08, 3.121483e-08, 2.996421e-08, 2.898199e-08, 
    2.854929e-08, 2.730864e-08, 2.572523e-08, 2.445045e-08, 2.387341e-08,
  2.233543e-08, 2.268878e-08, 2.273799e-08, 2.380582e-08, 2.127627e-08, 
    2.077312e-08, 2.573266e-08, 2.892581e-08, 2.794605e-08, 2.630157e-08, 
    2.547895e-08, 2.416935e-08, 2.336116e-08, 2.352992e-08, 2.371479e-08,
  2.360223e-08, 2.392458e-08, 2.390592e-08, 2.44317e-08, 2.469874e-08, 
    2.194175e-08, 1.952427e-08, 2.068692e-08, 2.196691e-08, 2.280528e-08, 
    2.322368e-08, 2.319485e-08, 2.389802e-08, 2.468125e-08, 2.504031e-08,
  2.431069e-08, 2.449199e-08, 2.486749e-08, 2.480756e-08, 2.494728e-08, 
    2.47492e-08, 2.333059e-08, 2.236645e-08, 2.30588e-08, 2.446479e-08, 
    2.486102e-08, 2.516167e-08, 2.561504e-08, 2.526586e-08, 2.492128e-08,
  2.472517e-08, 2.455042e-08, 2.460528e-08, 2.413578e-08, 2.441433e-08, 
    2.367985e-08, 2.425481e-08, 2.515596e-08, 2.583099e-08, 2.587414e-08, 
    2.594929e-08, 2.611649e-08, 2.588259e-08, 2.506179e-08, 2.423064e-08,
  2.305539e-08, 2.27974e-08, 2.282126e-08, 2.328706e-08, 2.373162e-08, 
    2.491262e-08, 2.658945e-08, 2.767961e-08, 2.770912e-08, 2.685503e-08, 
    2.651854e-08, 2.612133e-08, 2.509709e-08, 2.409549e-08, 2.372182e-08,
  2.182696e-08, 2.272661e-08, 2.384144e-08, 2.526474e-08, 2.692536e-08, 
    2.875262e-08, 2.990939e-08, 2.943117e-08, 2.787303e-08, 2.634494e-08, 
    2.512522e-08, 2.412181e-08, 2.357977e-08, 2.349471e-08, 2.413978e-08,
  2.419391e-08, 2.63166e-08, 2.817238e-08, 3.034319e-08, 3.096683e-08, 
    3.102786e-08, 2.981575e-08, 2.780049e-08, 2.527807e-08, 2.369369e-08, 
    2.306176e-08, 2.312031e-08, 2.341798e-08, 2.406014e-08, 2.44593e-08,
  2.318407e-08, 2.360037e-08, 2.391531e-08, 2.340833e-08, 2.304805e-08, 
    2.301738e-08, 2.303162e-08, 2.296205e-08, 2.315534e-08, 2.330582e-08, 
    2.374087e-08, 2.375177e-08, 2.360772e-08, 2.303487e-08, 2.29551e-08,
  2.360335e-08, 2.382771e-08, 2.359272e-08, 2.323003e-08, 2.318981e-08, 
    2.308067e-08, 2.317065e-08, 2.338281e-08, 2.36965e-08, 2.3596e-08, 
    2.336406e-08, 2.256357e-08, 2.242971e-08, 2.22633e-08, 2.267246e-08,
  2.341607e-08, 2.340403e-08, 2.331037e-08, 2.326639e-08, 2.344341e-08, 
    2.344113e-08, 2.368868e-08, 2.418156e-08, 2.413071e-08, 2.360167e-08, 
    2.289738e-08, 2.253288e-08, 2.276025e-08, 2.356146e-08, 2.472705e-08,
  2.331066e-08, 2.341891e-08, 2.331065e-08, 2.370886e-08, 2.378049e-08, 
    2.403446e-08, 2.445305e-08, 2.441444e-08, 2.373426e-08, 2.329119e-08, 
    2.325919e-08, 2.373005e-08, 2.481604e-08, 2.600155e-08, 2.697633e-08,
  2.308455e-08, 2.296188e-08, 2.337049e-08, 2.368761e-08, 2.454547e-08, 
    2.384192e-08, 2.448935e-08, 2.386239e-08, 2.340226e-08, 2.372196e-08, 
    2.452941e-08, 2.558431e-08, 2.642826e-08, 2.722647e-08, 2.704105e-08,
  2.283707e-08, 2.316797e-08, 2.354814e-08, 2.418854e-08, 2.409452e-08, 
    2.421132e-08, 2.381544e-08, 2.392162e-08, 2.479337e-08, 2.544458e-08, 
    2.609655e-08, 2.656482e-08, 2.677091e-08, 2.639584e-08, 2.596562e-08,
  2.30912e-08, 2.35599e-08, 2.403814e-08, 2.390497e-08, 2.385436e-08, 
    2.371185e-08, 2.386519e-08, 2.429291e-08, 2.492232e-08, 2.582855e-08, 
    2.619799e-08, 2.623625e-08, 2.54081e-08, 2.492879e-08, 2.4613e-08,
  2.376104e-08, 2.429931e-08, 2.427308e-08, 2.417269e-08, 2.410736e-08, 
    2.447744e-08, 2.504931e-08, 2.585181e-08, 2.662639e-08, 2.669084e-08, 
    2.601169e-08, 2.462345e-08, 2.404969e-08, 2.405792e-08, 2.475725e-08,
  2.438278e-08, 2.460989e-08, 2.460477e-08, 2.471728e-08, 2.525604e-08, 
    2.566884e-08, 2.616994e-08, 2.626742e-08, 2.580111e-08, 2.469281e-08, 
    2.353072e-08, 2.344689e-08, 2.385791e-08, 2.465582e-08, 2.506483e-08,
  2.428191e-08, 2.446987e-08, 2.456575e-08, 2.504581e-08, 2.514983e-08, 
    2.524017e-08, 2.479232e-08, 2.393847e-08, 2.348878e-08, 2.31578e-08, 
    2.356377e-08, 2.430298e-08, 2.474575e-08, 2.54266e-08, 2.522366e-08,
  2.194762e-08, 2.215272e-08, 2.220191e-08, 2.172122e-08, 2.254754e-08, 
    2.279579e-08, 2.283375e-08, 2.311752e-08, 2.361532e-08, 2.370641e-08, 
    2.364471e-08, 2.367217e-08, 2.367724e-08, 2.378125e-08, 2.345112e-08,
  2.229252e-08, 2.22624e-08, 2.202143e-08, 2.196083e-08, 2.286257e-08, 
    2.265818e-08, 2.287897e-08, 2.327068e-08, 2.343414e-08, 2.348524e-08, 
    2.374819e-08, 2.385582e-08, 2.406592e-08, 2.385923e-08, 2.395952e-08,
  2.222155e-08, 2.207505e-08, 2.206535e-08, 2.22382e-08, 2.263208e-08, 
    2.227945e-08, 2.265126e-08, 2.30071e-08, 2.320303e-08, 2.340291e-08, 
    2.365317e-08, 2.396841e-08, 2.401687e-08, 2.408313e-08, 2.462453e-08,
  2.23304e-08, 2.233046e-08, 2.255591e-08, 2.249859e-08, 2.235648e-08, 
    2.305402e-08, 2.270022e-08, 2.27178e-08, 2.265173e-08, 2.304958e-08, 
    2.364984e-08, 2.400077e-08, 2.409053e-08, 2.425287e-08, 2.448318e-08,
  2.243154e-08, 2.262297e-08, 2.278462e-08, 2.262221e-08, 2.274556e-08, 
    2.225529e-08, 2.283343e-08, 2.246257e-08, 2.24877e-08, 2.33093e-08, 
    2.397721e-08, 2.402762e-08, 2.412942e-08, 2.433795e-08, 2.442665e-08,
  2.28009e-08, 2.301267e-08, 2.314589e-08, 2.28901e-08, 2.24908e-08, 
    2.263511e-08, 2.27002e-08, 2.343987e-08, 2.43095e-08, 2.406013e-08, 
    2.416501e-08, 2.419728e-08, 2.442991e-08, 2.465368e-08, 2.493955e-08,
  2.325857e-08, 2.334102e-08, 2.331702e-08, 2.282079e-08, 2.306969e-08, 
    2.298015e-08, 2.322717e-08, 2.325841e-08, 2.325615e-08, 2.355493e-08, 
    2.430943e-08, 2.447787e-08, 2.468827e-08, 2.496608e-08, 2.51395e-08,
  2.380263e-08, 2.384635e-08, 2.379303e-08, 2.34701e-08, 2.337412e-08, 
    2.333289e-08, 2.340266e-08, 2.336834e-08, 2.364715e-08, 2.439342e-08, 
    2.47317e-08, 2.474124e-08, 2.496894e-08, 2.509868e-08, 2.545915e-08,
  2.455809e-08, 2.471882e-08, 2.410141e-08, 2.356599e-08, 2.365888e-08, 
    2.354626e-08, 2.345095e-08, 2.354581e-08, 2.383499e-08, 2.456652e-08, 
    2.481775e-08, 2.493713e-08, 2.493831e-08, 2.534878e-08, 2.535281e-08,
  2.540202e-08, 2.497374e-08, 2.403944e-08, 2.38918e-08, 2.434988e-08, 
    2.375975e-08, 2.363437e-08, 2.365569e-08, 2.417038e-08, 2.496262e-08, 
    2.50812e-08, 2.501455e-08, 2.520374e-08, 2.523587e-08, 2.550274e-08,
  2.337078e-08, 2.327679e-08, 2.408994e-08, 2.518972e-08, 2.530228e-08, 
    2.50103e-08, 2.504206e-08, 2.592268e-08, 2.540682e-08, 2.447724e-08, 
    2.416965e-08, 2.408449e-08, 2.420451e-08, 2.52144e-08, 2.601491e-08,
  2.353386e-08, 2.354538e-08, 2.465368e-08, 2.520764e-08, 2.5057e-08, 
    2.51728e-08, 2.532619e-08, 2.568742e-08, 2.531291e-08, 2.476753e-08, 
    2.418123e-08, 2.424248e-08, 2.468786e-08, 2.562939e-08, 2.631324e-08,
  2.394343e-08, 2.396218e-08, 2.514986e-08, 2.534365e-08, 2.479119e-08, 
    2.482371e-08, 2.552489e-08, 2.624919e-08, 2.564811e-08, 2.51876e-08, 
    2.504912e-08, 2.479375e-08, 2.499227e-08, 2.59905e-08, 2.691771e-08,
  2.415542e-08, 2.440876e-08, 2.545782e-08, 2.479792e-08, 2.45361e-08, 
    2.500444e-08, 2.600896e-08, 2.571961e-08, 2.522012e-08, 2.540851e-08, 
    2.505553e-08, 2.475377e-08, 2.532802e-08, 2.611938e-08, 2.685765e-08,
  2.447179e-08, 2.474108e-08, 2.52817e-08, 2.460635e-08, 2.488972e-08, 
    2.527985e-08, 2.60417e-08, 2.58311e-08, 2.549798e-08, 2.531223e-08, 
    2.514224e-08, 2.482079e-08, 2.490789e-08, 2.59783e-08, 2.693712e-08,
  2.433567e-08, 2.456005e-08, 2.495255e-08, 2.465479e-08, 2.506764e-08, 
    2.602721e-08, 2.617215e-08, 2.566737e-08, 2.525676e-08, 2.45327e-08, 
    2.468103e-08, 2.466571e-08, 2.501685e-08, 2.597721e-08, 2.673456e-08,
  2.397162e-08, 2.441377e-08, 2.472329e-08, 2.476793e-08, 2.551937e-08, 
    2.586306e-08, 2.602433e-08, 2.536084e-08, 2.443583e-08, 2.403628e-08, 
    2.456093e-08, 2.439447e-08, 2.478168e-08, 2.626297e-08, 2.684885e-08,
  2.340788e-08, 2.421874e-08, 2.460457e-08, 2.487307e-08, 2.544231e-08, 
    2.591129e-08, 2.561333e-08, 2.46108e-08, 2.407765e-08, 2.371622e-08, 
    2.406358e-08, 2.447467e-08, 2.535494e-08, 2.647938e-08, 2.651274e-08,
  2.380516e-08, 2.441671e-08, 2.44301e-08, 2.474673e-08, 2.547009e-08, 
    2.582009e-08, 2.535548e-08, 2.445559e-08, 2.388781e-08, 2.299751e-08, 
    2.404872e-08, 2.487107e-08, 2.572427e-08, 2.653569e-08, 2.663498e-08,
  2.410009e-08, 2.409553e-08, 2.419651e-08, 2.483824e-08, 2.570184e-08, 
    2.591072e-08, 2.509547e-08, 2.401585e-08, 2.324665e-08, 2.31045e-08, 
    2.432322e-08, 2.542319e-08, 2.650829e-08, 2.67366e-08, 2.655336e-08,
  2.19824e-08, 2.191661e-08, 2.207667e-08, 2.228143e-08, 2.286979e-08, 
    2.315635e-08, 2.319169e-08, 2.363369e-08, 2.406634e-08, 2.378882e-08, 
    2.422308e-08, 2.402303e-08, 2.486268e-08, 2.495155e-08, 2.403024e-08,
  2.199128e-08, 2.190525e-08, 2.226443e-08, 2.236664e-08, 2.270519e-08, 
    2.27096e-08, 2.297263e-08, 2.290676e-08, 2.290163e-08, 2.280928e-08, 
    2.362612e-08, 2.40189e-08, 2.493266e-08, 2.410485e-08, 2.325952e-08,
  2.195896e-08, 2.206848e-08, 2.232441e-08, 2.240987e-08, 2.251042e-08, 
    2.212957e-08, 2.242157e-08, 2.220602e-08, 2.198603e-08, 2.247731e-08, 
    2.345233e-08, 2.409977e-08, 2.474262e-08, 2.41373e-08, 2.344012e-08,
  2.223168e-08, 2.222674e-08, 2.229139e-08, 2.249394e-08, 2.227612e-08, 
    2.214932e-08, 2.19781e-08, 2.199351e-08, 2.230196e-08, 2.277316e-08, 
    2.353706e-08, 2.425737e-08, 2.451418e-08, 2.386923e-08, 2.361798e-08,
  2.249615e-08, 2.22835e-08, 2.231372e-08, 2.233197e-08, 2.24867e-08, 
    2.224658e-08, 2.249639e-08, 2.261311e-08, 2.291375e-08, 2.321839e-08, 
    2.391629e-08, 2.414668e-08, 2.391017e-08, 2.370937e-08, 2.399855e-08,
  2.241195e-08, 2.236251e-08, 2.233458e-08, 2.263565e-08, 2.271075e-08, 
    2.299151e-08, 2.309389e-08, 2.332668e-08, 2.327441e-08, 2.370718e-08, 
    2.391913e-08, 2.376018e-08, 2.36549e-08, 2.401814e-08, 2.415138e-08,
  2.261159e-08, 2.280193e-08, 2.293137e-08, 2.317225e-08, 2.338067e-08, 
    2.352379e-08, 2.369105e-08, 2.373397e-08, 2.352645e-08, 2.378427e-08, 
    2.396854e-08, 2.376981e-08, 2.404061e-08, 2.466721e-08, 2.406896e-08,
  2.300638e-08, 2.329421e-08, 2.340896e-08, 2.370816e-08, 2.390584e-08, 
    2.409388e-08, 2.419882e-08, 2.4113e-08, 2.413265e-08, 2.451471e-08, 
    2.457098e-08, 2.433401e-08, 2.48563e-08, 2.484527e-08, 2.347141e-08,
  2.37991e-08, 2.396804e-08, 2.399129e-08, 2.428629e-08, 2.444208e-08, 
    2.462992e-08, 2.471419e-08, 2.450845e-08, 2.475874e-08, 2.52576e-08, 
    2.500463e-08, 2.451411e-08, 2.496572e-08, 2.40797e-08, 2.276896e-08,
  2.435141e-08, 2.445165e-08, 2.450999e-08, 2.472631e-08, 2.478411e-08, 
    2.50864e-08, 2.503222e-08, 2.537751e-08, 2.5989e-08, 2.61916e-08, 
    2.521816e-08, 2.477624e-08, 2.439429e-08, 2.306156e-08, 2.230614e-08,
  2.361685e-08, 2.394272e-08, 2.375743e-08, 2.446385e-08, 2.316906e-08, 
    2.31601e-08, 2.32723e-08, 2.374375e-08, 2.396627e-08, 2.402972e-08, 
    2.360978e-08, 2.327426e-08, 2.286912e-08, 2.299702e-08, 2.33015e-08,
  2.434843e-08, 2.410741e-08, 2.383163e-08, 2.385334e-08, 2.30161e-08, 
    2.495473e-08, 2.557034e-08, 2.580707e-08, 2.577639e-08, 2.477919e-08, 
    2.451648e-08, 2.377092e-08, 2.333353e-08, 2.335737e-08, 2.366301e-08,
  2.337292e-08, 2.347558e-08, 2.291929e-08, 2.31937e-08, 2.297625e-08, 
    2.340208e-08, 2.835081e-08, 2.718887e-08, 2.647622e-08, 2.57385e-08, 
    2.481542e-08, 2.406511e-08, 2.359467e-08, 2.366498e-08, 2.400314e-08,
  2.317205e-08, 2.34029e-08, 2.412798e-08, 2.4406e-08, 2.4988e-08, 
    2.250493e-08, 2.324889e-08, 2.577749e-08, 2.534438e-08, 2.483755e-08, 
    2.436846e-08, 2.392401e-08, 2.390192e-08, 2.400395e-08, 2.416994e-08,
  2.658988e-08, 2.698622e-08, 2.694831e-08, 2.684616e-08, 2.708563e-08, 
    2.609668e-08, 2.151223e-08, 2.250259e-08, 2.357522e-08, 2.374679e-08, 
    2.383742e-08, 2.392956e-08, 2.415575e-08, 2.439211e-08, 2.47033e-08,
  2.673283e-08, 2.662211e-08, 2.617484e-08, 2.591147e-08, 2.55901e-08, 
    2.510183e-08, 2.496098e-08, 2.338441e-08, 2.345509e-08, 2.364784e-08, 
    2.386964e-08, 2.415846e-08, 2.443305e-08, 2.480978e-08, 2.5145e-08,
  2.442795e-08, 2.348786e-08, 2.293022e-08, 2.25112e-08, 2.241603e-08, 
    2.254599e-08, 2.262318e-08, 2.30045e-08, 2.350192e-08, 2.374762e-08, 
    2.421988e-08, 2.454656e-08, 2.508949e-08, 2.535077e-08, 2.525586e-08,
  2.197018e-08, 2.166516e-08, 2.16771e-08, 2.164277e-08, 2.181235e-08, 
    2.200938e-08, 2.24234e-08, 2.324546e-08, 2.38765e-08, 2.437637e-08, 
    2.489967e-08, 2.538571e-08, 2.566654e-08, 2.55652e-08, 2.58241e-08,
  2.365412e-08, 2.400637e-08, 2.438452e-08, 2.45755e-08, 2.445931e-08, 
    2.441165e-08, 2.450955e-08, 2.510066e-08, 2.547544e-08, 2.615934e-08, 
    2.594463e-08, 2.602314e-08, 2.575682e-08, 2.59424e-08, 2.580465e-08,
  2.654916e-08, 2.650706e-08, 2.655272e-08, 2.614305e-08, 2.599137e-08, 
    2.563028e-08, 2.543705e-08, 2.558596e-08, 2.555735e-08, 2.498448e-08, 
    2.512945e-08, 2.525326e-08, 2.568925e-08, 2.614365e-08, 2.591945e-08,
  2.439185e-08, 2.393192e-08, 2.35912e-08, 2.356917e-08, 2.330321e-08, 
    2.309768e-08, 2.295647e-08, 2.284546e-08, 2.343688e-08, 2.41956e-08, 
    2.593362e-08, 2.761421e-08, 2.798847e-08, 2.782921e-08, 2.821204e-08,
  2.528243e-08, 2.504565e-08, 2.48889e-08, 2.505063e-08, 2.461538e-08, 
    2.436486e-08, 2.429907e-08, 2.505196e-08, 2.608058e-08, 2.800967e-08, 
    2.951419e-08, 2.938517e-08, 2.865487e-08, 2.729186e-08, 2.63885e-08,
  2.48306e-08, 2.490686e-08, 2.481455e-08, 2.528887e-08, 2.437415e-08, 
    2.481078e-08, 2.964786e-08, 3.64555e-08, 3.727539e-08, 3.722055e-08, 
    3.541794e-08, 3.279382e-08, 3.062839e-08, 2.889043e-08, 2.603234e-08,
  2.466268e-08, 2.422486e-08, 2.400521e-08, 2.422829e-08, 2.328966e-08, 
    2.004897e-08, 2.0932e-08, 3.179421e-08, 3.282067e-08, 3.227677e-08, 
    3.068264e-08, 2.890248e-08, 2.745889e-08, 2.523835e-08, 2.316237e-08,
  2.542728e-08, 2.554749e-08, 2.48745e-08, 2.498346e-08, 2.477315e-08, 
    2.32129e-08, 1.595555e-08, 1.161963e-08, 1.545135e-08, 1.642726e-08, 
    1.759206e-08, 1.859768e-08, 1.938459e-08, 2.037507e-08, 2.075867e-08,
  2.574071e-08, 2.578843e-08, 2.540907e-08, 2.527785e-08, 2.511463e-08, 
    2.516221e-08, 2.462977e-08, 1.878358e-08, 1.648183e-08, 1.678895e-08, 
    1.648171e-08, 1.699069e-08, 1.797818e-08, 1.983948e-08, 2.130306e-08,
  2.641317e-08, 2.626342e-08, 2.604872e-08, 2.595411e-08, 2.566652e-08, 
    2.550705e-08, 2.523229e-08, 2.481889e-08, 2.361154e-08, 2.264446e-08, 
    2.141642e-08, 2.099558e-08, 2.162951e-08, 2.269643e-08, 2.330574e-08,
  2.635287e-08, 2.63728e-08, 2.62917e-08, 2.633169e-08, 2.598815e-08, 
    2.583553e-08, 2.527299e-08, 2.496153e-08, 2.470438e-08, 2.418515e-08, 
    2.372412e-08, 2.402736e-08, 2.451154e-08, 2.456583e-08, 2.388991e-08,
  2.475956e-08, 2.524592e-08, 2.553122e-08, 2.570961e-08, 2.584284e-08, 
    2.553316e-08, 2.487547e-08, 2.417155e-08, 2.378901e-08, 2.451083e-08, 
    2.44223e-08, 2.450537e-08, 2.446016e-08, 2.39984e-08, 2.368381e-08,
  2.336985e-08, 2.364787e-08, 2.404996e-08, 2.50056e-08, 2.5767e-08, 
    2.586014e-08, 2.60268e-08, 2.614188e-08, 2.592906e-08, 2.518747e-08, 
    2.438715e-08, 2.475918e-08, 2.477254e-08, 2.469253e-08, 2.459653e-08,
  2.597115e-08, 2.57151e-08, 2.558775e-08, 2.544792e-08, 2.533413e-08, 
    2.513667e-08, 2.487211e-08, 2.459798e-08, 2.433792e-08, 2.400889e-08, 
    2.377209e-08, 2.336795e-08, 2.298633e-08, 2.272317e-08, 2.237861e-08,
  2.601432e-08, 2.572791e-08, 2.554093e-08, 2.54951e-08, 2.537304e-08, 
    2.562338e-08, 2.557709e-08, 2.487425e-08, 2.441754e-08, 2.393205e-08, 
    2.367754e-08, 2.316615e-08, 2.308693e-08, 2.281846e-08, 2.260519e-08,
  2.618748e-08, 2.582348e-08, 2.554219e-08, 2.559828e-08, 2.495885e-08, 
    2.553307e-08, 2.728776e-08, 2.945082e-08, 2.798409e-08, 2.631091e-08, 
    2.520427e-08, 2.424136e-08, 2.397508e-08, 2.398989e-08, 2.480653e-08,
  2.587898e-08, 2.592736e-08, 2.557276e-08, 2.553993e-08, 2.493896e-08, 
    2.262649e-08, 2.430311e-08, 2.837509e-08, 2.879549e-08, 2.84224e-08, 
    2.825785e-08, 2.808356e-08, 2.868542e-08, 2.878482e-08, 2.96639e-08,
  2.589923e-08, 2.631003e-08, 2.613772e-08, 2.581801e-08, 2.555559e-08, 
    2.462605e-08, 2.143065e-08, 1.88809e-08, 2.251952e-08, 2.479229e-08, 
    2.646293e-08, 2.739819e-08, 2.801942e-08, 2.885107e-08, 2.940477e-08,
  2.541418e-08, 2.575934e-08, 2.604986e-08, 2.619095e-08, 2.605179e-08, 
    2.582743e-08, 2.507477e-08, 2.365062e-08, 2.19847e-08, 2.24873e-08, 
    2.256541e-08, 2.273153e-08, 2.261024e-08, 2.260765e-08, 2.224625e-08,
  2.398638e-08, 2.471384e-08, 2.505308e-08, 2.577639e-08, 2.621041e-08, 
    2.610602e-08, 2.597823e-08, 2.563871e-08, 2.534993e-08, 2.446409e-08, 
    2.394942e-08, 2.302156e-08, 2.258421e-08, 2.202705e-08, 2.132679e-08,
  2.326333e-08, 2.371064e-08, 2.403671e-08, 2.499745e-08, 2.551556e-08, 
    2.605138e-08, 2.639497e-08, 2.586246e-08, 2.620976e-08, 2.593659e-08, 
    2.579629e-08, 2.537031e-08, 2.451856e-08, 2.380187e-08, 2.313844e-08,
  2.292332e-08, 2.34953e-08, 2.338104e-08, 2.368793e-08, 2.457578e-08, 
    2.561935e-08, 2.572823e-08, 2.689711e-08, 2.78177e-08, 2.799203e-08, 
    2.804559e-08, 2.80311e-08, 2.79588e-08, 2.770255e-08, 2.73162e-08,
  2.358452e-08, 2.363553e-08, 2.361468e-08, 2.315129e-08, 2.344875e-08, 
    2.511246e-08, 2.568522e-08, 2.820093e-08, 2.740846e-08, 2.546195e-08, 
    2.412011e-08, 2.283136e-08, 2.315961e-08, 2.368875e-08, 2.439629e-08,
  2.631943e-08, 2.664627e-08, 2.696028e-08, 2.708822e-08, 2.713782e-08, 
    2.702882e-08, 2.689051e-08, 2.662999e-08, 2.660435e-08, 2.658868e-08, 
    2.668939e-08, 2.671507e-08, 2.673197e-08, 2.66564e-08, 2.66016e-08,
  2.552543e-08, 2.580895e-08, 2.614243e-08, 2.644891e-08, 2.665886e-08, 
    2.704469e-08, 2.721362e-08, 2.690951e-08, 2.649654e-08, 2.620603e-08, 
    2.618662e-08, 2.591327e-08, 2.622058e-08, 2.615723e-08, 2.636934e-08,
  2.480848e-08, 2.516436e-08, 2.545149e-08, 2.575279e-08, 2.584109e-08, 
    2.613495e-08, 2.655087e-08, 3.022327e-08, 3.011994e-08, 2.950719e-08, 
    2.870869e-08, 2.744898e-08, 2.654741e-08, 2.565744e-08, 2.551436e-08,
  2.459708e-08, 2.473067e-08, 2.493851e-08, 2.522277e-08, 2.563644e-08, 
    2.449313e-08, 2.424599e-08, 2.65358e-08, 2.889733e-08, 3.077649e-08, 
    3.137858e-08, 3.149841e-08, 3.109532e-08, 3.003801e-08, 2.906042e-08,
  2.408012e-08, 2.382096e-08, 2.382153e-08, 2.43257e-08, 2.506004e-08, 
    2.497398e-08, 2.446888e-08, 1.915632e-08, 1.827683e-08, 1.790552e-08, 
    1.976698e-08, 2.303409e-08, 2.609903e-08, 2.793615e-08, 2.889172e-08,
  2.400976e-08, 2.334009e-08, 2.278224e-08, 2.305434e-08, 2.342593e-08, 
    2.435319e-08, 2.520741e-08, 2.449028e-08, 2.30622e-08, 2.190653e-08, 
    2.074777e-08, 2.065779e-08, 2.105905e-08, 2.227049e-08, 2.400944e-08,
  2.440267e-08, 2.342984e-08, 2.243305e-08, 2.219776e-08, 2.236831e-08, 
    2.330688e-08, 2.443408e-08, 2.5352e-08, 2.579457e-08, 2.612339e-08, 
    2.539105e-08, 2.494772e-08, 2.383248e-08, 2.354327e-08, 2.318897e-08,
  2.488521e-08, 2.377364e-08, 2.251148e-08, 2.188057e-08, 2.1748e-08, 
    2.288019e-08, 2.370558e-08, 2.479112e-08, 2.585905e-08, 2.663041e-08, 
    2.73862e-08, 2.656564e-08, 2.653666e-08, 2.540135e-08, 2.438073e-08,
  2.558249e-08, 2.462822e-08, 2.316609e-08, 2.182437e-08, 2.152563e-08, 
    2.261918e-08, 2.392501e-08, 2.525033e-08, 2.704071e-08, 2.715352e-08, 
    2.797464e-08, 2.847336e-08, 2.859451e-08, 2.828016e-08, 2.65959e-08,
  2.583415e-08, 2.536521e-08, 2.398039e-08, 2.235743e-08, 2.185159e-08, 
    2.284402e-08, 2.429635e-08, 2.559672e-08, 2.596806e-08, 2.417632e-08, 
    2.322519e-08, 2.343294e-08, 2.507096e-08, 2.703052e-08, 2.651029e-08,
  2.489548e-08, 2.46542e-08, 2.488392e-08, 2.500107e-08, 2.575553e-08, 
    2.615451e-08, 2.704793e-08, 2.749926e-08, 2.773187e-08, 2.790481e-08, 
    2.742409e-08, 2.721499e-08, 2.665942e-08, 2.64073e-08, 2.639985e-08,
  2.505194e-08, 2.476446e-08, 2.45892e-08, 2.443805e-08, 2.463185e-08, 
    2.500125e-08, 2.57162e-08, 2.62832e-08, 2.677725e-08, 2.714593e-08, 
    2.75342e-08, 2.721618e-08, 2.750319e-08, 2.699804e-08, 2.689364e-08,
  2.498441e-08, 2.469503e-08, 2.450442e-08, 2.405307e-08, 2.423099e-08, 
    2.4474e-08, 2.580593e-08, 2.756942e-08, 2.778981e-08, 2.754722e-08, 
    2.7771e-08, 2.760986e-08, 2.765792e-08, 2.716028e-08, 2.701813e-08,
  2.506826e-08, 2.482877e-08, 2.441674e-08, 2.391278e-08, 2.318162e-08, 
    2.185102e-08, 2.230256e-08, 2.518274e-08, 2.655527e-08, 2.766638e-08, 
    2.80558e-08, 2.853887e-08, 2.897966e-08, 2.903282e-08, 2.918216e-08,
  2.487619e-08, 2.486437e-08, 2.486264e-08, 2.446879e-08, 2.356283e-08, 
    2.236072e-08, 2.038063e-08, 1.920426e-08, 2.093987e-08, 2.233667e-08, 
    2.421534e-08, 2.506147e-08, 2.601692e-08, 2.733142e-08, 2.837279e-08,
  2.564927e-08, 2.580772e-08, 2.612102e-08, 2.545226e-08, 2.432778e-08, 
    2.34849e-08, 2.247142e-08, 2.128806e-08, 2.086155e-08, 2.142413e-08, 
    2.223731e-08, 2.325655e-08, 2.325951e-08, 2.356096e-08, 2.413894e-08,
  2.593394e-08, 2.671036e-08, 2.705577e-08, 2.595382e-08, 2.47993e-08, 
    2.410155e-08, 2.359785e-08, 2.32778e-08, 2.277562e-08, 2.286958e-08, 
    2.285892e-08, 2.340529e-08, 2.346439e-08, 2.344047e-08, 2.340099e-08,
  2.609521e-08, 2.743181e-08, 2.722481e-08, 2.562612e-08, 2.458938e-08, 
    2.41567e-08, 2.42084e-08, 2.43957e-08, 2.424994e-08, 2.400168e-08, 
    2.358616e-08, 2.355849e-08, 2.363202e-08, 2.395084e-08, 2.292821e-08,
  2.607144e-08, 2.76386e-08, 2.740127e-08, 2.567948e-08, 2.438913e-08, 
    2.412842e-08, 2.481305e-08, 2.505913e-08, 2.633922e-08, 2.677261e-08, 
    2.636565e-08, 2.600226e-08, 2.537697e-08, 2.531636e-08, 2.493131e-08,
  2.609857e-08, 2.756368e-08, 2.750803e-08, 2.568463e-08, 2.406244e-08, 
    2.434004e-08, 2.554219e-08, 2.61716e-08, 2.74136e-08, 2.657988e-08, 
    2.608203e-08, 2.587132e-08, 2.624886e-08, 2.681432e-08, 2.674488e-08,
  2.55412e-08, 2.592279e-08, 2.60726e-08, 2.625742e-08, 2.614891e-08, 
    2.565743e-08, 2.51816e-08, 2.479829e-08, 2.473977e-08, 2.494424e-08, 
    2.544629e-08, 2.616848e-08, 2.640062e-08, 2.677201e-08, 2.673039e-08,
  2.548451e-08, 2.565576e-08, 2.587339e-08, 2.58412e-08, 2.588976e-08, 
    2.585175e-08, 2.552787e-08, 2.524673e-08, 2.48763e-08, 2.482781e-08, 
    2.488663e-08, 2.53416e-08, 2.621407e-08, 2.651537e-08, 2.681317e-08,
  2.595615e-08, 2.599766e-08, 2.634466e-08, 2.591864e-08, 2.59431e-08, 
    2.551362e-08, 2.576084e-08, 2.559643e-08, 2.538467e-08, 2.51564e-08, 
    2.503712e-08, 2.480854e-08, 2.535204e-08, 2.582254e-08, 2.648958e-08,
  2.61609e-08, 2.644547e-08, 2.640442e-08, 2.660194e-08, 2.605944e-08, 
    2.596065e-08, 2.523292e-08, 2.532123e-08, 2.545858e-08, 2.54208e-08, 
    2.582191e-08, 2.55084e-08, 2.542878e-08, 2.55748e-08, 2.590059e-08,
  2.652043e-08, 2.667631e-08, 2.689165e-08, 2.705675e-08, 2.727009e-08, 
    2.68106e-08, 2.62043e-08, 2.527623e-08, 2.449456e-08, 2.43489e-08, 
    2.5118e-08, 2.554727e-08, 2.560202e-08, 2.575687e-08, 2.574679e-08,
  2.675317e-08, 2.693749e-08, 2.725874e-08, 2.750254e-08, 2.795191e-08, 
    2.776356e-08, 2.749951e-08, 2.653123e-08, 2.520744e-08, 2.365214e-08, 
    2.324815e-08, 2.418474e-08, 2.516923e-08, 2.57826e-08, 2.620542e-08,
  2.661598e-08, 2.67287e-08, 2.680049e-08, 2.711007e-08, 2.699508e-08, 
    2.710281e-08, 2.683752e-08, 2.698447e-08, 2.647751e-08, 2.505477e-08, 
    2.311299e-08, 2.251929e-08, 2.337467e-08, 2.468947e-08, 2.556692e-08,
  2.636195e-08, 2.652678e-08, 2.65858e-08, 2.595426e-08, 2.550657e-08, 
    2.527251e-08, 2.530907e-08, 2.54827e-08, 2.559978e-08, 2.558074e-08, 
    2.457254e-08, 2.271421e-08, 2.223489e-08, 2.329419e-08, 2.428832e-08,
  2.613091e-08, 2.615627e-08, 2.593822e-08, 2.50651e-08, 2.449059e-08, 
    2.433041e-08, 2.440018e-08, 2.486807e-08, 2.479733e-08, 2.484613e-08, 
    2.452396e-08, 2.309559e-08, 2.188285e-08, 2.201912e-08, 2.279012e-08,
  2.595812e-08, 2.592321e-08, 2.58313e-08, 2.498368e-08, 2.442842e-08, 
    2.490851e-08, 2.59773e-08, 2.572255e-08, 2.555045e-08, 2.53622e-08, 
    2.527036e-08, 2.468637e-08, 2.287507e-08, 2.193825e-08, 2.227639e-08,
  2.407709e-08, 2.366265e-08, 2.378409e-08, 2.387676e-08, 2.463957e-08, 
    2.57284e-08, 2.651231e-08, 2.589314e-08, 2.420788e-08, 2.349591e-08, 
    2.408812e-08, 2.493722e-08, 2.541522e-08, 2.532966e-08, 2.519489e-08,
  2.318605e-08, 2.265071e-08, 2.272956e-08, 2.298295e-08, 2.299029e-08, 
    2.415708e-08, 2.54549e-08, 2.608827e-08, 2.590915e-08, 2.457715e-08, 
    2.425648e-08, 2.458614e-08, 2.542676e-08, 2.565657e-08, 2.53053e-08,
  2.281142e-08, 2.187059e-08, 2.148846e-08, 2.13671e-08, 2.283787e-08, 
    2.338132e-08, 2.448241e-08, 2.568306e-08, 2.612499e-08, 2.571864e-08, 
    2.492151e-08, 2.447196e-08, 2.477239e-08, 2.534119e-08, 2.568171e-08,
  2.171e-08, 2.139549e-08, 2.107832e-08, 2.149153e-08, 2.251159e-08, 
    2.400688e-08, 2.469589e-08, 2.555302e-08, 2.639321e-08, 2.654735e-08, 
    2.632661e-08, 2.563464e-08, 2.513372e-08, 2.50523e-08, 2.551664e-08,
  2.217229e-08, 2.263498e-08, 2.286343e-08, 2.347915e-08, 2.420716e-08, 
    2.509898e-08, 2.563199e-08, 2.614353e-08, 2.629241e-08, 2.633366e-08, 
    2.668613e-08, 2.642307e-08, 2.600519e-08, 2.555291e-08, 2.540283e-08,
  2.570477e-08, 2.56347e-08, 2.554253e-08, 2.567362e-08, 2.591496e-08, 
    2.610727e-08, 2.676027e-08, 2.634345e-08, 2.605281e-08, 2.652941e-08, 
    2.702648e-08, 2.711452e-08, 2.684847e-08, 2.64051e-08, 2.587058e-08,
  2.621814e-08, 2.604792e-08, 2.611191e-08, 2.601882e-08, 2.595703e-08, 
    2.605067e-08, 2.658569e-08, 2.702353e-08, 2.727759e-08, 2.709712e-08, 
    2.689623e-08, 2.686568e-08, 2.67594e-08, 2.654155e-08, 2.605248e-08,
  2.607532e-08, 2.607612e-08, 2.612484e-08, 2.584808e-08, 2.55188e-08, 
    2.527295e-08, 2.559952e-08, 2.621627e-08, 2.701255e-08, 2.754079e-08, 
    2.767363e-08, 2.716456e-08, 2.673012e-08, 2.67065e-08, 2.640988e-08,
  2.58915e-08, 2.599949e-08, 2.594611e-08, 2.55601e-08, 2.499804e-08, 
    2.486424e-08, 2.447957e-08, 2.493341e-08, 2.560061e-08, 2.671617e-08, 
    2.745529e-08, 2.730901e-08, 2.653656e-08, 2.611408e-08, 2.60733e-08,
  2.557013e-08, 2.55482e-08, 2.57089e-08, 2.569971e-08, 2.55672e-08, 
    2.528339e-08, 2.58947e-08, 2.525294e-08, 2.518608e-08, 2.592532e-08, 
    2.714622e-08, 2.730703e-08, 2.654651e-08, 2.604869e-08, 2.558667e-08,
  2.710386e-08, 2.678685e-08, 2.674612e-08, 2.714813e-08, 2.814203e-08, 
    2.89595e-08, 2.80934e-08, 2.762303e-08, 2.678191e-08, 2.569212e-08, 
    2.462848e-08, 2.480395e-08, 2.469641e-08, 2.476895e-08, 2.478821e-08,
  2.688652e-08, 2.682299e-08, 2.685341e-08, 2.717571e-08, 2.790383e-08, 
    2.760569e-08, 2.784e-08, 2.744972e-08, 2.761218e-08, 2.730247e-08, 
    2.61249e-08, 2.52935e-08, 2.556306e-08, 2.538863e-08, 2.494003e-08,
  2.62843e-08, 2.715872e-08, 2.780022e-08, 2.715678e-08, 2.68827e-08, 
    2.523322e-08, 2.511382e-08, 2.680743e-08, 2.771082e-08, 2.792114e-08, 
    2.729632e-08, 2.60378e-08, 2.56876e-08, 2.563765e-08, 2.556898e-08,
  2.576751e-08, 2.772295e-08, 2.868054e-08, 2.787606e-08, 2.638039e-08, 
    2.511869e-08, 2.405121e-08, 2.452266e-08, 2.779943e-08, 2.897621e-08, 
    2.858396e-08, 2.680398e-08, 2.573004e-08, 2.532431e-08, 2.538454e-08,
  2.41571e-08, 2.479831e-08, 2.64074e-08, 2.631983e-08, 2.514014e-08, 
    2.3944e-08, 2.33525e-08, 2.2484e-08, 2.332984e-08, 2.475039e-08, 
    2.740429e-08, 2.699724e-08, 2.56448e-08, 2.479469e-08, 2.490991e-08,
  2.604052e-08, 2.501714e-08, 2.428729e-08, 2.426241e-08, 2.387518e-08, 
    2.303235e-08, 2.281437e-08, 2.033098e-08, 1.997262e-08, 2.21463e-08, 
    2.579195e-08, 2.721593e-08, 2.624952e-08, 2.444729e-08, 2.398415e-08,
  2.605731e-08, 2.612114e-08, 2.568319e-08, 2.47916e-08, 2.432853e-08, 
    2.350496e-08, 2.328494e-08, 2.211888e-08, 2.036682e-08, 2.025123e-08, 
    2.197393e-08, 2.563174e-08, 2.661531e-08, 2.47412e-08, 2.344899e-08,
  2.559174e-08, 2.585534e-08, 2.612211e-08, 2.605773e-08, 2.562926e-08, 
    2.480227e-08, 2.420524e-08, 2.37377e-08, 2.298244e-08, 2.158336e-08, 
    2.15482e-08, 2.332392e-08, 2.606252e-08, 2.587618e-08, 2.416717e-08,
  2.505729e-08, 2.528029e-08, 2.554452e-08, 2.573736e-08, 2.569782e-08, 
    2.566241e-08, 2.532094e-08, 2.508948e-08, 2.502814e-08, 2.495392e-08, 
    2.408998e-08, 2.375051e-08, 2.527149e-08, 2.619387e-08, 2.542724e-08,
  2.465284e-08, 2.477985e-08, 2.49329e-08, 2.519828e-08, 2.536322e-08, 
    2.534447e-08, 2.543302e-08, 2.531089e-08, 2.525043e-08, 2.561018e-08, 
    2.575686e-08, 2.533078e-08, 2.57598e-08, 2.648667e-08, 2.639189e-08,
  2.63408e-08, 2.631594e-08, 2.641899e-08, 2.552579e-08, 2.586201e-08, 
    2.658994e-08, 2.611276e-08, 2.605205e-08, 2.589579e-08, 2.630353e-08, 
    2.664669e-08, 2.662904e-08, 2.634209e-08, 2.587337e-08, 2.555077e-08,
  2.599317e-08, 2.63528e-08, 2.657416e-08, 2.696357e-08, 2.57969e-08, 
    2.681473e-08, 2.688232e-08, 2.625286e-08, 2.575538e-08, 2.617051e-08, 
    2.65325e-08, 2.666106e-08, 2.663941e-08, 2.585564e-08, 2.541138e-08,
  2.55978e-08, 2.566828e-08, 2.630174e-08, 2.630248e-08, 2.709068e-08, 
    2.629456e-08, 2.713434e-08, 2.776945e-08, 2.637423e-08, 2.579785e-08, 
    2.606924e-08, 2.610961e-08, 2.618598e-08, 2.567003e-08, 2.529918e-08,
  2.550538e-08, 2.523465e-08, 2.586664e-08, 2.576188e-08, 2.662471e-08, 
    2.680949e-08, 2.624824e-08, 2.733181e-08, 2.860467e-08, 2.741156e-08, 
    2.666075e-08, 2.632767e-08, 2.622134e-08, 2.604998e-08, 2.570745e-08,
  2.567339e-08, 2.54585e-08, 2.55731e-08, 2.60902e-08, 2.642347e-08, 
    2.706355e-08, 2.633946e-08, 2.518708e-08, 2.594401e-08, 2.755264e-08, 
    2.754205e-08, 2.680453e-08, 2.690329e-08, 2.701745e-08, 2.68215e-08,
  2.529788e-08, 2.587046e-08, 2.549034e-08, 2.588967e-08, 2.691506e-08, 
    2.708204e-08, 2.752587e-08, 2.620021e-08, 2.488902e-08, 2.698804e-08, 
    2.912008e-08, 2.842263e-08, 2.77983e-08, 2.79275e-08, 2.761543e-08,
  2.484958e-08, 2.547496e-08, 2.598067e-08, 2.539051e-08, 2.612656e-08, 
    2.727416e-08, 2.76868e-08, 2.770564e-08, 2.665092e-08, 2.637477e-08, 
    2.743205e-08, 2.89682e-08, 2.867289e-08, 2.865439e-08, 2.784123e-08,
  2.445486e-08, 2.509668e-08, 2.553682e-08, 2.588499e-08, 2.576873e-08, 
    2.601274e-08, 2.69591e-08, 2.703951e-08, 2.592211e-08, 2.517116e-08, 
    2.597372e-08, 2.719664e-08, 2.845839e-08, 2.892494e-08, 2.813793e-08,
  2.414447e-08, 2.480973e-08, 2.513331e-08, 2.565719e-08, 2.582827e-08, 
    2.538015e-08, 2.598592e-08, 2.635286e-08, 2.571648e-08, 2.459194e-08, 
    2.409171e-08, 2.481139e-08, 2.694043e-08, 2.835539e-08, 2.817911e-08,
  2.371076e-08, 2.470336e-08, 2.506387e-08, 2.524401e-08, 2.555161e-08, 
    2.530333e-08, 2.533781e-08, 2.551035e-08, 2.514331e-08, 2.437534e-08, 
    2.355936e-08, 2.304877e-08, 2.463109e-08, 2.744069e-08, 2.790382e-08,
  2.588775e-08, 2.613216e-08, 2.521624e-08, 2.349732e-08, 2.285297e-08, 
    2.273112e-08, 2.36083e-08, 2.451479e-08, 2.564618e-08, 2.628686e-08, 
    2.689663e-08, 2.729237e-08, 2.735239e-08, 2.693019e-08, 2.655828e-08,
  2.58359e-08, 2.590767e-08, 2.552701e-08, 2.423069e-08, 2.294095e-08, 
    2.320846e-08, 2.339158e-08, 2.39988e-08, 2.516498e-08, 2.61634e-08, 
    2.678709e-08, 2.73634e-08, 2.733408e-08, 2.726939e-08, 2.760154e-08,
  2.559737e-08, 2.573677e-08, 2.583457e-08, 2.464107e-08, 2.350126e-08, 
    2.277028e-08, 2.377938e-08, 2.410743e-08, 2.463359e-08, 2.539878e-08, 
    2.611449e-08, 2.689047e-08, 2.758286e-08, 2.798778e-08, 2.795007e-08,
  2.531367e-08, 2.574122e-08, 2.587778e-08, 2.50486e-08, 2.363742e-08, 
    2.288029e-08, 2.370984e-08, 2.465786e-08, 2.519652e-08, 2.551679e-08, 
    2.600146e-08, 2.650432e-08, 2.704206e-08, 2.812638e-08, 2.813294e-08,
  2.523508e-08, 2.587155e-08, 2.586915e-08, 2.539707e-08, 2.420589e-08, 
    2.356187e-08, 2.35535e-08, 2.461151e-08, 2.566581e-08, 2.533729e-08, 
    2.532569e-08, 2.596699e-08, 2.652778e-08, 2.762519e-08, 2.807596e-08,
  2.521824e-08, 2.553767e-08, 2.593995e-08, 2.573183e-08, 2.460354e-08, 
    2.411752e-08, 2.450404e-08, 2.472242e-08, 2.39722e-08, 2.456708e-08, 
    2.667547e-08, 2.739569e-08, 2.698782e-08, 2.752752e-08, 2.81837e-08,
  2.548513e-08, 2.553012e-08, 2.590813e-08, 2.571486e-08, 2.496397e-08, 
    2.454357e-08, 2.475782e-08, 2.505627e-08, 2.424369e-08, 2.58324e-08, 
    2.762441e-08, 2.783977e-08, 2.712519e-08, 2.755033e-08, 2.796022e-08,
  2.578831e-08, 2.561464e-08, 2.552722e-08, 2.57943e-08, 2.53186e-08, 
    2.502384e-08, 2.492355e-08, 2.54478e-08, 2.459596e-08, 2.54893e-08, 
    2.720467e-08, 2.833899e-08, 2.813414e-08, 2.758743e-08, 2.778539e-08,
  2.593785e-08, 2.590243e-08, 2.565287e-08, 2.58807e-08, 2.572562e-08, 
    2.575693e-08, 2.550635e-08, 2.602634e-08, 2.549769e-08, 2.53409e-08, 
    2.602195e-08, 2.74113e-08, 2.796766e-08, 2.770919e-08, 2.748591e-08,
  2.604372e-08, 2.603395e-08, 2.564479e-08, 2.576554e-08, 2.594236e-08, 
    2.588473e-08, 2.598916e-08, 2.631193e-08, 2.579502e-08, 2.487575e-08, 
    2.536028e-08, 2.725123e-08, 2.777474e-08, 2.747536e-08, 2.723375e-08,
  2.45508e-08, 2.425458e-08, 2.34022e-08, 2.307081e-08, 2.336632e-08, 
    2.409798e-08, 2.463179e-08, 2.520075e-08, 2.55589e-08, 2.578417e-08, 
    2.615068e-08, 2.63973e-08, 2.64631e-08, 2.66013e-08, 2.623761e-08,
  2.428442e-08, 2.384396e-08, 2.334211e-08, 2.335334e-08, 2.387149e-08, 
    2.427876e-08, 2.469296e-08, 2.554992e-08, 2.607554e-08, 2.626026e-08, 
    2.636561e-08, 2.647856e-08, 2.637965e-08, 2.640187e-08, 2.656859e-08,
  2.423255e-08, 2.386487e-08, 2.350596e-08, 2.33941e-08, 2.348638e-08, 
    2.363033e-08, 2.450605e-08, 2.556087e-08, 2.631535e-08, 2.641642e-08, 
    2.656544e-08, 2.675401e-08, 2.704886e-08, 2.686066e-08, 2.700994e-08,
  2.41834e-08, 2.390239e-08, 2.37483e-08, 2.358839e-08, 2.387924e-08, 
    2.453205e-08, 2.58385e-08, 2.60786e-08, 2.63236e-08, 2.628222e-08, 
    2.687762e-08, 2.690211e-08, 2.654065e-08, 2.660538e-08, 2.664125e-08,
  2.423302e-08, 2.38825e-08, 2.406352e-08, 2.41722e-08, 2.529834e-08, 
    2.60798e-08, 2.625871e-08, 2.672595e-08, 2.63206e-08, 2.682477e-08, 
    2.703793e-08, 2.682329e-08, 2.685292e-08, 2.71831e-08, 2.662238e-08,
  2.459025e-08, 2.39427e-08, 2.379809e-08, 2.366438e-08, 2.425972e-08, 
    2.495825e-08, 2.515356e-08, 2.465532e-08, 2.612398e-08, 2.762177e-08, 
    2.710049e-08, 2.71321e-08, 2.729238e-08, 2.699579e-08, 2.633758e-08,
  2.484736e-08, 2.417229e-08, 2.387428e-08, 2.363968e-08, 2.408976e-08, 
    2.505485e-08, 2.601408e-08, 2.638213e-08, 2.745589e-08, 2.790187e-08, 
    2.72137e-08, 2.718792e-08, 2.62502e-08, 2.622949e-08, 2.627939e-08,
  2.549436e-08, 2.438761e-08, 2.376824e-08, 2.370745e-08, 2.369553e-08, 
    2.462162e-08, 2.565798e-08, 2.618519e-08, 2.655488e-08, 2.666521e-08, 
    2.668645e-08, 2.629442e-08, 2.588845e-08, 2.619191e-08, 2.631807e-08,
  2.582607e-08, 2.540939e-08, 2.432823e-08, 2.388018e-08, 2.360708e-08, 
    2.397496e-08, 2.470662e-08, 2.561752e-08, 2.63686e-08, 2.682704e-08, 
    2.674294e-08, 2.659713e-08, 2.659003e-08, 2.68027e-08, 2.694894e-08,
  2.54017e-08, 2.606627e-08, 2.534506e-08, 2.467813e-08, 2.403317e-08, 
    2.422266e-08, 2.425887e-08, 2.458785e-08, 2.530445e-08, 2.628897e-08, 
    2.659861e-08, 2.676464e-08, 2.715502e-08, 2.745817e-08, 2.775654e-08,
  2.598157e-08, 2.555016e-08, 2.489618e-08, 2.42067e-08, 2.425415e-08, 
    2.424789e-08, 2.44182e-08, 2.479185e-08, 2.510679e-08, 2.526873e-08, 
    2.532079e-08, 2.535088e-08, 2.557775e-08, 2.570641e-08, 2.598075e-08,
  2.63844e-08, 2.602519e-08, 2.535691e-08, 2.408663e-08, 2.372501e-08, 
    2.453249e-08, 2.489789e-08, 2.49807e-08, 2.514134e-08, 2.520971e-08, 
    2.532132e-08, 2.531514e-08, 2.537805e-08, 2.534669e-08, 2.535161e-08,
  2.670122e-08, 2.652712e-08, 2.627527e-08, 2.467034e-08, 2.27477e-08, 
    2.215842e-08, 2.366327e-08, 2.417536e-08, 2.539446e-08, 2.560765e-08, 
    2.556073e-08, 2.536781e-08, 2.528786e-08, 2.530986e-08, 2.540413e-08,
  2.667778e-08, 2.673166e-08, 2.670685e-08, 2.662123e-08, 2.525247e-08, 
    2.381585e-08, 2.300455e-08, 2.480878e-08, 2.595634e-08, 2.551076e-08, 
    2.567754e-08, 2.556995e-08, 2.551311e-08, 2.519572e-08, 2.497315e-08,
  2.706965e-08, 2.719333e-08, 2.661434e-08, 2.680521e-08, 2.688748e-08, 
    2.654976e-08, 2.727728e-08, 2.804615e-08, 2.52091e-08, 2.484491e-08, 
    2.553416e-08, 2.546476e-08, 2.523684e-08, 2.505453e-08, 2.523046e-08,
  2.688175e-08, 2.776542e-08, 2.739555e-08, 2.709554e-08, 2.697815e-08, 
    2.661245e-08, 2.654871e-08, 2.511295e-08, 2.493539e-08, 2.688727e-08, 
    2.647326e-08, 2.570907e-08, 2.539844e-08, 2.537316e-08, 2.556936e-08,
  2.525011e-08, 2.707473e-08, 2.815597e-08, 2.827391e-08, 2.837487e-08, 
    2.765458e-08, 2.754429e-08, 2.768741e-08, 2.790629e-08, 2.826308e-08, 
    2.595656e-08, 2.574858e-08, 2.567108e-08, 2.588162e-08, 2.603778e-08,
  2.517863e-08, 2.532325e-08, 2.64314e-08, 2.747225e-08, 2.816315e-08, 
    2.797419e-08, 2.736882e-08, 2.736175e-08, 2.705302e-08, 2.702335e-08, 
    2.605041e-08, 2.637838e-08, 2.608965e-08, 2.592661e-08, 2.566466e-08,
  2.579733e-08, 2.539984e-08, 2.573326e-08, 2.608195e-08, 2.677347e-08, 
    2.734137e-08, 2.724355e-08, 2.720397e-08, 2.696291e-08, 2.673609e-08, 
    2.660279e-08, 2.657077e-08, 2.590268e-08, 2.571148e-08, 2.557322e-08,
  2.555947e-08, 2.558713e-08, 2.559216e-08, 2.591785e-08, 2.568885e-08, 
    2.590364e-08, 2.594391e-08, 2.593932e-08, 2.58038e-08, 2.572766e-08, 
    2.574287e-08, 2.57152e-08, 2.579678e-08, 2.610814e-08, 2.657396e-08,
  2.458621e-08, 2.392765e-08, 2.335312e-08, 2.389876e-08, 2.419872e-08, 
    2.40365e-08, 2.419016e-08, 2.449961e-08, 2.47286e-08, 2.50812e-08, 
    2.532798e-08, 2.591625e-08, 2.538694e-08, 2.675032e-08, 2.654366e-08,
  2.602918e-08, 2.452624e-08, 2.292296e-08, 2.232649e-08, 2.324773e-08, 
    2.40756e-08, 2.436609e-08, 2.479225e-08, 2.490959e-08, 2.515123e-08, 
    2.526683e-08, 2.577517e-08, 2.565453e-08, 2.596971e-08, 2.6124e-08,
  2.710885e-08, 2.634617e-08, 2.485826e-08, 2.27702e-08, 2.210712e-08, 
    2.192531e-08, 2.359289e-08, 2.407918e-08, 2.499017e-08, 2.508122e-08, 
    2.505801e-08, 2.542256e-08, 2.574746e-08, 2.605613e-08, 2.585063e-08,
  2.736449e-08, 2.709819e-08, 2.695208e-08, 2.622466e-08, 2.499992e-08, 
    2.329699e-08, 2.238649e-08, 2.459321e-08, 2.524523e-08, 2.540586e-08, 
    2.543233e-08, 2.544815e-08, 2.563681e-08, 2.602819e-08, 2.625468e-08,
  2.750924e-08, 2.699354e-08, 2.720632e-08, 2.720721e-08, 2.7374e-08, 
    2.721416e-08, 2.715549e-08, 2.643392e-08, 2.414885e-08, 2.401049e-08, 
    2.496831e-08, 2.532846e-08, 2.556337e-08, 2.589421e-08, 2.623844e-08,
  2.783497e-08, 2.729686e-08, 2.698271e-08, 2.659165e-08, 2.645486e-08, 
    2.639495e-08, 2.600658e-08, 2.437469e-08, 2.391161e-08, 2.501045e-08, 
    2.584143e-08, 2.548903e-08, 2.545761e-08, 2.567825e-08, 2.595818e-08,
  2.714229e-08, 2.755426e-08, 2.714392e-08, 2.693423e-08, 2.659935e-08, 
    2.682888e-08, 2.693214e-08, 2.751056e-08, 2.771671e-08, 2.720019e-08, 
    2.575784e-08, 2.543389e-08, 2.543292e-08, 2.572773e-08, 2.597471e-08,
  2.665136e-08, 2.752421e-08, 2.767099e-08, 2.734038e-08, 2.649931e-08, 
    2.597832e-08, 2.562919e-08, 2.543076e-08, 2.552868e-08, 2.555864e-08, 
    2.529393e-08, 2.531798e-08, 2.537956e-08, 2.562182e-08, 2.575508e-08,
  2.57349e-08, 2.666147e-08, 2.776217e-08, 2.840154e-08, 2.778468e-08, 
    2.693799e-08, 2.615903e-08, 2.586814e-08, 2.52594e-08, 2.530004e-08, 
    2.515763e-08, 2.529567e-08, 2.541301e-08, 2.577189e-08, 2.590266e-08,
  2.533545e-08, 2.528848e-08, 2.643617e-08, 2.797869e-08, 2.84992e-08, 
    2.808039e-08, 2.708478e-08, 2.636682e-08, 2.593893e-08, 2.565915e-08, 
    2.546072e-08, 2.538748e-08, 2.554067e-08, 2.548193e-08, 2.551726e-08,
  2.455569e-08, 2.406786e-08, 2.398293e-08, 2.493089e-08, 2.584005e-08, 
    2.645433e-08, 2.550215e-08, 2.47899e-08, 2.443379e-08, 2.440044e-08, 
    2.502242e-08, 2.535954e-08, 2.523151e-08, 2.55557e-08, 2.488138e-08,
  2.572482e-08, 2.511884e-08, 2.414229e-08, 2.402941e-08, 2.477841e-08, 
    2.485912e-08, 2.465893e-08, 2.444119e-08, 2.422246e-08, 2.447494e-08, 
    2.499507e-08, 2.559603e-08, 2.535116e-08, 2.470943e-08, 2.441463e-08,
  2.60303e-08, 2.566158e-08, 2.52874e-08, 2.422501e-08, 2.39841e-08, 
    2.403979e-08, 2.463594e-08, 2.387668e-08, 2.390026e-08, 2.427424e-08, 
    2.483641e-08, 2.552446e-08, 2.548494e-08, 2.511246e-08, 2.516503e-08,
  2.651569e-08, 2.579109e-08, 2.579432e-08, 2.531576e-08, 2.461797e-08, 
    2.397611e-08, 2.398185e-08, 2.451346e-08, 2.425886e-08, 2.419612e-08, 
    2.472882e-08, 2.555069e-08, 2.553063e-08, 2.547258e-08, 2.578496e-08,
  2.718533e-08, 2.640247e-08, 2.573453e-08, 2.58239e-08, 2.547226e-08, 
    2.505053e-08, 2.427329e-08, 2.447472e-08, 2.401513e-08, 2.457974e-08, 
    2.472684e-08, 2.539455e-08, 2.562438e-08, 2.554098e-08, 2.590657e-08,
  2.773549e-08, 2.726988e-08, 2.636174e-08, 2.583945e-08, 2.555198e-08, 
    2.546071e-08, 2.506423e-08, 2.460342e-08, 2.416852e-08, 2.470044e-08, 
    2.47719e-08, 2.519358e-08, 2.551234e-08, 2.551401e-08, 2.581262e-08,
  2.746093e-08, 2.774395e-08, 2.736595e-08, 2.662223e-08, 2.60095e-08, 
    2.569091e-08, 2.550984e-08, 2.549776e-08, 2.486585e-08, 2.478427e-08, 
    2.472886e-08, 2.51349e-08, 2.547559e-08, 2.555951e-08, 2.55594e-08,
  2.547111e-08, 2.700578e-08, 2.742154e-08, 2.744043e-08, 2.671695e-08, 
    2.61605e-08, 2.542232e-08, 2.528627e-08, 2.535262e-08, 2.529431e-08, 
    2.514217e-08, 2.51281e-08, 2.530411e-08, 2.556009e-08, 2.535593e-08,
  2.476833e-08, 2.52683e-08, 2.645442e-08, 2.717855e-08, 2.754145e-08, 
    2.718986e-08, 2.653295e-08, 2.575178e-08, 2.542676e-08, 2.511819e-08, 
    2.501792e-08, 2.545557e-08, 2.536438e-08, 2.574866e-08, 2.522676e-08,
  2.471874e-08, 2.476699e-08, 2.521373e-08, 2.589419e-08, 2.64962e-08, 
    2.72517e-08, 2.726937e-08, 2.67109e-08, 2.606652e-08, 2.559024e-08, 
    2.527985e-08, 2.548933e-08, 2.535638e-08, 2.587402e-08, 2.525791e-08,
  2.473063e-08, 2.576881e-08, 2.691172e-08, 2.757696e-08, 2.785263e-08, 
    2.77705e-08, 2.743447e-08, 2.740244e-08, 2.741921e-08, 2.712228e-08, 
    2.726444e-08, 2.708512e-08, 2.72023e-08, 2.707952e-08, 2.689179e-08,
  2.427602e-08, 2.460921e-08, 2.490028e-08, 2.572532e-08, 2.631157e-08, 
    2.663909e-08, 2.689521e-08, 2.678521e-08, 2.694144e-08, 2.710726e-08, 
    2.693575e-08, 2.667547e-08, 2.679491e-08, 2.703622e-08, 2.687139e-08,
  2.49622e-08, 2.453752e-08, 2.458269e-08, 2.454774e-08, 2.507888e-08, 
    2.497008e-08, 2.584761e-08, 2.59505e-08, 2.632476e-08, 2.634737e-08, 
    2.652723e-08, 2.655101e-08, 2.641394e-08, 2.598889e-08, 2.613599e-08,
  2.607376e-08, 2.505039e-08, 2.476783e-08, 2.447682e-08, 2.449176e-08, 
    2.402661e-08, 2.413695e-08, 2.533914e-08, 2.503598e-08, 2.575086e-08, 
    2.599431e-08, 2.599414e-08, 2.566676e-08, 2.478948e-08, 2.485846e-08,
  2.66535e-08, 2.61116e-08, 2.52615e-08, 2.473801e-08, 2.462816e-08, 
    2.440941e-08, 2.390369e-08, 2.386479e-08, 2.51892e-08, 2.525203e-08, 
    2.524885e-08, 2.542034e-08, 2.497127e-08, 2.447137e-08, 2.513814e-08,
  2.549459e-08, 2.66341e-08, 2.634093e-08, 2.537232e-08, 2.48836e-08, 
    2.458701e-08, 2.426472e-08, 2.427889e-08, 2.425331e-08, 2.451304e-08, 
    2.4445e-08, 2.49565e-08, 2.454173e-08, 2.469026e-08, 2.521308e-08,
  2.405836e-08, 2.503406e-08, 2.656079e-08, 2.646484e-08, 2.545829e-08, 
    2.510199e-08, 2.43285e-08, 2.404289e-08, 2.382273e-08, 2.415389e-08, 
    2.400838e-08, 2.429935e-08, 2.427781e-08, 2.55449e-08, 2.593519e-08,
  2.497795e-08, 2.378829e-08, 2.438579e-08, 2.634451e-08, 2.64126e-08, 
    2.586158e-08, 2.53214e-08, 2.467592e-08, 2.403077e-08, 2.359155e-08, 
    2.339982e-08, 2.439816e-08, 2.46355e-08, 2.545092e-08, 2.575513e-08,
  2.698386e-08, 2.513082e-08, 2.356404e-08, 2.395062e-08, 2.568071e-08, 
    2.634976e-08, 2.594147e-08, 2.542898e-08, 2.468823e-08, 2.428177e-08, 
    2.448306e-08, 2.519408e-08, 2.559827e-08, 2.576516e-08, 2.584859e-08,
  2.695264e-08, 2.701103e-08, 2.485562e-08, 2.356488e-08, 2.376841e-08, 
    2.526043e-08, 2.638868e-08, 2.650357e-08, 2.56803e-08, 2.512907e-08, 
    2.483945e-08, 2.54457e-08, 2.570991e-08, 2.613489e-08, 2.596502e-08,
  2.363979e-08, 2.48419e-08, 2.471148e-08, 2.633508e-08, 2.708641e-08, 
    2.731507e-08, 2.695171e-08, 2.687312e-08, 2.656222e-08, 2.687053e-08, 
    2.707355e-08, 2.745028e-08, 2.767458e-08, 2.753924e-08, 2.746174e-08,
  2.35002e-08, 2.420382e-08, 2.447169e-08, 2.545567e-08, 2.649299e-08, 
    2.704685e-08, 2.782976e-08, 2.684529e-08, 2.711527e-08, 2.69688e-08, 
    2.719781e-08, 2.751634e-08, 2.773484e-08, 2.779753e-08, 2.753415e-08,
  2.371684e-08, 2.395204e-08, 2.440802e-08, 2.531684e-08, 2.610005e-08, 
    2.716265e-08, 2.712978e-08, 2.71979e-08, 2.720586e-08, 2.709785e-08, 
    2.703646e-08, 2.74645e-08, 2.780548e-08, 2.794439e-08, 2.7922e-08,
  2.467287e-08, 2.377786e-08, 2.427173e-08, 2.505116e-08, 2.584424e-08, 
    2.675129e-08, 2.71061e-08, 2.75043e-08, 2.763762e-08, 2.739128e-08, 
    2.748141e-08, 2.767985e-08, 2.783771e-08, 2.802842e-08, 2.77671e-08,
  2.576593e-08, 2.441686e-08, 2.424128e-08, 2.491828e-08, 2.549963e-08, 
    2.609143e-08, 2.622451e-08, 2.669976e-08, 2.662455e-08, 2.651465e-08, 
    2.638321e-08, 2.766092e-08, 2.794109e-08, 2.800006e-08, 2.77565e-08,
  2.55505e-08, 2.56014e-08, 2.4583e-08, 2.466253e-08, 2.515442e-08, 
    2.582822e-08, 2.586637e-08, 2.564724e-08, 2.549935e-08, 2.622344e-08, 
    2.783241e-08, 2.884804e-08, 2.765418e-08, 2.779891e-08, 2.75858e-08,
  2.491535e-08, 2.564789e-08, 2.562672e-08, 2.507223e-08, 2.49624e-08, 
    2.552862e-08, 2.651822e-08, 2.735944e-08, 2.808282e-08, 2.892098e-08, 
    2.929588e-08, 2.762976e-08, 2.760435e-08, 2.777026e-08, 2.755373e-08,
  2.412548e-08, 2.499231e-08, 2.555932e-08, 2.565401e-08, 2.519358e-08, 
    2.49692e-08, 2.535357e-08, 2.602239e-08, 2.676451e-08, 2.768106e-08, 
    2.761584e-08, 2.711647e-08, 2.761467e-08, 2.717834e-08, 2.739052e-08,
  2.40219e-08, 2.428728e-08, 2.524865e-08, 2.582466e-08, 2.583641e-08, 
    2.568664e-08, 2.54681e-08, 2.586242e-08, 2.610426e-08, 2.660674e-08, 
    2.650516e-08, 2.704729e-08, 2.691114e-08, 2.706567e-08, 2.725543e-08,
  2.417673e-08, 2.375416e-08, 2.392397e-08, 2.495774e-08, 2.548573e-08, 
    2.592443e-08, 2.586537e-08, 2.581984e-08, 2.612102e-08, 2.648604e-08, 
    2.628832e-08, 2.646566e-08, 2.666312e-08, 2.692183e-08, 2.686102e-08,
  2.515443e-08, 2.642891e-08, 2.734596e-08, 2.779095e-08, 2.77275e-08, 
    2.789508e-08, 2.753836e-08, 2.697056e-08, 2.639735e-08, 2.563417e-08, 
    2.543399e-08, 2.558078e-08, 2.578012e-08, 2.596835e-08, 2.636842e-08,
  2.63903e-08, 2.740363e-08, 2.779232e-08, 2.804217e-08, 2.779888e-08, 
    2.738569e-08, 2.783578e-08, 2.73025e-08, 2.678115e-08, 2.604597e-08, 
    2.589156e-08, 2.579259e-08, 2.594028e-08, 2.607271e-08, 2.6304e-08,
  2.674469e-08, 2.735073e-08, 2.768367e-08, 2.735866e-08, 2.801712e-08, 
    2.736159e-08, 2.754064e-08, 2.68437e-08, 2.661704e-08, 2.595411e-08, 
    2.577148e-08, 2.604323e-08, 2.628631e-08, 2.671224e-08, 2.702468e-08,
  2.708792e-08, 2.732939e-08, 2.745398e-08, 2.711016e-08, 2.720389e-08, 
    2.730382e-08, 2.717915e-08, 2.72904e-08, 2.664731e-08, 2.64686e-08, 
    2.641037e-08, 2.657839e-08, 2.653246e-08, 2.675494e-08, 2.688643e-08,
  2.705377e-08, 2.691388e-08, 2.700208e-08, 2.66928e-08, 2.657779e-08, 
    2.675418e-08, 2.670372e-08, 2.64708e-08, 2.559355e-08, 2.529206e-08, 
    2.654295e-08, 2.66876e-08, 2.700179e-08, 2.749458e-08, 2.74615e-08,
  2.73912e-08, 2.694302e-08, 2.702885e-08, 2.648948e-08, 2.582753e-08, 
    2.498566e-08, 2.47393e-08, 2.491838e-08, 2.532484e-08, 2.714067e-08, 
    2.794104e-08, 2.761116e-08, 2.768179e-08, 2.785042e-08, 2.763128e-08,
  2.748009e-08, 2.743127e-08, 2.779262e-08, 2.792043e-08, 2.762424e-08, 
    2.745651e-08, 2.737742e-08, 2.767583e-08, 2.832996e-08, 2.887809e-08, 
    2.741782e-08, 2.746697e-08, 2.750066e-08, 2.788317e-08, 2.760883e-08,
  2.717294e-08, 2.751707e-08, 2.777889e-08, 2.824635e-08, 2.870478e-08, 
    2.889513e-08, 2.915037e-08, 2.905764e-08, 2.898379e-08, 2.865732e-08, 
    2.808954e-08, 2.828239e-08, 2.814516e-08, 2.830498e-08, 2.758177e-08,
  2.633061e-08, 2.684785e-08, 2.704712e-08, 2.727636e-08, 2.74035e-08, 
    2.759455e-08, 2.770962e-08, 2.788571e-08, 2.782068e-08, 2.772452e-08, 
    2.766324e-08, 2.745293e-08, 2.726558e-08, 2.695145e-08, 2.648951e-08,
  2.527126e-08, 2.585044e-08, 2.650282e-08, 2.683159e-08, 2.709722e-08, 
    2.728602e-08, 2.751172e-08, 2.757578e-08, 2.780874e-08, 2.759265e-08, 
    2.778328e-08, 2.741814e-08, 2.726978e-08, 2.711104e-08, 2.687127e-08,
  2.750295e-08, 2.724872e-08, 2.748001e-08, 2.740448e-08, 2.775126e-08, 
    2.777264e-08, 2.780937e-08, 2.765552e-08, 2.767659e-08, 2.695656e-08, 
    2.673835e-08, 2.632242e-08, 2.67442e-08, 2.678197e-08, 2.733215e-08,
  2.791108e-08, 2.784275e-08, 2.777145e-08, 2.816397e-08, 2.779523e-08, 
    2.834392e-08, 2.806202e-08, 2.820659e-08, 2.79897e-08, 2.751729e-08, 
    2.70303e-08, 2.644064e-08, 2.66762e-08, 2.648349e-08, 2.663705e-08,
  2.679452e-08, 2.694943e-08, 2.729056e-08, 2.707053e-08, 2.804091e-08, 
    2.740176e-08, 2.843591e-08, 2.788938e-08, 2.779601e-08, 2.744412e-08, 
    2.697069e-08, 2.621117e-08, 2.623588e-08, 2.614249e-08, 2.63749e-08,
  2.638513e-08, 2.649693e-08, 2.721429e-08, 2.734168e-08, 2.759564e-08, 
    2.754176e-08, 2.757936e-08, 2.83486e-08, 2.759728e-08, 2.663497e-08, 
    2.595056e-08, 2.564503e-08, 2.547729e-08, 2.562387e-08, 2.581519e-08,
  2.64048e-08, 2.619335e-08, 2.686018e-08, 2.665327e-08, 2.679505e-08, 
    2.670216e-08, 2.66411e-08, 2.647702e-08, 2.612782e-08, 2.569559e-08, 
    2.517428e-08, 2.499132e-08, 2.517639e-08, 2.551229e-08, 2.582729e-08,
  2.694249e-08, 2.597871e-08, 2.625308e-08, 2.578381e-08, 2.618554e-08, 
    2.595307e-08, 2.604032e-08, 2.598998e-08, 2.601992e-08, 2.541199e-08, 
    2.527526e-08, 2.536947e-08, 2.568642e-08, 2.552214e-08, 2.596041e-08,
  2.816747e-08, 2.757623e-08, 2.73526e-08, 2.680604e-08, 2.66204e-08, 
    2.632424e-08, 2.622027e-08, 2.613759e-08, 2.603682e-08, 2.617044e-08, 
    2.591648e-08, 2.623818e-08, 2.593355e-08, 2.624262e-08, 2.63461e-08,
  2.72864e-08, 2.779917e-08, 2.782836e-08, 2.796406e-08, 2.774645e-08, 
    2.765208e-08, 2.750538e-08, 2.745013e-08, 2.738971e-08, 2.735593e-08, 
    2.738404e-08, 2.735624e-08, 2.720419e-08, 2.726671e-08, 2.699811e-08,
  2.483282e-08, 2.561845e-08, 2.622393e-08, 2.658627e-08, 2.692067e-08, 
    2.709259e-08, 2.744921e-08, 2.751846e-08, 2.76077e-08, 2.757004e-08, 
    2.746679e-08, 2.749342e-08, 2.734033e-08, 2.737081e-08, 2.701226e-08,
  2.326074e-08, 2.361477e-08, 2.406978e-08, 2.448023e-08, 2.499415e-08, 
    2.529944e-08, 2.574354e-08, 2.596459e-08, 2.633053e-08, 2.657869e-08, 
    2.678663e-08, 2.688079e-08, 2.710562e-08, 2.687538e-08, 2.711171e-08,
  2.685746e-08, 2.706585e-08, 2.707891e-08, 2.756391e-08, 2.757194e-08, 
    2.782464e-08, 2.825089e-08, 2.803962e-08, 2.83022e-08, 2.826844e-08, 
    2.841899e-08, 2.804403e-08, 2.809122e-08, 2.743732e-08, 2.702588e-08,
  2.656855e-08, 2.704394e-08, 2.727907e-08, 2.776667e-08, 2.804959e-08, 
    2.7767e-08, 2.833059e-08, 2.797235e-08, 2.831652e-08, 2.826166e-08, 
    2.847956e-08, 2.805187e-08, 2.831422e-08, 2.773131e-08, 2.729993e-08,
  2.685191e-08, 2.696114e-08, 2.789049e-08, 2.738183e-08, 2.822527e-08, 
    2.788043e-08, 2.820143e-08, 2.827815e-08, 2.831774e-08, 2.820837e-08, 
    2.837897e-08, 2.813022e-08, 2.786322e-08, 2.778644e-08, 2.730426e-08,
  2.697619e-08, 2.709028e-08, 2.804973e-08, 2.741782e-08, 2.842536e-08, 
    2.798509e-08, 2.780835e-08, 2.860068e-08, 2.864732e-08, 2.814945e-08, 
    2.8204e-08, 2.774552e-08, 2.74827e-08, 2.751905e-08, 2.702195e-08,
  2.673961e-08, 2.646626e-08, 2.695505e-08, 2.686699e-08, 2.743738e-08, 
    2.718378e-08, 2.671296e-08, 2.727746e-08, 2.767043e-08, 2.712682e-08, 
    2.62915e-08, 2.59848e-08, 2.600789e-08, 2.664098e-08, 2.649715e-08,
  2.683118e-08, 2.659835e-08, 2.675223e-08, 2.632761e-08, 2.641272e-08, 
    2.603473e-08, 2.645443e-08, 2.643078e-08, 2.588382e-08, 2.486821e-08, 
    2.531899e-08, 2.524861e-08, 2.548403e-08, 2.538454e-08, 2.583528e-08,
  2.64331e-08, 2.648095e-08, 2.653152e-08, 2.671401e-08, 2.668515e-08, 
    2.677311e-08, 2.634393e-08, 2.604535e-08, 2.560783e-08, 2.549846e-08, 
    2.537049e-08, 2.536903e-08, 2.535753e-08, 2.559567e-08, 2.608058e-08,
  2.580832e-08, 2.62015e-08, 2.620678e-08, 2.645467e-08, 2.658849e-08, 
    2.705434e-08, 2.745409e-08, 2.749031e-08, 2.747195e-08, 2.700655e-08, 
    2.661059e-08, 2.595512e-08, 2.600305e-08, 2.579202e-08, 2.568835e-08,
  2.642437e-08, 2.591866e-08, 2.572364e-08, 2.552409e-08, 2.547092e-08, 
    2.555446e-08, 2.6041e-08, 2.654993e-08, 2.729544e-08, 2.734753e-08, 
    2.732623e-08, 2.713804e-08, 2.652652e-08, 2.622932e-08, 2.575573e-08,
  2.72944e-08, 2.707508e-08, 2.652308e-08, 2.636122e-08, 2.60041e-08, 
    2.554473e-08, 2.51158e-08, 2.495718e-08, 2.59103e-08, 2.661586e-08, 
    2.727212e-08, 2.714692e-08, 2.65855e-08, 2.648329e-08, 2.660979e-08,
  2.667798e-08, 2.671768e-08, 2.672752e-08, 2.681319e-08, 2.672787e-08, 
    2.683339e-08, 2.677483e-08, 2.692777e-08, 2.701047e-08, 2.720695e-08, 
    2.727677e-08, 2.75078e-08, 2.769463e-08, 2.782313e-08, 2.774318e-08,
  2.700706e-08, 2.677506e-08, 2.720905e-08, 2.706209e-08, 2.732166e-08, 
    2.726942e-08, 2.77806e-08, 2.788607e-08, 2.797638e-08, 2.796698e-08, 
    2.805058e-08, 2.789778e-08, 2.812326e-08, 2.7999e-08, 2.790548e-08,
  2.681308e-08, 2.694994e-08, 2.71385e-08, 2.693143e-08, 2.73485e-08, 
    2.732056e-08, 2.74949e-08, 2.79051e-08, 2.791621e-08, 2.831581e-08, 
    2.820078e-08, 2.831024e-08, 2.828972e-08, 2.849243e-08, 2.848057e-08,
  2.723404e-08, 2.706862e-08, 2.712929e-08, 2.690103e-08, 2.709222e-08, 
    2.730137e-08, 2.637284e-08, 2.744087e-08, 2.821332e-08, 2.833037e-08, 
    2.84326e-08, 2.857599e-08, 2.836715e-08, 2.787192e-08, 2.785394e-08,
  2.715685e-08, 2.704067e-08, 2.699164e-08, 2.688911e-08, 2.662615e-08, 
    2.672943e-08, 2.680934e-08, 2.565358e-08, 2.789407e-08, 2.823978e-08, 
    2.738281e-08, 2.734196e-08, 2.703197e-08, 2.735061e-08, 2.710313e-08,
  2.720651e-08, 2.715209e-08, 2.720948e-08, 2.670365e-08, 2.6823e-08, 
    2.66941e-08, 2.677013e-08, 2.659037e-08, 2.524622e-08, 2.558614e-08, 
    2.615463e-08, 2.580215e-08, 2.614218e-08, 2.627536e-08, 2.646613e-08,
  2.708227e-08, 2.703765e-08, 2.713841e-08, 2.695374e-08, 2.634132e-08, 
    2.687988e-08, 2.648397e-08, 2.620865e-08, 2.584161e-08, 2.572401e-08, 
    2.54987e-08, 2.558931e-08, 2.580381e-08, 2.638142e-08, 2.647146e-08,
  2.700878e-08, 2.701189e-08, 2.749234e-08, 2.712612e-08, 2.651737e-08, 
    2.658743e-08, 2.732743e-08, 2.69316e-08, 2.635343e-08, 2.567999e-08, 
    2.554087e-08, 2.566779e-08, 2.617403e-08, 2.628711e-08, 2.671782e-08,
  2.691326e-08, 2.665718e-08, 2.756717e-08, 2.760307e-08, 2.658497e-08, 
    2.598256e-08, 2.584622e-08, 2.605985e-08, 2.537105e-08, 2.53119e-08, 
    2.580969e-08, 2.580085e-08, 2.582338e-08, 2.624652e-08, 2.68238e-08,
  2.698917e-08, 2.651836e-08, 2.718175e-08, 2.758471e-08, 2.707062e-08, 
    2.64033e-08, 2.622529e-08, 2.663233e-08, 2.735689e-08, 2.659714e-08, 
    2.581772e-08, 2.581617e-08, 2.60616e-08, 2.676035e-08, 2.730753e-08,
  2.398402e-08, 2.486742e-08, 2.548562e-08, 2.587679e-08, 2.626321e-08, 
    2.690645e-08, 2.722708e-08, 2.712466e-08, 2.691474e-08, 2.675697e-08, 
    2.698968e-08, 2.706954e-08, 2.7368e-08, 2.72473e-08, 2.729734e-08,
  2.506909e-08, 2.530312e-08, 2.578756e-08, 2.613871e-08, 2.704637e-08, 
    2.721641e-08, 2.719878e-08, 2.696768e-08, 2.684905e-08, 2.723731e-08, 
    2.756442e-08, 2.787297e-08, 2.832543e-08, 2.80613e-08, 2.803418e-08,
  2.511361e-08, 2.53222e-08, 2.605615e-08, 2.67819e-08, 2.746839e-08, 
    2.712619e-08, 2.657594e-08, 2.674832e-08, 2.687042e-08, 2.706413e-08, 
    2.727024e-08, 2.816586e-08, 2.827043e-08, 2.832279e-08, 2.843184e-08,
  2.546293e-08, 2.58249e-08, 2.674505e-08, 2.725135e-08, 2.768308e-08, 
    2.727813e-08, 2.642887e-08, 2.626705e-08, 2.62709e-08, 2.6957e-08, 
    2.729479e-08, 2.824558e-08, 2.852854e-08, 2.827506e-08, 2.829487e-08,
  2.602183e-08, 2.641385e-08, 2.72286e-08, 2.753846e-08, 2.713257e-08, 
    2.637323e-08, 2.714037e-08, 2.560307e-08, 2.577732e-08, 2.757905e-08, 
    2.664001e-08, 2.723716e-08, 2.729581e-08, 2.734564e-08, 2.687828e-08,
  2.683606e-08, 2.691162e-08, 2.737672e-08, 2.716047e-08, 2.689844e-08, 
    2.650356e-08, 2.606545e-08, 2.664424e-08, 2.668619e-08, 2.64003e-08, 
    2.645737e-08, 2.610343e-08, 2.635644e-08, 2.563068e-08, 2.523511e-08,
  2.692548e-08, 2.669427e-08, 2.700051e-08, 2.69908e-08, 2.695112e-08, 
    2.636597e-08, 2.580814e-08, 2.422962e-08, 2.620765e-08, 2.720668e-08, 
    2.657939e-08, 2.599391e-08, 2.501929e-08, 2.390393e-08, 2.315698e-08,
  2.707546e-08, 2.658179e-08, 2.716009e-08, 2.703859e-08, 2.742838e-08, 
    2.671661e-08, 2.499532e-08, 2.316357e-08, 2.329682e-08, 2.633466e-08, 
    2.676125e-08, 2.646859e-08, 2.572312e-08, 2.465291e-08, 2.432447e-08,
  2.632008e-08, 2.615627e-08, 2.690851e-08, 2.732899e-08, 2.817038e-08, 
    2.797197e-08, 2.426126e-08, 2.003168e-08, 2.014443e-08, 2.475544e-08, 
    2.673821e-08, 2.731903e-08, 2.716136e-08, 2.678658e-08, 2.663688e-08,
  2.627287e-08, 2.598081e-08, 2.68199e-08, 2.726999e-08, 2.932639e-08, 
    2.979768e-08, 2.936582e-08, 2.769169e-08, 2.772566e-08, 2.630973e-08, 
    2.688372e-08, 2.832448e-08, 2.843394e-08, 2.821664e-08, 2.782413e-08,
  2.166607e-08, 2.182344e-08, 2.213988e-08, 2.237832e-08, 2.2687e-08, 
    2.293918e-08, 2.352767e-08, 2.421116e-08, 2.505244e-08, 2.573423e-08, 
    2.598629e-08, 2.615088e-08, 2.625823e-08, 2.665262e-08, 2.696015e-08,
  2.335218e-08, 2.37548e-08, 2.397483e-08, 2.409567e-08, 2.422897e-08, 
    2.45481e-08, 2.495849e-08, 2.559934e-08, 2.607829e-08, 2.61297e-08, 
    2.612947e-08, 2.618541e-08, 2.651584e-08, 2.681292e-08, 2.703107e-08,
  2.513922e-08, 2.478403e-08, 2.44469e-08, 2.432746e-08, 2.462235e-08, 
    2.501677e-08, 2.533644e-08, 2.610406e-08, 2.614474e-08, 2.619123e-08, 
    2.623152e-08, 2.635016e-08, 2.650743e-08, 2.672837e-08, 2.70411e-08,
  2.405253e-08, 2.386605e-08, 2.419858e-08, 2.483886e-08, 2.537244e-08, 
    2.62232e-08, 2.610989e-08, 2.670314e-08, 2.581792e-08, 2.617809e-08, 
    2.624519e-08, 2.641421e-08, 2.603865e-08, 2.547437e-08, 2.576762e-08,
  2.459074e-08, 2.542916e-08, 2.625255e-08, 2.660175e-08, 2.668695e-08, 
    2.677299e-08, 2.740226e-08, 2.591756e-08, 2.496039e-08, 2.618921e-08, 
    2.66643e-08, 2.554384e-08, 2.359574e-08, 2.393603e-08, 2.499973e-08,
  2.620306e-08, 2.662131e-08, 2.65853e-08, 2.622221e-08, 2.65227e-08, 
    2.713866e-08, 2.689212e-08, 2.570287e-08, 2.590047e-08, 2.661131e-08, 
    2.598034e-08, 2.299867e-08, 2.293587e-08, 2.489614e-08, 2.654652e-08,
  2.705275e-08, 2.653941e-08, 2.616611e-08, 2.633024e-08, 2.774847e-08, 
    2.788967e-08, 2.625583e-08, 2.221358e-08, 2.436805e-08, 2.694103e-08, 
    2.494218e-08, 2.388334e-08, 2.480751e-08, 2.612975e-08, 2.71166e-08,
  2.562755e-08, 2.519207e-08, 2.6146e-08, 2.7517e-08, 2.88779e-08, 
    2.851607e-08, 2.395648e-08, 2.208461e-08, 2.541429e-08, 2.595082e-08, 
    2.518897e-08, 2.528291e-08, 2.622078e-08, 2.73127e-08, 2.824233e-08,
  2.509691e-08, 2.607086e-08, 2.728032e-08, 2.854641e-08, 3.029193e-08, 
    2.783711e-08, 2.290897e-08, 2.258095e-08, 2.574171e-08, 2.633555e-08, 
    2.611517e-08, 2.633738e-08, 2.712108e-08, 2.800573e-08, 2.846801e-08,
  2.557214e-08, 2.584975e-08, 2.734213e-08, 2.946475e-08, 3.126778e-08, 
    2.898657e-08, 2.784565e-08, 2.731652e-08, 2.675353e-08, 2.617028e-08, 
    2.621655e-08, 2.639227e-08, 2.69012e-08, 2.732117e-08, 2.727405e-08,
  2.445079e-08, 2.412195e-08, 2.351428e-08, 2.332559e-08, 2.300709e-08, 
    2.316153e-08, 2.309276e-08, 2.324087e-08, 2.320919e-08, 2.325321e-08, 
    2.338119e-08, 2.343882e-08, 2.380028e-08, 2.425379e-08, 2.470144e-08,
  2.534291e-08, 2.531908e-08, 2.516457e-08, 2.485449e-08, 2.458547e-08, 
    2.420106e-08, 2.436e-08, 2.412688e-08, 2.436726e-08, 2.432171e-08, 
    2.491259e-08, 2.477442e-08, 2.571953e-08, 2.570826e-08, 2.583513e-08,
  2.478948e-08, 2.504358e-08, 2.515134e-08, 2.512318e-08, 2.526026e-08, 
    2.513606e-08, 2.50835e-08, 2.498535e-08, 2.501498e-08, 2.510135e-08, 
    2.529182e-08, 2.535119e-08, 2.555655e-08, 2.547501e-08, 2.567343e-08,
  2.459247e-08, 2.437367e-08, 2.468073e-08, 2.440335e-08, 2.462238e-08, 
    2.475577e-08, 2.465135e-08, 2.494144e-08, 2.498466e-08, 2.532489e-08, 
    2.53996e-08, 2.548892e-08, 2.560829e-08, 2.553167e-08, 2.568927e-08,
  2.494778e-08, 2.506468e-08, 2.502965e-08, 2.519488e-08, 2.507973e-08, 
    2.543097e-08, 2.596875e-08, 2.621623e-08, 2.574655e-08, 2.635769e-08, 
    2.590158e-08, 2.619003e-08, 2.592159e-08, 2.520075e-08, 2.444639e-08,
  2.659919e-08, 2.654975e-08, 2.644863e-08, 2.629836e-08, 2.627757e-08, 
    2.631329e-08, 2.637396e-08, 2.654976e-08, 2.652203e-08, 2.580209e-08, 
    2.590961e-08, 2.510948e-08, 2.452798e-08, 2.446603e-08, 2.521345e-08,
  2.645806e-08, 2.596176e-08, 2.582733e-08, 2.573813e-08, 2.599431e-08, 
    2.65582e-08, 2.697941e-08, 2.628861e-08, 2.546166e-08, 2.520996e-08, 
    2.498861e-08, 2.52421e-08, 2.557036e-08, 2.66388e-08, 2.680349e-08,
  2.567229e-08, 2.533307e-08, 2.58132e-08, 2.708637e-08, 2.698356e-08, 
    2.755355e-08, 2.660412e-08, 2.54802e-08, 2.581744e-08, 2.508502e-08, 
    2.607113e-08, 2.660021e-08, 2.726006e-08, 2.796617e-08, 2.787765e-08,
  2.567822e-08, 2.663052e-08, 2.812935e-08, 2.976558e-08, 2.981848e-08, 
    2.736704e-08, 2.539046e-08, 2.505626e-08, 2.563343e-08, 2.691515e-08, 
    2.780986e-08, 2.849187e-08, 2.918582e-08, 2.898629e-08, 2.86798e-08,
  2.667972e-08, 2.8958e-08, 3.077385e-08, 3.086523e-08, 2.832154e-08, 
    2.584583e-08, 2.561669e-08, 2.587915e-08, 2.768947e-08, 2.88473e-08, 
    2.931354e-08, 2.987408e-08, 2.945862e-08, 2.922693e-08, 2.903467e-08,
  2.47803e-08, 2.502374e-08, 2.461913e-08, 2.388615e-08, 2.259742e-08, 
    2.186407e-08, 2.205293e-08, 2.244387e-08, 2.351061e-08, 2.385679e-08, 
    2.433926e-08, 2.452804e-08, 2.463916e-08, 2.475085e-08, 2.450539e-08,
  2.548122e-08, 2.494498e-08, 2.49348e-08, 2.479003e-08, 2.412468e-08, 
    2.332116e-08, 2.256462e-08, 2.222154e-08, 2.243087e-08, 2.294584e-08, 
    2.321197e-08, 2.351132e-08, 2.374345e-08, 2.386972e-08, 2.367501e-08,
  2.62799e-08, 2.548082e-08, 2.481982e-08, 2.452283e-08, 2.462601e-08, 
    2.406206e-08, 2.388461e-08, 2.380839e-08, 2.340251e-08, 2.3311e-08, 
    2.337529e-08, 2.342601e-08, 2.369454e-08, 2.370787e-08, 2.407079e-08,
  2.747557e-08, 2.622718e-08, 2.600779e-08, 2.437451e-08, 2.479766e-08, 
    2.440905e-08, 2.415496e-08, 2.437113e-08, 2.463714e-08, 2.451138e-08, 
    2.460713e-08, 2.449682e-08, 2.468437e-08, 2.447548e-08, 2.490749e-08,
  2.750624e-08, 2.67436e-08, 2.632241e-08, 2.536685e-08, 2.437841e-08, 
    2.458763e-08, 2.433632e-08, 2.368206e-08, 2.388121e-08, 2.405739e-08, 
    2.418746e-08, 2.446282e-08, 2.430405e-08, 2.497098e-08, 2.47728e-08,
  2.762831e-08, 2.731877e-08, 2.687054e-08, 2.646412e-08, 2.601388e-08, 
    2.489536e-08, 2.538702e-08, 2.505449e-08, 2.484304e-08, 2.470696e-08, 
    2.475333e-08, 2.502838e-08, 2.518642e-08, 2.543298e-08, 2.530932e-08,
  2.673456e-08, 2.663812e-08, 2.68923e-08, 2.643251e-08, 2.661161e-08, 
    2.586688e-08, 2.568564e-08, 2.572644e-08, 2.567299e-08, 2.576193e-08, 
    2.571064e-08, 2.575676e-08, 2.557928e-08, 2.558591e-08, 2.551154e-08,
  2.599855e-08, 2.601316e-08, 2.596094e-08, 2.601954e-08, 2.640611e-08, 
    2.593066e-08, 2.581816e-08, 2.579599e-08, 2.613664e-08, 2.604541e-08, 
    2.591674e-08, 2.592341e-08, 2.575067e-08, 2.586037e-08, 2.573325e-08,
  2.806648e-08, 2.803739e-08, 2.724952e-08, 2.748734e-08, 2.833593e-08, 
    2.750545e-08, 2.666963e-08, 2.642764e-08, 2.593319e-08, 2.600451e-08, 
    2.613628e-08, 2.648411e-08, 2.669605e-08, 2.717296e-08, 2.702639e-08,
  3.041054e-08, 2.992726e-08, 2.930744e-08, 2.981637e-08, 2.853506e-08, 
    2.623019e-08, 2.617142e-08, 2.603054e-08, 2.630688e-08, 2.709381e-08, 
    2.739882e-08, 2.769914e-08, 2.771179e-08, 2.813099e-08, 2.834476e-08,
  2.789711e-08, 2.793158e-08, 2.727986e-08, 2.66548e-08, 2.572529e-08, 
    2.401664e-08, 2.361642e-08, 2.332249e-08, 2.349745e-08, 2.358856e-08, 
    2.376726e-08, 2.423057e-08, 2.40728e-08, 2.410765e-08, 2.43643e-08,
  2.871518e-08, 2.88135e-08, 2.85752e-08, 2.741918e-08, 2.660551e-08, 
    2.570826e-08, 2.436389e-08, 2.323679e-08, 2.310539e-08, 2.319174e-08, 
    2.33589e-08, 2.360522e-08, 2.407736e-08, 2.419287e-08, 2.411874e-08,
  2.862804e-08, 2.949559e-08, 2.865935e-08, 2.886939e-08, 2.729194e-08, 
    2.563054e-08, 2.574868e-08, 2.454522e-08, 2.368803e-08, 2.338693e-08, 
    2.328021e-08, 2.313739e-08, 2.320213e-08, 2.330141e-08, 2.339426e-08,
  2.900901e-08, 2.883775e-08, 3.010154e-08, 2.82016e-08, 2.95553e-08, 
    2.767798e-08, 2.561171e-08, 2.533206e-08, 2.448561e-08, 2.390755e-08, 
    2.349572e-08, 2.31012e-08, 2.28499e-08, 2.278282e-08, 2.290081e-08,
  2.825178e-08, 2.802962e-08, 2.879165e-08, 2.897282e-08, 2.825388e-08, 
    2.902884e-08, 2.772508e-08, 2.625018e-08, 2.522772e-08, 2.487964e-08, 
    2.436276e-08, 2.395156e-08, 2.360802e-08, 2.341431e-08, 2.328221e-08,
  2.742907e-08, 2.83012e-08, 2.788669e-08, 2.888786e-08, 2.857786e-08, 
    2.815326e-08, 2.812802e-08, 2.711636e-08, 2.602449e-08, 2.51876e-08, 
    2.473375e-08, 2.429622e-08, 2.401728e-08, 2.384877e-08, 2.367316e-08,
  2.702384e-08, 2.733949e-08, 2.766873e-08, 2.785643e-08, 2.857615e-08, 
    2.817296e-08, 2.820444e-08, 2.78632e-08, 2.721635e-08, 2.661478e-08, 
    2.605046e-08, 2.560332e-08, 2.51291e-08, 2.487419e-08, 2.442452e-08,
  2.727686e-08, 2.70449e-08, 2.697174e-08, 2.722613e-08, 2.746247e-08, 
    2.75501e-08, 2.732263e-08, 2.71396e-08, 2.685097e-08, 2.672082e-08, 
    2.636249e-08, 2.612971e-08, 2.58337e-08, 2.571848e-08, 2.549465e-08,
  2.82814e-08, 2.816051e-08, 2.744716e-08, 2.713343e-08, 2.655278e-08, 
    2.701177e-08, 2.674724e-08, 2.670961e-08, 2.64741e-08, 2.649779e-08, 
    2.631992e-08, 2.637924e-08, 2.627498e-08, 2.603827e-08, 2.595629e-08,
  2.695048e-08, 2.724509e-08, 2.78985e-08, 2.878674e-08, 2.853145e-08, 
    2.782126e-08, 2.708712e-08, 2.686534e-08, 2.688739e-08, 2.674833e-08, 
    2.639982e-08, 2.649865e-08, 2.654847e-08, 2.668359e-08, 2.667993e-08,
  2.478506e-08, 2.525063e-08, 2.585217e-08, 2.643601e-08, 2.714635e-08, 
    2.732047e-08, 2.715584e-08, 2.669855e-08, 2.58624e-08, 2.494838e-08, 
    2.424074e-08, 2.393567e-08, 2.398759e-08, 2.420467e-08, 2.43256e-08,
  2.463018e-08, 2.530588e-08, 2.596286e-08, 2.628913e-08, 2.71369e-08, 
    2.755248e-08, 2.773838e-08, 2.701916e-08, 2.645615e-08, 2.5403e-08, 
    2.463624e-08, 2.388724e-08, 2.384362e-08, 2.39858e-08, 2.434208e-08,
  2.478989e-08, 2.537163e-08, 2.593869e-08, 2.591857e-08, 2.706932e-08, 
    2.73272e-08, 2.806058e-08, 2.786901e-08, 2.718416e-08, 2.652928e-08, 
    2.551116e-08, 2.455741e-08, 2.380624e-08, 2.361225e-08, 2.366731e-08,
  2.506679e-08, 2.549121e-08, 2.578438e-08, 2.617533e-08, 2.658055e-08, 
    2.77783e-08, 2.772332e-08, 2.826098e-08, 2.807545e-08, 2.75359e-08, 
    2.66097e-08, 2.549054e-08, 2.469608e-08, 2.379744e-08, 2.367063e-08,
  2.519475e-08, 2.538574e-08, 2.57301e-08, 2.630165e-08, 2.657805e-08, 
    2.663457e-08, 2.781504e-08, 2.816443e-08, 2.82617e-08, 2.881491e-08, 
    2.827952e-08, 2.716748e-08, 2.599815e-08, 2.485908e-08, 2.400505e-08,
  2.559095e-08, 2.560353e-08, 2.594977e-08, 2.607113e-08, 2.642692e-08, 
    2.631859e-08, 2.684725e-08, 2.802794e-08, 2.826983e-08, 2.845596e-08, 
    2.856662e-08, 2.811451e-08, 2.747416e-08, 2.64289e-08, 2.50999e-08,
  2.559471e-08, 2.562593e-08, 2.584865e-08, 2.578598e-08, 2.588413e-08, 
    2.622338e-08, 2.656857e-08, 2.714415e-08, 2.777043e-08, 2.832742e-08, 
    2.857351e-08, 2.856992e-08, 2.831429e-08, 2.780929e-08, 2.683037e-08,
  2.59405e-08, 2.560632e-08, 2.554125e-08, 2.558309e-08, 2.570618e-08, 
    2.59494e-08, 2.640797e-08, 2.691106e-08, 2.727507e-08, 2.785026e-08, 
    2.809838e-08, 2.846853e-08, 2.855734e-08, 2.865321e-08, 2.845495e-08,
  2.539082e-08, 2.494622e-08, 2.5122e-08, 2.525132e-08, 2.550668e-08, 
    2.575466e-08, 2.636728e-08, 2.663913e-08, 2.688114e-08, 2.723156e-08, 
    2.728507e-08, 2.744594e-08, 2.7477e-08, 2.757422e-08, 2.78181e-08,
  2.506161e-08, 2.468341e-08, 2.450997e-08, 2.468312e-08, 2.530759e-08, 
    2.607539e-08, 2.676383e-08, 2.719692e-08, 2.78249e-08, 2.80329e-08, 
    2.789515e-08, 2.746442e-08, 2.707356e-08, 2.685129e-08, 2.689949e-08,
  2.422515e-08, 2.361242e-08, 2.34856e-08, 2.337581e-08, 2.34195e-08, 
    2.341901e-08, 2.331157e-08, 2.36245e-08, 2.401935e-08, 2.467854e-08, 
    2.545999e-08, 2.579559e-08, 2.60762e-08, 2.604691e-08, 2.595883e-08,
  2.37493e-08, 2.342749e-08, 2.321199e-08, 2.319389e-08, 2.326048e-08, 
    2.319657e-08, 2.320864e-08, 2.349247e-08, 2.390575e-08, 2.446352e-08, 
    2.505266e-08, 2.575372e-08, 2.621784e-08, 2.637205e-08, 2.593744e-08,
  2.28862e-08, 2.295945e-08, 2.258572e-08, 2.284008e-08, 2.277982e-08, 
    2.3073e-08, 2.278618e-08, 2.363074e-08, 2.396881e-08, 2.441852e-08, 
    2.525187e-08, 2.605176e-08, 2.661237e-08, 2.654233e-08, 2.645176e-08,
  2.290971e-08, 2.271441e-08, 2.261092e-08, 2.268091e-08, 2.283502e-08, 
    2.349653e-08, 2.340704e-08, 2.396068e-08, 2.437917e-08, 2.495301e-08, 
    2.557268e-08, 2.625446e-08, 2.666785e-08, 2.658164e-08, 2.660404e-08,
  2.351789e-08, 2.312296e-08, 2.28181e-08, 2.30063e-08, 2.338354e-08, 
    2.379026e-08, 2.434593e-08, 2.388928e-08, 2.42479e-08, 2.49325e-08, 
    2.558555e-08, 2.615273e-08, 2.650618e-08, 2.668667e-08, 2.650154e-08,
  2.431014e-08, 2.410778e-08, 2.404e-08, 2.413551e-08, 2.425847e-08, 
    2.437499e-08, 2.436158e-08, 2.482113e-08, 2.528625e-08, 2.545679e-08, 
    2.562697e-08, 2.606563e-08, 2.602418e-08, 2.629094e-08, 2.641836e-08,
  2.442174e-08, 2.444851e-08, 2.455354e-08, 2.452871e-08, 2.443348e-08, 
    2.433057e-08, 2.463883e-08, 2.476243e-08, 2.523382e-08, 2.524794e-08, 
    2.563914e-08, 2.582544e-08, 2.579001e-08, 2.584514e-08, 2.622514e-08,
  2.608121e-08, 2.608999e-08, 2.556089e-08, 2.533907e-08, 2.52769e-08, 
    2.537767e-08, 2.532284e-08, 2.554136e-08, 2.560975e-08, 2.571134e-08, 
    2.585751e-08, 2.577643e-08, 2.585181e-08, 2.599442e-08, 2.632515e-08,
  2.581472e-08, 2.58227e-08, 2.589514e-08, 2.601087e-08, 2.616281e-08, 
    2.625412e-08, 2.601526e-08, 2.592278e-08, 2.580001e-08, 2.567177e-08, 
    2.582855e-08, 2.588685e-08, 2.59969e-08, 2.629922e-08, 2.688564e-08,
  2.44728e-08, 2.501873e-08, 2.582109e-08, 2.606906e-08, 2.640652e-08, 
    2.585737e-08, 2.577032e-08, 2.553378e-08, 2.564473e-08, 2.563804e-08, 
    2.583077e-08, 2.608956e-08, 2.648453e-08, 2.676986e-08, 2.707351e-08,
  2.538096e-08, 2.533565e-08, 2.504528e-08, 2.520436e-08, 2.516251e-08, 
    2.535807e-08, 2.523172e-08, 2.4876e-08, 2.451873e-08, 2.39563e-08, 
    2.365142e-08, 2.328671e-08, 2.317507e-08, 2.296689e-08, 2.311713e-08,
  2.551601e-08, 2.518654e-08, 2.51151e-08, 2.489977e-08, 2.508174e-08, 
    2.488887e-08, 2.519872e-08, 2.483463e-08, 2.446477e-08, 2.405467e-08, 
    2.368996e-08, 2.325797e-08, 2.331097e-08, 2.309704e-08, 2.305971e-08,
  2.556762e-08, 2.525246e-08, 2.527639e-08, 2.487611e-08, 2.50979e-08, 
    2.521566e-08, 2.509617e-08, 2.510955e-08, 2.450166e-08, 2.406185e-08, 
    2.364666e-08, 2.33491e-08, 2.348803e-08, 2.338483e-08, 2.368587e-08,
  2.554742e-08, 2.552422e-08, 2.526468e-08, 2.524182e-08, 2.457556e-08, 
    2.468091e-08, 2.475376e-08, 2.47869e-08, 2.441817e-08, 2.3976e-08, 
    2.36961e-08, 2.338519e-08, 2.366546e-08, 2.347625e-08, 2.399391e-08,
  2.58071e-08, 2.563603e-08, 2.54032e-08, 2.53266e-08, 2.487345e-08, 
    2.446379e-08, 2.417599e-08, 2.398713e-08, 2.439718e-08, 2.393904e-08, 
    2.401214e-08, 2.370157e-08, 2.375416e-08, 2.384056e-08, 2.41094e-08,
  2.577056e-08, 2.547598e-08, 2.543241e-08, 2.528515e-08, 2.533165e-08, 
    2.466361e-08, 2.468017e-08, 2.429441e-08, 2.430964e-08, 2.375472e-08, 
    2.328646e-08, 2.319265e-08, 2.346043e-08, 2.387132e-08, 2.432757e-08,
  2.555087e-08, 2.513387e-08, 2.52202e-08, 2.50683e-08, 2.532149e-08, 
    2.499023e-08, 2.476234e-08, 2.477358e-08, 2.461631e-08, 2.415818e-08, 
    2.391178e-08, 2.375525e-08, 2.408007e-08, 2.461524e-08, 2.472224e-08,
  2.526757e-08, 2.515074e-08, 2.516298e-08, 2.505354e-08, 2.534703e-08, 
    2.522476e-08, 2.511752e-08, 2.478166e-08, 2.443535e-08, 2.406042e-08, 
    2.411912e-08, 2.440045e-08, 2.492978e-08, 2.515132e-08, 2.513423e-08,
  2.498103e-08, 2.48643e-08, 2.497807e-08, 2.51486e-08, 2.540741e-08, 
    2.532011e-08, 2.525345e-08, 2.49662e-08, 2.473009e-08, 2.478052e-08, 
    2.485643e-08, 2.521979e-08, 2.532575e-08, 2.518358e-08, 2.556521e-08,
  2.529179e-08, 2.496271e-08, 2.473539e-08, 2.481257e-08, 2.495872e-08, 
    2.533687e-08, 2.516791e-08, 2.55306e-08, 2.516979e-08, 2.514484e-08, 
    2.520073e-08, 2.528764e-08, 2.526788e-08, 2.551545e-08, 2.578087e-08,
  2.704477e-08, 2.695066e-08, 2.718024e-08, 2.735169e-08, 2.716315e-08, 
    2.706183e-08, 2.671315e-08, 2.663462e-08, 2.637388e-08, 2.618502e-08, 
    2.589062e-08, 2.553458e-08, 2.553762e-08, 2.538848e-08, 2.52243e-08,
  2.707216e-08, 2.696212e-08, 2.744568e-08, 2.738147e-08, 2.735583e-08, 
    2.687611e-08, 2.664218e-08, 2.650586e-08, 2.616495e-08, 2.620731e-08, 
    2.572757e-08, 2.529151e-08, 2.520478e-08, 2.502626e-08, 2.508146e-08,
  2.711557e-08, 2.712755e-08, 2.743297e-08, 2.734887e-08, 2.719413e-08, 
    2.670914e-08, 2.663814e-08, 2.661152e-08, 2.626887e-08, 2.606219e-08, 
    2.588759e-08, 2.5383e-08, 2.527566e-08, 2.530273e-08, 2.524979e-08,
  2.706109e-08, 2.704429e-08, 2.757826e-08, 2.727729e-08, 2.693619e-08, 
    2.704052e-08, 2.642411e-08, 2.638549e-08, 2.613643e-08, 2.565684e-08, 
    2.539335e-08, 2.503113e-08, 2.489245e-08, 2.481507e-08, 2.477077e-08,
  2.706662e-08, 2.731349e-08, 2.753469e-08, 2.691436e-08, 2.668756e-08, 
    2.661869e-08, 2.667972e-08, 2.605538e-08, 2.64509e-08, 2.671799e-08, 
    2.629162e-08, 2.594117e-08, 2.547943e-08, 2.550294e-08, 2.51533e-08,
  2.715022e-08, 2.707142e-08, 2.68544e-08, 2.641307e-08, 2.638791e-08, 
    2.616856e-08, 2.619244e-08, 2.609152e-08, 2.480025e-08, 2.502743e-08, 
    2.512722e-08, 2.508824e-08, 2.506927e-08, 2.493219e-08, 2.465963e-08,
  2.691326e-08, 2.659572e-08, 2.638258e-08, 2.628786e-08, 2.605235e-08, 
    2.587587e-08, 2.58434e-08, 2.543972e-08, 2.529409e-08, 2.462379e-08, 
    2.480727e-08, 2.468455e-08, 2.491763e-08, 2.478328e-08, 2.47495e-08,
  2.676621e-08, 2.630233e-08, 2.62953e-08, 2.619325e-08, 2.604057e-08, 
    2.570583e-08, 2.553162e-08, 2.533164e-08, 2.512678e-08, 2.513558e-08, 
    2.491783e-08, 2.494633e-08, 2.474863e-08, 2.489142e-08, 2.469641e-08,
  2.633734e-08, 2.589431e-08, 2.6262e-08, 2.634144e-08, 2.617714e-08, 
    2.569096e-08, 2.52609e-08, 2.521962e-08, 2.488849e-08, 2.528501e-08, 
    2.505938e-08, 2.522424e-08, 2.518541e-08, 2.501684e-08, 2.480398e-08,
  2.54595e-08, 2.582664e-08, 2.639095e-08, 2.651242e-08, 2.640944e-08, 
    2.590085e-08, 2.565915e-08, 2.528812e-08, 2.474347e-08, 2.50414e-08, 
    2.48183e-08, 2.507816e-08, 2.507185e-08, 2.502327e-08, 2.487089e-08,
  2.527709e-08, 2.490828e-08, 2.525036e-08, 2.486876e-08, 2.541882e-08, 
    2.592297e-08, 2.630342e-08, 2.646893e-08, 2.667449e-08, 2.685427e-08, 
    2.688518e-08, 2.738194e-08, 2.692152e-08, 2.693366e-08, 2.650002e-08,
  2.492236e-08, 2.473095e-08, 2.48243e-08, 2.458437e-08, 2.603454e-08, 
    2.595105e-08, 2.607832e-08, 2.613383e-08, 2.64408e-08, 2.667054e-08, 
    2.691281e-08, 2.682249e-08, 2.709096e-08, 2.651306e-08, 2.601948e-08,
  2.438175e-08, 2.441877e-08, 2.424141e-08, 2.543803e-08, 2.617696e-08, 
    2.579524e-08, 2.553354e-08, 2.592697e-08, 2.615783e-08, 2.608236e-08, 
    2.690903e-08, 2.700425e-08, 2.72226e-08, 2.665501e-08, 2.649029e-08,
  2.43721e-08, 2.431805e-08, 2.508372e-08, 2.596988e-08, 2.551294e-08, 
    2.563661e-08, 2.573714e-08, 2.572753e-08, 2.606043e-08, 2.619762e-08, 
    2.63765e-08, 2.675668e-08, 2.666965e-08, 2.610727e-08, 2.610772e-08,
  2.423933e-08, 2.457924e-08, 2.531813e-08, 2.527104e-08, 2.521435e-08, 
    2.51089e-08, 2.589553e-08, 2.520039e-08, 2.575501e-08, 2.664939e-08, 
    2.714368e-08, 2.737958e-08, 2.743269e-08, 2.695396e-08, 2.642394e-08,
  2.445236e-08, 2.512799e-08, 2.519095e-08, 2.523168e-08, 2.496104e-08, 
    2.530899e-08, 2.516499e-08, 2.588814e-08, 2.535809e-08, 2.553639e-08, 
    2.614263e-08, 2.6731e-08, 2.689923e-08, 2.670904e-08, 2.640887e-08,
  2.524212e-08, 2.540992e-08, 2.517248e-08, 2.467401e-08, 2.471095e-08, 
    2.46763e-08, 2.497889e-08, 2.513915e-08, 2.528887e-08, 2.583041e-08, 
    2.592859e-08, 2.610895e-08, 2.608773e-08, 2.584921e-08, 2.578349e-08,
  2.543042e-08, 2.529387e-08, 2.459646e-08, 2.432144e-08, 2.429881e-08, 
    2.45489e-08, 2.495107e-08, 2.512662e-08, 2.569384e-08, 2.598542e-08, 
    2.60486e-08, 2.596537e-08, 2.562186e-08, 2.551285e-08, 2.523303e-08,
  2.528891e-08, 2.481146e-08, 2.446148e-08, 2.438614e-08, 2.465002e-08, 
    2.494504e-08, 2.531652e-08, 2.548409e-08, 2.590392e-08, 2.605283e-08, 
    2.600183e-08, 2.602405e-08, 2.566518e-08, 2.546127e-08, 2.519238e-08,
  2.50619e-08, 2.493625e-08, 2.52764e-08, 2.523199e-08, 2.522154e-08, 
    2.522283e-08, 2.525877e-08, 2.557793e-08, 2.576828e-08, 2.602217e-08, 
    2.58233e-08, 2.565688e-08, 2.549631e-08, 2.517861e-08, 2.501753e-08,
  2.48489e-08, 2.485785e-08, 2.483749e-08, 2.474377e-08, 2.45639e-08, 
    2.4523e-08, 2.451886e-08, 2.450987e-08, 2.454599e-08, 2.46845e-08, 
    2.471521e-08, 2.492123e-08, 2.481199e-08, 2.491176e-08, 2.532773e-08,
  2.478765e-08, 2.470103e-08, 2.481355e-08, 2.457352e-08, 2.485297e-08, 
    2.473096e-08, 2.486447e-08, 2.491313e-08, 2.508439e-08, 2.508354e-08, 
    2.508769e-08, 2.491349e-08, 2.520859e-08, 2.527515e-08, 2.537699e-08,
  2.503309e-08, 2.516566e-08, 2.523136e-08, 2.506003e-08, 2.54388e-08, 
    2.526166e-08, 2.504391e-08, 2.494192e-08, 2.505583e-08, 2.491437e-08, 
    2.488526e-08, 2.488744e-08, 2.505164e-08, 2.516985e-08, 2.536347e-08,
  2.556438e-08, 2.553052e-08, 2.544374e-08, 2.551616e-08, 2.525856e-08, 
    2.527504e-08, 2.49875e-08, 2.495415e-08, 2.492897e-08, 2.489086e-08, 
    2.484574e-08, 2.47749e-08, 2.52537e-08, 2.47183e-08, 2.560869e-08,
  2.579106e-08, 2.581133e-08, 2.576285e-08, 2.574381e-08, 2.559269e-08, 
    2.554991e-08, 2.564063e-08, 2.522453e-08, 2.493266e-08, 2.521847e-08, 
    2.493247e-08, 2.471629e-08, 2.484959e-08, 2.495336e-08, 2.488382e-08,
  2.626816e-08, 2.615265e-08, 2.624529e-08, 2.635337e-08, 2.636373e-08, 
    2.640822e-08, 2.617002e-08, 2.634626e-08, 2.605891e-08, 2.554719e-08, 
    2.514138e-08, 2.492816e-08, 2.48034e-08, 2.520257e-08, 2.501633e-08,
  2.636894e-08, 2.663148e-08, 2.701684e-08, 2.720058e-08, 2.727514e-08, 
    2.708804e-08, 2.687438e-08, 2.648696e-08, 2.60422e-08, 2.553737e-08, 
    2.515348e-08, 2.493078e-08, 2.493907e-08, 2.530474e-08, 2.522245e-08,
  2.696206e-08, 2.726732e-08, 2.755399e-08, 2.763912e-08, 2.75897e-08, 
    2.734675e-08, 2.719881e-08, 2.663662e-08, 2.615536e-08, 2.545658e-08, 
    2.506229e-08, 2.47882e-08, 2.48161e-08, 2.520923e-08, 2.530568e-08,
  2.730254e-08, 2.756875e-08, 2.799403e-08, 2.805607e-08, 2.808371e-08, 
    2.795504e-08, 2.784827e-08, 2.723808e-08, 2.665454e-08, 2.561756e-08, 
    2.486567e-08, 2.466568e-08, 2.462439e-08, 2.498653e-08, 2.531657e-08,
  2.751956e-08, 2.791506e-08, 2.828367e-08, 2.826738e-08, 2.816852e-08, 
    2.795295e-08, 2.793965e-08, 2.761584e-08, 2.657923e-08, 2.549907e-08, 
    2.476215e-08, 2.464827e-08, 2.456091e-08, 2.496092e-08, 2.534292e-08,
  2.719843e-08, 2.736714e-08, 2.75358e-08, 2.76341e-08, 2.748546e-08, 
    2.76308e-08, 2.755305e-08, 2.735171e-08, 2.716721e-08, 2.687825e-08, 
    2.643951e-08, 2.621894e-08, 2.586246e-08, 2.579213e-08, 2.54586e-08,
  2.726245e-08, 2.720397e-08, 2.73655e-08, 2.730652e-08, 2.768495e-08, 
    2.776015e-08, 2.76654e-08, 2.750333e-08, 2.733158e-08, 2.687313e-08, 
    2.643977e-08, 2.599502e-08, 2.587594e-08, 2.554284e-08, 2.534718e-08,
  2.677485e-08, 2.676756e-08, 2.694449e-08, 2.735985e-08, 2.781825e-08, 
    2.788004e-08, 2.788923e-08, 2.794546e-08, 2.772451e-08, 2.718936e-08, 
    2.668795e-08, 2.619655e-08, 2.57741e-08, 2.557413e-08, 2.546216e-08,
  2.672208e-08, 2.664941e-08, 2.686069e-08, 2.724415e-08, 2.780131e-08, 
    2.835158e-08, 2.820751e-08, 2.830969e-08, 2.776755e-08, 2.721293e-08, 
    2.676917e-08, 2.617552e-08, 2.574724e-08, 2.551554e-08, 2.567923e-08,
  2.662095e-08, 2.642066e-08, 2.654361e-08, 2.688335e-08, 2.750378e-08, 
    2.804501e-08, 2.855565e-08, 2.814801e-08, 2.733182e-08, 2.710863e-08, 
    2.673396e-08, 2.600145e-08, 2.576076e-08, 2.535314e-08, 2.547965e-08,
  2.656333e-08, 2.649236e-08, 2.641578e-08, 2.654355e-08, 2.702707e-08, 
    2.781197e-08, 2.815198e-08, 2.850011e-08, 2.805108e-08, 2.70866e-08, 
    2.67851e-08, 2.613895e-08, 2.586559e-08, 2.551844e-08, 2.545408e-08,
  2.657912e-08, 2.660058e-08, 2.633032e-08, 2.622909e-08, 2.645289e-08, 
    2.705642e-08, 2.783229e-08, 2.797733e-08, 2.76271e-08, 2.706151e-08, 
    2.64352e-08, 2.587257e-08, 2.566649e-08, 2.571661e-08, 2.549173e-08,
  2.657413e-08, 2.679175e-08, 2.663616e-08, 2.611503e-08, 2.583782e-08, 
    2.624323e-08, 2.715115e-08, 2.755466e-08, 2.747032e-08, 2.689891e-08, 
    2.642658e-08, 2.624973e-08, 2.598119e-08, 2.583983e-08, 2.512591e-08,
  2.647766e-08, 2.658924e-08, 2.671143e-08, 2.641096e-08, 2.584136e-08, 
    2.563926e-08, 2.625881e-08, 2.690982e-08, 2.711628e-08, 2.703159e-08, 
    2.647048e-08, 2.601914e-08, 2.564594e-08, 2.546174e-08, 2.46598e-08,
  2.640181e-08, 2.653596e-08, 2.665224e-08, 2.666126e-08, 2.597011e-08, 
    2.538427e-08, 2.548175e-08, 2.605288e-08, 2.632543e-08, 2.616852e-08, 
    2.61195e-08, 2.562841e-08, 2.526004e-08, 2.480963e-08, 2.469663e-08,
  2.503526e-08, 2.496801e-08, 2.560697e-08, 2.590942e-08, 2.633259e-08, 
    2.667133e-08, 2.694111e-08, 2.722131e-08, 2.778897e-08, 2.823877e-08, 
    2.829423e-08, 2.821602e-08, 2.815786e-08, 2.79285e-08, 2.793966e-08,
  2.566158e-08, 2.508189e-08, 2.557759e-08, 2.598157e-08, 2.615464e-08, 
    2.6264e-08, 2.662801e-08, 2.691601e-08, 2.738853e-08, 2.766467e-08, 
    2.78589e-08, 2.787585e-08, 2.797151e-08, 2.785838e-08, 2.759738e-08,
  2.613067e-08, 2.526872e-08, 2.526203e-08, 2.565739e-08, 2.600967e-08, 
    2.587119e-08, 2.59375e-08, 2.619423e-08, 2.650786e-08, 2.724894e-08, 
    2.744476e-08, 2.752599e-08, 2.767628e-08, 2.749566e-08, 2.727878e-08,
  2.661215e-08, 2.595828e-08, 2.543708e-08, 2.532634e-08, 2.611046e-08, 
    2.598333e-08, 2.572698e-08, 2.564048e-08, 2.581036e-08, 2.653851e-08, 
    2.699363e-08, 2.724732e-08, 2.730257e-08, 2.724273e-08, 2.710248e-08,
  2.608309e-08, 2.632302e-08, 2.586603e-08, 2.547042e-08, 2.532307e-08, 
    2.56508e-08, 2.578862e-08, 2.550696e-08, 2.531586e-08, 2.573293e-08, 
    2.601307e-08, 2.666522e-08, 2.683966e-08, 2.702847e-08, 2.705442e-08,
  2.584334e-08, 2.627947e-08, 2.612226e-08, 2.597295e-08, 2.584156e-08, 
    2.531424e-08, 2.533989e-08, 2.580544e-08, 2.561702e-08, 2.503911e-08, 
    2.545686e-08, 2.605208e-08, 2.637962e-08, 2.666945e-08, 2.700326e-08,
  2.550046e-08, 2.597781e-08, 2.597391e-08, 2.574164e-08, 2.615935e-08, 
    2.594859e-08, 2.512192e-08, 2.481691e-08, 2.518244e-08, 2.521165e-08, 
    2.477925e-08, 2.534869e-08, 2.576143e-08, 2.608559e-08, 2.60707e-08,
  2.528417e-08, 2.584541e-08, 2.583674e-08, 2.55462e-08, 2.595021e-08, 
    2.631242e-08, 2.606097e-08, 2.523426e-08, 2.506331e-08, 2.550629e-08, 
    2.53987e-08, 2.479142e-08, 2.478605e-08, 2.462023e-08, 2.419427e-08,
  2.51186e-08, 2.56112e-08, 2.584925e-08, 2.52193e-08, 2.545043e-08, 
    2.627139e-08, 2.620124e-08, 2.599455e-08, 2.488895e-08, 2.492412e-08, 
    2.547932e-08, 2.518263e-08, 2.500822e-08, 2.451038e-08, 2.438973e-08,
  2.488967e-08, 2.552512e-08, 2.563498e-08, 2.540185e-08, 2.496296e-08, 
    2.586872e-08, 2.63567e-08, 2.674968e-08, 2.599794e-08, 2.494036e-08, 
    2.510106e-08, 2.526725e-08, 2.539274e-08, 2.542709e-08, 2.573228e-08,
  2.440603e-08, 2.459385e-08, 2.543005e-08, 2.665101e-08, 2.608344e-08, 
    2.480273e-08, 2.564551e-08, 2.721971e-08, 2.761607e-08, 2.760092e-08, 
    2.800561e-08, 2.828966e-08, 2.815309e-08, 2.816203e-08, 2.82195e-08,
  2.450925e-08, 2.461674e-08, 2.505253e-08, 2.656397e-08, 2.657047e-08, 
    2.492446e-08, 2.518241e-08, 2.689288e-08, 2.752457e-08, 2.739213e-08, 
    2.773787e-08, 2.806748e-08, 2.806902e-08, 2.805145e-08, 2.804722e-08,
  2.444901e-08, 2.473044e-08, 2.477992e-08, 2.60292e-08, 2.689822e-08, 
    2.531377e-08, 2.497871e-08, 2.655065e-08, 2.74403e-08, 2.7361e-08, 
    2.733918e-08, 2.772936e-08, 2.783658e-08, 2.769264e-08, 2.741039e-08,
  2.423177e-08, 2.480634e-08, 2.477582e-08, 2.552216e-08, 2.694561e-08, 
    2.596902e-08, 2.485936e-08, 2.569906e-08, 2.722618e-08, 2.733523e-08, 
    2.71922e-08, 2.712246e-08, 2.716557e-08, 2.71073e-08, 2.705385e-08,
  2.410045e-08, 2.467549e-08, 2.491646e-08, 2.540195e-08, 2.639318e-08, 
    2.653819e-08, 2.56603e-08, 2.505346e-08, 2.653337e-08, 2.766959e-08, 
    2.743886e-08, 2.712041e-08, 2.696776e-08, 2.700002e-08, 2.705302e-08,
  2.404708e-08, 2.445791e-08, 2.480679e-08, 2.525632e-08, 2.629898e-08, 
    2.671237e-08, 2.559314e-08, 2.548543e-08, 2.593285e-08, 2.670135e-08, 
    2.786279e-08, 2.756829e-08, 2.725661e-08, 2.706724e-08, 2.706941e-08,
  2.387878e-08, 2.43752e-08, 2.485445e-08, 2.507947e-08, 2.59012e-08, 
    2.700878e-08, 2.620533e-08, 2.461136e-08, 2.478252e-08, 2.558156e-08, 
    2.629118e-08, 2.770195e-08, 2.741861e-08, 2.738733e-08, 2.698412e-08,
  2.376583e-08, 2.412882e-08, 2.472972e-08, 2.506579e-08, 2.566764e-08, 
    2.678281e-08, 2.705632e-08, 2.567391e-08, 2.466005e-08, 2.504441e-08, 
    2.502403e-08, 2.563091e-08, 2.619126e-08, 2.610239e-08, 2.591103e-08,
  2.370376e-08, 2.397939e-08, 2.452647e-08, 2.494501e-08, 2.544309e-08, 
    2.646144e-08, 2.717393e-08, 2.65625e-08, 2.535654e-08, 2.524072e-08, 
    2.510713e-08, 2.493456e-08, 2.511719e-08, 2.513131e-08, 2.528566e-08,
  2.369802e-08, 2.386404e-08, 2.43795e-08, 2.484023e-08, 2.526994e-08, 
    2.615752e-08, 2.754141e-08, 2.749021e-08, 2.616454e-08, 2.562889e-08, 
    2.546841e-08, 2.55018e-08, 2.528814e-08, 2.524312e-08, 2.532811e-08,
  2.584307e-08, 2.577101e-08, 2.601495e-08, 2.589129e-08, 2.559724e-08, 
    2.594493e-08, 2.677113e-08, 2.717948e-08, 2.760099e-08, 2.779243e-08, 
    2.808585e-08, 2.81398e-08, 2.819577e-08, 2.819202e-08, 2.805192e-08,
  2.594663e-08, 2.594714e-08, 2.591915e-08, 2.569935e-08, 2.578036e-08, 
    2.57971e-08, 2.677036e-08, 2.721946e-08, 2.739266e-08, 2.778779e-08, 
    2.805945e-08, 2.820491e-08, 2.819748e-08, 2.851972e-08, 2.834402e-08,
  2.623919e-08, 2.596845e-08, 2.590074e-08, 2.570485e-08, 2.576312e-08, 
    2.586362e-08, 2.64324e-08, 2.701586e-08, 2.735618e-08, 2.752969e-08, 
    2.812647e-08, 2.806074e-08, 2.823654e-08, 2.852102e-08, 2.850569e-08,
  2.64745e-08, 2.620258e-08, 2.602339e-08, 2.548483e-08, 2.585615e-08, 
    2.650432e-08, 2.636674e-08, 2.62337e-08, 2.690539e-08, 2.753077e-08, 
    2.799284e-08, 2.829778e-08, 2.843451e-08, 2.866927e-08, 2.866362e-08,
  2.674125e-08, 2.631212e-08, 2.634132e-08, 2.57136e-08, 2.512444e-08, 
    2.589729e-08, 2.710817e-08, 2.601568e-08, 2.666681e-08, 2.716994e-08, 
    2.770101e-08, 2.837493e-08, 2.847827e-08, 2.867893e-08, 2.857884e-08,
  2.704842e-08, 2.66132e-08, 2.617869e-08, 2.607399e-08, 2.559283e-08, 
    2.510554e-08, 2.641109e-08, 2.782828e-08, 2.729882e-08, 2.685128e-08, 
    2.741543e-08, 2.77981e-08, 2.810893e-08, 2.83513e-08, 2.817864e-08,
  2.721688e-08, 2.732628e-08, 2.676778e-08, 2.614576e-08, 2.572732e-08, 
    2.537021e-08, 2.529008e-08, 2.555851e-08, 2.650852e-08, 2.676929e-08, 
    2.697191e-08, 2.764892e-08, 2.777345e-08, 2.803429e-08, 2.797224e-08,
  2.713433e-08, 2.752202e-08, 2.727706e-08, 2.681303e-08, 2.598271e-08, 
    2.564269e-08, 2.567561e-08, 2.604633e-08, 2.621651e-08, 2.655576e-08, 
    2.643944e-08, 2.692053e-08, 2.743803e-08, 2.77108e-08, 2.756818e-08,
  2.70059e-08, 2.757269e-08, 2.787026e-08, 2.746433e-08, 2.672124e-08, 
    2.599953e-08, 2.542824e-08, 2.551552e-08, 2.60203e-08, 2.661342e-08, 
    2.660344e-08, 2.627342e-08, 2.66324e-08, 2.699698e-08, 2.703289e-08,
  2.644861e-08, 2.670068e-08, 2.75854e-08, 2.782009e-08, 2.714715e-08, 
    2.671297e-08, 2.61321e-08, 2.564754e-08, 2.543194e-08, 2.58083e-08, 
    2.665289e-08, 2.677489e-08, 2.637735e-08, 2.65846e-08, 2.683192e-08,
  2.591421e-08, 2.523725e-08, 2.507884e-08, 2.548425e-08, 2.60727e-08, 
    2.648551e-08, 2.637611e-08, 2.679902e-08, 2.749545e-08, 2.834117e-08, 
    2.820237e-08, 2.83323e-08, 2.771136e-08, 2.770571e-08, 2.709882e-08,
  2.590822e-08, 2.538254e-08, 2.511705e-08, 2.558974e-08, 2.59836e-08, 
    2.596627e-08, 2.643832e-08, 2.662672e-08, 2.736171e-08, 2.81582e-08, 
    2.857493e-08, 2.851562e-08, 2.812389e-08, 2.793265e-08, 2.723223e-08,
  2.584304e-08, 2.521426e-08, 2.494529e-08, 2.511282e-08, 2.560084e-08, 
    2.588884e-08, 2.576871e-08, 2.647726e-08, 2.755402e-08, 2.868632e-08, 
    2.909031e-08, 2.856688e-08, 2.810719e-08, 2.802557e-08, 2.74023e-08,
  2.585894e-08, 2.529537e-08, 2.502018e-08, 2.51745e-08, 2.562201e-08, 
    2.625141e-08, 2.59242e-08, 2.567644e-08, 2.649389e-08, 2.806368e-08, 
    2.897052e-08, 2.892504e-08, 2.852409e-08, 2.818144e-08, 2.775399e-08,
  2.562742e-08, 2.508763e-08, 2.493435e-08, 2.473183e-08, 2.490021e-08, 
    2.532636e-08, 2.609342e-08, 2.559053e-08, 2.621289e-08, 2.738441e-08, 
    2.866592e-08, 2.898109e-08, 2.890933e-08, 2.834006e-08, 2.802186e-08,
  2.54492e-08, 2.503758e-08, 2.476103e-08, 2.48098e-08, 2.493345e-08, 
    2.501305e-08, 2.534279e-08, 2.650453e-08, 2.651655e-08, 2.690411e-08, 
    2.812589e-08, 2.89483e-08, 2.90907e-08, 2.871363e-08, 2.804298e-08,
  2.520169e-08, 2.492044e-08, 2.448936e-08, 2.419458e-08, 2.450509e-08, 
    2.474292e-08, 2.480739e-08, 2.490606e-08, 2.535559e-08, 2.646748e-08, 
    2.730005e-08, 2.848207e-08, 2.848392e-08, 2.86778e-08, 2.83334e-08,
  2.4882e-08, 2.472131e-08, 2.461443e-08, 2.427062e-08, 2.426365e-08, 
    2.439261e-08, 2.463519e-08, 2.494872e-08, 2.512352e-08, 2.569585e-08, 
    2.657419e-08, 2.791404e-08, 2.836789e-08, 2.84222e-08, 2.800572e-08,
  2.491412e-08, 2.473109e-08, 2.464092e-08, 2.434773e-08, 2.436771e-08, 
    2.412875e-08, 2.394255e-08, 2.412537e-08, 2.442715e-08, 2.525896e-08, 
    2.613772e-08, 2.682356e-08, 2.811641e-08, 2.800493e-08, 2.829429e-08,
  2.499429e-08, 2.480732e-08, 2.49181e-08, 2.460553e-08, 2.448835e-08, 
    2.425324e-08, 2.398498e-08, 2.390834e-08, 2.391137e-08, 2.446643e-08, 
    2.567289e-08, 2.660931e-08, 2.680609e-08, 2.855876e-08, 2.766342e-08,
  2.499405e-08, 2.471767e-08, 2.447109e-08, 2.425298e-08, 2.409358e-08, 
    2.393029e-08, 2.398157e-08, 2.429408e-08, 2.453665e-08, 2.504512e-08, 
    2.530204e-08, 2.592599e-08, 2.624487e-08, 2.650783e-08, 2.687827e-08,
  2.493391e-08, 2.478578e-08, 2.463928e-08, 2.432229e-08, 2.441188e-08, 
    2.415686e-08, 2.453086e-08, 2.481355e-08, 2.493763e-08, 2.495358e-08, 
    2.537549e-08, 2.591938e-08, 2.668744e-08, 2.697077e-08, 2.704532e-08,
  2.504056e-08, 2.506763e-08, 2.504467e-08, 2.468286e-08, 2.491109e-08, 
    2.515102e-08, 2.517832e-08, 2.499586e-08, 2.478189e-08, 2.489276e-08, 
    2.524286e-08, 2.623202e-08, 2.664422e-08, 2.747014e-08, 2.758547e-08,
  2.54595e-08, 2.559439e-08, 2.525803e-08, 2.516235e-08, 2.527138e-08, 
    2.612711e-08, 2.531515e-08, 2.461997e-08, 2.453226e-08, 2.467447e-08, 
    2.52067e-08, 2.615549e-08, 2.687882e-08, 2.754217e-08, 2.818764e-08,
  2.578963e-08, 2.56897e-08, 2.548075e-08, 2.563358e-08, 2.583836e-08, 
    2.548081e-08, 2.53972e-08, 2.481361e-08, 2.415553e-08, 2.441136e-08, 
    2.505737e-08, 2.616466e-08, 2.725326e-08, 2.786046e-08, 2.829781e-08,
  2.602177e-08, 2.574458e-08, 2.572204e-08, 2.592448e-08, 2.584172e-08, 
    2.574779e-08, 2.51453e-08, 2.480211e-08, 2.45029e-08, 2.419496e-08, 
    2.50002e-08, 2.644162e-08, 2.755475e-08, 2.842123e-08, 2.835886e-08,
  2.606516e-08, 2.589984e-08, 2.600081e-08, 2.61063e-08, 2.602499e-08, 
    2.562496e-08, 2.513725e-08, 2.473127e-08, 2.421681e-08, 2.388614e-08, 
    2.485523e-08, 2.631515e-08, 2.753515e-08, 2.838753e-08, 2.837607e-08,
  2.628523e-08, 2.607937e-08, 2.616826e-08, 2.622052e-08, 2.596237e-08, 
    2.581693e-08, 2.543233e-08, 2.494074e-08, 2.428252e-08, 2.383677e-08, 
    2.475073e-08, 2.660617e-08, 2.785752e-08, 2.893762e-08, 2.844223e-08,
  2.611845e-08, 2.602377e-08, 2.615601e-08, 2.623313e-08, 2.614016e-08, 
    2.611393e-08, 2.587741e-08, 2.526595e-08, 2.447761e-08, 2.425112e-08, 
    2.442601e-08, 2.592827e-08, 2.742263e-08, 2.840636e-08, 2.851689e-08,
  2.612668e-08, 2.603464e-08, 2.62952e-08, 2.641043e-08, 2.632909e-08, 
    2.632953e-08, 2.641397e-08, 2.558897e-08, 2.453292e-08, 2.451749e-08, 
    2.418639e-08, 2.534216e-08, 2.766799e-08, 2.891895e-08, 2.849702e-08,
  2.532907e-08, 2.533568e-08, 2.54093e-08, 2.542397e-08, 2.553979e-08, 
    2.554333e-08, 2.558388e-08, 2.552947e-08, 2.555073e-08, 2.54927e-08, 
    2.551792e-08, 2.554588e-08, 2.551113e-08, 2.536426e-08, 2.516527e-08,
  2.607799e-08, 2.60938e-08, 2.617496e-08, 2.620833e-08, 2.633463e-08, 
    2.642618e-08, 2.643477e-08, 2.645891e-08, 2.650208e-08, 2.654673e-08, 
    2.672279e-08, 2.64794e-08, 2.66586e-08, 2.625509e-08, 2.58973e-08,
  2.627901e-08, 2.612183e-08, 2.636706e-08, 2.613339e-08, 2.662104e-08, 
    2.639835e-08, 2.631685e-08, 2.639765e-08, 2.643459e-08, 2.653842e-08, 
    2.646069e-08, 2.63594e-08, 2.62594e-08, 2.599713e-08, 2.598531e-08,
  2.584533e-08, 2.606567e-08, 2.589584e-08, 2.601564e-08, 2.581668e-08, 
    2.631434e-08, 2.598111e-08, 2.593871e-08, 2.59524e-08, 2.592697e-08, 
    2.587923e-08, 2.572532e-08, 2.572784e-08, 2.5394e-08, 2.56642e-08,
  2.593443e-08, 2.584368e-08, 2.598962e-08, 2.584106e-08, 2.619561e-08, 
    2.606695e-08, 2.642236e-08, 2.613786e-08, 2.594066e-08, 2.60258e-08, 
    2.594557e-08, 2.566576e-08, 2.548771e-08, 2.519427e-08, 2.512031e-08,
  2.590725e-08, 2.603577e-08, 2.600969e-08, 2.627877e-08, 2.642227e-08, 
    2.663612e-08, 2.657301e-08, 2.664356e-08, 2.667069e-08, 2.652007e-08, 
    2.614546e-08, 2.581398e-08, 2.53663e-08, 2.533576e-08, 2.524484e-08,
  2.600904e-08, 2.616944e-08, 2.654331e-08, 2.687987e-08, 2.721129e-08, 
    2.721607e-08, 2.705815e-08, 2.706646e-08, 2.681069e-08, 2.654854e-08, 
    2.593506e-08, 2.559371e-08, 2.519685e-08, 2.538683e-08, 2.555838e-08,
  2.624501e-08, 2.66636e-08, 2.714349e-08, 2.740039e-08, 2.757458e-08, 
    2.742874e-08, 2.754114e-08, 2.775376e-08, 2.730897e-08, 2.663622e-08, 
    2.589657e-08, 2.543757e-08, 2.51829e-08, 2.555183e-08, 2.607982e-08,
  2.639798e-08, 2.682413e-08, 2.71801e-08, 2.751454e-08, 2.771766e-08, 
    2.773957e-08, 2.810395e-08, 2.820602e-08, 2.726663e-08, 2.638425e-08, 
    2.615426e-08, 2.504407e-08, 2.468252e-08, 2.549302e-08, 2.605042e-08,
  2.654698e-08, 2.6923e-08, 2.725637e-08, 2.748954e-08, 2.765516e-08, 
    2.782327e-08, 2.823498e-08, 2.835589e-08, 2.650768e-08, 2.630818e-08, 
    2.473811e-08, 2.285091e-08, 2.41086e-08, 2.598231e-08, 2.704491e-08,
  2.591481e-08, 2.592944e-08, 2.596828e-08, 2.599384e-08, 2.598935e-08, 
    2.599568e-08, 2.599871e-08, 2.595775e-08, 2.5946e-08, 2.590358e-08, 
    2.5827e-08, 2.570596e-08, 2.561759e-08, 2.548832e-08, 2.533557e-08,
  2.607674e-08, 2.599942e-08, 2.606414e-08, 2.593501e-08, 2.604255e-08, 
    2.59669e-08, 2.596921e-08, 2.598229e-08, 2.60026e-08, 2.599068e-08, 
    2.607206e-08, 2.5974e-08, 2.617619e-08, 2.620339e-08, 2.602811e-08,
  2.591712e-08, 2.582511e-08, 2.58548e-08, 2.574357e-08, 2.605055e-08, 
    2.570098e-08, 2.57727e-08, 2.581941e-08, 2.588769e-08, 2.592026e-08, 
    2.594403e-08, 2.596516e-08, 2.596072e-08, 2.596996e-08, 2.610498e-08,
  2.600845e-08, 2.606412e-08, 2.60411e-08, 2.625045e-08, 2.606506e-08, 
    2.694314e-08, 2.64383e-08, 2.658865e-08, 2.666613e-08, 2.664343e-08, 
    2.661262e-08, 2.649833e-08, 2.643046e-08, 2.617616e-08, 2.636158e-08,
  2.630841e-08, 2.647093e-08, 2.672072e-08, 2.672846e-08, 2.722961e-08, 
    2.686589e-08, 2.785979e-08, 2.733495e-08, 2.680098e-08, 2.700077e-08, 
    2.695647e-08, 2.696131e-08, 2.685515e-08, 2.674769e-08, 2.643396e-08,
  2.669047e-08, 2.694821e-08, 2.70188e-08, 2.749565e-08, 2.71516e-08, 
    2.723433e-08, 2.682639e-08, 2.704652e-08, 2.728283e-08, 2.743926e-08, 
    2.722742e-08, 2.717293e-08, 2.720669e-08, 2.725258e-08, 2.705256e-08,
  2.687294e-08, 2.714158e-08, 2.714768e-08, 2.689949e-08, 2.648735e-08, 
    2.633236e-08, 2.665663e-08, 2.706319e-08, 2.743385e-08, 2.732414e-08, 
    2.727914e-08, 2.711508e-08, 2.722833e-08, 2.73454e-08, 2.734953e-08,
  2.713729e-08, 2.681252e-08, 2.587332e-08, 2.568373e-08, 2.526712e-08, 
    2.56302e-08, 2.612722e-08, 2.657066e-08, 2.668211e-08, 2.77248e-08, 
    2.785302e-08, 2.773523e-08, 2.765061e-08, 2.758227e-08, 2.749552e-08,
  2.646623e-08, 2.579891e-08, 2.530165e-08, 2.477131e-08, 2.460615e-08, 
    2.569163e-08, 2.630691e-08, 2.655181e-08, 2.734031e-08, 2.806322e-08, 
    2.735301e-08, 2.735342e-08, 2.747957e-08, 2.758399e-08, 2.736108e-08,
  2.618446e-08, 2.546502e-08, 2.49191e-08, 2.434001e-08, 2.471366e-08, 
    2.632703e-08, 2.634359e-08, 2.63805e-08, 2.678359e-08, 2.607377e-08, 
    2.519664e-08, 2.495213e-08, 2.485784e-08, 2.545504e-08, 2.618151e-08,
  2.623457e-08, 2.633463e-08, 2.623477e-08, 2.621711e-08, 2.60782e-08, 
    2.596137e-08, 2.591654e-08, 2.583937e-08, 2.577889e-08, 2.576705e-08, 
    2.568954e-08, 2.563359e-08, 2.562091e-08, 2.56111e-08, 2.562216e-08,
  2.637127e-08, 2.628033e-08, 2.624971e-08, 2.61425e-08, 2.60217e-08, 
    2.587144e-08, 2.576521e-08, 2.569443e-08, 2.573032e-08, 2.568451e-08, 
    2.578126e-08, 2.569056e-08, 2.585936e-08, 2.583219e-08, 2.5721e-08,
  2.616192e-08, 2.626977e-08, 2.635512e-08, 2.628333e-08, 2.644749e-08, 
    2.614724e-08, 2.621362e-08, 2.623583e-08, 2.630376e-08, 2.62602e-08, 
    2.62603e-08, 2.618514e-08, 2.623685e-08, 2.602809e-08, 2.612157e-08,
  2.646803e-08, 2.665779e-08, 2.669391e-08, 2.69521e-08, 2.672111e-08, 
    2.72892e-08, 2.653842e-08, 2.641641e-08, 2.630082e-08, 2.619862e-08, 
    2.643077e-08, 2.622375e-08, 2.672978e-08, 2.6557e-08, 2.682662e-08,
  2.701634e-08, 2.70932e-08, 2.694629e-08, 2.656164e-08, 2.572627e-08, 
    2.496963e-08, 2.51469e-08, 2.461193e-08, 2.390679e-08, 2.391723e-08, 
    2.40176e-08, 2.409167e-08, 2.447398e-08, 2.473941e-08, 2.508188e-08,
  2.712138e-08, 2.667842e-08, 2.615093e-08, 2.516537e-08, 2.397533e-08, 
    2.354339e-08, 2.290046e-08, 2.324652e-08, 2.357821e-08, 2.466325e-08, 
    2.49614e-08, 2.523467e-08, 2.534022e-08, 2.568885e-08, 2.528268e-08,
  2.656606e-08, 2.652153e-08, 2.592583e-08, 2.469237e-08, 2.394151e-08, 
    2.364766e-08, 2.464498e-08, 2.592162e-08, 2.624767e-08, 2.700168e-08, 
    2.658964e-08, 2.669095e-08, 2.67368e-08, 2.70578e-08, 2.663187e-08,
  2.72182e-08, 2.67641e-08, 2.588925e-08, 2.465858e-08, 2.459475e-08, 
    2.592484e-08, 2.664438e-08, 2.690931e-08, 2.646669e-08, 2.677955e-08, 
    2.636561e-08, 2.652363e-08, 2.656216e-08, 2.702571e-08, 2.671596e-08,
  2.733018e-08, 2.63856e-08, 2.499261e-08, 2.454756e-08, 2.583211e-08, 
    2.673171e-08, 2.658876e-08, 2.671636e-08, 2.672942e-08, 2.700453e-08, 
    2.700806e-08, 2.691112e-08, 2.70651e-08, 2.706427e-08, 2.690305e-08,
  2.68501e-08, 2.563559e-08, 2.474228e-08, 2.488963e-08, 2.661458e-08, 
    2.694648e-08, 2.681055e-08, 2.718177e-08, 2.736272e-08, 2.741737e-08, 
    2.744902e-08, 2.729123e-08, 2.681698e-08, 2.643718e-08, 2.620828e-08,
  2.621914e-08, 2.64479e-08, 2.657757e-08, 2.672456e-08, 2.679468e-08, 
    2.683373e-08, 2.685901e-08, 2.674593e-08, 2.68348e-08, 2.667282e-08, 
    2.670231e-08, 2.659336e-08, 2.655928e-08, 2.637567e-08, 2.621796e-08,
  2.635918e-08, 2.646131e-08, 2.657704e-08, 2.64238e-08, 2.66014e-08, 
    2.659226e-08, 2.665646e-08, 2.6888e-08, 2.693655e-08, 2.694583e-08, 
    2.688874e-08, 2.66441e-08, 2.670553e-08, 2.654068e-08, 2.635746e-08,
  2.643929e-08, 2.639349e-08, 2.644987e-08, 2.643412e-08, 2.709431e-08, 
    2.672155e-08, 2.702456e-08, 2.694936e-08, 2.707418e-08, 2.69811e-08, 
    2.691686e-08, 2.687409e-08, 2.688761e-08, 2.676355e-08, 2.677996e-08,
  2.64934e-08, 2.638947e-08, 2.656326e-08, 2.711801e-08, 2.705377e-08, 
    2.767846e-08, 2.710781e-08, 2.697355e-08, 2.67564e-08, 2.692969e-08, 
    2.666924e-08, 2.690755e-08, 2.67736e-08, 2.690461e-08, 2.697666e-08,
  2.61395e-08, 2.662149e-08, 2.730182e-08, 2.726834e-08, 2.742671e-08, 
    2.707273e-08, 2.763322e-08, 2.74925e-08, 2.728625e-08, 2.707103e-08, 
    2.646857e-08, 2.618981e-08, 2.590828e-08, 2.570018e-08, 2.54262e-08,
  2.71686e-08, 2.754738e-08, 2.749252e-08, 2.717972e-08, 2.697793e-08, 
    2.670196e-08, 2.669895e-08, 2.727648e-08, 2.791213e-08, 2.777625e-08, 
    2.771255e-08, 2.737486e-08, 2.736891e-08, 2.706492e-08, 2.681744e-08,
  2.750049e-08, 2.720802e-08, 2.684063e-08, 2.673602e-08, 2.683423e-08, 
    2.735551e-08, 2.870207e-08, 2.919725e-08, 2.892932e-08, 2.864027e-08, 
    2.813731e-08, 2.80758e-08, 2.786568e-08, 2.780683e-08, 2.761592e-08,
  2.713935e-08, 2.665086e-08, 2.731351e-08, 2.700463e-08, 2.777306e-08, 
    2.954157e-08, 2.973751e-08, 2.871505e-08, 2.785084e-08, 2.782821e-08, 
    2.767938e-08, 2.794271e-08, 2.765224e-08, 2.782165e-08, 2.748099e-08,
  2.699434e-08, 2.730885e-08, 2.751918e-08, 2.716528e-08, 3.052113e-08, 
    3.040736e-08, 2.857118e-08, 2.776635e-08, 2.805529e-08, 2.844979e-08, 
    2.845971e-08, 2.853701e-08, 2.84373e-08, 2.856836e-08, 2.846117e-08,
  2.740711e-08, 2.778551e-08, 2.748165e-08, 3.006889e-08, 3.205506e-08, 
    2.910654e-08, 2.732951e-08, 2.761318e-08, 2.811745e-08, 2.821517e-08, 
    2.796441e-08, 2.790308e-08, 2.77255e-08, 2.752963e-08, 2.787702e-08,
  2.762273e-08, 2.743007e-08, 2.729325e-08, 2.706516e-08, 2.720848e-08, 
    2.707514e-08, 2.714015e-08, 2.690101e-08, 2.679679e-08, 2.675185e-08, 
    2.696346e-08, 2.698833e-08, 2.74944e-08, 2.763345e-08, 2.780838e-08,
  2.700563e-08, 2.696327e-08, 2.691963e-08, 2.676645e-08, 2.688143e-08, 
    2.65611e-08, 2.683019e-08, 2.647711e-08, 2.706756e-08, 2.719236e-08, 
    2.780861e-08, 2.770473e-08, 2.839071e-08, 2.830895e-08, 2.839988e-08,
  2.63522e-08, 2.637021e-08, 2.635256e-08, 2.628789e-08, 2.665237e-08, 
    2.647698e-08, 2.669924e-08, 2.693323e-08, 2.788969e-08, 2.764623e-08, 
    2.80113e-08, 2.799286e-08, 2.850841e-08, 2.811091e-08, 2.850966e-08,
  2.639641e-08, 2.629154e-08, 2.632651e-08, 2.644824e-08, 2.653925e-08, 
    2.729296e-08, 2.721595e-08, 2.797306e-08, 2.800552e-08, 2.806138e-08, 
    2.865911e-08, 2.883975e-08, 2.893981e-08, 2.825619e-08, 2.829647e-08,
  2.66336e-08, 2.676751e-08, 2.687185e-08, 2.713014e-08, 2.76825e-08, 
    2.754306e-08, 2.855467e-08, 2.872623e-08, 2.852374e-08, 2.909493e-08, 
    2.951055e-08, 2.915292e-08, 2.828699e-08, 2.779878e-08, 2.729218e-08,
  2.706926e-08, 2.751655e-08, 2.761715e-08, 2.804938e-08, 2.82146e-08, 
    2.808059e-08, 2.830991e-08, 2.894538e-08, 2.985476e-08, 2.925392e-08, 
    2.801773e-08, 2.67409e-08, 2.646735e-08, 2.634158e-08, 2.65942e-08,
  2.802057e-08, 2.804644e-08, 2.830488e-08, 2.843006e-08, 2.820088e-08, 
    2.79127e-08, 2.964332e-08, 2.955001e-08, 2.843032e-08, 2.65134e-08, 
    2.581081e-08, 2.595928e-08, 2.621612e-08, 2.669252e-08, 2.71113e-08,
  2.784069e-08, 2.795753e-08, 2.82617e-08, 2.797162e-08, 2.771323e-08, 
    2.910858e-08, 2.965085e-08, 2.804304e-08, 2.60432e-08, 2.549962e-08, 
    2.573075e-08, 2.640962e-08, 2.662778e-08, 2.700724e-08, 2.698317e-08,
  2.774084e-08, 2.801777e-08, 2.8113e-08, 2.777063e-08, 2.878228e-08, 
    2.909061e-08, 2.686275e-08, 2.556078e-08, 2.541907e-08, 2.567452e-08, 
    2.664573e-08, 2.670268e-08, 2.685954e-08, 2.711539e-08, 2.700179e-08,
  2.789895e-08, 2.779805e-08, 2.74975e-08, 2.808344e-08, 2.845045e-08, 
    2.643956e-08, 2.531892e-08, 2.533443e-08, 2.60256e-08, 2.668812e-08, 
    2.694267e-08, 2.699531e-08, 2.748639e-08, 2.738802e-08, 2.710281e-08,
  2.688949e-08, 2.693802e-08, 2.687108e-08, 2.694873e-08, 2.668671e-08, 
    2.677226e-08, 2.678286e-08, 2.682541e-08, 2.683827e-08, 2.670177e-08, 
    2.695424e-08, 2.700944e-08, 2.723289e-08, 2.740566e-08, 2.749622e-08,
  2.677424e-08, 2.688121e-08, 2.680596e-08, 2.686315e-08, 2.672855e-08, 
    2.676829e-08, 2.681039e-08, 2.674909e-08, 2.662585e-08, 2.690709e-08, 
    2.711159e-08, 2.706658e-08, 2.745425e-08, 2.731814e-08, 2.760079e-08,
  2.69641e-08, 2.673167e-08, 2.7069e-08, 2.651215e-08, 2.680395e-08, 
    2.685647e-08, 2.643632e-08, 2.671435e-08, 2.672275e-08, 2.695571e-08, 
    2.703952e-08, 2.718901e-08, 2.7637e-08, 2.766249e-08, 2.817812e-08,
  2.686389e-08, 2.694232e-08, 2.680492e-08, 2.705881e-08, 2.650591e-08, 
    2.675574e-08, 2.668514e-08, 2.675963e-08, 2.732015e-08, 2.727656e-08, 
    2.77806e-08, 2.805596e-08, 2.801021e-08, 2.786643e-08, 2.739703e-08,
  2.690557e-08, 2.685017e-08, 2.724126e-08, 2.701075e-08, 2.749326e-08, 
    2.696927e-08, 2.741938e-08, 2.763688e-08, 2.765322e-08, 2.780852e-08, 
    2.815159e-08, 2.787887e-08, 2.743662e-08, 2.703006e-08, 2.645412e-08,
  2.67975e-08, 2.704134e-08, 2.727052e-08, 2.731802e-08, 2.75293e-08, 
    2.764886e-08, 2.770236e-08, 2.772848e-08, 2.762494e-08, 2.78595e-08, 
    2.746861e-08, 2.684085e-08, 2.676042e-08, 2.647977e-08, 2.713404e-08,
  2.681404e-08, 2.715831e-08, 2.710219e-08, 2.741443e-08, 2.747169e-08, 
    2.759597e-08, 2.752256e-08, 2.744012e-08, 2.714951e-08, 2.670893e-08, 
    2.647757e-08, 2.634239e-08, 2.704512e-08, 2.757792e-08, 2.861508e-08,
  2.65419e-08, 2.647701e-08, 2.663695e-08, 2.663514e-08, 2.675947e-08, 
    2.657226e-08, 2.655064e-08, 2.643447e-08, 2.630841e-08, 2.627418e-08, 
    2.672726e-08, 2.732055e-08, 2.826239e-08, 2.827133e-08, 2.825302e-08,
  2.625934e-08, 2.628063e-08, 2.632965e-08, 2.632326e-08, 2.608563e-08, 
    2.603344e-08, 2.582607e-08, 2.601519e-08, 2.639488e-08, 2.69545e-08, 
    2.792919e-08, 2.805993e-08, 2.811276e-08, 2.772593e-08, 2.754815e-08,
  2.638275e-08, 2.635131e-08, 2.61649e-08, 2.596757e-08, 2.591912e-08, 
    2.596983e-08, 2.643539e-08, 2.686059e-08, 2.752569e-08, 2.792517e-08, 
    2.79382e-08, 2.758784e-08, 2.740931e-08, 2.709107e-08, 2.756098e-08,
  2.564266e-08, 2.571579e-08, 2.577637e-08, 2.59461e-08, 2.597708e-08, 
    2.620575e-08, 2.635889e-08, 2.650515e-08, 2.66425e-08, 2.641838e-08, 
    2.614328e-08, 2.613105e-08, 2.573426e-08, 2.55381e-08, 2.593271e-08,
  2.567306e-08, 2.586926e-08, 2.581444e-08, 2.594754e-08, 2.590444e-08, 
    2.611479e-08, 2.626205e-08, 2.651722e-08, 2.668334e-08, 2.670738e-08, 
    2.683572e-08, 2.645149e-08, 2.679386e-08, 2.662877e-08, 2.707514e-08,
  2.619453e-08, 2.599416e-08, 2.624907e-08, 2.596472e-08, 2.617126e-08, 
    2.613658e-08, 2.624932e-08, 2.65176e-08, 2.667944e-08, 2.67326e-08, 
    2.69191e-08, 2.68396e-08, 2.706965e-08, 2.671622e-08, 2.69389e-08,
  2.643164e-08, 2.602707e-08, 2.63454e-08, 2.611414e-08, 2.619943e-08, 
    2.619346e-08, 2.606795e-08, 2.638897e-08, 2.669694e-08, 2.685614e-08, 
    2.689133e-08, 2.695794e-08, 2.697244e-08, 2.68486e-08, 2.69583e-08,
  2.641082e-08, 2.646322e-08, 2.629756e-08, 2.644491e-08, 2.617378e-08, 
    2.636103e-08, 2.633683e-08, 2.616138e-08, 2.659399e-08, 2.665112e-08, 
    2.689155e-08, 2.693642e-08, 2.710343e-08, 2.723124e-08, 2.738668e-08,
  2.692891e-08, 2.652683e-08, 2.672744e-08, 2.6465e-08, 2.648869e-08, 
    2.61824e-08, 2.632182e-08, 2.635497e-08, 2.604374e-08, 2.623625e-08, 
    2.654921e-08, 2.672217e-08, 2.69477e-08, 2.708559e-08, 2.714328e-08,
  2.715207e-08, 2.658047e-08, 2.708883e-08, 2.635371e-08, 2.66915e-08, 
    2.621619e-08, 2.641137e-08, 2.614139e-08, 2.634491e-08, 2.639204e-08, 
    2.645788e-08, 2.650644e-08, 2.649265e-08, 2.661297e-08, 2.663818e-08,
  2.695024e-08, 2.689998e-08, 2.6853e-08, 2.653693e-08, 2.643308e-08, 
    2.631432e-08, 2.621896e-08, 2.618006e-08, 2.611134e-08, 2.60892e-08, 
    2.608213e-08, 2.633393e-08, 2.649779e-08, 2.68512e-08, 2.687929e-08,
  2.698494e-08, 2.726855e-08, 2.696628e-08, 2.685731e-08, 2.678424e-08, 
    2.663039e-08, 2.6625e-08, 2.653552e-08, 2.6625e-08, 2.673178e-08, 
    2.694612e-08, 2.695201e-08, 2.692213e-08, 2.685674e-08, 2.677533e-08,
  2.686599e-08, 2.671896e-08, 2.706631e-08, 2.707992e-08, 2.689575e-08, 
    2.69135e-08, 2.686691e-08, 2.683956e-08, 2.684394e-08, 2.664786e-08, 
    2.654924e-08, 2.63774e-08, 2.648395e-08, 2.657388e-08, 2.693038e-08,
  2.645378e-08, 2.655583e-08, 2.668572e-08, 2.667194e-08, 2.667583e-08, 
    2.655881e-08, 2.655788e-08, 2.623121e-08, 2.657763e-08, 2.651516e-08, 
    2.658584e-08, 2.690464e-08, 2.682066e-08, 2.691381e-08, 2.688679e-08,
  2.669379e-08, 2.690097e-08, 2.704237e-08, 2.705586e-08, 2.704734e-08, 
    2.679174e-08, 2.681131e-08, 2.635725e-08, 2.616612e-08, 2.641367e-08, 
    2.653162e-08, 2.640205e-08, 2.681572e-08, 2.651866e-08, 2.686184e-08,
  2.702024e-08, 2.723326e-08, 2.728672e-08, 2.720134e-08, 2.73806e-08, 
    2.670291e-08, 2.649947e-08, 2.65773e-08, 2.617325e-08, 2.605089e-08, 
    2.630701e-08, 2.629284e-08, 2.663364e-08, 2.661841e-08, 2.647551e-08,
  2.729026e-08, 2.729104e-08, 2.715184e-08, 2.694702e-08, 2.686192e-08, 
    2.707155e-08, 2.631527e-08, 2.618589e-08, 2.624706e-08, 2.588597e-08, 
    2.5885e-08, 2.586645e-08, 2.624423e-08, 2.634093e-08, 2.665212e-08,
  2.728814e-08, 2.716129e-08, 2.697741e-08, 2.679513e-08, 2.689613e-08, 
    2.671778e-08, 2.693112e-08, 2.613168e-08, 2.610064e-08, 2.611573e-08, 
    2.610981e-08, 2.592342e-08, 2.60927e-08, 2.610496e-08, 2.642586e-08,
  2.74457e-08, 2.719808e-08, 2.709892e-08, 2.705105e-08, 2.703964e-08, 
    2.690129e-08, 2.701696e-08, 2.671829e-08, 2.620865e-08, 2.592724e-08, 
    2.602983e-08, 2.595444e-08, 2.584695e-08, 2.60091e-08, 2.59328e-08,
  2.715592e-08, 2.724847e-08, 2.731386e-08, 2.722139e-08, 2.705756e-08, 
    2.682801e-08, 2.679345e-08, 2.66754e-08, 2.649104e-08, 2.60886e-08, 
    2.595316e-08, 2.600629e-08, 2.586813e-08, 2.605375e-08, 2.569195e-08,
  2.719291e-08, 2.736642e-08, 2.735249e-08, 2.724727e-08, 2.722727e-08, 
    2.713166e-08, 2.704396e-08, 2.68594e-08, 2.677035e-08, 2.661077e-08, 
    2.641382e-08, 2.625208e-08, 2.594984e-08, 2.624282e-08, 2.599385e-08,
  2.703036e-08, 2.723939e-08, 2.742424e-08, 2.741293e-08, 2.754126e-08, 
    2.749333e-08, 2.74677e-08, 2.713577e-08, 2.700169e-08, 2.693317e-08, 
    2.676052e-08, 2.673313e-08, 2.647139e-08, 2.651138e-08, 2.643923e-08,
  2.686661e-08, 2.707794e-08, 2.721774e-08, 2.729617e-08, 2.751913e-08, 
    2.775274e-08, 2.787917e-08, 2.755609e-08, 2.751768e-08, 2.722163e-08, 
    2.70377e-08, 2.69616e-08, 2.679988e-08, 2.675758e-08, 2.667991e-08,
  2.607121e-08, 2.611674e-08, 2.629706e-08, 2.657907e-08, 2.685274e-08, 
    2.717532e-08, 2.735762e-08, 2.750016e-08, 2.758202e-08, 2.76055e-08, 
    2.756002e-08, 2.756977e-08, 2.723942e-08, 2.71033e-08, 2.686901e-08,
  2.642171e-08, 2.670865e-08, 2.713295e-08, 2.72211e-08, 2.769222e-08, 
    2.758249e-08, 2.76109e-08, 2.766062e-08, 2.765532e-08, 2.755524e-08, 
    2.77734e-08, 2.747383e-08, 2.773686e-08, 2.716011e-08, 2.706662e-08,
  2.670872e-08, 2.693034e-08, 2.706996e-08, 2.722354e-08, 2.774774e-08, 
    2.728785e-08, 2.734851e-08, 2.74745e-08, 2.751655e-08, 2.749388e-08, 
    2.75355e-08, 2.740837e-08, 2.730673e-08, 2.712039e-08, 2.705051e-08,
  2.67388e-08, 2.692801e-08, 2.716222e-08, 2.729142e-08, 2.726564e-08, 
    2.792583e-08, 2.751493e-08, 2.756204e-08, 2.733492e-08, 2.738058e-08, 
    2.739842e-08, 2.714865e-08, 2.699034e-08, 2.677086e-08, 2.70181e-08,
  2.69759e-08, 2.712431e-08, 2.725514e-08, 2.729627e-08, 2.763864e-08, 
    2.742389e-08, 2.817413e-08, 2.756924e-08, 2.737325e-08, 2.734141e-08, 
    2.712737e-08, 2.68649e-08, 2.660665e-08, 2.638606e-08, 2.636601e-08,
  2.679454e-08, 2.704235e-08, 2.726097e-08, 2.751947e-08, 2.762003e-08, 
    2.788227e-08, 2.772387e-08, 2.813984e-08, 2.82519e-08, 2.798558e-08, 
    2.768446e-08, 2.713647e-08, 2.682055e-08, 2.652264e-08, 2.622088e-08,
  2.673517e-08, 2.701122e-08, 2.728416e-08, 2.751473e-08, 2.79535e-08, 
    2.800276e-08, 2.831822e-08, 2.81976e-08, 2.804073e-08, 2.811059e-08, 
    2.778649e-08, 2.738068e-08, 2.689682e-08, 2.66017e-08, 2.613687e-08,
  2.672515e-08, 2.713059e-08, 2.737305e-08, 2.768596e-08, 2.795379e-08, 
    2.827157e-08, 2.850123e-08, 2.850559e-08, 2.865895e-08, 2.893296e-08, 
    2.848555e-08, 2.800734e-08, 2.716787e-08, 2.68505e-08, 2.624851e-08,
  2.690513e-08, 2.719477e-08, 2.747428e-08, 2.767301e-08, 2.795177e-08, 
    2.798514e-08, 2.836526e-08, 2.85886e-08, 2.915609e-08, 2.931647e-08, 
    2.841678e-08, 2.765157e-08, 2.707577e-08, 2.695071e-08, 2.653363e-08,
  2.692938e-08, 2.725427e-08, 2.757876e-08, 2.777752e-08, 2.775773e-08, 
    2.777121e-08, 2.795911e-08, 2.83469e-08, 2.930344e-08, 2.910898e-08, 
    2.757817e-08, 2.684948e-08, 2.708032e-08, 2.689126e-08, 2.663669e-08,
  2.432009e-08, 2.463862e-08, 2.508446e-08, 2.53944e-08, 2.572459e-08, 
    2.591047e-08, 2.606783e-08, 2.614449e-08, 2.62129e-08, 2.631404e-08, 
    2.651975e-08, 2.673657e-08, 2.699552e-08, 2.737082e-08, 2.743836e-08,
  2.516183e-08, 2.505945e-08, 2.523685e-08, 2.509287e-08, 2.550688e-08, 
    2.54946e-08, 2.597309e-08, 2.609467e-08, 2.659932e-08, 2.671914e-08, 
    2.73122e-08, 2.734054e-08, 2.804455e-08, 2.795661e-08, 2.78944e-08,
  2.638368e-08, 2.623696e-08, 2.657706e-08, 2.615617e-08, 2.65151e-08, 
    2.682582e-08, 2.709732e-08, 2.720122e-08, 2.752882e-08, 2.767023e-08, 
    2.791868e-08, 2.808466e-08, 2.834497e-08, 2.817598e-08, 2.837881e-08,
  2.734236e-08, 2.744303e-08, 2.732799e-08, 2.735534e-08, 2.716627e-08, 
    2.738458e-08, 2.764466e-08, 2.795815e-08, 2.813271e-08, 2.80646e-08, 
    2.827469e-08, 2.815732e-08, 2.839294e-08, 2.816899e-08, 2.850385e-08,
  2.792057e-08, 2.801185e-08, 2.779171e-08, 2.789195e-08, 2.806488e-08, 
    2.78671e-08, 2.816475e-08, 2.831539e-08, 2.813456e-08, 2.788894e-08, 
    2.783809e-08, 2.799316e-08, 2.820664e-08, 2.819004e-08, 2.800631e-08,
  2.787935e-08, 2.783764e-08, 2.788742e-08, 2.804666e-08, 2.781994e-08, 
    2.797022e-08, 2.766073e-08, 2.755222e-08, 2.755722e-08, 2.76874e-08, 
    2.770363e-08, 2.794369e-08, 2.806753e-08, 2.812058e-08, 2.803629e-08,
  2.757987e-08, 2.750099e-08, 2.74158e-08, 2.736953e-08, 2.728341e-08, 
    2.737407e-08, 2.725762e-08, 2.69982e-08, 2.691679e-08, 2.684206e-08, 
    2.73215e-08, 2.790312e-08, 2.811757e-08, 2.839252e-08, 2.825929e-08,
  2.765294e-08, 2.73202e-08, 2.723223e-08, 2.724203e-08, 2.718108e-08, 
    2.750698e-08, 2.707894e-08, 2.703169e-08, 2.719484e-08, 2.735636e-08, 
    2.79986e-08, 2.809013e-08, 2.814105e-08, 2.845005e-08, 2.8419e-08,
  2.762029e-08, 2.738464e-08, 2.742005e-08, 2.739526e-08, 2.751482e-08, 
    2.749727e-08, 2.675985e-08, 2.719112e-08, 2.747275e-08, 2.758557e-08, 
    2.787689e-08, 2.76736e-08, 2.779603e-08, 2.785394e-08, 2.800794e-08,
  2.798243e-08, 2.730297e-08, 2.711297e-08, 2.709683e-08, 2.726106e-08, 
    2.745405e-08, 2.698896e-08, 2.769166e-08, 2.790939e-08, 2.745257e-08, 
    2.790668e-08, 2.770361e-08, 2.806412e-08, 2.783294e-08, 2.780272e-08,
  2.556846e-08, 2.522563e-08, 2.566054e-08, 2.621417e-08, 2.683699e-08, 
    2.716861e-08, 2.615785e-08, 2.693337e-08, 2.751377e-08, 2.791946e-08, 
    2.804418e-08, 2.809201e-08, 2.78443e-08, 2.776357e-08, 2.755529e-08,
  2.562059e-08, 2.569148e-08, 2.529509e-08, 2.598918e-08, 2.560141e-08, 
    2.644957e-08, 2.634499e-08, 2.618128e-08, 2.651878e-08, 2.671143e-08, 
    2.666535e-08, 2.647291e-08, 2.669483e-08, 2.65038e-08, 2.668844e-08,
  2.668534e-08, 2.584559e-08, 2.57579e-08, 2.506272e-08, 2.595517e-08, 
    2.522348e-08, 2.572952e-08, 2.566802e-08, 2.57925e-08, 2.596598e-08, 
    2.622664e-08, 2.64605e-08, 2.691789e-08, 2.704681e-08, 2.778675e-08,
  2.721607e-08, 2.712981e-08, 2.695009e-08, 2.641186e-08, 2.567564e-08, 
    2.617749e-08, 2.561216e-08, 2.598921e-08, 2.648849e-08, 2.664461e-08, 
    2.687339e-08, 2.730853e-08, 2.749171e-08, 2.781235e-08, 2.813255e-08,
  2.696764e-08, 2.744117e-08, 2.777121e-08, 2.786124e-08, 2.784269e-08, 
    2.715196e-08, 2.773041e-08, 2.739223e-08, 2.781335e-08, 2.746459e-08, 
    2.768592e-08, 2.783855e-08, 2.7625e-08, 2.807714e-08, 2.762116e-08,
  2.718817e-08, 2.694034e-08, 2.714558e-08, 2.716473e-08, 2.770038e-08, 
    2.739509e-08, 2.770053e-08, 2.74639e-08, 2.745511e-08, 2.743383e-08, 
    2.775674e-08, 2.770289e-08, 2.789758e-08, 2.814509e-08, 2.835928e-08,
  2.761423e-08, 2.749355e-08, 2.735985e-08, 2.716565e-08, 2.730893e-08, 
    2.736897e-08, 2.768784e-08, 2.759227e-08, 2.773382e-08, 2.802448e-08, 
    2.816425e-08, 2.847161e-08, 2.878505e-08, 2.906583e-08, 2.928692e-08,
  2.752092e-08, 2.771354e-08, 2.782495e-08, 2.782529e-08, 2.795148e-08, 
    2.802695e-08, 2.806172e-08, 2.806243e-08, 2.822728e-08, 2.839606e-08, 
    2.879187e-08, 2.917803e-08, 2.924611e-08, 2.932974e-08, 2.91446e-08,
  2.700204e-08, 2.708703e-08, 2.700675e-08, 2.705292e-08, 2.717672e-08, 
    2.743979e-08, 2.746004e-08, 2.795364e-08, 2.829721e-08, 2.967839e-08, 
    2.956224e-08, 2.928404e-08, 2.910468e-08, 2.914724e-08, 2.849086e-08,
  2.671577e-08, 2.67189e-08, 2.652265e-08, 2.649243e-08, 2.68647e-08, 
    2.735976e-08, 2.775269e-08, 2.815888e-08, 2.95303e-08, 2.905825e-08, 
    2.830442e-08, 2.812613e-08, 2.821802e-08, 2.813164e-08, 2.782598e-08,
  2.757743e-08, 2.744714e-08, 2.672049e-08, 2.737448e-08, 2.632587e-08, 
    2.472859e-08, 2.255716e-08, 2.583592e-08, 2.908011e-08, 2.94001e-08, 
    2.919009e-08, 2.920342e-08, 2.900687e-08, 2.79039e-08, 2.745324e-08,
  2.741917e-08, 2.750597e-08, 2.630289e-08, 2.626685e-08, 2.747976e-08, 
    2.569823e-08, 2.21228e-08, 2.668438e-08, 2.924021e-08, 3.00517e-08, 
    3.000722e-08, 2.958083e-08, 2.830484e-08, 2.771529e-08, 2.897204e-08,
  2.708286e-08, 2.715356e-08, 2.666238e-08, 2.632745e-08, 2.613652e-08, 
    2.557102e-08, 2.482824e-08, 2.4345e-08, 2.728835e-08, 2.883923e-08, 
    2.85545e-08, 2.795678e-08, 2.76771e-08, 2.867882e-08, 3.01693e-08,
  2.667493e-08, 2.68445e-08, 2.699363e-08, 2.604657e-08, 2.625853e-08, 
    2.553785e-08, 2.3906e-08, 2.603197e-08, 2.792595e-08, 2.674963e-08, 
    2.733196e-08, 2.776467e-08, 2.810654e-08, 2.936666e-08, 2.954798e-08,
  2.705409e-08, 2.68917e-08, 2.715061e-08, 2.668308e-08, 2.628234e-08, 
    2.582162e-08, 2.400832e-08, 2.735051e-08, 2.699365e-08, 2.680253e-08, 
    2.931928e-08, 2.822821e-08, 2.83112e-08, 2.837428e-08, 2.778468e-08,
  2.714271e-08, 2.714636e-08, 2.733596e-08, 2.697369e-08, 2.666919e-08, 
    2.621214e-08, 2.55221e-08, 2.592398e-08, 2.556513e-08, 2.839717e-08, 
    2.971173e-08, 2.900758e-08, 2.813137e-08, 2.765311e-08, 2.692231e-08,
  2.662728e-08, 2.687198e-08, 2.742925e-08, 2.731234e-08, 2.754586e-08, 
    2.687915e-08, 2.596985e-08, 2.609447e-08, 2.5404e-08, 2.688721e-08, 
    2.816416e-08, 2.798749e-08, 2.746041e-08, 2.714277e-08, 2.684993e-08,
  2.633714e-08, 2.644984e-08, 2.695031e-08, 2.721661e-08, 2.751627e-08, 
    2.812247e-08, 2.772011e-08, 2.729634e-08, 2.655785e-08, 2.650404e-08, 
    2.667477e-08, 2.668949e-08, 2.669998e-08, 2.688602e-08, 2.720991e-08,
  2.662243e-08, 2.6724e-08, 2.687536e-08, 2.717943e-08, 2.717531e-08, 
    2.752483e-08, 2.798187e-08, 2.839408e-08, 2.799409e-08, 2.766976e-08, 
    2.733771e-08, 2.738766e-08, 2.73936e-08, 2.762001e-08, 2.778343e-08,
  2.692089e-08, 2.695641e-08, 2.689808e-08, 2.725327e-08, 2.741759e-08, 
    2.740701e-08, 2.737226e-08, 2.763802e-08, 2.826119e-08, 2.828536e-08, 
    2.863949e-08, 2.797534e-08, 2.824052e-08, 2.837013e-08, 2.867061e-08,
  2.654809e-08, 2.685703e-08, 2.702924e-08, 2.722332e-08, 2.725823e-08, 
    2.711358e-08, 2.617914e-08, 2.450815e-08, 2.489927e-08, 2.443063e-08, 
    2.435566e-08, 2.599008e-08, 2.755649e-08, 2.657789e-08, 2.419926e-08,
  2.627487e-08, 2.654025e-08, 2.665688e-08, 2.688381e-08, 2.710129e-08, 
    2.684786e-08, 2.509094e-08, 2.479566e-08, 2.452432e-08, 2.457814e-08, 
    2.440833e-08, 2.657826e-08, 2.77557e-08, 2.511353e-08, 2.324684e-08,
  2.588883e-08, 2.611795e-08, 2.624788e-08, 2.670928e-08, 2.693813e-08, 
    2.631963e-08, 2.466298e-08, 2.286891e-08, 2.435235e-08, 2.497716e-08, 
    2.503944e-08, 2.686203e-08, 2.572246e-08, 2.372247e-08, 2.444715e-08,
  2.553216e-08, 2.578136e-08, 2.622324e-08, 2.651197e-08, 2.699464e-08, 
    2.602733e-08, 2.439026e-08, 2.380435e-08, 2.54581e-08, 2.503338e-08, 
    2.516539e-08, 2.614975e-08, 2.49475e-08, 2.448208e-08, 2.51916e-08,
  2.539459e-08, 2.562242e-08, 2.631163e-08, 2.646407e-08, 2.704707e-08, 
    2.644171e-08, 2.438664e-08, 2.492349e-08, 2.531851e-08, 2.250044e-08, 
    2.548436e-08, 2.551997e-08, 2.476114e-08, 2.558251e-08, 2.657376e-08,
  2.510258e-08, 2.53249e-08, 2.602345e-08, 2.636648e-08, 2.71099e-08, 
    2.676663e-08, 2.464433e-08, 2.28358e-08, 1.942982e-08, 2.370082e-08, 
    2.757286e-08, 2.588985e-08, 2.582007e-08, 2.800967e-08, 3.001856e-08,
  2.513372e-08, 2.507315e-08, 2.547139e-08, 2.652636e-08, 2.666999e-08, 
    2.766052e-08, 2.507816e-08, 2.380015e-08, 2.169539e-08, 3.041847e-08, 
    3.084858e-08, 2.657146e-08, 2.708318e-08, 2.989068e-08, 3.149828e-08,
  2.534065e-08, 2.506812e-08, 2.519891e-08, 2.648639e-08, 2.633096e-08, 
    2.796317e-08, 2.621034e-08, 2.426541e-08, 2.267447e-08, 3.197972e-08, 
    3.138382e-08, 2.738171e-08, 2.834043e-08, 3.044332e-08, 2.940419e-08,
  2.514525e-08, 2.539687e-08, 2.556252e-08, 2.592866e-08, 2.651416e-08, 
    2.765518e-08, 2.708858e-08, 2.55807e-08, 2.354662e-08, 3.127125e-08, 
    3.128151e-08, 2.859116e-08, 2.929088e-08, 2.957566e-08, 2.758489e-08,
  2.497065e-08, 2.578209e-08, 2.647513e-08, 2.608692e-08, 2.65383e-08, 
    2.737004e-08, 2.771465e-08, 2.639954e-08, 2.382663e-08, 2.953812e-08, 
    3.181677e-08, 2.982566e-08, 2.960704e-08, 2.891949e-08, 2.66853e-08,
  2.436566e-08, 2.453815e-08, 2.440285e-08, 2.451291e-08, 2.460665e-08, 
    2.467585e-08, 2.488082e-08, 2.501872e-08, 2.540575e-08, 2.572664e-08, 
    2.584943e-08, 2.594654e-08, 2.611209e-08, 2.636157e-08, 2.657288e-08,
  2.490923e-08, 2.498555e-08, 2.480033e-08, 2.484945e-08, 2.485888e-08, 
    2.503619e-08, 2.526357e-08, 2.562357e-08, 2.574154e-08, 2.591413e-08, 
    2.595449e-08, 2.586399e-08, 2.622684e-08, 2.646203e-08, 2.606897e-08,
  2.521367e-08, 2.530923e-08, 2.512814e-08, 2.512955e-08, 2.510194e-08, 
    2.515102e-08, 2.564912e-08, 2.585497e-08, 2.608532e-08, 2.571334e-08, 
    2.605388e-08, 2.580008e-08, 2.675542e-08, 2.554299e-08, 2.598191e-08,
  2.553324e-08, 2.574708e-08, 2.534802e-08, 2.547527e-08, 2.517197e-08, 
    2.54371e-08, 2.573777e-08, 2.610424e-08, 2.577421e-08, 2.561109e-08, 
    2.599217e-08, 2.635879e-08, 2.649276e-08, 2.63205e-08, 2.541431e-08,
  2.557552e-08, 2.599127e-08, 2.547161e-08, 2.557852e-08, 2.51896e-08, 
    2.559859e-08, 2.562463e-08, 2.601367e-08, 2.668323e-08, 2.560286e-08, 
    2.479048e-08, 2.566764e-08, 2.680027e-08, 2.512336e-08, 2.396972e-08,
  2.579692e-08, 2.636939e-08, 2.574009e-08, 2.581755e-08, 2.545863e-08, 
    2.532935e-08, 2.657004e-08, 2.578258e-08, 2.379964e-08, 2.411622e-08, 
    2.61014e-08, 2.794529e-08, 2.548769e-08, 2.30143e-08, 2.704294e-08,
  2.583828e-08, 2.663913e-08, 2.607599e-08, 2.606937e-08, 2.547732e-08, 
    2.564866e-08, 2.668767e-08, 2.561537e-08, 2.423888e-08, 2.526299e-08, 
    2.752855e-08, 2.691762e-08, 2.353677e-08, 2.683372e-08, 2.991592e-08,
  2.596017e-08, 2.677232e-08, 2.646733e-08, 2.652443e-08, 2.541005e-08, 
    2.598551e-08, 2.679794e-08, 2.474963e-08, 2.357635e-08, 2.600773e-08, 
    2.753933e-08, 2.526361e-08, 2.601422e-08, 2.973456e-08, 2.771566e-08,
  2.604132e-08, 2.698112e-08, 2.685232e-08, 2.685368e-08, 2.572681e-08, 
    2.585146e-08, 2.710245e-08, 2.391328e-08, 2.418864e-08, 2.451927e-08, 
    2.391563e-08, 2.544108e-08, 2.885447e-08, 2.910996e-08, 2.792676e-08,
  2.61898e-08, 2.708136e-08, 2.697126e-08, 2.694859e-08, 2.627133e-08, 
    2.599358e-08, 2.711836e-08, 2.34493e-08, 2.103781e-08, 2.079651e-08, 
    2.719681e-08, 3.040003e-08, 2.859879e-08, 2.807739e-08, 2.797004e-08,
  2.665836e-08, 2.710594e-08, 2.655362e-08, 2.665462e-08, 2.651376e-08, 
    2.614796e-08, 2.577872e-08, 2.589023e-08, 2.553763e-08, 2.492253e-08, 
    2.426515e-08, 2.425745e-08, 2.427809e-08, 2.489032e-08, 2.515911e-08,
  2.681329e-08, 2.734963e-08, 2.67193e-08, 2.674738e-08, 2.644376e-08, 
    2.606511e-08, 2.598481e-08, 2.592229e-08, 2.554683e-08, 2.510809e-08, 
    2.428228e-08, 2.395214e-08, 2.408845e-08, 2.427325e-08, 2.471342e-08,
  2.685575e-08, 2.728608e-08, 2.656093e-08, 2.663385e-08, 2.623876e-08, 
    2.562042e-08, 2.574487e-08, 2.487726e-08, 2.526772e-08, 2.500881e-08, 
    2.480346e-08, 2.4352e-08, 2.434475e-08, 2.447128e-08, 2.465799e-08,
  2.66572e-08, 2.748651e-08, 2.659982e-08, 2.640933e-08, 2.626811e-08, 
    2.588353e-08, 2.515221e-08, 2.532185e-08, 2.436475e-08, 2.471095e-08, 
    2.513569e-08, 2.544716e-08, 2.612806e-08, 2.567738e-08, 2.578253e-08,
  2.607041e-08, 2.753263e-08, 2.687301e-08, 2.597385e-08, 2.563506e-08, 
    2.529885e-08, 2.498508e-08, 2.592511e-08, 2.738905e-08, 2.590794e-08, 
    2.581026e-08, 2.542961e-08, 2.545887e-08, 2.564557e-08, 2.591121e-08,
  2.544942e-08, 2.718497e-08, 2.725801e-08, 2.593718e-08, 2.537688e-08, 
    2.52501e-08, 2.592666e-08, 2.638366e-08, 2.611301e-08, 2.610227e-08, 
    2.684726e-08, 2.713468e-08, 2.702173e-08, 2.649262e-08, 2.611875e-08,
  2.478311e-08, 2.686793e-08, 2.735942e-08, 2.611944e-08, 2.51101e-08, 
    2.482062e-08, 2.517067e-08, 2.697619e-08, 2.834394e-08, 2.917717e-08, 
    2.822842e-08, 2.707055e-08, 2.586833e-08, 2.682159e-08, 2.726242e-08,
  2.449821e-08, 2.60888e-08, 2.705519e-08, 2.66152e-08, 2.565549e-08, 
    2.500374e-08, 2.492251e-08, 2.650107e-08, 2.821346e-08, 2.822384e-08, 
    2.730503e-08, 2.672141e-08, 2.683165e-08, 2.724607e-08, 2.726693e-08,
  2.445232e-08, 2.552787e-08, 2.657834e-08, 2.701572e-08, 2.600395e-08, 
    2.513446e-08, 2.448175e-08, 2.544692e-08, 2.708349e-08, 2.729752e-08, 
    2.757833e-08, 2.680383e-08, 2.588414e-08, 2.73218e-08, 2.773295e-08,
  2.407518e-08, 2.505244e-08, 2.610846e-08, 2.714044e-08, 2.63201e-08, 
    2.534973e-08, 2.379735e-08, 2.348169e-08, 2.757427e-08, 2.993654e-08, 
    2.873133e-08, 2.724117e-08, 2.733398e-08, 2.796244e-08, 2.839478e-08,
  2.482677e-08, 2.524408e-08, 2.521356e-08, 2.523631e-08, 2.62049e-08, 
    2.697859e-08, 2.721746e-08, 2.645847e-08, 2.629083e-08, 2.63732e-08, 
    2.597072e-08, 2.591076e-08, 2.533859e-08, 2.506389e-08, 2.490385e-08,
  2.449735e-08, 2.504167e-08, 2.517166e-08, 2.526354e-08, 2.595638e-08, 
    2.676588e-08, 2.751491e-08, 2.652744e-08, 2.62098e-08, 2.629717e-08, 
    2.609026e-08, 2.582141e-08, 2.580264e-08, 2.532181e-08, 2.479653e-08,
  2.384805e-08, 2.452416e-08, 2.495862e-08, 2.483073e-08, 2.572176e-08, 
    2.672451e-08, 2.754011e-08, 2.723065e-08, 2.637143e-08, 2.622764e-08, 
    2.602224e-08, 2.551799e-08, 2.528141e-08, 2.530666e-08, 2.513276e-08,
  2.335249e-08, 2.392546e-08, 2.473896e-08, 2.482498e-08, 2.51289e-08, 
    2.712667e-08, 2.836975e-08, 2.838605e-08, 2.69678e-08, 2.672215e-08, 
    2.640487e-08, 2.600424e-08, 2.552775e-08, 2.47896e-08, 2.513382e-08,
  2.301418e-08, 2.315175e-08, 2.42257e-08, 2.473234e-08, 2.513457e-08, 
    2.56775e-08, 2.850096e-08, 2.895846e-08, 2.826956e-08, 2.727604e-08, 
    2.68303e-08, 2.703904e-08, 2.688716e-08, 2.605235e-08, 2.516277e-08,
  2.283121e-08, 2.266884e-08, 2.349557e-08, 2.465019e-08, 2.537445e-08, 
    2.604119e-08, 2.700384e-08, 2.941762e-08, 2.836941e-08, 2.725378e-08, 
    2.679365e-08, 2.702146e-08, 2.702474e-08, 2.714357e-08, 2.698596e-08,
  2.278698e-08, 2.250539e-08, 2.296775e-08, 2.406255e-08, 2.536533e-08, 
    2.623432e-08, 2.700474e-08, 2.716333e-08, 2.713084e-08, 2.699867e-08, 
    2.67199e-08, 2.681437e-08, 2.695613e-08, 2.676411e-08, 2.673612e-08,
  2.283285e-08, 2.24763e-08, 2.282153e-08, 2.366987e-08, 2.507286e-08, 
    2.633823e-08, 2.684128e-08, 2.724581e-08, 2.697661e-08, 2.636916e-08, 
    2.639986e-08, 2.684947e-08, 2.73165e-08, 2.763309e-08, 2.798744e-08,
  2.284665e-08, 2.261474e-08, 2.305267e-08, 2.362374e-08, 2.471216e-08, 
    2.646701e-08, 2.703276e-08, 2.657529e-08, 2.704439e-08, 2.693751e-08, 
    2.697331e-08, 2.776951e-08, 2.831296e-08, 2.842282e-08, 2.886647e-08,
  2.276285e-08, 2.242839e-08, 2.313375e-08, 2.412177e-08, 2.472196e-08, 
    2.636708e-08, 2.713831e-08, 2.670232e-08, 2.662512e-08, 2.713476e-08, 
    2.699378e-08, 2.74314e-08, 2.838052e-08, 2.900458e-08, 2.96873e-08,
  2.316479e-08, 2.284906e-08, 2.318959e-08, 2.48485e-08, 2.672943e-08, 
    2.820564e-08, 2.878599e-08, 2.868494e-08, 2.816658e-08, 2.779591e-08, 
    2.774333e-08, 2.713351e-08, 2.67178e-08, 2.607096e-08, 2.62895e-08,
  2.324195e-08, 2.291683e-08, 2.304178e-08, 2.437725e-08, 2.63687e-08, 
    2.84979e-08, 2.932308e-08, 2.914881e-08, 2.795744e-08, 2.759911e-08, 
    2.747739e-08, 2.738799e-08, 2.702164e-08, 2.623078e-08, 2.59146e-08,
  2.324381e-08, 2.298071e-08, 2.287063e-08, 2.413124e-08, 2.646564e-08, 
    2.892839e-08, 2.918861e-08, 2.870267e-08, 2.856938e-08, 2.745179e-08, 
    2.716305e-08, 2.728168e-08, 2.675857e-08, 2.66382e-08, 2.640722e-08,
  2.324277e-08, 2.312297e-08, 2.293769e-08, 2.407029e-08, 2.652486e-08, 
    2.996676e-08, 2.918e-08, 2.828279e-08, 2.775958e-08, 2.769699e-08, 
    2.710042e-08, 2.670712e-08, 2.69375e-08, 2.671697e-08, 2.675585e-08,
  2.331899e-08, 2.342606e-08, 2.303992e-08, 2.400274e-08, 2.682486e-08, 
    2.943535e-08, 2.95808e-08, 2.831305e-08, 2.774355e-08, 2.669916e-08, 
    2.672361e-08, 2.649889e-08, 2.687386e-08, 2.705871e-08, 2.679512e-08,
  2.339836e-08, 2.359446e-08, 2.352741e-08, 2.443966e-08, 2.679394e-08, 
    2.95408e-08, 2.917012e-08, 2.82056e-08, 2.775431e-08, 2.709224e-08, 
    2.693681e-08, 2.670614e-08, 2.699212e-08, 2.690505e-08, 2.674997e-08,
  2.345667e-08, 2.367745e-08, 2.397925e-08, 2.509987e-08, 2.705493e-08, 
    2.90798e-08, 2.926711e-08, 2.770366e-08, 2.663449e-08, 2.646558e-08, 
    2.672493e-08, 2.660908e-08, 2.693919e-08, 2.728991e-08, 2.69074e-08,
  2.355466e-08, 2.352929e-08, 2.43742e-08, 2.600472e-08, 2.720124e-08, 
    2.863522e-08, 2.85977e-08, 2.752503e-08, 2.742211e-08, 2.738012e-08, 
    2.730611e-08, 2.675797e-08, 2.702065e-08, 2.717089e-08, 2.687184e-08,
  2.362362e-08, 2.317032e-08, 2.420406e-08, 2.675648e-08, 2.772597e-08, 
    2.811787e-08, 2.806195e-08, 2.725027e-08, 2.692056e-08, 2.709605e-08, 
    2.682369e-08, 2.678379e-08, 2.716228e-08, 2.721117e-08, 2.690323e-08,
  2.382441e-08, 2.314546e-08, 2.399527e-08, 2.754993e-08, 2.820364e-08, 
    2.769929e-08, 2.787964e-08, 2.731878e-08, 2.722952e-08, 2.734722e-08, 
    2.736479e-08, 2.724942e-08, 2.711528e-08, 2.679157e-08, 2.680421e-08,
  2.551299e-08, 2.561679e-08, 2.667689e-08, 2.752667e-08, 2.825653e-08, 
    2.878161e-08, 2.903914e-08, 2.874587e-08, 2.801743e-08, 2.741517e-08, 
    2.705454e-08, 2.718694e-08, 2.740292e-08, 2.767731e-08, 2.79335e-08,
  2.543958e-08, 2.591583e-08, 2.672196e-08, 2.754609e-08, 2.841431e-08, 
    2.878718e-08, 2.908082e-08, 2.903237e-08, 2.755504e-08, 2.613022e-08, 
    2.590478e-08, 2.595199e-08, 2.658981e-08, 2.621936e-08, 2.661147e-08,
  2.509823e-08, 2.59656e-08, 2.676405e-08, 2.757618e-08, 2.876893e-08, 
    2.865183e-08, 2.879237e-08, 2.857727e-08, 2.725552e-08, 2.590104e-08, 
    2.617322e-08, 2.628575e-08, 2.640695e-08, 2.631448e-08, 2.629315e-08,
  2.453348e-08, 2.571308e-08, 2.693025e-08, 2.748439e-08, 2.841121e-08, 
    2.897487e-08, 2.872467e-08, 2.854955e-08, 2.6655e-08, 2.577288e-08, 
    2.64392e-08, 2.643849e-08, 2.661448e-08, 2.64212e-08, 2.646272e-08,
  2.431271e-08, 2.525982e-08, 2.68452e-08, 2.76178e-08, 2.815725e-08, 
    2.757029e-08, 2.892102e-08, 2.878394e-08, 2.688295e-08, 2.600771e-08, 
    2.688556e-08, 2.723211e-08, 2.684382e-08, 2.701144e-08, 2.621531e-08,
  2.415091e-08, 2.490799e-08, 2.63236e-08, 2.751222e-08, 2.822791e-08, 
    2.805361e-08, 2.795983e-08, 2.950012e-08, 2.852453e-08, 2.734283e-08, 
    2.721452e-08, 2.767348e-08, 2.676145e-08, 2.715346e-08, 2.702585e-08,
  2.455479e-08, 2.487501e-08, 2.578326e-08, 2.734086e-08, 2.80736e-08, 
    2.756993e-08, 2.808073e-08, 2.787361e-08, 2.772048e-08, 2.763495e-08, 
    2.762418e-08, 2.793421e-08, 2.702063e-08, 2.762221e-08, 2.795059e-08,
  2.474601e-08, 2.530507e-08, 2.540211e-08, 2.661205e-08, 2.812445e-08, 
    2.758755e-08, 2.769995e-08, 2.85641e-08, 2.856521e-08, 2.804172e-08, 
    2.777673e-08, 2.804507e-08, 2.766669e-08, 2.851354e-08, 2.8439e-08,
  2.478946e-08, 2.564451e-08, 2.578661e-08, 2.61935e-08, 2.769727e-08, 
    2.752529e-08, 2.738383e-08, 2.779346e-08, 2.840178e-08, 2.835261e-08, 
    2.793434e-08, 2.817534e-08, 2.805965e-08, 2.852162e-08, 2.83912e-08,
  2.448255e-08, 2.58051e-08, 2.612752e-08, 2.596131e-08, 2.762302e-08, 
    2.761605e-08, 2.705172e-08, 2.756848e-08, 2.819342e-08, 2.859714e-08, 
    2.847787e-08, 2.836127e-08, 2.812295e-08, 2.839312e-08, 2.792248e-08,
  2.520327e-08, 2.619528e-08, 2.745209e-08, 2.67138e-08, 2.498826e-08, 
    2.577339e-08, 2.606277e-08, 2.661686e-08, 2.700375e-08, 2.788384e-08, 
    2.775151e-08, 2.668313e-08, 2.763907e-08, 2.753802e-08, 2.758236e-08,
  2.517127e-08, 2.608862e-08, 2.66802e-08, 2.685555e-08, 2.502896e-08, 
    2.499089e-08, 2.581319e-08, 2.574679e-08, 2.680986e-08, 2.714377e-08, 
    2.813408e-08, 2.733453e-08, 2.724575e-08, 2.802347e-08, 2.777111e-08,
  2.526975e-08, 2.644778e-08, 2.642483e-08, 2.673148e-08, 2.460868e-08, 
    2.434389e-08, 2.538511e-08, 2.50164e-08, 2.547942e-08, 2.665125e-08, 
    2.778482e-08, 2.788451e-08, 2.725761e-08, 2.815877e-08, 2.792244e-08,
  2.499456e-08, 2.656756e-08, 2.644949e-08, 2.621671e-08, 2.446458e-08, 
    2.437681e-08, 2.448354e-08, 2.438814e-08, 2.472244e-08, 2.60439e-08, 
    2.686482e-08, 2.837003e-08, 2.764779e-08, 2.757412e-08, 2.836326e-08,
  2.489327e-08, 2.61885e-08, 2.646216e-08, 2.626608e-08, 2.452914e-08, 
    2.352014e-08, 2.400575e-08, 2.423828e-08, 2.406161e-08, 2.497849e-08, 
    2.61704e-08, 2.779597e-08, 2.811968e-08, 2.787811e-08, 2.790316e-08,
  2.480804e-08, 2.572273e-08, 2.635112e-08, 2.609399e-08, 2.449772e-08, 
    2.373385e-08, 2.306088e-08, 2.403608e-08, 2.405102e-08, 2.406927e-08, 
    2.583555e-08, 2.701911e-08, 2.831011e-08, 2.794752e-08, 2.826506e-08,
  2.455159e-08, 2.507841e-08, 2.582002e-08, 2.598143e-08, 2.438002e-08, 
    2.375143e-08, 2.230939e-08, 2.202158e-08, 2.261229e-08, 2.350375e-08, 
    2.522121e-08, 2.643384e-08, 2.813482e-08, 2.813298e-08, 2.801651e-08,
  2.41289e-08, 2.470287e-08, 2.507725e-08, 2.547586e-08, 2.432463e-08, 
    2.393646e-08, 2.220968e-08, 2.136158e-08, 2.207782e-08, 2.307592e-08, 
    2.50192e-08, 2.609045e-08, 2.763569e-08, 2.804632e-08, 2.782851e-08,
  2.389024e-08, 2.440966e-08, 2.430285e-08, 2.498023e-08, 2.357415e-08, 
    2.370411e-08, 2.179205e-08, 2.055393e-08, 2.148648e-08, 2.284132e-08, 
    2.481269e-08, 2.602638e-08, 2.723798e-08, 2.783058e-08, 2.794186e-08,
  2.373652e-08, 2.413047e-08, 2.40715e-08, 2.419837e-08, 2.297246e-08, 
    2.312427e-08, 2.160689e-08, 2.066941e-08, 2.116222e-08, 2.252324e-08, 
    2.476348e-08, 2.619246e-08, 2.686622e-08, 2.759468e-08, 2.767432e-08,
  2.249316e-08, 2.283925e-08, 2.243122e-08, 2.2206e-08, 2.201486e-08, 
    2.226721e-08, 2.191449e-08, 2.152491e-08, 2.068315e-08, 2.05061e-08, 
    2.110659e-08, 2.225767e-08, 2.400093e-08, 2.474255e-08, 2.562891e-08,
  2.324091e-08, 2.311933e-08, 2.263447e-08, 2.234228e-08, 2.200085e-08, 
    2.206159e-08, 2.210879e-08, 2.141299e-08, 2.063565e-08, 2.100518e-08, 
    2.139632e-08, 2.255788e-08, 2.418238e-08, 2.486338e-08, 2.536624e-08,
  2.367456e-08, 2.356541e-08, 2.306822e-08, 2.253178e-08, 2.205889e-08, 
    2.188107e-08, 2.143408e-08, 2.124682e-08, 2.108215e-08, 2.166139e-08, 
    2.211771e-08, 2.2867e-08, 2.392586e-08, 2.521068e-08, 2.556465e-08,
  2.379566e-08, 2.405988e-08, 2.371302e-08, 2.303311e-08, 2.251336e-08, 
    2.209361e-08, 2.088931e-08, 2.112767e-08, 2.147745e-08, 2.233507e-08, 
    2.270929e-08, 2.327936e-08, 2.45443e-08, 2.549439e-08, 2.551096e-08,
  2.396215e-08, 2.44051e-08, 2.439733e-08, 2.362353e-08, 2.26335e-08, 
    2.185468e-08, 2.166309e-08, 2.081215e-08, 2.147462e-08, 2.348334e-08, 
    2.341134e-08, 2.387062e-08, 2.502533e-08, 2.574573e-08, 2.574081e-08,
  2.420237e-08, 2.46119e-08, 2.491636e-08, 2.428099e-08, 2.316727e-08, 
    2.270212e-08, 2.184354e-08, 2.253615e-08, 2.280325e-08, 2.370583e-08, 
    2.380582e-08, 2.461525e-08, 2.550779e-08, 2.580902e-08, 2.567304e-08,
  2.447232e-08, 2.475224e-08, 2.51881e-08, 2.472634e-08, 2.367575e-08, 
    2.28845e-08, 2.300488e-08, 2.213629e-08, 2.241633e-08, 2.446909e-08, 
    2.461228e-08, 2.510063e-08, 2.554378e-08, 2.568751e-08, 2.559391e-08,
  2.468991e-08, 2.476117e-08, 2.526582e-08, 2.506614e-08, 2.423019e-08, 
    2.345219e-08, 2.318574e-08, 2.294034e-08, 2.308927e-08, 2.508056e-08, 
    2.503832e-08, 2.557807e-08, 2.572349e-08, 2.576553e-08, 2.553751e-08,
  2.476843e-08, 2.491882e-08, 2.538354e-08, 2.53681e-08, 2.453853e-08, 
    2.375902e-08, 2.37913e-08, 2.328085e-08, 2.328455e-08, 2.499959e-08, 
    2.54436e-08, 2.589388e-08, 2.566866e-08, 2.567627e-08, 2.531634e-08,
  2.471432e-08, 2.500685e-08, 2.534338e-08, 2.538044e-08, 2.475793e-08, 
    2.416129e-08, 2.400295e-08, 2.365094e-08, 2.347288e-08, 2.504358e-08, 
    2.573181e-08, 2.611281e-08, 2.569197e-08, 2.569453e-08, 2.518498e-08,
  2.247443e-08, 2.341913e-08, 2.431577e-08, 2.448741e-08, 2.476976e-08, 
    2.469245e-08, 2.476717e-08, 2.513981e-08, 2.490757e-08, 2.54622e-08, 
    2.571552e-08, 2.56821e-08, 2.602706e-08, 2.56462e-08, 2.50592e-08,
  2.205134e-08, 2.292853e-08, 2.400593e-08, 2.434744e-08, 2.475666e-08, 
    2.517517e-08, 2.498382e-08, 2.522904e-08, 2.508056e-08, 2.542337e-08, 
    2.571601e-08, 2.59201e-08, 2.629336e-08, 2.564465e-08, 2.553288e-08,
  2.155319e-08, 2.224606e-08, 2.347143e-08, 2.398999e-08, 2.424962e-08, 
    2.492855e-08, 2.513974e-08, 2.52909e-08, 2.500189e-08, 2.530391e-08, 
    2.559907e-08, 2.600823e-08, 2.604944e-08, 2.606055e-08, 2.635637e-08,
  2.144494e-08, 2.169417e-08, 2.287583e-08, 2.385419e-08, 2.405521e-08, 
    2.491282e-08, 2.520227e-08, 2.548125e-08, 2.505791e-08, 2.517551e-08, 
    2.538292e-08, 2.592041e-08, 2.600762e-08, 2.612951e-08, 2.580228e-08,
  2.133673e-08, 2.143208e-08, 2.211549e-08, 2.34363e-08, 2.361052e-08, 
    2.383347e-08, 2.503141e-08, 2.461402e-08, 2.437407e-08, 2.516646e-08, 
    2.499315e-08, 2.564909e-08, 2.587459e-08, 2.585985e-08, 2.590444e-08,
  2.156716e-08, 2.139111e-08, 2.163702e-08, 2.294525e-08, 2.356789e-08, 
    2.409852e-08, 2.446004e-08, 2.525525e-08, 2.499786e-08, 2.509741e-08, 
    2.48166e-08, 2.532783e-08, 2.589087e-08, 2.582249e-08, 2.576468e-08,
  2.18562e-08, 2.153348e-08, 2.143079e-08, 2.255624e-08, 2.315594e-08, 
    2.339213e-08, 2.471457e-08, 2.459684e-08, 2.430106e-08, 2.498433e-08, 
    2.476751e-08, 2.506766e-08, 2.578689e-08, 2.586382e-08, 2.563633e-08,
  2.214342e-08, 2.173824e-08, 2.137232e-08, 2.231246e-08, 2.302708e-08, 
    2.330543e-08, 2.427828e-08, 2.481795e-08, 2.423338e-08, 2.472706e-08, 
    2.480764e-08, 2.501172e-08, 2.564338e-08, 2.582853e-08, 2.566975e-08,
  2.24593e-08, 2.18443e-08, 2.144171e-08, 2.216653e-08, 2.280865e-08, 
    2.29967e-08, 2.412642e-08, 2.452107e-08, 2.402168e-08, 2.442952e-08, 
    2.470513e-08, 2.498354e-08, 2.564249e-08, 2.581706e-08, 2.556247e-08,
  2.281081e-08, 2.187103e-08, 2.152319e-08, 2.207216e-08, 2.272292e-08, 
    2.310786e-08, 2.361092e-08, 2.447631e-08, 2.398374e-08, 2.414041e-08, 
    2.458852e-08, 2.522506e-08, 2.553696e-08, 2.579411e-08, 2.565647e-08,
  2.429006e-08, 2.341383e-08, 2.268305e-08, 2.238878e-08, 2.220795e-08, 
    2.252185e-08, 2.279256e-08, 2.349557e-08, 2.336445e-08, 2.347355e-08, 
    2.372684e-08, 2.451494e-08, 2.524222e-08, 2.570633e-08, 2.565571e-08,
  2.467381e-08, 2.347686e-08, 2.288156e-08, 2.268883e-08, 2.231218e-08, 
    2.246908e-08, 2.296724e-08, 2.326156e-08, 2.333336e-08, 2.343535e-08, 
    2.358464e-08, 2.413319e-08, 2.488204e-08, 2.548784e-08, 2.568866e-08,
  2.468858e-08, 2.364734e-08, 2.297082e-08, 2.282621e-08, 2.244368e-08, 
    2.233378e-08, 2.32074e-08, 2.326843e-08, 2.33796e-08, 2.35112e-08, 
    2.339472e-08, 2.389698e-08, 2.440104e-08, 2.573657e-08, 2.586547e-08,
  2.504698e-08, 2.415005e-08, 2.319304e-08, 2.292562e-08, 2.285514e-08, 
    2.265425e-08, 2.27024e-08, 2.375712e-08, 2.369197e-08, 2.377501e-08, 
    2.349848e-08, 2.369897e-08, 2.404098e-08, 2.460848e-08, 2.516703e-08,
  2.542281e-08, 2.434496e-08, 2.346331e-08, 2.299414e-08, 2.303696e-08, 
    2.275071e-08, 2.307994e-08, 2.272494e-08, 2.29147e-08, 2.409855e-08, 
    2.368236e-08, 2.372019e-08, 2.390449e-08, 2.471445e-08, 2.524075e-08,
  2.599223e-08, 2.466093e-08, 2.386509e-08, 2.315176e-08, 2.321771e-08, 
    2.322745e-08, 2.347619e-08, 2.373188e-08, 2.33602e-08, 2.353262e-08, 
    2.354624e-08, 2.374559e-08, 2.381503e-08, 2.430113e-08, 2.481192e-08,
  2.64936e-08, 2.476492e-08, 2.413454e-08, 2.341792e-08, 2.329646e-08, 
    2.327631e-08, 2.365404e-08, 2.371909e-08, 2.309966e-08, 2.349405e-08, 
    2.340826e-08, 2.367763e-08, 2.382161e-08, 2.443648e-08, 2.477245e-08,
  2.677508e-08, 2.500289e-08, 2.430051e-08, 2.359126e-08, 2.346206e-08, 
    2.355217e-08, 2.36845e-08, 2.404603e-08, 2.351491e-08, 2.327439e-08, 
    2.309069e-08, 2.345962e-08, 2.377238e-08, 2.447136e-08, 2.46546e-08,
  2.682212e-08, 2.506213e-08, 2.438032e-08, 2.374027e-08, 2.358015e-08, 
    2.359584e-08, 2.380223e-08, 2.390408e-08, 2.346051e-08, 2.33327e-08, 
    2.303759e-08, 2.328581e-08, 2.379152e-08, 2.449806e-08, 2.481515e-08,
  2.69305e-08, 2.537154e-08, 2.436635e-08, 2.376738e-08, 2.362292e-08, 
    2.387927e-08, 2.388074e-08, 2.401907e-08, 2.36744e-08, 2.296209e-08, 
    2.271086e-08, 2.339018e-08, 2.377192e-08, 2.451838e-08, 2.517046e-08,
  2.440014e-08, 2.506947e-08, 2.473695e-08, 2.394572e-08, 2.456354e-08, 
    2.404172e-08, 2.411996e-08, 2.39529e-08, 2.426358e-08, 2.442654e-08, 
    2.441787e-08, 2.380365e-08, 2.353133e-08, 2.354175e-08, 2.40095e-08,
  2.4509e-08, 2.539069e-08, 2.564424e-08, 2.431969e-08, 2.456786e-08, 
    2.424924e-08, 2.426615e-08, 2.39229e-08, 2.440258e-08, 2.442852e-08, 
    2.452344e-08, 2.416224e-08, 2.3649e-08, 2.309826e-08, 2.369483e-08,
  2.420166e-08, 2.495549e-08, 2.643352e-08, 2.467039e-08, 2.465305e-08, 
    2.436704e-08, 2.436275e-08, 2.412893e-08, 2.437724e-08, 2.430049e-08, 
    2.475191e-08, 2.444053e-08, 2.388003e-08, 2.338195e-08, 2.37059e-08,
  2.399947e-08, 2.45932e-08, 2.68067e-08, 2.498656e-08, 2.452878e-08, 
    2.455235e-08, 2.420896e-08, 2.424261e-08, 2.461513e-08, 2.413922e-08, 
    2.460204e-08, 2.427658e-08, 2.412689e-08, 2.345464e-08, 2.350654e-08,
  2.345852e-08, 2.439815e-08, 2.707562e-08, 2.52405e-08, 2.457726e-08, 
    2.428922e-08, 2.410929e-08, 2.382946e-08, 2.438516e-08, 2.455061e-08, 
    2.448713e-08, 2.446642e-08, 2.403764e-08, 2.405693e-08, 2.3732e-08,
  2.347453e-08, 2.45601e-08, 2.703201e-08, 2.528798e-08, 2.451231e-08, 
    2.463692e-08, 2.4297e-08, 2.447103e-08, 2.459908e-08, 2.460722e-08, 
    2.450644e-08, 2.428059e-08, 2.432095e-08, 2.4337e-08, 2.414031e-08,
  2.350567e-08, 2.464861e-08, 2.652379e-08, 2.522511e-08, 2.468931e-08, 
    2.442031e-08, 2.434548e-08, 2.442414e-08, 2.449665e-08, 2.449369e-08, 
    2.485125e-08, 2.511277e-08, 2.503205e-08, 2.494981e-08, 2.465669e-08,
  2.346777e-08, 2.479343e-08, 2.627121e-08, 2.513667e-08, 2.47338e-08, 
    2.467487e-08, 2.464725e-08, 2.496292e-08, 2.532797e-08, 2.571353e-08, 
    2.579741e-08, 2.611209e-08, 2.575278e-08, 2.569918e-08, 2.504014e-08,
  2.367865e-08, 2.506532e-08, 2.587911e-08, 2.499278e-08, 2.486426e-08, 
    2.463839e-08, 2.485374e-08, 2.528551e-08, 2.56655e-08, 2.601149e-08, 
    2.613132e-08, 2.681883e-08, 2.692095e-08, 2.648829e-08, 2.620439e-08,
  2.418708e-08, 2.52878e-08, 2.571242e-08, 2.499717e-08, 2.490598e-08, 
    2.479894e-08, 2.526915e-08, 2.567335e-08, 2.629863e-08, 2.644474e-08, 
    2.71861e-08, 2.770972e-08, 2.760157e-08, 2.750931e-08, 2.6969e-08,
  2.536505e-08, 2.44964e-08, 2.475156e-08, 2.539551e-08, 2.567627e-08, 
    2.59503e-08, 2.623392e-08, 2.591444e-08, 2.562394e-08, 2.571946e-08, 
    2.543628e-08, 2.528526e-08, 2.484644e-08, 2.469678e-08, 2.445871e-08,
  2.52536e-08, 2.493337e-08, 2.495925e-08, 2.552039e-08, 2.586688e-08, 
    2.60451e-08, 2.635105e-08, 2.594314e-08, 2.607059e-08, 2.584175e-08, 
    2.580291e-08, 2.547847e-08, 2.529416e-08, 2.47993e-08, 2.396965e-08,
  2.512466e-08, 2.497978e-08, 2.496706e-08, 2.556907e-08, 2.596724e-08, 
    2.624232e-08, 2.641401e-08, 2.621568e-08, 2.663061e-08, 2.628256e-08, 
    2.6446e-08, 2.610146e-08, 2.581097e-08, 2.515118e-08, 2.430973e-08,
  2.502004e-08, 2.540678e-08, 2.529874e-08, 2.580999e-08, 2.631203e-08, 
    2.656715e-08, 2.662937e-08, 2.655322e-08, 2.720656e-08, 2.69e-08, 
    2.708328e-08, 2.666282e-08, 2.649202e-08, 2.549591e-08, 2.518618e-08,
  2.494463e-08, 2.559362e-08, 2.544388e-08, 2.587046e-08, 2.647197e-08, 
    2.666915e-08, 2.674785e-08, 2.675166e-08, 2.749264e-08, 2.776854e-08, 
    2.789131e-08, 2.795511e-08, 2.74831e-08, 2.635485e-08, 2.590438e-08,
  2.498356e-08, 2.591379e-08, 2.581381e-08, 2.606978e-08, 2.673357e-08, 
    2.707186e-08, 2.704479e-08, 2.753797e-08, 2.817657e-08, 2.83268e-08, 
    2.861163e-08, 2.817662e-08, 2.81345e-08, 2.716626e-08, 2.635434e-08,
  2.50504e-08, 2.609844e-08, 2.591751e-08, 2.613722e-08, 2.681662e-08, 
    2.725577e-08, 2.767503e-08, 2.777131e-08, 2.788851e-08, 2.799883e-08, 
    2.822935e-08, 2.805301e-08, 2.818359e-08, 2.780024e-08, 2.681656e-08,
  2.517832e-08, 2.62147e-08, 2.621336e-08, 2.627216e-08, 2.690021e-08, 
    2.755643e-08, 2.781464e-08, 2.819727e-08, 2.840973e-08, 2.825318e-08, 
    2.83569e-08, 2.810282e-08, 2.875544e-08, 2.837561e-08, 2.749265e-08,
  2.54062e-08, 2.625467e-08, 2.635207e-08, 2.632992e-08, 2.706193e-08, 
    2.778866e-08, 2.811289e-08, 2.814039e-08, 2.835844e-08, 2.757686e-08, 
    2.739817e-08, 2.728748e-08, 2.830452e-08, 2.860596e-08, 2.788457e-08,
  2.568554e-08, 2.626517e-08, 2.642949e-08, 2.638445e-08, 2.706095e-08, 
    2.801247e-08, 2.805047e-08, 2.822435e-08, 2.803582e-08, 2.721172e-08, 
    2.778017e-08, 2.76625e-08, 2.824845e-08, 2.859074e-08, 2.799259e-08,
  2.621034e-08, 2.54033e-08, 2.617157e-08, 2.689826e-08, 2.666695e-08, 
    2.726716e-08, 2.751245e-08, 2.774308e-08, 2.758585e-08, 2.764948e-08, 
    2.738584e-08, 2.731804e-08, 2.702933e-08, 2.638645e-08, 2.569293e-08,
  2.628369e-08, 2.574966e-08, 2.646892e-08, 2.719452e-08, 2.700887e-08, 
    2.75753e-08, 2.809395e-08, 2.81065e-08, 2.807693e-08, 2.793371e-08, 
    2.785761e-08, 2.740387e-08, 2.754136e-08, 2.664888e-08, 2.549806e-08,
  2.628579e-08, 2.602119e-08, 2.671918e-08, 2.744991e-08, 2.70653e-08, 
    2.772487e-08, 2.832036e-08, 2.825462e-08, 2.835288e-08, 2.805671e-08, 
    2.828924e-08, 2.759914e-08, 2.777094e-08, 2.734106e-08, 2.550868e-08,
  2.636613e-08, 2.631122e-08, 2.69887e-08, 2.758091e-08, 2.735263e-08, 
    2.804607e-08, 2.83535e-08, 2.832455e-08, 2.916351e-08, 2.862991e-08, 
    2.850459e-08, 2.819866e-08, 2.782598e-08, 2.783369e-08, 2.615227e-08,
  2.646656e-08, 2.644844e-08, 2.706392e-08, 2.754527e-08, 2.749932e-08, 
    2.811192e-08, 2.86052e-08, 2.82506e-08, 2.851075e-08, 2.781302e-08, 
    2.825388e-08, 2.810419e-08, 2.80995e-08, 2.798331e-08, 2.668601e-08,
  2.674753e-08, 2.651037e-08, 2.707919e-08, 2.75204e-08, 2.779906e-08, 
    2.856277e-08, 2.884682e-08, 2.883809e-08, 2.898727e-08, 2.840272e-08, 
    2.857312e-08, 2.855134e-08, 2.819674e-08, 2.820673e-08, 2.717279e-08,
  2.681951e-08, 2.635764e-08, 2.707342e-08, 2.754089e-08, 2.795878e-08, 
    2.87684e-08, 2.901825e-08, 2.847828e-08, 2.854911e-08, 2.760102e-08, 
    2.764237e-08, 2.845539e-08, 2.833007e-08, 2.818878e-08, 2.742981e-08,
  2.679812e-08, 2.635139e-08, 2.724948e-08, 2.737301e-08, 2.796361e-08, 
    2.86708e-08, 2.84673e-08, 2.847405e-08, 2.872271e-08, 2.854214e-08, 
    2.810742e-08, 2.859737e-08, 2.82357e-08, 2.809371e-08, 2.762269e-08,
  2.642561e-08, 2.625316e-08, 2.72622e-08, 2.761874e-08, 2.834732e-08, 
    2.861019e-08, 2.829381e-08, 2.828865e-08, 2.83632e-08, 2.81548e-08, 
    2.763573e-08, 2.826314e-08, 2.832985e-08, 2.810071e-08, 2.762451e-08,
  2.6807e-08, 2.626835e-08, 2.706265e-08, 2.738391e-08, 2.78956e-08, 
    2.828203e-08, 2.770958e-08, 2.755863e-08, 2.751974e-08, 2.772012e-08, 
    2.829263e-08, 2.841554e-08, 2.817694e-08, 2.810705e-08, 2.737223e-08,
  2.772224e-08, 2.735007e-08, 2.689752e-08, 2.667288e-08, 2.659838e-08, 
    2.678673e-08, 2.680262e-08, 2.692663e-08, 2.698184e-08, 2.731603e-08, 
    2.75448e-08, 2.775776e-08, 2.754658e-08, 2.718122e-08, 2.670164e-08,
  2.785893e-08, 2.716708e-08, 2.681187e-08, 2.695523e-08, 2.706321e-08, 
    2.717968e-08, 2.738006e-08, 2.755236e-08, 2.753465e-08, 2.769607e-08, 
    2.762738e-08, 2.79941e-08, 2.765512e-08, 2.752212e-08, 2.686804e-08,
  2.712673e-08, 2.668258e-08, 2.662254e-08, 2.714902e-08, 2.716676e-08, 
    2.769069e-08, 2.78831e-08, 2.813318e-08, 2.789791e-08, 2.818463e-08, 
    2.774354e-08, 2.805014e-08, 2.787219e-08, 2.738571e-08, 2.67927e-08,
  2.686828e-08, 2.686494e-08, 2.702741e-08, 2.753669e-08, 2.7657e-08, 
    2.822647e-08, 2.786484e-08, 2.83541e-08, 2.767021e-08, 2.829412e-08, 
    2.818866e-08, 2.83584e-08, 2.793721e-08, 2.754488e-08, 2.685649e-08,
  2.65278e-08, 2.679456e-08, 2.741718e-08, 2.768083e-08, 2.796522e-08, 
    2.763174e-08, 2.860024e-08, 2.8491e-08, 2.820397e-08, 2.783484e-08, 
    2.837948e-08, 2.839874e-08, 2.780711e-08, 2.753651e-08, 2.690572e-08,
  2.612607e-08, 2.691221e-08, 2.783922e-08, 2.784519e-08, 2.772117e-08, 
    2.823533e-08, 2.699185e-08, 2.478809e-08, 2.831943e-08, 2.926767e-08, 
    2.912354e-08, 2.882604e-08, 2.787784e-08, 2.751196e-08, 2.683129e-08,
  2.637733e-08, 2.69781e-08, 2.814545e-08, 2.80482e-08, 2.790407e-08, 
    2.825569e-08, 2.822413e-08, 2.84605e-08, 2.94797e-08, 3.025436e-08, 
    2.933569e-08, 2.874976e-08, 2.767195e-08, 2.75532e-08, 2.668348e-08,
  2.646772e-08, 2.696842e-08, 2.831119e-08, 2.822164e-08, 2.79088e-08, 
    2.834966e-08, 2.900482e-08, 2.909396e-08, 2.956689e-08, 3.024208e-08, 
    2.906216e-08, 2.830861e-08, 2.776773e-08, 2.755506e-08, 2.638582e-08,
  2.685723e-08, 2.666549e-08, 2.809147e-08, 2.845427e-08, 2.805109e-08, 
    2.788511e-08, 2.89986e-08, 2.882993e-08, 2.973188e-08, 2.928961e-08, 
    2.845263e-08, 2.830862e-08, 2.759874e-08, 2.737596e-08, 2.610693e-08,
  2.731792e-08, 2.666135e-08, 2.755739e-08, 2.843401e-08, 2.836243e-08, 
    2.793319e-08, 2.809969e-08, 2.847166e-08, 2.88056e-08, 2.834726e-08, 
    2.880252e-08, 2.802734e-08, 2.754377e-08, 2.723486e-08, 2.579706e-08,
  2.761031e-08, 2.774212e-08, 2.830704e-08, 2.856136e-08, 2.809332e-08, 
    2.788156e-08, 2.779421e-08, 2.802797e-08, 2.798205e-08, 2.735363e-08, 
    2.711703e-08, 2.706548e-08, 2.755976e-08, 2.792837e-08, 2.836169e-08,
  2.757753e-08, 2.820064e-08, 2.886794e-08, 2.860147e-08, 2.799693e-08, 
    2.737485e-08, 2.777754e-08, 2.813833e-08, 2.831971e-08, 2.751396e-08, 
    2.694408e-08, 2.676204e-08, 2.721479e-08, 2.825577e-08, 2.838446e-08,
  2.761e-08, 2.831092e-08, 2.871734e-08, 2.843261e-08, 2.782347e-08, 
    2.704697e-08, 2.822399e-08, 2.832691e-08, 2.868862e-08, 2.76441e-08, 
    2.668859e-08, 2.657806e-08, 2.699638e-08, 2.76523e-08, 2.813685e-08,
  2.769866e-08, 2.849731e-08, 2.905417e-08, 2.870796e-08, 2.780556e-08, 
    2.778414e-08, 2.641416e-08, 2.837933e-08, 2.818768e-08, 2.766516e-08, 
    2.671827e-08, 2.643025e-08, 2.712241e-08, 2.759929e-08, 2.781748e-08,
  2.762585e-08, 2.842025e-08, 2.892523e-08, 2.893138e-08, 2.778841e-08, 
    2.690909e-08, 2.787769e-08, 2.925653e-08, 2.833329e-08, 2.729942e-08, 
    2.658949e-08, 2.668858e-08, 2.721121e-08, 2.761064e-08, 2.789736e-08,
  2.768593e-08, 2.85314e-08, 2.912932e-08, 2.936463e-08, 2.884825e-08, 
    2.650723e-08, 2.665649e-08, 2.663887e-08, 2.687768e-08, 2.757502e-08, 
    2.663584e-08, 2.669894e-08, 2.739789e-08, 2.758187e-08, 2.770613e-08,
  2.756403e-08, 2.823572e-08, 2.899093e-08, 2.936132e-08, 2.986988e-08, 
    2.85622e-08, 2.703208e-08, 2.809474e-08, 2.795625e-08, 2.727625e-08, 
    2.653072e-08, 2.722307e-08, 2.760369e-08, 2.761001e-08, 2.764047e-08,
  2.750884e-08, 2.812565e-08, 2.892807e-08, 2.919708e-08, 2.971875e-08, 
    2.993093e-08, 2.859878e-08, 2.860159e-08, 2.789065e-08, 2.752797e-08, 
    2.713754e-08, 2.745923e-08, 2.761527e-08, 2.763705e-08, 2.757391e-08,
  2.732436e-08, 2.773051e-08, 2.872763e-08, 2.909514e-08, 2.945506e-08, 
    2.992633e-08, 3.00364e-08, 2.890285e-08, 2.901185e-08, 2.780712e-08, 
    2.738089e-08, 2.794122e-08, 2.778126e-08, 2.759813e-08, 2.728333e-08,
  2.716725e-08, 2.744924e-08, 2.822917e-08, 2.881769e-08, 2.906838e-08, 
    2.92602e-08, 2.950149e-08, 2.910419e-08, 2.862763e-08, 2.743106e-08, 
    2.790117e-08, 2.803457e-08, 2.760459e-08, 2.7458e-08, 2.701795e-08,
  2.757308e-08, 2.810201e-08, 2.930495e-08, 2.966698e-08, 2.858552e-08, 
    2.762469e-08, 2.7631e-08, 2.814707e-08, 2.881805e-08, 2.889223e-08, 
    2.894567e-08, 2.839576e-08, 2.827496e-08, 2.741539e-08, 2.673177e-08,
  2.786209e-08, 2.859223e-08, 2.943581e-08, 2.913281e-08, 2.850888e-08, 
    2.68426e-08, 2.76285e-08, 2.798848e-08, 2.811827e-08, 2.813643e-08, 
    2.854346e-08, 2.849852e-08, 2.841748e-08, 2.787271e-08, 2.722883e-08,
  2.790975e-08, 2.864662e-08, 2.922405e-08, 2.899143e-08, 2.808003e-08, 
    2.728148e-08, 2.773566e-08, 2.794159e-08, 2.855236e-08, 2.860132e-08, 
    2.847131e-08, 2.831984e-08, 2.78498e-08, 2.691256e-08, 2.644179e-08,
  2.792583e-08, 2.86442e-08, 2.895971e-08, 2.856409e-08, 2.817609e-08, 
    2.829943e-08, 2.795999e-08, 2.921392e-08, 2.817756e-08, 2.789939e-08, 
    2.793266e-08, 2.814957e-08, 2.766951e-08, 2.696332e-08, 2.638469e-08,
  2.790712e-08, 2.845208e-08, 2.87124e-08, 2.83157e-08, 2.800332e-08, 
    2.867121e-08, 2.876625e-08, 2.914489e-08, 2.796998e-08, 2.822526e-08, 
    2.7976e-08, 2.74484e-08, 2.740858e-08, 2.715179e-08, 2.650276e-08,
  2.792951e-08, 2.825261e-08, 2.850118e-08, 2.802326e-08, 2.757531e-08, 
    2.795331e-08, 2.838764e-08, 2.808503e-08, 2.83183e-08, 2.814032e-08, 
    2.758566e-08, 2.726246e-08, 2.753637e-08, 2.77399e-08, 2.75083e-08,
  2.78688e-08, 2.803041e-08, 2.827078e-08, 2.79144e-08, 2.740015e-08, 
    2.761613e-08, 2.769951e-08, 2.809178e-08, 2.794581e-08, 2.787319e-08, 
    2.750034e-08, 2.731832e-08, 2.752062e-08, 2.777396e-08, 2.762052e-08,
  2.771411e-08, 2.783506e-08, 2.810783e-08, 2.774817e-08, 2.71155e-08, 
    2.695427e-08, 2.73431e-08, 2.722279e-08, 2.727465e-08, 2.727414e-08, 
    2.739662e-08, 2.764342e-08, 2.772054e-08, 2.789976e-08, 2.804912e-08,
  2.724392e-08, 2.762453e-08, 2.78636e-08, 2.806274e-08, 2.714118e-08, 
    2.668033e-08, 2.661783e-08, 2.675471e-08, 2.676588e-08, 2.690567e-08, 
    2.726414e-08, 2.766622e-08, 2.785835e-08, 2.816461e-08, 2.818796e-08,
  2.66093e-08, 2.745552e-08, 2.758683e-08, 2.815387e-08, 2.775757e-08, 
    2.697047e-08, 2.661253e-08, 2.661823e-08, 2.680937e-08, 2.70755e-08, 
    2.754467e-08, 2.794128e-08, 2.826468e-08, 2.852286e-08, 2.858129e-08,
  2.771167e-08, 2.745369e-08, 2.741929e-08, 2.820437e-08, 2.90785e-08, 
    2.872379e-08, 2.813515e-08, 2.843046e-08, 2.892612e-08, 2.770023e-08, 
    2.776333e-08, 2.714028e-08, 2.741438e-08, 2.688031e-08, 2.780072e-08,
  2.768969e-08, 2.763204e-08, 2.744748e-08, 2.827522e-08, 2.90755e-08, 
    2.871615e-08, 2.819215e-08, 2.789536e-08, 2.821382e-08, 2.785308e-08, 
    2.733769e-08, 2.669574e-08, 2.625519e-08, 2.561391e-08, 2.604213e-08,
  2.725373e-08, 2.753899e-08, 2.744014e-08, 2.796278e-08, 2.904097e-08, 
    2.889076e-08, 2.768684e-08, 2.814312e-08, 2.828586e-08, 2.730869e-08, 
    2.789092e-08, 2.711485e-08, 2.710948e-08, 2.689306e-08, 2.594236e-08,
  2.714428e-08, 2.758368e-08, 2.750371e-08, 2.766683e-08, 2.871509e-08, 
    2.825528e-08, 2.751661e-08, 2.780016e-08, 2.835968e-08, 2.750546e-08, 
    2.701346e-08, 2.690869e-08, 2.589878e-08, 2.582622e-08, 2.514864e-08,
  2.650594e-08, 2.749342e-08, 2.762411e-08, 2.755078e-08, 2.791534e-08, 
    2.823163e-08, 2.83003e-08, 2.800393e-08, 2.617381e-08, 2.650339e-08, 
    2.536937e-08, 2.434349e-08, 2.372246e-08, 2.360938e-08, 2.322089e-08,
  2.61769e-08, 2.708932e-08, 2.772105e-08, 2.768538e-08, 2.779524e-08, 
    2.793451e-08, 2.779332e-08, 2.808311e-08, 2.670637e-08, 2.608326e-08, 
    2.453096e-08, 2.294406e-08, 2.256192e-08, 2.193574e-08, 2.144868e-08,
  2.544317e-08, 2.657556e-08, 2.759932e-08, 2.788834e-08, 2.775303e-08, 
    2.789388e-08, 2.784088e-08, 2.815026e-08, 2.781887e-08, 2.621349e-08, 
    2.451738e-08, 2.32273e-08, 2.301584e-08, 2.26561e-08, 2.273115e-08,
  2.486839e-08, 2.587775e-08, 2.719213e-08, 2.798586e-08, 2.79708e-08, 
    2.792048e-08, 2.761661e-08, 2.779926e-08, 2.796346e-08, 2.670527e-08, 
    2.534853e-08, 2.437619e-08, 2.403498e-08, 2.368801e-08, 2.376416e-08,
  2.433172e-08, 2.51515e-08, 2.645763e-08, 2.767037e-08, 2.807002e-08, 
    2.810996e-08, 2.785737e-08, 2.741314e-08, 2.755962e-08, 2.685401e-08, 
    2.600356e-08, 2.536806e-08, 2.454935e-08, 2.435022e-08, 2.486778e-08,
  2.421904e-08, 2.442976e-08, 2.563492e-08, 2.719826e-08, 2.81151e-08, 
    2.828618e-08, 2.845007e-08, 2.749064e-08, 2.773636e-08, 2.750333e-08, 
    2.685107e-08, 2.598595e-08, 2.550289e-08, 2.570527e-08, 2.586265e-08,
  2.442054e-08, 2.534449e-08, 2.718586e-08, 2.866238e-08, 2.9188e-08, 
    2.816266e-08, 2.633107e-08, 2.460951e-08, 2.393378e-08, 2.396253e-08, 
    2.500687e-08, 2.601353e-08, 2.648308e-08, 2.74197e-08, 2.89764e-08,
  2.431758e-08, 2.512106e-08, 2.699458e-08, 2.850066e-08, 2.897101e-08, 
    2.784428e-08, 2.612764e-08, 2.481238e-08, 2.331402e-08, 2.372512e-08, 
    2.44169e-08, 2.534247e-08, 2.593806e-08, 2.645454e-08, 2.833828e-08,
  2.422723e-08, 2.470161e-08, 2.664713e-08, 2.819483e-08, 2.881503e-08, 
    2.810404e-08, 2.529588e-08, 2.397042e-08, 2.288e-08, 2.326496e-08, 
    2.396371e-08, 2.491531e-08, 2.572982e-08, 2.658687e-08, 2.805422e-08,
  2.423332e-08, 2.442433e-08, 2.619516e-08, 2.772307e-08, 2.88385e-08, 
    2.758138e-08, 2.743568e-08, 2.380425e-08, 2.23574e-08, 2.282977e-08, 
    2.360787e-08, 2.423598e-08, 2.459242e-08, 2.491526e-08, 2.589318e-08,
  2.434521e-08, 2.418818e-08, 2.568726e-08, 2.736912e-08, 2.886772e-08, 
    2.813493e-08, 2.772765e-08, 2.5945e-08, 2.205515e-08, 2.216926e-08, 
    2.351741e-08, 2.42895e-08, 2.498602e-08, 2.531577e-08, 2.575715e-08,
  2.451305e-08, 2.404934e-08, 2.507503e-08, 2.671708e-08, 2.866475e-08, 
    2.881306e-08, 2.781386e-08, 2.555613e-08, 2.238741e-08, 2.235239e-08, 
    2.348106e-08, 2.481061e-08, 2.50371e-08, 2.466383e-08, 2.448647e-08,
  2.474945e-08, 2.399497e-08, 2.464459e-08, 2.600532e-08, 2.834508e-08, 
    2.88644e-08, 2.851159e-08, 2.752428e-08, 2.396599e-08, 2.242808e-08, 
    2.345773e-08, 2.510787e-08, 2.627923e-08, 2.584828e-08, 2.474103e-08,
  2.510204e-08, 2.412296e-08, 2.43372e-08, 2.518801e-08, 2.789097e-08, 
    2.880287e-08, 2.848016e-08, 2.731246e-08, 2.571863e-08, 2.301386e-08, 
    2.341814e-08, 2.465967e-08, 2.639941e-08, 2.706078e-08, 2.621004e-08,
  2.545187e-08, 2.437895e-08, 2.421791e-08, 2.444015e-08, 2.70956e-08, 
    2.862397e-08, 2.895623e-08, 2.717921e-08, 2.74268e-08, 2.439971e-08, 
    2.410629e-08, 2.456993e-08, 2.602486e-08, 2.730192e-08, 2.770224e-08,
  2.583983e-08, 2.458603e-08, 2.42731e-08, 2.392038e-08, 2.620584e-08, 
    2.822914e-08, 2.913865e-08, 2.748316e-08, 2.700107e-08, 2.614501e-08, 
    2.497944e-08, 2.481458e-08, 2.554905e-08, 2.654194e-08, 2.696787e-08,
  2.616531e-08, 2.597086e-08, 2.550336e-08, 2.50161e-08, 2.557608e-08, 
    2.64617e-08, 2.759975e-08, 2.831865e-08, 2.575177e-08, 2.45882e-08, 
    2.601642e-08, 2.619118e-08, 2.547884e-08, 2.808389e-08, 2.961943e-08,
  2.627303e-08, 2.609396e-08, 2.532986e-08, 2.494055e-08, 2.547576e-08, 
    2.680655e-08, 2.843689e-08, 2.896694e-08, 2.575221e-08, 2.43793e-08, 
    2.613673e-08, 2.648832e-08, 2.514015e-08, 2.673403e-08, 3.002765e-08,
  2.640203e-08, 2.605037e-08, 2.520768e-08, 2.486425e-08, 2.542019e-08, 
    2.762515e-08, 2.859207e-08, 2.870929e-08, 2.553704e-08, 2.428506e-08, 
    2.603226e-08, 2.686384e-08, 2.541095e-08, 2.533202e-08, 2.925096e-08,
  2.656534e-08, 2.635674e-08, 2.517072e-08, 2.474714e-08, 2.54514e-08, 
    2.78685e-08, 2.963935e-08, 2.84354e-08, 2.56979e-08, 2.420165e-08, 
    2.582412e-08, 2.710631e-08, 2.593838e-08, 2.458516e-08, 2.743937e-08,
  2.667828e-08, 2.649179e-08, 2.512507e-08, 2.469464e-08, 2.560646e-08, 
    2.773164e-08, 2.958503e-08, 2.941857e-08, 2.663569e-08, 2.41882e-08, 
    2.555933e-08, 2.720587e-08, 2.676772e-08, 2.468123e-08, 2.560209e-08,
  2.657964e-08, 2.675232e-08, 2.535752e-08, 2.454845e-08, 2.57424e-08, 
    2.76284e-08, 2.884794e-08, 2.858168e-08, 2.698902e-08, 2.469241e-08, 
    2.534245e-08, 2.687852e-08, 2.711731e-08, 2.564302e-08, 2.473814e-08,
  2.647844e-08, 2.68916e-08, 2.557578e-08, 2.452567e-08, 2.562094e-08, 
    2.751378e-08, 2.882575e-08, 2.852733e-08, 2.722913e-08, 2.626399e-08, 
    2.533484e-08, 2.653519e-08, 2.732719e-08, 2.640797e-08, 2.482777e-08,
  2.617572e-08, 2.696341e-08, 2.602811e-08, 2.453395e-08, 2.563501e-08, 
    2.736216e-08, 2.848676e-08, 2.866816e-08, 2.790839e-08, 2.695175e-08, 
    2.527471e-08, 2.591315e-08, 2.68258e-08, 2.687801e-08, 2.603704e-08,
  2.604051e-08, 2.692598e-08, 2.630866e-08, 2.468078e-08, 2.515146e-08, 
    2.707121e-08, 2.829832e-08, 2.904929e-08, 2.75463e-08, 2.715871e-08, 
    2.528004e-08, 2.575745e-08, 2.66377e-08, 2.659918e-08, 2.617199e-08,
  2.586302e-08, 2.693738e-08, 2.677182e-08, 2.484918e-08, 2.523226e-08, 
    2.679771e-08, 2.775193e-08, 2.852879e-08, 2.810955e-08, 2.641615e-08, 
    2.445866e-08, 2.580448e-08, 2.652211e-08, 2.649786e-08, 2.616894e-08,
  2.499156e-08, 2.609396e-08, 2.689792e-08, 2.563746e-08, 2.482207e-08, 
    2.670812e-08, 2.872121e-08, 2.938395e-08, 3.123701e-08, 2.851244e-08, 
    2.505876e-08, 2.523305e-08, 2.659251e-08, 2.654695e-08, 2.668216e-08,
  2.503936e-08, 2.633904e-08, 2.688922e-08, 2.566285e-08, 2.519043e-08, 
    2.69537e-08, 2.871842e-08, 3.0122e-08, 3.123127e-08, 2.690338e-08, 
    2.399987e-08, 2.499099e-08, 2.670281e-08, 2.613725e-08, 2.643803e-08,
  2.500888e-08, 2.615209e-08, 2.67334e-08, 2.568171e-08, 2.540386e-08, 
    2.776628e-08, 2.862483e-08, 2.929823e-08, 3.072484e-08, 2.59909e-08, 
    2.299649e-08, 2.49734e-08, 2.661741e-08, 2.596515e-08, 2.701562e-08,
  2.505842e-08, 2.632415e-08, 2.680508e-08, 2.58833e-08, 2.549333e-08, 
    2.808404e-08, 2.721858e-08, 2.934303e-08, 3.004238e-08, 2.436082e-08, 
    2.218006e-08, 2.496284e-08, 2.649699e-08, 2.617063e-08, 2.696185e-08,
  2.518156e-08, 2.625467e-08, 2.680165e-08, 2.584865e-08, 2.568728e-08, 
    2.615068e-08, 2.705618e-08, 3.202501e-08, 2.982781e-08, 2.137834e-08, 
    2.18891e-08, 2.53545e-08, 2.647817e-08, 2.599953e-08, 2.737961e-08,
  2.523259e-08, 2.639406e-08, 2.693431e-08, 2.598012e-08, 2.549559e-08, 
    2.615703e-08, 2.702352e-08, 2.929501e-08, 2.738002e-08, 2.290502e-08, 
    2.37423e-08, 2.572524e-08, 2.636544e-08, 2.616027e-08, 2.758901e-08,
  2.547648e-08, 2.620868e-08, 2.701076e-08, 2.601698e-08, 2.539485e-08, 
    2.576741e-08, 2.66784e-08, 2.773087e-08, 2.757388e-08, 2.583223e-08, 
    2.45472e-08, 2.63597e-08, 2.631243e-08, 2.606481e-08, 2.738509e-08,
  2.569962e-08, 2.632808e-08, 2.705595e-08, 2.625656e-08, 2.543152e-08, 
    2.573747e-08, 2.610137e-08, 2.754236e-08, 2.786284e-08, 2.588776e-08, 
    2.469199e-08, 2.634408e-08, 2.628052e-08, 2.631052e-08, 2.738633e-08,
  2.616923e-08, 2.618582e-08, 2.688968e-08, 2.634229e-08, 2.533148e-08, 
    2.551868e-08, 2.587163e-08, 2.682628e-08, 2.759477e-08, 2.624062e-08, 
    2.479499e-08, 2.64413e-08, 2.646242e-08, 2.626364e-08, 2.724968e-08,
  2.640876e-08, 2.626307e-08, 2.679935e-08, 2.650214e-08, 2.553475e-08, 
    2.556469e-08, 2.562053e-08, 2.659304e-08, 2.751091e-08, 2.744469e-08, 
    2.599437e-08, 2.613471e-08, 2.692198e-08, 2.677439e-08, 2.686358e-08,
  2.620038e-08, 2.636678e-08, 2.680301e-08, 2.707094e-08, 2.650974e-08, 
    2.630966e-08, 2.572695e-08, 2.672787e-08, 2.949646e-08, 2.991334e-08, 
    2.553076e-08, 2.213199e-08, 2.299998e-08, 2.46226e-08, 2.518481e-08,
  2.627188e-08, 2.668473e-08, 2.703767e-08, 2.709376e-08, 2.661749e-08, 
    2.629906e-08, 2.583138e-08, 2.739167e-08, 2.968468e-08, 2.874839e-08, 
    2.302572e-08, 2.224728e-08, 2.443516e-08, 2.540273e-08, 2.543202e-08,
  2.64915e-08, 2.710099e-08, 2.694895e-08, 2.706408e-08, 2.657551e-08, 
    2.650377e-08, 2.542271e-08, 2.755439e-08, 2.950344e-08, 2.762512e-08, 
    2.258709e-08, 2.367366e-08, 2.565361e-08, 2.607605e-08, 2.674219e-08,
  2.657024e-08, 2.734826e-08, 2.691394e-08, 2.71513e-08, 2.646602e-08, 
    2.651173e-08, 2.609086e-08, 2.759591e-08, 2.891035e-08, 2.623306e-08, 
    2.294166e-08, 2.476916e-08, 2.630067e-08, 2.648579e-08, 2.757519e-08,
  2.697222e-08, 2.758429e-08, 2.678486e-08, 2.726413e-08, 2.651953e-08, 
    2.622026e-08, 2.614945e-08, 2.797735e-08, 2.86749e-08, 2.482052e-08, 
    2.339297e-08, 2.6002e-08, 2.682841e-08, 2.70304e-08, 2.791787e-08,
  2.722634e-08, 2.757189e-08, 2.675992e-08, 2.735862e-08, 2.655534e-08, 
    2.640954e-08, 2.550358e-08, 2.695841e-08, 2.80031e-08, 2.58991e-08, 
    2.513135e-08, 2.652146e-08, 2.710778e-08, 2.710331e-08, 2.760794e-08,
  2.741373e-08, 2.755537e-08, 2.661938e-08, 2.741057e-08, 2.671478e-08, 
    2.634607e-08, 2.563449e-08, 2.656249e-08, 2.730883e-08, 2.583686e-08, 
    2.551175e-08, 2.732024e-08, 2.736318e-08, 2.699643e-08, 2.655443e-08,
  2.768041e-08, 2.736051e-08, 2.647737e-08, 2.745148e-08, 2.682587e-08, 
    2.653503e-08, 2.560171e-08, 2.641834e-08, 2.719942e-08, 2.611518e-08, 
    2.584875e-08, 2.731955e-08, 2.758709e-08, 2.668025e-08, 2.553962e-08,
  2.773101e-08, 2.718579e-08, 2.63758e-08, 2.768004e-08, 2.711992e-08, 
    2.677394e-08, 2.567456e-08, 2.626499e-08, 2.715084e-08, 2.601063e-08, 
    2.57223e-08, 2.761421e-08, 2.771344e-08, 2.652681e-08, 2.485341e-08,
  2.796563e-08, 2.705951e-08, 2.639927e-08, 2.767935e-08, 2.719939e-08, 
    2.707593e-08, 2.592348e-08, 2.608467e-08, 2.740801e-08, 2.619281e-08, 
    2.567558e-08, 2.763191e-08, 2.793485e-08, 2.621246e-08, 2.471256e-08,
  2.726608e-08, 2.709745e-08, 2.689179e-08, 2.737184e-08, 2.654208e-08, 
    2.673837e-08, 2.666043e-08, 2.820258e-08, 2.935372e-08, 2.699148e-08, 
    2.36747e-08, 2.393728e-08, 2.587051e-08, 2.655062e-08, 2.650822e-08,
  2.748397e-08, 2.735322e-08, 2.698012e-08, 2.762761e-08, 2.657245e-08, 
    2.627823e-08, 2.677721e-08, 2.806298e-08, 2.967607e-08, 2.704615e-08, 
    2.345854e-08, 2.434114e-08, 2.683685e-08, 2.727312e-08, 2.740513e-08,
  2.74116e-08, 2.711239e-08, 2.681325e-08, 2.766661e-08, 2.657945e-08, 
    2.628151e-08, 2.632382e-08, 2.824021e-08, 2.973444e-08, 2.668512e-08, 
    2.329843e-08, 2.486227e-08, 2.718169e-08, 2.767762e-08, 2.785478e-08,
  2.742497e-08, 2.717704e-08, 2.680783e-08, 2.772097e-08, 2.68139e-08, 
    2.65968e-08, 2.609153e-08, 2.736308e-08, 2.958888e-08, 2.638774e-08, 
    2.324545e-08, 2.536582e-08, 2.782117e-08, 2.766237e-08, 2.712284e-08,
  2.709209e-08, 2.705918e-08, 2.656147e-08, 2.764152e-08, 2.678959e-08, 
    2.617265e-08, 2.647111e-08, 2.705384e-08, 2.860565e-08, 2.506954e-08, 
    2.346642e-08, 2.595089e-08, 2.795038e-08, 2.734378e-08, 2.651599e-08,
  2.676057e-08, 2.711477e-08, 2.65229e-08, 2.761479e-08, 2.709038e-08, 
    2.650077e-08, 2.601686e-08, 2.666107e-08, 2.716799e-08, 2.55302e-08, 
    2.514523e-08, 2.6268e-08, 2.810806e-08, 2.735731e-08, 2.662574e-08,
  2.661255e-08, 2.705096e-08, 2.643001e-08, 2.766516e-08, 2.728097e-08, 
    2.626986e-08, 2.62589e-08, 2.641378e-08, 2.678888e-08, 2.614975e-08, 
    2.579264e-08, 2.711859e-08, 2.815937e-08, 2.714236e-08, 2.670151e-08,
  2.666968e-08, 2.702067e-08, 2.666559e-08, 2.819873e-08, 2.781073e-08, 
    2.644645e-08, 2.605498e-08, 2.640269e-08, 2.678222e-08, 2.686644e-08, 
    2.647157e-08, 2.696909e-08, 2.796207e-08, 2.702397e-08, 2.720144e-08,
  2.652203e-08, 2.676567e-08, 2.722328e-08, 2.894785e-08, 2.813212e-08, 
    2.588826e-08, 2.584296e-08, 2.644135e-08, 2.67139e-08, 2.642806e-08, 
    2.620055e-08, 2.705686e-08, 2.785072e-08, 2.682759e-08, 2.740635e-08,
  2.645374e-08, 2.683368e-08, 2.852608e-08, 2.981291e-08, 2.807205e-08, 
    2.503575e-08, 2.533067e-08, 2.647281e-08, 2.68693e-08, 2.610411e-08, 
    2.62385e-08, 2.70104e-08, 2.771948e-08, 2.680397e-08, 2.740385e-08,
  3.108387e-08, 2.912149e-08, 2.728888e-08, 2.697366e-08, 2.673714e-08, 
    2.720153e-08, 2.865059e-08, 2.890375e-08, 2.762983e-08, 2.714477e-08, 
    2.601444e-08, 2.568147e-08, 2.609783e-08, 2.707436e-08, 2.715159e-08,
  3.097505e-08, 2.879802e-08, 2.71991e-08, 2.713214e-08, 2.699955e-08, 
    2.750747e-08, 2.906538e-08, 2.918246e-08, 2.773803e-08, 2.720197e-08, 
    2.64438e-08, 2.573445e-08, 2.61756e-08, 2.673861e-08, 2.674122e-08,
  3.043689e-08, 2.831157e-08, 2.712273e-08, 2.704952e-08, 2.714711e-08, 
    2.826753e-08, 2.92203e-08, 2.911918e-08, 2.724145e-08, 2.720026e-08, 
    2.653042e-08, 2.567402e-08, 2.567355e-08, 2.645308e-08, 2.671517e-08,
  2.938886e-08, 2.779871e-08, 2.697127e-08, 2.697979e-08, 2.731901e-08, 
    2.868515e-08, 2.930025e-08, 2.813203e-08, 2.70872e-08, 2.743932e-08, 
    2.657336e-08, 2.538393e-08, 2.5242e-08, 2.571597e-08, 2.621971e-08,
  2.838927e-08, 2.750387e-08, 2.683671e-08, 2.68112e-08, 2.779343e-08, 
    2.905935e-08, 2.962729e-08, 2.781934e-08, 2.760738e-08, 2.747073e-08, 
    2.611654e-08, 2.496655e-08, 2.484792e-08, 2.568531e-08, 2.577205e-08,
  2.751058e-08, 2.70278e-08, 2.668327e-08, 2.68548e-08, 2.845822e-08, 
    3.078648e-08, 2.980798e-08, 2.796149e-08, 2.745358e-08, 2.601953e-08, 
    2.468523e-08, 2.473428e-08, 2.566928e-08, 2.654631e-08, 2.689106e-08,
  2.685661e-08, 2.717702e-08, 2.688974e-08, 2.717112e-08, 2.952204e-08, 
    3.102689e-08, 2.950244e-08, 2.755831e-08, 2.615521e-08, 2.463889e-08, 
    2.53905e-08, 2.666305e-08, 2.713671e-08, 2.710928e-08, 2.71075e-08,
  2.791594e-08, 2.744538e-08, 2.67097e-08, 2.767642e-08, 3.025562e-08, 
    3.15125e-08, 2.86929e-08, 2.639294e-08, 2.524061e-08, 2.634305e-08, 
    2.71251e-08, 2.681718e-08, 2.677857e-08, 2.673513e-08, 2.69253e-08,
  2.806705e-08, 2.654205e-08, 2.702833e-08, 2.825804e-08, 3.06869e-08, 
    3.073892e-08, 2.734962e-08, 2.5606e-08, 2.608339e-08, 2.662346e-08, 
    2.660461e-08, 2.653223e-08, 2.676272e-08, 2.68427e-08, 2.713204e-08,
  2.62499e-08, 2.662303e-08, 2.767078e-08, 2.897202e-08, 3.006899e-08, 
    2.881501e-08, 2.675356e-08, 2.649051e-08, 2.649908e-08, 2.668759e-08, 
    2.670567e-08, 2.651572e-08, 2.664695e-08, 2.69741e-08, 2.725965e-08,
  2.935515e-08, 2.972414e-08, 2.981151e-08, 3.026435e-08, 3.00616e-08, 
    2.885287e-08, 2.770468e-08, 2.806967e-08, 2.858931e-08, 2.911334e-08, 
    2.798941e-08, 2.736834e-08, 2.665164e-08, 2.686672e-08, 2.653916e-08,
  2.943036e-08, 2.94927e-08, 2.97531e-08, 2.99182e-08, 2.941042e-08, 
    2.805977e-08, 2.763755e-08, 2.850131e-08, 2.86544e-08, 2.790553e-08, 
    2.79126e-08, 2.759804e-08, 2.693619e-08, 2.619813e-08, 2.619142e-08,
  2.918687e-08, 2.921567e-08, 2.929437e-08, 2.917616e-08, 2.855934e-08, 
    2.813239e-08, 2.770142e-08, 2.894838e-08, 2.843105e-08, 2.730418e-08, 
    2.750066e-08, 2.770693e-08, 2.726972e-08, 2.657145e-08, 2.57421e-08,
  2.890192e-08, 2.867138e-08, 2.860544e-08, 2.868843e-08, 2.81421e-08, 
    2.768758e-08, 2.824913e-08, 2.902022e-08, 2.751749e-08, 2.721495e-08, 
    2.73135e-08, 2.730083e-08, 2.726e-08, 2.688927e-08, 2.624279e-08,
  2.836132e-08, 2.807588e-08, 2.831875e-08, 2.810183e-08, 2.74799e-08, 
    2.723976e-08, 2.819562e-08, 2.85163e-08, 2.759813e-08, 2.684033e-08, 
    2.700735e-08, 2.698923e-08, 2.689452e-08, 2.677768e-08, 2.682839e-08,
  2.78379e-08, 2.800961e-08, 2.813504e-08, 2.764292e-08, 2.72694e-08, 
    2.806738e-08, 2.713564e-08, 2.712604e-08, 2.672094e-08, 2.71533e-08, 
    2.729736e-08, 2.716333e-08, 2.702474e-08, 2.674405e-08, 2.680219e-08,
  2.839559e-08, 2.79135e-08, 2.750137e-08, 2.726497e-08, 2.737461e-08, 
    2.799996e-08, 2.796564e-08, 2.754552e-08, 2.685583e-08, 2.723418e-08, 
    2.679301e-08, 2.698082e-08, 2.671144e-08, 2.667611e-08, 2.628752e-08,
  2.805712e-08, 2.683407e-08, 2.735389e-08, 2.734602e-08, 2.776956e-08, 
    2.842914e-08, 2.748916e-08, 2.740934e-08, 2.719383e-08, 2.71034e-08, 
    2.692548e-08, 2.701032e-08, 2.676978e-08, 2.645257e-08, 2.590955e-08,
  2.685817e-08, 2.65269e-08, 2.763684e-08, 2.747117e-08, 2.814752e-08, 
    2.808629e-08, 2.780806e-08, 2.759929e-08, 2.703062e-08, 2.697941e-08, 
    2.661866e-08, 2.65616e-08, 2.606154e-08, 2.570583e-08, 2.55283e-08,
  2.678215e-08, 2.655866e-08, 2.807558e-08, 2.738746e-08, 2.820634e-08, 
    2.806516e-08, 2.762069e-08, 2.740726e-08, 2.681603e-08, 2.644364e-08, 
    2.639482e-08, 2.620476e-08, 2.57981e-08, 2.579546e-08, 2.578218e-08,
  2.722838e-08, 2.670785e-08, 2.724778e-08, 2.743082e-08, 2.764499e-08, 
    2.792537e-08, 2.730308e-08, 2.747351e-08, 2.798279e-08, 2.798553e-08, 
    2.726636e-08, 2.704936e-08, 2.696207e-08, 2.703678e-08, 2.743174e-08,
  2.705109e-08, 2.667919e-08, 2.725019e-08, 2.757378e-08, 2.798943e-08, 
    2.803081e-08, 2.761677e-08, 2.795046e-08, 2.777135e-08, 2.684858e-08, 
    2.628732e-08, 2.661567e-08, 2.656771e-08, 2.715287e-08, 2.641498e-08,
  2.68977e-08, 2.657192e-08, 2.739939e-08, 2.770523e-08, 2.832707e-08, 
    2.845438e-08, 2.72733e-08, 2.80637e-08, 2.726257e-08, 2.593184e-08, 
    2.579219e-08, 2.625715e-08, 2.658233e-08, 2.637416e-08, 2.621474e-08,
  2.700615e-08, 2.672072e-08, 2.752564e-08, 2.77521e-08, 2.835433e-08, 
    2.903464e-08, 2.781214e-08, 2.809746e-08, 2.636429e-08, 2.484142e-08, 
    2.537524e-08, 2.617599e-08, 2.672272e-08, 2.657317e-08, 2.686949e-08,
  2.698713e-08, 2.67349e-08, 2.763585e-08, 2.776732e-08, 2.811814e-08, 
    2.781669e-08, 2.840448e-08, 2.923032e-08, 2.607044e-08, 2.404844e-08, 
    2.535637e-08, 2.606605e-08, 2.66513e-08, 2.686089e-08, 2.68573e-08,
  2.705061e-08, 2.684407e-08, 2.770886e-08, 2.781615e-08, 2.81983e-08, 
    2.787948e-08, 2.747062e-08, 2.76351e-08, 2.606821e-08, 2.536863e-08, 
    2.549042e-08, 2.559144e-08, 2.613694e-08, 2.638545e-08, 2.659438e-08,
  2.701894e-08, 2.68787e-08, 2.77475e-08, 2.781653e-08, 2.812797e-08, 
    2.74844e-08, 2.76271e-08, 2.750877e-08, 2.584146e-08, 2.499758e-08, 
    2.534295e-08, 2.529232e-08, 2.560748e-08, 2.616417e-08, 2.67557e-08,
  2.714179e-08, 2.693709e-08, 2.777595e-08, 2.789742e-08, 2.822324e-08, 
    2.751727e-08, 2.74702e-08, 2.754286e-08, 2.568543e-08, 2.479285e-08, 
    2.527813e-08, 2.524468e-08, 2.510963e-08, 2.553544e-08, 2.64354e-08,
  2.715321e-08, 2.696295e-08, 2.771846e-08, 2.796148e-08, 2.853711e-08, 
    2.748863e-08, 2.744666e-08, 2.755771e-08, 2.564514e-08, 2.462532e-08, 
    2.50991e-08, 2.521258e-08, 2.487856e-08, 2.49284e-08, 2.559258e-08,
  2.722825e-08, 2.696454e-08, 2.76839e-08, 2.796583e-08, 2.873683e-08, 
    2.775048e-08, 2.742028e-08, 2.761893e-08, 2.59787e-08, 2.48083e-08, 
    2.514256e-08, 2.525908e-08, 2.480519e-08, 2.492448e-08, 2.516475e-08,
  2.75952e-08, 2.766894e-08, 2.824285e-08, 2.82701e-08, 2.87359e-08, 
    2.83856e-08, 2.897386e-08, 2.76216e-08, 2.643974e-08, 2.559999e-08, 
    2.520412e-08, 2.524981e-08, 2.569835e-08, 2.662055e-08, 2.71404e-08,
  2.763358e-08, 2.771004e-08, 2.815944e-08, 2.808748e-08, 2.885134e-08, 
    2.836516e-08, 2.897975e-08, 2.814297e-08, 2.707415e-08, 2.594317e-08, 
    2.540136e-08, 2.526079e-08, 2.566216e-08, 2.651063e-08, 2.617764e-08,
  2.769659e-08, 2.749281e-08, 2.797949e-08, 2.810518e-08, 2.900172e-08, 
    2.836832e-08, 2.881334e-08, 2.746619e-08, 2.747224e-08, 2.653202e-08, 
    2.572488e-08, 2.532444e-08, 2.552882e-08, 2.594921e-08, 2.620472e-08,
  2.78475e-08, 2.753849e-08, 2.794852e-08, 2.809253e-08, 2.886448e-08, 
    2.892455e-08, 2.795876e-08, 2.726327e-08, 2.78684e-08, 2.672579e-08, 
    2.625298e-08, 2.536275e-08, 2.540614e-08, 2.556871e-08, 2.638678e-08,
  2.779602e-08, 2.743962e-08, 2.770323e-08, 2.795948e-08, 2.887039e-08, 
    2.848822e-08, 2.824836e-08, 2.89912e-08, 2.84053e-08, 2.620973e-08, 
    2.616135e-08, 2.568052e-08, 2.539897e-08, 2.543852e-08, 2.59448e-08,
  2.78166e-08, 2.755725e-08, 2.77357e-08, 2.805272e-08, 2.881634e-08, 
    2.831116e-08, 2.86628e-08, 2.849579e-08, 2.822381e-08, 2.680327e-08, 
    2.624272e-08, 2.592911e-08, 2.571013e-08, 2.52993e-08, 2.546979e-08,
  2.786171e-08, 2.754441e-08, 2.760133e-08, 2.805324e-08, 2.88705e-08, 
    2.836e-08, 2.852829e-08, 2.809714e-08, 2.780071e-08, 2.687612e-08, 
    2.653572e-08, 2.632122e-08, 2.616691e-08, 2.554675e-08, 2.56392e-08,
  2.79259e-08, 2.773927e-08, 2.770936e-08, 2.832304e-08, 2.890818e-08, 
    2.833858e-08, 2.806095e-08, 2.797752e-08, 2.784844e-08, 2.724022e-08, 
    2.638818e-08, 2.660541e-08, 2.665829e-08, 2.612444e-08, 2.556082e-08,
  2.829483e-08, 2.773883e-08, 2.749781e-08, 2.826334e-08, 2.884248e-08, 
    2.839339e-08, 2.784302e-08, 2.787544e-08, 2.779449e-08, 2.707176e-08, 
    2.650408e-08, 2.704581e-08, 2.714226e-08, 2.661629e-08, 2.573756e-08,
  2.83252e-08, 2.754135e-08, 2.769209e-08, 2.845523e-08, 2.894047e-08, 
    2.822065e-08, 2.773642e-08, 2.752296e-08, 2.731701e-08, 2.7083e-08, 
    2.678288e-08, 2.741464e-08, 2.730774e-08, 2.716023e-08, 2.62918e-08,
  2.763392e-08, 2.773371e-08, 2.771611e-08, 2.734472e-08, 2.75944e-08, 
    2.837819e-08, 2.899097e-08, 2.646632e-08, 2.640788e-08, 2.688187e-08, 
    2.715549e-08, 2.677717e-08, 2.644201e-08, 2.614069e-08, 2.626323e-08,
  2.756066e-08, 2.752978e-08, 2.741591e-08, 2.726161e-08, 2.716873e-08, 
    2.793619e-08, 2.847826e-08, 2.677184e-08, 2.620307e-08, 2.622358e-08, 
    2.745976e-08, 2.676691e-08, 2.65243e-08, 2.606086e-08, 2.586034e-08,
  2.748744e-08, 2.68505e-08, 2.696633e-08, 2.706379e-08, 2.684117e-08, 
    2.761716e-08, 2.764919e-08, 2.539885e-08, 2.591816e-08, 2.672228e-08, 
    2.741189e-08, 2.678697e-08, 2.661911e-08, 2.616731e-08, 2.578775e-08,
  2.723969e-08, 2.662287e-08, 2.667052e-08, 2.66375e-08, 2.645338e-08, 
    2.732152e-08, 2.51598e-08, 2.550529e-08, 2.61592e-08, 2.659493e-08, 
    2.67147e-08, 2.621283e-08, 2.66677e-08, 2.638014e-08, 2.626216e-08,
  2.693465e-08, 2.629038e-08, 2.626623e-08, 2.614746e-08, 2.651571e-08, 
    2.623027e-08, 2.544529e-08, 2.701085e-08, 2.67545e-08, 2.605552e-08, 
    2.645392e-08, 2.661297e-08, 2.679701e-08, 2.659326e-08, 2.670465e-08,
  2.682336e-08, 2.603662e-08, 2.591687e-08, 2.566375e-08, 2.587049e-08, 
    2.666753e-08, 2.603412e-08, 2.599709e-08, 2.6179e-08, 2.648692e-08, 
    2.6367e-08, 2.634094e-08, 2.671887e-08, 2.68007e-08, 2.69455e-08,
  2.686698e-08, 2.56113e-08, 2.542476e-08, 2.513025e-08, 2.616698e-08, 
    2.638317e-08, 2.628243e-08, 2.617816e-08, 2.602069e-08, 2.650291e-08, 
    2.630562e-08, 2.673367e-08, 2.674318e-08, 2.713661e-08, 2.710493e-08,
  2.66602e-08, 2.524259e-08, 2.500371e-08, 2.505919e-08, 2.60714e-08, 
    2.611465e-08, 2.623143e-08, 2.656712e-08, 2.654137e-08, 2.65613e-08, 
    2.669104e-08, 2.678978e-08, 2.680313e-08, 2.710274e-08, 2.721296e-08,
  2.630402e-08, 2.475428e-08, 2.478111e-08, 2.488656e-08, 2.601253e-08, 
    2.615681e-08, 2.659308e-08, 2.676229e-08, 2.685652e-08, 2.695307e-08, 
    2.688869e-08, 2.705634e-08, 2.704316e-08, 2.719765e-08, 2.727528e-08,
  2.58366e-08, 2.444935e-08, 2.470582e-08, 2.491405e-08, 2.600012e-08, 
    2.617398e-08, 2.678472e-08, 2.699694e-08, 2.690516e-08, 2.696219e-08, 
    2.714308e-08, 2.737808e-08, 2.740965e-08, 2.744622e-08, 2.749083e-08,
  2.493053e-08, 2.463687e-08, 2.472175e-08, 2.461994e-08, 2.459241e-08, 
    2.475591e-08, 2.523203e-08, 2.595983e-08, 2.612583e-08, 2.603208e-08, 
    2.578788e-08, 2.530725e-08, 2.493687e-08, 2.536775e-08, 2.568108e-08,
  2.482454e-08, 2.478142e-08, 2.476238e-08, 2.48885e-08, 2.51916e-08, 
    2.580969e-08, 2.678386e-08, 2.678144e-08, 2.706838e-08, 2.645135e-08, 
    2.627838e-08, 2.544356e-08, 2.596616e-08, 2.503908e-08, 2.553782e-08,
  2.487597e-08, 2.464333e-08, 2.480236e-08, 2.516072e-08, 2.585351e-08, 
    2.712497e-08, 2.755787e-08, 2.756773e-08, 2.753253e-08, 2.671526e-08, 
    2.636505e-08, 2.572183e-08, 2.597635e-08, 2.568478e-08, 2.517122e-08,
  2.480896e-08, 2.447855e-08, 2.495399e-08, 2.547119e-08, 2.668394e-08, 
    2.823391e-08, 2.880166e-08, 2.836939e-08, 2.793088e-08, 2.718015e-08, 
    2.648544e-08, 2.604931e-08, 2.574813e-08, 2.570973e-08, 2.579533e-08,
  2.478812e-08, 2.441754e-08, 2.511547e-08, 2.58583e-08, 2.734892e-08, 
    2.811042e-08, 2.966076e-08, 2.971223e-08, 2.877814e-08, 2.735483e-08, 
    2.620977e-08, 2.611993e-08, 2.613472e-08, 2.52037e-08, 2.612048e-08,
  2.469279e-08, 2.432464e-08, 2.526621e-08, 2.631044e-08, 2.758721e-08, 
    2.866599e-08, 2.886919e-08, 3.039811e-08, 2.983184e-08, 2.728255e-08, 
    2.668629e-08, 2.605386e-08, 2.641391e-08, 2.522086e-08, 2.620106e-08,
  2.456548e-08, 2.440758e-08, 2.553313e-08, 2.663518e-08, 2.78637e-08, 
    2.866618e-08, 2.928478e-08, 2.92398e-08, 2.87662e-08, 2.822183e-08, 
    2.760406e-08, 2.655158e-08, 2.646857e-08, 2.543908e-08, 2.632718e-08,
  2.442672e-08, 2.441946e-08, 2.562126e-08, 2.678883e-08, 2.761927e-08, 
    2.871148e-08, 2.914967e-08, 2.931617e-08, 2.876295e-08, 2.811655e-08, 
    2.803815e-08, 2.740302e-08, 2.691346e-08, 2.576892e-08, 2.637224e-08,
  2.416778e-08, 2.443971e-08, 2.564836e-08, 2.680392e-08, 2.750271e-08, 
    2.843353e-08, 2.890302e-08, 2.893745e-08, 2.854891e-08, 2.752119e-08, 
    2.757855e-08, 2.783935e-08, 2.728475e-08, 2.621415e-08, 2.632499e-08,
  2.403757e-08, 2.441409e-08, 2.551171e-08, 2.654767e-08, 2.718531e-08, 
    2.77658e-08, 2.84663e-08, 2.896067e-08, 2.881103e-08, 2.7647e-08, 
    2.694635e-08, 2.762461e-08, 2.770166e-08, 2.679788e-08, 2.642018e-08,
  2.30926e-08, 2.508561e-08, 2.647016e-08, 2.695777e-08, 2.822894e-08, 
    2.89934e-08, 2.912425e-08, 2.970489e-08, 2.97463e-08, 2.924876e-08, 
    2.836201e-08, 2.792317e-08, 2.629393e-08, 2.519938e-08, 2.554777e-08,
  2.308146e-08, 2.515134e-08, 2.652353e-08, 2.695426e-08, 2.833655e-08, 
    2.898529e-08, 2.926219e-08, 2.998311e-08, 2.967929e-08, 3.061897e-08, 
    2.94444e-08, 2.861265e-08, 2.780446e-08, 2.646562e-08, 2.511717e-08,
  2.283357e-08, 2.442397e-08, 2.650679e-08, 2.68616e-08, 2.82884e-08, 
    2.875282e-08, 2.883482e-08, 2.923187e-08, 2.907281e-08, 2.994318e-08, 
    3.041432e-08, 2.927677e-08, 2.847246e-08, 2.727963e-08, 2.580918e-08,
  2.276695e-08, 2.40124e-08, 2.628683e-08, 2.674429e-08, 2.767958e-08, 
    2.908107e-08, 2.870934e-08, 2.797257e-08, 2.764398e-08, 2.961867e-08, 
    2.934443e-08, 2.897437e-08, 2.828609e-08, 2.774808e-08, 2.633051e-08,
  2.280952e-08, 2.312422e-08, 2.594956e-08, 2.664651e-08, 2.747372e-08, 
    2.813819e-08, 2.784867e-08, 2.921798e-08, 2.816118e-08, 2.787813e-08, 
    2.828835e-08, 2.838439e-08, 2.820016e-08, 2.777434e-08, 2.638274e-08,
  2.309931e-08, 2.259743e-08, 2.53708e-08, 2.640222e-08, 2.718799e-08, 
    2.809722e-08, 2.761881e-08, 2.839642e-08, 2.697037e-08, 2.60993e-08, 
    2.770763e-08, 2.752055e-08, 2.762639e-08, 2.731809e-08, 2.61425e-08,
  2.372928e-08, 2.189821e-08, 2.456675e-08, 2.610267e-08, 2.678216e-08, 
    2.786838e-08, 2.743473e-08, 2.787566e-08, 2.766461e-08, 2.751173e-08, 
    2.701095e-08, 2.693412e-08, 2.701542e-08, 2.667204e-08, 2.575983e-08,
  2.469216e-08, 2.177614e-08, 2.357949e-08, 2.572918e-08, 2.639254e-08, 
    2.776613e-08, 2.75021e-08, 2.770002e-08, 2.750192e-08, 2.68705e-08, 
    2.686684e-08, 2.636944e-08, 2.666671e-08, 2.578421e-08, 2.53486e-08,
  2.615579e-08, 2.196703e-08, 2.240142e-08, 2.520108e-08, 2.607347e-08, 
    2.723746e-08, 2.748366e-08, 2.765987e-08, 2.785791e-08, 2.692843e-08, 
    2.695282e-08, 2.655132e-08, 2.633763e-08, 2.527606e-08, 2.507802e-08,
  2.721027e-08, 2.271985e-08, 2.115222e-08, 2.433699e-08, 2.544768e-08, 
    2.701555e-08, 2.750659e-08, 2.711175e-08, 2.802552e-08, 2.741654e-08, 
    2.679585e-08, 2.656715e-08, 2.586995e-08, 2.522911e-08, 2.529156e-08,
  2.489534e-08, 2.415621e-08, 2.452026e-08, 2.774938e-08, 2.830217e-08, 
    2.814752e-08, 2.686333e-08, 2.682504e-08, 2.895089e-08, 3.039942e-08, 
    2.792048e-08, 2.598946e-08, 2.518666e-08, 2.601444e-08, 2.479199e-08,
  2.508488e-08, 2.42481e-08, 2.437377e-08, 2.776311e-08, 2.836244e-08, 
    2.833653e-08, 2.699145e-08, 2.693917e-08, 2.803886e-08, 3.023596e-08, 
    2.868646e-08, 2.697451e-08, 2.552766e-08, 2.574751e-08, 2.5043e-08,
  2.51384e-08, 2.430051e-08, 2.387581e-08, 2.761067e-08, 2.818314e-08, 
    2.827052e-08, 2.695699e-08, 2.641956e-08, 2.812934e-08, 2.977824e-08, 
    2.958467e-08, 2.83965e-08, 2.639656e-08, 2.583883e-08, 2.500506e-08,
  2.539993e-08, 2.443491e-08, 2.363791e-08, 2.736282e-08, 2.807739e-08, 
    2.847025e-08, 2.75501e-08, 2.659013e-08, 2.756044e-08, 3.032886e-08, 
    3.01813e-08, 2.962752e-08, 2.74244e-08, 2.656565e-08, 2.584101e-08,
  2.553355e-08, 2.456367e-08, 2.316363e-08, 2.701738e-08, 2.777446e-08, 
    2.70354e-08, 2.82647e-08, 2.77439e-08, 2.738564e-08, 2.905123e-08, 
    3.03978e-08, 2.995216e-08, 2.807162e-08, 2.714807e-08, 2.651246e-08,
  2.56512e-08, 2.474434e-08, 2.287281e-08, 2.6414e-08, 2.786907e-08, 
    2.713088e-08, 2.667193e-08, 2.803773e-08, 2.840914e-08, 2.785277e-08, 
    2.932854e-08, 2.905781e-08, 2.879068e-08, 2.784109e-08, 2.695543e-08,
  2.564458e-08, 2.492168e-08, 2.276082e-08, 2.564217e-08, 2.764026e-08, 
    2.729415e-08, 2.653841e-08, 2.616793e-08, 2.691957e-08, 2.760043e-08, 
    2.837722e-08, 2.882531e-08, 2.885452e-08, 2.799223e-08, 2.704989e-08,
  2.558271e-08, 2.514891e-08, 2.285758e-08, 2.476469e-08, 2.74682e-08, 
    2.708238e-08, 2.661131e-08, 2.615144e-08, 2.640098e-08, 2.626863e-08, 
    2.675701e-08, 2.725683e-08, 2.784144e-08, 2.756559e-08, 2.71317e-08,
  2.548973e-08, 2.531861e-08, 2.313934e-08, 2.373001e-08, 2.699325e-08, 
    2.727236e-08, 2.647461e-08, 2.577287e-08, 2.587459e-08, 2.5939e-08, 
    2.56943e-08, 2.543146e-08, 2.585943e-08, 2.612327e-08, 2.627715e-08,
  2.548181e-08, 2.553759e-08, 2.369776e-08, 2.309168e-08, 2.635801e-08, 
    2.720232e-08, 2.679705e-08, 2.579929e-08, 2.5489e-08, 2.550423e-08, 
    2.526197e-08, 2.499281e-08, 2.453248e-08, 2.447854e-08, 2.423374e-08,
  2.364392e-08, 2.435217e-08, 2.428195e-08, 2.517708e-08, 2.658023e-08, 
    2.667801e-08, 2.751607e-08, 2.945131e-08, 3.006239e-08, 2.728143e-08, 
    2.452592e-08, 2.492777e-08, 2.527154e-08, 2.505622e-08, 2.543209e-08,
  2.379044e-08, 2.481047e-08, 2.432297e-08, 2.544679e-08, 2.672635e-08, 
    2.693396e-08, 2.799053e-08, 2.945641e-08, 2.983808e-08, 2.791281e-08, 
    2.458616e-08, 2.512268e-08, 2.465328e-08, 2.451068e-08, 2.613783e-08,
  2.44789e-08, 2.494732e-08, 2.377507e-08, 2.588224e-08, 2.664729e-08, 
    2.639793e-08, 2.798139e-08, 2.947214e-08, 3.005086e-08, 2.739376e-08, 
    2.486756e-08, 2.514746e-08, 2.505781e-08, 2.487601e-08, 2.598183e-08,
  2.503241e-08, 2.429421e-08, 2.402406e-08, 2.650215e-08, 2.627519e-08, 
    2.626927e-08, 2.759709e-08, 2.813167e-08, 2.94172e-08, 2.765755e-08, 
    2.489904e-08, 2.510476e-08, 2.510259e-08, 2.471828e-08, 2.549694e-08,
  2.502042e-08, 2.387547e-08, 2.432917e-08, 2.670284e-08, 2.598359e-08, 
    2.526562e-08, 2.774325e-08, 2.747638e-08, 2.877954e-08, 2.910823e-08, 
    2.642579e-08, 2.534837e-08, 2.53046e-08, 2.504036e-08, 2.508712e-08,
  2.469008e-08, 2.367956e-08, 2.479226e-08, 2.681149e-08, 2.603948e-08, 
    2.500114e-08, 2.557441e-08, 2.709685e-08, 2.803748e-08, 2.896999e-08, 
    2.860451e-08, 2.606604e-08, 2.540098e-08, 2.53874e-08, 2.506912e-08,
  2.471856e-08, 2.37542e-08, 2.462436e-08, 2.662278e-08, 2.617028e-08, 
    2.514341e-08, 2.540316e-08, 2.52979e-08, 2.57167e-08, 2.854603e-08, 
    2.887434e-08, 2.751559e-08, 2.585622e-08, 2.557056e-08, 2.516386e-08,
  2.503976e-08, 2.37092e-08, 2.42893e-08, 2.615862e-08, 2.651019e-08, 
    2.531788e-08, 2.560783e-08, 2.538155e-08, 2.467032e-08, 2.490524e-08, 
    2.812808e-08, 2.836383e-08, 2.695052e-08, 2.563223e-08, 2.568385e-08,
  2.51938e-08, 2.422158e-08, 2.364397e-08, 2.530616e-08, 2.648171e-08, 
    2.600748e-08, 2.599936e-08, 2.65047e-08, 2.574309e-08, 2.413014e-08, 
    2.473686e-08, 2.653959e-08, 2.768609e-08, 2.690861e-08, 2.494632e-08,
  2.533323e-08, 2.48005e-08, 2.363049e-08, 2.430607e-08, 2.573857e-08, 
    2.618868e-08, 2.615626e-08, 2.689012e-08, 2.755385e-08, 2.658588e-08, 
    2.487719e-08, 2.503897e-08, 2.535097e-08, 2.59505e-08, 2.532411e-08,
  2.423883e-08, 2.452416e-08, 2.472687e-08, 2.499863e-08, 2.554559e-08, 
    2.553023e-08, 2.588482e-08, 2.67884e-08, 2.872935e-08, 2.746564e-08, 
    2.549368e-08, 2.499763e-08, 2.513577e-08, 2.630203e-08, 2.77921e-08,
  2.460569e-08, 2.437601e-08, 2.465991e-08, 2.541993e-08, 2.579346e-08, 
    2.548e-08, 2.588099e-08, 2.710061e-08, 2.868798e-08, 2.679308e-08, 
    2.508735e-08, 2.483917e-08, 2.517381e-08, 2.795005e-08, 2.892178e-08,
  2.431232e-08, 2.384437e-08, 2.497234e-08, 2.628651e-08, 2.587491e-08, 
    2.502724e-08, 2.603231e-08, 2.734204e-08, 2.868423e-08, 2.559451e-08, 
    2.520118e-08, 2.529709e-08, 2.622661e-08, 2.908823e-08, 2.915725e-08,
  2.387305e-08, 2.37739e-08, 2.592155e-08, 2.678595e-08, 2.523235e-08, 
    2.59656e-08, 2.57453e-08, 2.650116e-08, 2.795457e-08, 2.505718e-08, 
    2.513835e-08, 2.51254e-08, 2.581772e-08, 2.843316e-08, 2.904318e-08,
  2.402716e-08, 2.397248e-08, 2.553471e-08, 2.651036e-08, 2.611796e-08, 
    2.587666e-08, 2.653047e-08, 2.581442e-08, 2.68963e-08, 2.767811e-08, 
    2.453461e-08, 2.51536e-08, 2.530243e-08, 2.76323e-08, 2.87827e-08,
  2.454146e-08, 2.387183e-08, 2.485352e-08, 2.633891e-08, 2.642316e-08, 
    2.647294e-08, 2.619869e-08, 2.654645e-08, 2.786514e-08, 2.816695e-08, 
    2.476884e-08, 2.506732e-08, 2.544673e-08, 2.627277e-08, 2.796749e-08,
  2.469116e-08, 2.399412e-08, 2.431244e-08, 2.555277e-08, 2.669539e-08, 
    2.707655e-08, 2.708964e-08, 2.583793e-08, 2.600486e-08, 2.823723e-08, 
    2.690125e-08, 2.48928e-08, 2.558924e-08, 2.576904e-08, 2.6545e-08,
  2.49734e-08, 2.446394e-08, 2.389553e-08, 2.460969e-08, 2.586267e-08, 
    2.717065e-08, 2.794031e-08, 2.758116e-08, 2.561162e-08, 2.658945e-08, 
    2.80221e-08, 2.594402e-08, 2.530241e-08, 2.549526e-08, 2.625404e-08,
  2.494281e-08, 2.48029e-08, 2.419586e-08, 2.387259e-08, 2.483564e-08, 
    2.600439e-08, 2.76978e-08, 2.852254e-08, 2.735228e-08, 2.554832e-08, 
    2.669831e-08, 2.712741e-08, 2.601644e-08, 2.520715e-08, 2.567068e-08,
  2.484001e-08, 2.495617e-08, 2.480049e-08, 2.410303e-08, 2.403179e-08, 
    2.467321e-08, 2.617106e-08, 2.804811e-08, 2.871639e-08, 2.769666e-08, 
    2.632038e-08, 2.631095e-08, 2.637631e-08, 2.606704e-08, 2.565286e-08,
  2.459292e-08, 2.369321e-08, 2.358254e-08, 2.487347e-08, 2.620404e-08, 
    2.673036e-08, 2.640379e-08, 2.552016e-08, 2.627442e-08, 2.75207e-08, 
    2.766497e-08, 2.62102e-08, 2.512689e-08, 2.657601e-08, 2.849417e-08,
  2.44529e-08, 2.383821e-08, 2.436257e-08, 2.561569e-08, 2.669124e-08, 
    2.676049e-08, 2.641183e-08, 2.592528e-08, 2.706704e-08, 2.743218e-08, 
    2.652929e-08, 2.512282e-08, 2.576924e-08, 2.780896e-08, 2.903808e-08,
  2.462023e-08, 2.407502e-08, 2.445154e-08, 2.528096e-08, 2.676532e-08, 
    2.704908e-08, 2.67631e-08, 2.605283e-08, 2.739878e-08, 2.693147e-08, 
    2.586212e-08, 2.522119e-08, 2.597831e-08, 2.847289e-08, 2.910311e-08,
  2.470274e-08, 2.426997e-08, 2.415839e-08, 2.516881e-08, 2.669408e-08, 
    2.784753e-08, 2.678407e-08, 2.635222e-08, 2.742079e-08, 2.669181e-08, 
    2.573264e-08, 2.522663e-08, 2.597333e-08, 2.783172e-08, 2.887702e-08,
  2.488349e-08, 2.45705e-08, 2.425041e-08, 2.465278e-08, 2.590901e-08, 
    2.734189e-08, 2.759694e-08, 2.592045e-08, 2.560551e-08, 2.805613e-08, 
    2.570834e-08, 2.532895e-08, 2.609802e-08, 2.738818e-08, 2.895199e-08,
  2.481799e-08, 2.47403e-08, 2.43915e-08, 2.420758e-08, 2.54637e-08, 
    2.718204e-08, 2.75846e-08, 2.697151e-08, 2.72712e-08, 2.806853e-08, 
    2.578161e-08, 2.532189e-08, 2.590645e-08, 2.687906e-08, 2.880827e-08,
  2.47967e-08, 2.485793e-08, 2.456327e-08, 2.400761e-08, 2.431278e-08, 
    2.608036e-08, 2.766833e-08, 2.695676e-08, 2.645237e-08, 2.706674e-08, 
    2.689247e-08, 2.557777e-08, 2.588889e-08, 2.688561e-08, 3.022833e-08,
  2.472919e-08, 2.504127e-08, 2.501605e-08, 2.437873e-08, 2.383172e-08, 
    2.448767e-08, 2.675756e-08, 2.745294e-08, 2.699698e-08, 2.699371e-08, 
    2.716811e-08, 2.600705e-08, 2.599311e-08, 2.694879e-08, 3.070375e-08,
  2.437759e-08, 2.497642e-08, 2.504404e-08, 2.484808e-08, 2.396888e-08, 
    2.379814e-08, 2.522875e-08, 2.637495e-08, 2.717754e-08, 2.712296e-08, 
    2.683534e-08, 2.654325e-08, 2.602815e-08, 2.669662e-08, 2.964314e-08,
  2.393209e-08, 2.490342e-08, 2.511484e-08, 2.518174e-08, 2.469388e-08, 
    2.368627e-08, 2.410519e-08, 2.509796e-08, 2.613645e-08, 2.741183e-08, 
    2.715523e-08, 2.643022e-08, 2.611195e-08, 2.643276e-08, 2.772373e-08,
  2.411767e-08, 2.468128e-08, 2.485716e-08, 2.424688e-08, 2.413202e-08, 
    2.562423e-08, 2.743576e-08, 2.703685e-08, 2.63218e-08, 2.648681e-08, 
    2.722271e-08, 2.769114e-08, 2.641033e-08, 2.584819e-08, 2.652872e-08,
  2.458176e-08, 2.500935e-08, 2.467142e-08, 2.422848e-08, 2.432446e-08, 
    2.635353e-08, 2.736998e-08, 2.641239e-08, 2.63204e-08, 2.677645e-08, 
    2.740231e-08, 2.666949e-08, 2.57287e-08, 2.606165e-08, 2.669141e-08,
  2.47508e-08, 2.486622e-08, 2.462975e-08, 2.420874e-08, 2.441884e-08, 
    2.636029e-08, 2.680456e-08, 2.606084e-08, 2.652805e-08, 2.690963e-08, 
    2.715915e-08, 2.653544e-08, 2.56789e-08, 2.60201e-08, 2.772428e-08,
  2.481431e-08, 2.501568e-08, 2.479456e-08, 2.444611e-08, 2.435427e-08, 
    2.594865e-08, 2.627912e-08, 2.596902e-08, 2.688727e-08, 2.654991e-08, 
    2.697707e-08, 2.624359e-08, 2.595048e-08, 2.608285e-08, 2.712467e-08,
  2.486378e-08, 2.504461e-08, 2.483627e-08, 2.452937e-08, 2.445748e-08, 
    2.476876e-08, 2.595039e-08, 2.67655e-08, 2.660884e-08, 2.645604e-08, 
    2.712845e-08, 2.632236e-08, 2.622397e-08, 2.602581e-08, 2.7671e-08,
  2.497083e-08, 2.523356e-08, 2.51419e-08, 2.488903e-08, 2.466509e-08, 
    2.488626e-08, 2.518509e-08, 2.581431e-08, 2.643141e-08, 2.633834e-08, 
    2.688359e-08, 2.627907e-08, 2.585395e-08, 2.609765e-08, 2.758054e-08,
  2.522116e-08, 2.547005e-08, 2.544734e-08, 2.526911e-08, 2.505564e-08, 
    2.483822e-08, 2.511728e-08, 2.516711e-08, 2.576005e-08, 2.622407e-08, 
    2.708942e-08, 2.666786e-08, 2.611333e-08, 2.649609e-08, 2.824065e-08,
  2.563181e-08, 2.57622e-08, 2.590312e-08, 2.59038e-08, 2.566083e-08, 
    2.537206e-08, 2.531512e-08, 2.514156e-08, 2.549411e-08, 2.598143e-08, 
    2.634238e-08, 2.62308e-08, 2.609036e-08, 2.703677e-08, 2.879928e-08,
  2.611016e-08, 2.59799e-08, 2.606815e-08, 2.639985e-08, 2.628443e-08, 
    2.584247e-08, 2.56093e-08, 2.540092e-08, 2.521477e-08, 2.519671e-08, 
    2.545662e-08, 2.597347e-08, 2.567837e-08, 2.73571e-08, 2.894939e-08,
  2.689969e-08, 2.630452e-08, 2.608371e-08, 2.657571e-08, 2.681277e-08, 
    2.654077e-08, 2.629107e-08, 2.61125e-08, 2.555716e-08, 2.495887e-08, 
    2.414289e-08, 2.546468e-08, 2.590279e-08, 2.754132e-08, 2.854009e-08,
  2.545814e-08, 2.56156e-08, 2.587658e-08, 2.618894e-08, 2.630085e-08, 
    2.64315e-08, 2.653482e-08, 2.621958e-08, 2.610943e-08, 2.605734e-08, 
    2.636629e-08, 2.677212e-08, 2.694923e-08, 2.717266e-08, 2.689071e-08,
  2.580753e-08, 2.595981e-08, 2.642323e-08, 2.662112e-08, 2.685204e-08, 
    2.727635e-08, 2.696742e-08, 2.653603e-08, 2.653473e-08, 2.620421e-08, 
    2.642605e-08, 2.663392e-08, 2.710683e-08, 2.74657e-08, 2.637861e-08,
  2.613605e-08, 2.618608e-08, 2.649933e-08, 2.678166e-08, 2.726638e-08, 
    2.763308e-08, 2.703661e-08, 2.659946e-08, 2.640921e-08, 2.566011e-08, 
    2.580649e-08, 2.63705e-08, 2.704355e-08, 2.609341e-08, 2.612996e-08,
  2.653905e-08, 2.643948e-08, 2.67185e-08, 2.715754e-08, 2.738708e-08, 
    2.788559e-08, 2.650545e-08, 2.606404e-08, 2.620113e-08, 2.528784e-08, 
    2.53322e-08, 2.616586e-08, 2.657231e-08, 2.613254e-08, 2.697831e-08,
  2.708501e-08, 2.705643e-08, 2.741742e-08, 2.786964e-08, 2.77548e-08, 
    2.632801e-08, 2.716738e-08, 2.774439e-08, 2.647293e-08, 2.401961e-08, 
    2.474271e-08, 2.612375e-08, 2.669637e-08, 2.617476e-08, 2.688828e-08,
  2.792594e-08, 2.785731e-08, 2.832629e-08, 2.874871e-08, 2.771127e-08, 
    2.808475e-08, 2.843754e-08, 2.746082e-08, 2.575755e-08, 2.418713e-08, 
    2.467105e-08, 2.550406e-08, 2.585876e-08, 2.595564e-08, 2.736581e-08,
  2.888724e-08, 2.896489e-08, 2.88916e-08, 2.847791e-08, 2.777333e-08, 
    2.784133e-08, 2.858209e-08, 2.774975e-08, 2.604022e-08, 2.411434e-08, 
    2.454002e-08, 2.60602e-08, 2.594967e-08, 2.605847e-08, 2.815511e-08,
  2.996961e-08, 2.957434e-08, 2.872523e-08, 2.794449e-08, 2.774299e-08, 
    2.871598e-08, 2.829554e-08, 2.755374e-08, 2.600741e-08, 2.466141e-08, 
    2.478713e-08, 2.621694e-08, 2.652173e-08, 2.803943e-08, 2.850573e-08,
  3.091107e-08, 3.017e-08, 2.803409e-08, 2.698657e-08, 2.759266e-08, 
    2.861836e-08, 2.822771e-08, 2.745626e-08, 2.573886e-08, 2.465263e-08, 
    2.541478e-08, 2.693529e-08, 2.770649e-08, 2.857696e-08, 2.674914e-08,
  3.111682e-08, 3.017977e-08, 2.724408e-08, 2.588759e-08, 2.727471e-08, 
    2.895404e-08, 2.806313e-08, 2.697885e-08, 2.574953e-08, 2.544757e-08, 
    2.630205e-08, 2.769182e-08, 2.748129e-08, 2.598962e-08, 2.217705e-08,
  2.904424e-08, 2.913936e-08, 2.858479e-08, 2.880239e-08, 2.848067e-08, 
    2.98622e-08, 3.151138e-08, 3.187727e-08, 3.152891e-08, 3.053957e-08, 
    2.857754e-08, 2.674712e-08, 2.609904e-08, 2.649056e-08, 2.702715e-08,
  2.846445e-08, 2.824661e-08, 2.902999e-08, 2.930015e-08, 2.903935e-08, 
    3.154542e-08, 3.232158e-08, 3.21384e-08, 3.097715e-08, 2.982769e-08, 
    2.832052e-08, 2.629757e-08, 2.608893e-08, 2.722381e-08, 2.757105e-08,
  2.863339e-08, 2.895159e-08, 2.96939e-08, 2.880524e-08, 2.93249e-08, 
    2.835049e-08, 2.90871e-08, 3.002971e-08, 2.82908e-08, 2.762077e-08, 
    2.672923e-08, 2.559237e-08, 2.577839e-08, 2.671892e-08, 2.704841e-08,
  2.862051e-08, 2.933362e-08, 2.919569e-08, 2.850749e-08, 2.828605e-08, 
    2.568684e-08, 2.379937e-08, 2.279757e-08, 2.368923e-08, 2.496894e-08, 
    2.626326e-08, 2.569837e-08, 2.549778e-08, 2.675303e-08, 2.699404e-08,
  2.816321e-08, 2.866891e-08, 2.806541e-08, 2.768728e-08, 2.713569e-08, 
    2.552563e-08, 2.344714e-08, 2.345126e-08, 2.552366e-08, 2.451248e-08, 
    2.504622e-08, 2.491078e-08, 2.591486e-08, 2.643693e-08, 2.704004e-08,
  2.745192e-08, 2.679993e-08, 2.634703e-08, 2.653996e-08, 2.58976e-08, 
    2.64179e-08, 2.731914e-08, 2.596635e-08, 2.629971e-08, 2.69486e-08, 
    2.601726e-08, 2.430629e-08, 2.547279e-08, 2.675879e-08, 2.690367e-08,
  2.662757e-08, 2.513587e-08, 2.477483e-08, 2.55137e-08, 2.613098e-08, 
    2.647047e-08, 2.663256e-08, 2.666004e-08, 2.571241e-08, 2.404597e-08, 
    2.410459e-08, 2.500009e-08, 2.53715e-08, 2.624467e-08, 2.709275e-08,
  2.754874e-08, 2.411016e-08, 2.336375e-08, 2.467931e-08, 2.579018e-08, 
    2.632572e-08, 2.646107e-08, 2.629353e-08, 2.583905e-08, 2.520677e-08, 
    2.519111e-08, 2.551877e-08, 2.583182e-08, 2.654371e-08, 2.765087e-08,
  2.904766e-08, 2.483735e-08, 2.232677e-08, 2.35302e-08, 2.565301e-08, 
    2.607537e-08, 2.572757e-08, 2.635871e-08, 2.728334e-08, 2.731453e-08, 
    2.69126e-08, 2.652389e-08, 2.649099e-08, 2.695327e-08, 2.808614e-08,
  3.122967e-08, 2.763627e-08, 2.166324e-08, 2.166974e-08, 2.493879e-08, 
    2.611591e-08, 2.553186e-08, 2.534759e-08, 2.714925e-08, 2.80254e-08, 
    2.764662e-08, 2.707447e-08, 2.687901e-08, 2.696947e-08, 2.775663e-08,
  2.659456e-08, 2.66651e-08, 2.620145e-08, 2.55791e-08, 2.50619e-08, 
    2.507138e-08, 2.577161e-08, 2.664236e-08, 2.751289e-08, 2.796171e-08, 
    2.855149e-08, 2.931555e-08, 2.894937e-08, 2.851692e-08, 2.849441e-08,
  2.829598e-08, 2.843398e-08, 2.792118e-08, 2.61851e-08, 2.470925e-08, 
    2.404177e-08, 2.420841e-08, 2.524589e-08, 2.617723e-08, 2.689861e-08, 
    2.757781e-08, 2.916138e-08, 2.92252e-08, 2.854887e-08, 2.826039e-08,
  3.031017e-08, 3.073637e-08, 2.920687e-08, 2.594263e-08, 2.368195e-08, 
    2.215995e-08, 2.357859e-08, 2.493958e-08, 2.582013e-08, 2.58338e-08, 
    2.618476e-08, 2.805051e-08, 2.890649e-08, 2.800109e-08, 2.784797e-08,
  3.170878e-08, 3.153285e-08, 2.893423e-08, 2.47409e-08, 2.075859e-08, 
    2.156975e-08, 2.350309e-08, 2.343506e-08, 2.450844e-08, 2.359729e-08, 
    2.382443e-08, 2.669025e-08, 2.816939e-08, 2.772847e-08, 2.757653e-08,
  3.255721e-08, 3.205184e-08, 2.719204e-08, 2.090429e-08, 1.961527e-08, 
    2.208389e-08, 2.285221e-08, 2.409298e-08, 2.559008e-08, 2.344734e-08, 
    2.224828e-08, 2.515991e-08, 2.700083e-08, 2.722686e-08, 2.775163e-08,
  3.356743e-08, 3.226847e-08, 2.423955e-08, 1.880984e-08, 2.007238e-08, 
    2.399407e-08, 2.500725e-08, 2.531089e-08, 2.51705e-08, 2.593965e-08, 
    2.372183e-08, 2.509487e-08, 2.622687e-08, 2.732511e-08, 2.841229e-08,
  3.513449e-08, 3.27956e-08, 2.176775e-08, 1.869786e-08, 2.239818e-08, 
    2.53776e-08, 2.547832e-08, 2.597927e-08, 2.627222e-08, 2.5387e-08, 
    2.431089e-08, 2.531622e-08, 2.599209e-08, 2.813078e-08, 2.865634e-08,
  3.561674e-08, 3.238952e-08, 2.089671e-08, 1.936498e-08, 2.350941e-08, 
    2.541181e-08, 2.476618e-08, 2.597662e-08, 2.681592e-08, 2.52869e-08, 
    2.466939e-08, 2.533015e-08, 2.627576e-08, 2.850463e-08, 2.856322e-08,
  3.412699e-08, 3.324844e-08, 2.092601e-08, 2.010442e-08, 2.44568e-08, 
    2.505595e-08, 2.445556e-08, 2.675672e-08, 2.688662e-08, 2.458543e-08, 
    2.467791e-08, 2.548674e-08, 2.676375e-08, 2.879655e-08, 2.78858e-08,
  3.30294e-08, 3.272056e-08, 2.160957e-08, 2.039552e-08, 2.443068e-08, 
    2.515263e-08, 2.488841e-08, 2.586444e-08, 2.584144e-08, 2.503577e-08, 
    2.566537e-08, 2.606693e-08, 2.742659e-08, 2.856572e-08, 2.719148e-08,
  2.934158e-08, 2.978261e-08, 3.025422e-08, 3.155601e-08, 3.209646e-08, 
    3.243652e-08, 3.155021e-08, 3.027716e-08, 2.798515e-08, 2.654435e-08, 
    2.588815e-08, 2.55493e-08, 2.58392e-08, 2.578104e-08, 2.628015e-08,
  2.943602e-08, 2.979355e-08, 3.127646e-08, 3.36916e-08, 3.479567e-08, 
    3.498675e-08, 3.322817e-08, 3.013555e-08, 2.666846e-08, 2.419782e-08, 
    2.382652e-08, 2.429232e-08, 2.52e-08, 2.636547e-08, 2.71119e-08,
  2.941237e-08, 2.957111e-08, 3.167697e-08, 3.302967e-08, 3.33623e-08, 
    3.03384e-08, 2.843633e-08, 2.712744e-08, 2.411356e-08, 2.203224e-08, 
    2.200441e-08, 2.323407e-08, 2.50072e-08, 2.667932e-08, 2.770169e-08,
  2.901191e-08, 2.934268e-08, 3.006324e-08, 2.973862e-08, 2.556364e-08, 
    2.144446e-08, 1.992748e-08, 2.03149e-08, 2.160636e-08, 2.070491e-08, 
    2.123071e-08, 2.290473e-08, 2.536787e-08, 2.72915e-08, 2.79993e-08,
  2.86338e-08, 2.870537e-08, 2.864207e-08, 2.436858e-08, 2.225028e-08, 
    2.09656e-08, 2.021668e-08, 1.992975e-08, 2.156774e-08, 2.092009e-08, 
    2.114198e-08, 2.276676e-08, 2.624891e-08, 2.771568e-08, 2.795096e-08,
  2.710008e-08, 2.757925e-08, 2.490335e-08, 2.231851e-08, 2.213652e-08, 
    2.264785e-08, 2.393114e-08, 2.312615e-08, 2.199912e-08, 2.293727e-08, 
    2.297788e-08, 2.422787e-08, 2.703893e-08, 2.784653e-08, 2.804267e-08,
  2.638195e-08, 2.691356e-08, 2.40174e-08, 2.169924e-08, 2.319514e-08, 
    2.409485e-08, 2.467805e-08, 2.503915e-08, 2.319621e-08, 2.420727e-08, 
    2.384713e-08, 2.547572e-08, 2.780654e-08, 2.811063e-08, 2.814612e-08,
  2.606818e-08, 2.666083e-08, 2.205184e-08, 2.105502e-08, 2.405543e-08, 
    2.507455e-08, 2.466747e-08, 2.49638e-08, 2.442445e-08, 2.501153e-08, 
    2.4644e-08, 2.640224e-08, 2.827457e-08, 2.828351e-08, 2.807282e-08,
  2.61747e-08, 2.702643e-08, 2.111788e-08, 2.162698e-08, 2.574616e-08, 
    2.593427e-08, 2.569544e-08, 2.585316e-08, 2.529983e-08, 2.512299e-08, 
    2.535516e-08, 2.756546e-08, 2.82902e-08, 2.841138e-08, 2.782873e-08,
  2.607456e-08, 2.694591e-08, 2.10078e-08, 2.286206e-08, 2.663021e-08, 
    2.640367e-08, 2.614736e-08, 2.620751e-08, 2.503858e-08, 2.529042e-08, 
    2.662499e-08, 2.807812e-08, 2.859987e-08, 2.843401e-08, 2.716505e-08,
  2.870217e-08, 2.966751e-08, 2.972266e-08, 2.972065e-08, 2.902379e-08, 
    2.882634e-08, 2.882156e-08, 2.936768e-08, 3.027585e-08, 3.065734e-08, 
    3.036083e-08, 2.897625e-08, 2.723423e-08, 2.684678e-08, 2.814318e-08,
  3.006055e-08, 3.00661e-08, 2.988159e-08, 2.867359e-08, 2.868674e-08, 
    2.779017e-08, 2.80872e-08, 2.96665e-08, 3.180115e-08, 3.35025e-08, 
    3.279312e-08, 3.049768e-08, 2.706113e-08, 2.692132e-08, 2.77434e-08,
  2.979172e-08, 2.939081e-08, 2.842233e-08, 2.716488e-08, 2.72061e-08, 
    2.722233e-08, 2.581819e-08, 2.808791e-08, 3.09231e-08, 3.384542e-08, 
    3.356159e-08, 3.055098e-08, 2.683645e-08, 2.633144e-08, 2.707781e-08,
  2.93916e-08, 2.773279e-08, 2.602565e-08, 2.572291e-08, 2.529541e-08, 
    2.513819e-08, 2.478244e-08, 2.180393e-08, 2.783794e-08, 3.153043e-08, 
    3.141524e-08, 2.918001e-08, 2.588284e-08, 2.577892e-08, 2.66082e-08,
  2.618811e-08, 2.468071e-08, 2.448786e-08, 2.460342e-08, 2.48204e-08, 
    2.434567e-08, 2.363785e-08, 2.128906e-08, 2.299643e-08, 2.708762e-08, 
    2.753772e-08, 2.592832e-08, 2.469287e-08, 2.55163e-08, 2.661301e-08,
  2.405328e-08, 2.423767e-08, 2.494413e-08, 2.529277e-08, 2.475287e-08, 
    2.363811e-08, 2.35179e-08, 2.004322e-08, 1.941489e-08, 2.445726e-08, 
    2.467968e-08, 2.384658e-08, 2.377824e-08, 2.538791e-08, 2.641304e-08,
  2.411957e-08, 2.527253e-08, 2.567559e-08, 2.518444e-08, 2.389452e-08, 
    2.290209e-08, 2.31707e-08, 2.181816e-08, 2.106154e-08, 2.355447e-08, 
    2.277416e-08, 2.229104e-08, 2.352584e-08, 2.558528e-08, 2.661027e-08,
  2.526241e-08, 2.594721e-08, 2.577285e-08, 2.324703e-08, 2.190551e-08, 
    2.29125e-08, 2.33833e-08, 2.321831e-08, 2.248383e-08, 2.281584e-08, 
    2.179053e-08, 2.178829e-08, 2.420797e-08, 2.623319e-08, 2.696826e-08,
  2.555074e-08, 2.596233e-08, 2.400348e-08, 2.278827e-08, 2.333721e-08, 
    2.429724e-08, 2.423238e-08, 2.43466e-08, 2.321212e-08, 2.191287e-08, 
    2.163558e-08, 2.313517e-08, 2.567525e-08, 2.703718e-08, 2.75886e-08,
  2.55583e-08, 2.48085e-08, 2.350335e-08, 2.514384e-08, 2.568024e-08, 
    2.549385e-08, 2.493726e-08, 2.448828e-08, 2.270574e-08, 2.198543e-08, 
    2.362173e-08, 2.515577e-08, 2.673151e-08, 2.760668e-08, 2.775839e-08,
  2.855155e-08, 2.849008e-08, 2.897454e-08, 2.956652e-08, 3.049576e-08, 
    2.996656e-08, 2.980859e-08, 2.953555e-08, 2.992253e-08, 2.989064e-08, 
    2.948253e-08, 2.889457e-08, 2.846016e-08, 2.838487e-08, 2.909374e-08,
  2.877263e-08, 2.988227e-08, 3.043989e-08, 3.003908e-08, 2.933796e-08, 
    2.834932e-08, 2.745155e-08, 2.793995e-08, 2.782451e-08, 2.745525e-08, 
    2.784787e-08, 2.842621e-08, 2.810085e-08, 2.883213e-08, 2.964117e-08,
  3.0246e-08, 2.919967e-08, 2.824016e-08, 2.701333e-08, 2.662204e-08, 
    2.624801e-08, 2.523266e-08, 2.593697e-08, 2.629939e-08, 2.66504e-08, 
    2.734996e-08, 2.861557e-08, 2.878279e-08, 2.914686e-08, 3.000473e-08,
  2.878483e-08, 2.701514e-08, 2.546208e-08, 2.486672e-08, 2.382792e-08, 
    2.363973e-08, 2.381226e-08, 2.371103e-08, 2.49692e-08, 2.588664e-08, 
    2.831639e-08, 2.964461e-08, 2.904999e-08, 2.93092e-08, 2.857051e-08,
  2.594633e-08, 2.471382e-08, 2.441248e-08, 2.408611e-08, 2.403281e-08, 
    2.402654e-08, 2.355158e-08, 2.377315e-08, 2.536877e-08, 2.605395e-08, 
    2.934651e-08, 3.056812e-08, 2.972661e-08, 2.955539e-08, 2.826381e-08,
  2.492303e-08, 2.486958e-08, 2.517316e-08, 2.53313e-08, 2.551355e-08, 
    2.527892e-08, 2.473163e-08, 2.386393e-08, 2.290012e-08, 2.686383e-08, 
    3.077088e-08, 3.172344e-08, 2.981506e-08, 2.866769e-08, 2.802217e-08,
  2.603467e-08, 2.613261e-08, 2.618367e-08, 2.617914e-08, 2.61917e-08, 
    2.559578e-08, 2.472115e-08, 2.335477e-08, 2.27857e-08, 2.828222e-08, 
    3.22798e-08, 3.180298e-08, 2.927118e-08, 2.829089e-08, 2.861287e-08,
  2.65442e-08, 2.606068e-08, 2.591652e-08, 2.578426e-08, 2.512234e-08, 
    2.482321e-08, 2.409323e-08, 2.22231e-08, 2.301374e-08, 2.98541e-08, 
    3.232405e-08, 3.080361e-08, 2.798966e-08, 2.778255e-08, 2.851856e-08,
  2.507052e-08, 2.473519e-08, 2.385683e-08, 2.330377e-08, 2.344402e-08, 
    2.374289e-08, 2.307307e-08, 2.199352e-08, 2.455175e-08, 2.966668e-08, 
    3.107449e-08, 2.89317e-08, 2.711599e-08, 2.785425e-08, 2.890163e-08,
  2.359226e-08, 2.378121e-08, 2.34996e-08, 2.301386e-08, 2.280269e-08, 
    2.300999e-08, 2.225462e-08, 2.260346e-08, 2.573716e-08, 2.902022e-08, 
    2.939565e-08, 2.750205e-08, 2.663771e-08, 2.785254e-08, 2.876937e-08,
  2.889447e-08, 2.946099e-08, 2.948122e-08, 2.913713e-08, 2.894245e-08, 
    2.873388e-08, 2.837429e-08, 2.824159e-08, 2.804653e-08, 2.811549e-08, 
    2.804579e-08, 2.83875e-08, 2.77758e-08, 2.806052e-08, 2.763742e-08,
  2.942114e-08, 2.933021e-08, 2.993943e-08, 2.863697e-08, 2.904061e-08, 
    2.756931e-08, 2.715684e-08, 2.744139e-08, 2.70661e-08, 2.694379e-08, 
    2.704277e-08, 2.782489e-08, 2.80901e-08, 2.83444e-08, 2.822602e-08,
  2.959203e-08, 2.96507e-08, 2.927223e-08, 2.869775e-08, 2.880777e-08, 
    2.839491e-08, 2.800469e-08, 2.676764e-08, 2.522409e-08, 2.536652e-08, 
    2.601187e-08, 2.721731e-08, 2.885266e-08, 2.864058e-08, 2.851922e-08,
  2.952519e-08, 2.894064e-08, 2.866379e-08, 2.847532e-08, 2.70744e-08, 
    2.678701e-08, 2.616131e-08, 2.233978e-08, 2.255731e-08, 2.411454e-08, 
    2.640224e-08, 2.826488e-08, 2.958998e-08, 2.91645e-08, 2.86696e-08,
  2.942324e-08, 2.945208e-08, 2.91619e-08, 2.789877e-08, 2.684824e-08, 
    2.573716e-08, 2.282546e-08, 2.172566e-08, 2.491933e-08, 2.641605e-08, 
    2.725233e-08, 2.905838e-08, 2.971147e-08, 2.915979e-08, 2.838757e-08,
  2.994542e-08, 2.92392e-08, 2.782163e-08, 2.655014e-08, 2.602724e-08, 
    2.597598e-08, 2.561013e-08, 2.321432e-08, 2.424355e-08, 2.775227e-08, 
    2.814606e-08, 2.990926e-08, 3.001757e-08, 2.893537e-08, 2.613626e-08,
  2.891485e-08, 2.739882e-08, 2.614285e-08, 2.585623e-08, 2.631405e-08, 
    2.611552e-08, 2.478133e-08, 2.400352e-08, 2.654224e-08, 2.827568e-08, 
    2.896185e-08, 3.039634e-08, 2.895244e-08, 2.658858e-08, 2.662057e-08,
  2.72875e-08, 2.576508e-08, 2.465214e-08, 2.562317e-08, 2.61189e-08, 
    2.500142e-08, 2.401767e-08, 2.505629e-08, 2.765462e-08, 2.913671e-08, 
    3.007081e-08, 2.991512e-08, 2.714795e-08, 2.740286e-08, 2.924014e-08,
  2.469552e-08, 2.377833e-08, 2.380422e-08, 2.563079e-08, 2.545305e-08, 
    2.445806e-08, 2.473131e-08, 2.691779e-08, 2.869865e-08, 3.023162e-08, 
    3.014537e-08, 2.782928e-08, 2.710054e-08, 2.912797e-08, 3.185529e-08,
  2.347327e-08, 2.352022e-08, 2.395217e-08, 2.469949e-08, 2.454456e-08, 
    2.46047e-08, 2.610506e-08, 2.823624e-08, 2.991622e-08, 3.063871e-08, 
    2.872584e-08, 2.727076e-08, 2.889429e-08, 3.237711e-08, 3.323159e-08,
  2.772364e-08, 2.809575e-08, 2.907119e-08, 2.936837e-08, 3.041101e-08, 
    3.099224e-08, 3.137781e-08, 3.112199e-08, 3.000009e-08, 2.924699e-08, 
    2.797658e-08, 2.740169e-08, 2.644898e-08, 2.603752e-08, 2.652647e-08,
  2.825991e-08, 2.863036e-08, 2.949402e-08, 2.987665e-08, 3.18282e-08, 
    3.153355e-08, 3.100023e-08, 3.046711e-08, 2.886645e-08, 2.774734e-08, 
    2.66317e-08, 2.524401e-08, 2.457114e-08, 2.498427e-08, 2.552561e-08,
  2.853026e-08, 2.928924e-08, 3.000234e-08, 3.195329e-08, 3.233101e-08, 
    3.167285e-08, 3.053606e-08, 2.899193e-08, 2.772183e-08, 2.588117e-08, 
    2.431642e-08, 2.352762e-08, 2.348427e-08, 2.410142e-08, 2.538176e-08,
  2.823513e-08, 2.915758e-08, 3.083002e-08, 3.231795e-08, 3.044575e-08, 
    3.021384e-08, 2.847473e-08, 2.708255e-08, 2.529382e-08, 2.423973e-08, 
    2.377414e-08, 2.407774e-08, 2.506626e-08, 2.546425e-08, 2.604122e-08,
  2.89669e-08, 3.043575e-08, 3.201304e-08, 3.073149e-08, 2.927573e-08, 
    2.72793e-08, 2.671063e-08, 2.735274e-08, 2.507273e-08, 2.446821e-08, 
    2.544923e-08, 2.715264e-08, 2.758385e-08, 2.733437e-08, 2.724613e-08,
  2.975701e-08, 3.04151e-08, 2.990624e-08, 2.808251e-08, 2.664533e-08, 
    2.646535e-08, 2.589061e-08, 2.553248e-08, 2.575924e-08, 2.714057e-08, 
    2.848235e-08, 2.961731e-08, 2.89206e-08, 2.80995e-08, 2.798856e-08,
  2.919691e-08, 2.924697e-08, 2.779102e-08, 2.615516e-08, 2.585881e-08, 
    2.591959e-08, 2.611687e-08, 2.621263e-08, 2.78404e-08, 2.909647e-08, 
    2.971859e-08, 2.994551e-08, 2.813941e-08, 2.791935e-08, 2.734235e-08,
  2.832767e-08, 2.706733e-08, 2.567593e-08, 2.529267e-08, 2.53793e-08, 
    2.585292e-08, 2.610779e-08, 2.776755e-08, 2.79529e-08, 2.801957e-08, 
    2.810932e-08, 2.706738e-08, 2.707772e-08, 2.719954e-08, 2.677485e-08,
  2.701093e-08, 2.559779e-08, 2.495186e-08, 2.509642e-08, 2.500616e-08, 
    2.716395e-08, 2.822739e-08, 2.80155e-08, 2.778051e-08, 2.704515e-08, 
    2.66206e-08, 2.651985e-08, 2.734956e-08, 2.715968e-08, 2.752189e-08,
  2.482588e-08, 2.43889e-08, 2.436645e-08, 2.45631e-08, 2.651651e-08, 
    2.844662e-08, 2.852554e-08, 2.825154e-08, 2.820359e-08, 2.734923e-08, 
    2.772508e-08, 2.765763e-08, 2.80831e-08, 2.817768e-08, 2.867667e-08,
  2.875948e-08, 2.848266e-08, 2.822021e-08, 2.795456e-08, 2.731373e-08, 
    2.737894e-08, 2.749126e-08, 2.803646e-08, 2.83964e-08, 2.839086e-08, 
    2.813836e-08, 2.807258e-08, 2.872503e-08, 2.876726e-08, 2.780268e-08,
  2.897224e-08, 2.85633e-08, 2.831875e-08, 2.775405e-08, 2.732901e-08, 
    2.765627e-08, 2.771492e-08, 2.798192e-08, 2.854996e-08, 2.798122e-08, 
    2.783532e-08, 2.822895e-08, 2.894099e-08, 2.8329e-08, 2.750319e-08,
  2.857705e-08, 2.803287e-08, 2.762671e-08, 2.709007e-08, 2.739387e-08, 
    2.813127e-08, 2.825712e-08, 2.841442e-08, 2.829235e-08, 2.822726e-08, 
    2.834021e-08, 2.884263e-08, 2.879065e-08, 2.821203e-08, 2.760598e-08,
  2.8286e-08, 2.805839e-08, 2.751594e-08, 2.760396e-08, 2.794523e-08, 
    2.790891e-08, 2.789987e-08, 2.875985e-08, 2.906155e-08, 2.94526e-08, 
    2.935561e-08, 2.949789e-08, 2.918891e-08, 2.84453e-08, 2.737837e-08,
  2.841718e-08, 2.79178e-08, 2.816373e-08, 2.821126e-08, 2.824334e-08, 
    2.737191e-08, 2.825028e-08, 2.920358e-08, 2.932122e-08, 2.848533e-08, 
    2.83542e-08, 2.865313e-08, 2.835833e-08, 2.818776e-08, 2.722626e-08,
  2.85368e-08, 2.851209e-08, 2.857638e-08, 2.835703e-08, 2.739701e-08, 
    2.782149e-08, 2.788136e-08, 2.779362e-08, 2.788897e-08, 2.85625e-08, 
    2.924661e-08, 2.906585e-08, 2.86769e-08, 2.80125e-08, 2.764671e-08,
  2.836044e-08, 2.82344e-08, 2.810392e-08, 2.747984e-08, 2.749008e-08, 
    2.7626e-08, 2.813695e-08, 2.794239e-08, 2.806589e-08, 2.880751e-08, 
    2.828095e-08, 2.766026e-08, 2.751674e-08, 2.734828e-08, 2.740087e-08,
  2.839201e-08, 2.799431e-08, 2.766823e-08, 2.749582e-08, 2.725126e-08, 
    2.71879e-08, 2.736539e-08, 2.873908e-08, 3.060775e-08, 2.914786e-08, 
    2.73204e-08, 2.741291e-08, 2.787128e-08, 2.771828e-08, 2.7409e-08,
  2.891534e-08, 2.806327e-08, 2.771738e-08, 2.726113e-08, 2.676652e-08, 
    2.606675e-08, 2.770533e-08, 3.172029e-08, 3.138859e-08, 2.811795e-08, 
    2.655777e-08, 2.736179e-08, 2.765822e-08, 2.74362e-08, 2.736705e-08,
  2.843191e-08, 2.756457e-08, 2.714635e-08, 2.597279e-08, 2.535091e-08, 
    2.604052e-08, 3.165732e-08, 3.469806e-08, 3.166988e-08, 2.71209e-08, 
    2.666266e-08, 2.691391e-08, 2.731509e-08, 2.666937e-08, 2.744376e-08,
  2.883253e-08, 2.891858e-08, 2.913035e-08, 2.930309e-08, 2.944237e-08, 
    2.958614e-08, 2.971395e-08, 2.958318e-08, 2.961971e-08, 2.935232e-08, 
    2.931204e-08, 2.8777e-08, 2.836469e-08, 2.827538e-08, 2.81954e-08,
  2.914551e-08, 2.913331e-08, 2.943292e-08, 2.961948e-08, 3.004514e-08, 
    2.997444e-08, 2.991044e-08, 2.951645e-08, 2.944023e-08, 2.910716e-08, 
    2.897373e-08, 2.862027e-08, 2.850833e-08, 2.853229e-08, 2.805099e-08,
  2.92471e-08, 2.94385e-08, 2.980738e-08, 3.026165e-08, 3.027417e-08, 
    2.94061e-08, 2.920669e-08, 2.92461e-08, 2.900488e-08, 2.90058e-08, 
    2.881584e-08, 2.88344e-08, 2.867505e-08, 2.824317e-08, 2.753887e-08,
  2.948465e-08, 2.988634e-08, 3.041559e-08, 3.048823e-08, 2.971782e-08, 
    2.984898e-08, 2.912436e-08, 2.91755e-08, 2.926566e-08, 2.894776e-08, 
    2.876742e-08, 2.870962e-08, 2.856008e-08, 2.814556e-08, 2.800777e-08,
  3.020652e-08, 3.048149e-08, 3.058092e-08, 2.988252e-08, 2.948117e-08, 
    2.954591e-08, 2.946138e-08, 2.86352e-08, 2.833529e-08, 2.858545e-08, 
    2.834476e-08, 2.823739e-08, 2.805923e-08, 2.800039e-08, 2.758278e-08,
  3.045965e-08, 3.038353e-08, 2.985936e-08, 2.926778e-08, 2.962835e-08, 
    2.922273e-08, 2.850864e-08, 2.840886e-08, 2.784903e-08, 2.831939e-08, 
    2.847307e-08, 2.853587e-08, 2.871746e-08, 2.886426e-08, 2.826767e-08,
  3.018399e-08, 2.963382e-08, 2.919602e-08, 2.913444e-08, 2.89042e-08, 
    2.836044e-08, 2.828947e-08, 2.792995e-08, 2.764693e-08, 2.853401e-08, 
    2.844379e-08, 2.945528e-08, 2.892808e-08, 2.859524e-08, 2.80821e-08,
  2.938884e-08, 2.891607e-08, 2.873706e-08, 2.866709e-08, 2.830217e-08, 
    2.755855e-08, 2.779803e-08, 2.670925e-08, 2.869553e-08, 2.908875e-08, 
    3.002853e-08, 2.952816e-08, 2.957101e-08, 2.881701e-08, 2.890994e-08,
  2.86514e-08, 2.927744e-08, 2.876361e-08, 2.859566e-08, 2.768951e-08, 
    2.704668e-08, 2.74146e-08, 2.935729e-08, 3.082062e-08, 3.104069e-08, 
    3.020491e-08, 2.964296e-08, 2.947299e-08, 2.932901e-08, 2.902434e-08,
  2.929142e-08, 2.875821e-08, 2.811456e-08, 2.817128e-08, 2.679458e-08, 
    2.729906e-08, 2.933699e-08, 3.041739e-08, 3.078268e-08, 2.819591e-08, 
    2.799575e-08, 2.854637e-08, 2.882959e-08, 2.895671e-08, 2.849773e-08,
  2.961516e-08, 3.013898e-08, 3.025662e-08, 3.039899e-08, 3.000875e-08, 
    2.977895e-08, 2.955526e-08, 2.965701e-08, 2.954734e-08, 2.962597e-08, 
    2.980855e-08, 2.998736e-08, 3.013353e-08, 2.978999e-08, 2.965227e-08,
  3.103478e-08, 3.052613e-08, 3.015459e-08, 2.952994e-08, 2.953349e-08, 
    2.935824e-08, 2.914019e-08, 2.932867e-08, 2.94946e-08, 2.95326e-08, 
    2.994717e-08, 3.004538e-08, 2.995214e-08, 2.956494e-08, 2.979757e-08,
  2.917798e-08, 2.911713e-08, 2.869374e-08, 2.841032e-08, 2.904195e-08, 
    2.939202e-08, 2.894792e-08, 2.892508e-08, 2.960009e-08, 2.954639e-08, 
    2.997663e-08, 2.971782e-08, 2.95046e-08, 2.978912e-08, 3.00169e-08,
  2.757409e-08, 2.743379e-08, 2.775611e-08, 2.806348e-08, 2.8694e-08, 
    2.938806e-08, 2.940877e-08, 3.003848e-08, 3.006964e-08, 3.015799e-08, 
    2.991229e-08, 2.92634e-08, 2.955138e-08, 2.980022e-08, 3.020332e-08,
  2.553095e-08, 2.590597e-08, 2.664999e-08, 2.725244e-08, 2.810853e-08, 
    2.817686e-08, 2.975512e-08, 3.046053e-08, 3.111658e-08, 2.920457e-08, 
    2.781352e-08, 2.815915e-08, 2.891077e-08, 2.969315e-08, 3.014839e-08,
  2.480921e-08, 2.53116e-08, 2.58027e-08, 2.700951e-08, 2.76673e-08, 
    2.926262e-08, 2.834308e-08, 2.836462e-08, 2.80978e-08, 2.711534e-08, 
    2.723791e-08, 2.785885e-08, 2.853752e-08, 2.906956e-08, 2.922235e-08,
  2.399391e-08, 2.448547e-08, 2.553655e-08, 2.687416e-08, 2.809054e-08, 
    2.841091e-08, 2.844923e-08, 2.774248e-08, 2.692522e-08, 2.649111e-08, 
    2.718514e-08, 2.920763e-08, 2.929563e-08, 2.877715e-08, 2.857529e-08,
  2.497561e-08, 2.534352e-08, 2.656988e-08, 2.784415e-08, 2.868292e-08, 
    2.879365e-08, 2.809929e-08, 2.832718e-08, 2.765034e-08, 2.723757e-08, 
    2.681622e-08, 2.892937e-08, 2.945524e-08, 2.84447e-08, 2.828078e-08,
  2.534318e-08, 2.68287e-08, 2.801991e-08, 2.884437e-08, 2.94423e-08, 
    2.84969e-08, 2.849401e-08, 2.810576e-08, 2.827086e-08, 2.84849e-08, 
    2.77749e-08, 2.912494e-08, 2.908585e-08, 2.812156e-08, 2.780954e-08,
  2.767303e-08, 2.87489e-08, 2.890816e-08, 3.003089e-08, 2.888033e-08, 
    2.806248e-08, 2.782308e-08, 2.76926e-08, 2.931958e-08, 2.893935e-08, 
    2.86317e-08, 2.961121e-08, 2.890182e-08, 2.785416e-08, 2.766905e-08,
  3.107975e-08, 2.980567e-08, 2.923522e-08, 2.930911e-08, 2.897795e-08, 
    2.911547e-08, 2.902691e-08, 2.945728e-08, 3.010556e-08, 3.036167e-08, 
    3.002906e-08, 2.927415e-08, 2.932791e-08, 2.97746e-08, 3.013064e-08,
  2.886677e-08, 2.786716e-08, 2.790224e-08, 2.81073e-08, 2.806864e-08, 
    2.878904e-08, 2.936891e-08, 3.040852e-08, 3.112416e-08, 3.068497e-08, 
    2.999542e-08, 2.965909e-08, 2.965947e-08, 3.005952e-08, 2.943369e-08,
  2.650586e-08, 2.595626e-08, 2.6575e-08, 2.628559e-08, 2.704218e-08, 
    2.707246e-08, 2.813802e-08, 2.924061e-08, 3.01199e-08, 3.010699e-08, 
    2.993848e-08, 2.979656e-08, 2.96108e-08, 2.897012e-08, 2.889885e-08,
  2.605609e-08, 2.615913e-08, 2.56445e-08, 2.588204e-08, 2.52602e-08, 
    2.623874e-08, 2.621021e-08, 2.753312e-08, 2.754421e-08, 2.793545e-08, 
    2.910694e-08, 2.937255e-08, 2.904467e-08, 2.825693e-08, 2.81037e-08,
  2.596607e-08, 2.586527e-08, 2.568366e-08, 2.5444e-08, 2.525857e-08, 
    2.487413e-08, 2.530219e-08, 2.63282e-08, 2.704684e-08, 2.777269e-08, 
    2.861616e-08, 2.81334e-08, 2.723294e-08, 2.702892e-08, 2.818113e-08,
  2.63895e-08, 2.658848e-08, 2.632279e-08, 2.552841e-08, 2.507106e-08, 
    2.396698e-08, 2.406509e-08, 2.396808e-08, 2.46174e-08, 2.701735e-08, 
    2.711062e-08, 2.549353e-08, 2.531661e-08, 2.648651e-08, 2.915842e-08,
  2.732535e-08, 2.731606e-08, 2.659818e-08, 2.56698e-08, 2.499175e-08, 
    2.405559e-08, 2.384428e-08, 2.434637e-08, 2.576376e-08, 2.576413e-08, 
    2.52507e-08, 2.522848e-08, 2.587385e-08, 2.789696e-08, 2.923959e-08,
  2.806695e-08, 2.780531e-08, 2.715582e-08, 2.707374e-08, 2.675553e-08, 
    2.708229e-08, 2.687679e-08, 2.702579e-08, 2.675934e-08, 2.686886e-08, 
    2.625583e-08, 2.566365e-08, 2.713901e-08, 2.896182e-08, 2.810854e-08,
  2.805552e-08, 2.781521e-08, 2.79921e-08, 2.801257e-08, 2.840775e-08, 
    2.857819e-08, 2.822984e-08, 2.819037e-08, 2.787378e-08, 2.80555e-08, 
    2.681196e-08, 2.712429e-08, 2.829487e-08, 2.869476e-08, 2.660364e-08,
  2.79744e-08, 2.843196e-08, 2.844131e-08, 2.829963e-08, 2.816146e-08, 
    2.810448e-08, 2.832134e-08, 2.74017e-08, 2.840348e-08, 2.821627e-08, 
    2.715281e-08, 2.852828e-08, 2.875502e-08, 2.803509e-08, 2.715975e-08,
  3.242571e-08, 3.193747e-08, 3.061869e-08, 2.986565e-08, 2.960266e-08, 
    2.862021e-08, 2.66892e-08, 2.523348e-08, 2.664365e-08, 2.79192e-08, 
    2.857298e-08, 2.935374e-08, 2.987832e-08, 3.153406e-08, 3.109249e-08,
  3.207869e-08, 3.10784e-08, 3.021437e-08, 2.968038e-08, 2.974023e-08, 
    2.847826e-08, 2.681955e-08, 2.604507e-08, 2.665013e-08, 2.792048e-08, 
    2.968464e-08, 3.096623e-08, 3.135208e-08, 3.099203e-08, 3.098612e-08,
  3.11969e-08, 3.075514e-08, 2.995916e-08, 2.928802e-08, 2.9518e-08, 
    2.83292e-08, 2.588635e-08, 2.599591e-08, 2.739979e-08, 2.94314e-08, 
    3.222992e-08, 3.228097e-08, 3.181928e-08, 3.154264e-08, 3.080028e-08,
  3.125262e-08, 3.04102e-08, 2.984354e-08, 2.900572e-08, 2.841159e-08, 
    2.829444e-08, 2.696866e-08, 2.663496e-08, 2.708161e-08, 2.792532e-08, 
    3.162649e-08, 3.21082e-08, 3.219513e-08, 2.966356e-08, 2.880088e-08,
  3.075166e-08, 3.024804e-08, 2.957548e-08, 2.843108e-08, 2.848918e-08, 
    2.806113e-08, 2.732754e-08, 2.446318e-08, 2.789536e-08, 2.986564e-08, 
    2.930292e-08, 2.99911e-08, 2.847185e-08, 2.728631e-08, 2.62462e-08,
  3.050181e-08, 2.98206e-08, 2.890759e-08, 2.846579e-08, 2.849649e-08, 
    2.832629e-08, 2.716513e-08, 2.71432e-08, 2.481779e-08, 2.719457e-08, 
    2.810916e-08, 2.774283e-08, 2.687708e-08, 2.619853e-08, 2.766524e-08,
  3.013817e-08, 2.941312e-08, 2.88565e-08, 2.808846e-08, 2.828739e-08, 
    2.833522e-08, 2.743256e-08, 2.659133e-08, 2.447005e-08, 2.532618e-08, 
    2.701828e-08, 2.712134e-08, 2.612023e-08, 2.693643e-08, 2.904871e-08,
  2.941659e-08, 2.904075e-08, 2.795892e-08, 2.824844e-08, 2.832458e-08, 
    2.804114e-08, 2.843629e-08, 2.670766e-08, 2.391769e-08, 2.464542e-08, 
    2.61571e-08, 2.59111e-08, 2.641541e-08, 2.845351e-08, 2.863687e-08,
  2.863e-08, 2.859627e-08, 2.846707e-08, 2.793471e-08, 2.761356e-08, 
    2.809577e-08, 2.848428e-08, 2.754772e-08, 2.497321e-08, 2.47392e-08, 
    2.608473e-08, 2.577223e-08, 2.699517e-08, 2.740048e-08, 2.634153e-08,
  2.877566e-08, 2.931852e-08, 2.754232e-08, 2.637521e-08, 2.675009e-08, 
    2.741649e-08, 2.851536e-08, 2.777896e-08, 2.541722e-08, 2.527258e-08, 
    2.590102e-08, 2.62037e-08, 2.667853e-08, 2.603914e-08, 2.651831e-08,
  3.090186e-08, 3.084597e-08, 3.149239e-08, 3.1587e-08, 3.154898e-08, 
    3.01415e-08, 2.9082e-08, 2.87128e-08, 2.84684e-08, 2.781021e-08, 
    2.90199e-08, 3.043368e-08, 3.008921e-08, 3.036541e-08, 3.028191e-08,
  3.074487e-08, 3.154684e-08, 3.176997e-08, 3.152718e-08, 3.135412e-08, 
    2.998398e-08, 2.899598e-08, 2.850578e-08, 2.811155e-08, 2.761756e-08, 
    2.920516e-08, 2.96697e-08, 2.916644e-08, 2.991172e-08, 2.992793e-08,
  3.116529e-08, 3.216935e-08, 3.16607e-08, 3.099876e-08, 3.060405e-08, 
    2.99321e-08, 2.866322e-08, 2.809945e-08, 2.800086e-08, 2.767651e-08, 
    2.893572e-08, 2.895913e-08, 2.832408e-08, 2.821102e-08, 2.849916e-08,
  3.242257e-08, 3.214101e-08, 3.10666e-08, 3.060524e-08, 3.008103e-08, 
    2.965489e-08, 2.852209e-08, 2.778162e-08, 2.785676e-08, 2.765628e-08, 
    2.844867e-08, 2.802285e-08, 2.762368e-08, 2.731309e-08, 2.730228e-08,
  3.261398e-08, 3.147707e-08, 3.036989e-08, 3.054789e-08, 3.003302e-08, 
    2.800575e-08, 2.757463e-08, 2.756971e-08, 2.63439e-08, 2.786444e-08, 
    2.807325e-08, 2.754635e-08, 2.734867e-08, 2.767598e-08, 2.759215e-08,
  3.214252e-08, 3.035813e-08, 3.033472e-08, 3.062773e-08, 2.882064e-08, 
    2.793447e-08, 2.66829e-08, 2.79017e-08, 2.965426e-08, 2.786517e-08, 
    2.762053e-08, 2.699925e-08, 2.687601e-08, 2.642286e-08, 2.678228e-08,
  3.117754e-08, 2.998848e-08, 3.094895e-08, 2.947318e-08, 2.799905e-08, 
    2.66646e-08, 2.64661e-08, 2.806663e-08, 2.811755e-08, 2.644308e-08, 
    2.774412e-08, 2.713126e-08, 2.695513e-08, 2.549265e-08, 2.424946e-08,
  2.989736e-08, 2.987584e-08, 3.053708e-08, 2.8359e-08, 2.682586e-08, 
    2.617073e-08, 2.681757e-08, 2.871228e-08, 2.700427e-08, 2.662504e-08, 
    2.778436e-08, 2.807514e-08, 2.844775e-08, 2.762579e-08, 2.633091e-08,
  2.917229e-08, 3.068335e-08, 3.005749e-08, 2.72301e-08, 2.635599e-08, 
    2.603638e-08, 2.768569e-08, 2.88291e-08, 2.607625e-08, 2.693379e-08, 
    2.821698e-08, 2.862755e-08, 2.926059e-08, 2.920394e-08, 2.848721e-08,
  2.900853e-08, 3.080405e-08, 2.860644e-08, 2.688678e-08, 2.67864e-08, 
    2.655993e-08, 2.837412e-08, 2.795506e-08, 2.608386e-08, 2.742875e-08, 
    2.829344e-08, 2.821985e-08, 2.816689e-08, 2.762962e-08, 2.651949e-08,
  2.885762e-08, 2.871125e-08, 3.086355e-08, 3.267009e-08, 3.592763e-08, 
    3.39604e-08, 3.070691e-08, 2.93274e-08, 2.754535e-08, 2.732026e-08, 
    2.700455e-08, 2.663618e-08, 2.681181e-08, 2.737699e-08, 2.824193e-08,
  2.772418e-08, 2.998891e-08, 3.233909e-08, 3.50738e-08, 3.49746e-08, 
    3.260402e-08, 2.972639e-08, 2.821002e-08, 2.726011e-08, 2.735534e-08, 
    2.720908e-08, 2.635957e-08, 2.64253e-08, 2.681621e-08, 2.786215e-08,
  2.817605e-08, 3.239694e-08, 3.448954e-08, 3.508785e-08, 3.341414e-08, 
    3.099741e-08, 2.87339e-08, 2.732742e-08, 2.700643e-08, 2.792244e-08, 
    2.699467e-08, 2.617544e-08, 2.612955e-08, 2.664941e-08, 2.684038e-08,
  3.073706e-08, 3.497483e-08, 3.459253e-08, 3.391849e-08, 3.13104e-08, 
    2.954e-08, 2.81103e-08, 2.67527e-08, 2.680616e-08, 2.835173e-08, 
    2.724392e-08, 2.563636e-08, 2.538821e-08, 2.560336e-08, 2.612204e-08,
  3.429821e-08, 3.540452e-08, 3.326048e-08, 3.254209e-08, 2.997889e-08, 
    2.785938e-08, 2.801223e-08, 2.690056e-08, 2.771568e-08, 2.8862e-08, 
    2.735463e-08, 2.590574e-08, 2.535297e-08, 2.540313e-08, 2.546577e-08,
  3.516579e-08, 3.354349e-08, 3.284122e-08, 3.115141e-08, 2.839184e-08, 
    2.826766e-08, 2.663393e-08, 2.877143e-08, 2.994225e-08, 2.804697e-08, 
    2.776849e-08, 2.643362e-08, 2.577436e-08, 2.509561e-08, 2.52851e-08,
  3.442253e-08, 3.25676e-08, 3.159325e-08, 2.922493e-08, 2.812571e-08, 
    2.741196e-08, 2.769966e-08, 2.709216e-08, 2.764409e-08, 2.833708e-08, 
    2.797302e-08, 2.732596e-08, 2.707598e-08, 2.620445e-08, 2.558493e-08,
  3.330357e-08, 3.141479e-08, 3.023467e-08, 2.856745e-08, 2.791853e-08, 
    2.768396e-08, 2.747992e-08, 2.840244e-08, 2.81201e-08, 2.797369e-08, 
    2.763001e-08, 2.744576e-08, 2.748149e-08, 2.676807e-08, 2.672589e-08,
  3.195424e-08, 3.029528e-08, 2.957422e-08, 2.786484e-08, 2.802397e-08, 
    2.750274e-08, 2.758584e-08, 2.755457e-08, 2.799717e-08, 2.754751e-08, 
    2.682644e-08, 2.689094e-08, 2.709109e-08, 2.670724e-08, 2.708673e-08,
  3.068753e-08, 2.952386e-08, 2.903311e-08, 2.797834e-08, 2.792789e-08, 
    2.713333e-08, 2.744555e-08, 2.779725e-08, 2.77799e-08, 2.667501e-08, 
    2.623212e-08, 2.66409e-08, 2.719765e-08, 2.707865e-08, 2.757711e-08,
  2.523895e-08, 2.584821e-08, 2.772914e-08, 3.066388e-08, 3.214042e-08, 
    3.173944e-08, 2.996642e-08, 2.866211e-08, 2.85126e-08, 2.81922e-08, 
    2.709373e-08, 2.748929e-08, 2.780586e-08, 2.658918e-08, 2.61852e-08,
  2.508323e-08, 2.665322e-08, 2.896454e-08, 3.14719e-08, 3.224971e-08, 
    3.11669e-08, 2.953581e-08, 2.822394e-08, 2.847937e-08, 2.776027e-08, 
    2.699612e-08, 2.782527e-08, 2.772327e-08, 2.671488e-08, 2.607618e-08,
  2.621366e-08, 2.858625e-08, 2.98926e-08, 3.133678e-08, 3.191258e-08, 
    3.082141e-08, 2.847846e-08, 2.835628e-08, 2.859317e-08, 2.70269e-08, 
    2.668901e-08, 2.794165e-08, 2.73749e-08, 2.665587e-08, 2.62402e-08,
  2.842356e-08, 2.941684e-08, 3.014064e-08, 3.217088e-08, 3.10169e-08, 
    3.026582e-08, 2.777054e-08, 2.883662e-08, 2.863076e-08, 2.622095e-08, 
    2.681753e-08, 2.789225e-08, 2.72052e-08, 2.621377e-08, 2.543567e-08,
  2.965903e-08, 2.95965e-08, 3.151412e-08, 3.184137e-08, 3.049738e-08, 
    2.860516e-08, 2.753737e-08, 2.919694e-08, 2.800495e-08, 2.52532e-08, 
    2.680555e-08, 2.784327e-08, 2.707681e-08, 2.619409e-08, 2.519735e-08,
  2.952956e-08, 3.005358e-08, 3.202515e-08, 3.132234e-08, 2.969909e-08, 
    2.83762e-08, 2.728516e-08, 2.822229e-08, 2.719492e-08, 2.600383e-08, 
    2.695209e-08, 2.775615e-08, 2.677329e-08, 2.57219e-08, 2.477782e-08,
  2.983753e-08, 3.151092e-08, 3.22151e-08, 3.021147e-08, 2.901596e-08, 
    2.727285e-08, 2.759514e-08, 2.782691e-08, 2.640889e-08, 2.56971e-08, 
    2.781892e-08, 2.768403e-08, 2.641854e-08, 2.575736e-08, 2.496753e-08,
  3.129301e-08, 3.22387e-08, 3.121637e-08, 2.92406e-08, 2.844708e-08, 
    2.741076e-08, 2.762936e-08, 2.736573e-08, 2.635945e-08, 2.66429e-08, 
    2.754594e-08, 2.710901e-08, 2.597041e-08, 2.601723e-08, 2.535496e-08,
  3.204013e-08, 3.143286e-08, 3.016359e-08, 2.866708e-08, 2.814736e-08, 
    2.692677e-08, 2.788253e-08, 2.709248e-08, 2.651625e-08, 2.653416e-08, 
    2.731029e-08, 2.674815e-08, 2.593849e-08, 2.642118e-08, 2.612676e-08,
  3.182917e-08, 3.075473e-08, 2.95151e-08, 2.815367e-08, 2.792768e-08, 
    2.714595e-08, 2.759578e-08, 2.65806e-08, 2.661113e-08, 2.708148e-08, 
    2.695968e-08, 2.671577e-08, 2.612959e-08, 2.61244e-08, 2.61117e-08,
  2.877808e-08, 3.100693e-08, 3.147646e-08, 3.064067e-08, 3.041199e-08, 
    3.046371e-08, 2.996703e-08, 2.892246e-08, 2.938125e-08, 2.819906e-08, 
    2.617371e-08, 2.588001e-08, 2.613785e-08, 2.625213e-08, 2.467956e-08,
  3.066082e-08, 3.176269e-08, 3.128506e-08, 3.044596e-08, 3.075872e-08, 
    3.041696e-08, 2.916426e-08, 2.885279e-08, 2.920981e-08, 2.674729e-08, 
    2.570453e-08, 2.576942e-08, 2.604672e-08, 2.545267e-08, 2.415134e-08,
  3.197952e-08, 3.197536e-08, 3.106921e-08, 3.063061e-08, 3.03651e-08, 
    2.937741e-08, 2.801961e-08, 2.859682e-08, 2.845101e-08, 2.582743e-08, 
    2.550839e-08, 2.566453e-08, 2.579224e-08, 2.529044e-08, 2.495583e-08,
  3.197452e-08, 3.161891e-08, 3.099332e-08, 3.051019e-08, 2.955187e-08, 
    2.881385e-08, 2.786133e-08, 2.82833e-08, 2.745562e-08, 2.510633e-08, 
    2.547599e-08, 2.584252e-08, 2.615926e-08, 2.580505e-08, 2.569314e-08,
  3.196471e-08, 3.140446e-08, 3.10428e-08, 3.00101e-08, 2.884594e-08, 
    2.765119e-08, 2.774684e-08, 2.792682e-08, 2.698573e-08, 2.464673e-08, 
    2.553469e-08, 2.613123e-08, 2.65597e-08, 2.638326e-08, 2.611739e-08,
  3.22182e-08, 3.115448e-08, 3.072902e-08, 2.904653e-08, 2.794163e-08, 
    2.746031e-08, 2.717257e-08, 2.662529e-08, 2.66739e-08, 2.551406e-08, 
    2.601999e-08, 2.639925e-08, 2.697511e-08, 2.704155e-08, 2.651856e-08,
  3.191209e-08, 3.077938e-08, 2.995966e-08, 2.834348e-08, 2.763363e-08, 
    2.712097e-08, 2.693033e-08, 2.630413e-08, 2.667224e-08, 2.585805e-08, 
    2.605811e-08, 2.654507e-08, 2.719571e-08, 2.758189e-08, 2.711344e-08,
  3.154932e-08, 3.031361e-08, 2.927607e-08, 2.775104e-08, 2.709411e-08, 
    2.694821e-08, 2.651003e-08, 2.645462e-08, 2.686489e-08, 2.609793e-08, 
    2.592982e-08, 2.649728e-08, 2.735392e-08, 2.789618e-08, 2.816943e-08,
  3.092022e-08, 2.994361e-08, 2.863219e-08, 2.727216e-08, 2.713515e-08, 
    2.661424e-08, 2.627421e-08, 2.660551e-08, 2.669861e-08, 2.603081e-08, 
    2.577789e-08, 2.622568e-08, 2.699463e-08, 2.755253e-08, 2.857074e-08,
  3.057134e-08, 2.966284e-08, 2.797579e-08, 2.702274e-08, 2.707142e-08, 
    2.631065e-08, 2.639472e-08, 2.688626e-08, 2.641812e-08, 2.548451e-08, 
    2.511549e-08, 2.598903e-08, 2.664575e-08, 2.72148e-08, 2.834001e-08,
  2.829175e-08, 2.938576e-08, 3.123763e-08, 3.006516e-08, 2.851477e-08, 
    2.771303e-08, 2.869142e-08, 2.77214e-08, 2.669762e-08, 2.634671e-08, 
    2.559999e-08, 2.562494e-08, 2.620218e-08, 2.660689e-08, 2.594688e-08,
  2.869695e-08, 3.013868e-08, 3.124974e-08, 2.923679e-08, 2.824476e-08, 
    2.820661e-08, 2.905765e-08, 2.762269e-08, 2.655448e-08, 2.616535e-08, 
    2.594476e-08, 2.615884e-08, 2.706765e-08, 2.72182e-08, 2.651304e-08,
  2.922537e-08, 3.063561e-08, 3.065455e-08, 2.896084e-08, 2.791088e-08, 
    2.760114e-08, 2.901704e-08, 2.633844e-08, 2.615596e-08, 2.613944e-08, 
    2.621081e-08, 2.662949e-08, 2.735268e-08, 2.784233e-08, 2.730064e-08,
  2.966191e-08, 3.081357e-08, 3.017877e-08, 2.864222e-08, 2.726261e-08, 
    2.847494e-08, 2.566125e-08, 2.569934e-08, 2.645541e-08, 2.597529e-08, 
    2.627032e-08, 2.641329e-08, 2.701385e-08, 2.75658e-08, 2.692133e-08,
  3.049594e-08, 3.104206e-08, 2.973412e-08, 2.872063e-08, 2.707835e-08, 
    2.631041e-08, 2.589789e-08, 2.679809e-08, 2.609109e-08, 2.578373e-08, 
    2.592433e-08, 2.569413e-08, 2.650325e-08, 2.759033e-08, 2.725343e-08,
  3.094281e-08, 3.102407e-08, 2.948187e-08, 2.863051e-08, 2.617957e-08, 
    2.68681e-08, 2.691755e-08, 2.573029e-08, 2.709326e-08, 2.635475e-08, 
    2.464816e-08, 2.490475e-08, 2.635863e-08, 2.75838e-08, 2.780446e-08,
  3.129718e-08, 3.118222e-08, 2.930533e-08, 2.789921e-08, 2.558059e-08, 
    2.641578e-08, 2.725066e-08, 2.680306e-08, 2.669233e-08, 2.574276e-08, 
    2.497208e-08, 2.576871e-08, 2.677698e-08, 2.77096e-08, 2.875831e-08,
  3.124126e-08, 3.10938e-08, 2.922447e-08, 2.702345e-08, 2.516909e-08, 
    2.66449e-08, 2.709251e-08, 2.687724e-08, 2.723506e-08, 2.66054e-08, 
    2.611582e-08, 2.689422e-08, 2.786667e-08, 2.857434e-08, 2.906172e-08,
  3.121566e-08, 3.116011e-08, 2.909586e-08, 2.654408e-08, 2.494706e-08, 
    2.660992e-08, 2.735751e-08, 2.680769e-08, 2.702601e-08, 2.669166e-08, 
    2.696873e-08, 2.834086e-08, 2.923469e-08, 2.98264e-08, 2.997113e-08,
  3.099402e-08, 3.117643e-08, 2.942703e-08, 2.6132e-08, 2.466797e-08, 
    2.6591e-08, 2.711094e-08, 2.682158e-08, 2.722538e-08, 2.693023e-08, 
    2.750987e-08, 2.879175e-08, 2.996932e-08, 3.052103e-08, 3.026946e-08,
  2.854473e-08, 2.99799e-08, 3.345023e-08, 3.183747e-08, 2.847094e-08, 
    2.646508e-08, 2.739169e-08, 2.686733e-08, 2.531084e-08, 2.4965e-08, 
    2.532491e-08, 2.573894e-08, 2.665612e-08, 2.742584e-08, 2.571121e-08,
  2.893366e-08, 3.131489e-08, 3.315754e-08, 3.022106e-08, 2.727815e-08, 
    2.69132e-08, 2.786867e-08, 2.651326e-08, 2.493684e-08, 2.462375e-08, 
    2.547503e-08, 2.545837e-08, 2.621289e-08, 2.754927e-08, 2.594649e-08,
  3.055021e-08, 3.172162e-08, 3.21323e-08, 2.868816e-08, 2.594209e-08, 
    2.718675e-08, 2.810559e-08, 2.546488e-08, 2.51749e-08, 2.541721e-08, 
    2.562948e-08, 2.509133e-08, 2.561281e-08, 2.733588e-08, 2.619107e-08,
  3.09718e-08, 3.152042e-08, 3.115516e-08, 2.69197e-08, 2.50391e-08, 
    2.788111e-08, 2.675073e-08, 2.520664e-08, 2.598718e-08, 2.610828e-08, 
    2.610058e-08, 2.51293e-08, 2.528265e-08, 2.736446e-08, 2.645009e-08,
  3.113265e-08, 3.10771e-08, 2.990004e-08, 2.581953e-08, 2.558905e-08, 
    2.689779e-08, 2.674174e-08, 2.691445e-08, 2.653242e-08, 2.704538e-08, 
    2.703204e-08, 2.521553e-08, 2.49988e-08, 2.702761e-08, 2.665655e-08,
  3.055442e-08, 3.054397e-08, 2.898454e-08, 2.525941e-08, 2.625539e-08, 
    2.803384e-08, 2.755435e-08, 2.633604e-08, 2.770004e-08, 2.843106e-08, 
    2.80407e-08, 2.544874e-08, 2.481297e-08, 2.687728e-08, 2.692093e-08,
  2.988875e-08, 2.987247e-08, 2.809134e-08, 2.530521e-08, 2.732931e-08, 
    2.822152e-08, 2.761869e-08, 2.750949e-08, 2.752706e-08, 2.772267e-08, 
    2.93372e-08, 2.831584e-08, 2.612828e-08, 2.667418e-08, 2.720513e-08,
  2.914629e-08, 2.92892e-08, 2.779553e-08, 2.600575e-08, 2.812039e-08, 
    2.880993e-08, 2.785614e-08, 2.724528e-08, 2.714835e-08, 2.785204e-08, 
    2.956317e-08, 2.954363e-08, 2.755117e-08, 2.72496e-08, 2.740017e-08,
  2.864965e-08, 2.86447e-08, 2.781655e-08, 2.635583e-08, 2.86746e-08, 
    2.94633e-08, 2.792812e-08, 2.73737e-08, 2.698568e-08, 2.706686e-08, 
    2.855686e-08, 2.999345e-08, 2.888443e-08, 2.802873e-08, 2.710216e-08,
  2.830016e-08, 2.849247e-08, 2.82651e-08, 2.654679e-08, 2.773561e-08, 
    2.995415e-08, 2.879988e-08, 2.746959e-08, 2.712067e-08, 2.74945e-08, 
    2.807336e-08, 2.957022e-08, 2.942272e-08, 2.864625e-08, 2.717962e-08,
  3.005707e-08, 3.013023e-08, 2.939173e-08, 2.806273e-08, 2.910113e-08, 
    2.950934e-08, 2.896262e-08, 2.862959e-08, 2.808283e-08, 2.715423e-08, 
    2.685035e-08, 2.564094e-08, 2.59538e-08, 2.819995e-08, 2.994698e-08,
  3.06826e-08, 2.931938e-08, 2.880001e-08, 2.848981e-08, 2.999602e-08, 
    2.868509e-08, 2.910328e-08, 2.88718e-08, 2.682353e-08, 2.611497e-08, 
    2.674845e-08, 2.590677e-08, 2.605351e-08, 2.892947e-08, 3.010699e-08,
  3.022518e-08, 2.864743e-08, 2.90856e-08, 2.925171e-08, 2.899654e-08, 
    2.91705e-08, 2.862489e-08, 2.460531e-08, 2.495281e-08, 2.612161e-08, 
    2.712037e-08, 2.618493e-08, 2.669454e-08, 2.894766e-08, 3.014754e-08,
  2.942086e-08, 2.881989e-08, 2.953506e-08, 2.874904e-08, 2.796282e-08, 
    2.898516e-08, 2.594459e-08, 2.357817e-08, 2.526479e-08, 2.628827e-08, 
    2.740627e-08, 2.624009e-08, 2.677951e-08, 2.911858e-08, 2.982891e-08,
  2.919027e-08, 2.91006e-08, 2.965684e-08, 2.856061e-08, 2.833746e-08, 
    2.830756e-08, 2.513827e-08, 2.668756e-08, 2.669117e-08, 2.643195e-08, 
    2.744418e-08, 2.640549e-08, 2.690763e-08, 2.917626e-08, 3.010755e-08,
  2.893808e-08, 2.942182e-08, 2.961592e-08, 2.778052e-08, 2.82421e-08, 
    2.836923e-08, 2.708144e-08, 2.666064e-08, 2.64966e-08, 2.724243e-08, 
    2.796364e-08, 2.634407e-08, 2.703403e-08, 2.897202e-08, 2.993041e-08,
  2.884181e-08, 2.964983e-08, 2.913362e-08, 2.72466e-08, 2.818521e-08, 
    2.849566e-08, 2.762605e-08, 2.682276e-08, 2.669324e-08, 2.796625e-08, 
    2.814436e-08, 2.629902e-08, 2.712722e-08, 2.880121e-08, 2.963216e-08,
  2.85461e-08, 2.972803e-08, 2.903336e-08, 2.709097e-08, 2.800129e-08, 
    2.85045e-08, 2.872344e-08, 2.796095e-08, 2.777714e-08, 2.869646e-08, 
    2.778785e-08, 2.593582e-08, 2.70677e-08, 2.855639e-08, 2.933863e-08,
  2.79329e-08, 2.96206e-08, 2.900158e-08, 2.704026e-08, 2.789213e-08, 
    2.844457e-08, 2.912982e-08, 2.890741e-08, 2.851033e-08, 2.873302e-08, 
    2.682711e-08, 2.612363e-08, 2.704624e-08, 2.828367e-08, 2.904109e-08,
  2.756495e-08, 2.955403e-08, 2.940727e-08, 2.707859e-08, 2.789862e-08, 
    2.820683e-08, 2.924325e-08, 2.968054e-08, 2.900965e-08, 2.79429e-08, 
    2.67985e-08, 2.626607e-08, 2.682938e-08, 2.783322e-08, 2.866081e-08,
  3.249047e-08, 3.433899e-08, 3.341519e-08, 3.170981e-08, 3.137514e-08, 
    2.803773e-08, 2.73762e-08, 2.693413e-08, 2.6769e-08, 2.693193e-08, 
    2.616514e-08, 2.749931e-08, 2.688228e-08, 3.012119e-08, 2.79062e-08,
  3.39222e-08, 3.470632e-08, 3.305474e-08, 3.173028e-08, 3.015093e-08, 
    2.793456e-08, 2.806842e-08, 2.784333e-08, 2.714043e-08, 2.645088e-08, 
    2.623849e-08, 2.700003e-08, 2.691986e-08, 3.086789e-08, 2.72587e-08,
  3.451101e-08, 3.418702e-08, 3.261663e-08, 3.072268e-08, 2.844428e-08, 
    2.917042e-08, 2.827401e-08, 2.737906e-08, 2.620743e-08, 2.603096e-08, 
    2.632816e-08, 2.741175e-08, 2.791661e-08, 3.055371e-08, 2.608127e-08,
  3.496915e-08, 3.34602e-08, 3.197494e-08, 2.895894e-08, 2.794119e-08, 
    2.936129e-08, 2.947153e-08, 2.7863e-08, 2.557805e-08, 2.531089e-08, 
    2.66234e-08, 2.801335e-08, 2.894718e-08, 2.950183e-08, 2.497952e-08,
  3.470772e-08, 3.208914e-08, 3.079681e-08, 2.809966e-08, 2.846927e-08, 
    2.927939e-08, 2.936928e-08, 2.675159e-08, 2.597469e-08, 2.509773e-08, 
    2.747142e-08, 2.860788e-08, 2.966561e-08, 2.860052e-08, 2.451099e-08,
  3.302487e-08, 3.04754e-08, 2.973741e-08, 2.74135e-08, 2.871452e-08, 
    3.01897e-08, 2.828641e-08, 2.509433e-08, 2.313632e-08, 2.595849e-08, 
    2.87591e-08, 2.920379e-08, 2.970616e-08, 2.749268e-08, 2.427112e-08,
  3.113235e-08, 2.94975e-08, 2.89597e-08, 2.721482e-08, 2.920221e-08, 
    2.959067e-08, 2.794431e-08, 2.499022e-08, 2.454921e-08, 2.838515e-08, 
    2.917267e-08, 2.930631e-08, 2.956733e-08, 2.682967e-08, 2.488577e-08,
  2.937515e-08, 2.899784e-08, 2.840093e-08, 2.702778e-08, 2.889148e-08, 
    2.884286e-08, 2.721286e-08, 2.50139e-08, 2.645197e-08, 2.888613e-08, 
    2.887652e-08, 2.912668e-08, 2.891434e-08, 2.682456e-08, 2.625173e-08,
  2.828235e-08, 2.880078e-08, 2.771572e-08, 2.683412e-08, 2.892446e-08, 
    2.851632e-08, 2.715982e-08, 2.64848e-08, 2.768314e-08, 2.902656e-08, 
    2.836406e-08, 2.882303e-08, 2.891509e-08, 2.734955e-08, 2.782067e-08,
  2.756775e-08, 2.833735e-08, 2.717175e-08, 2.646066e-08, 2.770869e-08, 
    2.784676e-08, 2.724691e-08, 2.703571e-08, 2.811831e-08, 2.906917e-08, 
    2.789689e-08, 2.888027e-08, 2.874116e-08, 2.769986e-08, 2.909004e-08,
  2.964989e-08, 2.978612e-08, 3.126504e-08, 3.21138e-08, 3.325924e-08, 
    3.340299e-08, 3.163888e-08, 3.057735e-08, 2.960829e-08, 2.779287e-08, 
    2.76143e-08, 2.79772e-08, 2.902966e-08, 3.059078e-08, 3.150303e-08,
  2.940744e-08, 3.063948e-08, 3.194187e-08, 3.282967e-08, 3.334484e-08, 
    3.352386e-08, 3.035769e-08, 3.093416e-08, 2.859346e-08, 2.767793e-08, 
    2.721512e-08, 2.83973e-08, 2.975984e-08, 3.117471e-08, 3.219202e-08,
  2.921337e-08, 3.083436e-08, 3.209819e-08, 3.331566e-08, 3.247051e-08, 
    3.244848e-08, 2.927079e-08, 2.876975e-08, 2.799203e-08, 2.80226e-08, 
    2.746857e-08, 2.921404e-08, 3.096347e-08, 3.163487e-08, 3.219571e-08,
  3.053981e-08, 3.18263e-08, 3.290176e-08, 3.27122e-08, 3.060097e-08, 
    3.062089e-08, 3.061903e-08, 2.880183e-08, 2.842603e-08, 2.741715e-08, 
    2.786561e-08, 2.990005e-08, 3.123447e-08, 3.170623e-08, 3.176564e-08,
  3.177086e-08, 3.21627e-08, 3.235371e-08, 3.053491e-08, 3.000671e-08, 
    2.767691e-08, 2.9403e-08, 2.950733e-08, 2.882055e-08, 2.771821e-08, 
    2.867892e-08, 3.062213e-08, 3.132846e-08, 3.207434e-08, 3.1773e-08,
  3.216599e-08, 3.16602e-08, 3.066575e-08, 2.915489e-08, 2.75976e-08, 
    2.892511e-08, 2.782723e-08, 2.818518e-08, 2.769046e-08, 2.768829e-08, 
    2.951218e-08, 3.080158e-08, 3.133839e-08, 3.145744e-08, 3.068844e-08,
  3.20829e-08, 3.026813e-08, 2.905406e-08, 2.721781e-08, 2.797572e-08, 
    2.858272e-08, 2.747279e-08, 2.730293e-08, 2.648729e-08, 2.811779e-08, 
    3.0174e-08, 3.096643e-08, 3.09514e-08, 3.038731e-08, 2.973658e-08,
  3.007562e-08, 2.813594e-08, 2.716316e-08, 2.709876e-08, 2.823636e-08, 
    2.784441e-08, 2.632726e-08, 2.627917e-08, 2.7337e-08, 2.945535e-08, 
    3.064033e-08, 3.019688e-08, 2.9541e-08, 2.949974e-08, 2.873507e-08,
  2.76978e-08, 2.729364e-08, 2.669109e-08, 2.708306e-08, 2.752747e-08, 
    2.589365e-08, 2.544865e-08, 2.587854e-08, 2.835843e-08, 3.026282e-08, 
    2.992357e-08, 2.902712e-08, 2.831843e-08, 2.809825e-08, 2.838709e-08,
  2.686022e-08, 2.651558e-08, 2.635332e-08, 2.70297e-08, 2.628291e-08, 
    2.547711e-08, 2.565492e-08, 2.692846e-08, 2.981193e-08, 2.982758e-08, 
    2.885221e-08, 2.776992e-08, 2.703042e-08, 2.727054e-08, 2.906201e-08,
  2.81134e-08, 2.779776e-08, 2.711859e-08, 2.829406e-08, 2.825829e-08, 
    2.885729e-08, 2.937979e-08, 2.946866e-08, 3.082685e-08, 3.134955e-08, 
    2.999303e-08, 2.844572e-08, 2.685741e-08, 2.846041e-08, 3.11898e-08,
  2.825405e-08, 2.804692e-08, 2.812234e-08, 2.89082e-08, 2.910596e-08, 
    2.990587e-08, 2.997978e-08, 3.089434e-08, 3.11803e-08, 2.978155e-08, 
    2.892274e-08, 2.71399e-08, 2.658887e-08, 3.118099e-08, 3.207421e-08,
  2.864592e-08, 2.863088e-08, 2.866529e-08, 2.959599e-08, 2.965544e-08, 
    3.076973e-08, 3.054267e-08, 3.042814e-08, 3.036196e-08, 2.935736e-08, 
    2.77031e-08, 2.681496e-08, 2.877595e-08, 3.286801e-08, 3.019418e-08,
  2.954229e-08, 2.996349e-08, 2.956476e-08, 3.056184e-08, 2.997639e-08, 
    3.036991e-08, 3.271939e-08, 3.039583e-08, 2.817092e-08, 2.793186e-08, 
    2.77139e-08, 2.813935e-08, 3.159093e-08, 3.067825e-08, 2.858447e-08,
  2.985577e-08, 2.96018e-08, 3.064652e-08, 2.997111e-08, 3.163697e-08, 
    2.990875e-08, 3.064607e-08, 3.246979e-08, 3.061341e-08, 2.737292e-08, 
    2.790368e-08, 3.043847e-08, 3.233991e-08, 2.968207e-08, 2.904144e-08,
  2.962174e-08, 3.067478e-08, 3.078986e-08, 3.231745e-08, 3.095925e-08, 
    3.082737e-08, 2.822215e-08, 2.854566e-08, 2.892391e-08, 2.8073e-08, 
    2.928155e-08, 3.208446e-08, 3.085291e-08, 2.865826e-08, 2.844482e-08,
  3.063978e-08, 3.157445e-08, 3.212424e-08, 3.178e-08, 3.066727e-08, 
    2.995889e-08, 2.886587e-08, 2.785414e-08, 2.777148e-08, 2.869436e-08, 
    3.172167e-08, 3.205182e-08, 2.997451e-08, 2.87922e-08, 2.827727e-08,
  3.239249e-08, 3.22179e-08, 3.1688e-08, 3.084357e-08, 2.977565e-08, 
    2.909074e-08, 2.840211e-08, 2.809201e-08, 2.842002e-08, 3.075666e-08, 
    3.287836e-08, 3.15806e-08, 2.980978e-08, 2.810333e-08, 2.632211e-08,
  3.146525e-08, 3.007673e-08, 2.942646e-08, 2.856833e-08, 2.801717e-08, 
    2.783566e-08, 2.787902e-08, 2.825325e-08, 2.979497e-08, 3.294419e-08, 
    3.341608e-08, 3.013894e-08, 2.887517e-08, 2.753067e-08, 2.788589e-08,
  2.873111e-08, 2.773967e-08, 2.751157e-08, 2.738306e-08, 2.740607e-08, 
    2.798757e-08, 2.881267e-08, 2.984368e-08, 3.296843e-08, 3.395398e-08, 
    3.067818e-08, 2.986965e-08, 3.027203e-08, 3.21836e-08, 3.68708e-08,
  2.946441e-08, 2.994474e-08, 2.961754e-08, 2.894213e-08, 2.747514e-08, 
    2.72512e-08, 2.747437e-08, 2.719431e-08, 2.798969e-08, 2.905088e-08, 
    3.120179e-08, 3.126972e-08, 3.070495e-08, 2.693342e-08, 2.555326e-08,
  2.961833e-08, 3.02362e-08, 2.950984e-08, 2.919921e-08, 2.661781e-08, 
    2.709265e-08, 2.730381e-08, 2.817844e-08, 2.885544e-08, 2.915711e-08, 
    3.161166e-08, 3.1935e-08, 2.855788e-08, 2.964955e-08, 2.758443e-08,
  2.924154e-08, 2.996277e-08, 2.925635e-08, 2.872868e-08, 2.617682e-08, 
    2.646483e-08, 2.716095e-08, 2.789965e-08, 2.818484e-08, 2.976145e-08, 
    3.324555e-08, 3.031678e-08, 2.924949e-08, 3.103392e-08, 2.943634e-08,
  2.864111e-08, 2.974902e-08, 2.90764e-08, 2.883201e-08, 2.636662e-08, 
    2.625027e-08, 2.929827e-08, 2.891307e-08, 2.84032e-08, 3.153173e-08, 
    3.282933e-08, 2.939941e-08, 3.094433e-08, 3.049263e-08, 2.983822e-08,
  2.811964e-08, 2.9664e-08, 2.878077e-08, 2.855298e-08, 2.703017e-08, 
    2.841857e-08, 2.862578e-08, 3.157024e-08, 3.43257e-08, 3.304334e-08, 
    3.043878e-08, 3.009442e-08, 3.046858e-08, 2.995099e-08, 3.009951e-08,
  2.780066e-08, 3.003825e-08, 2.926395e-08, 2.88762e-08, 2.772859e-08, 
    2.855825e-08, 2.826542e-08, 2.778851e-08, 3.072394e-08, 3.020367e-08, 
    2.846988e-08, 3.080062e-08, 2.906794e-08, 2.897292e-08, 2.984858e-08,
  2.794989e-08, 2.988094e-08, 2.95159e-08, 2.922592e-08, 2.819283e-08, 
    2.823681e-08, 2.899108e-08, 3.022515e-08, 3.142346e-08, 2.953767e-08, 
    3.053303e-08, 2.920665e-08, 2.712765e-08, 2.759833e-08, 2.908711e-08,
  2.787647e-08, 2.952502e-08, 2.963565e-08, 2.946411e-08, 2.886807e-08, 
    2.842305e-08, 2.938918e-08, 3.141232e-08, 3.026097e-08, 2.874974e-08, 
    2.95247e-08, 2.717833e-08, 2.640366e-08, 2.697711e-08, 2.736523e-08,
  2.850533e-08, 2.973018e-08, 3.009788e-08, 3.02887e-08, 2.965524e-08, 
    2.917345e-08, 2.979482e-08, 3.06338e-08, 2.873108e-08, 2.907542e-08, 
    2.874878e-08, 2.495068e-08, 2.369974e-08, 2.369728e-08, 2.406525e-08,
  2.966071e-08, 3.06237e-08, 3.042021e-08, 3.001233e-08, 2.929273e-08, 
    2.90305e-08, 2.931626e-08, 2.941315e-08, 2.861654e-08, 2.886962e-08, 
    2.44708e-08, 2.306636e-08, 2.363583e-08, 2.41907e-08, 2.58865e-08,
  3.012244e-08, 3.023927e-08, 3.012845e-08, 2.930912e-08, 2.849415e-08, 
    2.823656e-08, 2.825043e-08, 2.843981e-08, 2.867726e-08, 2.755148e-08, 
    2.7698e-08, 2.77217e-08, 3.162079e-08, 2.994754e-08, 2.832263e-08,
  3.014759e-08, 3.014138e-08, 3.007412e-08, 2.96248e-08, 2.755921e-08, 
    2.830072e-08, 2.779594e-08, 2.816706e-08, 2.855706e-08, 2.791895e-08, 
    2.817249e-08, 2.935114e-08, 3.110934e-08, 3.083147e-08, 2.838613e-08,
  2.98794e-08, 2.994021e-08, 2.970515e-08, 2.812122e-08, 2.671136e-08, 
    2.780011e-08, 2.787008e-08, 2.751318e-08, 2.763917e-08, 2.819761e-08, 
    2.92487e-08, 3.090455e-08, 3.039738e-08, 3.130451e-08, 3.001854e-08,
  2.990847e-08, 2.979975e-08, 2.924272e-08, 2.813381e-08, 2.865762e-08, 
    2.707098e-08, 2.75173e-08, 2.741167e-08, 2.748943e-08, 2.843038e-08, 
    3.021738e-08, 3.079312e-08, 3.142392e-08, 3.182923e-08, 3.163379e-08,
  2.998579e-08, 2.993759e-08, 2.892145e-08, 2.848076e-08, 2.863279e-08, 
    2.732433e-08, 2.642233e-08, 2.839e-08, 3.001897e-08, 3.051217e-08, 
    3.133436e-08, 3.168637e-08, 3.149653e-08, 3.161937e-08, 3.067537e-08,
  2.985922e-08, 2.955511e-08, 2.889203e-08, 2.912505e-08, 2.795002e-08, 
    2.722677e-08, 2.871096e-08, 2.898352e-08, 3.030522e-08, 3.181913e-08, 
    3.126955e-08, 3.133019e-08, 3.04707e-08, 2.916472e-08, 2.918611e-08,
  2.949854e-08, 2.95369e-08, 2.898215e-08, 2.93137e-08, 2.696525e-08, 
    2.590556e-08, 2.927379e-08, 3.069134e-08, 3.154914e-08, 3.195937e-08, 
    3.108542e-08, 3.05608e-08, 2.904163e-08, 2.736416e-08, 2.816688e-08,
  2.941183e-08, 2.959379e-08, 2.914033e-08, 2.938104e-08, 2.627949e-08, 
    2.523015e-08, 2.989337e-08, 3.006184e-08, 3.064034e-08, 2.959033e-08, 
    3.053418e-08, 2.923511e-08, 2.632682e-08, 2.594492e-08, 2.783146e-08,
  2.928885e-08, 2.95456e-08, 2.87368e-08, 2.887678e-08, 2.547334e-08, 
    2.580068e-08, 2.884163e-08, 2.97541e-08, 3.042932e-08, 3.064921e-08, 
    3.226462e-08, 2.792034e-08, 2.403194e-08, 2.667551e-08, 2.870958e-08,
  2.870422e-08, 2.898634e-08, 2.919067e-08, 2.969167e-08, 2.620431e-08, 
    2.822205e-08, 2.833394e-08, 3.057281e-08, 3.112749e-08, 3.36953e-08, 
    3.326171e-08, 2.617454e-08, 2.259639e-08, 2.675644e-08, 2.927728e-08,
  2.969811e-08, 2.975976e-08, 3.027121e-08, 2.991554e-08, 2.989431e-08, 
    3.05674e-08, 3.082664e-08, 3.080108e-08, 2.992301e-08, 2.944322e-08, 
    2.791191e-08, 2.67449e-08, 2.669605e-08, 2.753879e-08, 2.809375e-08,
  3.008703e-08, 2.98067e-08, 3.046483e-08, 3.008775e-08, 2.916722e-08, 
    3.004109e-08, 3.060303e-08, 3.065137e-08, 3.018711e-08, 2.951962e-08, 
    2.861645e-08, 2.744036e-08, 2.784097e-08, 2.85722e-08, 2.848167e-08,
  3.035229e-08, 3.029418e-08, 3.062713e-08, 3.032447e-08, 2.899388e-08, 
    2.892754e-08, 2.992399e-08, 3.078266e-08, 2.977873e-08, 2.919623e-08, 
    2.868754e-08, 2.831938e-08, 2.851858e-08, 2.858214e-08, 2.856012e-08,
  3.109895e-08, 3.05282e-08, 2.998038e-08, 2.872566e-08, 2.721834e-08, 
    2.799148e-08, 2.91813e-08, 2.945223e-08, 3.00411e-08, 2.949204e-08, 
    2.898081e-08, 2.88464e-08, 2.901898e-08, 2.897208e-08, 2.915771e-08,
  3.097625e-08, 2.996179e-08, 2.769667e-08, 2.73397e-08, 2.775998e-08, 
    2.875511e-08, 2.847213e-08, 2.988512e-08, 2.941691e-08, 2.900324e-08, 
    2.928573e-08, 2.933645e-08, 2.924004e-08, 2.932524e-08, 2.948298e-08,
  2.807781e-08, 2.692869e-08, 2.611351e-08, 2.659057e-08, 2.809176e-08, 
    2.998044e-08, 3.021591e-08, 2.710689e-08, 2.632366e-08, 2.875147e-08, 
    2.930763e-08, 2.962335e-08, 2.990801e-08, 2.978418e-08, 2.975481e-08,
  2.718613e-08, 2.625045e-08, 2.683669e-08, 2.818576e-08, 2.963479e-08, 
    2.944835e-08, 2.80226e-08, 2.644476e-08, 2.716169e-08, 2.897875e-08, 
    2.972061e-08, 3.025447e-08, 3.035911e-08, 3.052115e-08, 3.075663e-08,
  2.783925e-08, 2.813531e-08, 2.98947e-08, 3.071892e-08, 3.029384e-08, 
    2.849981e-08, 2.7821e-08, 2.752475e-08, 2.85697e-08, 2.939416e-08, 
    2.957859e-08, 3.02111e-08, 3.083614e-08, 3.075692e-08, 3.014276e-08,
  2.86318e-08, 2.908696e-08, 2.945505e-08, 2.857363e-08, 2.623364e-08, 
    2.467275e-08, 2.801039e-08, 2.802993e-08, 2.935018e-08, 3.039368e-08, 
    3.160481e-08, 3.295654e-08, 3.246326e-08, 3.095355e-08, 3.015695e-08,
  2.892518e-08, 2.913474e-08, 2.899877e-08, 2.672639e-08, 2.439638e-08, 
    2.661052e-08, 2.886741e-08, 3.033007e-08, 3.312108e-08, 3.303296e-08, 
    3.512296e-08, 3.392629e-08, 2.994725e-08, 2.815379e-08, 2.73933e-08,
  2.942881e-08, 3.002296e-08, 3.036858e-08, 3.057067e-08, 3.027095e-08, 
    3.235202e-08, 3.37351e-08, 3.403532e-08, 2.912308e-08, 2.454769e-08, 
    2.320501e-08, 2.275821e-08, 2.341642e-08, 2.446843e-08, 2.47693e-08,
  2.956913e-08, 3.022257e-08, 3.090373e-08, 3.08488e-08, 3.036219e-08, 
    3.289508e-08, 3.367272e-08, 3.462155e-08, 2.985727e-08, 2.589737e-08, 
    2.350694e-08, 2.278579e-08, 2.295919e-08, 2.331093e-08, 2.383944e-08,
  3.036611e-08, 3.078172e-08, 3.128584e-08, 3.028852e-08, 2.968219e-08, 
    3.268213e-08, 3.574334e-08, 3.651078e-08, 2.997485e-08, 2.65901e-08, 
    2.420312e-08, 2.283989e-08, 2.246004e-08, 2.278064e-08, 2.353092e-08,
  3.08628e-08, 3.06642e-08, 3.054915e-08, 3.112907e-08, 3.066014e-08, 
    3.167673e-08, 3.532832e-08, 3.746206e-08, 3.246899e-08, 2.721183e-08, 
    2.521433e-08, 2.361513e-08, 2.292485e-08, 2.386009e-08, 2.479611e-08,
  2.987095e-08, 2.956191e-08, 2.923126e-08, 3.096024e-08, 3.054859e-08, 
    2.990042e-08, 3.227543e-08, 3.410901e-08, 3.545907e-08, 2.93633e-08, 
    2.600648e-08, 2.493461e-08, 2.431588e-08, 2.505016e-08, 2.580204e-08,
  3.02441e-08, 3.021857e-08, 2.97958e-08, 3.094064e-08, 3.079011e-08, 
    2.96387e-08, 3.156067e-08, 3.306764e-08, 3.206039e-08, 2.777351e-08, 
    2.672026e-08, 2.652535e-08, 2.536732e-08, 2.537338e-08, 2.622514e-08,
  2.874036e-08, 2.905655e-08, 2.947909e-08, 3.059946e-08, 3.011624e-08, 
    2.853569e-08, 3.088392e-08, 3.186026e-08, 3.056618e-08, 2.919634e-08, 
    2.820182e-08, 2.784579e-08, 2.698291e-08, 2.719654e-08, 2.791102e-08,
  2.799763e-08, 2.813908e-08, 2.882841e-08, 2.93352e-08, 2.957067e-08, 
    2.83969e-08, 2.953762e-08, 3.032225e-08, 2.930468e-08, 2.882667e-08, 
    2.819871e-08, 2.810274e-08, 2.815239e-08, 2.858004e-08, 2.925987e-08,
  2.879078e-08, 2.910202e-08, 2.910853e-08, 2.918507e-08, 2.947255e-08, 
    2.873969e-08, 2.855933e-08, 2.940209e-08, 2.873263e-08, 2.865174e-08, 
    2.875625e-08, 2.832405e-08, 2.856576e-08, 2.889207e-08, 2.971642e-08,
  2.906994e-08, 2.860323e-08, 2.766734e-08, 2.684867e-08, 2.754803e-08, 
    2.844159e-08, 2.861129e-08, 2.904077e-08, 2.91711e-08, 2.935138e-08, 
    2.986858e-08, 2.979124e-08, 3.061395e-08, 3.161498e-08, 3.227361e-08,
  2.760511e-08, 2.833469e-08, 2.82143e-08, 2.916064e-08, 2.952548e-08, 
    2.991793e-08, 2.96943e-08, 2.993765e-08, 3.031018e-08, 3.069374e-08, 
    3.059151e-08, 2.909189e-08, 3.030203e-08, 2.964707e-08, 2.96863e-08,
  2.963351e-08, 2.991742e-08, 3.033229e-08, 2.965669e-08, 2.994104e-08, 
    3.062603e-08, 3.029686e-08, 3.042726e-08, 3.075733e-08, 3.121256e-08, 
    3.067757e-08, 2.90566e-08, 2.952933e-08, 2.897075e-08, 2.91361e-08,
  3.006703e-08, 3.019048e-08, 3.078206e-08, 3.032773e-08, 3.01373e-08, 
    3.077162e-08, 3.09185e-08, 3.100137e-08, 3.094255e-08, 3.183191e-08, 
    3.098211e-08, 2.94397e-08, 2.975611e-08, 2.89583e-08, 2.829667e-08,
  3.008144e-08, 3.049054e-08, 3.021174e-08, 3.028894e-08, 2.974107e-08, 
    2.997553e-08, 3.151787e-08, 3.057155e-08, 3.114969e-08, 3.206304e-08, 
    3.13882e-08, 3.005146e-08, 2.991215e-08, 2.868315e-08, 2.672951e-08,
  2.974781e-08, 3.036614e-08, 3.091828e-08, 3.115611e-08, 2.974649e-08, 
    3.019633e-08, 2.94983e-08, 3.023799e-08, 3.653646e-08, 3.259448e-08, 
    3.129956e-08, 3.011997e-08, 2.950557e-08, 2.75916e-08, 2.556898e-08,
  3.157561e-08, 3.214594e-08, 3.285325e-08, 3.298645e-08, 3.059482e-08, 
    3.089251e-08, 3.000735e-08, 3.31174e-08, 3.596179e-08, 3.146613e-08, 
    3.072427e-08, 2.955307e-08, 2.834495e-08, 2.633898e-08, 2.446443e-08,
  3.219592e-08, 3.354903e-08, 3.306069e-08, 3.22265e-08, 3.157279e-08, 
    3.107003e-08, 3.125636e-08, 3.347635e-08, 3.432387e-08, 3.010373e-08, 
    2.923846e-08, 2.844358e-08, 2.684052e-08, 2.493884e-08, 2.385089e-08,
  3.151647e-08, 3.331516e-08, 3.257732e-08, 3.237732e-08, 3.248971e-08, 
    3.12906e-08, 3.117505e-08, 3.374366e-08, 3.407433e-08, 2.980316e-08, 
    2.829995e-08, 2.77677e-08, 2.608523e-08, 2.470047e-08, 2.364634e-08,
  3.085334e-08, 3.158446e-08, 3.202148e-08, 3.202865e-08, 3.177177e-08, 
    3.123212e-08, 3.214656e-08, 3.357827e-08, 3.288253e-08, 2.833241e-08, 
    2.725243e-08, 2.615515e-08, 2.50866e-08, 2.456391e-08, 2.438851e-08,
  3.02812e-08, 3.061275e-08, 3.09417e-08, 3.078877e-08, 3.155577e-08, 
    3.046156e-08, 3.177208e-08, 3.331151e-08, 3.230225e-08, 2.71796e-08, 
    2.632168e-08, 2.563903e-08, 2.534082e-08, 2.525459e-08, 2.538922e-08,
  2.874764e-08, 2.849205e-08, 2.795673e-08, 2.769733e-08, 2.719344e-08, 
    2.703269e-08, 2.670561e-08, 2.719525e-08, 2.834209e-08, 2.967592e-08, 
    3.140506e-08, 3.246309e-08, 3.219816e-08, 3.10121e-08, 3.051611e-08,
  2.907038e-08, 2.87814e-08, 2.91942e-08, 2.900871e-08, 2.89045e-08, 
    2.808044e-08, 2.753226e-08, 2.736795e-08, 2.805448e-08, 2.894516e-08, 
    3.063974e-08, 3.158975e-08, 3.181884e-08, 3.124778e-08, 3.074714e-08,
  2.92519e-08, 2.902754e-08, 2.95557e-08, 2.932211e-08, 3.001847e-08, 
    2.904407e-08, 2.80739e-08, 2.777043e-08, 2.805696e-08, 2.94142e-08, 
    3.079053e-08, 3.145698e-08, 3.178089e-08, 3.172178e-08, 3.139754e-08,
  2.914175e-08, 2.947869e-08, 2.997323e-08, 2.983333e-08, 2.928059e-08, 
    2.92291e-08, 2.867242e-08, 2.803237e-08, 2.84728e-08, 2.953665e-08, 
    3.102046e-08, 3.152688e-08, 3.176602e-08, 3.173399e-08, 3.116672e-08,
  2.955266e-08, 3.087685e-08, 3.14133e-08, 3.113174e-08, 3.041215e-08, 
    2.951434e-08, 2.846185e-08, 2.809313e-08, 2.990493e-08, 3.053794e-08, 
    3.11951e-08, 3.146621e-08, 3.1646e-08, 3.226584e-08, 3.176276e-08,
  2.999425e-08, 3.206434e-08, 3.241137e-08, 3.279419e-08, 3.041885e-08, 
    2.915977e-08, 2.85456e-08, 2.769446e-08, 2.906608e-08, 3.110856e-08, 
    3.135765e-08, 3.147297e-08, 3.189341e-08, 3.223448e-08, 3.145507e-08,
  2.973511e-08, 3.143295e-08, 3.094902e-08, 3.349764e-08, 3.183314e-08, 
    3.040742e-08, 2.862007e-08, 2.845542e-08, 2.99799e-08, 3.09275e-08, 
    3.123379e-08, 3.145141e-08, 3.205129e-08, 3.228629e-08, 3.061062e-08,
  2.962025e-08, 3.141387e-08, 3.181777e-08, 3.209684e-08, 3.196799e-08, 
    3.04075e-08, 2.875524e-08, 2.91668e-08, 3.070874e-08, 3.117949e-08, 
    3.120767e-08, 3.15632e-08, 3.203109e-08, 3.175331e-08, 2.918868e-08,
  2.835349e-08, 3.005484e-08, 3.094292e-08, 3.083617e-08, 3.115516e-08, 
    3.002397e-08, 2.901258e-08, 2.993393e-08, 3.09263e-08, 3.074418e-08, 
    3.134549e-08, 3.200848e-08, 3.241272e-08, 3.072624e-08, 2.645657e-08,
  2.888071e-08, 3.000722e-08, 3.005904e-08, 2.969164e-08, 3.110069e-08, 
    2.934832e-08, 2.984074e-08, 3.060633e-08, 3.143894e-08, 3.082069e-08, 
    3.1823e-08, 3.228987e-08, 3.193684e-08, 2.951106e-08, 2.51548e-08,
  3.15409e-08, 3.138732e-08, 3.071176e-08, 3.0257e-08, 2.968808e-08, 
    2.960248e-08, 2.91621e-08, 2.867799e-08, 2.882672e-08, 2.980941e-08, 
    3.042686e-08, 3.133922e-08, 3.248254e-08, 3.240716e-08, 3.344307e-08,
  3.057675e-08, 3.032943e-08, 3.031534e-08, 3.001065e-08, 2.991359e-08, 
    3.033015e-08, 3.122747e-08, 3.111422e-08, 3.008354e-08, 2.964653e-08, 
    2.973782e-08, 3.132477e-08, 3.263487e-08, 3.23069e-08, 3.241156e-08,
  2.982829e-08, 3.039476e-08, 3.011307e-08, 2.97016e-08, 2.915682e-08, 
    3.008422e-08, 3.313538e-08, 3.410186e-08, 3.182121e-08, 2.941823e-08, 
    2.86597e-08, 3.08536e-08, 3.309563e-08, 3.224381e-08, 3.186186e-08,
  2.981727e-08, 2.964576e-08, 2.864508e-08, 2.852473e-08, 2.736681e-08, 
    2.545973e-08, 2.838335e-08, 3.093272e-08, 3.090498e-08, 2.849986e-08, 
    2.806882e-08, 3.083152e-08, 3.344726e-08, 3.237323e-08, 3.139374e-08,
  2.835209e-08, 2.74552e-08, 2.712886e-08, 2.71137e-08, 2.844644e-08, 
    2.557056e-08, 2.190887e-08, 2.57191e-08, 2.767179e-08, 2.693045e-08, 
    2.850632e-08, 3.169866e-08, 3.389261e-08, 3.263428e-08, 3.194431e-08,
  2.541573e-08, 2.686504e-08, 2.869156e-08, 2.990291e-08, 3.10205e-08, 
    3.000643e-08, 2.56828e-08, 2.559905e-08, 2.693412e-08, 2.764203e-08, 
    2.984959e-08, 3.301561e-08, 3.349497e-08, 3.252866e-08, 3.143962e-08,
  2.724767e-08, 2.886523e-08, 3.093891e-08, 3.122747e-08, 3.131366e-08, 
    3.050087e-08, 2.821037e-08, 2.702896e-08, 2.763077e-08, 2.904222e-08, 
    3.215055e-08, 3.357915e-08, 3.299438e-08, 3.212271e-08, 3.254147e-08,
  2.810338e-08, 3.004488e-08, 3.164072e-08, 3.292653e-08, 3.218415e-08, 
    3.090966e-08, 2.830319e-08, 2.818718e-08, 2.893189e-08, 3.123751e-08, 
    3.343943e-08, 3.323844e-08, 3.260889e-08, 3.312784e-08, 3.096591e-08,
  2.760534e-08, 3.05865e-08, 3.094189e-08, 3.292051e-08, 3.107641e-08, 
    2.987235e-08, 2.829586e-08, 2.89439e-08, 3.066576e-08, 3.30968e-08, 
    3.353111e-08, 3.314365e-08, 3.2386e-08, 3.039898e-08, 2.344307e-08,
  2.753345e-08, 3.038594e-08, 3.006977e-08, 3.021621e-08, 2.924835e-08, 
    2.917009e-08, 2.850915e-08, 3.038053e-08, 3.290249e-08, 3.359346e-08, 
    3.336047e-08, 3.25308e-08, 3.102759e-08, 2.712857e-08, 2.60295e-08,
  3.240653e-08, 3.280581e-08, 3.231275e-08, 3.190654e-08, 3.146928e-08, 
    3.174416e-08, 3.19578e-08, 3.211117e-08, 3.187121e-08, 3.22732e-08, 
    3.261734e-08, 3.17833e-08, 3.145889e-08, 3.158938e-08, 3.183482e-08,
  3.103376e-08, 3.191631e-08, 3.216369e-08, 3.213872e-08, 3.235296e-08, 
    3.290904e-08, 3.266329e-08, 3.241248e-08, 3.276697e-08, 3.245934e-08, 
    3.267026e-08, 3.141841e-08, 3.112501e-08, 3.113612e-08, 3.131534e-08,
  3.021062e-08, 3.04015e-08, 3.04173e-08, 3.079476e-08, 3.197468e-08, 
    3.250613e-08, 3.327215e-08, 3.223587e-08, 3.254298e-08, 3.250944e-08, 
    3.184264e-08, 3.065994e-08, 3.158357e-08, 3.148843e-08, 3.049967e-08,
  2.956466e-08, 3.001106e-08, 3.031982e-08, 3.125691e-08, 3.143042e-08, 
    3.182862e-08, 3.142495e-08, 3.089135e-08, 2.988331e-08, 3.098419e-08, 
    3.084494e-08, 3.060361e-08, 3.172316e-08, 3.053836e-08, 3.057566e-08,
  2.969939e-08, 3.021036e-08, 3.079013e-08, 3.078629e-08, 3.103837e-08, 
    3.004022e-08, 2.91289e-08, 2.818572e-08, 2.816305e-08, 2.543716e-08, 
    2.695816e-08, 2.968027e-08, 3.191737e-08, 3.057498e-08, 3.011042e-08,
  3.071342e-08, 3.011323e-08, 2.936171e-08, 2.921382e-08, 2.921492e-08, 
    2.929859e-08, 2.861456e-08, 2.474069e-08, 2.413491e-08, 2.670406e-08, 
    2.772919e-08, 3.069246e-08, 3.256356e-08, 3.033037e-08, 2.994145e-08,
  2.692754e-08, 2.723415e-08, 2.709762e-08, 2.796945e-08, 2.890106e-08, 
    2.860126e-08, 2.857389e-08, 2.671291e-08, 2.43015e-08, 2.575777e-08, 
    2.74009e-08, 3.228041e-08, 3.239307e-08, 3.007225e-08, 3.086109e-08,
  2.710503e-08, 2.790139e-08, 2.850385e-08, 2.961827e-08, 3.066311e-08, 
    3.045646e-08, 2.96099e-08, 2.827691e-08, 2.574631e-08, 2.548595e-08, 
    2.877628e-08, 3.378099e-08, 3.229977e-08, 3.073498e-08, 2.947264e-08,
  3.11398e-08, 3.009578e-08, 2.94369e-08, 3.027914e-08, 3.053974e-08, 
    3.176299e-08, 3.061935e-08, 2.893509e-08, 2.675762e-08, 2.63512e-08, 
    3.083809e-08, 3.473137e-08, 3.239138e-08, 2.99053e-08, 2.642722e-08,
  2.79958e-08, 2.910292e-08, 2.890127e-08, 3.00821e-08, 2.991376e-08, 
    3.070017e-08, 3.010683e-08, 2.92875e-08, 2.75918e-08, 2.805456e-08, 
    3.397965e-08, 3.52115e-08, 3.175091e-08, 2.658263e-08, 2.852783e-08,
  2.814966e-08, 2.974767e-08, 3.037241e-08, 3.154075e-08, 3.185507e-08, 
    3.2362e-08, 3.174157e-08, 3.111279e-08, 3.004185e-08, 2.941848e-08, 
    2.89861e-08, 2.900224e-08, 3.048386e-08, 3.201048e-08, 3.120169e-08,
  2.784973e-08, 2.920347e-08, 3.026282e-08, 3.096054e-08, 3.05772e-08, 
    3.122729e-08, 3.101619e-08, 3.10689e-08, 3.015836e-08, 2.898489e-08, 
    2.885387e-08, 2.934575e-08, 3.132519e-08, 3.113091e-08, 3.039287e-08,
  2.74662e-08, 2.886529e-08, 2.993699e-08, 2.948832e-08, 2.942099e-08, 
    3.044719e-08, 3.177342e-08, 3.187415e-08, 3.089381e-08, 2.96443e-08, 
    2.959631e-08, 3.006949e-08, 3.097859e-08, 3.001306e-08, 3.041417e-08,
  2.858133e-08, 2.789982e-08, 2.880764e-08, 2.882454e-08, 2.96671e-08, 
    2.904774e-08, 3.063527e-08, 3.155319e-08, 3.081866e-08, 3.022972e-08, 
    2.993123e-08, 3.093551e-08, 3.047439e-08, 2.939289e-08, 2.95418e-08,
  2.913681e-08, 2.822364e-08, 2.797084e-08, 2.816664e-08, 2.911258e-08, 
    2.932635e-08, 2.921073e-08, 3.0198e-08, 3.070009e-08, 3.067744e-08, 
    3.027433e-08, 2.975367e-08, 2.903623e-08, 2.902274e-08, 2.913831e-08,
  2.991043e-08, 2.909059e-08, 2.799287e-08, 2.777246e-08, 2.830655e-08, 
    2.922533e-08, 2.939759e-08, 2.863809e-08, 2.88607e-08, 3.014947e-08, 
    3.015776e-08, 2.91775e-08, 2.849616e-08, 2.868879e-08, 2.893267e-08,
  3.049703e-08, 3.129142e-08, 3.084756e-08, 2.954968e-08, 2.917412e-08, 
    2.896399e-08, 2.874507e-08, 2.842946e-08, 2.829449e-08, 2.876674e-08, 
    2.850951e-08, 2.780567e-08, 2.768271e-08, 2.868445e-08, 2.934114e-08,
  2.508627e-08, 2.7898e-08, 2.948862e-08, 2.952489e-08, 2.939586e-08, 
    2.894451e-08, 2.856031e-08, 2.861723e-08, 2.83433e-08, 2.815546e-08, 
    2.762617e-08, 2.729142e-08, 2.789177e-08, 2.849419e-08, 2.948139e-08,
  2.716858e-08, 2.676356e-08, 2.802242e-08, 2.879923e-08, 2.906755e-08, 
    2.855432e-08, 2.847221e-08, 2.808137e-08, 2.787021e-08, 2.756885e-08, 
    2.610257e-08, 2.649081e-08, 2.839509e-08, 2.87407e-08, 3.01308e-08,
  3.193288e-08, 2.998219e-08, 2.905766e-08, 2.921055e-08, 2.931865e-08, 
    2.921081e-08, 2.90837e-08, 2.84477e-08, 2.785458e-08, 2.652444e-08, 
    2.591135e-08, 2.821082e-08, 2.85758e-08, 2.95744e-08, 2.914137e-08,
  3.181338e-08, 3.161432e-08, 3.179102e-08, 3.04241e-08, 2.873092e-08, 
    2.894277e-08, 3.208191e-08, 3.056212e-08, 3.214281e-08, 3.181277e-08, 
    3.161846e-08, 2.884852e-08, 2.64502e-08, 2.633078e-08, 2.82143e-08,
  3.178331e-08, 3.152299e-08, 3.149168e-08, 3.077727e-08, 2.971348e-08, 
    2.967209e-08, 2.830926e-08, 3.104634e-08, 3.080563e-08, 3.031015e-08, 
    2.966319e-08, 2.7091e-08, 2.717748e-08, 2.899882e-08, 3.071399e-08,
  3.179552e-08, 3.090308e-08, 3.104409e-08, 3.007285e-08, 2.889421e-08, 
    3.091131e-08, 2.840267e-08, 2.84283e-08, 2.921364e-08, 2.785262e-08, 
    2.721343e-08, 2.702181e-08, 2.8895e-08, 3.006229e-08, 3.174867e-08,
  3.191993e-08, 3.137642e-08, 3.098283e-08, 2.976425e-08, 3.078824e-08, 
    3.117913e-08, 3.073295e-08, 3.01506e-08, 2.918284e-08, 2.748503e-08, 
    2.822349e-08, 2.999023e-08, 3.13398e-08, 3.275228e-08, 3.311895e-08,
  3.228492e-08, 3.195322e-08, 3.124403e-08, 2.947794e-08, 2.996958e-08, 
    2.997561e-08, 3.017248e-08, 3.12346e-08, 3.110713e-08, 3.007743e-08, 
    3.053131e-08, 3.220202e-08, 3.244871e-08, 3.206259e-08, 2.955428e-08,
  3.285013e-08, 3.239485e-08, 3.108303e-08, 2.948345e-08, 2.973634e-08, 
    2.985436e-08, 2.9781e-08, 2.959812e-08, 2.958722e-08, 3.164997e-08, 
    3.288494e-08, 3.242658e-08, 3.157977e-08, 2.912907e-08, 2.70879e-08,
  3.260341e-08, 3.123889e-08, 3.101304e-08, 3.03938e-08, 2.967847e-08, 
    2.924176e-08, 2.944733e-08, 2.908812e-08, 3.051889e-08, 3.072192e-08, 
    3.043793e-08, 2.999908e-08, 2.887205e-08, 2.649053e-08, 2.770225e-08,
  3.132076e-08, 2.96726e-08, 2.990394e-08, 3.039689e-08, 2.958016e-08, 
    2.887452e-08, 2.822113e-08, 2.825449e-08, 2.865693e-08, 2.900766e-08, 
    2.895681e-08, 2.932617e-08, 2.652442e-08, 2.671559e-08, 2.931666e-08,
  3.203642e-08, 3.060082e-08, 2.949711e-08, 2.984113e-08, 2.959475e-08, 
    2.951712e-08, 2.883637e-08, 2.868855e-08, 2.890068e-08, 2.905795e-08, 
    2.900363e-08, 2.684701e-08, 2.610113e-08, 2.830768e-08, 2.973776e-08,
  3.276981e-08, 3.171363e-08, 2.955614e-08, 2.821431e-08, 2.813599e-08, 
    2.876427e-08, 2.871056e-08, 2.881616e-08, 2.862626e-08, 2.799296e-08, 
    2.758991e-08, 2.602762e-08, 2.707047e-08, 3.006538e-08, 2.909518e-08,
  2.098579e-08, 2.191387e-08, 2.419731e-08, 2.578508e-08, 2.785293e-08, 
    2.860723e-08, 2.867426e-08, 2.942478e-08, 3.087844e-08, 3.247131e-08, 
    3.03214e-08, 2.991089e-08, 2.918775e-08, 2.857724e-08, 2.697614e-08,
  2.086051e-08, 2.172567e-08, 2.381614e-08, 2.565035e-08, 2.674447e-08, 
    2.801244e-08, 2.805402e-08, 2.910389e-08, 2.94495e-08, 2.953087e-08, 
    2.954594e-08, 2.907628e-08, 2.896357e-08, 2.939343e-08, 3.030656e-08,
  2.208099e-08, 2.299199e-08, 2.465164e-08, 2.586215e-08, 2.666713e-08, 
    2.817973e-08, 2.752099e-08, 2.834665e-08, 2.92298e-08, 2.86083e-08, 
    2.852953e-08, 2.86892e-08, 2.916319e-08, 3.0207e-08, 3.152904e-08,
  2.534456e-08, 2.600145e-08, 2.695807e-08, 2.746618e-08, 2.770964e-08, 
    2.79834e-08, 2.820932e-08, 2.905378e-08, 3.002205e-08, 2.918257e-08, 
    2.967488e-08, 3.060433e-08, 3.129773e-08, 3.28419e-08, 3.243324e-08,
  2.984829e-08, 2.977706e-08, 2.96987e-08, 2.890702e-08, 2.93527e-08, 
    2.824345e-08, 2.82436e-08, 3.057582e-08, 3.032158e-08, 3.020023e-08, 
    3.110054e-08, 3.12925e-08, 3.103669e-08, 3.083388e-08, 2.958926e-08,
  3.056518e-08, 3.04237e-08, 3.029441e-08, 2.985078e-08, 2.955442e-08, 
    2.967815e-08, 2.900441e-08, 2.872801e-08, 2.945747e-08, 3.168228e-08, 
    3.097397e-08, 3.012749e-08, 2.982819e-08, 2.880761e-08, 2.785007e-08,
  3.255169e-08, 3.240686e-08, 3.21044e-08, 3.132935e-08, 3.051663e-08, 
    3.139911e-08, 3.063744e-08, 2.988423e-08, 3.088379e-08, 3.110397e-08, 
    2.985631e-08, 2.980843e-08, 2.914695e-08, 2.80964e-08, 2.964017e-08,
  3.138662e-08, 3.091611e-08, 3.069746e-08, 3.076053e-08, 3.160269e-08, 
    3.273984e-08, 3.167111e-08, 3.071475e-08, 3.078446e-08, 3.014328e-08, 
    3.024275e-08, 2.941044e-08, 2.817387e-08, 2.896098e-08, 3.066386e-08,
  3.076377e-08, 3.037274e-08, 3.033445e-08, 3.138277e-08, 3.265829e-08, 
    3.248924e-08, 3.113523e-08, 3.078775e-08, 3.10114e-08, 3.05248e-08, 
    2.975066e-08, 2.786913e-08, 2.822147e-08, 2.973114e-08, 3.088528e-08,
  3.042479e-08, 3.056842e-08, 3.063395e-08, 3.096359e-08, 3.110059e-08, 
    3.075824e-08, 2.966202e-08, 2.978521e-08, 3.033141e-08, 2.96482e-08, 
    2.827631e-08, 2.717886e-08, 2.884238e-08, 3.004041e-08, 3.163686e-08,
  2.415171e-08, 2.256135e-08, 2.144222e-08, 2.099011e-08, 2.123135e-08, 
    2.211712e-08, 2.316492e-08, 2.410184e-08, 2.504214e-08, 2.599628e-08, 
    2.694425e-08, 2.808882e-08, 2.856922e-08, 2.898599e-08, 2.953782e-08,
  2.322048e-08, 2.232966e-08, 2.20972e-08, 2.274896e-08, 2.406085e-08, 
    2.540129e-08, 2.584273e-08, 2.62715e-08, 2.658037e-08, 2.668714e-08, 
    2.768537e-08, 2.880791e-08, 2.930005e-08, 2.902513e-08, 2.940453e-08,
  2.350527e-08, 2.404587e-08, 2.52309e-08, 2.685958e-08, 2.847853e-08, 
    2.926351e-08, 2.892147e-08, 2.812118e-08, 2.76856e-08, 2.796888e-08, 
    2.859806e-08, 2.968157e-08, 2.983969e-08, 2.963898e-08, 3.016816e-08,
  2.627369e-08, 2.792146e-08, 2.926331e-08, 3.106659e-08, 3.092356e-08, 
    3.132933e-08, 3.132656e-08, 3.044545e-08, 2.961083e-08, 2.907545e-08, 
    2.957507e-08, 3.044325e-08, 3.079485e-08, 3.052606e-08, 3.019278e-08,
  2.913891e-08, 3.084558e-08, 3.209086e-08, 3.232689e-08, 3.343398e-08, 
    3.264577e-08, 3.270095e-08, 3.203191e-08, 3.229363e-08, 3.07919e-08, 
    3.056782e-08, 3.110614e-08, 3.109533e-08, 3.065206e-08, 3.022049e-08,
  3.145953e-08, 3.215147e-08, 3.288326e-08, 3.374458e-08, 3.317258e-08, 
    3.272174e-08, 3.201559e-08, 3.051546e-08, 2.967324e-08, 3.169191e-08, 
    3.235181e-08, 3.244967e-08, 3.194266e-08, 3.06727e-08, 3.026033e-08,
  3.288959e-08, 3.365488e-08, 3.29781e-08, 3.170654e-08, 3.148956e-08, 
    3.124335e-08, 3.119217e-08, 3.059021e-08, 3.039464e-08, 3.068478e-08, 
    3.075733e-08, 3.084696e-08, 3.007807e-08, 2.946252e-08, 2.975705e-08,
  3.398576e-08, 3.306593e-08, 3.191912e-08, 3.065501e-08, 3.063744e-08, 
    3.054735e-08, 3.055624e-08, 3.02775e-08, 3.018724e-08, 2.972665e-08, 
    3.013797e-08, 3.053099e-08, 2.984074e-08, 2.966294e-08, 3.040272e-08,
  3.206667e-08, 2.983845e-08, 2.896126e-08, 2.850915e-08, 2.882348e-08, 
    2.961552e-08, 3.088766e-08, 3.051786e-08, 3.058193e-08, 3.064923e-08, 
    3.113927e-08, 3.01421e-08, 2.993103e-08, 2.970881e-08, 3.051251e-08,
  2.812161e-08, 2.752974e-08, 2.791241e-08, 2.895775e-08, 2.979803e-08, 
    2.96131e-08, 3.029324e-08, 2.964189e-08, 2.908396e-08, 3.052743e-08, 
    3.082588e-08, 3.021336e-08, 3.012617e-08, 3.022645e-08, 3.102262e-08,
  2.743903e-08, 2.770383e-08, 2.655379e-08, 2.527331e-08, 2.442356e-08, 
    2.409223e-08, 2.424851e-08, 2.438301e-08, 2.492677e-08, 2.63225e-08, 
    2.780257e-08, 2.908849e-08, 3.02432e-08, 3.018305e-08, 2.9879e-08,
  2.653618e-08, 2.606317e-08, 2.562023e-08, 2.481048e-08, 2.531144e-08, 
    2.543477e-08, 2.49108e-08, 2.545665e-08, 2.657757e-08, 2.770784e-08, 
    2.928426e-08, 3.04441e-08, 3.149065e-08, 3.114733e-08, 2.988957e-08,
  2.556676e-08, 2.548645e-08, 2.548702e-08, 2.517219e-08, 2.553668e-08, 
    2.561188e-08, 2.569024e-08, 2.7004e-08, 2.824529e-08, 2.972953e-08, 
    3.094507e-08, 3.136376e-08, 3.135201e-08, 3.056651e-08, 3.036223e-08,
  2.531836e-08, 2.527491e-08, 2.504501e-08, 2.515793e-08, 2.52854e-08, 
    2.61631e-08, 2.794035e-08, 2.917322e-08, 3.108396e-08, 3.13e-08, 
    3.174437e-08, 3.15258e-08, 3.124214e-08, 3.101556e-08, 3.04694e-08,
  2.452192e-08, 2.457246e-08, 2.514936e-08, 2.622236e-08, 2.758148e-08, 
    2.854403e-08, 3.010331e-08, 3.173197e-08, 3.217855e-08, 3.19594e-08, 
    3.195656e-08, 3.158925e-08, 3.118177e-08, 3.110484e-08, 3.024549e-08,
  2.534712e-08, 2.631044e-08, 2.751144e-08, 2.877249e-08, 2.993877e-08, 
    3.160265e-08, 3.300349e-08, 3.25749e-08, 3.263109e-08, 3.36837e-08, 
    3.351844e-08, 3.29448e-08, 3.252053e-08, 3.1921e-08, 3.120823e-08,
  2.813177e-08, 2.870423e-08, 2.989567e-08, 3.117285e-08, 3.23616e-08, 
    3.319368e-08, 3.386139e-08, 3.291541e-08, 3.141258e-08, 3.062534e-08, 
    2.97345e-08, 2.983677e-08, 2.99288e-08, 2.982677e-08, 2.965338e-08,
  2.945042e-08, 3.079065e-08, 3.146687e-08, 3.179327e-08, 3.137841e-08, 
    3.090338e-08, 3.04513e-08, 2.963935e-08, 2.920192e-08, 2.866693e-08, 
    2.846757e-08, 2.84752e-08, 2.863359e-08, 2.880733e-08, 2.961141e-08,
  3.110894e-08, 3.157703e-08, 3.06515e-08, 2.997229e-08, 2.964305e-08, 
    2.930349e-08, 2.903623e-08, 2.847374e-08, 2.855997e-08, 2.894798e-08, 
    2.89213e-08, 2.876958e-08, 2.928403e-08, 2.927615e-08, 2.913466e-08,
  3.058106e-08, 2.963178e-08, 2.887883e-08, 2.868173e-08, 2.896228e-08, 
    2.84624e-08, 2.821213e-08, 2.836582e-08, 2.885348e-08, 2.705593e-08, 
    2.830662e-08, 2.936553e-08, 2.994234e-08, 2.947675e-08, 2.937135e-08,
  3.449478e-08, 3.406345e-08, 3.355748e-08, 3.232542e-08, 3.067747e-08, 
    2.897971e-08, 2.737531e-08, 2.608349e-08, 2.49771e-08, 2.398743e-08, 
    2.319534e-08, 2.291129e-08, 2.350662e-08, 2.419175e-08, 2.487643e-08,
  3.243364e-08, 3.270382e-08, 3.237252e-08, 3.205792e-08, 3.099449e-08, 
    3.088566e-08, 2.91766e-08, 2.765608e-08, 2.618104e-08, 2.472535e-08, 
    2.407595e-08, 2.378324e-08, 2.465809e-08, 2.492351e-08, 2.616387e-08,
  2.900815e-08, 2.930756e-08, 2.960656e-08, 2.858893e-08, 2.896697e-08, 
    2.815503e-08, 2.78609e-08, 2.716908e-08, 2.659555e-08, 2.60722e-08, 
    2.606789e-08, 2.635099e-08, 2.652772e-08, 2.644141e-08, 2.745766e-08,
  2.755963e-08, 2.812029e-08, 2.825196e-08, 2.845207e-08, 2.831479e-08, 
    2.812837e-08, 2.771383e-08, 2.77847e-08, 2.796219e-08, 2.729064e-08, 
    2.73492e-08, 2.835151e-08, 2.851029e-08, 2.846126e-08, 2.892559e-08,
  2.676488e-08, 2.729441e-08, 2.766405e-08, 2.804702e-08, 2.800822e-08, 
    2.776403e-08, 2.731836e-08, 2.774008e-08, 2.85974e-08, 2.839518e-08, 
    2.851388e-08, 2.923968e-08, 2.983717e-08, 3.054145e-08, 3.026815e-08,
  2.597942e-08, 2.557046e-08, 2.562163e-08, 2.601525e-08, 2.680492e-08, 
    2.712028e-08, 2.764748e-08, 2.735995e-08, 2.729289e-08, 2.903013e-08, 
    2.992896e-08, 3.072787e-08, 3.103818e-08, 3.063715e-08, 2.991598e-08,
  2.687449e-08, 2.596459e-08, 2.510918e-08, 2.454857e-08, 2.408523e-08, 
    2.431055e-08, 2.484805e-08, 2.604103e-08, 2.754552e-08, 2.939491e-08, 
    3.040958e-08, 3.058424e-08, 3.002884e-08, 2.920741e-08, 2.839816e-08,
  2.846842e-08, 2.791629e-08, 2.69581e-08, 2.627031e-08, 2.57701e-08, 
    2.566811e-08, 2.613017e-08, 2.720435e-08, 2.832649e-08, 2.887805e-08, 
    2.93388e-08, 2.893424e-08, 2.839364e-08, 2.787015e-08, 2.792669e-08,
  2.895072e-08, 2.910004e-08, 2.91973e-08, 2.909362e-08, 2.906419e-08, 
    2.907607e-08, 2.958213e-08, 2.962216e-08, 2.978078e-08, 2.997799e-08, 
    2.997852e-08, 2.957487e-08, 2.923403e-08, 2.92428e-08, 2.984036e-08,
  2.916179e-08, 2.909603e-08, 2.911858e-08, 2.909083e-08, 2.93269e-08, 
    2.967123e-08, 3.022066e-08, 2.966757e-08, 3.062179e-08, 3.086814e-08, 
    3.088283e-08, 3.021465e-08, 2.975306e-08, 2.974888e-08, 2.968722e-08,
  3.009568e-08, 3.086636e-08, 3.17527e-08, 3.224504e-08, 3.2223e-08, 
    3.232811e-08, 3.215775e-08, 3.296277e-08, 3.355197e-08, 3.546767e-08, 
    3.581731e-08, 3.550947e-08, 3.522555e-08, 3.354493e-08, 3.194931e-08,
  3.042311e-08, 3.09477e-08, 3.153763e-08, 3.160658e-08, 3.181145e-08, 
    3.165332e-08, 3.120656e-08, 3.164561e-08, 3.244672e-08, 3.214792e-08, 
    3.232535e-08, 3.317545e-08, 3.314858e-08, 3.260223e-08, 3.132545e-08,
  2.931684e-08, 2.958115e-08, 3.004975e-08, 2.986988e-08, 3.016719e-08, 
    2.978646e-08, 3.018323e-08, 3.00185e-08, 3.028854e-08, 3.058814e-08, 
    3.075556e-08, 3.026835e-08, 3.020168e-08, 3.005555e-08, 2.991408e-08,
  2.926746e-08, 2.92638e-08, 2.884855e-08, 2.866147e-08, 2.82601e-08, 
    2.91861e-08, 2.999681e-08, 2.945269e-08, 2.940818e-08, 2.919425e-08, 
    2.926228e-08, 2.904565e-08, 2.943001e-08, 2.988632e-08, 3.022756e-08,
  2.9294e-08, 2.932054e-08, 2.926492e-08, 2.934876e-08, 2.948253e-08, 
    2.962262e-08, 2.920282e-08, 3.093916e-08, 3.034088e-08, 2.962555e-08, 
    2.998145e-08, 3.007882e-08, 2.984509e-08, 3.030431e-08, 3.116484e-08,
  3.065125e-08, 3.032055e-08, 3.023765e-08, 3.015913e-08, 3.026934e-08, 
    3.035318e-08, 3.011161e-08, 2.933553e-08, 2.903392e-08, 2.898751e-08, 
    2.871846e-08, 2.81609e-08, 2.861456e-08, 2.935153e-08, 3.011606e-08,
  3.190711e-08, 3.154943e-08, 3.134033e-08, 3.10868e-08, 3.073103e-08, 
    3.05358e-08, 2.990777e-08, 2.890883e-08, 2.823296e-08, 2.781835e-08, 
    2.793678e-08, 2.819487e-08, 2.912817e-08, 2.963921e-08, 2.980462e-08,
  2.836968e-08, 2.863758e-08, 2.872995e-08, 2.87377e-08, 2.866806e-08, 
    2.86022e-08, 2.851193e-08, 2.845225e-08, 2.811428e-08, 2.793443e-08, 
    2.738132e-08, 2.717568e-08, 2.700619e-08, 2.745569e-08, 2.777912e-08,
  2.818126e-08, 2.840883e-08, 2.847501e-08, 2.87072e-08, 2.884002e-08, 
    2.904889e-08, 2.90702e-08, 2.908608e-08, 2.885091e-08, 2.867439e-08, 
    2.830779e-08, 2.73389e-08, 2.695871e-08, 2.623176e-08, 2.588686e-08,
  2.912517e-08, 2.920285e-08, 2.931987e-08, 2.935278e-08, 2.951147e-08, 
    2.935962e-08, 2.962064e-08, 2.935284e-08, 2.95178e-08, 2.939475e-08, 
    2.968038e-08, 2.914268e-08, 2.859744e-08, 2.792807e-08, 2.678544e-08,
  2.548163e-08, 2.537375e-08, 2.626343e-08, 2.662396e-08, 2.660379e-08, 
    2.653718e-08, 2.467961e-08, 2.309826e-08, 2.283882e-08, 2.357782e-08, 
    2.634897e-08, 2.887104e-08, 3.068498e-08, 3.342232e-08, 3.218997e-08,
  2.565553e-08, 2.557869e-08, 2.558783e-08, 2.658387e-08, 2.630796e-08, 
    2.660197e-08, 2.597361e-08, 2.492734e-08, 2.497597e-08, 2.552784e-08, 
    2.749998e-08, 2.846527e-08, 3.109154e-08, 3.080762e-08, 3.134634e-08,
  2.649126e-08, 2.615543e-08, 2.656301e-08, 2.660166e-08, 2.744632e-08, 
    2.764278e-08, 2.641861e-08, 2.651799e-08, 2.605253e-08, 2.663e-08, 
    2.751781e-08, 2.885854e-08, 2.959458e-08, 3.013696e-08, 3.157156e-08,
  2.69562e-08, 2.73865e-08, 2.729683e-08, 2.7731e-08, 2.686572e-08, 
    2.689861e-08, 2.672844e-08, 2.679511e-08, 2.702592e-08, 2.657318e-08, 
    2.751441e-08, 2.882466e-08, 2.982161e-08, 3.11718e-08, 3.094165e-08,
  2.651443e-08, 2.772722e-08, 2.816813e-08, 2.803814e-08, 2.818766e-08, 
    2.697917e-08, 2.751777e-08, 2.832642e-08, 2.87505e-08, 2.767745e-08, 
    2.883573e-08, 3.026474e-08, 3.058447e-08, 3.045225e-08, 2.964222e-08,
  2.605595e-08, 2.640698e-08, 2.726013e-08, 2.737316e-08, 2.769888e-08, 
    2.751255e-08, 2.726266e-08, 2.675597e-08, 2.689626e-08, 2.874335e-08, 
    3.02034e-08, 3.025797e-08, 2.962126e-08, 2.90114e-08, 2.946176e-08,
  2.751565e-08, 2.703638e-08, 2.72266e-08, 2.778883e-08, 2.826989e-08, 
    2.860614e-08, 2.898528e-08, 2.904861e-08, 2.960977e-08, 2.994982e-08, 
    3.023159e-08, 2.987448e-08, 2.922833e-08, 2.916414e-08, 2.914961e-08,
  2.967239e-08, 2.933511e-08, 2.909299e-08, 2.908322e-08, 2.929562e-08, 
    2.953644e-08, 2.972102e-08, 2.97301e-08, 2.990407e-08, 2.948398e-08, 
    2.95662e-08, 2.926379e-08, 2.895015e-08, 2.86615e-08, 2.871809e-08,
  2.994288e-08, 2.967658e-08, 2.966232e-08, 2.952244e-08, 2.947075e-08, 
    2.947284e-08, 2.9658e-08, 2.974183e-08, 2.982905e-08, 2.986541e-08, 
    2.972964e-08, 2.90457e-08, 2.902418e-08, 2.835487e-08, 2.849735e-08,
  2.985641e-08, 2.986965e-08, 2.983345e-08, 2.991942e-08, 2.989496e-08, 
    2.997515e-08, 2.989405e-08, 2.988513e-08, 2.984094e-08, 2.972638e-08, 
    2.930243e-08, 2.877193e-08, 2.817825e-08, 2.851583e-08, 2.765599e-08,
  2.8983e-08, 2.803065e-08, 2.808484e-08, 2.700992e-08, 2.471309e-08, 
    2.384814e-08, 2.420842e-08, 2.367145e-08, 2.404176e-08, 2.356889e-08, 
    2.281665e-08, 2.20299e-08, 2.254692e-08, 2.33353e-08, 2.404987e-08,
  2.931301e-08, 2.845873e-08, 2.812784e-08, 2.8452e-08, 2.561755e-08, 
    2.456599e-08, 2.428052e-08, 2.362598e-08, 2.35177e-08, 2.22659e-08, 
    2.182527e-08, 2.168429e-08, 2.276547e-08, 2.334733e-08, 2.447111e-08,
  2.91229e-08, 2.877183e-08, 2.846489e-08, 2.845338e-08, 2.787637e-08, 
    2.538469e-08, 2.532084e-08, 2.467657e-08, 2.45305e-08, 2.345473e-08, 
    2.259431e-08, 2.273712e-08, 2.336229e-08, 2.43408e-08, 2.48915e-08,
  2.924191e-08, 2.881439e-08, 2.865766e-08, 2.872329e-08, 2.809078e-08, 
    2.700562e-08, 2.512528e-08, 2.562389e-08, 2.616175e-08, 2.538557e-08, 
    2.531999e-08, 2.576612e-08, 2.553067e-08, 2.483525e-08, 2.488362e-08,
  2.927317e-08, 2.874923e-08, 2.846121e-08, 2.901094e-08, 2.89392e-08, 
    2.790668e-08, 2.678346e-08, 2.556492e-08, 2.560886e-08, 2.423169e-08, 
    2.430505e-08, 2.409741e-08, 2.380578e-08, 2.412465e-08, 2.545563e-08,
  2.882326e-08, 2.891771e-08, 2.840921e-08, 2.872061e-08, 2.921598e-08, 
    2.883531e-08, 2.828947e-08, 2.666589e-08, 2.592193e-08, 2.56896e-08, 
    2.521971e-08, 2.493888e-08, 2.491852e-08, 2.55834e-08, 2.631105e-08,
  2.791137e-08, 2.814537e-08, 2.823184e-08, 2.772419e-08, 2.856879e-08, 
    2.854973e-08, 2.88443e-08, 2.793524e-08, 2.690809e-08, 2.682862e-08, 
    2.58217e-08, 2.571037e-08, 2.55697e-08, 2.577546e-08, 2.61338e-08,
  2.781558e-08, 2.777536e-08, 2.802747e-08, 2.750076e-08, 2.754972e-08, 
    2.756483e-08, 2.770622e-08, 2.810809e-08, 2.769223e-08, 2.682752e-08, 
    2.610951e-08, 2.573946e-08, 2.56194e-08, 2.577787e-08, 2.670435e-08,
  2.794156e-08, 2.768061e-08, 2.777143e-08, 2.761523e-08, 2.706108e-08, 
    2.671764e-08, 2.6749e-08, 2.673635e-08, 2.660598e-08, 2.666381e-08, 
    2.661982e-08, 2.617166e-08, 2.615936e-08, 2.668284e-08, 2.75177e-08,
  3.161915e-08, 2.921653e-08, 2.829493e-08, 2.789102e-08, 2.759034e-08, 
    2.680633e-08, 2.654023e-08, 2.659624e-08, 2.668387e-08, 2.672255e-08, 
    2.675917e-08, 2.662325e-08, 2.70291e-08, 2.721379e-08, 2.732019e-08,
  3.210391e-08, 3.063131e-08, 2.939664e-08, 2.834106e-08, 2.616228e-08, 
    2.456137e-08, 2.491387e-08, 2.581744e-08, 2.58695e-08, 2.649627e-08, 
    2.662073e-08, 2.648335e-08, 2.598801e-08, 2.603763e-08, 2.570151e-08,
  3.362729e-08, 3.217103e-08, 3.035572e-08, 3.034948e-08, 2.797942e-08, 
    2.61666e-08, 2.482007e-08, 2.476607e-08, 2.514952e-08, 2.544906e-08, 
    2.639516e-08, 2.608866e-08, 2.560137e-08, 2.521865e-08, 2.504324e-08,
  3.469792e-08, 3.418506e-08, 3.239978e-08, 3.076591e-08, 3.041849e-08, 
    2.726658e-08, 2.670195e-08, 2.542946e-08, 2.50602e-08, 2.525486e-08, 
    2.557119e-08, 2.499295e-08, 2.419205e-08, 2.415672e-08, 2.502613e-08,
  3.390546e-08, 3.514058e-08, 3.451096e-08, 3.350431e-08, 3.201468e-08, 
    3.038422e-08, 2.685865e-08, 2.757263e-08, 2.758672e-08, 2.65166e-08, 
    2.617876e-08, 2.498921e-08, 2.443188e-08, 2.472347e-08, 2.482324e-08,
  3.275469e-08, 3.434213e-08, 3.470486e-08, 3.45523e-08, 3.402702e-08, 
    3.334009e-08, 3.047019e-08, 2.713505e-08, 2.541429e-08, 2.504501e-08, 
    2.491333e-08, 2.445655e-08, 2.421186e-08, 2.440967e-08, 2.400762e-08,
  3.052564e-08, 3.291114e-08, 3.418504e-08, 3.447055e-08, 3.429304e-08, 
    3.415413e-08, 3.436933e-08, 3.070152e-08, 2.735144e-08, 2.562146e-08, 
    2.441588e-08, 2.392612e-08, 2.387264e-08, 2.386923e-08, 2.35697e-08,
  2.99015e-08, 3.055535e-08, 3.244428e-08, 3.3846e-08, 3.427179e-08, 
    3.376606e-08, 3.397011e-08, 3.457439e-08, 3.174571e-08, 2.923422e-08, 
    2.635082e-08, 2.465684e-08, 2.400271e-08, 2.36097e-08, 2.374738e-08,
  2.952049e-08, 2.9857e-08, 3.028301e-08, 3.160578e-08, 3.306997e-08, 
    3.364089e-08, 3.332059e-08, 3.332307e-08, 3.388203e-08, 3.236369e-08, 
    2.953544e-08, 2.75224e-08, 2.579013e-08, 2.498611e-08, 2.485599e-08,
  2.982359e-08, 2.93438e-08, 2.949928e-08, 3.010364e-08, 3.11444e-08, 
    3.189206e-08, 3.298003e-08, 3.276381e-08, 3.250552e-08, 3.239909e-08, 
    3.144777e-08, 2.931025e-08, 2.751617e-08, 2.597872e-08, 2.542019e-08,
  3.003975e-08, 2.942494e-08, 2.875487e-08, 2.887565e-08, 2.99935e-08, 
    3.082018e-08, 3.164389e-08, 3.226374e-08, 3.277087e-08, 3.198102e-08, 
    3.176907e-08, 3.121595e-08, 2.986487e-08, 2.776849e-08, 2.664349e-08,
  2.441174e-08, 2.286401e-08, 2.246853e-08, 2.646473e-08, 2.642772e-08, 
    2.573734e-08, 2.687567e-08, 2.934375e-08, 3.155358e-08, 3.126347e-08, 
    2.870896e-08, 2.70741e-08, 2.603885e-08, 2.607668e-08, 2.524736e-08,
  2.593085e-08, 2.376647e-08, 2.284723e-08, 2.590326e-08, 2.600712e-08, 
    2.633992e-08, 2.584579e-08, 2.868919e-08, 3.131523e-08, 3.312769e-08, 
    3.114752e-08, 2.865361e-08, 2.718627e-08, 2.623681e-08, 2.523172e-08,
  2.769985e-08, 2.543456e-08, 2.359134e-08, 2.563399e-08, 2.596859e-08, 
    2.538243e-08, 2.603459e-08, 2.779933e-08, 2.990226e-08, 3.280109e-08, 
    3.214507e-08, 2.976981e-08, 2.756514e-08, 2.608199e-08, 2.532444e-08,
  3.045476e-08, 2.77882e-08, 2.55503e-08, 2.51301e-08, 2.609608e-08, 
    2.539975e-08, 2.62666e-08, 2.781543e-08, 2.957946e-08, 3.147287e-08, 
    3.244062e-08, 3.062136e-08, 2.814669e-08, 2.662636e-08, 2.601426e-08,
  3.407158e-08, 3.031737e-08, 2.8485e-08, 2.686184e-08, 2.607892e-08, 
    2.62418e-08, 2.546076e-08, 2.670755e-08, 2.85931e-08, 2.948402e-08, 
    2.98873e-08, 3.009714e-08, 2.897113e-08, 2.771401e-08, 2.678925e-08,
  3.597837e-08, 3.412213e-08, 3.170129e-08, 2.943583e-08, 2.717788e-08, 
    2.631309e-08, 2.621944e-08, 2.512192e-08, 2.665712e-08, 2.907323e-08, 
    2.87762e-08, 2.839651e-08, 2.818025e-08, 2.761623e-08, 2.688989e-08,
  3.589199e-08, 3.65839e-08, 3.550815e-08, 3.383019e-08, 3.108096e-08, 
    2.791723e-08, 2.616519e-08, 2.561068e-08, 2.62331e-08, 2.739838e-08, 
    2.783435e-08, 2.746466e-08, 2.749906e-08, 2.754973e-08, 2.694427e-08,
  3.447903e-08, 3.591472e-08, 3.679541e-08, 3.603395e-08, 3.501747e-08, 
    3.301925e-08, 3.023004e-08, 2.770774e-08, 2.686905e-08, 2.648274e-08, 
    2.670253e-08, 2.644935e-08, 2.645645e-08, 2.649569e-08, 2.594887e-08,
  3.600826e-08, 3.562626e-08, 3.571827e-08, 3.624672e-08, 3.59461e-08, 
    3.476385e-08, 3.331177e-08, 3.170817e-08, 3.017674e-08, 2.947411e-08, 
    2.916161e-08, 2.866089e-08, 2.833793e-08, 2.782083e-08, 2.705174e-08,
  3.410367e-08, 3.613636e-08, 3.694376e-08, 3.574662e-08, 3.548015e-08, 
    3.564822e-08, 3.524343e-08, 3.427353e-08, 3.401143e-08, 3.399802e-08, 
    3.385351e-08, 3.332754e-08, 3.258634e-08, 3.111947e-08, 2.945107e-08,
  3.056116e-08, 2.963985e-08, 2.996692e-08, 2.872397e-08, 2.651377e-08, 
    2.326231e-08, 2.23872e-08, 2.152461e-08, 2.053349e-08, 1.927812e-08, 
    1.522983e-08, 1.483834e-08, 1.745819e-08, 2.334845e-08, 2.68382e-08,
  2.918487e-08, 2.880067e-08, 2.946342e-08, 2.832971e-08, 2.597591e-08, 
    2.345637e-08, 2.1704e-08, 2.109009e-08, 2.074067e-08, 2.069278e-08, 
    1.725908e-08, 1.6205e-08, 1.802328e-08, 2.177953e-08, 2.618846e-08,
  2.878255e-08, 2.792937e-08, 2.850054e-08, 2.768301e-08, 2.533947e-08, 
    2.283298e-08, 2.181113e-08, 2.141254e-08, 2.088691e-08, 2.132981e-08, 
    1.939851e-08, 1.78326e-08, 1.889296e-08, 2.12193e-08, 2.511996e-08,
  2.763744e-08, 2.740345e-08, 2.731661e-08, 2.758977e-08, 2.444386e-08, 
    2.262334e-08, 2.065324e-08, 2.112299e-08, 2.208257e-08, 2.183662e-08, 
    2.13826e-08, 2.074424e-08, 2.076362e-08, 2.203512e-08, 2.442298e-08,
  2.745721e-08, 2.754552e-08, 2.577062e-08, 2.66041e-08, 2.458369e-08, 
    2.398775e-08, 1.983138e-08, 2.205941e-08, 2.28459e-08, 2.197757e-08, 
    2.245317e-08, 2.276992e-08, 2.270425e-08, 2.372156e-08, 2.55024e-08,
  2.635585e-08, 2.79512e-08, 2.566527e-08, 2.589614e-08, 2.475713e-08, 
    2.464068e-08, 2.397577e-08, 2.315912e-08, 2.222789e-08, 2.217472e-08, 
    2.321822e-08, 2.391468e-08, 2.45682e-08, 2.539193e-08, 2.619603e-08,
  2.646824e-08, 2.754406e-08, 2.604421e-08, 2.525533e-08, 2.451726e-08, 
    2.429987e-08, 2.558539e-08, 2.47805e-08, 2.321223e-08, 2.321854e-08, 
    2.394607e-08, 2.525586e-08, 2.632046e-08, 2.729878e-08, 2.760988e-08,
  2.802765e-08, 2.785102e-08, 2.742221e-08, 2.541465e-08, 2.445303e-08, 
    2.409142e-08, 2.486835e-08, 2.590796e-08, 2.469792e-08, 2.369336e-08, 
    2.377374e-08, 2.480656e-08, 2.603384e-08, 2.719186e-08, 2.776561e-08,
  3.199679e-08, 2.819102e-08, 2.806315e-08, 2.793296e-08, 2.55629e-08, 
    2.44699e-08, 2.399502e-08, 2.520976e-08, 2.480952e-08, 2.407288e-08, 
    2.380982e-08, 2.449767e-08, 2.542535e-08, 2.642441e-08, 2.716246e-08,
  3.699081e-08, 3.297781e-08, 2.912598e-08, 2.805689e-08, 2.844221e-08, 
    2.781337e-08, 2.608514e-08, 2.549926e-08, 2.606349e-08, 2.566137e-08, 
    2.46326e-08, 2.440573e-08, 2.48029e-08, 2.545037e-08, 2.599762e-08,
  3.338124e-08, 3.048969e-08, 3.089513e-08, 3.310792e-08, 3.319752e-08, 
    3.140012e-08, 2.749989e-08, 2.169222e-08, 2.065906e-08, 2.117875e-08, 
    2.293633e-08, 2.434937e-08, 2.688718e-08, 2.871604e-08, 3.024612e-08,
  3.361362e-08, 3.104332e-08, 3.099319e-08, 3.318072e-08, 3.323268e-08, 
    3.199893e-08, 2.697048e-08, 2.138905e-08, 2.098873e-08, 2.117457e-08, 
    2.138062e-08, 2.182712e-08, 2.408227e-08, 2.619469e-08, 2.800313e-08,
  3.291004e-08, 3.156881e-08, 3.09734e-08, 3.274228e-08, 3.226141e-08, 
    3.223417e-08, 2.807461e-08, 2.15405e-08, 2.057411e-08, 2.056432e-08, 
    1.962622e-08, 1.940578e-08, 2.187486e-08, 2.410324e-08, 2.639921e-08,
  3.161505e-08, 3.203192e-08, 3.099656e-08, 3.254517e-08, 3.191036e-08, 
    3.187236e-08, 2.710824e-08, 2.290712e-08, 2.121008e-08, 2.033214e-08, 
    1.837028e-08, 1.804958e-08, 2.00346e-08, 2.226242e-08, 2.557688e-08,
  3.031941e-08, 3.25219e-08, 3.089426e-08, 3.176211e-08, 3.229948e-08, 
    3.220705e-08, 2.617648e-08, 2.163061e-08, 2.12311e-08, 1.997838e-08, 
    1.731865e-08, 1.69073e-08, 1.861416e-08, 2.004785e-08, 2.300168e-08,
  2.951684e-08, 3.242127e-08, 3.095683e-08, 3.086064e-08, 3.150716e-08, 
    3.111693e-08, 2.754959e-08, 2.257793e-08, 2.106397e-08, 1.940917e-08, 
    1.696159e-08, 1.637188e-08, 1.75832e-08, 1.826828e-08, 2.100181e-08,
  2.853192e-08, 3.157207e-08, 3.100214e-08, 3.002791e-08, 3.080575e-08, 
    2.991109e-08, 2.977328e-08, 2.389102e-08, 2.08758e-08, 1.995772e-08, 
    1.766366e-08, 1.628182e-08, 1.734065e-08, 1.814119e-08, 2.020602e-08,
  2.971232e-08, 3.063572e-08, 3.131294e-08, 2.970493e-08, 3.035524e-08, 
    2.892479e-08, 2.916429e-08, 2.564143e-08, 2.18781e-08, 2.098518e-08, 
    1.988629e-08, 1.792769e-08, 1.784093e-08, 1.847551e-08, 1.993139e-08,
  3.049947e-08, 2.911079e-08, 3.144058e-08, 2.995884e-08, 2.993124e-08, 
    2.888492e-08, 2.823202e-08, 2.762806e-08, 2.273023e-08, 2.124208e-08, 
    2.069711e-08, 1.900204e-08, 1.825011e-08, 1.867986e-08, 1.952975e-08,
  3.376796e-08, 2.967347e-08, 3.04375e-08, 3.070971e-08, 2.96291e-08, 
    2.933334e-08, 2.799028e-08, 2.705334e-08, 2.506364e-08, 2.154471e-08, 
    2.065991e-08, 1.938708e-08, 1.896861e-08, 1.923699e-08, 1.974764e-08,
  3.114812e-08, 3.105382e-08, 3.174237e-08, 3.201535e-08, 3.071357e-08, 
    3.29044e-08, 3.365183e-08, 3.074175e-08, 2.564663e-08, 2.335449e-08, 
    2.684572e-08, 2.948291e-08, 3.113991e-08, 3.088613e-08, 3.341173e-08,
  3.223078e-08, 3.126605e-08, 3.06991e-08, 3.168029e-08, 3.123816e-08, 
    3.332451e-08, 3.216608e-08, 3.032186e-08, 2.642442e-08, 2.492573e-08, 
    2.720114e-08, 2.947526e-08, 3.137983e-08, 3.085561e-08, 3.327104e-08,
  3.256572e-08, 3.207309e-08, 3.038767e-08, 3.164086e-08, 3.165642e-08, 
    3.368394e-08, 3.258116e-08, 2.97857e-08, 2.691236e-08, 2.553802e-08, 
    2.69949e-08, 2.897514e-08, 3.127545e-08, 3.130905e-08, 3.148046e-08,
  3.255029e-08, 3.235684e-08, 3.075133e-08, 3.163385e-08, 3.207919e-08, 
    3.295149e-08, 3.137604e-08, 3.070157e-08, 2.94665e-08, 2.68636e-08, 
    2.728378e-08, 2.926461e-08, 3.126566e-08, 3.113064e-08, 2.95617e-08,
  3.190689e-08, 3.196389e-08, 3.055893e-08, 3.13967e-08, 3.252977e-08, 
    3.232566e-08, 3.008389e-08, 2.949842e-08, 3.050674e-08, 2.765042e-08, 
    2.683557e-08, 2.922227e-08, 3.091908e-08, 3.055747e-08, 2.860831e-08,
  3.141671e-08, 3.152007e-08, 3.041114e-08, 3.104346e-08, 3.264698e-08, 
    3.23984e-08, 3.044537e-08, 2.922378e-08, 3.001611e-08, 2.643544e-08, 
    2.713106e-08, 3.002068e-08, 3.054999e-08, 2.989106e-08, 2.865579e-08,
  3.113984e-08, 3.135946e-08, 3.02813e-08, 3.138966e-08, 3.255319e-08, 
    3.222249e-08, 3.030203e-08, 2.904165e-08, 2.872632e-08, 2.624171e-08, 
    2.762491e-08, 2.945342e-08, 2.971914e-08, 2.896297e-08, 2.843803e-08,
  3.121126e-08, 3.115654e-08, 3.043881e-08, 3.202377e-08, 3.332922e-08, 
    3.207127e-08, 2.974199e-08, 2.857452e-08, 2.86197e-08, 2.649266e-08, 
    2.728857e-08, 2.843484e-08, 2.840415e-08, 2.741065e-08, 2.731272e-08,
  3.095983e-08, 3.104789e-08, 3.018619e-08, 3.231673e-08, 3.333309e-08, 
    3.17234e-08, 2.92133e-08, 2.791573e-08, 2.716387e-08, 2.546037e-08, 
    2.631912e-08, 2.692123e-08, 2.700218e-08, 2.647393e-08, 2.646105e-08,
  3.097438e-08, 3.103425e-08, 3.003163e-08, 3.269289e-08, 3.402467e-08, 
    3.204391e-08, 2.83732e-08, 2.722337e-08, 2.635307e-08, 2.459948e-08, 
    2.594676e-08, 2.565047e-08, 2.537984e-08, 2.489281e-08, 2.511201e-08,
  3.172492e-08, 3.208314e-08, 3.416216e-08, 3.2454e-08, 2.98018e-08, 
    2.695259e-08, 2.577384e-08, 2.540986e-08, 2.362589e-08, 2.300162e-08, 
    2.525755e-08, 2.87839e-08, 3.357216e-08, 3.247877e-08, 3.120024e-08,
  3.122418e-08, 3.258831e-08, 3.266971e-08, 3.427461e-08, 3.316395e-08, 
    3.244879e-08, 2.802643e-08, 2.604298e-08, 2.540641e-08, 2.467396e-08, 
    2.56945e-08, 2.847692e-08, 3.291224e-08, 3.218722e-08, 2.979106e-08,
  3.045396e-08, 3.177475e-08, 3.216456e-08, 3.333952e-08, 3.35275e-08, 
    3.197762e-08, 3.437034e-08, 2.861959e-08, 2.536404e-08, 2.402724e-08, 
    2.440816e-08, 2.783547e-08, 3.17949e-08, 3.079365e-08, 2.851219e-08,
  3.081691e-08, 3.078838e-08, 3.112739e-08, 3.234366e-08, 3.361244e-08, 
    3.368406e-08, 3.26845e-08, 3.507207e-08, 3.272749e-08, 2.761e-08, 
    2.583435e-08, 2.772243e-08, 3.141513e-08, 2.909223e-08, 2.689332e-08,
  2.954638e-08, 3.039905e-08, 3.108896e-08, 3.150951e-08, 3.296308e-08, 
    3.310681e-08, 3.238188e-08, 3.095088e-08, 3.104497e-08, 2.860947e-08, 
    2.613749e-08, 2.741042e-08, 3.086346e-08, 2.820103e-08, 2.677404e-08,
  2.277983e-08, 2.609083e-08, 2.957965e-08, 3.046156e-08, 3.235762e-08, 
    3.263708e-08, 3.301678e-08, 3.144282e-08, 3.123947e-08, 2.984698e-08, 
    2.768225e-08, 2.747237e-08, 3.062264e-08, 2.704816e-08, 2.704323e-08,
  2.33478e-08, 2.579298e-08, 2.827699e-08, 2.947629e-08, 3.075474e-08, 
    3.197222e-08, 3.315599e-08, 3.086803e-08, 3.143941e-08, 3.08994e-08, 
    2.799023e-08, 2.737564e-08, 3.046196e-08, 2.619856e-08, 2.69399e-08,
  3.044716e-08, 3.069202e-08, 3.04033e-08, 3.008966e-08, 3.066606e-08, 
    3.143053e-08, 3.279323e-08, 3.142932e-08, 3.159311e-08, 3.052264e-08, 
    2.875889e-08, 2.80313e-08, 3.045882e-08, 2.598844e-08, 2.644915e-08,
  3.061523e-08, 3.071894e-08, 3.098281e-08, 3.03408e-08, 3.055305e-08, 
    3.132003e-08, 3.227796e-08, 3.132289e-08, 3.156877e-08, 3.047746e-08, 
    2.899145e-08, 2.860788e-08, 3.041562e-08, 2.560631e-08, 2.536518e-08,
  3.063601e-08, 3.094008e-08, 3.06408e-08, 3.06616e-08, 3.055077e-08, 
    3.135827e-08, 3.202903e-08, 3.185582e-08, 3.21167e-08, 3.122158e-08, 
    3.080973e-08, 2.961576e-08, 3.059013e-08, 2.567941e-08, 2.511149e-08,
  3.31734e-08, 3.233372e-08, 3.136161e-08, 2.851325e-08, 2.854491e-08, 
    2.812425e-08, 2.748611e-08, 2.758276e-08, 2.629986e-08, 2.683974e-08, 
    2.802558e-08, 2.894499e-08, 2.886553e-08, 2.817537e-08, 3.048904e-08,
  3.308382e-08, 3.34219e-08, 3.241924e-08, 3.309695e-08, 2.945143e-08, 
    3.056915e-08, 2.88687e-08, 2.769955e-08, 2.730924e-08, 2.633129e-08, 
    2.844827e-08, 2.890365e-08, 2.890498e-08, 2.818764e-08, 3.06561e-08,
  3.214578e-08, 3.274215e-08, 3.261547e-08, 3.291936e-08, 3.297324e-08, 
    3.062164e-08, 3.254531e-08, 3.036329e-08, 2.747343e-08, 2.5383e-08, 
    2.68044e-08, 2.897643e-08, 2.946621e-08, 2.839165e-08, 2.980644e-08,
  3.190482e-08, 3.221191e-08, 3.242829e-08, 3.291185e-08, 3.335098e-08, 
    3.272002e-08, 3.118497e-08, 3.503368e-08, 3.406588e-08, 2.845638e-08, 
    2.613856e-08, 2.852692e-08, 2.976375e-08, 2.919404e-08, 2.951405e-08,
  3.292329e-08, 3.286612e-08, 3.286935e-08, 3.220992e-08, 3.259707e-08, 
    3.200604e-08, 3.097149e-08, 3.103442e-08, 3.371425e-08, 3.068446e-08, 
    2.660634e-08, 2.724876e-08, 2.926994e-08, 2.958331e-08, 2.964259e-08,
  2.617838e-08, 2.686951e-08, 3.006336e-08, 3.160108e-08, 3.266506e-08, 
    3.348621e-08, 3.24924e-08, 3.091389e-08, 3.214315e-08, 3.286346e-08, 
    2.76773e-08, 2.736427e-08, 2.863255e-08, 2.96291e-08, 3.002909e-08,
  2.762113e-08, 2.558193e-08, 2.43456e-08, 2.500679e-08, 2.704185e-08, 
    3.111119e-08, 3.349672e-08, 3.220135e-08, 3.130055e-08, 3.308852e-08, 
    3.042387e-08, 2.770399e-08, 2.799036e-08, 2.911036e-08, 3.061819e-08,
  3.159075e-08, 3.150862e-08, 2.966648e-08, 2.721973e-08, 2.611992e-08, 
    2.636694e-08, 3.11158e-08, 3.249709e-08, 3.16973e-08, 3.22694e-08, 
    3.102544e-08, 2.853842e-08, 2.839361e-08, 2.772418e-08, 3.069583e-08,
  3.272838e-08, 3.095147e-08, 3.089473e-08, 3.048938e-08, 2.874911e-08, 
    2.697834e-08, 2.756011e-08, 3.133449e-08, 3.158438e-08, 3.243635e-08, 
    3.167294e-08, 2.948835e-08, 2.882532e-08, 2.707253e-08, 3.012186e-08,
  3.342907e-08, 3.291683e-08, 3.201913e-08, 3.101839e-08, 3.098218e-08, 
    2.94575e-08, 2.826967e-08, 2.940215e-08, 3.13526e-08, 3.195494e-08, 
    3.190062e-08, 3.002067e-08, 2.984517e-08, 2.680757e-08, 2.876421e-08 ;

 scalar_axis = 0 ;


 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

}
