netcdf \00010101.atmos_daily.tile3.sfcWind {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float sfcWind(time, grid_yt, grid_xt) ;
		sfcWind:_FillValue = 1.e+20f ;
		sfcWind:missing_value = 1.e+20f ;
		sfcWind:units = "m s-1" ;
		sfcWind:long_name = "Near-Surface Wind Speed" ;
		sfcWind:cell_methods = "time: mean" ;
		sfcWind:cell_measures = "area: area" ;
		sfcWind:coordinates = "height10m" ;
		sfcWind:time_avg_info = "average_T1,average_T2,average_DT" ;
		sfcWind:standard_name = "wind_speed" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 sfcWind =
  2.676566, 2.237342, 5.129944, 7.198593, 6.214886, 5.142076, 5.013721, 
    5.342939, 6.598415, 5.693856, 5.622478, 6.245234, 5.875058, 4.904199, 
    3.53325,
  4.973601, 3.771099, 2.270533, 4.682699, 4.716466, 3.74073, 3.092965, 
    2.75934, 4.598237, 6.578317, 6.022286, 7.330775, 8.256284, 5.240748, 
    3.802712,
  3.855431, 4.546868, 4.164764, 4.210362, 5.43315, 3.403949, 2.89205, 
    2.496255, 3.092183, 5.056227, 5.617712, 6.300957, 7.660041, 7.941545, 
    6.479714,
  4.966655, 3.692921, 4.051068, 4.372036, 5.392989, 5.326138, 3.071459, 
    3.252526, 3.983122, 3.772166, 3.66767, 4.688342, 6.245932, 7.456203, 
    7.870568,
  6.941166, 5.303833, 4.264295, 4.282642, 4.536706, 5.419481, 5.606862, 
    3.205959, 3.065808, 2.628367, 2.589093, 3.915194, 5.625845, 7.472782, 
    8.621073,
  6.914999, 6.719146, 5.562489, 5.138032, 4.985198, 5.011254, 4.617621, 
    5.058997, 4.676475, 3.63218, 3.231067, 4.280926, 5.34482, 6.706551, 
    7.588317,
  9.013399, 7.674922, 7.054093, 6.491871, 6.205678, 6.325101, 6.473647, 
    6.381407, 5.742992, 5.384028, 5.266144, 5.39699, 5.844362, 6.443192, 
    6.876163,
  9.911755, 8.970157, 7.891126, 7.512885, 7.266252, 7.245043, 7.303005, 
    7.178771, 6.706326, 6.703771, 6.623506, 6.165756, 5.999803, 6.194599, 
    6.206333,
  9.474393, 8.770818, 8.020311, 7.724492, 7.492144, 7.401909, 7.316968, 
    7.447396, 7.518128, 7.371616, 7.084847, 6.765952, 6.731335, 6.728504, 
    6.175414,
  8.760885, 8.395451, 7.938554, 7.524782, 7.155605, 6.99757, 7.205554, 
    7.41612, 6.877507, 5.53698, 5.705801, 6.498296, 6.262331, 5.886835, 
    5.061543,
  2.257151, 5.220962, 2.838068, 5.205431, 7.995394, 8.675356, 12.3755, 
    12.16394, 9.63312, 6.776289, 7.7875, 10.9948, 11.65955, 11.14645, 9.620898,
  6.575763, 3.195955, 3.783875, 4.753549, 5.461802, 6.3886, 11.69327, 
    12.63624, 11.23887, 9.071395, 8.776546, 12.63033, 15.14775, 10.10787, 
    9.168555,
  9.825434, 8.260166, 5.910193, 6.02725, 5.475399, 4.058213, 8.986619, 
    11.64125, 12.21465, 10.91617, 10.77696, 12.52533, 14.3524, 14.37023, 
    11.27739,
  9.613156, 9.986547, 9.359886, 7.890607, 6.406147, 5.643474, 4.02662, 
    8.926245, 12.59436, 11.11136, 10.61069, 11.91677, 13.18163, 13.46354, 
    11.86341,
  8.719664, 9.149869, 8.963287, 8.571285, 7.586767, 7.009469, 6.3846, 
    4.072005, 6.221241, 7.142079, 9.444481, 11.08412, 12.78644, 13.3361, 
    12.57618,
  8.102984, 8.586874, 8.554405, 8.527715, 8.346902, 8.044715, 7.519625, 
    7.674266, 6.548102, 6.508625, 7.037171, 10.19614, 11.75675, 12.38341, 
    11.58002,
  7.718087, 8.182459, 8.219266, 8.237362, 8.095512, 8.13272, 8.097324, 
    7.947407, 7.666409, 8.414713, 9.074242, 9.720152, 10.88356, 11.79967, 
    11.81977,
  7.406002, 7.906741, 8.040468, 8.198955, 7.919717, 7.556585, 7.210545, 
    7.276116, 7.86842, 8.847655, 9.213075, 9.113804, 9.718444, 10.59703, 
    10.84272,
  7.047329, 7.428276, 7.635486, 7.996443, 8.128611, 8.19648, 8.190429, 
    8.373331, 8.649445, 8.615705, 8.546315, 8.317041, 8.571449, 9.340138, 
    9.252439,
  6.512143, 7.03782, 7.28215, 7.445424, 7.638267, 8.044954, 8.534299, 
    8.747893, 7.853069, 6.394479, 6.732209, 7.410385, 7.223111, 7.695226, 
    7.827901,
  5.2674, 6.090342, 4.273342, 4.695629, 5.963855, 6.601816, 9.700163, 
    8.839339, 4.408764, 4.888645, 7.647266, 9.11939, 7.477998, 6.660182, 
    5.65778,
  7.376053, 7.084338, 6.645313, 5.6377, 4.264649, 4.704199, 7.366572, 
    6.447047, 3.591378, 7.363238, 8.841674, 11.42346, 12.37407, 6.711712, 
    5.602903,
  7.002623, 7.223259, 7.447055, 7.105412, 5.579566, 2.889048, 4.97482, 
    4.887989, 5.290305, 9.661407, 11.16408, 12.30538, 12.62315, 12.27331, 
    8.131632,
  6.779916, 7.027283, 7.68712, 8.320389, 8.39426, 5.063607, 2.30301, 4.77946, 
    7.664616, 9.082118, 11.29782, 12.74012, 12.96855, 12.42451, 10.32566,
  7.003661, 7.18357, 7.739654, 8.730014, 9.6057, 8.085889, 5.086749, 
    3.858768, 4.708672, 6.181781, 10.56187, 12.95168, 13.85486, 13.73399, 
    11.98227,
  7.190763, 7.525041, 7.971897, 8.841977, 9.917504, 9.57567, 7.988483, 
    8.191723, 7.275955, 7.621949, 8.440189, 12.91563, 13.96324, 13.85624, 
    12.28858,
  7.590819, 8.147516, 8.477576, 9.163658, 9.901878, 9.979602, 9.673445, 
    9.855131, 10.36388, 11.52177, 12.55323, 13.404, 14.15667, 14.21286, 
    13.99304,
  7.690682, 8.564265, 9.11147, 9.726278, 10.06819, 10.18854, 10.45117, 11.34, 
    12.16793, 13.05649, 13.66135, 13.88352, 14.39873, 15.1386, 15.81145,
  7.743967, 8.592483, 9.317517, 10.08936, 10.42586, 10.41197, 10.68605, 
    11.79595, 12.81554, 13.49295, 14.13357, 14.40852, 15.1885, 16.49484, 
    15.8692,
  7.814574, 8.838723, 9.433667, 10.10335, 10.7061, 10.80058, 10.87085, 
    11.531, 11.3141, 9.841432, 11.23683, 14.59071, 15.215, 15.92125, 14.18395,
  6.447871, 7.524941, 5.377026, 5.605843, 3.546718, 4.462369, 8.367403, 
    9.377589, 8.617589, 5.697855, 5.959538, 8.122555, 6.950385, 5.233516, 
    3.040021,
  7.524348, 5.896281, 4.61349, 3.876809, 2.26205, 2.81425, 5.574991, 
    8.084692, 8.62747, 8.144123, 7.985967, 10.98124, 11.21346, 5.011013, 
    3.149437,
  6.077006, 4.283867, 3.865932, 3.927748, 3.240459, 2.807011, 4.499547, 
    7.008015, 9.320097, 10.77663, 11.45693, 12.13805, 11.06287, 8.004298, 
    4.837331,
  4.338677, 3.42979, 4.02746, 4.361959, 4.085223, 3.814719, 4.605927, 
    6.672979, 9.320237, 10.54159, 11.94661, 12.12127, 10.63051, 7.872997, 
    5.833707,
  3.107805, 3.288079, 4.085297, 4.329671, 3.96828, 4.846987, 9.073192, 
    6.597667, 6.34355, 7.193169, 11.26338, 11.68129, 10.17512, 8.067396, 
    6.273265,
  2.924794, 3.588563, 4.257727, 4.096549, 3.301427, 5.112312, 10.82116, 
    11.65729, 9.809886, 9.038532, 8.636379, 11.24989, 9.57517, 7.713228, 
    7.299282,
  3.108172, 3.866643, 4.332938, 3.621466, 2.941133, 6.060406, 10.66759, 
    11.48594, 12.27331, 12.94169, 12.5756, 11.21897, 9.468002, 8.899949, 
    10.09713,
  3.731552, 4.201309, 4.585914, 3.565553, 4.426233, 8.388972, 12.18073, 
    13.04066, 13.55182, 13.761, 13.02012, 11.20898, 10.19947, 11.06676, 
    12.36287,
  4.420626, 4.695058, 4.820432, 4.634914, 6.892412, 10.66267, 12.92259, 
    13.07367, 13.46644, 13.76475, 13.00175, 11.66208, 11.86162, 13.21751, 
    12.70554,
  4.693767, 5.056462, 5.263218, 6.935612, 9.315482, 11.67645, 13.21455, 
    13.63159, 12.586, 10.19555, 10.17276, 12.55049, 13.14847, 13.50118, 
    12.12362,
  6.325981, 8.535336, 7.156028, 8.130208, 4.946604, 3.856562, 8.939967, 
    10.14307, 8.974958, 6.010798, 5.467537, 6.258366, 4.408255, 2.792312, 
    2.056079,
  8.544291, 8.670268, 7.81982, 6.617763, 4.499989, 6.793281, 9.647645, 
    9.339651, 8.252845, 7.621101, 6.863775, 7.981449, 6.083217, 2.233597, 
    1.348033,
  7.892917, 7.673219, 6.197774, 6.376148, 8.280169, 6.66054, 7.824824, 
    8.572418, 8.987446, 9.30792, 9.303471, 8.356108, 5.227978, 2.933376, 
    2.071805,
  7.849223, 7.122646, 5.945812, 7.706151, 11.17471, 9.253628, 6.610838, 
    7.079964, 7.523088, 8.569442, 9.465666, 8.113613, 5.307953, 3.403818, 
    2.429037,
  8.026664, 7.136493, 6.356838, 7.939669, 10.44839, 11.81648, 11.78, 6.93401, 
    5.026925, 5.933441, 8.810946, 7.68448, 5.09288, 3.252682, 2.30711,
  7.995856, 7.40433, 6.731279, 7.801232, 9.22723, 11.02446, 13.07906, 
    12.26688, 9.225309, 8.261337, 6.971602, 7.685919, 4.953757, 3.11988, 
    3.113241,
  8.33755, 8.01079, 7.149076, 7.741569, 8.425085, 10.21242, 12.07219, 
    11.27063, 11.53649, 11.76125, 10.37759, 7.978199, 4.845638, 3.327373, 
    3.760747,
  9.004086, 8.522618, 7.219384, 7.366332, 8.171852, 10.60426, 12.94846, 
    12.6138, 12.71908, 12.15754, 10.71072, 7.910759, 4.674873, 3.887438, 
    4.306443,
  9.652769, 8.848811, 7.380692, 7.215401, 8.516116, 11.84339, 13.68478, 
    12.59656, 12.19985, 11.86709, 10.66808, 7.587941, 4.962209, 4.835042, 
    4.517015,
  9.903681, 8.538985, 7.028929, 7.673536, 9.786084, 12.6415, 13.79149, 
    12.84947, 11.31579, 8.714995, 7.878811, 7.371952, 5.691524, 5.308788, 
    4.424294,
  5.648944, 7.451566, 6.595611, 7.659402, 6.957153, 5.203731, 6.895168, 
    8.268055, 6.855992, 3.383074, 2.653455, 3.469206, 3.159338, 3.478807, 
    2.94666,
  7.869815, 8.445765, 8.713507, 9.067552, 6.369481, 5.176528, 7.400589, 
    7.656099, 5.889519, 4.048784, 2.698423, 3.797035, 4.388642, 2.820866, 
    1.782141,
  7.768455, 8.741469, 9.274922, 10.21344, 8.982773, 5.953169, 7.003803, 
    7.199245, 6.483496, 4.939179, 3.403181, 3.535324, 4.540225, 3.84253, 
    1.42375,
  8.141805, 9.059665, 9.545518, 10.89802, 12.88613, 10.00992, 6.201511, 
    5.616955, 4.704871, 4.431619, 3.403067, 3.140164, 4.077629, 3.665161, 
    1.837633,
  8.89572, 9.37854, 9.695147, 10.61628, 13.06314, 13.25169, 11.38473, 
    6.015388, 4.074206, 3.812463, 3.627328, 2.721015, 3.454533, 3.453539, 
    2.663993,
  9.692572, 9.641799, 9.672244, 10.3666, 12.69099, 13.40254, 12.7555, 
    11.70638, 7.921458, 6.358003, 4.037633, 2.381596, 2.592621, 3.203698, 
    3.366425,
  10.57005, 10.03754, 9.708907, 10.56092, 12.43096, 12.83623, 11.76435, 
    10.32878, 9.198935, 8.692348, 6.088489, 2.421711, 2.026601, 2.744389, 
    2.936467,
  11.02349, 10.1719, 9.70274, 10.85414, 12.54398, 12.49629, 12.07457, 11.788, 
    11.20112, 9.749838, 6.728385, 2.936096, 1.908122, 2.581881, 2.930777,
  11.27106, 10.30248, 9.952607, 11.28555, 12.69612, 12.39971, 12.10446, 
    11.68048, 10.85529, 9.645205, 7.402756, 3.751693, 2.025494, 2.305043, 
    2.577282,
  11.04034, 10.1821, 9.97564, 11.34453, 12.63061, 12.30932, 12.23036, 
    12.00477, 10.11852, 7.220146, 6.185321, 4.447738, 2.273983, 1.88907, 
    2.342562,
  4.865697, 6.946022, 6.659752, 7.505806, 6.493139, 4.50583, 3.923552, 
    3.803232, 4.072763, 3.807205, 4.5029, 3.919564, 3.122314, 3.640477, 
    3.138391,
  7.859253, 8.060833, 8.839211, 8.832809, 6.302575, 4.117329, 4.175149, 
    3.41256, 3.635052, 4.900749, 4.873224, 5.487565, 4.252197, 2.717789, 
    2.437264,
  8.577957, 8.598182, 9.484961, 10.02961, 7.932535, 4.025171, 4.044272, 
    2.976579, 2.731307, 3.933542, 5.861169, 6.042147, 4.908083, 3.722207, 
    3.336406,
  9.322439, 9.422224, 10.09943, 10.8244, 10.51439, 7.352609, 3.6781, 
    2.532501, 2.294263, 3.093576, 4.923769, 5.627968, 4.973802, 3.761924, 
    3.055209,
  10.53913, 10.4858, 10.89901, 11.47842, 10.78724, 8.982109, 7.367062, 
    3.067693, 2.53794, 2.292643, 3.247794, 5.076087, 4.816714, 4.126807, 
    2.782353,
  11.71333, 11.29907, 11.57267, 11.97376, 11.2571, 9.226321, 7.417449, 
    5.357789, 3.129664, 2.415121, 1.782175, 4.241781, 4.979162, 4.791076, 
    4.009931,
  12.67599, 12.215, 12.35065, 12.7049, 12.00957, 10.05194, 7.794874, 
    5.149667, 3.968252, 3.932776, 2.677155, 3.632612, 4.643477, 4.741834, 
    4.45203,
  12.94792, 12.73088, 12.81961, 13.19706, 12.63462, 10.64016, 8.589883, 
    7.21865, 6.432206, 5.038966, 3.09832, 2.716768, 4.277606, 4.623248, 
    4.440538,
  12.55187, 12.90599, 13.28834, 13.69524, 13.22708, 11.21588, 8.94953, 
    7.688651, 7.050154, 5.662179, 4.046185, 1.935966, 3.464253, 4.373347, 
    4.46021,
  11.93983, 12.59039, 13.1751, 13.59477, 13.2299, 11.31537, 8.767681, 
    8.029303, 7.682194, 5.419854, 4.442766, 2.194334, 2.191396, 3.465152, 
    4.08339,
  5.532729, 7.869373, 6.965435, 7.248662, 5.007086, 1.861451, 3.498797, 
    5.180386, 5.762467, 3.985022, 3.565114, 3.635799, 3.410076, 3.598775, 
    3.04056,
  8.692351, 9.978804, 10.16274, 9.027081, 5.458793, 2.150165, 2.780995, 
    4.400072, 5.292077, 5.036636, 4.095773, 4.66457, 4.93212, 3.237766, 
    2.679876,
  9.006564, 10.8081, 11.28459, 10.2476, 6.843683, 2.55808, 1.830363, 
    2.981696, 4.216638, 5.110519, 5.186659, 5.087273, 4.85446, 4.846385, 
    3.920353,
  8.646903, 10.92272, 11.78848, 10.97309, 8.614044, 5.314394, 2.336986, 
    2.855181, 3.981485, 4.298725, 4.915589, 5.190724, 5.03905, 4.786297, 
    4.252375,
  7.900221, 10.88533, 11.97751, 11.24175, 8.696708, 5.949118, 5.043592, 
    2.421004, 2.060235, 2.489384, 4.108311, 4.955101, 4.880614, 4.698464, 
    4.339772,
  7.364312, 10.7949, 11.93108, 11.19884, 9.150743, 6.488184, 4.372681, 
    2.714844, 2.729831, 3.39158, 3.609378, 4.779891, 4.608314, 4.077835, 
    3.246785,
  8.028172, 10.58799, 11.6433, 11.24037, 9.649682, 7.112318, 4.976859, 
    2.925723, 3.262817, 4.389073, 4.787179, 4.680481, 4.533529, 4.027202, 
    3.190645,
  8.864995, 10.33363, 11.26102, 11.2088, 10.19687, 8.14972, 5.688583, 
    4.055049, 4.133268, 4.792703, 4.890965, 4.729079, 4.714757, 4.41777, 
    3.769854,
  9.207134, 10.243, 11.18481, 11.36409, 10.726, 9.207776, 7.137011, 4.92128, 
    4.538311, 5.034261, 4.75001, 4.655538, 4.961062, 4.881531, 4.16797,
  11.30646, 11.12191, 11.21317, 11.45155, 11.10684, 9.853225, 8.191512, 
    6.33043, 5.333071, 4.657636, 4.402446, 4.652347, 5.018022, 4.986595, 
    4.335745,
  4.706368, 8.607952, 8.798394, 10.00335, 7.598094, 5.279632, 6.941613, 
    6.780446, 5.610685, 3.636719, 3.487492, 3.297128, 3.714339, 4.293313, 
    3.737277,
  5.393965, 9.687178, 11.89757, 11.49464, 6.851958, 4.507771, 6.845479, 
    6.841622, 5.465273, 4.201134, 2.976569, 3.255254, 3.641246, 3.098551, 
    3.00237,
  4.38359, 9.442265, 12.49169, 12.16739, 8.50324, 4.267771, 5.856414, 
    6.503351, 6.164331, 4.744919, 3.579711, 2.960504, 2.957498, 3.192905, 
    2.583782,
  4.580482, 9.290597, 12.56672, 12.31447, 10.71015, 7.545235, 4.362595, 
    4.606547, 4.2617, 4.484294, 3.758394, 2.784984, 2.521631, 2.631073, 
    2.478955,
  5.020181, 9.36693, 12.40666, 11.90942, 10.11958, 9.14231, 8.503239, 
    4.519539, 3.605686, 3.90701, 4.745904, 3.436862, 2.561419, 2.439025, 
    2.74065,
  5.16722, 9.50814, 12.04795, 11.34085, 9.588134, 8.449897, 8.604783, 
    8.472171, 6.05292, 5.275027, 5.041353, 4.552317, 2.930045, 2.525478, 
    2.683289,
  5.806234, 9.719622, 11.59535, 10.67478, 8.810568, 7.547213, 7.140622, 
    6.324478, 5.939044, 7.113808, 7.010445, 5.213098, 3.277083, 2.29127, 
    1.90135,
  5.72582, 9.446876, 10.81135, 9.930005, 8.276264, 7.074458, 6.523122, 
    6.374712, 6.916414, 7.601491, 7.005937, 5.618233, 3.745972, 2.358782, 
    2.072212,
  5.371377, 8.806076, 10.15647, 9.318643, 7.784125, 6.807949, 6.043951, 
    5.317929, 5.843452, 6.940423, 7.041921, 5.992015, 4.473422, 3.438213, 
    3.073272,
  6.160585, 7.876328, 9.300264, 8.953384, 7.664724, 6.621761, 6.029016, 
    5.416363, 5.647261, 5.387189, 5.987144, 6.207534, 5.140503, 4.49659, 
    3.948613,
  5.901932, 8.184597, 6.70495, 6.817003, 5.85981, 4.29058, 5.23857, 5.53484, 
    6.083797, 4.484345, 4.752928, 5.067269, 4.0532, 3.829602, 3.35907,
  9.213236, 9.503554, 9.356365, 8.175788, 5.426669, 3.788155, 4.943905, 
    5.219836, 5.590844, 5.775627, 5.097376, 6.60453, 6.779786, 3.848913, 
    3.394642,
  9.045356, 9.46045, 9.669355, 8.647976, 6.430966, 3.013605, 3.846889, 
    3.847132, 3.905388, 4.917331, 6.233069, 6.93413, 7.218227, 6.908862, 
    4.653176,
  8.799802, 9.466289, 9.605604, 8.509484, 7.296633, 5.226601, 2.38944, 
    3.387752, 3.913159, 3.81198, 4.935904, 6.198584, 6.754334, 6.932894, 
    5.694706,
  9.001707, 9.387442, 9.370314, 8.295838, 6.885045, 5.628635, 4.645867, 
    2.149518, 3.062454, 2.701612, 3.019207, 4.983314, 6.1453, 6.561931, 
    6.907558,
  8.876091, 9.236551, 9.239599, 8.231499, 7.206998, 5.910779, 4.709842, 
    3.716892, 2.430038, 1.905288, 2.328661, 3.699276, 5.232233, 6.177033, 
    7.15176,
  8.075912, 8.943159, 9.204719, 8.438302, 7.404428, 6.294295, 5.105021, 
    3.602925, 2.508403, 2.794819, 2.912813, 3.009692, 4.118124, 5.602052, 
    7.251866,
  7.109616, 8.495394, 9.023877, 8.506646, 7.710736, 6.942384, 6.150697, 
    4.70458, 3.534071, 3.47896, 3.379005, 2.81764, 3.377841, 4.836395, 
    6.278863,
  6.588718, 8.276615, 9.152003, 8.673676, 7.828351, 7.073381, 6.441782, 
    5.631338, 4.440187, 4.445053, 4.876651, 3.60818, 3.121245, 4.086595, 
    4.972872,
  7.456804, 8.054016, 8.939194, 8.805348, 8.053878, 7.227547, 6.637617, 
    6.1798, 5.608046, 4.959473, 5.400912, 4.682501, 3.641682, 3.629661, 
    4.108955,
  4.057718, 4.371275, 2.583485, 2.475929, 3.639771, 4.135655, 5.386626, 
    5.768576, 6.612471, 4.741183, 4.480164, 4.21019, 2.950642, 2.987876, 
    2.428247,
  6.228278, 4.617505, 3.064959, 2.304882, 2.33133, 3.898491, 5.703063, 
    6.055915, 6.789916, 6.554974, 5.012808, 5.560711, 4.942787, 3.210776, 
    3.072376,
  5.919842, 4.378007, 3.093019, 2.084568, 1.782703, 2.19023, 4.689634, 
    4.91202, 5.513291, 6.878586, 6.900951, 6.269884, 6.241178, 5.913092, 
    3.993778,
  5.833354, 4.431814, 3.399728, 1.997557, 1.40587, 1.695324, 1.763151, 
    5.070348, 7.712199, 7.662927, 7.60447, 6.966374, 6.751788, 6.658394, 
    5.361024,
  6.071954, 5.111403, 4.319631, 3.075709, 1.661733, 1.445701, 1.718597, 
    2.187094, 3.515337, 4.843382, 6.473742, 7.001587, 7.270809, 7.111843, 
    7.560399,
  7.513063, 6.697297, 5.876964, 4.677046, 3.117821, 1.399025, 1.643669, 
    2.990526, 1.624298, 2.617321, 4.317072, 6.173604, 6.969302, 7.510973, 
    8.47315,
  9.668384, 9.265064, 8.387494, 7.26918, 5.637989, 3.206583, 1.463917, 
    2.285893, 2.813554, 3.355157, 4.496603, 5.564673, 6.489243, 7.075838, 
    8.42579,
  11.39547, 11.53982, 10.93149, 9.607867, 7.860511, 5.932543, 4.202165, 
    3.15324, 3.586293, 3.70659, 3.610765, 4.652383, 5.772137, 6.71996, 
    7.737216,
  12.74179, 13.27917, 13.23897, 12.03491, 9.779819, 7.459118, 5.297348, 
    4.03539, 4.656116, 4.698279, 3.003331, 3.43322, 4.623632, 6.010536, 
    6.512589,
  10.11545, 11.7453, 12.61547, 12.84353, 11.54505, 9.010182, 6.624331, 
    5.468206, 5.928007, 5.03204, 3.944818, 3.272702, 3.348186, 4.426528, 
    5.709217,
  3.185826, 3.055042, 3.471933, 2.63087, 2.034699, 3.048089, 4.567438, 
    5.192883, 5.315899, 4.059145, 4.250091, 4.739316, 3.802477, 3.624555, 
    3.229285,
  5.394598, 3.540131, 1.932818, 1.44765, 1.414552, 1.892757, 4.212577, 
    4.996297, 5.373487, 5.458049, 5.1103, 6.792465, 6.849403, 4.021681, 
    3.837011,
  5.737999, 4.479711, 2.679182, 2.177775, 2.01553, 1.583456, 2.796303, 
    4.210442, 4.726451, 5.598093, 6.516964, 7.556244, 8.372944, 8.069737, 
    6.138281,
  6.437821, 5.411855, 4.379252, 3.606569, 2.508438, 2.805431, 1.821997, 
    3.815066, 5.464559, 5.756902, 6.345576, 7.372863, 8.594738, 9.102748, 
    8.004222,
  8.106486, 7.105046, 6.180076, 4.860508, 2.989393, 1.734942, 4.675584, 
    2.247838, 2.707774, 3.884666, 5.173265, 6.78941, 8.206013, 9.280378, 
    10.17847,
  10.83737, 9.498386, 8.259811, 6.471676, 4.735497, 2.520827, 3.651876, 
    4.102962, 1.059525, 2.204585, 3.622113, 5.758455, 7.519471, 9.036531, 
    10.81539,
  13.65419, 12.30894, 10.41555, 8.271766, 6.330012, 4.755146, 5.049638, 
    4.533054, 1.990492, 1.799071, 2.824561, 4.5877, 6.635709, 8.319914, 
    10.41706,
  11.21804, 13.10268, 13.07813, 11.36737, 9.074532, 7.144638, 7.012515, 
    7.083934, 4.88706, 2.432069, 1.915253, 3.251232, 5.392658, 7.328416, 
    9.565567,
  4.60875, 5.104574, 8.724586, 11.55767, 11.74736, 9.918619, 8.464067, 
    8.039197, 7.270212, 5.148034, 3.022098, 1.92587, 3.554624, 5.947112, 
    8.429029,
  5.540038, 4.502351, 3.325431, 5.258508, 9.687979, 11.10509, 9.941257, 
    8.68248, 7.785678, 5.764583, 4.813913, 2.726784, 1.816953, 4.148333, 
    7.104447,
  4.132129, 4.190121, 4.445381, 5.242248, 3.410038, 1.618947, 2.467774, 
    4.130494, 5.46928, 4.89977, 5.705835, 7.154598, 5.961607, 5.341382, 
    4.002805,
  7.236729, 4.574401, 2.974372, 2.521932, 3.092771, 1.774487, 2.069048, 
    3.413501, 4.889832, 6.028249, 6.836507, 9.555165, 9.542266, 5.07928, 
    4.593153,
  8.347221, 5.767514, 3.693038, 4.104083, 1.997216, 2.385365, 1.844831, 
    1.975224, 2.582121, 4.97908, 7.798064, 10.23283, 10.93173, 9.661461, 
    6.603491,
  8.720086, 7.366376, 5.184095, 4.739166, 2.774497, 3.692121, 1.55974, 
    2.319139, 4.30456, 5.328059, 6.905702, 9.183935, 10.95638, 11.06059, 
    8.624543,
  9.067961, 8.179012, 6.997211, 5.602832, 4.630503, 2.805287, 5.121317, 
    2.067151, 2.924722, 4.100009, 5.620687, 7.650841, 9.727874, 11.00855, 
    10.79067,
  10.6328, 9.281037, 8.231966, 6.70366, 5.562225, 3.164154, 4.393656, 
    5.007274, 3.440015, 2.901199, 3.905541, 6.046314, 8.158278, 9.975264, 
    11.03907,
  12.26688, 10.59166, 9.171172, 7.771753, 6.599313, 4.765627, 4.72074, 
    4.743708, 4.209733, 3.566037, 4.142251, 4.85421, 6.230748, 8.182841, 
    10.17257,
  12.17749, 11.4874, 10.45289, 9.425303, 8.519662, 7.1299, 6.562028, 
    6.745748, 6.642476, 5.960617, 5.242468, 4.383014, 4.525999, 5.877561, 
    8.096663,
  8.811747, 10.01343, 10.56852, 10.50257, 10.17618, 9.205239, 8.513628, 
    8.463898, 8.297946, 7.074645, 6.335875, 5.377788, 4.010439, 4.185956, 
    5.822001,
  5.614242, 6.755966, 8.06176, 8.928264, 9.627161, 9.617815, 9.465493, 
    9.229988, 8.074474, 5.927775, 6.33911, 7.293045, 5.763407, 4.377142, 
    3.999093,
  8.790821, 10.87337, 8.46753, 8.785545, 6.555889, 3.54414, 2.79087, 
    2.143156, 2.559009, 2.936082, 4.382288, 5.513359, 4.911601, 4.525085, 
    2.934867,
  12.28042, 11.11881, 10.16081, 8.855936, 4.731696, 1.740695, 2.071971, 
    2.324667, 3.472674, 3.847155, 4.50854, 6.382427, 6.880147, 4.29682, 
    3.539824,
  11.5064, 9.930027, 9.541972, 8.758312, 5.654658, 2.094641, 1.045757, 
    1.436186, 2.324188, 3.020412, 4.573555, 6.315518, 7.81246, 7.228889, 
    4.996949,
  10.33953, 8.739219, 8.396926, 7.843716, 6.390952, 4.623681, 1.753466, 
    1.895514, 3.333144, 3.056047, 3.977402, 5.842175, 7.632548, 7.73905, 
    6.041926,
  9.61808, 8.353555, 7.229459, 6.034119, 4.830643, 3.825262, 4.848138, 
    2.309733, 2.964124, 3.397388, 3.753645, 5.898321, 7.228621, 7.136908, 
    6.475379,
  9.157559, 8.37231, 7.231927, 5.838188, 4.61514, 3.576902, 4.036478, 
    4.589216, 3.992766, 3.78842, 4.012321, 6.477111, 7.250192, 6.302297, 
    5.4636,
  9.003205, 8.432755, 7.584352, 6.570775, 5.79601, 5.36318, 5.40706, 
    5.422512, 4.715438, 5.854287, 6.815829, 7.634896, 7.137312, 5.3649, 
    4.19745,
  9.252961, 8.697984, 8.199452, 7.631521, 7.456653, 7.466616, 7.685243, 
    7.623724, 7.432156, 6.981265, 7.907895, 7.823179, 6.482633, 4.563443, 
    3.507407,
  9.589992, 9.230744, 9.193387, 9.134091, 9.252168, 9.344498, 9.422462, 
    9.379038, 9.11223, 7.048235, 7.185032, 7.045774, 6.237112, 4.996377, 
    3.920979,
  9.955256, 9.843093, 9.929488, 10.12981, 10.40565, 10.63203, 10.7732, 
    10.45473, 8.285835, 5.697019, 6.571977, 8.016209, 7.074212, 6.35814, 
    5.282373,
  6.600402, 10.54861, 9.614014, 11.27806, 9.895319, 6.053406, 5.60976, 
    3.416738, 1.239037, 2.302795, 4.047443, 5.57227, 5.828889, 5.388053, 
    3.453009,
  10.25315, 12.41531, 13.29077, 12.61887, 7.921637, 4.503846, 4.859607, 
    2.786997, 2.440202, 4.134914, 4.760657, 6.778001, 7.864617, 4.61875, 
    3.090457,
  10.65678, 12.71357, 13.91716, 13.07893, 8.988732, 4.248497, 3.151658, 
    2.580873, 3.546522, 4.48299, 5.288293, 7.269625, 8.072322, 6.327062, 
    3.597196,
  10.72483, 12.59216, 13.63029, 12.7891, 11.02571, 7.111084, 2.670691, 
    1.308923, 2.363042, 2.057381, 4.402522, 6.980067, 7.753511, 5.378855, 
    3.608131,
  10.91134, 12.3572, 12.93251, 11.96897, 10.17422, 8.414868, 6.38381, 
    2.437881, 1.570135, 2.528992, 4.353723, 6.4067, 7.159794, 4.267031, 
    3.116444,
  10.99601, 11.92786, 12.16169, 11.1583, 9.852296, 8.293519, 7.125976, 
    5.185888, 3.034508, 3.780077, 3.916987, 5.769063, 6.433319, 4.17279, 
    2.136413,
  10.87025, 11.34649, 11.23286, 10.31251, 9.107751, 7.947078, 6.822543, 
    5.811627, 5.084004, 5.273932, 5.195084, 5.604811, 5.717566, 4.48113, 
    1.660885,
  10.28854, 10.4046, 10.00429, 9.152997, 8.284471, 7.46148, 6.952074, 
    6.623979, 6.408046, 5.483312, 5.52109, 5.420407, 5.346097, 4.662166, 
    1.969588,
  9.276164, 9.180963, 8.823153, 8.173213, 7.593825, 7.300504, 7.351593, 
    7.546215, 7.555023, 5.931969, 5.976445, 6.218277, 5.945007, 5.247193, 
    3.174367,
  7.804911, 7.570743, 7.384935, 7.308066, 7.412013, 7.714617, 8.177129, 
    8.451207, 7.099526, 5.002565, 6.039537, 7.670609, 7.142905, 6.473494, 
    5.11342,
  7.779065, 10.28309, 8.312889, 9.222607, 7.619728, 4.541872, 3.736452, 
    2.162892, 3.583177, 3.825232, 2.868859, 3.356904, 3.5267, 3.150054, 
    2.902898,
  12.2899, 12.23329, 11.41615, 10.28042, 6.139679, 3.602959, 3.353292, 
    1.81876, 3.885079, 5.13553, 4.070677, 3.441026, 4.651532, 3.175937, 
    2.862447,
  12.39379, 12.13965, 11.75815, 10.94002, 7.634396, 3.815625, 2.360785, 
    1.224043, 3.278378, 4.558833, 5.292083, 4.615663, 4.196691, 5.097429, 
    4.138512,
  11.78435, 11.49554, 11.32784, 11.05305, 10.22526, 6.982447, 2.836514, 
    1.493469, 2.283121, 3.139354, 4.644488, 5.715745, 4.725369, 5.17896, 
    4.868449,
  10.66312, 10.67112, 10.6809, 10.61881, 10.05158, 9.013443, 7.230655, 
    3.287742, 1.749566, 2.032218, 4.130989, 5.333416, 6.280163, 5.36647, 
    6.058136,
  9.701818, 10.09103, 10.26375, 10.30695, 10.13969, 9.365982, 8.448495, 
    6.895845, 3.541111, 2.189843, 3.199386, 4.779752, 6.064791, 5.506523, 
    6.188756,
  8.898491, 9.635915, 10.12279, 10.08555, 9.985076, 9.447248, 8.493336, 
    7.246181, 5.44777, 3.483685, 3.763382, 4.721004, 5.656883, 6.149603, 
    6.314033,
  7.980174, 8.985055, 9.796532, 9.902767, 9.893684, 9.6695, 9.039845, 8.3488, 
    7.315285, 5.038881, 4.236465, 4.599754, 5.51258, 6.243146, 6.028043,
  6.993393, 8.092615, 9.034041, 9.317954, 9.383353, 9.392653, 9.080052, 
    8.485266, 7.640584, 6.207294, 4.955919, 5.032342, 5.786574, 6.02323, 
    5.479634,
  5.520275, 6.512891, 7.290069, 7.694093, 8.040358, 8.284212, 8.358141, 
    8.083543, 6.943491, 4.755005, 5.18048, 5.648964, 5.739019, 5.9289, 
    5.294306,
  6.208655, 7.860638, 6.183523, 6.169946, 4.426025, 2.446849, 2.639277, 
    4.700215, 5.861772, 4.878762, 5.271228, 7.393245, 6.601018, 5.119331, 
    4.304044,
  9.865131, 9.415935, 8.619508, 7.147533, 3.93151, 1.526987, 1.788892, 
    3.801583, 5.694224, 5.957235, 5.967283, 9.262547, 9.981906, 5.22755, 
    3.367647,
  10.48023, 9.703243, 9.081619, 8.147436, 5.809135, 2.486163, 2.603033, 
    2.995728, 3.90908, 4.892782, 6.314673, 9.486029, 10.89107, 8.631336, 
    4.973754,
  10.69067, 9.884067, 9.260694, 8.520702, 7.9258, 5.899059, 2.390339, 
    2.928794, 4.307277, 4.220223, 4.992903, 8.241857, 10.38847, 9.385479, 
    6.088859,
  10.65756, 10.11478, 9.39032, 8.552647, 8.003577, 7.494781, 6.528172, 
    2.815077, 3.521907, 3.54797, 3.869617, 6.502421, 9.421911, 9.520658, 
    7.258307,
  10.12363, 10.11917, 9.403863, 8.693191, 8.341862, 8.076038, 8.114335, 
    7.539656, 5.486383, 3.608963, 2.646888, 4.944909, 8.195824, 8.918081, 
    7.747339,
  9.269541, 9.579055, 9.235055, 8.709579, 8.429191, 8.170969, 8.04326, 
    7.688241, 6.800319, 4.917179, 3.265575, 3.282548, 6.492876, 8.161367, 
    7.646123,
  8.511911, 8.787011, 8.793075, 8.638118, 8.513451, 8.222715, 7.930278, 
    7.395638, 6.781555, 5.766769, 4.886623, 3.087098, 4.474138, 6.565992, 
    6.924812,
  7.259303, 8.052204, 8.611817, 8.955153, 9.169142, 9.001657, 8.577769, 
    7.935912, 7.023608, 6.189635, 5.957713, 4.475176, 3.067577, 4.531682, 
    5.858045,
  3.855883, 4.996433, 6.162229, 7.064224, 7.714062, 7.922819, 7.865478, 
    7.56415, 6.338286, 4.79563, 5.92213, 6.060116, 3.799678, 3.045186, 
    4.270118,
  5.538321, 6.928534, 5.165935, 4.636313, 3.589536, 3.308949, 3.905955, 
    4.328326, 4.690073, 4.07587, 4.135221, 4.517647, 4.133694, 4.129585, 
    3.565378,
  8.694207, 7.691854, 6.034854, 3.427622, 1.794847, 3.520948, 4.731143, 
    4.703241, 4.700067, 4.500423, 4.262011, 5.11848, 5.078627, 3.102984, 
    2.628716,
  8.221943, 6.661803, 4.823211, 3.169821, 2.556093, 2.565756, 4.52587, 
    4.423487, 3.143924, 4.058448, 4.660714, 5.201233, 5.002546, 4.277793, 
    3.129071,
  7.231881, 5.590473, 4.308237, 3.800709, 4.172708, 4.120535, 3.147422, 
    3.954995, 3.147432, 3.835295, 4.576429, 5.096415, 5.170827, 4.116301, 
    3.174313,
  7.031541, 5.645036, 4.912419, 4.921131, 5.735627, 6.292629, 5.842523, 
    3.105677, 2.750785, 3.052114, 4.561458, 5.04932, 5.53528, 4.384102, 
    2.941453,
  6.977317, 6.516152, 6.371337, 6.623405, 7.291189, 7.601111, 7.012694, 
    5.882077, 3.720795, 3.406317, 3.903628, 4.755113, 5.844177, 5.00506, 
    3.053619,
  7.571508, 7.652897, 7.959709, 8.255311, 8.490312, 7.946927, 6.596362, 
    4.847347, 2.736068, 4.507984, 6.181194, 4.45472, 6.058308, 5.877079, 
    4.02465,
  8.804162, 8.378914, 8.41048, 8.473766, 8.265303, 7.019855, 5.232838, 
    3.736575, 2.683532, 4.288515, 6.726446, 5.042481, 5.728564, 6.514235, 
    4.923511,
  9.407605, 8.783781, 8.372358, 7.782663, 6.843114, 5.508269, 4.797223, 
    4.579159, 4.364179, 4.411908, 6.901412, 6.654984, 5.162101, 6.454079, 
    6.145304,
  7.515796, 6.328261, 5.440392, 4.669532, 4.095718, 3.837441, 3.875902, 
    4.043617, 4.05636, 3.97724, 5.931068, 8.112292, 5.994048, 5.279871, 
    6.199364,
  3.7332, 3.188526, 1.917853, 3.516217, 4.450903, 4.513604, 3.846476, 
    4.666885, 6.436342, 4.048989, 2.998586, 2.869503, 3.359715, 4.248571, 
    4.609026,
  5.846456, 3.298204, 1.77943, 3.03361, 4.148382, 4.995658, 5.6269, 3.923486, 
    6.521902, 5.794692, 3.784827, 3.451952, 3.643369, 3.541471, 4.511229,
  5.578584, 3.172982, 1.773531, 3.623852, 4.570025, 4.592739, 5.952552, 
    3.537456, 6.023265, 6.753618, 5.054025, 3.631426, 3.292591, 4.782893, 
    5.605975,
  5.404241, 3.278581, 2.852871, 4.856116, 7.266408, 6.425317, 4.372542, 
    3.216207, 3.263551, 6.761625, 5.724566, 4.014306, 3.26175, 4.670812, 
    5.573116,
  5.433076, 4.204302, 4.408788, 6.176658, 8.464708, 8.844225, 6.015908, 
    2.616592, 2.91746, 4.745517, 5.321003, 4.380907, 3.284158, 4.183375, 
    6.197893,
  5.965694, 5.686504, 5.80012, 7.05486, 8.530952, 8.57658, 6.243464, 
    3.533121, 2.25743, 3.083743, 3.817334, 4.457064, 3.497009, 3.736851, 
    5.64944,
  6.316249, 6.243423, 6.430296, 7.12244, 8.177827, 7.457987, 5.52041, 
    3.308109, 1.919146, 4.014184, 5.674351, 4.784585, 3.911544, 3.245439, 
    4.442399,
  7.984393, 7.284372, 7.122775, 7.477304, 7.889085, 6.358296, 4.445759, 
    3.064151, 2.826475, 4.507936, 6.134165, 5.389099, 4.249737, 3.016643, 
    3.379075,
  9.764737, 8.97428, 8.358998, 8.012813, 6.947641, 5.042644, 4.187864, 
    3.777682, 4.427526, 4.698042, 6.364714, 6.415745, 5.244319, 3.540995, 
    2.271768,
  10.40785, 9.566898, 8.42308, 7.227278, 5.601775, 4.879311, 4.642848, 
    4.496539, 4.442057, 4.221063, 5.815458, 7.491629, 6.839461, 4.976956, 
    2.447393,
  4.004686, 3.9972, 3.926405, 5.871718, 6.978483, 7.183959, 8.592108, 
    6.662881, 4.486709, 3.762302, 4.300552, 4.685695, 4.269891, 4.203556, 
    3.529917,
  7.432558, 5.794902, 4.989845, 5.8897, 5.396309, 6.106268, 8.134979, 
    6.92132, 5.505276, 4.849803, 4.438756, 5.074315, 4.403376, 3.489138, 
    3.278916,
  8.319006, 6.906734, 6.07531, 6.662998, 5.950323, 5.157122, 6.678599, 
    6.177904, 4.984344, 4.965694, 5.069549, 4.808229, 4.189233, 5.037021, 
    4.017788,
  8.717314, 7.672441, 7.114904, 7.361767, 8.833053, 6.741039, 4.735421, 
    5.367511, 6.31132, 5.603374, 4.514411, 4.035382, 3.934308, 5.106784, 
    3.928055,
  7.965442, 7.936872, 7.85575, 8.141917, 9.27262, 8.875995, 6.427486, 
    3.798233, 5.258554, 5.220373, 4.173136, 3.693727, 3.429929, 4.292402, 
    4.582441,
  7.251875, 7.476181, 7.864942, 8.342365, 8.772647, 8.718006, 7.947182, 
    6.049993, 5.169336, 4.438258, 3.510909, 4.13133, 2.977497, 3.197732, 
    4.098057,
  8.585588, 8.203096, 8.263187, 8.500107, 8.741938, 8.792173, 8.80838, 
    8.293805, 6.388485, 5.018813, 4.937958, 4.449498, 2.283275, 1.593873, 
    3.398224,
  10.02994, 9.565112, 9.44702, 9.375648, 9.520269, 9.516201, 9.122515, 
    8.343999, 6.675958, 5.572744, 4.776005, 4.080215, 2.147667, 1.124103, 
    2.753455,
  10.12261, 10.30658, 10.32753, 10.20971, 10.19173, 10.03105, 9.601027, 
    8.643242, 7.788082, 5.242677, 4.387582, 4.002018, 2.606608, 2.373556, 
    1.807525,
  9.240671, 9.853199, 10.2597, 10.57051, 10.8434, 10.55248, 9.591677, 
    9.296779, 6.62746, 4.02224, 4.584779, 4.041582, 2.873266, 4.081994, 
    2.100235,
  5.21099, 6.832413, 6.028667, 7.288939, 6.944037, 6.644565, 9.463963, 
    10.37342, 9.721254, 7.405952, 7.142209, 6.789349, 5.045526, 2.170166, 
    3.198397,
  9.13701, 9.640193, 9.494046, 9.713114, 5.763348, 5.774864, 9.868049, 
    10.54449, 10.31626, 8.500834, 7.108144, 7.587493, 5.663706, 2.397803, 
    4.46736,
  8.319671, 9.681117, 9.995657, 10.51609, 7.945249, 5.576315, 8.427629, 
    9.736564, 9.64211, 9.270798, 8.546647, 7.989081, 5.571936, 3.79693, 
    7.117565,
  7.023778, 8.357069, 9.371741, 10.29999, 10.90227, 8.621248, 5.733505, 
    6.61775, 8.122284, 8.564598, 8.487993, 7.955941, 5.133623, 4.219114, 
    8.631398,
  6.553926, 7.683639, 9.069385, 10.33825, 11.38407, 11.71075, 9.960735, 
    5.763523, 6.772356, 6.675237, 7.858179, 7.918599, 4.992414, 5.311128, 
    10.42083,
  6.912235, 7.971724, 9.484607, 10.90057, 12.0091, 12.83558, 13.01872, 
    12.2983, 8.912442, 7.263432, 6.78143, 8.05863, 5.00456, 5.793779, 9.951278,
  9.030939, 10.19122, 11.4454, 12.44734, 13.36172, 13.86631, 14.32468, 
    13.99535, 12.91015, 10.66728, 9.561544, 8.33426, 5.262682, 7.68783, 
    10.92901,
  10.98353, 11.92223, 12.73871, 13.09886, 13.82556, 14.12327, 13.55818, 
    12.86476, 11.92045, 10.00703, 9.117327, 7.601912, 6.121493, 10.05697, 
    12.49416,
  11.30817, 11.79304, 12.39173, 12.65334, 13.32368, 12.80299, 11.69232, 
    11.15589, 10.96466, 8.822965, 7.927328, 6.869347, 6.746801, 12.30256, 
    13.67844,
  11.17074, 11.2759, 12.03142, 12.93336, 13.18796, 11.00337, 9.625662, 
    10.24475, 8.881919, 6.30594, 6.512885, 6.333402, 7.595559, 13.65282, 
    13.42782,
  6.625301, 8.89212, 7.762812, 9.343493, 8.273619, 7.272513, 10.20242, 
    10.92672, 11.35407, 8.286463, 8.800984, 10.05715, 9.141253, 6.413385, 
    5.857602,
  11.10184, 12.00258, 11.83468, 11.82875, 6.744306, 6.225551, 10.95487, 
    11.0813, 12.19482, 10.82752, 11.37563, 13.4892, 11.75282, 6.688187, 
    7.140174,
  11.88845, 12.88545, 12.77495, 12.72132, 8.948559, 6.742779, 9.718802, 
    11.55487, 12.49443, 13.21125, 14.10242, 13.10239, 10.99843, 9.067344, 
    9.269227,
  13.14564, 13.50783, 13.33776, 13.10167, 13.04648, 10.38811, 6.174309, 
    7.634704, 11.5601, 12.82986, 12.53022, 10.33705, 9.426074, 8.110437, 
    12.27608,
  14.83334, 14.87486, 14.55936, 14.15139, 14.04841, 13.9235, 11.71986, 
    7.566143, 8.73385, 8.845694, 9.396373, 7.51696, 8.353271, 7.984799, 
    16.57927,
  15.78078, 16.24002, 16.06326, 15.56691, 15.24172, 15.12242, 15.08667, 
    14.58747, 10.03122, 6.683281, 4.61202, 6.281215, 7.817996, 8.154986, 
    17.41802,
  15.89349, 16.76593, 17.30622, 16.98684, 16.26775, 15.31625, 14.71073, 
    13.51446, 10.43163, 6.561673, 4.962882, 5.907629, 5.955707, 10.04854, 
    19.08859,
  15.50494, 16.3693, 17.20816, 17.122, 16.04718, 14.72211, 13.14512, 
    10.50895, 7.604319, 5.194164, 5.005634, 5.334955, 4.294208, 13.39679, 
    19.90398,
  15.78803, 16.1156, 16.29513, 16.08952, 15.34313, 14.1254, 11.85753, 
    9.233651, 6.788835, 5.104608, 4.974497, 4.271122, 5.723792, 17.44167, 
    18.82686,
  15.85969, 15.39067, 14.74842, 14.57602, 14.61853, 13.11474, 10.55615, 
    7.927144, 5.695101, 4.255054, 4.615034, 3.92905, 9.318294, 19.58301, 
    16.78276,
  9.933788, 12.65821, 11.24257, 13.80145, 12.30111, 10.08295, 12.54598, 
    11.56654, 10.57273, 7.667469, 7.511876, 8.302069, 8.129296, 8.534555, 
    6.823736,
  16.15931, 16.56067, 15.89706, 15.84477, 9.499352, 9.026053, 13.88717, 
    13.06617, 12.47969, 10.59854, 8.487925, 11.12936, 11.6029, 7.479361, 
    2.55328,
  15.4835, 17.55622, 17.14722, 16.82355, 12.34301, 8.675146, 12.11704, 
    13.85755, 13.45998, 12.26984, 12.2892, 12.11115, 10.7215, 5.914349, 
    3.309682,
  13.7468, 16.60781, 17.45683, 17.52727, 17.82786, 13.94304, 7.889194, 
    8.076578, 11.69442, 13.14598, 12.52414, 11.35028, 8.017682, 3.895845, 
    6.594779,
  12.15267, 14.20153, 16.06777, 17.17419, 18.1621, 18.51372, 14.7685, 
    8.730231, 7.611857, 8.051073, 10.17735, 9.59194, 5.900697, 4.94134, 
    8.950442,
  9.621774, 11.27717, 13.23008, 15.38003, 17.06361, 18.53966, 19.33559, 
    18.5282, 11.33856, 7.180701, 6.454403, 7.563016, 4.965694, 7.783786, 
    9.817017,
  7.978712, 8.655012, 10.13874, 12.26461, 14.48778, 16.51826, 18.21248, 
    18.66756, 16.13875, 12.36249, 10.16054, 7.253964, 7.470158, 10.66985, 
    11.75867,
  7.375381, 6.939651, 7.243153, 8.736205, 11.58589, 14.15222, 15.54365, 
    16.90335, 16.99602, 14.59442, 11.42233, 8.803438, 10.56639, 12.66793, 
    12.79961,
  7.669841, 8.342712, 8.449548, 8.015173, 9.424589, 12.14788, 14.49074, 
    15.75236, 16.25492, 15.90559, 13.44574, 11.72932, 13.44596, 14.57518, 
    12.67763,
  8.459513, 9.074997, 9.088686, 8.666931, 8.753317, 9.885716, 12.61034, 
    14.35803, 13.47221, 10.88045, 11.18572, 13.90406, 15.6469, 15.80281, 
    13.18674,
  10.53507, 13.81213, 11.94574, 14.3952, 12.73112, 10.17842, 12.92113, 
    11.11664, 9.548328, 6.529075, 5.274692, 5.081461, 3.634202, 2.739154, 
    2.182731,
  15.88103, 16.93533, 16.54018, 15.95482, 9.688957, 8.857731, 13.07265, 
    12.26188, 10.79427, 9.190517, 6.549015, 6.665135, 5.678386, 3.274041, 
    2.123763,
  14.51711, 16.92414, 17.12539, 16.95072, 12.38702, 7.468158, 11.18184, 
    12.92618, 12.55586, 10.66068, 9.277595, 8.236989, 6.963293, 5.707336, 
    4.160754,
  11.50323, 15.65891, 16.74015, 17.42009, 17.0694, 11.99293, 6.821496, 
    8.061968, 11.27119, 13.50099, 11.65208, 9.751763, 7.753398, 6.101208, 
    5.971642,
  4.800111, 12.37525, 15.17382, 16.45342, 16.83398, 15.63193, 12.92802, 
    8.206007, 7.456984, 8.786765, 12.1961, 11.90345, 9.43098, 8.065584, 
    8.629401,
  7.556304, 7.119095, 11.91586, 14.09033, 15.33095, 15.31718, 15.27237, 
    14.98405, 10.06956, 6.930941, 8.036343, 12.0801, 10.76402, 9.751755, 
    9.75551,
  11.18257, 7.292825, 7.969949, 11.25805, 13.42761, 14.13599, 14.1624, 
    13.62214, 11.94475, 10.55749, 10.73747, 10.97221, 11.14944, 11.41392, 
    11.37503,
  13.31545, 10.85856, 7.345004, 7.14051, 9.458675, 11.70789, 13.12237, 
    13.88353, 13.821, 12.61928, 11.03799, 10.44546, 11.52128, 12.06113, 
    12.64196,
  13.23089, 13.32898, 11.66756, 8.843334, 6.047236, 5.511981, 8.925636, 
    11.92062, 13.35341, 13.57493, 13.1056, 12.09149, 12.5753, 13.88732, 
    11.87183,
  10.99145, 11.42238, 11.36731, 10.74871, 9.464702, 7.189464, 4.998818, 
    8.141022, 10.02725, 9.570415, 11.05, 13.82693, 14.06514, 14.96818, 
    13.41595,
  8.795207, 12.3782, 10.89248, 13.71418, 12.61192, 10.3549, 13.1943, 
    11.38179, 9.047009, 5.209124, 3.878651, 3.363887, 2.812159, 2.923683, 
    2.908672,
  13.57544, 14.47375, 14.58335, 14.82623, 9.584759, 8.970145, 12.83235, 
    11.14922, 8.948199, 6.950897, 4.525833, 4.094559, 3.826272, 2.797491, 
    2.421081,
  14.05471, 14.63443, 15.32202, 15.64238, 11.73754, 7.908601, 10.26578, 
    11.25372, 9.197636, 7.852002, 6.289787, 4.660839, 3.808365, 3.942512, 
    3.802051,
  13.94312, 14.36011, 15.37662, 16.20254, 16.25041, 11.95909, 7.943214, 
    7.244525, 7.271747, 7.945628, 7.153072, 5.404304, 4.246294, 4.124661, 
    4.658284,
  12.78901, 13.7561, 14.86176, 15.85335, 15.79478, 15.06526, 13.60314, 
    8.286252, 5.778946, 6.321294, 8.165607, 7.062024, 5.470775, 5.08245, 
    5.468802,
  11.04743, 12.896, 14.12504, 15.1419, 15.4835, 15.11995, 15.32292, 14.94946, 
    9.743924, 7.137143, 7.198562, 8.634337, 7.022544, 5.930345, 5.518452,
  10.00281, 11.135, 12.74005, 13.94611, 14.36927, 14.13364, 13.92173, 
    13.12603, 11.91427, 11.57045, 11.51969, 10.12653, 8.581532, 7.280389, 
    6.559559,
  10.19691, 10.12998, 11.04492, 12.45471, 13.19777, 13.14301, 13.00797, 
    13.01015, 12.85564, 12.44147, 11.85908, 10.4292, 9.298297, 8.161758, 
    7.383453,
  11.15831, 10.26686, 9.981817, 10.82934, 11.82113, 12.27713, 12.41076, 
    12.09671, 11.74651, 11.4739, 11.02807, 10.45074, 9.405952, 8.903625, 
    8.04292,
  11.82749, 10.92708, 10.01278, 9.484623, 9.426197, 9.796538, 10.91043, 
    11.42128, 9.927733, 7.379477, 8.896763, 10.52864, 9.722097, 9.78341, 
    8.922286,
  9.452599, 12.98006, 11.6285, 13.74614, 11.21945, 8.323005, 10.39841, 
    9.045219, 7.354128, 4.862386, 4.209572, 4.464723, 4.251711, 4.472836, 
    3.95018,
  14.68249, 15.29392, 15.18658, 14.50186, 9.284927, 7.911421, 9.568761, 
    8.608979, 6.996227, 5.93079, 4.581549, 4.976616, 5.162025, 3.393904, 
    2.955565,
  15.65843, 15.90995, 15.74732, 15.16291, 10.55319, 7.731636, 7.76302, 
    7.647485, 7.589968, 6.457348, 5.883146, 5.090735, 4.775623, 4.110782, 
    3.120192,
  15.7864, 15.86171, 15.671, 15.11966, 14.49463, 10.68209, 7.240678, 
    6.459886, 5.947434, 4.614757, 5.072705, 4.649437, 4.386581, 4.128977, 
    3.533457,
  15.53266, 15.64848, 15.46731, 14.98409, 13.98057, 13.34422, 11.72714, 
    6.799212, 3.811605, 3.125094, 4.233134, 3.89051, 3.52036, 3.435049, 
    3.333896,
  15.19481, 15.19095, 15.03527, 14.55538, 13.93547, 12.97927, 12.02971, 
    11.04047, 6.953694, 4.986242, 3.9025, 3.738689, 2.898864, 2.619579, 
    2.61129,
  14.81435, 14.86941, 14.7503, 14.32115, 13.58946, 12.62997, 11.27038, 
    9.582026, 8.569566, 7.472483, 5.619496, 3.9083, 2.744471, 2.205692, 
    2.341427,
  14.33465, 14.34855, 14.22182, 13.92814, 13.3228, 12.35214, 11.18641, 
    10.34942, 9.994767, 8.680429, 5.91241, 4.007444, 2.755853, 2.246205, 
    2.374239,
  13.72146, 13.95815, 13.943, 13.61053, 12.97936, 12.15688, 11.19174, 
    10.09951, 9.495514, 8.352731, 6.295392, 4.728595, 3.320777, 2.583535, 
    2.408039,
  12.72478, 13.10186, 13.16407, 12.87173, 12.30914, 11.48973, 10.63854, 
    9.692298, 7.320133, 5.634081, 5.824599, 5.748517, 4.659431, 3.534706, 
    2.900959,
  8.821611, 12.31769, 10.91889, 12.86038, 10.02252, 6.705121, 7.797811, 
    6.838418, 6.829792, 4.689189, 4.53544, 4.800196, 4.31883, 4.469801, 
    3.947755,
  14.1002, 15.03809, 14.99109, 13.73376, 8.286025, 6.528049, 7.763775, 
    7.005268, 6.589719, 6.592489, 5.292912, 6.296979, 6.513326, 3.79323, 
    3.08339,
  15.51298, 15.78437, 15.20941, 13.27638, 9.417426, 5.962482, 6.610176, 
    7.226419, 7.431693, 6.928678, 7.032168, 6.816864, 6.865025, 5.400682, 
    3.295785,
  16.01206, 15.57276, 14.39143, 12.77821, 11.33545, 8.847858, 5.48155, 
    6.614786, 8.295982, 6.737206, 6.354203, 6.196559, 6.254618, 5.917451, 
    4.459803,
  15.89236, 15.08462, 13.54441, 12.17549, 10.63714, 9.866091, 8.73347, 
    5.114034, 3.683734, 3.748237, 5.405107, 5.957911, 6.099414, 6.15745, 
    5.76349,
  15.65649, 14.56016, 13.05368, 11.74521, 10.68734, 9.122016, 7.828803, 
    7.622077, 5.297106, 4.338067, 4.369934, 5.679711, 5.942047, 6.066928, 
    5.988472,
  15.17448, 14.17878, 12.96048, 11.78843, 10.61898, 9.733332, 8.56543, 
    7.376866, 6.768492, 6.00803, 5.178163, 5.336498, 5.786472, 5.984608, 
    5.962976,
  14.46385, 13.51296, 12.48295, 11.53366, 10.68401, 9.919669, 9.342472, 
    8.780301, 7.472868, 5.586813, 4.350157, 4.666945, 5.391687, 5.798042, 
    5.94753,
  13.98966, 13.12837, 12.21381, 11.18881, 10.35981, 9.577111, 8.726908, 
    7.862006, 6.530579, 4.198808, 2.948997, 3.542589, 4.680887, 5.480787, 
    5.507384,
  13.50019, 12.63887, 11.64283, 10.6234, 9.752617, 8.827191, 8.00005, 
    7.216578, 5.085736, 2.495184, 1.612204, 2.128819, 3.494503, 4.711443, 
    4.975122,
  6.728757, 8.147712, 6.170547, 6.799247, 5.704941, 4.880224, 5.902358, 
    5.139315, 5.369965, 3.555717, 2.672221, 2.823961, 2.475358, 2.263283, 
    1.219485,
  11.03688, 10.1212, 8.786245, 7.359347, 4.823533, 5.052986, 6.324285, 
    5.454534, 4.548089, 4.201579, 2.75328, 2.762166, 2.601413, 1.713213, 
    1.72956,
  12.3827, 11.12186, 9.588739, 7.516456, 5.782145, 3.898915, 5.880213, 
    6.28347, 6.118073, 5.070289, 3.999526, 3.133857, 2.641419, 2.422504, 
    2.123543,
  13.29441, 11.89831, 9.998307, 7.939179, 6.252542, 5.361948, 3.260715, 
    6.116264, 9.001148, 6.937958, 5.038215, 3.855915, 3.361399, 3.151822, 
    3.096666,
  13.93069, 12.5054, 10.48552, 8.830971, 7.104262, 6.040783, 5.534213, 
    3.859468, 4.419138, 4.70421, 5.775234, 5.449029, 4.844855, 4.581464, 
    4.610788,
  14.50081, 12.94758, 10.98328, 9.564906, 8.760123, 8.071887, 7.582042, 
    7.867118, 5.221982, 5.173984, 5.091115, 6.64377, 6.575989, 6.054911, 
    6.063668,
  15.11964, 13.5637, 11.73321, 10.30744, 9.303561, 9.088362, 9.097093, 
    8.970995, 8.714294, 8.694756, 8.147498, 7.800386, 7.445484, 6.974812, 
    6.829509,
  15.49419, 13.94308, 12.15519, 10.64832, 9.582995, 9.07359, 8.966394, 
    9.03823, 8.727248, 8.380873, 8.323791, 8.23402, 7.806643, 7.170681, 
    6.938352,
  15.55497, 14.17484, 12.66005, 11.07614, 9.805412, 9.103462, 8.609062, 
    8.14728, 7.362037, 6.406685, 7.636694, 8.296654, 7.964424, 7.547935, 
    6.777685,
  15.28154, 13.9483, 12.46241, 11.06001, 9.786561, 8.774542, 8.040922, 
    6.83439, 4.53103, 3.571654, 5.006527, 6.917425, 7.355923, 7.532188, 
    6.948447,
  2.877916, 3.887151, 4.358409, 5.219018, 5.125987, 3.933498, 4.422589, 
    4.066279, 3.946617, 3.118062, 3.024786, 3.201781, 3.427574, 4.051334, 
    3.923789,
  4.574678, 4.477252, 5.093381, 4.943259, 3.993018, 3.217078, 3.495749, 
    3.420838, 3.000762, 3.160627, 3.072101, 3.616342, 4.245287, 2.848728, 
    2.283664,
  5.453144, 4.988551, 5.161579, 4.788857, 4.436731, 2.8831, 2.556519, 
    2.87751, 3.632665, 3.648766, 3.570765, 3.51329, 3.574361, 3.303128, 
    2.77497,
  6.068575, 5.389724, 4.995412, 4.573144, 4.157423, 3.996412, 2.447966, 
    2.865775, 3.140942, 2.987136, 3.410201, 3.172933, 3.106349, 3.27422, 
    3.366542,
  6.255103, 5.311456, 4.642572, 4.860518, 4.581818, 4.386791, 4.829395, 
    3.106485, 2.432781, 2.629051, 3.312728, 2.789299, 2.640357, 3.063554, 
    3.509854,
  6.742918, 5.675108, 5.306985, 5.710961, 6.147413, 6.150396, 5.453024, 
    5.349364, 4.320163, 4.259852, 3.510707, 3.650672, 3.484182, 3.487159, 
    3.298296,
  7.626903, 6.969211, 7.04009, 7.374471, 7.448542, 7.836269, 7.713606, 
    7.24923, 6.960192, 6.748695, 5.917163, 5.269191, 5.013624, 4.637047, 
    4.016048,
  8.948431, 8.401247, 8.36723, 8.566689, 8.687982, 8.835045, 8.905384, 
    9.047201, 8.748063, 8.120332, 7.305586, 6.819829, 6.133954, 5.496637, 
    5.058713,
  10.34517, 9.777559, 9.673077, 9.543628, 9.553405, 9.775242, 9.861247, 
    9.802382, 9.420077, 8.744149, 8.186292, 7.742255, 6.93927, 6.160931, 
    5.751076,
  11.57132, 10.84821, 10.53247, 10.07726, 9.8829, 9.933119, 9.846784, 
    9.436724, 7.898309, 6.036477, 6.95455, 8.381855, 7.622452, 7.221158, 
    6.963759,
  3.335619, 4.470774, 4.240438, 4.475117, 4.404743, 3.656412, 4.307695, 
    4.945157, 6.081208, 4.609704, 4.137146, 4.379149, 4.53878, 4.615223, 
    3.663192,
  5.104657, 5.293906, 5.612199, 5.084558, 3.922319, 3.767744, 5.58571, 
    5.893099, 6.321672, 6.353576, 5.263125, 6.200865, 6.651719, 3.993236, 
    3.11519,
  6.093085, 5.862292, 6.258246, 5.651607, 4.881969, 3.391047, 5.123896, 
    6.239788, 7.04435, 7.132771, 7.258382, 6.98734, 7.069365, 5.985178, 
    4.283758,
  6.492162, 6.360064, 6.672876, 6.128659, 5.419173, 5.007086, 3.319345, 
    5.481227, 7.113928, 6.227323, 6.47865, 6.409046, 7.118417, 6.70739, 
    5.280425,
  6.309049, 6.368866, 6.675573, 6.663342, 5.698852, 5.427164, 5.721449, 
    3.501919, 2.826425, 3.196538, 5.173428, 5.659424, 6.515531, 7.043604, 
    6.241021,
  6.00472, 6.080722, 6.370679, 6.673189, 6.560117, 6.045398, 4.833586, 
    4.659303, 4.52387, 4.547173, 4.093446, 5.594453, 6.514779, 6.96488, 
    6.897085,
  5.49628, 6.112801, 6.659997, 6.842581, 6.745775, 6.799117, 5.843897, 
    4.935636, 5.962698, 6.091784, 5.652363, 6.026951, 6.635975, 6.838905, 
    7.421294,
  5.266018, 6.45886, 7.065618, 7.290513, 7.159855, 7.001899, 6.609081, 
    7.192396, 7.460733, 6.396111, 5.988758, 6.387019, 6.768728, 6.961679, 
    7.244202,
  6.233857, 6.781129, 7.282741, 7.737492, 7.827112, 7.68272, 7.212209, 
    7.383795, 7.258308, 6.232535, 6.040255, 6.433602, 6.614677, 6.409842, 
    6.276367,
  7.832005, 7.525564, 7.666486, 7.796147, 7.842931, 7.84158, 7.868649, 
    8.127973, 6.695982, 4.71712, 5.111824, 6.397648, 6.084348, 6.121185, 
    6.106122,
  2.727513, 3.057782, 2.41794, 1.614102, 1.070556, 1.344373, 1.845106, 
    3.387569, 3.627873, 2.347124, 2.639998, 3.669566, 4.852737, 5.349071, 
    5.263632,
  4.787024, 4.027852, 3.274884, 2.3795, 1.338347, 1.15243, 2.746649, 
    4.049634, 3.349849, 3.141841, 3.93171, 5.652477, 7.869774, 5.383318, 
    5.544972,
  5.800302, 4.758123, 4.084091, 3.597857, 3.541863, 2.168608, 3.242952, 
    4.555606, 4.826348, 4.607606, 5.934554, 7.274, 8.70306, 9.089025, 6.792384,
  5.839255, 4.787525, 4.250532, 4.435947, 5.194077, 5.141035, 3.571761, 
    4.254959, 4.587669, 4.453236, 6.733381, 8.143724, 9.258108, 8.752545, 
    7.420877,
  5.576928, 4.419581, 3.893764, 4.812487, 6.240184, 7.158648, 7.160936, 
    4.12572, 2.772563, 3.476779, 6.8266, 8.240338, 8.938691, 8.399037, 
    7.210883,
  5.835958, 4.199329, 3.567139, 4.569503, 6.695174, 7.511875, 6.948668, 
    6.925098, 5.686877, 5.928953, 5.977744, 8.414628, 8.409579, 7.936109, 
    6.888884,
  6.596471, 4.598547, 3.828641, 4.777802, 6.320497, 7.555854, 7.326709, 
    6.288394, 7.013359, 8.691356, 9.186293, 8.917722, 8.206024, 7.627962, 
    6.975707,
  7.031204, 5.470532, 4.50556, 4.962167, 5.860204, 6.641663, 7.308558, 
    8.009643, 8.761809, 9.192736, 9.427551, 9.031349, 8.093757, 7.439781, 
    6.734225,
  7.407891, 6.876673, 5.996043, 5.741712, 5.793577, 6.157464, 6.596757, 
    7.247196, 8.008742, 8.454264, 9.010232, 9.04809, 8.247993, 7.366148, 
    6.395943,
  7.071911, 7.25576, 6.71623, 6.238706, 5.799571, 5.756391, 6.326362, 
    7.334568, 6.877538, 5.821237, 6.786254, 8.737785, 8.092598, 7.340611, 
    6.065463,
  2.302125, 1.851819, 1.43337, 1.691342, 2.821304, 2.905954, 2.475193, 
    3.020563, 4.95934, 4.303277, 4.319345, 5.07442, 5.149148, 4.769101, 
    3.759285,
  4.739063, 3.616827, 2.412315, 1.511436, 1.163516, 2.656148, 3.461298, 
    3.600093, 4.990138, 5.762995, 5.622266, 7.177761, 8.256675, 5.00168, 
    4.465124,
  6.193068, 5.320297, 3.821065, 2.925823, 2.113084, 1.456936, 3.406395, 
    4.024582, 5.810246, 7.030046, 7.70363, 8.194421, 8.619103, 8.818347, 
    6.642051,
  6.804006, 6.302518, 5.159836, 4.158542, 4.140164, 3.680923, 2.364603, 
    4.352736, 5.78902, 6.133068, 7.670924, 8.103686, 8.545318, 8.763005, 
    7.892977,
  7.286888, 7.079848, 6.58071, 5.592402, 5.037032, 5.361502, 5.66861, 
    3.163067, 3.014385, 3.962035, 6.896755, 8.268991, 8.837288, 9.00011, 
    8.475509,
  7.603891, 7.391159, 7.330003, 6.611641, 5.831407, 5.834344, 5.295797, 
    5.904655, 6.131726, 6.150195, 5.943997, 8.27549, 8.476727, 8.073443, 
    6.993065,
  7.932022, 7.27595, 7.272453, 6.955346, 6.542816, 6.659534, 6.152423, 
    5.440571, 7.164161, 8.774301, 8.975342, 8.684999, 8.175191, 7.517272, 
    6.867205,
  7.65209, 6.693993, 6.514706, 6.553618, 6.734885, 7.141614, 7.672427, 
    7.74411, 9.04628, 9.599806, 9.044706, 8.639642, 7.784476, 6.970946, 
    6.329457,
  6.939447, 5.886223, 5.239722, 5.541336, 6.292967, 7.104992, 8.107007, 
    8.360312, 9.058558, 9.206329, 9.018354, 8.927591, 7.918163, 7.128999, 
    6.280744,
  6.156184, 5.009859, 3.903802, 3.960182, 4.915304, 6.042461, 7.509832, 
    8.810735, 8.05848, 6.597198, 7.559814, 9.487432, 8.642241, 7.841495, 
    6.766576,
  4.24707, 3.894601, 2.257605, 1.412062, 2.418081, 2.684268, 3.729996, 
    5.40864, 5.728465, 4.12135, 3.710292, 4.140296, 3.732939, 3.581819, 
    2.639356,
  8.12765, 6.287553, 4.109758, 2.954367, 2.078735, 2.182733, 2.738638, 
    4.900996, 5.494711, 5.157476, 4.463889, 5.383476, 5.670745, 3.448851, 
    2.755323,
  10.33105, 8.737659, 6.290479, 5.302821, 4.870192, 2.495605, 1.982876, 
    3.61882, 5.748445, 5.827265, 5.881162, 5.886376, 5.488771, 5.081911, 
    4.41057,
  11.70905, 10.31925, 8.457672, 6.828404, 7.219581, 6.255108, 3.200402, 
    2.874284, 4.292223, 5.46237, 6.106308, 5.568045, 4.932693, 5.041993, 
    5.623415,
  12.81311, 11.34177, 9.970357, 8.445135, 7.387453, 8.007514, 8.260699, 
    4.547458, 3.926958, 4.71793, 6.519042, 6.688731, 6.061857, 6.183039, 
    6.51305,
  13.5727, 12.16886, 10.83936, 9.274436, 7.57396, 6.111149, 9.093417, 
    10.30744, 7.611401, 6.44903, 6.466471, 7.923512, 7.025536, 6.41455, 
    5.949041,
  14.08243, 12.77255, 11.45234, 9.920246, 8.217665, 5.936601, 6.751862, 
    9.201102, 8.607762, 8.500299, 9.558154, 8.859536, 8.173466, 7.32053, 
    6.803397,
  14.10242, 12.61978, 11.36535, 10.1908, 8.88888, 7.12106, 6.104572, 
    7.712955, 9.149765, 8.956078, 8.876501, 8.931355, 8.661837, 7.889489, 
    7.344817,
  13.38115, 12.0087, 11.02439, 10.13095, 9.152685, 7.759895, 6.759411, 
    7.353514, 8.462098, 8.745256, 9.002451, 9.384735, 9.079586, 8.502905, 
    7.934688,
  11.8581, 10.80887, 9.990682, 8.969954, 8.243933, 7.219577, 6.477086, 
    6.94279, 7.350188, 6.579314, 7.762341, 9.787004, 9.474783, 9.361604, 
    8.47613,
  7.861219, 10.5078, 8.471923, 8.400023, 6.682885, 5.462821, 6.454357, 
    6.100238, 5.567243, 3.306887, 2.40759, 2.524601, 2.903514, 3.035965, 
    2.369992,
  12.62517, 13.22704, 12.46056, 10.48392, 6.135742, 4.325557, 6.030329, 
    5.75934, 5.084354, 4.414742, 3.101997, 3.356293, 3.722476, 2.903048, 
    2.515958,
  13.7513, 14.7249, 14.31552, 12.68136, 8.395199, 4.696376, 4.678191, 
    5.187902, 5.561729, 5.330248, 4.680349, 3.756874, 3.046133, 3.941985, 
    4.013772,
  14.32669, 15.53174, 15.44537, 14.62682, 12.93435, 8.589915, 4.747694, 
    3.435293, 2.637201, 5.240236, 5.310302, 4.241799, 3.399225, 3.822554, 
    4.871112,
  14.45116, 16.05655, 16.33157, 15.6313, 13.86455, 12.19911, 10.36315, 
    5.691713, 4.058506, 4.801772, 6.707791, 6.262732, 4.632974, 4.543796, 
    5.110238,
  14.08505, 16.17109, 16.81497, 16.18398, 14.60804, 12.85464, 12.27267, 
    11.49351, 7.336947, 5.568216, 6.701585, 8.143634, 6.276954, 5.205665, 
    4.583521,
  13.49644, 16.1312, 17.20774, 16.71897, 15.21474, 13.13933, 11.26567, 
    10.11699, 8.095286, 7.411946, 9.263832, 8.865833, 7.799305, 6.675035, 
    5.731863,
  12.27765, 15.29707, 17.11963, 16.93466, 15.59037, 13.58174, 11.26251, 
    9.902955, 9.419246, 8.843742, 8.69659, 8.580898, 8.261411, 7.652758, 
    6.772656,
  11.14595, 14.46136, 16.71124, 16.83452, 15.69238, 13.86314, 11.63424, 
    9.066199, 7.607964, 8.788702, 9.423533, 9.392904, 8.729736, 8.148793, 
    7.375465,
  9.550482, 12.98909, 15.63576, 15.93984, 15.07193, 13.63776, 11.61937, 
    8.308141, 5.834369, 5.739212, 7.644213, 10.06318, 9.610602, 9.158321, 
    8.066476,
  5.880562, 7.871939, 8.559533, 12.18568, 10.73283, 7.551363, 7.985775, 
    6.77611, 5.537259, 3.423825, 3.319194, 3.994794, 3.937322, 3.663971, 
    2.818582,
  8.382029, 9.589155, 11.22013, 13.06451, 8.473191, 5.651058, 7.6521, 
    6.743192, 5.300725, 4.45689, 3.800104, 5.020876, 5.765537, 3.504958, 
    2.935683,
  8.732265, 10.3868, 12.72569, 14.28921, 10.89351, 6.518816, 6.19315, 
    6.32078, 6.163787, 5.505935, 4.944619, 5.135676, 5.280081, 5.081861, 
    4.327011,
  8.631247, 10.54086, 13.77115, 15.75401, 15.44275, 10.9664, 6.69433, 
    4.40503, 3.296028, 5.060137, 5.050373, 4.901776, 4.837355, 4.9508, 
    5.269675,
  8.216253, 10.10795, 14.13444, 16.02445, 15.68628, 14.50348, 12.58171, 
    6.979485, 4.281396, 4.338681, 6.006359, 5.717394, 4.86169, 5.377679, 
    5.791367,
  7.993406, 9.435381, 13.91115, 15.94281, 15.80567, 15.08393, 14.66297, 
    13.06109, 7.54801, 5.775455, 6.06388, 7.001246, 5.644043, 5.120922, 
    5.01706,
  7.832979, 8.726234, 13.52898, 15.82017, 15.61249, 14.94724, 13.60779, 
    10.98956, 7.971509, 8.085602, 8.849312, 7.707707, 6.729415, 5.781129, 
    5.259496,
  7.020667, 7.584414, 12.65632, 15.48968, 15.3851, 14.603, 13.72872, 
    12.59349, 10.83363, 9.218384, 8.306968, 7.637958, 7.177593, 6.33272, 
    5.621321,
  5.649923, 6.157523, 11.53938, 15.08162, 15.04088, 14.37391, 13.61662, 
    12.40011, 10.34799, 8.445848, 8.114645, 7.95319, 7.461242, 6.895094, 
    5.935649,
  3.973242, 4.921639, 9.674673, 14.16089, 14.29818, 13.77507, 13.29327, 
    12.29614, 8.465993, 6.195182, 6.8126, 8.296908, 7.963631, 7.447773, 
    6.617007,
  5.839097, 7.767067, 6.047562, 8.16014, 8.389047, 6.858011, 8.918523, 
    8.824747, 7.849889, 4.907332, 4.257459, 4.700275, 4.332245, 3.822458, 
    3.123525,
  8.57812, 7.813663, 7.729199, 9.821604, 8.290367, 6.076345, 7.797724, 
    8.15948, 7.359007, 6.110617, 5.054885, 6.243737, 6.857506, 3.950485, 
    3.143384,
  9.900608, 7.370914, 8.703374, 12.52251, 10.64708, 6.789098, 6.474343, 
    7.229965, 7.674582, 6.851814, 6.458362, 6.531173, 6.5347, 6.245239, 
    4.849757,
  10.4972, 7.538527, 9.588696, 14.31067, 15.01069, 11.05813, 7.145831, 
    5.249508, 4.627479, 5.675888, 6.382882, 6.348921, 6.022473, 5.894065, 
    5.997695,
  9.857825, 7.175072, 9.06354, 14.13899, 14.86155, 13.90774, 12.71368, 
    7.19388, 4.194857, 4.342322, 6.510937, 6.731597, 6.415232, 6.547609, 
    6.578607,
  8.305125, 6.5877, 7.867459, 13.48471, 14.54837, 13.34579, 13.56544, 
    12.67198, 7.794148, 6.374915, 6.18995, 7.289944, 6.682051, 6.120767, 
    5.595904,
  5.672099, 5.25224, 6.219098, 12.86172, 14.40201, 12.93868, 11.71488, 
    9.769508, 8.350676, 9.261846, 9.066932, 7.861595, 7.076093, 6.15863, 
    5.58787,
  3.738698, 4.179608, 4.831912, 12.17375, 14.30728, 12.95924, 12.34227, 
    11.58175, 10.6146, 9.909423, 8.912461, 7.995789, 7.123761, 6.01428, 
    5.319082,
  3.130254, 4.366344, 4.399421, 11.86948, 14.13635, 12.96502, 12.4774, 
    11.53084, 10.33734, 8.777138, 8.348053, 8.068311, 7.26598, 6.141002, 
    5.261745,
  3.652116, 4.310866, 4.322384, 12.66872, 13.48687, 12.11084, 12.26486, 
    11.7888, 8.271675, 6.189666, 6.871573, 8.341354, 7.598471, 6.713354, 
    5.589857,
  8.895617, 11.38966, 8.437229, 8.980242, 5.85453, 4.797215, 7.165349, 
    8.685318, 9.496642, 6.152259, 4.874162, 4.739924, 3.610005, 2.940481, 
    2.718281,
  12.79487, 12.96796, 11.34474, 9.246323, 5.169561, 5.484601, 6.446891, 
    7.884461, 8.797247, 7.950727, 5.817205, 6.381366, 5.921828, 2.993968, 
    2.228096,
  11.50912, 12.07256, 11.53891, 10.7661, 8.332661, 7.602123, 5.812239, 
    6.428265, 8.347151, 8.636318, 7.682037, 6.959749, 5.89752, 4.802031, 
    3.591634,
  10.78272, 11.02136, 11.39592, 12.45963, 13.62328, 11.37059, 7.9446, 
    5.261195, 4.767939, 6.745978, 7.358379, 6.827299, 5.76002, 4.903977, 
    4.677398,
  9.663803, 10.40054, 11.07242, 12.66924, 14.51031, 14.50291, 12.71087, 
    8.289728, 5.069082, 5.230855, 7.314806, 7.401412, 6.655904, 6.010241, 
    5.314946,
  5.4956, 7.731597, 9.98372, 12.24633, 14.15051, 13.64473, 12.47402, 
    11.47059, 8.851384, 8.02397, 6.855247, 8.097767, 7.098215, 6.003314, 
    5.126198,
  2.54684, 4.237545, 7.729001, 11.44271, 13.75696, 12.41875, 9.129221, 
    7.125559, 9.310932, 11.48629, 10.0748, 8.735577, 7.600688, 6.394137, 
    5.689399,
  4.073161, 4.041876, 7.026491, 11.28358, 13.64359, 12.39177, 10.56406, 
    10.03975, 11.10972, 11.0615, 9.562682, 8.575883, 7.554519, 6.400938, 
    5.500429,
  5.368705, 5.658418, 7.867544, 11.95021, 13.60579, 12.06443, 10.71421, 
    10.69934, 11.34084, 9.716097, 8.813335, 8.267971, 7.362853, 6.392867, 
    5.272295,
  5.807045, 6.55253, 9.296298, 12.76416, 13.11293, 11.49898, 11.24824, 
    11.68311, 9.168622, 6.423991, 6.920878, 8.01168, 7.195494, 6.48683, 
    5.480461,
  9.291058, 12.6029, 9.72068, 11.29859, 9.830462, 7.362054, 8.742034, 
    7.910439, 7.81055, 6.245427, 5.82114, 6.334308, 5.197194, 3.533327, 
    2.995494,
  11.67847, 12.56745, 11.64202, 10.31243, 5.870804, 4.919988, 6.371441, 
    6.902138, 7.734049, 7.708408, 6.875756, 8.280399, 7.468118, 3.794744, 
    3.267843,
  9.08332, 10.18539, 10.596, 9.688328, 6.556779, 4.855489, 4.662786, 
    5.437953, 7.717808, 9.073013, 9.047544, 8.824284, 7.244364, 4.534768, 
    3.155366,
  7.839289, 8.524514, 9.525136, 10.26561, 10.41453, 8.062525, 6.287494, 
    5.128244, 4.979869, 6.755024, 8.511065, 7.955365, 6.137851, 3.429316, 
    2.466045,
  7.205176, 7.768897, 8.898479, 10.4172, 11.3647, 11.17158, 10.10961, 
    6.809333, 3.978314, 4.667311, 7.792432, 7.922721, 6.306642, 3.604276, 
    2.234044,
  5.135448, 5.317132, 7.815398, 10.49615, 11.88845, 10.96343, 10.04997, 
    9.58745, 7.125926, 6.965603, 7.141756, 8.548489, 6.697217, 3.627453, 
    2.214212,
  3.720038, 2.995456, 6.83181, 11.45037, 11.87531, 10.42301, 8.164786, 
    6.084878, 7.255379, 10.48711, 10.73178, 9.220748, 7.064221, 4.111246, 
    2.42021,
  4.525662, 4.006391, 8.51537, 12.11833, 11.50779, 10.14535, 8.81671, 
    8.219898, 9.059975, 10.51993, 10.22009, 9.176188, 7.078311, 4.452853, 
    2.974844,
  11.18315, 10.35657, 12.1575, 12.22811, 10.79515, 9.742363, 8.796161, 
    8.866441, 9.581351, 9.558532, 9.443902, 8.78937, 7.111765, 4.914725, 
    3.346168,
  15.72618, 14.60607, 13.19917, 11.69217, 10.55463, 10.35034, 10.64956, 
    10.78821, 8.928448, 6.748058, 7.247637, 8.431788, 6.941093, 5.148037, 
    3.639045,
  8.589997, 11.78567, 10.0555, 12.18091, 10.93116, 8.742011, 10.64785, 
    9.916585, 8.767631, 5.483337, 5.229387, 5.723007, 5.447008, 5.721446, 
    5.715511,
  11.5929, 13.7112, 13.7077, 13.22782, 7.594492, 6.703971, 9.822159, 
    8.844158, 8.311103, 7.037801, 5.685511, 7.407275, 8.260503, 5.675547, 
    5.141064,
  9.134246, 11.14571, 12.67955, 12.8151, 9.315285, 5.681967, 6.687533, 
    6.752685, 6.417387, 6.853599, 7.074884, 7.50953, 8.448064, 8.927131, 
    7.419007,
  7.92367, 8.435283, 9.386366, 10.50418, 12.03665, 8.716913, 4.013165, 
    3.181226, 3.471663, 4.726052, 6.151625, 7.18096, 7.810943, 8.376506, 
    7.987623,
  7.768876, 7.023847, 6.758883, 7.732458, 10.01978, 10.77923, 8.24627, 
    4.712191, 2.912263, 3.305221, 5.742612, 7.766065, 8.578366, 9.026924, 
    9.467457,
  8.026958, 6.629237, 4.766871, 4.721602, 7.286209, 9.039314, 7.932282, 
    7.077328, 5.747453, 5.27871, 5.786669, 8.64974, 8.842858, 8.27484, 7.5942,
  9.521709, 9.884056, 7.862948, 7.938314, 10.39852, 9.393473, 6.712989, 
    5.056853, 6.138112, 7.704525, 8.675035, 9.544795, 8.906872, 7.777997, 
    6.620601,
  9.171968, 10.70298, 11.74608, 11.92285, 10.6961, 8.724646, 7.630558, 
    7.811148, 7.778371, 7.67639, 8.721936, 9.435916, 8.222692, 6.625766, 
    5.230736,
  8.279612, 8.629157, 9.079409, 9.292394, 8.696535, 8.028303, 7.783595, 
    8.094641, 7.934926, 7.464917, 8.389536, 8.553215, 7.236615, 5.42321, 
    4.210852,
  9.51403, 9.460857, 9.243361, 8.917013, 8.542821, 8.141731, 8.344992, 
    8.312265, 6.763889, 5.415628, 6.555961, 7.809352, 6.354362, 4.13155, 
    3.657389,
  4.924578, 8.218732, 7.665888, 10.22308, 9.291537, 8.051071, 10.20482, 
    9.919801, 9.420779, 6.198598, 5.819244, 6.649394, 5.992643, 5.422652, 
    5.311869,
  4.712364, 7.123869, 8.710311, 10.18235, 6.763952, 6.801691, 10.05799, 
    9.172796, 8.810289, 7.581461, 6.409682, 8.067238, 8.446638, 5.423975, 
    4.793713,
  6.018211, 6.621734, 7.272404, 8.267639, 6.977053, 5.637906, 7.290514, 
    8.411089, 8.305216, 8.209365, 8.273726, 7.923851, 8.260628, 7.646031, 
    5.975302,
  7.110886, 8.343338, 8.297446, 7.132611, 7.996524, 7.014221, 3.947145, 
    3.494801, 5.256433, 7.730227, 7.902313, 7.068445, 6.711743, 6.818763, 
    7.054543,
  6.882226, 8.661888, 8.744613, 7.475801, 5.886613, 8.050939, 7.289742, 
    4.132585, 4.068218, 5.472119, 7.814561, 7.538503, 6.865985, 7.391201, 
    9.048898,
  6.253427, 8.661381, 9.426735, 9.349397, 7.296642, 5.802363, 5.80281, 
    4.755908, 4.210639, 4.723291, 6.479745, 8.211772, 7.675992, 7.749981, 
    8.702809,
  4.802395, 7.674612, 9.2999, 10.24239, 10.25261, 8.476569, 5.87923, 
    3.868314, 3.147388, 5.692359, 8.553767, 9.054599, 8.923697, 9.099156, 
    9.845649,
  3.735114, 5.886822, 7.553457, 8.544281, 8.772363, 8.291295, 7.579453, 
    7.283876, 5.980511, 5.638488, 8.120025, 9.492843, 9.794854, 10.18993, 
    10.43624,
  4.103688, 5.058459, 6.402925, 7.305828, 7.569199, 7.382584, 7.3166, 
    7.731902, 7.325851, 7.121349, 8.334328, 9.650839, 10.50718, 10.80243, 
    9.225475,
  5.148306, 5.288192, 6.032767, 6.820711, 6.936125, 6.431073, 6.383383, 
    6.604459, 5.640278, 5.014345, 6.750042, 9.667536, 10.47979, 10.50399, 
    8.6068,
  1.95126, 3.890397, 4.051109, 6.340527, 6.635725, 5.884193, 7.102674, 
    6.331611, 5.718166, 3.907724, 3.707589, 4.440774, 4.510697, 4.802792, 
    5.128998,
  1.769526, 3.281513, 4.447633, 5.645931, 4.275019, 4.691635, 6.945122, 
    6.373693, 6.035481, 5.593698, 4.790101, 5.63553, 6.571523, 4.523042, 
    4.5352,
  2.206552, 4.477715, 4.977884, 5.231035, 4.082056, 3.339027, 4.740393, 
    4.749286, 4.704863, 5.785641, 6.461643, 6.334168, 6.871462, 7.17376, 
    5.92737,
  1.969861, 4.398706, 6.527816, 7.318563, 5.658043, 3.605853, 2.392074, 
    3.187484, 3.720573, 4.900344, 6.06636, 6.188241, 6.313978, 6.724384, 
    7.244533,
  1.766885, 3.409473, 5.979143, 7.531456, 7.716484, 6.451503, 4.047099, 
    2.146026, 3.305344, 4.022179, 5.598476, 6.611527, 6.785377, 7.393089, 
    8.226617,
  2.470508, 2.939265, 5.46442, 7.371833, 7.892899, 7.405473, 5.982249, 
    4.300996, 4.43799, 3.859216, 4.019189, 6.051015, 6.858758, 6.993656, 
    7.319333,
  3.649887, 3.237666, 5.532919, 7.331959, 7.814179, 7.246213, 6.534157, 
    6.159909, 5.902369, 3.881433, 3.854581, 5.718704, 6.918921, 7.358212, 
    7.650434,
  4.196799, 4.030068, 6.416598, 7.516764, 7.732657, 6.993893, 6.082221, 
    5.950402, 5.647569, 4.024989, 3.68268, 5.865267, 7.199618, 7.901174, 
    8.293525,
  4.169679, 5.468691, 7.406497, 7.557376, 7.442039, 6.573332, 5.397388, 
    5.285844, 4.713102, 3.797276, 3.286231, 6.07333, 7.617061, 8.96474, 
    8.74495,
  5.296374, 7.82111, 8.597513, 7.720603, 7.167897, 6.21358, 4.338688, 
    4.059829, 3.152551, 2.286671, 3.198566, 6.610484, 8.616172, 9.653437, 
    8.51845,
  2.605921, 2.152991, 2.667245, 4.733387, 5.964045, 6.086497, 8.830505, 
    8.851597, 6.895988, 4.395713, 4.221075, 4.419935, 3.600956, 3.304041, 
    3.609279,
  3.967503, 3.060782, 4.043332, 6.257998, 5.386803, 6.337051, 9.039639, 
    9.378992, 8.286767, 5.508854, 4.569724, 5.076075, 4.771149, 3.155638, 
    3.102716,
  4.883531, 4.695889, 5.820492, 7.738281, 6.622588, 6.066204, 8.121935, 
    8.857442, 7.501038, 5.633254, 5.301751, 5.028364, 4.227845, 4.383569, 
    3.657127,
  5.051993, 5.955008, 8.491395, 11.17093, 11.52007, 8.760118, 7.145154, 
    6.51173, 5.978065, 5.476351, 5.283985, 4.543087, 3.434781, 3.594624, 
    4.314188,
  5.141493, 7.360495, 10.25823, 13.07317, 14.48495, 13.3618, 9.465333, 
    4.293832, 3.858016, 3.912107, 4.677895, 3.837749, 3.33803, 4.033847, 
    5.15419,
  6.537518, 9.169109, 11.9389, 13.99374, 14.61854, 13.00986, 9.094267, 
    5.639819, 3.797319, 3.758581, 3.287241, 2.518277, 2.402032, 4.338387, 
    4.97391,
  7.878586, 10.62354, 12.73755, 13.73209, 12.687, 10.12236, 7.938677, 
    5.098709, 3.666939, 4.572064, 3.155543, 1.473099, 1.757583, 4.831894, 
    5.528393,
  8.262756, 11.2311, 12.79678, 12.91387, 10.1517, 7.558726, 7.357684, 
    5.419947, 3.784616, 3.817076, 1.943574, 0.9700216, 2.655376, 5.023011, 
    5.88532,
  9.11334, 11.79431, 12.54489, 11.75776, 8.048891, 6.170735, 6.861265, 
    4.905568, 4.232346, 3.060604, 1.275396, 1.914632, 4.01428, 5.865089, 
    6.191621,
  9.620073, 11.26613, 11.43688, 10.61592, 7.250388, 5.604003, 6.091016, 
    3.278339, 3.314796, 2.395619, 1.560881, 3.050135, 4.746294, 6.057144, 
    5.730482,
  3.36732, 2.298503, 4.128647, 7.360623, 8.161851, 8.024634, 11.03662, 
    12.94737, 12.80564, 9.44072, 9.476556, 9.381746, 7.894847, 6.343388, 
    5.755483,
  3.05326, 4.09707, 6.818953, 8.70939, 7.010116, 7.46797, 10.52843, 11.25533, 
    11.40607, 10.35702, 8.728272, 9.287934, 6.870952, 4.606439, 5.24388,
  3.345664, 7.161252, 8.99044, 9.110828, 6.141913, 5.43284, 7.96771, 
    8.841794, 9.769118, 10.03628, 9.240612, 8.441886, 9.568735, 9.221061, 
    7.130671,
  5.735354, 8.31814, 9.355413, 9.501351, 7.326774, 4.098248, 4.029028, 
    6.614467, 10.14433, 10.15284, 9.145062, 9.825917, 8.899934, 7.672088, 
    6.020428,
  7.180729, 7.858589, 8.262321, 8.783969, 7.75483, 6.568194, 4.46289, 
    3.620692, 5.405038, 6.067145, 7.953315, 6.877335, 5.138144, 4.553028, 
    4.597962,
  7.092477, 6.553257, 6.954412, 8.028013, 7.528071, 6.568806, 6.288574, 
    4.847325, 3.785006, 4.761351, 4.66331, 5.18966, 3.216179, 3.274454, 
    4.389734,
  6.538945, 6.017395, 6.542206, 7.480423, 7.250793, 6.50151, 6.302023, 
    5.407474, 5.128536, 5.694758, 5.065716, 3.987578, 2.949985, 4.077959, 
    5.235933,
  5.991771, 6.407711, 7.070031, 7.723953, 7.494708, 6.845462, 6.316929, 
    5.400907, 4.552996, 4.438726, 4.038702, 3.466898, 3.225496, 4.288692, 
    4.79916,
  5.381413, 6.362178, 7.367427, 7.923941, 7.50081, 6.759041, 6.51658, 
    5.525671, 4.060938, 3.658225, 3.424579, 3.083719, 3.485289, 4.12358, 
    4.018316,
  4.759393, 6.104749, 7.458272, 8.288696, 8.233918, 7.360497, 6.770483, 
    6.004455, 3.867804, 3.482753, 3.233229, 3.349771, 3.362241, 3.635033, 
    3.099082,
  4.97754, 5.372701, 3.099575, 3.802004, 4.489738, 5.195583, 7.567156, 
    7.399602, 5.28963, 4.298879, 5.276932, 7.665074, 6.493046, 4.04879, 
    2.420708,
  7.631038, 4.996937, 2.834424, 3.59098, 3.373286, 4.983339, 7.767824, 
    8.191584, 6.044715, 5.225369, 5.015223, 8.278605, 9.412121, 5.016244, 
    2.856391,
  8.248001, 4.964729, 2.694964, 3.296103, 3.160893, 4.147873, 7.206414, 
    7.497314, 4.826772, 4.75615, 4.51346, 6.683093, 8.340954, 7.848657, 
    5.369947,
  7.573234, 4.239823, 2.51434, 3.535111, 4.098195, 4.028389, 5.00175, 
    6.608928, 7.003411, 3.773843, 4.675604, 4.241382, 5.67295, 6.525344, 
    5.556519,
  6.374149, 3.214161, 2.700632, 4.26806, 5.613776, 6.391734, 6.427222, 
    5.082153, 5.782652, 3.384846, 5.294734, 2.86115, 3.176065, 4.254694, 
    4.690302,
  4.808226, 2.295161, 2.865, 4.714081, 6.403734, 7.692542, 8.429973, 
    8.873991, 7.979944, 4.228271, 4.622608, 4.094793, 2.568057, 2.860465, 
    3.575516,
  4.235516, 3.046867, 3.362824, 4.585654, 6.420014, 7.820775, 9.439979, 
    10.25758, 11.64391, 7.378737, 6.221971, 5.429905, 3.94698, 3.492823, 
    3.086294,
  4.096029, 3.128742, 3.654599, 5.323676, 6.706697, 7.586792, 8.970536, 
    10.2316, 11.66951, 9.837398, 7.146096, 6.690623, 6.171566, 5.278289, 
    3.838128,
  3.428097, 2.586069, 3.92366, 5.92962, 6.962903, 7.051828, 8.778952, 
    10.47261, 11.78475, 10.04272, 8.100296, 7.686262, 8.059292, 7.02034, 
    5.354798,
  2.576032, 2.800481, 5.039061, 7.055212, 7.865094, 8.051758, 8.481507, 
    9.964593, 10.07739, 6.96226, 6.988136, 9.160413, 8.72201, 8.604092, 
    7.039433,
  6.461444, 5.995696, 2.963517, 4.262152, 4.536984, 4.63354, 6.520946, 
    3.150526, 1.734185, 2.008384, 4.06732, 5.01922, 4.229353, 4.333174, 
    4.080698,
  8.99523, 5.595871, 3.656477, 3.865836, 3.244337, 4.17437, 7.554466, 
    6.580654, 1.714878, 1.108767, 2.596858, 4.758885, 4.641344, 2.983372, 
    2.734708,
  8.894064, 5.476086, 3.856565, 3.259222, 2.81267, 2.78745, 6.058961, 
    7.136121, 3.611036, 1.703856, 1.8589, 3.082912, 3.943363, 3.73033, 
    2.846953,
  7.897395, 4.995766, 3.736276, 3.370725, 2.442301, 2.162895, 3.124631, 
    5.530218, 7.959625, 3.158257, 2.976697, 2.757921, 3.136174, 3.10453, 
    2.870035,
  6.522305, 4.024882, 2.940112, 2.592863, 2.283457, 3.291406, 3.406497, 
    3.411052, 5.28479, 3.858845, 3.608674, 4.013934, 4.235393, 3.56607, 
    3.283715,
  5.231599, 3.16124, 2.261882, 1.930981, 2.571181, 3.868414, 4.7988, 4.7023, 
    5.197456, 5.51382, 3.828821, 4.204152, 5.642905, 5.344779, 4.388505,
  4.32422, 2.922448, 2.175699, 2.272446, 3.804487, 4.970246, 6.009185, 
    5.950684, 6.962451, 7.84767, 7.176057, 4.634639, 5.499825, 6.631464, 
    6.147568,
  4.561878, 4.037528, 3.933532, 4.607664, 5.934269, 6.544913, 6.680161, 
    6.634634, 7.127656, 7.942959, 7.889876, 5.850307, 5.196702, 6.984777, 
    7.363868,
  5.633444, 5.815431, 6.072745, 6.53737, 7.166964, 7.661928, 8.057818, 
    7.937157, 8.068979, 8.305924, 8.138157, 7.29882, 5.676492, 6.613069, 
    7.28002,
  7.001377, 7.120262, 6.877158, 7.946825, 8.7561, 9.249374, 9.165827, 
    8.424098, 7.76005, 6.300441, 6.731203, 8.020354, 6.941205, 6.011815, 
    7.102108,
  8.065275, 8.646607, 5.933161, 5.357009, 3.889817, 2.772856, 3.312241, 
    3.961234, 4.837741, 3.772869, 3.648563, 3.806012, 3.285856, 3.099118, 
    3.201274,
  10.8015, 9.033883, 6.302083, 4.447338, 2.864153, 2.103127, 2.885189, 
    3.791091, 4.829357, 5.420571, 5.216301, 5.813585, 5.649034, 3.85088, 
    3.672226,
  10.42886, 8.46696, 6.364297, 3.978868, 2.636075, 2.077927, 3.666857, 
    5.011136, 5.5253, 6.304181, 7.217472, 7.717963, 8.10497, 8.278874, 
    6.058067,
  8.917574, 7.344297, 6.054513, 5.043814, 4.670925, 4.157118, 3.679348, 
    5.147419, 6.549631, 6.861212, 7.458726, 8.568681, 9.25921, 9.504897, 
    8.438663,
  7.064256, 5.960095, 5.832644, 6.470734, 7.661632, 8.382626, 7.03648, 
    4.924456, 6.157115, 5.886672, 7.950924, 9.601405, 10.13413, 10.55552, 
    10.91035,
  5.683478, 5.638901, 6.889125, 8.323494, 9.776981, 10.72546, 11.18878, 
    10.76433, 9.935609, 8.288198, 8.049425, 11.47964, 11.74066, 11.8857, 
    11.77859,
  5.888927, 6.983333, 8.765258, 10.17808, 11.60277, 12.56751, 13.4185, 
    13.72743, 13.70856, 13.63859, 13.51841, 13.62643, 13.32716, 12.78143, 
    12.6909,
  7.755212, 9.411577, 11.11612, 12.32632, 13.68209, 14.62486, 15.11186, 
    15.3877, 16.06118, 15.73315, 15.82093, 15.21832, 14.51656, 13.63211, 
    12.99297,
  10.70226, 12.26831, 13.59181, 14.53593, 15.22424, 16.10616, 17.05745, 
    17.41052, 17.45589, 15.64286, 15.55822, 15.61883, 15.02923, 13.63632, 
    11.65026,
  13.39646, 14.65394, 15.8561, 16.3577, 17.20862, 17.74561, 18.69611, 
    16.92273, 15.87807, 10.97716, 11.5425, 15.25607, 14.16348, 11.02382, 
    9.505904,
  4.589754, 7.08382, 5.952003, 6.647703, 5.555925, 4.90057, 7.311667, 
    8.610833, 9.344582, 7.667127, 9.15028, 10.51501, 10.26118, 9.541093, 
    9.827024,
  7.633014, 7.913537, 7.207823, 6.096901, 3.830373, 4.069031, 7.352252, 
    8.664817, 11.04484, 10.74454, 10.18261, 12.20675, 13.0843, 9.831044, 
    10.31079,
  8.524915, 8.453454, 7.694353, 6.701498, 4.812936, 3.518308, 6.933348, 
    9.043306, 11.5895, 13.33203, 13.5577, 14.2273, 14.23368, 14.56336, 
    12.73197,
  8.746974, 8.595675, 8.188046, 7.993624, 8.118217, 6.090369, 5.666656, 
    8.324142, 11.97648, 12.24062, 13.87514, 16.04006, 16.02773, 16.28972, 
    14.59611,
  8.793663, 8.431553, 8.325192, 8.615528, 9.688123, 10.59728, 9.368897, 
    8.193244, 11.00892, 10.29006, 15.15225, 17.38431, 17.48172, 18.01437, 
    18.15504,
  8.750056, 8.482159, 8.733485, 9.446156, 10.67778, 12.1433, 13.48311, 
    14.0825, 14.55972, 12.66253, 12.2297, 17.43657, 18.46261, 19.24906, 
    19.29802,
  8.486227, 8.825687, 9.598787, 10.54722, 11.84281, 13.4142, 15.03031, 
    16.8589, 17.78467, 15.68351, 16.04142, 17.70607, 18.83356, 19.46054, 
    20.01875,
  8.183181, 9.175594, 10.39141, 11.55324, 13.04301, 14.61801, 15.50814, 
    15.90091, 15.61952, 15.154, 16.25766, 17.84289, 18.95739, 19.70515, 20.482,
  8.386169, 9.806472, 11.30004, 12.64402, 13.94754, 14.92912, 15.92788, 
    14.83153, 13.59725, 14.61379, 15.70954, 17.61357, 18.69223, 19.64177, 
    19.41017,
  9.425107, 10.81575, 12.53734, 13.79062, 15.14483, 14.79, 13.31916, 12.312, 
    11.09076, 9.819706, 12.07896, 17.52671, 18.77538, 19.72611, 18.56501,
  4.907539, 6.944307, 6.425174, 8.459392, 7.383606, 6.191475, 8.284791, 
    8.061208, 7.860134, 6.2276, 6.497819, 7.202978, 6.5139, 5.725469, 5.596255,
  7.284283, 8.05917, 7.778505, 7.813025, 4.851676, 4.656235, 8.06778, 
    8.01769, 8.732933, 7.99911, 7.618636, 8.896794, 8.17002, 5.791728, 
    5.977933,
  8.16967, 8.787725, 8.691195, 8.8709, 6.434834, 3.651825, 6.38932, 7.962315, 
    9.498778, 10.02045, 9.741449, 9.420407, 8.59265, 8.63098, 7.024489,
  9.032202, 9.450165, 9.741198, 10.17743, 10.94883, 7.93666, 3.636772, 
    4.804811, 7.095157, 8.716683, 9.426886, 9.285622, 8.24012, 8.203367, 
    7.238749,
  9.695542, 9.650736, 9.874179, 10.1305, 10.83536, 11.767, 9.794992, 
    5.335646, 5.335075, 5.629405, 8.265936, 8.681805, 8.548452, 9.156713, 
    9.693992,
  10.03445, 9.906662, 10.03547, 10.12955, 10.45042, 11.25704, 12.50634, 
    13.04246, 10.26301, 8.831516, 7.895225, 10.61472, 11.02504, 11.19607, 
    11.47012,
  9.756432, 9.752199, 9.928717, 10.01798, 10.40428, 10.86546, 11.73826, 
    12.83747, 13.23845, 13.29863, 12.56344, 11.96219, 11.52672, 11.44749, 
    11.53214,
  8.760397, 8.936779, 9.338573, 9.758771, 10.43108, 11.06172, 11.6159, 
    12.17061, 12.61485, 12.53203, 12.59248, 11.828, 11.69479, 11.51533, 
    11.75812,
  8.04698, 8.006783, 8.317191, 8.549935, 9.252556, 10.074, 11.25757, 
    12.27521, 12.36997, 12.58703, 12.82486, 12.30455, 11.73081, 11.6769, 
    11.39631,
  7.328394, 6.654385, 6.442967, 6.752027, 7.659811, 9.253445, 10.95024, 
    11.63048, 11.00762, 8.800835, 9.969233, 12.59687, 12.28914, 12.06994, 
    11.4049,
  5.632582, 8.013103, 7.070198, 9.111292, 8.102086, 6.310418, 8.084504, 
    7.28156, 6.043377, 4.397289, 4.484409, 5.106802, 4.487449, 4.345492, 
    5.137443,
  8.116549, 8.807858, 8.867144, 9.215082, 5.750497, 4.862683, 7.093439, 
    6.203499, 6.059912, 5.663074, 5.413603, 6.895892, 6.928577, 5.188092, 
    5.719394,
  9.644295, 9.295216, 8.913316, 8.783309, 6.000756, 3.928626, 5.385315, 
    5.49767, 6.077214, 6.764528, 7.287745, 8.040941, 8.477276, 8.783764, 
    6.674435,
  9.657825, 9.454304, 9.464175, 9.277369, 7.961195, 5.725778, 3.380029, 
    3.642488, 5.15096, 6.280447, 6.6518, 6.9691, 6.840179, 6.952892, 6.342839,
  8.97808, 9.258945, 9.363728, 9.035834, 8.55458, 7.697242, 6.486232, 
    3.465809, 3.790431, 4.352829, 5.289487, 5.694154, 6.619588, 7.225214, 
    7.493439,
  9.012897, 9.505297, 9.199256, 8.495121, 7.773428, 6.970999, 7.233263, 
    7.491719, 5.62365, 4.631305, 4.235062, 7.079431, 7.928417, 8.005767, 
    9.032051,
  10.05647, 9.791106, 8.830452, 7.459492, 6.632951, 5.809059, 6.125558, 
    6.498305, 5.710815, 5.480597, 6.518417, 7.537048, 7.490439, 8.235303, 
    9.575067,
  10.43816, 9.096024, 7.564416, 6.442621, 5.630524, 5.399734, 5.292477, 
    4.844778, 4.320035, 5.978598, 6.961492, 6.693306, 7.361582, 8.665261, 
    10.05957,
  9.536826, 8.136032, 6.661068, 5.089463, 4.367864, 4.312202, 4.639758, 
    4.170678, 5.391892, 6.303363, 6.734145, 6.825578, 7.80101, 9.214664, 
    10.24604,
  7.905557, 6.456662, 5.172566, 4.064262, 3.847535, 4.497144, 4.121133, 
    5.08877, 5.565697, 4.598684, 5.642163, 6.910814, 7.740183, 9.324182, 
    9.993925,
  3.966881, 5.757541, 5.624527, 8.527819, 8.726269, 7.955436, 10.16301, 
    10.20953, 8.279534, 4.703174, 4.332859, 4.392266, 3.763209, 3.517688, 
    3.985496,
  5.444806, 6.126239, 7.022631, 8.609432, 6.617291, 6.614872, 9.994211, 
    9.837117, 8.58295, 5.966787, 5.022641, 5.526935, 5.498663, 4.063727, 
    4.250309,
  6.641526, 6.713795, 7.447269, 9.197515, 7.108441, 6.310119, 8.286802, 
    8.665269, 7.744537, 6.86899, 6.358835, 6.114986, 6.499959, 7.104738, 
    5.803327,
  7.390232, 7.638204, 8.787926, 9.758463, 9.904513, 7.081066, 6.503247, 
    6.878013, 6.988294, 6.407273, 6.207407, 6.298368, 6.600472, 7.253205, 
    6.423577,
  7.566547, 7.900764, 8.981761, 9.690468, 10.07508, 9.414853, 7.251514, 
    5.502158, 6.057775, 5.585142, 6.450126, 7.227382, 7.56303, 7.634594, 
    7.172334,
  8.03075, 8.751756, 9.186185, 9.325825, 9.599879, 9.797177, 9.161345, 
    8.380027, 7.241158, 6.247975, 5.580977, 8.179564, 8.405831, 7.589909, 
    7.31732,
  8.786489, 8.996142, 9.077247, 9.062965, 9.477909, 9.775964, 10.12078, 
    10.10261, 8.946314, 8.316951, 8.028964, 8.737837, 7.282291, 7.039179, 
    7.339139,
  9.298402, 9.189827, 9.211653, 9.375534, 9.874307, 10.49462, 10.64458, 
    10.43954, 9.500745, 9.395203, 9.28778, 6.760854, 6.883211, 7.296303, 
    6.280485,
  9.256129, 9.600507, 9.926404, 10.08833, 10.71813, 10.93428, 11.37983, 
    11.06881, 10.47432, 9.774623, 7.130588, 7.445878, 7.428695, 6.047299, 
    6.166179,
  9.41323, 9.954017, 10.62161, 11.30707, 11.88957, 12.16035, 11.99688, 
    11.35092, 9.232738, 5.009841, 6.455523, 8.129824, 5.938131, 5.422133, 
    5.836925,
  4.775323, 6.93188, 5.784063, 7.721228, 7.35574, 6.336759, 9.493462, 
    10.87782, 9.768135, 7.393202, 7.505285, 8.159516, 7.537706, 7.38461, 
    7.503653,
  7.463597, 8.093822, 7.576242, 7.893085, 5.269836, 6.109254, 9.791971, 
    10.70368, 11.53484, 10.08314, 8.549201, 9.645884, 9.991165, 7.840322, 
    8.096815,
  10.14068, 10.06385, 9.341694, 9.168849, 6.510934, 5.788563, 9.642544, 
    10.00339, 10.455, 10.72887, 10.95689, 11.75162, 12.52257, 12.37758, 
    10.06725,
  11.8344, 11.58417, 11.25619, 10.55121, 9.486598, 7.851147, 7.283763, 
    8.892419, 11.00501, 10.60543, 11.64806, 13.61481, 14.23229, 13.40781, 
    9.933846,
  13.06832, 12.51322, 11.87846, 11.35872, 11.24359, 11.01668, 9.330772, 
    7.611208, 9.430731, 9.815365, 13.60762, 15.49498, 15.35206, 13.23065, 
    10.83526,
  13.38029, 12.66196, 11.8567, 11.38459, 11.52344, 11.64766, 11.6597, 
    12.34801, 11.60343, 11.58106, 11.58005, 15.58658, 15.12705, 12.29594, 
    9.953204,
  11.89587, 11.64167, 11.44814, 11.16613, 11.74809, 11.85046, 12.57042, 
    13.56988, 14.7378, 15.13478, 14.98195, 15.51466, 13.27136, 9.871435, 
    7.589566,
  11.12915, 11.43394, 11.55765, 11.64102, 11.88998, 12.44739, 12.97803, 
    13.45803, 14.41286, 14.92225, 14.99733, 14.19674, 9.968064, 7.120341, 
    5.459701,
  12.20708, 12.29741, 12.2916, 11.6102, 12.15119, 12.53138, 13.27058, 
    13.70231, 13.79541, 13.71918, 13.71213, 11.4124, 6.650217, 5.860879, 
    5.192508,
  12.90528, 12.55723, 12.596, 12.44257, 12.40148, 13.10829, 13.57481, 
    13.03213, 10.97064, 8.915184, 9.265345, 6.991678, 6.199343, 5.365197, 
    3.649051,
  7.341906, 10.49476, 8.892182, 10.7143, 9.485789, 7.753011, 11.01424, 
    12.17919, 12.41286, 9.20507, 9.081838, 9.834546, 9.039924, 8.399747, 
    7.876414,
  11.5803, 12.76347, 11.49442, 10.86124, 7.038514, 7.086524, 11.20128, 
    11.89894, 12.74125, 11.23498, 9.684829, 11.342, 10.13175, 7.53705, 
    7.593989,
  13.80291, 14.64935, 14.25878, 12.70125, 9.43778, 7.10761, 10.64758, 
    11.15339, 11.38459, 11.58669, 11.17493, 11.03386, 10.27872, 10.15384, 
    8.816453,
  15.01682, 15.1584, 14.90321, 14.32632, 12.9609, 9.380743, 7.508859, 
    9.401525, 9.64398, 9.053165, 10.05169, 10.97336, 11.13041, 11.51748, 
    8.863223,
  16.13871, 15.70477, 15.05437, 14.34807, 13.63943, 12.41833, 10.36436, 
    7.117217, 7.273443, 6.803825, 9.723221, 11.35951, 11.4981, 11.50883, 
    9.572118,
  15.83627, 15.1221, 14.36612, 13.63805, 12.96855, 12.2749, 11.96371, 
    12.06271, 9.776066, 8.669621, 8.554097, 11.74091, 11.86138, 11.31951, 
    8.111616,
  13.47161, 13.12642, 12.77562, 12.09644, 11.88077, 11.5934, 11.74674, 
    11.66906, 11.95294, 12.04257, 11.83022, 11.90035, 11.53766, 9.93153, 
    6.706125,
  12.42001, 12.37835, 12.33983, 11.89201, 11.7882, 11.93957, 11.68039, 
    11.55552, 11.96778, 12.04927, 12.04346, 11.70715, 11.0304, 8.447457, 
    7.746727,
  14.54957, 14.30994, 14.06657, 13.26523, 13.27674, 12.50485, 12.85668, 
    12.76877, 12.4495, 11.8119, 11.46576, 11.30999, 10.28031, 8.607561, 
    7.818399,
  16.79136, 16.36722, 15.9435, 14.78991, 14.39614, 13.97718, 13.97504, 
    13.49794, 10.76876, 8.643887, 8.777, 10.73292, 9.424251, 9.478948, 
    7.419141,
  8.663574, 12.04714, 10.27772, 13.57296, 12.70426, 9.898085, 12.38502, 
    12.12765, 11.65235, 9.09772, 8.856795, 9.149226, 8.465245, 7.724981, 
    7.526527,
  13.36772, 15.10272, 13.40902, 13.55432, 9.14475, 8.511754, 14.54745, 
    13.89457, 13.42849, 11.86622, 9.889562, 11.17946, 11.40621, 8.055403, 
    7.696053,
  15.30925, 16.36048, 15.97681, 14.87396, 11.23856, 8.43725, 12.3991, 
    12.86554, 12.77742, 12.49117, 11.68031, 11.47792, 11.39529, 10.80559, 
    8.664862,
  16.09891, 16.8919, 16.94312, 16.76452, 15.97914, 11.20575, 8.086926, 
    9.448102, 11.38651, 11.47369, 11.76913, 10.89407, 9.756338, 9.643085, 
    8.04821,
  16.57775, 16.8897, 16.80466, 16.35005, 15.90426, 14.8998, 12.46563, 
    7.889956, 7.235853, 6.654891, 9.846677, 9.818428, 8.697864, 8.889918, 
    8.888384,
  15.55007, 15.7209, 15.7103, 15.46084, 14.92861, 14.31325, 14.06364, 
    14.02854, 9.967444, 7.365764, 6.999464, 9.316428, 9.016885, 9.440075, 
    9.953072,
  12.74086, 12.99337, 13.19962, 13.2697, 13.3265, 13.09557, 12.96424, 
    12.74356, 12.19037, 10.76665, 10.33911, 10.11157, 10.05489, 9.939396, 
    9.867867,
  11.22703, 11.63509, 12.03704, 11.97801, 12.08656, 12.39666, 12.2804, 
    11.95751, 11.73994, 10.68386, 10.49429, 10.18372, 9.915276, 9.686652, 
    9.763459,
  10.75965, 11.16269, 11.48836, 11.37791, 11.39563, 11.43497, 12.1767, 
    12.6884, 12.01979, 10.68419, 10.79193, 10.4448, 10.27741, 10.4497, 9.71771,
  8.830853, 9.364546, 9.805141, 9.711924, 9.617078, 9.724428, 9.806045, 
    9.849158, 9.303368, 8.324406, 8.720638, 11.07602, 10.57308, 10.11204, 
    9.336377,
  7.994765, 11.33155, 9.236082, 12.216, 10.30365, 9.083072, 11.70503, 
    10.99381, 10.43845, 8.678534, 8.428713, 8.997336, 7.769568, 6.69565, 
    6.534934,
  11.87981, 13.54423, 12.65143, 11.88999, 7.414193, 7.639849, 13.22342, 
    11.87672, 11.77137, 11.22798, 9.871661, 11.03488, 10.62575, 7.288893, 
    7.004771,
  11.77174, 13.78466, 14.20521, 14.10404, 9.339788, 7.26328, 11.76514, 
    12.89533, 12.93035, 11.83277, 12.70317, 12.93871, 12.01396, 11.23957, 
    8.552814,
  10.22183, 12.37981, 14.06613, 14.83362, 14.50087, 11.35233, 6.892925, 
    8.75951, 11.228, 12.62028, 13.0998, 13.08751, 12.74861, 11.78372, 9.522237,
  7.057811, 7.770425, 9.691849, 11.69031, 13.18303, 14.97981, 13.01854, 
    8.127806, 7.705493, 7.390484, 11.09801, 11.86355, 10.76197, 9.90717, 
    9.654879,
  5.371058, 4.406931, 4.479873, 5.108244, 6.29831, 8.344103, 11.40439, 
    14.15012, 9.928927, 7.251176, 7.202673, 10.34983, 9.927858, 9.45672, 
    9.342295,
  5.732053, 4.911368, 4.686472, 4.806464, 5.578444, 6.540004, 8.14242, 
    9.950212, 10.73959, 9.54291, 9.72089, 10.10792, 9.940026, 9.718131, 
    9.703918,
  7.359737, 6.670643, 6.33172, 6.441312, 7.07798, 7.532363, 7.475904, 
    7.445293, 8.244545, 7.511616, 8.578312, 9.09361, 9.357041, 9.342032, 
    9.458412,
  8.441084, 8.039426, 7.337409, 6.687409, 6.372502, 5.928829, 5.545047, 
    6.251218, 7.539355, 8.291124, 9.711678, 9.667569, 9.758489, 9.520528, 
    9.104902,
  8.716559, 8.611614, 8.130584, 7.246423, 6.252102, 5.309008, 5.548575, 
    6.036343, 5.791883, 5.529872, 6.149316, 6.439639, 5.332125, 4.580302, 
    4.15126,
  7.926132, 11.53982, 9.966699, 13.00688, 10.85432, 9.50803, 13.50087, 
    12.19413, 11.65613, 8.943577, 8.238787, 9.082815, 7.56053, 6.686445, 
    6.545029,
  11.24237, 13.75457, 13.79372, 13.2685, 7.578278, 8.302008, 14.07668, 
    13.83216, 12.79304, 11.82152, 10.32747, 12.24644, 11.45861, 7.775909, 
    7.078757,
  9.178668, 11.9137, 13.97236, 15.26425, 10.53859, 7.846483, 11.70148, 
    13.14493, 12.98818, 12.20791, 13.14618, 13.32776, 12.9176, 12.10754, 
    8.939709,
  5.808053, 5.919355, 7.481746, 10.12245, 13.36023, 11.47319, 6.728641, 
    7.882558, 10.74176, 11.69564, 12.52108, 13.53196, 12.91938, 12.69916, 
    10.16552,
  4.38201, 3.772671, 4.030073, 4.890412, 6.351172, 11.0052, 11.20362, 
    6.296522, 5.908024, 6.745683, 9.381012, 10.5516, 10.44345, 10.76547, 
    11.10524,
  5.376784, 4.224195, 4.186141, 4.550744, 5.127196, 4.239688, 7.920691, 
    10.55273, 6.844709, 4.256399, 4.911076, 7.425514, 7.977898, 8.701768, 
    9.520775,
  6.234181, 5.285413, 4.343836, 4.151442, 4.419007, 5.003121, 4.217373, 
    4.533627, 4.297369, 3.561443, 4.125385, 4.829304, 5.065878, 5.622617, 
    6.526359,
  6.441652, 6.279205, 5.43468, 4.740715, 4.378609, 4.152784, 3.762094, 
    3.165291, 3.050644, 2.826123, 3.706691, 4.03187, 4.732415, 5.65955, 
    6.566969,
  5.870571, 6.20538, 5.806958, 5.34035, 5.296319, 5.123976, 4.843025, 
    4.932444, 4.839251, 5.189277, 6.347566, 5.120063, 5.821865, 6.908258, 
    8.320672,
  5.207568, 6.121751, 6.142336, 5.774269, 6.035481, 5.858891, 5.007393, 
    4.475603, 4.112211, 3.846956, 4.389255, 4.655527, 4.474283, 4.76727, 
    4.938929,
  6.918136, 10.02486, 8.489274, 10.46282, 8.320137, 7.826704, 10.89137, 
    10.85588, 10.36577, 8.24132, 8.709214, 9.840137, 8.978568, 7.837048, 
    7.91839,
  9.420902, 11.70944, 11.84859, 11.28796, 5.980603, 7.051376, 11.33163, 
    11.58043, 11.36178, 10.61195, 10.16879, 12.48136, 12.52858, 8.361846, 
    7.828475,
  8.591183, 9.906183, 11.53893, 13.06239, 9.169972, 6.882656, 10.17841, 
    11.60633, 12.13202, 12.31451, 13.60725, 14.08297, 14.03851, 13.79228, 
    9.384964,
  7.20944, 6.440169, 7.06363, 8.467301, 10.91241, 10.08443, 6.052303, 
    7.076087, 9.593836, 11.15609, 13.43975, 14.8776, 14.85104, 14.81966, 
    11.53715,
  5.552757, 4.533463, 4.406484, 4.621559, 5.247386, 8.23674, 8.853203, 
    5.542877, 5.686531, 7.008614, 10.60432, 12.54752, 13.32349, 13.47293, 
    14.01616,
  5.423586, 4.495244, 3.780025, 3.327708, 3.072092, 3.68924, 5.687346, 
    7.786209, 5.112791, 3.789542, 4.962769, 7.979461, 8.929288, 10.38687, 
    11.57547,
  5.993237, 5.262032, 4.595596, 4.436851, 4.181571, 4.139256, 4.340569, 
    4.531144, 3.754132, 2.20206, 2.478877, 3.773983, 5.011126, 6.031296, 
    6.724302,
  7.311162, 6.944034, 6.441803, 6.6978, 6.535512, 6.187756, 5.519081, 
    5.111628, 4.492574, 3.371371, 2.671863, 2.171845, 2.753861, 3.437135, 
    3.941323,
  8.22169, 8.014817, 7.533977, 7.699752, 7.269883, 6.809836, 6.167861, 
    5.502224, 4.553516, 3.979915, 3.509241, 1.777504, 2.055371, 2.600999, 
    3.169652,
  7.498715, 7.726908, 7.603349, 7.616731, 7.374992, 6.818921, 6.285107, 
    5.620216, 4.645057, 3.784507, 3.213393, 2.069803, 1.398749, 1.498108, 
    2.529433,
  7.006031, 10.24924, 8.92412, 10.6759, 8.390185, 7.452877, 10.03468, 
    9.057471, 8.533552, 6.06228, 6.639796, 7.776071, 7.299487, 6.63395, 
    7.167916,
  8.599765, 10.83796, 11.8746, 11.75425, 7.188746, 7.377628, 11.05442, 
    10.25516, 9.519897, 8.169953, 7.944502, 9.642612, 9.908898, 6.699843, 
    6.726335,
  7.174895, 8.071877, 10.44559, 12.86479, 10.19774, 7.2323, 9.886349, 
    11.36304, 11.4353, 9.866199, 10.85051, 10.77131, 10.58875, 10.52299, 
    7.586085,
  5.685074, 5.449182, 6.810699, 7.525985, 12.59769, 11.36321, 6.451606, 
    7.359145, 10.54559, 11.43935, 12.39793, 12.35731, 11.10741, 10.8601, 
    9.411854,
  5.36727, 5.914389, 6.486267, 7.365334, 5.545304, 9.761511, 10.23814, 
    6.452518, 6.926855, 8.40978, 12.32577, 13.3127, 12.48339, 12.0299, 
    12.13444,
  5.815313, 6.314986, 6.371386, 7.371893, 8.684986, 5.869844, 5.039331, 
    7.547489, 4.800012, 4.187159, 6.836758, 10.80788, 11.50053, 11.60747, 
    11.66542,
  5.498315, 5.619778, 5.174541, 6.012064, 7.351456, 9.090627, 8.813745, 
    6.479463, 4.234925, 2.86841, 4.47894, 6.773468, 8.399676, 9.389131, 
    10.35398,
  5.129647, 4.214808, 3.386335, 3.812048, 4.490149, 5.295952, 6.003269, 
    6.812887, 7.254392, 6.086573, 3.239693, 3.023862, 3.908889, 5.226842, 
    6.7613,
  5.603343, 3.728987, 2.730119, 2.863148, 3.387181, 4.020356, 4.018888, 
    3.649492, 3.245123, 3.4232, 3.576055, 4.081785, 3.22915, 2.636678, 
    3.155168,
  7.543195, 4.846857, 3.586866, 3.015412, 3.34138, 3.792654, 3.775384, 
    3.142384, 2.389662, 2.369592, 2.086066, 2.319512, 2.630766, 2.456403, 
    1.586817,
  8.41614, 10.80358, 8.690897, 10.70745, 8.582168, 8.060695, 10.63265, 
    9.849052, 9.020896, 6.230458, 5.932719, 6.745738, 6.013844, 5.384382, 
    5.421659,
  11.83375, 11.98555, 10.66483, 10.31169, 5.951675, 6.819415, 10.69208, 
    10.23846, 9.967419, 8.705914, 7.479095, 8.752672, 9.060072, 5.988956, 
    5.845898,
  9.844406, 10.18568, 8.691715, 8.021039, 6.622321, 5.406794, 8.374403, 
    9.852211, 10.04634, 10.05829, 10.42241, 9.811371, 9.467305, 9.162641, 
    6.780938,
  7.469975, 7.414132, 5.446503, 4.41408, 6.518598, 6.361928, 3.9101, 
    5.447662, 7.600817, 10.10319, 11.34346, 10.35735, 9.428762, 9.027519, 
    8.072526,
  9.794755, 9.223598, 5.974895, 3.917845, 3.049935, 4.775267, 5.233277, 
    2.796766, 3.279208, 4.666019, 9.556993, 10.95734, 10.32213, 9.898237, 
    10.19241,
  12.7021, 10.83592, 6.41649, 3.56427, 4.307945, 4.240978, 4.104814, 
    4.587831, 2.967997, 2.904171, 3.627338, 8.060287, 9.790917, 9.790559, 
    9.722826,
  13.3927, 10.52332, 6.167932, 3.077475, 3.339198, 5.597589, 7.288008, 
    7.506471, 6.197301, 5.369491, 4.679679, 5.912416, 8.200921, 9.704959, 
    10.02542,
  12.27549, 8.695733, 4.086173, 3.881066, 4.249318, 4.940921, 5.581526, 
    4.85133, 3.718749, 4.019516, 5.135986, 4.595884, 7.069961, 9.211696, 
    9.72423,
  12.50381, 9.821888, 6.987216, 5.634136, 5.221043, 4.514585, 3.853451, 
    3.077951, 2.219937, 2.780174, 4.969094, 5.995456, 4.413427, 8.127573, 
    8.975019,
  12.84492, 10.72856, 9.350798, 9.352737, 9.376216, 7.334558, 4.821069, 
    2.275774, 1.162336, 1.914391, 3.737747, 6.225011, 5.198403, 6.068448, 
    8.340454,
  6.125191, 9.243629, 8.252221, 11.70309, 10.94531, 9.284458, 11.30307, 
    9.332506, 8.878311, 6.189525, 5.718972, 5.890442, 4.620955, 3.926888, 
    3.609342,
  7.246834, 9.011479, 9.038326, 9.213657, 6.68137, 7.551662, 11.02849, 
    9.94908, 9.673506, 8.639371, 7.167788, 8.121687, 7.966005, 4.727671, 
    3.957521,
  7.166672, 8.826312, 9.248557, 8.594337, 7.045533, 5.294721, 8.566237, 
    10.35103, 9.817625, 9.387334, 9.841292, 9.484324, 9.449425, 8.373607, 
    5.882167,
  6.964635, 8.170289, 8.991039, 9.472919, 9.911841, 6.781621, 3.855163, 
    6.031063, 8.344953, 9.974833, 10.42072, 9.466505, 9.357623, 8.972085, 
    7.489356,
  8.141449, 10.11059, 9.946653, 8.874425, 8.092104, 8.625385, 6.893522, 
    4.600459, 5.010869, 6.192439, 9.594114, 10.02908, 9.61557, 9.972809, 
    10.30792,
  13.22034, 12.38782, 10.53089, 7.983847, 5.072946, 4.506749, 7.306881, 
    8.870315, 5.666564, 4.595253, 4.915902, 7.18577, 8.422196, 9.164972, 
    9.427046,
  14.44245, 12.97699, 10.90955, 7.711246, 5.030205, 4.227388, 5.558386, 
    8.249209, 8.104679, 7.411481, 6.39844, 5.622386, 4.73445, 5.523359, 
    7.178075,
  16.02467, 14.24608, 12.24198, 9.918852, 8.876146, 8.263943, 9.308054, 
    10.6902, 11.06146, 8.681739, 6.119808, 4.961356, 4.808645, 3.97346, 
    4.012646,
  17.06454, 14.88157, 12.39638, 10.42016, 10.15723, 10.98689, 8.268681, 
    9.526078, 10.92635, 9.097545, 6.631729, 4.949448, 4.548931, 4.146641, 
    3.383058,
  14.16861, 12.2336, 10.50686, 9.414855, 9.323755, 10.88393, 12.68971, 
    10.5422, 7.20204, 5.372768, 4.736567, 4.993361, 4.938401, 5.009414, 
    4.318545,
  3.124835, 5.009633, 4.898648, 7.813118, 7.784956, 7.741634, 10.64822, 
    10.55241, 9.869846, 6.63827, 5.496022, 5.530376, 4.231553, 3.363661, 
    3.831719,
  5.025331, 5.033085, 5.486198, 6.386228, 4.804728, 5.853378, 9.461428, 
    10.21963, 9.996264, 8.430034, 6.392724, 7.042452, 6.088778, 3.260238, 
    3.052416,
  4.813605, 6.057136, 6.422193, 6.740529, 5.750445, 4.71711, 6.918292, 
    9.221786, 10.26856, 9.966555, 8.945482, 7.957417, 6.432559, 4.842874, 
    3.058125,
  2.797315, 3.197209, 5.588875, 6.784421, 7.549508, 5.575066, 4.515642, 
    6.010225, 7.913672, 9.253654, 8.977026, 7.966863, 6.327118, 4.78518, 
    3.374217,
  7.769537, 8.899569, 8.053387, 7.200591, 6.205252, 6.505454, 6.365842, 
    4.847955, 4.623837, 6.045368, 8.609871, 8.072249, 6.8497, 5.654285, 
    4.121358,
  12.03768, 11.42532, 10.4558, 9.442932, 7.987475, 6.135656, 5.809166, 
    7.230727, 5.724924, 5.675894, 6.360046, 8.340475, 7.634799, 6.382027, 
    4.73167,
  12.55409, 12.36794, 11.85874, 11.44026, 10.2458, 8.708429, 5.94775, 
    3.723347, 4.812312, 8.586658, 9.432415, 8.867268, 8.133629, 7.241541, 
    5.867773,
  11.67158, 11.83834, 11.46947, 11.27478, 10.24597, 9.137996, 7.955299, 
    6.611323, 5.03154, 4.366658, 8.784206, 9.48259, 8.623542, 7.779967, 
    6.674906,
  9.733024, 9.656174, 9.369434, 8.991346, 8.308368, 7.599203, 7.092296, 
    7.095933, 6.162048, 4.862097, 6.524266, 9.261983, 9.127145, 8.250257, 
    6.830996,
  8.152355, 8.019052, 7.686921, 7.025869, 6.57982, 6.621836, 6.862376, 
    7.10763, 5.544075, 4.115241, 5.56547, 8.929018, 9.186124, 8.688392, 
    7.290181,
  2.753623, 4.602363, 4.707425, 6.618659, 6.404032, 6.146551, 8.755889, 
    9.30365, 9.039429, 7.101398, 7.444187, 8.775519, 8.383475, 7.413267, 
    6.672776,
  5.650109, 5.839239, 5.35974, 5.871241, 4.426733, 5.567955, 8.492505, 
    9.071499, 9.358581, 8.968619, 8.363191, 11.2477, 11.69753, 7.323828, 
    6.242078,
  4.472658, 6.661644, 7.321323, 6.839839, 5.119354, 4.179793, 6.858679, 
    8.964841, 10.07041, 10.51914, 11.10788, 11.53487, 12.07874, 10.65066, 
    7.459824,
  4.635715, 2.532458, 4.270802, 7.841187, 8.543081, 6.021083, 3.702208, 
    5.264395, 7.999933, 10.33012, 10.8878, 11.0138, 10.71832, 9.896152, 
    7.924004,
  10.99875, 10.39365, 7.345465, 3.280034, 7.125709, 9.000741, 6.899289, 
    4.96115, 5.274234, 6.496629, 10.33381, 10.69294, 10.3261, 9.868205, 
    8.779789,
  10.57602, 12.00061, 13.00896, 10.99362, 7.014787, 5.735965, 7.522892, 
    8.452374, 6.216481, 6.34679, 7.740251, 10.88361, 10.40728, 9.399941, 
    7.919319,
  8.648606, 9.614352, 11.3322, 13.12145, 13.61526, 11.7295, 7.367898, 
    5.819263, 7.141265, 9.441898, 10.95653, 10.96432, 10.71584, 9.558194, 
    7.911439,
  7.068779, 7.412221, 8.355783, 9.797224, 10.9417, 11.72305, 11.42307, 
    8.661677, 5.743363, 7.245043, 9.919738, 10.93092, 10.76229, 9.727194, 
    8.39765,
  6.652332, 6.876401, 7.609805, 8.378008, 8.794291, 9.041407, 9.422804, 
    9.648304, 7.433936, 5.504736, 7.951591, 10.55326, 10.59713, 10.0869, 
    8.310847,
  7.75372, 6.885871, 7.012293, 6.712972, 6.667916, 6.967369, 7.215663, 
    7.315251, 6.380817, 4.308013, 4.88621, 9.197021, 10.2743, 10.02819, 
    8.386638,
  2.046262, 1.935232, 1.613695, 3.056677, 3.338199, 3.163897, 4.314057, 
    4.875574, 7.818687, 7.356246, 8.074167, 10.23819, 10.01199, 8.804729, 
    7.703516,
  4.282676, 3.258535, 1.770269, 2.706413, 2.791684, 3.918282, 5.411696, 
    5.596682, 7.418353, 9.244013, 9.171255, 12.52084, 13.10673, 8.613863, 
    7.875501,
  7.646522, 3.830935, 4.847346, 2.840457, 3.038169, 2.989741, 5.536727, 
    6.610081, 8.537676, 10.18043, 11.47501, 12.3732, 12.81522, 12.27248, 
    9.928728,
  11.8749, 6.825361, 4.051771, 5.97823, 4.620021, 3.815391, 3.526927, 
    6.241296, 7.881002, 8.401297, 10.56906, 11.84482, 12.52564, 12.33458, 
    10.61964,
  11.08436, 12.65411, 6.666608, 4.689046, 7.280972, 6.150502, 5.568507, 
    4.586266, 4.657198, 5.662213, 9.924659, 11.79759, 12.46183, 12.19841, 
    11.53347,
  8.090278, 10.99609, 13.06784, 7.078585, 6.113657, 7.887335, 7.460114, 
    7.767378, 6.291453, 6.558193, 7.841592, 11.73588, 11.8552, 10.84852, 
    9.819549,
  7.038412, 8.538788, 11.79374, 12.42898, 7.934934, 7.156164, 6.625026, 
    7.80589, 8.59823, 9.724263, 10.86956, 11.44114, 11.06097, 10.7276, 
    10.06377,
  6.896848, 7.439422, 9.395768, 11.38433, 11.3498, 9.577136, 7.829947, 
    6.238678, 8.683788, 9.641728, 10.06818, 10.94841, 10.82444, 10.40881, 
    10.39563,
  8.52721, 8.200041, 8.565865, 9.670375, 10.73642, 10.75487, 9.150397, 
    6.755408, 5.059507, 8.405321, 9.490151, 10.35012, 10.46752, 10.50189, 
    10.05719,
  8.7249, 8.350951, 7.923244, 7.958899, 8.314026, 8.899194, 8.5003, 6.707024, 
    3.821482, 4.889319, 7.062862, 9.966773, 10.30786, 10.98728, 9.787642,
  5.430339, 5.667033, 4.542571, 7.455359, 8.110503, 6.896481, 8.629191, 
    8.36188, 9.251388, 7.115257, 7.088131, 7.473067, 6.406602, 5.470098, 
    4.811154,
  9.856898, 6.175679, 5.517942, 6.449395, 3.94778, 2.767044, 3.457728, 
    5.488703, 7.862203, 8.920415, 7.804753, 9.848071, 9.761844, 5.435277, 
    4.703709,
  12.45741, 9.679731, 5.795285, 4.438346, 3.61749, 2.505532, 4.071552, 
    5.647927, 8.127137, 9.537881, 9.818081, 9.323881, 9.25399, 8.608319, 
    6.504304,
  12.37016, 12.24374, 8.801517, 6.293118, 5.143125, 4.10913, 3.680037, 
    6.028337, 7.182637, 7.301754, 8.490506, 8.574835, 8.345718, 8.716149, 
    8.104975,
  11.63299, 12.68005, 10.79872, 7.838345, 6.8672, 5.863629, 6.193138, 
    4.937071, 4.588082, 4.679272, 7.535711, 8.447741, 8.777122, 9.406423, 
    9.57737,
  11.20863, 12.88227, 12.47861, 9.645444, 7.680282, 7.108093, 6.196747, 
    6.940438, 6.301047, 6.587919, 6.618929, 9.059555, 9.202303, 8.843834, 
    8.848527,
  10.79904, 12.84641, 13.59628, 12.03315, 9.313472, 8.464104, 8.011597, 
    7.664349, 8.183096, 9.599447, 10.15356, 10.34337, 10.14636, 9.979152, 
    10.61456,
  10.80433, 12.59138, 13.70135, 13.69187, 11.73235, 9.803362, 9.106781, 
    9.261095, 9.379016, 10.04533, 11.11642, 11.66286, 12.38678, 12.40338, 
    12.24391,
  11.14369, 12.60471, 13.4639, 13.7451, 12.86369, 11.08553, 9.937767, 
    9.930904, 9.993778, 10.71029, 11.98598, 13.21297, 13.67093, 13.13074, 
    11.51605,
  10.14607, 11.4706, 12.65016, 13.16134, 12.69377, 11.14238, 9.868936, 
    9.947495, 8.917809, 7.649108, 9.693225, 13.34825, 12.85854, 11.90249, 
    10.71062,
  6.77118, 8.041276, 4.689914, 4.09279, 3.188748, 7.384395, 13.46854, 
    13.25512, 10.82323, 7.021139, 6.722671, 7.392819, 6.624201, 5.689495, 
    4.561367,
  9.561997, 6.718038, 4.978483, 3.685384, 3.35315, 3.554666, 12.64255, 
    14.31952, 11.56209, 9.654725, 7.758338, 9.265641, 9.194431, 5.245401, 
    4.289484,
  10.04604, 7.026825, 4.486609, 3.586159, 3.867593, 4.477468, 9.262283, 
    12.81619, 12.09043, 10.83935, 9.634307, 8.952485, 8.548989, 7.612966, 
    5.714382,
  11.34038, 9.239757, 7.797303, 7.311958, 7.524203, 8.509294, 8.458971, 
    8.766582, 9.364092, 8.561193, 8.471504, 7.755666, 7.182194, 7.241573, 
    6.561892,
  12.33867, 11.02152, 9.923008, 9.833643, 10.49343, 11.80503, 11.5408, 
    8.143855, 5.633473, 4.813231, 7.280922, 7.265155, 6.921313, 6.862079, 
    7.015183,
  12.97737, 12.08481, 11.15347, 10.75266, 11.38174, 11.68812, 11.29314, 
    10.84297, 7.778862, 6.779126, 5.705063, 7.019043, 6.347729, 5.661335, 
    5.187773,
  13.47257, 12.81489, 11.98616, 11.28646, 11.37773, 11.73614, 11.19413, 
    10.08091, 9.282883, 8.983205, 7.73091, 6.550955, 5.533137, 4.390108, 
    4.041677,
  13.83633, 13.21997, 12.52316, 11.90211, 11.18851, 11.10629, 10.8977, 
    10.35418, 8.54961, 7.37377, 6.427352, 5.198428, 4.571035, 4.881497, 
    5.403453,
  13.54289, 13.15103, 12.49966, 11.81767, 10.67932, 10.10196, 9.614981, 
    8.764876, 7.317331, 5.890547, 5.177976, 5.446314, 5.999284, 6.347046, 
    6.019304,
  11.96201, 12.04261, 11.62898, 10.86778, 9.302081, 8.139674, 7.63348, 
    7.644833, 5.674323, 4.182939, 4.702157, 7.015374, 7.577833, 7.385654, 
    7.097704,
  3.324945, 4.661197, 3.58685, 5.18865, 5.990315, 5.035372, 5.03194, 
    4.519783, 4.076797, 2.620807, 2.850103, 4.580425, 5.266807, 5.14102, 
    4.120699,
  7.026899, 6.076353, 5.938957, 5.74843, 4.487033, 4.424012, 6.437444, 
    6.399878, 4.109198, 2.204661, 3.192816, 6.166247, 8.40239, 5.561035, 
    4.333514,
  11.41306, 9.694257, 8.736979, 8.14789, 7.970681, 6.687906, 7.927919, 
    7.867574, 6.589664, 5.802066, 5.810363, 6.641816, 9.637486, 10.01274, 
    6.652562,
  13.13645, 12.72431, 12.16792, 11.52611, 10.92968, 8.586721, 5.288869, 
    6.085059, 8.407784, 8.042767, 7.856328, 7.027654, 8.487322, 10.39392, 
    8.891323,
  11.7069, 12.0062, 11.93356, 11.63192, 10.23944, 8.624166, 7.152623, 
    4.152034, 4.251839, 5.1143, 7.682769, 7.358636, 7.846739, 10.61115, 
    10.73487,
  9.691937, 10.05785, 9.944374, 9.652772, 8.980604, 7.60631, 6.143782, 
    6.27997, 4.688306, 5.323975, 6.055204, 8.206379, 8.162006, 9.787657, 
    9.704897,
  7.962752, 8.15694, 8.041018, 7.807797, 7.718844, 7.713162, 7.011883, 
    6.384545, 6.125504, 7.03317, 7.964237, 8.467962, 8.961399, 9.321864, 
    9.22926,
  6.995246, 7.499608, 7.568061, 7.48751, 7.097023, 6.901573, 6.684433, 6.398, 
    5.729642, 5.762889, 6.294121, 6.923497, 7.442172, 7.677914, 7.426886,
  6.287759, 6.948289, 7.221578, 7.057464, 6.215367, 5.660274, 5.265417, 
    4.775769, 4.002716, 3.66809, 3.942865, 4.523659, 5.186311, 5.70668, 
    5.859753,
  4.817498, 5.224532, 5.583289, 5.383502, 4.875451, 4.341858, 3.76087, 
    3.270866, 2.782217, 2.370946, 2.857739, 3.754956, 4.181449, 4.42557, 
    4.514952,
  4.063093, 5.52918, 4.693204, 5.078868, 4.189802, 3.678061, 5.187124, 
    6.854042, 8.103045, 7.128722, 8.002794, 8.378294, 6.507639, 5.818626, 
    5.292125,
  7.161475, 6.141449, 5.543669, 4.788356, 3.650604, 3.988451, 6.079613, 
    7.067529, 8.247313, 8.584629, 8.108314, 9.598722, 9.12369, 5.460778, 
    4.511392,
  7.537874, 6.420023, 5.83829, 4.819464, 4.400695, 3.357798, 5.48945, 
    6.406963, 7.128817, 8.267559, 8.664932, 8.606221, 8.415209, 6.841357, 
    5.414375,
  7.897155, 7.481236, 7.170998, 6.38531, 5.255733, 4.160327, 2.365238, 
    4.944489, 7.7049, 8.288102, 7.98448, 7.353884, 7.114559, 6.755639, 
    5.396346,
  6.875486, 7.004159, 6.859826, 6.579339, 5.502967, 4.75954, 3.963162, 
    2.762068, 4.313725, 5.297597, 6.946974, 5.945016, 6.013834, 6.624986, 
    5.732248,
  4.375096, 4.703048, 4.668834, 4.614788, 4.616342, 4.920135, 4.862081, 
    5.068837, 4.561892, 5.628444, 5.092865, 4.996941, 4.522886, 6.608604, 
    6.041259,
  2.626914, 2.845414, 2.645634, 2.826238, 3.610639, 4.508487, 4.787837, 
    5.644962, 6.885816, 8.350297, 8.11008, 5.790379, 3.842766, 6.278813, 
    5.934032,
  2.382569, 2.704163, 2.648276, 3.024342, 3.538852, 3.593828, 3.527346, 
    4.001101, 4.871687, 6.847753, 8.030437, 7.251878, 5.104017, 6.214923, 
    5.94204,
  3.327787, 3.900385, 3.509055, 3.362324, 2.780252, 2.523487, 2.344489, 
    2.109015, 2.794287, 4.931823, 6.683977, 7.181183, 5.573553, 5.528216, 
    5.648085,
  3.187274, 3.011022, 2.686061, 1.943461, 1.677308, 1.73945, 2.296683, 
    1.886146, 0.9870979, 2.128285, 3.721301, 5.710023, 5.171721, 4.274569, 
    4.519774,
  2.463506, 4.039179, 4.305976, 6.034028, 5.914042, 5.308556, 7.993198, 
    9.083668, 9.617331, 7.452503, 6.78626, 8.113035, 10.18038, 8.804582, 
    6.976809,
  3.24172, 3.34972, 4.434185, 5.026849, 4.302467, 4.804021, 8.654188, 
    10.08146, 11.39578, 10.60198, 6.739723, 9.48319, 13.82394, 8.872798, 
    6.718905,
  3.476893, 2.771883, 3.080269, 3.622725, 4.21594, 3.969602, 7.70493, 
    9.124776, 10.95845, 11.85746, 8.721631, 9.981004, 14.23397, 13.30076, 
    9.010524,
  4.184581, 3.108205, 2.780439, 3.832949, 5.197693, 5.714309, 4.659194, 
    8.033169, 14.56778, 14.36623, 10.72937, 10.48071, 12.83917, 12.7441, 
    10.75559,
  5.206693, 4.147093, 3.005223, 2.991695, 4.246911, 6.793689, 7.165829, 
    5.642301, 7.977856, 9.081412, 10.48469, 10.88466, 11.97862, 11.92139, 
    12.12517,
  7.617042, 6.904759, 5.647019, 3.840427, 2.639913, 4.71749, 7.562216, 
    8.480468, 6.816887, 7.580768, 7.803361, 10.97612, 10.40281, 9.744331, 
    9.718484,
  8.141341, 7.896224, 7.53949, 6.165953, 3.627471, 2.359604, 5.713424, 
    8.564301, 10.56435, 11.48607, 10.80645, 10.59728, 9.847662, 9.073619, 
    8.565985,
  6.696235, 5.69837, 5.267569, 4.476182, 4.121151, 3.542518, 3.926772, 
    5.899568, 8.090914, 9.884747, 10.1409, 9.662423, 8.986651, 8.236636, 
    7.326674,
  6.468043, 4.681486, 4.142505, 4.538822, 4.835237, 5.192509, 4.413657, 
    4.073026, 5.843755, 8.023082, 8.604777, 8.165546, 7.508235, 6.990059, 
    6.544864,
  8.141651, 5.882261, 5.838133, 5.25644, 5.194846, 5.281798, 5.287919, 
    4.679672, 3.588427, 4.144383, 5.266311, 6.90426, 5.968462, 5.412266, 
    5.368721,
  6.007084, 7.539449, 6.245363, 7.886899, 7.61016, 6.348398, 8.824435, 
    7.864081, 6.327886, 5.150867, 5.163828, 4.594299, 3.951895, 3.942212, 
    3.548551,
  9.836522, 9.147225, 8.603543, 8.969646, 6.423924, 5.879911, 8.444431, 
    7.477467, 6.020135, 6.612463, 6.695105, 7.477695, 7.510789, 4.311496, 
    3.716669,
  9.514306, 9.267067, 8.908349, 9.354999, 7.808288, 6.037019, 6.428018, 
    4.729482, 4.940657, 6.86012, 8.843998, 9.203848, 8.835074, 7.759616, 
    6.027698,
  8.476702, 7.734901, 8.052903, 9.229112, 7.756389, 3.596658, 2.522702, 
    4.254344, 4.953768, 5.486028, 8.88323, 10.29218, 9.581718, 8.247446, 
    7.32965,
  7.467896, 5.677696, 6.920628, 7.651481, 5.602736, 4.270687, 3.864279, 
    2.651498, 3.256828, 3.991648, 8.561984, 10.56033, 10.34031, 8.959089, 
    8.188246,
  7.194434, 5.345214, 7.491236, 8.088925, 5.814638, 5.156504, 4.932249, 
    4.543606, 4.516096, 6.551526, 7.872529, 10.94283, 9.422538, 9.120632, 
    8.095545,
  8.056532, 6.880251, 8.32515, 8.160312, 7.95522, 7.453392, 7.720872, 
    7.94453, 8.7523, 10.83594, 11.43651, 10.88295, 9.436029, 9.563075, 
    8.741739,
  8.704347, 7.604408, 8.50326, 9.76717, 10.44617, 9.912295, 10.15338, 
    10.66499, 10.96731, 11.31661, 11.26324, 10.02467, 9.828753, 9.300145, 
    8.25456,
  9.24428, 8.65496, 10.38088, 12.05016, 11.41801, 10.84824, 10.93837, 
    11.28222, 11.19732, 10.51444, 10.17968, 9.586059, 9.380065, 8.51025, 
    7.093587,
  10.53145, 11.13988, 12.51499, 11.55982, 10.67438, 10.11968, 10.19351, 
    10.52472, 8.25924, 6.292176, 6.348064, 8.100892, 7.39935, 6.330917, 
    5.183959,
  7.650518, 12.20802, 10.84851, 12.98872, 10.74376, 8.124389, 9.968848, 
    9.711125, 9.36817, 6.506998, 6.001859, 6.072195, 4.799609, 4.308477, 
    4.419899,
  5.705524, 8.620122, 10.85404, 12.02848, 7.70952, 6.261999, 9.568454, 
    9.736969, 9.76605, 8.423285, 6.428238, 6.077674, 5.232408, 3.25658, 
    3.141626,
  4.02464, 5.500645, 8.242646, 10.9309, 8.7826, 5.946659, 7.710866, 7.580417, 
    6.450057, 6.838816, 5.931027, 3.28228, 2.887136, 3.976663, 3.600745,
  4.115305, 5.553671, 8.411047, 10.7197, 9.488341, 6.088063, 3.268903, 
    2.810126, 4.11876, 4.847726, 4.54446, 1.981103, 2.106177, 2.800617, 
    3.520234,
  3.516226, 4.370674, 6.028726, 7.415572, 8.021212, 6.022747, 5.286959, 
    4.503026, 3.720922, 3.3567, 3.653085, 2.686882, 2.767017, 2.638469, 
    2.648893,
  7.520443, 7.403225, 7.891272, 8.413143, 7.240082, 5.319914, 5.714954, 
    8.120917, 6.589386, 5.05024, 3.924739, 4.66406, 4.780559, 4.721537, 
    4.349187,
  10.672, 10.43814, 10.10994, 9.653752, 9.072618, 9.51789, 10.21122, 
    9.873931, 8.884652, 7.566541, 6.963684, 6.608361, 6.361864, 5.957064, 
    5.615534,
  12.7837, 13.02895, 12.98156, 12.74645, 12.50359, 12.87629, 12.78964, 
    11.64539, 9.887609, 8.456223, 7.731195, 7.112883, 6.395843, 5.687741, 
    5.005826,
  14.82227, 15.19453, 15.09516, 14.7492, 14.1454, 13.46896, 12.38451, 
    11.0602, 9.130594, 7.959527, 7.293401, 6.979262, 6.418846, 5.809186, 
    5.130359,
  14.85753, 15.07567, 14.81936, 13.98446, 12.83553, 11.38444, 10.03172, 
    9.400653, 6.914542, 5.060616, 5.086132, 6.278331, 5.995584, 5.578815, 
    5.193089,
  3.288126, 6.546033, 8.691699, 12.96469, 11.14573, 8.101997, 9.154812, 
    7.670301, 6.414485, 4.273284, 3.828339, 4.623392, 4.414782, 4.340955, 
    4.970497,
  4.014085, 5.273526, 8.49763, 11.69076, 8.341431, 6.74712, 9.013269, 
    7.882494, 6.320963, 5.35135, 4.537971, 5.993142, 7.07395, 5.076458, 
    5.095068,
  3.47171, 4.107701, 6.975731, 10.46323, 9.305791, 6.351601, 6.437128, 
    6.723073, 5.901901, 5.88487, 6.330989, 6.728478, 7.331079, 7.882483, 
    5.995027,
  3.45053, 4.853343, 7.726731, 10.66658, 12.05624, 8.745826, 5.235968, 
    3.32319, 2.48374, 4.206813, 4.887958, 5.248831, 5.455517, 5.757924, 
    4.958866,
  7.059029, 7.795032, 9.606691, 11.13224, 10.62507, 9.426773, 8.317603, 
    4.153512, 2.935398, 3.154444, 2.616132, 3.289755, 3.827099, 4.056417, 
    3.98061,
  10.50705, 11.01562, 11.40469, 11.42217, 10.22717, 8.006063, 6.468365, 
    5.663372, 3.071362, 1.327618, 1.057067, 2.298086, 3.025126, 3.006505, 
    2.774384,
  11.36248, 11.76425, 11.34451, 10.73006, 9.858697, 8.879578, 6.894938, 
    4.922043, 3.901877, 2.939642, 1.889001, 2.383472, 2.356346, 2.153875, 
    1.807775,
  11.35931, 11.60947, 11.16093, 10.70754, 10.15585, 9.588464, 8.375355, 
    6.75699, 4.86021, 3.644274, 3.114264, 2.963476, 2.654941, 2.233335, 
    1.926197,
  12.44788, 12.50515, 11.86807, 11.06083, 9.929377, 8.755733, 7.055882, 
    5.275887, 3.87925, 3.452933, 3.775861, 3.905756, 3.617913, 3.20663, 
    2.852906,
  12.33415, 11.96827, 10.97019, 9.362766, 7.555505, 6.088203, 4.571867, 
    3.823238, 2.671819, 2.191586, 2.804679, 3.811215, 3.859599, 3.589478, 
    3.266977,
  3.724024, 4.734351, 4.015353, 5.823142, 6.277359, 6.386002, 8.985866, 
    9.473833, 8.178412, 4.811536, 3.302145, 3.265589, 3.067654, 2.941719, 
    2.959477,
  4.866862, 3.690666, 3.547935, 5.72679, 6.00079, 6.168383, 8.71302, 
    8.874709, 6.822147, 5.12965, 3.443239, 3.666867, 4.048068, 3.403849, 
    3.430607,
  5.067159, 4.677657, 4.762616, 7.71773, 8.215933, 6.940046, 6.962729, 
    6.639726, 5.654957, 4.581093, 3.797457, 4.131487, 5.193696, 6.152781, 
    4.613594,
  5.205319, 5.764443, 6.659311, 9.239985, 10.63865, 8.770657, 6.229157, 
    4.052139, 1.593624, 3.160047, 4.18325, 4.917655, 5.46232, 5.457083, 
    4.037433,
  6.616492, 7.204059, 8.434149, 10.26839, 9.8043, 9.172959, 8.169889, 
    4.353103, 2.567197, 3.528427, 2.850871, 3.324821, 3.495812, 3.558246, 
    3.249512,
  8.359628, 8.81375, 9.584289, 10.28391, 9.24628, 7.282617, 6.350183, 
    5.271881, 2.200549, 1.147725, 1.069049, 1.486019, 2.47833, 2.662822, 
    2.62312,
  9.665668, 9.867461, 9.66452, 9.390837, 8.324152, 7.171093, 5.317752, 
    3.463836, 3.451741, 3.223553, 1.940684, 1.989976, 2.09551, 1.985329, 
    1.901598,
  9.620554, 9.291242, 8.393673, 7.871654, 7.212345, 6.71454, 6.177634, 
    5.275591, 3.874201, 2.359642, 2.098184, 2.317351, 2.436782, 2.38147, 
    2.225358,
  9.927986, 9.336452, 8.251928, 7.307794, 6.194212, 5.596499, 5.102601, 
    4.155066, 2.905432, 2.09942, 2.334165, 2.765225, 2.905003, 2.94988, 
    2.899883,
  9.523639, 9.156234, 8.116011, 6.389078, 4.79739, 3.976336, 3.896054, 
    3.626161, 2.555354, 1.258042, 1.307616, 2.460298, 2.988733, 3.032491, 
    3.160733,
  2.377323, 3.324789, 2.654313, 3.131397, 2.223197, 1.82025, 2.785603, 
    3.263569, 4.856977, 5.3222, 5.662945, 6.191155, 5.558879, 4.313589, 
    3.390664,
  2.62938, 1.854817, 1.552319, 2.230764, 2.716184, 3.349885, 4.80113, 
    6.607621, 8.447064, 8.615907, 7.149622, 7.108994, 5.779792, 3.350193, 
    2.985818,
  2.996348, 2.766411, 2.96158, 4.008781, 4.733012, 3.966421, 6.738122, 
    8.900436, 9.816621, 9.100948, 7.113141, 4.888041, 3.293997, 2.91595, 
    2.999497,
  4.003637, 4.239846, 4.845367, 5.714641, 5.99264, 6.030674, 4.950457, 
    6.886593, 7.883101, 5.659951, 4.418493, 2.969966, 2.43499, 2.710471, 
    2.434892,
  5.81096, 6.081522, 6.698955, 7.640128, 6.703606, 6.810206, 7.164852, 
    4.437575, 3.374688, 2.322455, 2.575337, 2.082636, 2.235031, 2.731896, 
    3.529291,
  6.241228, 7.116601, 7.836869, 8.427878, 7.748, 6.218494, 5.089957, 5.34856, 
    3.768525, 2.807863, 2.985573, 2.903576, 3.118748, 3.410064, 4.320805,
  5.909877, 7.047361, 7.480958, 7.760295, 7.615301, 7.461253, 6.36391, 
    5.425925, 5.056397, 4.666674, 3.865915, 3.336189, 3.434301, 3.850242, 
    4.667091,
  5.318964, 6.298123, 6.468415, 6.699001, 7.04322, 7.506001, 7.430766, 
    6.835417, 5.702538, 4.784174, 3.952062, 3.650365, 3.696484, 4.210918, 
    4.743052,
  5.410142, 6.238715, 6.421603, 6.788876, 7.336728, 7.572669, 6.98873, 
    6.082913, 5.257689, 4.600412, 4.20757, 4.158679, 4.251076, 4.565887, 
    4.856019,
  7.004964, 7.543252, 8.011435, 7.608167, 7.39236, 7.191501, 6.568009, 
    5.70717, 4.371089, 3.368517, 3.614686, 4.571617, 4.71652, 4.90143, 
    5.139664,
  2.604736, 3.164532, 3.268926, 4.120303, 4.311902, 4.584155, 5.613937, 
    5.031392, 4.258307, 3.406353, 3.573194, 4.104302, 4.016783, 3.847035, 
    3.079958,
  4.436202, 3.7448, 4.447227, 4.082877, 3.661724, 5.2749, 8.205246, 8.212709, 
    8.189522, 7.209296, 5.461368, 5.571701, 4.926123, 2.940957, 1.98823,
  5.176639, 4.188649, 4.581109, 3.734842, 3.667003, 3.582677, 6.496487, 
    7.911553, 8.261163, 7.789128, 6.71627, 5.600736, 4.683542, 2.593828, 
    1.370219,
  5.750343, 4.974338, 5.054529, 4.472768, 3.731646, 3.306556, 2.502589, 
    5.915532, 9.465473, 8.164799, 6.941185, 6.267991, 6.269579, 5.433208, 
    3.820894,
  6.077724, 5.451712, 5.398916, 5.185925, 4.06176, 3.964228, 3.441005, 
    3.197201, 4.09271, 4.730156, 6.133584, 6.468391, 7.068055, 7.208547, 
    6.926483,
  6.741251, 6.081148, 5.789247, 5.137516, 4.725662, 5.177565, 5.302907, 
    4.810399, 3.065775, 3.811877, 4.384554, 6.292449, 6.833614, 6.965579, 
    7.518078,
  7.546416, 7.170853, 6.315218, 5.352635, 5.377681, 6.396506, 6.852753, 
    6.698181, 6.010795, 6.102026, 5.957236, 6.195266, 6.354801, 6.32725, 
    6.847486,
  8.36742, 7.635324, 6.500051, 6.124116, 6.522049, 6.895284, 6.927755, 
    6.553693, 6.178686, 5.937274, 5.877733, 5.843189, 5.864657, 6.000105, 
    6.433581,
  9.196681, 8.333322, 8.051425, 8.015608, 7.821414, 7.433978, 6.625197, 
    5.998456, 5.840734, 5.654291, 5.705967, 5.723771, 5.749143, 5.626181, 
    5.656345,
  10.59894, 10.62177, 10.64707, 9.359697, 7.526596, 6.503716, 5.683999, 
    5.578397, 4.739279, 3.887856, 4.163688, 5.543253, 5.432811, 5.334173, 
    5.114191,
  6.807353, 9.124041, 7.113951, 8.122395, 6.005073, 4.372156, 4.796605, 
    3.997174, 3.687266, 2.687089, 2.733318, 3.366975, 3.050505, 2.904996, 
    2.983591,
  8.831664, 8.361941, 7.168569, 5.536273, 3.867169, 3.537392, 4.473014, 
    4.369362, 4.197387, 3.903658, 3.274778, 4.115681, 3.92576, 2.66155, 
    2.193841,
  8.072029, 6.77035, 4.964127, 3.032902, 2.550826, 2.128685, 3.096367, 
    3.60364, 3.714895, 4.107339, 4.59217, 4.922691, 4.922778, 3.589652, 
    1.42828,
  6.717324, 5.488729, 4.102933, 2.783672, 1.847437, 2.264378, 1.496587, 
    3.188708, 5.302355, 4.765328, 4.90771, 5.156133, 5.191102, 4.385972, 
    2.659636,
  5.9424, 4.594004, 4.060941, 4.076907, 3.777309, 3.228359, 2.540616, 
    2.228524, 2.560252, 3.196076, 4.252009, 5.033411, 5.483032, 5.481641, 
    4.992775,
  6.335068, 4.723277, 4.26685, 4.19932, 4.341737, 4.770409, 4.400479, 
    2.78123, 1.514744, 2.435818, 3.135594, 4.629334, 5.375052, 5.880297, 
    6.57367,
  7.181074, 5.045915, 4.306807, 4.241221, 4.438647, 4.526045, 4.717887, 
    4.477593, 3.892189, 3.919939, 3.959473, 4.375764, 5.042978, 5.43095, 
    6.088218,
  7.688771, 5.032829, 4.674617, 4.924415, 4.900226, 4.361449, 3.883674, 
    3.449731, 3.4598, 3.739686, 3.766874, 3.848321, 4.163296, 4.508969, 
    4.916742,
  7.671663, 6.150377, 6.692809, 6.165352, 5.613476, 4.685407, 3.675915, 
    2.897419, 2.947943, 3.236629, 3.327361, 3.27059, 3.180697, 3.213784, 
    3.052262,
  8.947272, 8.731135, 8.634392, 6.93815, 5.409757, 4.211857, 3.241178, 
    2.540363, 2.216949, 1.798685, 1.813828, 2.209969, 2.144483, 1.938732, 
    1.757054,
  8.933265, 12.63888, 10.64474, 13.9363, 12.15591, 9.355865, 11.19816, 
    10.089, 8.628136, 5.115265, 3.688205, 2.742298, 2.204127, 1.982841, 
    1.935941,
  10.98292, 11.38388, 11.49973, 11.15157, 7.909095, 6.552531, 8.956481, 
    7.807144, 6.462614, 4.603543, 2.552436, 1.927439, 2.266265, 2.567001, 
    2.683758,
  8.907149, 8.684194, 8.822289, 8.083841, 6.019164, 4.331905, 5.463171, 
    5.598244, 4.871892, 3.527794, 1.920926, 1.869841, 2.652546, 3.239308, 
    2.685951,
  6.213506, 6.554322, 6.714542, 5.664972, 4.70944, 4.610734, 3.128763, 
    3.931854, 3.823419, 2.728544, 2.338439, 2.696074, 2.491395, 1.767868, 
    1.979356,
  4.763286, 5.413214, 5.699361, 5.214414, 3.619991, 3.207037, 4.485005, 
    2.670512, 0.9432118, 1.376331, 2.727388, 3.193958, 2.400407, 1.906397, 
    2.583785,
  4.482621, 4.857017, 4.93811, 4.446016, 3.839671, 3.122361, 2.598891, 
    3.279921, 2.574504, 1.747135, 2.628631, 3.532408, 3.865379, 3.684774, 
    3.382041,
  4.800951, 4.607007, 4.407052, 3.804446, 3.631621, 4.3687, 4.683091, 
    4.462212, 3.677396, 2.95159, 2.77546, 3.343428, 3.531154, 3.084197, 
    2.328977,
  4.945456, 3.955348, 3.934414, 3.23446, 3.473798, 4.631608, 4.991404, 
    4.31945, 3.033527, 2.1451, 2.19438, 2.684177, 3.115558, 3.230621, 3.059644,
  3.716348, 2.692842, 3.942521, 3.734946, 4.14483, 5.034891, 4.877035, 
    3.465399, 2.287026, 1.93058, 2.194803, 2.804352, 3.550802, 4.408499, 
    4.940699,
  5.190265, 5.662534, 5.546874, 4.937419, 4.519971, 4.388822, 3.917203, 
    3.053207, 2.377297, 1.739889, 2.289557, 3.801101, 5.134641, 6.716304, 
    7.874723,
  9.181049, 13.11982, 11.72984, 15.31936, 14.79456, 12.0352, 15.77458, 
    15.53963, 15.13514, 10.10958, 9.10917, 9.21134, 8.770933, 7.786312, 
    5.733503,
  11.00777, 12.98553, 14.50397, 14.92954, 11.90034, 11.91155, 17.22258, 
    16.18213, 15.02888, 12.42273, 9.41427, 9.916623, 9.205894, 5.815994, 
    4.271616,
  8.753013, 10.24861, 12.11851, 12.30142, 9.274858, 7.565269, 11.07024, 
    13.42954, 12.61765, 11.36473, 9.644917, 8.208684, 7.045415, 6.034934, 
    4.62219,
  6.797002, 8.314024, 9.549659, 9.843519, 9.037498, 6.487185, 4.377428, 
    7.755252, 9.232929, 7.278325, 6.06655, 4.852654, 4.542503, 4.470607, 
    4.387825,
  5.70842, 6.582566, 7.510178, 7.888657, 6.914118, 5.644403, 4.900199, 
    3.332385, 2.963447, 2.867899, 3.606115, 2.889714, 2.465987, 2.610399, 
    3.296868,
  5.010841, 5.262913, 6.140001, 5.977821, 5.707853, 4.605525, 3.750579, 
    3.919556, 3.078466, 1.702433, 2.013566, 1.713802, 1.65304, 1.549415, 
    1.885185,
  6.566417, 5.238867, 4.261615, 3.750982, 3.879555, 4.261562, 3.845536, 
    2.986428, 1.79664, 1.483126, 1.80403, 2.161171, 2.243519, 2.171316, 
    1.89843,
  9.305581, 9.294168, 6.827005, 4.588328, 3.053024, 3.112835, 2.632316, 
    2.767666, 3.089704, 4.201698, 5.098217, 5.591687, 5.609611, 5.363031, 
    4.688654,
  6.971587, 8.490836, 5.8252, 4.36876, 4.439495, 3.278146, 2.933362, 
    3.925439, 5.864307, 7.298258, 8.079697, 9.01154, 8.966953, 8.838226, 
    7.590121,
  4.840448, 5.812581, 6.651137, 7.568285, 5.516306, 4.093489, 4.426734, 
    6.198977, 7.198628, 6.172516, 7.896704, 11.91826, 12.38097, 12.46356, 
    11.12653,
  6.714076, 11.56013, 10.68688, 13.00597, 12.69321, 10.22493, 9.857308, 
    7.138762, 7.123812, 5.275975, 5.209972, 6.883826, 7.826876, 7.184661, 
    5.730278,
  7.222783, 10.48148, 12.80395, 13.09474, 9.999922, 11.44134, 15.61011, 
    12.98468, 10.86195, 8.743242, 6.966595, 8.798603, 10.16635, 6.884584, 
    5.635273,
  7.067636, 8.235501, 10.79074, 12.22121, 9.216439, 7.332664, 11.73979, 
    15.15478, 14.44071, 12.23922, 10.61191, 10.15979, 10.30419, 9.609786, 
    7.083537,
  6.750349, 7.837406, 9.041272, 10.00671, 10.34359, 6.484506, 4.329642, 
    10.54856, 14.42114, 12.40777, 11.18395, 10.78628, 10.56819, 9.179466, 
    7.172898,
  5.807842, 6.177511, 6.852155, 6.670012, 7.28719, 7.66071, 5.171988, 
    4.066459, 5.329873, 6.116657, 7.960858, 8.328808, 9.050336, 8.398044, 
    7.089611,
  6.298443, 4.976714, 4.435468, 3.882715, 2.982712, 3.572549, 4.275075, 
    3.75982, 2.048203, 2.043362, 3.586778, 5.260587, 6.30233, 6.749297, 
    6.745426,
  8.363139, 5.94104, 3.54805, 2.579353, 2.397321, 2.07099, 1.523731, 
    2.288153, 2.726691, 2.35889, 2.643382, 3.672399, 4.556922, 5.180971, 
    5.642932,
  7.505007, 5.496239, 4.653592, 3.390452, 3.357453, 4.031478, 4.404677, 
    4.058021, 6.202883, 6.958578, 6.459185, 5.870418, 5.407043, 5.1408, 
    5.349922,
  6.559212, 6.295129, 4.640364, 3.787896, 4.005131, 5.093758, 5.305789, 
    5.283677, 5.70785, 6.545276, 8.631816, 9.164701, 8.356159, 7.472453, 
    6.129193,
  7.920549, 7.411219, 6.486041, 5.106052, 5.087946, 5.736691, 5.519982, 
    4.617361, 3.850082, 3.331241, 4.830999, 9.901758, 10.94197, 10.10206, 
    7.987736,
  4.180389, 6.168169, 5.668745, 8.351419, 8.721951, 7.778723, 8.894515, 
    3.787718, 1.941056, 2.448217, 2.739174, 3.704023, 3.854388, 3.754405, 
    3.095796,
  5.763111, 6.162735, 5.67428, 6.624306, 5.872149, 6.546904, 10.59215, 
    9.521228, 5.833081, 2.697208, 1.61934, 3.976188, 6.0842, 4.086301, 
    3.373453,
  7.071506, 6.040445, 3.908087, 4.200082, 4.587101, 4.217044, 7.424599, 
    10.03207, 10.5731, 9.288918, 6.257605, 3.52582, 3.810812, 5.696108, 
    4.890101,
  8.550479, 7.991414, 4.162094, 2.526881, 3.871739, 3.447041, 2.555683, 
    7.146793, 11.23398, 10.95975, 9.297104, 7.2772, 4.865152, 3.172613, 
    4.647818,
  9.170203, 8.36085, 4.590378, 2.444665, 1.920238, 2.958726, 2.230921, 
    2.622861, 4.48647, 5.734901, 7.170362, 7.018778, 6.389301, 4.70876, 
    3.336484,
  9.113062, 7.32044, 2.924424, 1.702448, 2.011428, 1.110661, 1.565956, 
    1.532612, 0.7297996, 2.500839, 4.047672, 5.680657, 6.035442, 5.62008, 
    4.881455,
  7.8207, 4.648525, 2.985725, 2.268956, 1.616414, 1.996624, 1.498075, 
    0.9579957, 0.7784835, 1.469261, 2.531255, 4.028845, 5.264916, 5.664977, 
    6.515962,
  5.203276, 4.436409, 4.905917, 2.869181, 2.16095, 2.360906, 2.085, 1.676523, 
    1.302011, 1.46636, 1.403993, 2.283638, 3.763879, 4.906043, 6.003836,
  4.46609, 4.859188, 5.186096, 3.119179, 2.131431, 2.02635, 1.646249, 
    1.288973, 1.945724, 2.114513, 1.337048, 2.30304, 3.10746, 4.063775, 
    4.713543,
  4.507638, 4.828298, 4.334645, 2.343944, 2.18489, 2.22384, 1.926804, 
    1.211731, 1.251309, 1.074523, 1.29796, 1.773316, 3.458335, 3.982415, 
    4.208992,
  4.299973, 4.572807, 3.216139, 2.746847, 2.192267, 2.655215, 5.019428, 
    5.766331, 4.517214, 2.09637, 1.403433, 1.239388, 1.972906, 2.800297, 
    2.631286,
  7.750441, 6.449234, 4.483675, 3.530564, 2.296478, 1.928893, 4.139105, 
    5.712608, 6.498797, 5.358572, 3.154016, 2.170493, 1.77562, 0.9898524, 
    1.005877,
  9.556479, 8.456779, 6.097873, 4.506954, 3.415371, 1.688359, 2.081042, 
    3.21687, 5.09072, 6.667306, 6.776878, 5.650879, 3.392694, 2.60707, 
    1.736146,
  10.40697, 10.42517, 8.404405, 5.579846, 4.735682, 3.390818, 1.493101, 
    2.241912, 5.336684, 5.880439, 6.139112, 6.574358, 6.431525, 4.718031, 
    2.759752,
  10.58465, 10.94737, 9.612772, 6.718136, 5.052522, 3.780158, 3.258166, 
    1.80189, 2.196025, 2.648139, 4.288968, 5.351207, 6.078061, 6.28203, 
    4.716318,
  10.33187, 10.82676, 9.823875, 7.187252, 5.505502, 3.860728, 1.999046, 
    1.835453, 2.187688, 1.767677, 2.611942, 4.087735, 5.242029, 5.938504, 
    6.237403,
  9.858362, 10.30295, 9.76491, 7.497544, 5.86605, 4.774475, 3.344147, 
    2.84036, 2.964615, 2.333542, 2.347682, 3.043882, 4.221778, 5.176788, 
    5.850594,
  9.21613, 9.752844, 9.677572, 7.701788, 5.387705, 4.723897, 4.611523, 
    3.733225, 2.956976, 2.226747, 2.095664, 2.406821, 3.521655, 4.746377, 
    5.580483,
  8.698319, 9.329983, 9.479807, 7.7833, 5.277115, 4.854648, 5.133233, 
    4.178118, 3.363662, 2.531107, 2.090187, 2.050376, 3.138815, 4.470817, 
    5.303863,
  8.49652, 9.290187, 9.222922, 6.962132, 5.359644, 5.300233, 5.252917, 
    4.792628, 3.743461, 1.963314, 1.593533, 1.984758, 2.647186, 3.983359, 
    4.975543,
  2.655463, 3.413733, 3.682619, 6.057751, 5.765499, 2.972319, 2.176325, 
    2.229636, 2.957948, 2.222842, 1.611277, 1.417403, 1.408452, 2.106115, 
    1.930278,
  5.037313, 4.153607, 4.854711, 6.774251, 5.321348, 2.717974, 1.823143, 
    2.275056, 3.057496, 3.5418, 3.085677, 3.309287, 2.469192, 1.928035, 
    1.687955,
  6.636138, 6.431565, 6.237018, 7.605649, 6.384414, 3.078604, 1.490473, 
    1.706368, 2.266664, 3.028497, 3.915357, 4.793106, 4.744298, 3.962957, 
    2.917556,
  7.783188, 8.292048, 8.298461, 8.724997, 8.777021, 5.658094, 2.685153, 
    2.146304, 2.279774, 1.679173, 2.880729, 3.604036, 4.30567, 4.545714, 
    4.029346,
  8.492778, 8.924681, 9.224543, 9.588288, 8.777426, 7.363444, 5.993827, 
    2.671385, 1.870795, 1.894027, 2.350773, 2.465878, 3.279184, 3.75984, 
    3.901818,
  9.117317, 9.499712, 9.713428, 10.12562, 9.560122, 7.435246, 5.949619, 
    4.068042, 2.423132, 3.441428, 3.095746, 2.696088, 2.834047, 3.665516, 
    4.499185,
  8.866316, 9.544811, 9.925311, 10.34565, 10.24671, 8.447514, 5.500404, 
    3.186479, 3.724685, 4.91357, 4.517084, 3.181378, 2.700478, 3.717192, 
    5.069798,
  7.075018, 8.455081, 9.559328, 10.28053, 10.28511, 8.921043, 6.610458, 
    5.657071, 5.238514, 4.782473, 4.494323, 3.291362, 2.836208, 4.226069, 
    5.740092,
  5.093663, 6.819864, 8.347121, 9.596598, 9.519036, 8.001059, 7.419577, 
    6.984467, 5.897707, 4.97144, 4.317304, 3.482777, 3.082431, 4.485919, 
    5.881731,
  4.911364, 6.031469, 7.395377, 7.908233, 7.703626, 7.713835, 8.245022, 
    7.835506, 5.295374, 3.534148, 3.537743, 3.774185, 3.280375, 4.349156, 
    5.727548,
  3.213648, 3.131639, 1.819071, 1.52105, 3.13458, 3.775473, 4.201134, 
    3.332879, 4.4622, 3.588292, 3.389316, 3.628006, 2.937365, 2.645608, 
    1.770232,
  3.688361, 2.935173, 2.534641, 3.128959, 3.213398, 3.744381, 4.821379, 
    3.514113, 3.477027, 3.861848, 3.37558, 4.196087, 3.809705, 2.46497, 
    1.420357,
  3.46019, 4.185769, 4.112935, 3.922202, 3.73186, 2.629889, 4.052079, 
    4.410627, 4.414268, 4.471204, 4.661388, 5.054501, 4.349944, 3.503078, 
    2.372346,
  3.802916, 5.717462, 5.603534, 4.601357, 4.18013, 3.265981, 2.547529, 
    4.303767, 5.13151, 4.561037, 5.52612, 5.691565, 5.057652, 3.952034, 
    2.825493,
  3.627936, 6.093613, 6.218638, 5.111734, 3.67424, 3.098307, 4.528083, 
    2.849633, 2.257366, 2.940844, 4.666784, 4.903395, 4.222312, 2.968188, 
    1.840898,
  3.284883, 6.6545, 7.232192, 5.987168, 5.03033, 3.649756, 3.215405, 
    2.978044, 3.644505, 4.276067, 3.810409, 4.426199, 3.357457, 2.666203, 
    2.812813,
  2.8058, 6.958509, 7.656582, 6.466801, 6.090472, 4.865005, 3.325897, 
    2.343074, 5.147399, 6.329541, 5.707022, 4.371098, 3.02133, 3.032267, 
    3.55914,
  3.064147, 7.318744, 8.073634, 6.611314, 6.376267, 5.774895, 4.880862, 
    4.976156, 6.371394, 6.595588, 5.789921, 4.010737, 3.09404, 3.611454, 
    4.231545,
  3.430907, 7.569471, 8.826347, 7.162249, 6.603192, 6.466393, 5.687428, 
    5.70614, 6.415429, 6.219902, 5.253743, 3.697103, 3.26188, 3.97651, 
    4.348477,
  3.543499, 6.672317, 8.730539, 7.164937, 6.099807, 6.485456, 6.75035, 
    6.685686, 5.567986, 4.081356, 3.844059, 3.609652, 3.329228, 4.125678, 
    4.507218,
  5.530205, 6.250065, 4.348656, 5.028918, 3.465563, 3.113167, 4.669001, 
    4.159874, 3.053542, 2.165881, 2.246592, 3.311704, 4.011841, 3.921091, 
    3.050169,
  7.496229, 6.639652, 6.162572, 5.741653, 3.341407, 2.552392, 3.916958, 
    3.622379, 2.638955, 2.581893, 2.580409, 4.142756, 5.568186, 3.466331, 
    2.979677,
  7.065361, 6.448265, 6.710683, 6.460086, 4.060613, 2.181515, 2.866496, 
    3.311291, 3.272834, 3.507001, 3.9653, 4.592401, 5.165792, 5.228354, 
    4.232298,
  6.601122, 7.022759, 7.980389, 6.646387, 4.034545, 2.486001, 1.256644, 
    3.483155, 5.516728, 5.026339, 5.47837, 5.946182, 6.105325, 5.5905, 
    4.489399,
  6.133731, 8.226214, 9.265897, 6.4002, 2.597295, 1.619999, 2.767957, 
    2.196144, 2.065088, 3.254878, 5.371854, 6.271091, 6.350683, 5.74043, 
    4.285623,
  7.587534, 9.924611, 9.43838, 5.767109, 2.925173, 1.288329, 1.320519, 
    3.510117, 4.0756, 3.935264, 4.222139, 5.655923, 5.390379, 4.995909, 
    3.897138,
  9.796251, 10.78021, 9.05715, 5.352292, 3.052191, 2.905793, 4.147434, 
    4.916526, 5.79678, 6.215475, 5.996344, 5.381734, 4.585981, 4.088945, 
    3.392522,
  10.91321, 10.7186, 8.23959, 4.897991, 4.121412, 5.346821, 6.29471, 
    6.645581, 6.933332, 6.632696, 5.719083, 4.606791, 3.883716, 3.659122, 
    3.385519,
  11.08407, 10.25726, 7.473332, 5.732379, 6.331406, 6.832181, 6.519651, 
    6.534908, 6.616066, 5.59047, 4.618542, 3.863083, 3.631714, 3.796288, 
    3.47271,
  10.72166, 9.865647, 7.898799, 6.86658, 6.473637, 6.4201, 6.210479, 
    6.097027, 4.808072, 3.218984, 3.11221, 3.365847, 3.394247, 3.565579, 
    3.545329,
  4.596758, 7.02112, 6.321066, 8.583488, 7.562239, 5.153273, 6.62885, 
    6.338374, 5.428856, 4.032948, 3.921038, 4.498856, 4.344049, 4.164762, 
    3.797297,
  6.850652, 7.587802, 7.619163, 7.542422, 3.696209, 4.091378, 5.576503, 
    5.268101, 4.731496, 3.871149, 3.340271, 4.710061, 6.019967, 4.17311, 
    3.660585,
  7.34382, 6.752494, 6.624101, 5.669584, 5.653619, 4.955882, 4.655605, 
    4.385701, 3.722146, 2.697479, 2.222432, 3.455669, 5.511128, 6.330976, 
    5.380731,
  7.493269, 6.854589, 6.634005, 7.727946, 7.845821, 5.024106, 3.578867, 
    3.875199, 4.157333, 3.028644, 1.491765, 2.339915, 4.595984, 6.045479, 
    6.486456,
  7.568204, 7.88624, 9.152049, 9.383375, 7.926709, 5.580814, 4.554688, 
    2.926377, 1.571719, 1.575846, 2.274393, 2.497187, 5.118585, 6.732787, 
    7.266587,
  9.109754, 9.38274, 9.212757, 8.582067, 7.573466, 6.298562, 5.041969, 
    4.065621, 2.797183, 2.355834, 2.61148, 4.153255, 5.950121, 7.287766, 
    7.521283,
  9.616075, 9.240609, 8.668174, 7.796725, 7.020594, 6.937008, 6.700441, 
    5.974594, 5.257016, 5.051615, 5.17659, 6.219406, 7.424488, 8.384464, 
    8.97604,
  9.218278, 8.968129, 8.574813, 8.124071, 7.723718, 7.590091, 7.194547, 
    6.853125, 6.600998, 6.383423, 6.657809, 7.352658, 7.977158, 8.701903, 
    8.909435,
  8.254478, 8.528157, 8.495124, 8.372562, 8.143888, 7.73815, 7.00154, 
    6.784594, 6.769297, 6.408043, 6.749629, 7.390018, 7.67099, 7.898256, 
    6.787302,
  6.646924, 7.065726, 7.137675, 6.542143, 6.077387, 6.201035, 5.930054, 
    5.81261, 5.102727, 4.006207, 4.624669, 6.530742, 6.547353, 6.357418, 
    5.608847,
  4.007155, 5.212507, 5.177567, 7.215271, 6.579455, 4.389714, 5.370503, 
    5.787821, 5.068422, 3.472503, 3.30725, 3.705398, 3.80897, 4.288052, 
    4.824895,
  5.116595, 4.980296, 5.272219, 7.030739, 5.247229, 4.136146, 5.405674, 
    5.523267, 5.261274, 4.743004, 3.836553, 4.042168, 4.071477, 2.866246, 
    3.819068,
  5.365892, 4.036645, 4.229584, 6.145126, 5.745682, 3.749592, 4.845569, 
    4.911935, 4.454433, 4.74206, 4.610852, 4.172168, 4.050005, 4.65553, 
    5.458092,
  6.866332, 7.43815, 7.417689, 6.704844, 7.601987, 5.881294, 3.287648, 
    4.402752, 6.297812, 5.413006, 4.163486, 2.880849, 3.660437, 4.984319, 
    6.126682,
  7.018579, 7.821485, 8.38773, 7.578844, 7.049031, 7.795364, 5.964621, 
    3.170521, 3.717753, 3.822631, 3.673659, 2.063841, 3.662388, 5.564099, 
    6.71393,
  6.822623, 7.631293, 8.534897, 8.25275, 7.346864, 7.811225, 8.083214, 
    6.447409, 4.757772, 3.989417, 2.395247, 2.48888, 4.297789, 5.793304, 
    6.278193,
  6.38152, 7.224325, 8.207752, 8.809416, 8.530273, 8.174342, 8.317059, 
    8.310685, 7.585647, 6.242518, 4.327268, 4.301663, 5.464783, 6.245535, 
    7.112971,
  5.830729, 6.456906, 7.16512, 8.373369, 9.102818, 8.846511, 8.128154, 
    7.993776, 8.201088, 7.835663, 6.661909, 6.602293, 7.029846, 7.711701, 
    8.42747,
  5.774872, 5.771883, 5.631555, 6.324038, 7.556821, 8.005405, 7.59142, 
    7.664025, 8.04439, 8.296699, 8.058366, 8.086936, 8.264865, 8.349346, 
    7.289204,
  5.987809, 5.355644, 4.446199, 3.745453, 4.82732, 6.337551, 6.847159, 
    6.866543, 6.283371, 5.215593, 5.598852, 7.855842, 7.804135, 7.541958, 
    6.300257,
  4.397202, 4.348351, 3.685079, 4.917318, 5.086413, 4.203467, 5.908451, 
    6.195679, 5.350577, 3.995894, 4.262474, 4.604365, 3.553554, 2.907412, 
    2.558155,
  6.138947, 4.404757, 4.055943, 4.496314, 4.198717, 4.08277, 6.136395, 
    6.610194, 6.33562, 5.261529, 4.26008, 4.500748, 2.860173, 1.974155, 
    2.163019,
  6.350414, 4.131943, 3.741776, 3.870939, 4.200151, 3.509809, 5.647336, 
    6.296444, 5.68375, 5.520862, 5.259545, 4.35856, 3.001687, 2.549492, 
    4.428608,
  7.365188, 6.076111, 6.139303, 4.460297, 5.167321, 4.686858, 3.502344, 
    5.60323, 8.751656, 8.184301, 6.744844, 5.583506, 5.10619, 5.625607, 
    6.435296,
  7.599554, 5.96784, 6.529662, 6.094005, 4.819973, 5.665895, 4.960911, 
    3.405502, 4.937439, 5.581117, 6.81768, 6.765988, 6.845968, 7.414542, 
    7.778358,
  8.253222, 5.801217, 6.313159, 6.499375, 5.525357, 5.164592, 5.766839, 
    5.148915, 3.967426, 4.50115, 4.677162, 7.321852, 8.024026, 8.539442, 
    8.580484,
  8.73038, 6.051154, 5.864623, 6.831719, 5.855355, 5.205044, 5.331966, 
    6.107622, 6.524114, 6.936315, 6.60336, 7.337554, 7.976656, 8.525998, 
    9.07717,
  9.563788, 7.033384, 5.342176, 7.385615, 6.370974, 5.294985, 4.927736, 
    5.211631, 5.980787, 6.539163, 6.78172, 7.041519, 7.434502, 7.959757, 
    8.209147,
  10.44634, 8.086143, 5.03802, 8.079563, 7.519607, 5.663121, 4.636438, 
    4.348542, 5.148601, 5.785421, 6.193146, 6.407738, 6.617872, 6.735303, 
    6.167296,
  10.94412, 8.846152, 5.763844, 7.82883, 9.725867, 6.679091, 4.613615, 
    4.119566, 3.909941, 3.453247, 3.990667, 5.312953, 5.180909, 4.949526, 
    4.504261,
  7.017314, 6.009379, 7.635952, 8.175966, 4.726665, 2.758483, 3.002658, 
    3.54646, 3.760348, 3.095459, 3.409144, 3.983519, 4.019845, 3.400181, 
    2.683553,
  10.5929, 6.593845, 10.63129, 8.389393, 4.097288, 3.164072, 4.323673, 
    4.805409, 5.228672, 3.881326, 2.098542, 2.897654, 4.514848, 3.29515, 
    2.638412,
  10.27293, 6.940237, 11.30731, 8.464349, 4.750302, 2.522837, 4.505389, 
    5.681637, 6.182662, 5.84776, 4.810209, 4.444657, 4.400125, 4.521682, 
    3.553662,
  9.971231, 7.170192, 11.41359, 8.83647, 5.420275, 3.700067, 2.225171, 
    5.516699, 9.897442, 8.92067, 7.134856, 6.104386, 5.207756, 4.203278, 
    3.795086,
  9.964257, 7.883896, 10.8931, 10.61452, 6.698012, 5.379653, 4.320599, 
    3.385959, 5.002897, 5.697402, 6.892425, 6.665791, 6.254649, 5.299433, 
    4.567837,
  10.11054, 9.026964, 10.16592, 12.48347, 9.224872, 7.702087, 6.723919, 
    6.10544, 3.723334, 4.858142, 5.449049, 7.941567, 8.209489, 7.987656, 
    7.73316,
  10.23565, 10.34508, 10.41031, 13.59895, 10.57414, 9.156338, 7.801009, 
    7.422705, 7.495994, 8.225508, 8.028272, 8.728455, 8.854885, 8.778734, 
    8.676483,
  10.39291, 10.91601, 10.68856, 13.80491, 11.32786, 9.812711, 8.284776, 
    7.950888, 7.833326, 8.068604, 8.167875, 8.397985, 8.33637, 8.461627, 
    7.993256,
  10.33517, 10.72343, 10.9563, 14.1122, 12.26036, 10.45848, 8.524474, 
    7.787858, 7.557091, 7.366313, 7.536875, 7.698954, 7.75028, 8.036801, 
    7.741229,
  10.18066, 10.16878, 10.95395, 13.70377, 12.52752, 10.31137, 8.619662, 
    7.590051, 5.877256, 4.754426, 5.285691, 7.503208, 7.404661, 7.767132, 
    7.784039,
  6.735251, 8.593094, 6.013465, 6.656524, 5.788588, 5.206618, 5.580133, 
    2.941958, 1.478409, 1.994853, 2.88095, 3.835838, 4.170156, 4.037362, 
    3.563703,
  9.845153, 8.685614, 7.374119, 5.922732, 4.40455, 4.934627, 7.174548, 
    5.847574, 3.217604, 1.744008, 2.760353, 4.304909, 5.443959, 3.794063, 
    3.428433,
  10.25306, 8.598551, 7.873216, 6.98143, 5.215424, 3.633089, 6.102593, 
    6.48616, 4.983178, 3.019213, 3.13136, 4.249056, 5.251079, 5.586034, 
    4.691283,
  10.02292, 9.255935, 8.896137, 8.479557, 8.347184, 5.829399, 3.224273, 
    6.009656, 8.737659, 5.669368, 2.830338, 3.524357, 5.117895, 5.941002, 
    5.910652,
  10.06864, 9.760349, 9.649944, 9.68277, 9.721323, 9.395734, 7.140353, 
    4.225637, 5.087614, 4.727176, 4.091534, 3.255225, 4.458701, 6.014872, 
    7.369195,
  10.12117, 9.958644, 9.906973, 9.904728, 10.21417, 10.79558, 10.61357, 
    9.025954, 6.006954, 5.775167, 3.851494, 3.652087, 3.973213, 4.928133, 
    6.116441,
  10.07072, 10.15192, 10.1473, 10.28801, 10.63437, 10.88567, 10.9017, 
    11.0077, 11.44601, 11.41365, 8.950985, 5.433736, 4.15829, 4.265644, 
    5.180583,
  10.20623, 10.45019, 10.5681, 10.90765, 11.25677, 11.163, 10.98646, 
    11.27961, 11.78936, 12.53364, 12.19423, 9.361794, 6.112007, 4.87158, 
    4.988081,
  10.42565, 10.72374, 10.87278, 11.0466, 11.12784, 10.94328, 10.95766, 
    11.3565, 11.83988, 12.38731, 13.22483, 12.68684, 9.539623, 7.122937, 
    6.134631,
  10.7664, 10.99806, 10.98173, 10.76848, 10.50628, 10.46523, 10.13439, 
    10.66608, 9.389489, 7.996468, 9.643641, 13.62806, 12.4796, 9.916165, 
    7.694248,
  3.147098, 4.506719, 4.803689, 5.872737, 4.279723, 3.562809, 4.405045, 
    3.463586, 2.279666, 1.883888, 1.804398, 2.814018, 2.970123, 3.106664, 
    3.64239,
  3.600337, 4.009491, 6.37694, 6.675806, 4.443701, 3.692502, 5.256959, 
    4.339206, 2.111879, 2.341742, 1.383815, 2.400036, 3.511693, 2.765628, 
    3.14451,
  5.283635, 4.120203, 5.925281, 7.935366, 6.283111, 3.599502, 5.318992, 
    5.039168, 2.175535, 2.10182, 2.85414, 2.309388, 3.543442, 3.910249, 
    3.698262,
  6.671097, 7.085452, 7.676769, 8.470203, 9.161263, 6.648427, 3.763818, 
    4.909752, 6.232865, 1.794448, 3.014253, 3.239023, 3.658469, 4.600595, 
    4.441005,
  7.334021, 8.115564, 8.454964, 8.476722, 9.135614, 9.538419, 6.943838, 
    3.632034, 4.185579, 2.855028, 1.906628, 4.01066, 4.112788, 4.779595, 
    5.282991,
  7.671347, 8.523319, 8.85862, 9.001515, 9.290334, 9.77247, 9.335911, 
    7.042622, 5.06898, 3.802109, 1.45116, 4.151901, 4.732996, 4.856647, 
    5.412839,
  8.016011, 8.920809, 9.479537, 9.883525, 10.25152, 10.27199, 9.917336, 
    9.290854, 9.017709, 7.466576, 2.401215, 3.510498, 4.633615, 5.139052, 
    5.425382,
  8.080739, 9.138443, 9.9752, 10.75331, 11.08182, 10.97369, 10.4092, 
    9.425683, 9.234733, 9.246675, 6.089331, 2.182959, 4.512594, 5.289927, 
    5.625956,
  8.065344, 8.998033, 9.836545, 10.60917, 10.9677, 11.11761, 11.17597, 
    10.50808, 10.04063, 9.811533, 8.703123, 4.022555, 3.16284, 5.394681, 
    5.881886,
  7.768325, 8.628949, 9.336848, 10.02389, 10.5492, 11.08869, 11.30782, 
    11.12834, 8.949922, 6.616657, 6.68038, 7.405001, 2.958947, 4.261409, 
    5.757795,
  2.863268, 3.500072, 3.324294, 3.64834, 2.21959, 1.985795, 3.16348, 
    3.676548, 3.354009, 3.006743, 3.149232, 3.289993, 2.927173, 2.542456, 
    2.563128,
  2.188134, 2.052257, 3.99236, 4.410567, 2.820272, 2.558352, 3.828746, 
    4.141441, 3.696092, 3.321012, 3.256749, 3.479881, 3.457672, 2.702554, 
    2.815333,
  3.318106, 2.265729, 3.003447, 4.913236, 4.359295, 2.992944, 4.319507, 
    3.97901, 2.825653, 2.385048, 3.500928, 3.329794, 3.503647, 4.052084, 
    3.646657,
  5.23635, 4.588008, 4.616124, 4.995283, 6.020556, 4.952785, 3.213931, 
    4.148595, 5.496555, 2.947039, 2.358164, 2.857767, 3.056464, 3.91417, 
    3.395072,
  6.322681, 6.42601, 6.163143, 5.857523, 6.08138, 6.702093, 5.313141, 
    2.92154, 3.630798, 3.391545, 2.479411, 2.357944, 2.051855, 3.632978, 
    3.932232,
  6.993645, 7.262748, 7.259206, 7.104339, 7.125558, 7.489276, 6.862209, 
    4.749669, 4.354042, 3.721075, 1.950926, 2.125671, 1.200917, 3.153314, 
    4.776194,
  7.371143, 7.819649, 8.312229, 8.760053, 8.971271, 8.602974, 8.007187, 
    6.857643, 6.425264, 5.089179, 1.251872, 2.215588, 1.127777, 2.770377, 
    4.798377,
  7.404276, 8.14269, 8.951765, 9.792616, 10.20751, 9.861816, 8.982486, 
    7.671893, 7.249698, 6.502784, 2.976, 1.749632, 1.782964, 2.745982, 
    4.665901,
  7.357185, 7.915068, 8.591231, 9.332996, 9.790495, 10.08805, 10.19658, 
    9.66558, 9.10239, 8.302744, 5.989112, 1.396327, 2.467186, 2.916835, 
    4.229303,
  7.074299, 7.277792, 7.48632, 7.786295, 8.498025, 9.62723, 10.49227, 
    10.67502, 8.909922, 6.88395, 5.896163, 3.741861, 1.89032, 3.055609, 
    3.966806,
  5.137158, 6.365047, 4.707055, 5.01077, 4.281831, 3.216679, 2.936878, 
    2.35254, 2.161019, 2.249683, 2.839856, 3.677411, 3.540861, 3.200533, 
    2.7742,
  5.233267, 4.855487, 5.086246, 4.099685, 2.806047, 2.481276, 2.963236, 
    2.641284, 2.712123, 3.171139, 3.639381, 4.765402, 5.33513, 3.443403, 
    2.959581,
  4.328739, 2.721827, 4.080815, 4.449905, 3.564614, 2.416791, 3.341309, 
    2.939027, 2.398381, 3.060131, 4.074055, 4.831275, 5.787648, 6.081452, 
    4.269075,
  4.269543, 3.961187, 4.153632, 4.199409, 5.376405, 3.899087, 2.638022, 
    3.629593, 4.276242, 3.03948, 2.753759, 3.408386, 4.542792, 5.457705, 
    5.333923,
  4.603538, 4.682399, 4.736611, 4.117258, 4.694311, 5.424877, 3.902256, 
    2.674179, 3.301537, 3.381633, 3.233692, 2.820757, 3.53933, 4.339622, 
    5.664928,
  3.952327, 4.299052, 4.650633, 4.705749, 5.145071, 5.742414, 5.377385, 
    3.94045, 3.683973, 3.503963, 2.672848, 2.50108, 2.553194, 3.322163, 
    4.525619,
  3.320659, 4.008035, 4.623409, 5.383753, 6.14418, 6.055136, 6.190962, 
    5.670473, 5.241075, 4.605243, 3.293227, 2.152986, 2.117156, 3.150353, 
    4.610837,
  2.995064, 3.823109, 4.775092, 5.664287, 6.385307, 6.408453, 6.65487, 
    6.105189, 5.639097, 5.269191, 4.285251, 3.010025, 3.019356, 4.107893, 
    5.284472,
  2.612879, 3.232167, 4.212482, 5.075799, 5.768156, 6.415647, 7.239879, 
    7.22192, 6.749896, 6.029038, 5.627769, 4.51883, 3.658047, 4.286097, 
    5.043276,
  2.72939, 3.143926, 4.311642, 5.283004, 6.288626, 6.978086, 7.469135, 
    7.928956, 6.624732, 4.796696, 4.923618, 5.732574, 4.264913, 4.175828, 
    4.5286,
  3.768456, 4.621556, 3.378977, 3.269908, 2.310895, 2.13436, 3.195608, 
    3.693029, 3.643469, 3.378, 3.852706, 4.242917, 4.168421, 4.359154, 
    4.204696,
  2.600227, 2.53545, 2.866326, 3.120301, 2.764094, 3.197452, 4.72927, 
    4.981407, 4.978683, 4.22099, 3.457133, 3.703867, 3.640863, 2.786051, 
    2.984635,
  3.491566, 4.149375, 4.830566, 5.830877, 4.894716, 3.731752, 5.207658, 
    5.764956, 5.583993, 5.784593, 5.819061, 5.560789, 5.244434, 4.826178, 
    3.420279,
  4.922343, 6.101369, 7.080131, 7.426317, 8.547017, 7.302141, 5.381006, 
    5.306284, 7.23508, 7.611067, 7.475981, 7.192229, 6.704388, 6.476033, 
    5.7402,
  6.323097, 8.002919, 8.860147, 8.267013, 9.50502, 9.415774, 8.610518, 
    5.869024, 6.139829, 6.370485, 8.37359, 9.190074, 7.948299, 7.827123, 
    8.077088,
  8.956412, 9.948202, 9.384739, 8.391082, 9.618307, 10.27569, 10.90193, 
    10.69389, 9.00298, 7.137362, 6.74073, 9.319983, 8.810594, 8.542075, 
    8.372696,
  10.63777, 9.821877, 8.805327, 8.929187, 9.903095, 9.532039, 10.24756, 
    11.05608, 10.39455, 10.08818, 9.748589, 10.13, 9.633837, 8.942726, 
    8.371419,
  10.14092, 8.636889, 8.772447, 9.358495, 9.734528, 9.287442, 9.409169, 
    10.25744, 10.64065, 10.83538, 10.71886, 10.49794, 9.796032, 9.192084, 
    8.593546,
  8.477361, 8.1551, 8.916659, 9.266773, 9.245569, 9.1369, 9.978216, 11.21163, 
    11.39443, 10.82667, 10.52868, 10.09307, 10.05104, 9.512473, 8.381189,
  7.119902, 7.764457, 8.729387, 8.769807, 9.111691, 9.376992, 10.24539, 
    11.1869, 9.919512, 7.434291, 7.98271, 10.34896, 9.526193, 9.462411, 
    8.137463,
  3.349769, 4.781948, 4.717046, 5.013167, 3.261989, 2.457854, 3.671098, 
    4.209255, 4.3258, 3.576613, 3.602702, 4.256979, 3.584373, 2.944923, 
    2.806767,
  5.760389, 6.737896, 7.62235, 7.819958, 4.909075, 4.325331, 6.775561, 
    7.347939, 7.739737, 7.250622, 6.356989, 7.639456, 7.541894, 5.026417, 
    4.633189,
  8.281878, 8.610403, 10.01808, 10.16963, 6.40217, 4.395743, 5.415417, 
    6.689916, 7.469416, 7.880731, 8.462403, 9.33154, 10.23667, 10.53653, 
    7.301083,
  10.66541, 12.48549, 12.74699, 10.03253, 6.095386, 4.233013, 3.669071, 
    4.487644, 5.296177, 6.166537, 7.858568, 8.825026, 9.484912, 10.72883, 
    9.481247,
  12.37977, 13.99111, 12.72311, 6.185439, 5.253111, 4.966657, 4.742967, 
    3.806627, 4.555583, 5.132082, 7.390146, 8.832026, 8.841529, 9.601233, 
    11.49835,
  13.6906, 12.94321, 7.447946, 4.816825, 6.414325, 7.45016, 7.093992, 
    6.180014, 5.254102, 5.017708, 5.874152, 9.637832, 10.05476, 10.55991, 
    11.01712,
  12.9959, 8.698565, 5.31636, 6.240417, 7.628657, 5.924661, 5.745175, 
    6.349652, 7.157805, 8.426644, 9.544491, 10.83799, 11.82892, 11.95403, 
    11.78069,
  9.257873, 6.737713, 6.618832, 7.399226, 6.71425, 6.698296, 6.203581, 
    6.696828, 8.678884, 10.15802, 10.89472, 11.41223, 11.9355, 11.6193, 
    11.49109,
  7.692203, 7.296361, 6.88837, 6.502803, 6.612267, 5.939624, 7.215243, 
    9.500479, 10.82331, 11.54622, 11.15829, 10.40753, 9.86008, 9.696324, 
    9.089722,
  7.550208, 7.178907, 6.732379, 6.408842, 5.961302, 6.695157, 8.769803, 
    10.40981, 9.940824, 8.105594, 8.260255, 9.357061, 7.23542, 6.962642, 
    6.685326,
  3.381097, 5.654964, 6.567787, 9.298553, 9.583117, 7.233143, 7.301142, 
    5.416293, 4.925996, 3.710887, 3.49655, 3.454714, 2.38713, 2.163035, 
    2.307427,
  6.311053, 7.807475, 9.369683, 10.60509, 7.618958, 4.857646, 4.57462, 
    5.916036, 6.676645, 6.109573, 5.686225, 6.546392, 5.956516, 2.99464, 
    2.02417,
  8.943481, 9.336801, 10.85186, 11.84486, 6.266838, 2.941783, 4.966224, 
    5.168726, 5.327308, 6.461246, 7.389677, 7.836381, 7.723239, 6.880043, 
    4.36256,
  10.4014, 12.14177, 13.19997, 7.780651, 3.143768, 3.005662, 3.227947, 
    4.81672, 5.314606, 6.62155, 7.94249, 8.147317, 8.030183, 8.036681, 
    6.443399,
  11.20665, 12.60025, 9.636737, 4.194529, 5.549096, 4.158841, 3.17538, 
    3.065865, 4.498383, 5.635445, 7.897432, 8.305407, 7.847022, 8.197412, 
    8.676125,
  11.22621, 8.6589, 3.404835, 6.244145, 3.896364, 3.975118, 4.778515, 
    4.432303, 5.131704, 5.257406, 5.230126, 7.274816, 7.125096, 7.375922, 
    7.997086,
  7.596602, 3.164748, 5.119858, 2.559513, 3.639392, 3.247909, 5.36969, 
    6.934583, 7.439285, 7.136899, 6.762051, 6.816481, 6.960735, 7.268905, 
    7.922257,
  3.911257, 4.881298, 2.650887, 3.160273, 4.145364, 4.762133, 6.239089, 
    7.390624, 7.816797, 7.374683, 6.853887, 7.083786, 7.96844, 8.509641, 
    9.403666,
  6.452739, 4.044165, 3.170352, 3.628217, 4.683999, 6.195495, 7.920039, 
    8.785092, 8.255791, 7.401836, 6.569639, 7.192877, 8.812731, 9.52625, 
    8.968075,
  6.842703, 4.555626, 4.043464, 4.400224, 5.577618, 7.412194, 8.397295, 
    8.393729, 6.649351, 4.708823, 5.622563, 8.018125, 8.554915, 8.471377, 
    6.446541,
  4.877141, 6.097232, 5.26614, 6.321538, 6.279653, 5.822381, 8.285276, 
    6.905836, 4.762, 2.6403, 3.095186, 4.04387, 4.708833, 4.868396, 4.734977,
  7.524161, 7.491811, 7.396045, 7.681952, 5.045675, 4.749011, 6.357161, 
    4.619868, 2.878788, 2.92235, 3.790129, 5.210786, 6.148961, 4.922032, 
    5.360183,
  8.352903, 8.326014, 8.277662, 8.831391, 6.553121, 4.317513, 3.984531, 
    3.349994, 3.18241, 4.176192, 5.579005, 6.581509, 7.144022, 7.480835, 
    6.418639,
  8.025884, 9.111281, 9.704985, 9.341156, 7.699974, 5.22292, 2.379769, 
    2.522862, 3.469652, 4.617725, 6.160417, 7.330284, 7.71543, 8.112208, 
    6.710906,
  7.917638, 8.778609, 9.501494, 7.393722, 6.286183, 5.371848, 4.764415, 
    2.863457, 4.05484, 4.642933, 6.465098, 8.010402, 8.14242, 8.682849, 
    8.617391,
  8.192232, 8.730947, 8.03092, 6.850433, 5.970149, 5.019116, 4.834066, 
    5.218452, 5.019958, 4.698425, 5.417342, 8.489943, 8.868702, 8.937844, 
    8.790593,
  8.716963, 8.483632, 7.5194, 5.802631, 4.882894, 3.017133, 2.786722, 
    3.835255, 5.658218, 7.106773, 7.976122, 8.568663, 8.527312, 8.509609, 
    8.702507,
  9.174378, 8.057794, 7.344306, 5.772896, 4.660107, 3.839241, 3.408458, 
    4.690281, 6.78792, 7.406372, 7.036882, 7.200563, 7.750978, 8.29135, 
    8.990889,
  6.897754, 8.452795, 7.913337, 5.86986, 4.546245, 3.956599, 4.473063, 
    6.178144, 7.10669, 6.646144, 5.68856, 6.77549, 8.029216, 8.907675, 
    8.929192,
  7.330835, 7.723237, 7.000081, 6.152135, 4.359185, 3.78284, 4.488925, 
    6.136101, 5.670326, 4.192778, 5.025443, 7.133782, 8.040771, 9.142536, 
    8.789962,
  3.716071, 5.88463, 6.006604, 7.98495, 7.587369, 6.341441, 7.766815, 
    8.160785, 7.568537, 5.459877, 5.131597, 5.426785, 4.532355, 4.094138, 
    4.253998,
  5.24329, 6.412721, 7.369294, 8.018457, 5.774964, 4.754699, 7.756246, 
    8.103565, 8.005587, 7.239934, 5.941856, 6.528536, 6.597935, 4.59907, 
    4.348785,
  5.656244, 6.76145, 7.709749, 8.668441, 6.937169, 4.480491, 5.817256, 
    7.782506, 7.883132, 7.793018, 7.550595, 7.469329, 7.802547, 7.847431, 
    6.075355,
  5.904345, 7.450434, 8.942603, 9.935773, 10.24259, 7.482007, 4.291843, 
    4.370042, 6.020327, 8.112254, 8.448177, 8.363579, 7.996899, 8.147392, 
    7.199672,
  6.319826, 7.343106, 9.046626, 10.19127, 9.96945, 10.18134, 8.086107, 
    5.243581, 4.730884, 5.333842, 7.142734, 8.094687, 7.8167, 8.396537, 8.4989,
  6.492655, 6.775328, 8.21066, 9.540665, 10.04251, 9.723605, 10.32377, 
    9.899494, 6.612349, 3.826364, 3.82108, 6.068512, 6.364768, 6.796319, 
    7.46663,
  6.280407, 6.182994, 7.055225, 8.337295, 9.552208, 8.950044, 8.520253, 
    7.938957, 6.567246, 5.341694, 4.685809, 4.815875, 5.575642, 6.268142, 
    7.153998,
  5.427825, 5.324474, 5.915055, 7.121586, 8.398583, 7.697282, 7.515631, 
    6.843037, 5.143019, 4.380856, 4.503246, 4.97539, 5.474617, 6.517367, 
    8.539714,
  4.394516, 4.936242, 6.133009, 6.89051, 5.829907, 5.811954, 5.841555, 
    5.109279, 4.780968, 4.643316, 4.348553, 4.559, 6.019354, 8.162159, 
    9.677949,
  5.036506, 4.503013, 5.017933, 5.610029, 7.127327, 8.795297, 8.461867, 
    6.657609, 4.764401, 3.197883, 3.087732, 5.199017, 7.351007, 9.645195, 
    10.66413,
  5.279352, 7.398857, 6.188842, 8.062771, 7.384412, 6.053782, 7.648091, 
    8.288631, 8.20425, 6.49378, 6.804005, 8.064036, 7.63795, 7.05282, 6.772824,
  7.058001, 7.279212, 6.978424, 7.205485, 4.98578, 4.810221, 7.089266, 
    7.989904, 8.432391, 8.030289, 7.813762, 10.40615, 11.04038, 7.5378, 
    6.811099,
  6.494901, 5.353679, 5.699671, 6.06222, 5.026644, 4.067032, 4.666127, 
    6.030793, 7.697678, 8.366125, 8.606699, 10.12122, 11.47316, 10.60749, 
    7.66106,
  4.743029, 4.357486, 4.618295, 4.268599, 5.514885, 4.864006, 3.808489, 
    3.50191, 4.481721, 6.749999, 7.757684, 8.557752, 9.801394, 9.77701, 
    8.704462,
  3.808903, 3.942549, 3.423982, 3.490527, 4.009559, 5.299709, 5.992938, 
    4.41227, 2.82022, 3.897577, 6.652672, 7.689423, 8.315649, 9.381671, 
    10.69269,
  3.627918, 3.506987, 3.407693, 4.574921, 5.373312, 4.836806, 5.28457, 
    5.400009, 3.719802, 3.323335, 4.021486, 6.168681, 6.922062, 7.753381, 
    8.537244,
  4.698017, 4.154902, 4.503836, 5.863219, 6.716462, 6.398791, 5.475893, 
    4.459192, 4.093088, 4.260278, 4.475525, 4.340611, 3.771081, 3.58563, 
    3.553741,
  7.107863, 6.678009, 7.067274, 7.847039, 8.120215, 7.597869, 6.986395, 
    6.708508, 6.030072, 5.49147, 5.231965, 5.354787, 5.267434, 4.21556, 
    3.204587,
  9.936207, 9.538785, 9.461057, 9.49991, 9.224304, 8.845977, 8.577232, 
    8.59208, 8.706805, 8.615043, 8.193873, 7.180003, 5.174729, 3.652605, 
    3.261007,
  12.3043, 12.28582, 12.03778, 11.63656, 11.5283, 11.31019, 10.84826, 
    9.92223, 7.297513, 4.674092, 3.763805, 3.100143, 2.440162, 3.252425, 
    4.187578,
  6.218492, 8.260777, 7.567139, 10.05772, 9.331735, 7.956689, 10.04462, 
    10.36215, 9.886511, 6.80656, 5.966089, 6.206025, 4.847787, 4.316322, 
    4.269813,
  7.809103, 7.865151, 8.184283, 8.143619, 5.783537, 5.858934, 8.822469, 
    8.97148, 9.19402, 8.262157, 6.883191, 7.565322, 7.105604, 4.392684, 
    3.985159,
  8.104725, 7.068769, 6.936589, 6.905678, 5.111057, 4.487309, 6.026703, 
    6.670161, 6.462053, 7.014635, 7.159947, 6.657639, 6.806518, 6.189365, 
    4.763966,
  8.672322, 8.627823, 8.313741, 7.513737, 6.265177, 4.175173, 2.601961, 
    2.880095, 3.523701, 4.352267, 4.794472, 5.240045, 5.388599, 5.55148, 
    5.094715,
  9.136581, 9.135276, 9.152264, 8.647245, 8.171873, 6.483603, 4.242887, 
    2.361805, 2.102326, 2.239404, 2.76441, 3.162105, 3.471588, 4.040023, 
    4.841073,
  9.686349, 9.550535, 9.597262, 9.625074, 9.831469, 9.835409, 8.103793, 
    5.556935, 3.866637, 4.102674, 3.528312, 3.835112, 3.773268, 3.792274, 
    3.807334,
  9.788415, 9.762583, 9.8189, 10.12546, 10.50639, 10.78176, 10.80564, 
    10.32678, 9.85638, 9.656783, 9.128321, 8.752936, 8.135353, 7.325096, 
    6.461607,
  9.362477, 9.463734, 9.440029, 9.835176, 10.26302, 10.35559, 10.7943, 
    11.41951, 11.74155, 11.84751, 11.76143, 11.71607, 11.13553, 10.22344, 
    8.659704,
  8.695656, 8.449901, 7.894839, 7.623851, 7.91382, 8.273017, 8.725917, 
    9.532962, 9.831021, 9.316591, 8.962348, 8.676834, 8.06601, 7.225804, 
    5.845362,
  7.745787, 7.385979, 6.532128, 5.638867, 5.17563, 5.312193, 5.952312, 
    6.681969, 5.852228, 4.433482, 4.475496, 5.452068, 4.765945, 4.064925, 
    3.359379,
  2.730413, 4.298683, 4.452045, 6.290372, 6.833196, 6.636867, 8.539001, 
    9.283224, 8.920192, 7.171221, 8.035291, 8.92959, 8.18732, 7.723514, 
    7.607666,
  4.852492, 5.539942, 5.751392, 6.126348, 4.997643, 5.675241, 7.74816, 
    7.965709, 7.489945, 6.486352, 6.510343, 8.239676, 8.470304, 5.994435, 
    6.23617,
  7.478673, 6.252262, 5.831138, 5.713232, 4.794509, 4.870783, 7.029787, 
    6.773781, 5.414629, 5.624399, 6.198441, 6.811258, 7.305794, 7.550668, 
    6.175549,
  9.200929, 8.515507, 7.408032, 5.999131, 6.067992, 4.882903, 4.283884, 
    5.16574, 6.669788, 7.36276, 7.033288, 6.536077, 6.507965, 6.739386, 
    5.75983,
  10.21765, 9.162952, 7.95601, 6.241696, 6.041399, 5.712588, 4.481283, 
    2.848784, 4.439811, 5.795312, 7.51135, 7.447412, 6.749879, 6.244253, 
    5.848955,
  10.70724, 9.855535, 8.617102, 6.838993, 5.672985, 5.112078, 4.484664, 
    3.893818, 4.069847, 5.112128, 5.90446, 8.513177, 8.45834, 7.750915, 
    6.644266,
  10.69885, 10.30833, 9.058816, 5.969345, 6.84469, 4.891295, 3.90883, 
    4.625544, 6.074009, 7.38951, 8.170013, 8.576854, 8.77139, 8.739826, 
    8.261137,
  8.795982, 8.002669, 7.107451, 9.702911, 7.618424, 4.334849, 3.221849, 
    4.033188, 5.177459, 6.051948, 6.589668, 6.957914, 7.165312, 7.642409, 
    7.707292,
  8.148254, 8.37419, 11.77126, 12.32016, 7.767972, 4.243204, 3.340025, 
    4.170277, 5.036476, 5.578979, 5.758654, 5.902825, 5.982474, 6.492385, 
    6.54647,
  10.34008, 10.7223, 12.8397, 12.09335, 7.377153, 4.666506, 4.281938, 
    4.918084, 4.718578, 3.825527, 4.108209, 5.324973, 5.384952, 5.992739, 
    6.072619,
  2.023928, 3.256519, 3.667361, 5.161232, 5.158569, 4.398436, 5.937185, 
    6.433596, 6.398063, 5.082932, 5.166198, 5.826021, 5.516366, 5.21405, 
    5.270184,
  3.166847, 3.83606, 4.603246, 5.483035, 4.362402, 3.823222, 5.559821, 
    6.116671, 6.608421, 6.079669, 5.441498, 6.71223, 7.100056, 5.103991, 
    5.148989,
  4.861131, 4.962968, 5.345423, 5.83863, 4.70127, 3.551538, 4.440444, 
    5.991869, 6.200151, 5.771774, 6.118149, 6.795235, 7.298179, 7.175822, 
    6.022288,
  6.756408, 6.619703, 6.751022, 6.565979, 6.258886, 5.232737, 3.533093, 
    3.842737, 5.264035, 5.784602, 5.816951, 6.017201, 6.348107, 6.534168, 
    5.345121,
  6.755268, 7.083167, 7.726489, 7.699749, 7.188234, 6.805088, 4.581202, 
    3.138113, 3.27585, 3.684333, 4.703134, 5.243156, 5.256104, 5.81257, 
    6.067114,
  8.061091, 9.050199, 9.547561, 9.150732, 8.368183, 8.031854, 8.091585, 
    6.029166, 3.152646, 2.405059, 2.838741, 4.443328, 4.651592, 4.983613, 
    5.633725,
  11.79048, 12.35993, 12.62966, 12.96398, 12.93331, 11.88955, 8.587932, 
    5.930949, 3.718925, 3.321434, 3.943575, 4.029003, 3.835489, 4.26249, 
    5.053755,
  14.26106, 13.83113, 13.11605, 12.12137, 9.659561, 6.984595, 4.841742, 
    3.951305, 4.506318, 5.025992, 5.00833, 4.809124, 4.77358, 5.261751, 
    5.551317,
  13.21972, 12.3126, 10.64938, 8.721289, 6.595242, 5.387743, 5.311005, 
    5.931079, 6.518827, 6.493073, 6.552054, 6.84, 6.600441, 6.406583, 5.865828,
  10.04868, 9.035789, 7.652828, 6.198454, 5.610036, 5.912658, 6.556132, 
    7.657242, 7.044956, 5.603863, 6.329926, 8.364647, 7.545133, 6.93834, 
    6.078799,
  6.699501, 10.02985, 10.77024, 13.8799, 10.94565, 8.231762, 10.85701, 
    11.13067, 10.56882, 8.019631, 7.483054, 8.359339, 7.682897, 6.700788, 
    5.595259,
  9.108404, 10.6878, 12.8321, 14.14556, 11.57475, 10.28595, 12.21335, 
    11.41225, 10.90746, 9.569546, 7.971438, 9.216963, 9.035531, 6.058027, 
    5.371757,
  8.806067, 9.91919, 11.68054, 12.4943, 10.03939, 8.771832, 11.78661, 
    12.80958, 11.93629, 11.3143, 9.941688, 8.800355, 7.957819, 7.051359, 
    5.821899,
  7.575396, 9.172131, 10.39032, 10.70961, 9.904722, 7.073596, 6.504238, 
    10.318, 12.60715, 10.63876, 10.32425, 9.163946, 8.117757, 6.863415, 
    5.276506,
  7.511653, 8.579481, 9.441186, 9.639093, 8.818645, 7.371912, 5.735042, 
    5.232053, 5.06747, 5.369792, 7.609172, 7.194927, 6.354584, 5.43537, 
    4.787763,
  8.245001, 8.684514, 9.33623, 9.825264, 9.878939, 9.097858, 6.941346, 
    6.491057, 4.342207, 3.092962, 3.615374, 5.15697, 5.439825, 5.507167, 
    5.197381,
  5.93326, 6.184446, 6.419726, 6.566968, 6.747757, 7.159425, 6.955881, 
    5.283577, 3.306625, 3.943858, 4.885287, 5.929276, 6.801542, 7.440961, 
    7.615554,
  4.102269, 3.894984, 3.535352, 2.982111, 2.260982, 1.84542, 1.931828, 
    2.914172, 4.525929, 6.013017, 7.30837, 8.498918, 9.773647, 10.74596, 
    10.78892,
  5.320076, 4.987888, 4.688984, 4.301133, 4.352338, 5.328163, 6.081006, 
    6.833988, 7.777022, 8.740318, 10.25389, 11.52255, 12.39547, 12.74073, 
    11.85894,
  8.040432, 7.843603, 7.739113, 6.400361, 7.144625, 8.457851, 8.817469, 
    9.466858, 8.639012, 7.281658, 8.77114, 12.18526, 12.33147, 12.18993, 
    10.9528,
  6.926449, 12.27375, 14.04768, 17.96508, 9.362514, 3.356735, 5.343076, 
    7.448446, 9.015299, 8.289425, 8.311369, 8.829939, 8.247941, 6.688984, 
    5.311761,
  8.596939, 12.1743, 16.25671, 18.50144, 11.39791, 4.98357, 3.913612, 
    7.978913, 9.77195, 10.09135, 8.705906, 10.73315, 10.14178, 6.321767, 
    5.682052,
  9.099792, 11.0954, 14.37413, 17.16403, 12.70991, 6.802546, 5.493988, 
    7.349094, 10.76904, 11.2327, 10.7521, 10.84692, 10.34538, 9.583691, 
    7.940386,
  7.741561, 9.997177, 12.90167, 15.62731, 16.30569, 9.575233, 4.299725, 
    7.817464, 9.917912, 9.139556, 10.34698, 10.02863, 9.514692, 9.456431, 
    9.120317,
  6.010683, 7.303818, 9.979209, 12.3689, 15.63619, 15.48942, 8.922228, 
    5.622292, 5.28204, 5.660793, 8.984491, 9.61538, 9.760948, 10.09733, 
    10.2128,
  5.092283, 5.173232, 6.619413, 8.014247, 11.25803, 14.97628, 14.61213, 
    9.057079, 6.04258, 6.272152, 6.780329, 9.600322, 9.906316, 10.07637, 
    9.809115,
  6.263931, 5.266447, 4.287856, 3.072221, 5.067585, 8.921745, 11.89199, 
    12.16628, 10.36584, 9.853608, 9.269517, 9.802654, 9.842295, 10.21947, 
    10.33379,
  9.07042, 8.788432, 7.91859, 5.14671, 3.100112, 3.38141, 6.022742, 8.545395, 
    9.130862, 8.856745, 9.129297, 9.363003, 9.646588, 10.42999, 10.76287,
  12.21105, 12.98921, 12.61707, 10.6317, 8.688389, 6.734744, 4.574211, 
    5.245054, 6.781189, 7.255335, 7.603944, 8.594125, 9.373068, 9.874765, 
    9.678651,
  8.262482, 7.45354, 7.245455, 8.417222, 10.34507, 11.57305, 9.011393, 
    6.629673, 5.455518, 4.53375, 5.650297, 8.01076, 8.623528, 8.95739, 
    7.847092,
  3.7614, 5.416264, 5.879829, 9.602655, 12.44172, 8.079916, 4.446569, 
    2.795774, 3.231327, 3.23276, 4.533813, 5.333292, 4.998843, 4.228204, 
    3.913955,
  6.048334, 6.485603, 7.018987, 9.420158, 8.987215, 5.381797, 2.881387, 
    3.521544, 3.102229, 4.585931, 5.298749, 6.19052, 5.883113, 3.798962, 
    3.725809,
  6.629481, 6.224563, 6.413977, 8.188482, 7.747436, 4.658936, 2.034494, 
    3.138722, 4.557278, 6.389605, 6.748473, 6.000259, 5.694283, 5.623442, 
    4.990471,
  7.659088, 6.401256, 6.362383, 6.468809, 9.097452, 5.963131, 1.648032, 
    3.71556, 5.145907, 6.342779, 6.41697, 5.752365, 6.066769, 5.996162, 
    5.337361,
  8.782578, 6.66251, 5.545297, 4.44093, 7.604704, 9.118731, 3.160414, 
    4.82861, 4.172633, 4.090621, 5.51255, 5.828027, 6.240751, 6.074116, 
    6.311269,
  9.413311, 7.8647, 5.50071, 3.239861, 4.892034, 8.816462, 5.020744, 5.50523, 
    5.247863, 4.792101, 4.302744, 6.517119, 6.489888, 6.641144, 7.664474,
  9.860023, 9.180005, 7.182028, 3.848681, 2.325056, 5.488831, 6.253259, 
    5.23977, 6.819709, 7.058067, 6.511698, 7.116712, 7.198833, 8.228992, 
    9.9012,
  10.6469, 10.28075, 9.208417, 6.170085, 3.271909, 1.823803, 4.940078, 
    5.555861, 6.402454, 6.952536, 7.14187, 7.724471, 8.128371, 9.602488, 
    11.29666,
  10.63143, 10.24185, 9.453642, 6.605247, 4.818685, 4.099123, 3.379204, 
    4.998713, 5.536707, 5.604992, 6.944857, 8.109056, 8.921733, 10.44555, 
    10.55841,
  11.24035, 11.62121, 9.971588, 7.323823, 3.3014, 5.962692, 4.495204, 
    4.253775, 4.18349, 3.386153, 4.840205, 8.154481, 9.41072, 10.69779, 
    10.29821,
  5.954861, 7.372508, 5.443836, 6.301877, 4.24969, 2.896143, 3.248931, 
    2.206113, 2.902217, 1.342932, 1.352409, 2.735332, 3.69835, 4.085977, 
    3.836759,
  9.082234, 8.806593, 8.151716, 6.308257, 3.429083, 2.451253, 1.833603, 
    2.285528, 1.887809, 0.7843283, 1.379102, 3.229883, 5.193675, 3.861139, 
    3.729956,
  11.37474, 10.23582, 8.60186, 7.049553, 3.740357, 2.025737, 0.9158511, 
    1.341452, 1.466837, 1.237742, 2.514571, 3.913942, 5.348858, 5.920148, 
    5.73176,
  11.59492, 12.17432, 10.35664, 7.977229, 5.625549, 2.839925, 0.8107606, 
    0.9113466, 0.9526374, 2.089209, 3.840278, 4.721329, 5.72604, 6.577114, 
    6.630123,
  11.23475, 12.57381, 11.30675, 8.169507, 6.066802, 4.330575, 2.912696, 
    2.468521, 1.521814, 2.079396, 4.715918, 5.488698, 6.252747, 6.558113, 
    6.623132,
  11.18716, 12.51977, 11.91346, 8.710414, 6.467676, 5.599241, 2.921767, 
    3.727603, 2.809539, 3.416971, 4.150976, 6.275698, 5.920831, 5.761989, 
    7.523404,
  11.46542, 12.69534, 12.12515, 9.752422, 6.572253, 4.026724, 1.64241, 
    2.289578, 3.577638, 5.804459, 6.155358, 6.371515, 6.493234, 8.981426, 
    12.30402,
  11.71815, 13.1515, 12.67315, 11.31354, 7.330547, 2.84264, 1.400873, 
    3.714786, 4.645341, 6.557366, 6.876244, 7.438605, 9.667562, 13.3706, 
    13.91578,
  11.55522, 13.26301, 12.95784, 12.34397, 8.102937, 2.382027, 2.632094, 
    4.387681, 5.687434, 7.004736, 7.700405, 9.947825, 13.05869, 14.11721, 
    12.32745,
  10.3841, 11.9312, 12.47033, 12.80395, 8.852984, 3.893921, 3.938221, 
    5.270272, 5.381377, 5.207002, 7.162687, 12.10789, 13.43116, 12.87607, 
    11.32223,
  4.900963, 5.308014, 4.703533, 6.703769, 8.183158, 4.331439, 2.412306, 
    4.179758, 5.214477, 4.178637, 4.607205, 5.100274, 5.809648, 6.793358, 
    7.069689,
  7.057414, 5.426917, 5.021613, 5.793402, 6.064347, 3.771308, 2.565938, 
    3.662931, 4.894256, 4.381749, 3.938743, 5.43741, 7.576514, 6.191633, 
    7.196302,
  10.53851, 7.996851, 4.904456, 4.545931, 5.000851, 3.978018, 3.125626, 
    3.182744, 3.903961, 3.969655, 4.509861, 6.027673, 8.084514, 9.300667, 
    8.558343,
  11.18979, 10.61083, 8.42439, 5.586777, 6.047787, 4.809714, 2.466869, 
    3.159467, 5.532567, 5.193178, 5.35416, 6.90018, 8.979195, 10.38759, 
    10.0731,
  11.1211, 11.15661, 9.524488, 6.117795, 6.069551, 6.661215, 3.526954, 
    2.066236, 3.222182, 3.721336, 6.313526, 8.463223, 10.09519, 11.28714, 
    11.77997,
  10.80879, 11.38789, 10.42063, 7.451927, 6.334538, 6.41457, 5.76625, 
    4.440547, 4.017562, 4.85898, 5.912575, 9.965575, 11.2414, 12.49363, 
    13.09037,
  10.12915, 11.3519, 11.47967, 9.687855, 6.435893, 5.235565, 5.962829, 
    6.921439, 7.39897, 8.002995, 9.372372, 11.064, 12.38991, 13.16741, 
    13.25343,
  9.120262, 10.65645, 11.62754, 11.34165, 7.913357, 4.93718, 5.625947, 
    6.997928, 7.450372, 9.189251, 10.39232, 11.77244, 12.35902, 12.16436, 
    11.09466,
  8.169032, 9.579942, 10.64473, 11.54723, 9.201951, 5.04329, 5.051394, 
    6.379103, 8.181237, 8.760863, 9.934697, 11.24998, 11.0233, 10.22029, 
    8.876083,
  6.70822, 8.220192, 8.916462, 10.41554, 10.68534, 6.281641, 4.24401, 
    6.009867, 6.619737, 6.060287, 7.436767, 10.08617, 9.59558, 9.066276, 
    8.097672,
  4.15569, 5.220757, 5.832652, 8.278697, 6.893951, 5.3102, 7.052245, 
    8.118551, 8.3042, 6.244497, 6.43747, 6.909864, 4.447735, 2.800673, 
    1.860646,
  5.50771, 4.766739, 6.52172, 8.202251, 5.451418, 4.543163, 7.311135, 
    8.548594, 9.066199, 9.018328, 8.286896, 10.45642, 9.662517, 4.818551, 
    3.481284,
  6.830308, 5.624654, 6.360645, 8.096553, 5.68866, 3.87663, 5.522971, 
    7.877743, 9.081367, 10.27754, 11.14838, 12.71248, 13.39935, 11.71467, 
    8.276373,
  6.234872, 6.495163, 6.910457, 7.722161, 8.006001, 4.835666, 2.848227, 
    6.071673, 10.83496, 10.73334, 10.74005, 11.8617, 13.56396, 14.03915, 
    11.81215,
  5.450272, 5.82921, 5.776482, 5.787095, 7.039165, 7.757727, 4.50403, 
    3.316483, 4.963561, 6.045592, 8.990299, 10.29601, 11.55749, 12.59676, 
    12.67436,
  5.023657, 5.412645, 5.235502, 4.964688, 5.357789, 6.562976, 6.615752, 
    5.263433, 3.36465, 4.198753, 5.383499, 8.500986, 9.271973, 9.795913, 
    10.4387,
  4.707724, 5.248526, 5.508842, 4.834965, 4.626709, 5.153038, 5.286741, 
    5.662423, 5.908147, 6.206519, 6.238449, 6.844602, 7.322115, 7.494636, 
    7.651744,
  4.536314, 4.974341, 5.816924, 5.552305, 4.667476, 4.607123, 4.688547, 
    5.026202, 5.015625, 5.201132, 5.161439, 5.257002, 5.472457, 5.754834, 
    5.782894,
  4.866104, 5.031948, 5.625663, 5.835775, 4.995297, 4.283738, 4.746807, 
    4.552235, 4.203468, 3.906923, 3.898513, 4.001139, 4.154923, 4.624987, 
    4.811815,
  5.565936, 5.375542, 5.541885, 5.801471, 6.177599, 4.870497, 5.301524, 
    5.100564, 3.65181, 2.606859, 2.706017, 3.395961, 3.461683, 4.024002, 
    4.609127,
  4.488751, 6.087145, 5.533736, 7.433467, 6.801384, 5.956373, 8.154728, 
    8.722865, 8.854111, 6.971456, 6.915949, 7.270044, 5.288756, 3.84597, 
    2.041229,
  6.533156, 7.610296, 7.450725, 7.546472, 5.605305, 5.321685, 8.024883, 
    8.439001, 9.11004, 8.287993, 7.384586, 8.113754, 7.475264, 4.172941, 
    3.269105,
  6.977688, 7.961829, 8.195388, 7.943889, 5.915702, 5.24248, 7.329676, 
    8.113153, 8.125317, 8.056179, 8.165917, 8.205976, 7.707887, 6.288254, 
    4.178811,
  7.466661, 8.208101, 8.781422, 8.264216, 8.325502, 6.933171, 5.72655, 
    6.122144, 8.107431, 8.933128, 7.906032, 7.471612, 7.082344, 6.122005, 
    5.141019,
  8.141976, 8.473555, 9.035369, 8.408813, 9.414382, 9.856582, 8.482275, 
    5.897025, 6.188719, 6.343122, 7.704875, 7.33339, 6.632485, 5.517546, 
    5.365922,
  8.628342, 8.975595, 9.466785, 9.126837, 10.795, 12.02234, 12.14174, 
    12.02358, 9.543623, 7.095761, 6.389116, 7.71306, 6.698452, 5.328975, 
    4.305028,
  8.680593, 9.390144, 10.12327, 10.55982, 11.63668, 12.81289, 14.44653, 
    14.34187, 12.54002, 10.41873, 9.01278, 8.465728, 7.381705, 5.892504, 
    4.588767,
  8.857987, 9.610674, 10.49378, 11.22656, 12.44649, 13.58879, 14.83804, 
    15.00222, 13.02052, 10.53973, 9.209797, 9.073251, 8.296965, 6.515563, 
    4.985296,
  9.001642, 9.588625, 10.60221, 11.15771, 12.63092, 14.42981, 15.80052, 
    15.23647, 12.48432, 9.480052, 8.834542, 10.13869, 9.271288, 7.081638, 
    5.42928,
  8.438832, 9.094535, 10.24549, 10.68488, 12.79954, 15.30346, 16.55298, 
    14.65277, 10.13862, 6.464263, 7.552165, 10.57434, 9.018094, 6.990366, 
    5.480607,
  5.593488, 8.06286, 7.353003, 10.02815, 9.664703, 8.488304, 11.71885, 
    12.03023, 9.85885, 6.680262, 6.775606, 7.043602, 6.218967, 6.278816, 
    6.732489,
  8.172467, 8.538612, 9.196442, 10.2011, 8.038859, 8.284203, 12.21061, 
    13.30608, 12.0552, 8.497497, 6.280676, 6.756769, 7.155055, 5.556152, 
    5.909313,
  9.105819, 9.768388, 10.42836, 11.17774, 8.558034, 8.027821, 12.03327, 
    12.72849, 11.12329, 8.781956, 6.567148, 5.809264, 6.811903, 7.622413, 
    6.961539,
  8.965528, 10.04455, 11.28572, 12.16544, 12.30103, 9.669764, 8.60815, 
    11.43507, 13.54197, 9.441135, 6.70147, 5.04102, 5.259702, 6.987663, 
    8.056849,
  8.196916, 9.244289, 10.6824, 11.58403, 13.43045, 14.40753, 11.44786, 
    8.791684, 9.049562, 7.57456, 6.886267, 5.440176, 6.237312, 9.353239, 
    8.910859,
  7.407897, 8.559823, 9.975427, 11.39822, 13.56163, 15.05717, 15.34212, 
    13.34404, 8.886059, 6.991748, 5.594456, 6.578373, 9.016994, 10.57764, 
    8.530391,
  6.538937, 7.634353, 9.026264, 10.9165, 12.68798, 13.7793, 14.85872, 
    14.74787, 12.86884, 9.700654, 8.186818, 8.098665, 10.01342, 10.32489, 
    8.777458,
  5.787495, 6.809218, 8.118066, 9.884195, 11.67432, 12.70376, 13.63718, 
    13.78044, 12.78725, 10.70888, 7.977609, 8.710603, 9.749504, 9.157674, 
    8.061359,
  5.269555, 5.966418, 6.853259, 8.160256, 10.01572, 11.22683, 12.4088, 
    13.0089, 12.94326, 11.55725, 9.557902, 9.103176, 8.690768, 7.166345, 
    5.649909,
  4.977449, 5.340729, 6.205247, 7.293159, 9.122457, 10.01307, 10.69036, 
    11.07357, 9.85561, 7.936159, 7.320745, 8.521041, 7.118302, 5.625388, 
    4.025198,
  4.05439, 5.499039, 5.651557, 8.831993, 8.212473, 6.287442, 8.886549, 
    9.25975, 8.508864, 5.991523, 4.548458, 3.372696, 2.609318, 2.76133, 
    2.321473,
  5.643249, 6.315533, 6.924856, 8.465354, 6.519024, 5.843796, 9.188891, 
    9.960848, 9.774113, 8.122522, 5.549376, 4.816123, 3.481185, 2.288177, 
    1.782069,
  7.10793, 7.606851, 7.857297, 8.224813, 6.102499, 5.582763, 7.926403, 
    8.412895, 8.960748, 9.00797, 8.263024, 6.767416, 5.285684, 3.752728, 
    2.147972,
  7.641052, 8.206672, 8.647191, 8.327172, 8.016385, 6.209985, 5.370532, 
    6.72393, 9.714854, 10.12437, 9.313501, 8.36861, 6.934584, 5.40928, 
    3.621052,
  8.471297, 8.514209, 8.808757, 7.995518, 8.377095, 8.354856, 6.939215, 
    5.029393, 5.855522, 6.799616, 8.34349, 8.235311, 7.533815, 6.459296, 
    5.038871,
  9.421611, 9.02944, 8.87307, 8.359725, 8.910513, 8.904449, 9.017295, 
    8.905935, 7.194924, 6.012856, 5.699669, 7.285141, 6.700143, 6.026933, 
    5.4383,
  10.15445, 9.719569, 9.563461, 9.061027, 9.276185, 9.192432, 9.300815, 
    9.402899, 9.202537, 8.452343, 7.947373, 7.117301, 5.888076, 5.142167, 
    4.486298,
  10.80046, 10.35692, 9.833623, 9.575286, 10.14684, 9.872824, 9.430689, 
    9.196363, 9.071821, 8.736063, 8.310905, 7.046378, 5.461505, 4.314538, 
    3.453932,
  11.57847, 11.30082, 10.58282, 10.18393, 10.61803, 10.48992, 10.08308, 
    9.659781, 9.078125, 8.085342, 8.039546, 7.273574, 5.488567, 4.250993, 
    3.259363,
  12.09172, 11.57831, 10.83687, 10.64499, 10.69644, 10.58293, 10.2215, 
    9.640037, 7.929002, 5.526898, 5.922418, 7.167124, 5.446254, 4.178081, 
    3.46633,
  7.876667, 10.51197, 8.807687, 10.17775, 8.795548, 6.714339, 8.529855, 
    9.469645, 9.228305, 7.822615, 8.514099, 8.636744, 6.99633, 5.515326, 
    4.507407,
  11.35686, 12.06196, 11.50532, 10.1993, 5.83861, 4.948026, 7.908394, 
    8.273156, 7.99271, 8.555492, 9.073599, 10.9148, 10.26999, 6.548621, 
    5.012214,
  11.36891, 11.41677, 11.23619, 10.42671, 6.02451, 4.494877, 6.181764, 
    7.330166, 7.256877, 8.011367, 9.732965, 11.47789, 12.26941, 10.9426, 
    7.218622,
  11.98131, 11.79725, 11.37602, 10.54894, 8.764813, 5.473118, 4.416515, 
    4.996928, 6.140122, 7.414011, 9.207355, 10.81819, 11.92515, 11.2763, 
    8.365538,
  12.21201, 11.6743, 11.30488, 10.36834, 9.421535, 8.048417, 6.095859, 
    4.319929, 4.738457, 5.230673, 8.00718, 10.0831, 11.24082, 11.75906, 
    10.53156,
  12.15128, 11.38709, 10.73851, 10.21424, 9.45735, 9.190211, 8.581426, 
    7.563458, 6.27125, 5.638865, 5.970404, 9.458275, 10.32862, 10.7194, 
    9.964663,
  11.70484, 10.92586, 10.22726, 9.756738, 9.354618, 9.187424, 9.354053, 
    9.626579, 9.429798, 9.054906, 8.720992, 8.838733, 8.521822, 10.48119, 
    9.859196,
  11.24429, 10.45224, 9.626987, 9.235958, 9.175964, 9.312007, 9.186576, 
    9.557216, 10.17597, 10.57995, 9.589372, 8.504317, 11.70327, 12.10366, 
    9.23213,
  10.89376, 9.908236, 8.933686, 8.487325, 8.622918, 8.95496, 9.398642, 
    9.882589, 10.51005, 10.62039, 9.434822, 12.06434, 13.90866, 11.18946, 
    7.548073,
  10.32333, 9.212391, 8.353323, 8.862226, 9.199131, 8.993453, 8.984384, 
    9.182862, 8.47204, 6.977021, 7.921102, 12.17805, 10.95012, 8.179531, 
    5.545743,
  6.471545, 8.354462, 7.033316, 8.322896, 6.837212, 4.690313, 5.833926, 
    5.816845, 5.012103, 4.214959, 5.074752, 5.933212, 6.838181, 7.580469, 
    7.718194,
  9.209978, 8.81733, 8.591742, 7.584839, 4.965464, 4.200938, 5.852379, 
    6.105105, 5.823089, 5.156921, 4.993867, 6.163682, 7.285954, 6.869452, 
    7.424492,
  9.402581, 8.637018, 8.054487, 6.757031, 4.509642, 3.92842, 5.496034, 
    5.151974, 4.958455, 6.046637, 6.677182, 6.199225, 6.840617, 9.146613, 
    8.264415,
  9.526074, 8.771851, 8.060595, 6.571509, 5.373141, 4.288056, 3.694878, 
    4.768753, 6.574939, 8.006137, 8.507703, 7.075112, 5.796536, 7.444214, 
    8.59991,
  9.911901, 8.679172, 7.986476, 6.350246, 5.637116, 5.712099, 4.76186, 
    3.332533, 4.708402, 6.586174, 9.202026, 8.32281, 5.863571, 6.210266, 
    9.682719,
  10.30013, 9.026123, 7.889543, 6.733202, 6.244021, 6.051563, 6.182519, 
    5.311611, 4.439581, 4.981909, 6.236722, 8.791049, 6.647761, 3.911378, 
    5.104253,
  10.49735, 9.531001, 8.390411, 7.412739, 6.818542, 6.319212, 6.40119, 
    6.141756, 6.156184, 6.946125, 8.543134, 9.534191, 8.572868, 7.609184, 
    8.585183,
  11.0606, 10.19154, 9.228089, 8.228224, 7.308575, 6.694461, 6.594733, 
    6.440218, 5.85102, 6.04248, 7.033429, 8.285522, 9.901028, 10.95464, 
    10.80439,
  11.3715, 10.73739, 9.759086, 8.708261, 7.616619, 7.087141, 7.076797, 
    6.9388, 6.374691, 5.542613, 5.470099, 5.744291, 5.992554, 6.365892, 
    6.123429,
  10.95901, 10.48842, 10.15837, 9.588516, 7.976598, 7.287607, 7.783485, 
    7.875065, 6.896825, 5.089215, 4.323542, 5.1778, 4.482603, 4.221744, 
    3.855775,
  8.886944, 11.23397, 9.044133, 8.287483, 4.11628, 2.845541, 3.89294, 
    4.779144, 4.444775, 2.942602, 2.477704, 2.983084, 2.58762, 1.783648, 
    3.506462,
  12.56162, 12.52314, 11.71357, 9.033828, 3.708484, 2.588165, 4.354779, 
    4.866256, 5.002882, 4.213793, 3.619086, 3.956537, 3.215575, 1.888296, 
    2.531859,
  12.64713, 11.96731, 11.21366, 9.674581, 4.89374, 2.714203, 3.548989, 
    5.146468, 5.656065, 5.235523, 5.323958, 5.427471, 4.596286, 3.938587, 
    3.116015,
  13.10595, 12.53059, 11.56991, 10.04478, 7.428977, 4.370364, 2.482666, 
    2.389452, 4.191025, 6.367186, 6.550302, 6.176183, 5.222133, 4.345975, 
    4.154614,
  13.76225, 12.50482, 11.24753, 9.760297, 8.153539, 6.516434, 4.637578, 
    3.064593, 3.296997, 4.299376, 5.708221, 6.362148, 5.457904, 4.326061, 
    5.431409,
  14.37421, 12.31032, 10.68272, 9.351507, 8.254795, 7.351451, 6.544735, 
    6.396448, 4.789531, 3.485084, 3.552557, 5.476594, 5.523129, 4.766326, 
    4.498114,
  14.67574, 12.56475, 10.38744, 8.737782, 8.247668, 7.472528, 6.721631, 
    6.458539, 6.107975, 6.035869, 5.728198, 5.190442, 5.213181, 5.124749, 
    3.406827,
  14.73722, 12.56262, 9.692386, 8.171042, 8.359533, 7.773421, 6.710371, 
    6.434093, 6.810291, 7.352857, 7.357646, 6.488923, 5.256828, 4.586759, 
    4.026456,
  14.7042, 11.99566, 8.381892, 6.735209, 7.277021, 7.52939, 7.24344, 
    7.086017, 7.231136, 7.827792, 8.736023, 8.77392, 7.282205, 5.692508, 
    4.119646,
  13.10729, 10.66675, 6.90357, 5.699414, 6.750176, 7.415307, 7.480627, 
    7.407702, 6.489807, 5.566195, 6.979995, 9.7927, 8.659669, 7.253363, 
    5.335776,
  8.735644, 10.40433, 7.405, 8.908333, 7.258971, 4.754297, 5.262037, 
    5.105028, 5.234237, 4.551244, 4.204492, 3.595767, 2.525035, 1.923848, 
    1.682624,
  12.02994, 10.71605, 8.755972, 8.29305, 5.928795, 5.021801, 6.508492, 
    5.939787, 5.725978, 5.330823, 5.157833, 6.111233, 4.813625, 2.419232, 
    1.363088,
  11.50717, 10.22494, 8.676508, 7.48851, 6.210741, 5.366949, 6.670069, 
    6.156997, 6.170626, 6.580809, 6.639017, 7.100982, 7.643258, 5.689656, 
    2.952108,
  11.46724, 10.40241, 8.786702, 7.396243, 7.685075, 6.057148, 5.018999, 
    4.97524, 6.751382, 7.988094, 8.184909, 7.93961, 8.139157, 8.479893, 
    6.232254,
  11.671, 9.830035, 8.394338, 6.874412, 7.882476, 8.252765, 6.418165, 4.4721, 
    4.927631, 5.918146, 7.597567, 7.983165, 7.549824, 8.042828, 9.345209,
  11.78092, 9.768629, 7.882009, 6.917819, 8.163097, 8.51563, 7.89732, 
    6.130666, 4.361438, 4.902651, 5.124476, 6.967165, 7.32582, 6.98919, 
    7.667581,
  11.10363, 9.64821, 7.662778, 7.101743, 7.970222, 8.271297, 7.969742, 
    7.757124, 7.191893, 7.274165, 7.555294, 7.614722, 7.340298, 7.316772, 
    6.47155,
  10.48746, 9.351181, 7.708759, 7.461562, 8.023391, 8.139438, 7.661125, 
    7.34929, 7.346257, 7.52963, 8.037963, 8.56827, 8.322143, 7.637168, 
    6.725583,
  9.743064, 8.521679, 7.234226, 7.126099, 7.326521, 8.153402, 8.045933, 
    7.668775, 7.249084, 7.237519, 7.523588, 8.164729, 8.592405, 8.148974, 
    6.795491,
  8.514677, 7.10219, 6.431729, 6.778811, 7.510027, 8.326104, 8.19096, 
    8.02453, 6.719144, 4.883125, 5.325156, 7.469192, 7.969676, 8.308082, 
    7.116552,
  4.895745, 6.619992, 6.856863, 8.606681, 7.089405, 6.22975, 8.424249, 
    9.214838, 10.15913, 8.027913, 7.632987, 7.492661, 4.841619, 2.975988, 
    1.980081,
  7.04321, 6.728611, 8.133873, 8.431044, 5.698224, 5.186177, 8.077895, 
    8.893528, 10.03564, 10.38888, 9.247399, 9.462342, 7.881031, 4.11244, 
    2.656034,
  7.801558, 7.639779, 8.250813, 8.168321, 6.354294, 4.878517, 6.645821, 
    6.815059, 7.716058, 9.852848, 11.24086, 11.10969, 8.99471, 7.607923, 
    4.33582,
  7.982491, 7.794591, 7.729874, 7.09739, 7.726202, 5.639592, 4.536414, 
    6.004493, 8.43394, 8.878334, 9.625147, 10.59704, 10.09329, 8.291101, 
    6.243723,
  8.100611, 7.727673, 7.345656, 6.141373, 6.795271, 6.728909, 5.673229, 
    4.120403, 5.228672, 6.410332, 8.001139, 8.639421, 9.446372, 8.976495, 
    7.156723,
  8.595629, 8.020708, 7.385828, 6.71996, 7.242015, 6.355734, 6.798099, 
    6.344288, 5.431177, 5.034659, 4.890437, 6.919161, 7.861528, 9.302105, 
    7.718401,
  9.144824, 8.435331, 7.563068, 7.229502, 7.492734, 6.901594, 7.385154, 
    7.515635, 7.119051, 6.513867, 6.299146, 6.182454, 6.536656, 7.795881, 
    9.870391,
  9.701232, 9.103498, 8.285733, 7.628793, 8.133608, 7.963315, 7.711889, 
    7.26615, 6.722321, 5.88064, 5.554147, 5.234489, 5.438498, 6.872614, 
    9.477059,
  10.03615, 9.359219, 8.551148, 7.107073, 7.465578, 8.574001, 8.705123, 
    8.193077, 6.726885, 5.235723, 4.611546, 4.463654, 4.291228, 5.830158, 
    8.056696,
  9.924532, 9.0684, 8.654039, 7.557353, 7.867325, 9.289444, 9.185931, 
    8.41406, 5.934314, 3.373283, 3.433856, 3.979964, 3.195274, 4.600444, 
    7.048283,
  6.943941, 9.45974, 8.265703, 10.31325, 8.576743, 6.090276, 7.888267, 
    6.427649, 4.57967, 3.08284, 3.894108, 6.299458, 6.90445, 5.709614, 
    3.366674,
  11.0456, 10.24206, 9.575996, 8.902641, 5.487318, 5.145285, 8.006429, 
    6.663682, 5.074492, 3.547152, 2.490617, 5.209481, 7.092147, 5.008973, 
    4.21649,
  12.27701, 11.29246, 9.815669, 7.320168, 5.241891, 4.045168, 6.065686, 
    6.59969, 5.958681, 4.488541, 3.029002, 2.84817, 5.563114, 6.504182, 
    5.657956,
  12.43608, 11.44182, 9.524088, 6.375175, 5.756579, 4.331347, 3.903757, 
    4.169518, 4.98556, 5.510732, 4.630979, 2.324742, 3.166033, 5.74716, 
    6.535131,
  12.23096, 11.18995, 9.054278, 5.294122, 4.680415, 4.274677, 5.317487, 
    4.064439, 3.699226, 4.144971, 5.40584, 4.124956, 1.940109, 4.026444, 
    7.023339,
  12.24718, 11.26856, 8.990433, 5.431946, 4.181664, 2.432795, 3.850813, 
    5.787661, 4.302445, 3.391382, 4.134708, 5.304479, 3.131647, 2.454464, 
    5.850441,
  12.32659, 11.57489, 9.564316, 6.566139, 4.096422, 2.284784, 2.507053, 
    3.959004, 4.323151, 4.345227, 5.589909, 6.10781, 4.268013, 1.927874, 
    4.621753,
  12.41912, 12.02537, 10.58258, 8.057496, 5.811327, 3.580263, 4.092482, 
    4.430723, 4.392878, 3.934225, 5.113002, 6.407794, 4.866919, 1.954516, 
    4.152006,
  12.21307, 11.9075, 10.90142, 8.502921, 6.533328, 4.927823, 4.691582, 
    4.814841, 4.196366, 3.594224, 4.854043, 6.482013, 5.073493, 2.026823, 
    3.65446,
  11.67108, 11.33895, 11.38265, 10.04674, 8.083236, 6.342342, 4.495068, 
    4.129875, 3.698045, 2.963322, 4.07108, 6.478892, 4.651683, 1.874066, 
    3.597867,
  6.235058, 7.310905, 6.322994, 8.187187, 8.648587, 7.031651, 6.724217, 
    8.183472, 8.773394, 6.102549, 3.747475, 2.805973, 3.668271, 3.562579, 
    3.068126,
  11.10532, 9.420387, 8.206757, 8.221266, 6.00788, 3.621668, 3.828984, 
    8.286696, 9.937363, 7.573442, 4.176386, 3.173924, 4.217481, 3.361649, 
    3.121175,
  12.1377, 11.25266, 10.23205, 7.492525, 4.116024, 2.899827, 5.704461, 
    10.42644, 11.13022, 7.786112, 4.788429, 3.158921, 4.824502, 4.890994, 
    3.702994,
  12.37492, 11.48817, 9.805054, 6.103563, 5.480298, 3.901076, 5.759575, 
    8.637135, 7.95506, 6.062168, 4.377696, 3.07881, 4.804433, 4.750496, 
    3.881448,
  12.4789, 11.39116, 9.183859, 4.951307, 4.113454, 3.886304, 6.623165, 
    6.529733, 4.252656, 4.134331, 4.129059, 3.395496, 4.693578, 4.883433, 
    3.901873,
  12.59293, 11.82133, 9.792376, 6.07578, 3.671856, 3.42732, 5.193328, 
    8.966925, 6.062925, 4.971031, 3.578078, 4.069685, 4.409632, 5.009241, 
    4.361728,
  12.58959, 12.60588, 11.40217, 8.448568, 5.102826, 4.122042, 5.187008, 
    8.251019, 8.061745, 7.293776, 5.937484, 5.035676, 4.607326, 4.907867, 
    5.497127,
  12.26801, 13.1051, 12.99335, 11.47725, 8.531289, 7.438081, 9.511434, 
    9.879354, 8.728963, 7.552365, 6.387392, 5.674956, 5.0727, 5.228567, 
    5.906221,
  10.8958, 12.09889, 12.28382, 12.00942, 11.01879, 10.00051, 9.82144, 
    9.092261, 7.788741, 6.813842, 6.331918, 6.249318, 5.655723, 5.537612, 
    5.319595,
  7.923519, 9.590316, 10.43369, 10.57411, 10.16294, 9.341429, 8.353385, 
    7.968114, 5.99972, 4.429864, 4.850245, 6.5389, 5.900251, 5.826276, 
    5.253123,
  5.1829, 5.561595, 5.411452, 9.047524, 10.58254, 7.267153, 7.084814, 
    6.204123, 5.429786, 3.580496, 7.186674, 8.852221, 8.070936, 6.214831, 
    4.179255,
  8.722227, 7.078452, 7.125458, 9.215744, 7.991054, 5.863528, 3.530707, 
    6.452127, 6.007947, 6.294598, 8.150336, 9.639408, 9.191658, 5.131351, 
    3.750796,
  8.848653, 8.399355, 9.380424, 9.748466, 8.230823, 6.312757, 6.295262, 
    6.664488, 7.484307, 8.322175, 9.513011, 8.73648, 7.533957, 6.433614, 
    4.592819,
  8.241585, 8.027596, 8.960412, 9.949958, 10.99567, 8.207698, 5.804432, 
    8.760221, 10.0094, 8.827831, 8.263949, 6.25483, 5.898805, 5.947799, 
    5.101046,
  7.662321, 7.184024, 7.90002, 8.65556, 10.38734, 10.48519, 7.373779, 
    5.015408, 5.36179, 5.069868, 5.053619, 4.01431, 4.741367, 5.384888, 
    5.963712,
  7.518757, 6.884744, 7.232691, 8.182008, 9.273029, 9.709245, 9.204886, 
    6.734554, 3.100603, 2.420022, 2.155753, 3.516844, 4.203985, 5.267178, 
    5.899731,
  7.827893, 7.661288, 7.449476, 7.648603, 8.08998, 8.003314, 7.721817, 
    6.689058, 4.945522, 3.094506, 3.157206, 3.894297, 4.18539, 5.918336, 
    6.327093,
  7.482641, 8.09177, 7.933784, 7.506267, 7.501739, 7.397828, 6.797164, 
    5.63697, 4.443689, 4.313993, 4.155162, 3.732513, 4.876189, 6.324624, 
    6.301627,
  6.563354, 7.403, 7.353052, 7.014168, 6.762234, 7.141145, 6.969525, 6.33912, 
    5.495527, 4.935384, 4.18118, 4.774114, 5.900884, 5.866412, 4.83525,
  4.857814, 5.868044, 6.107352, 6.404912, 6.380527, 7.046111, 7.408241, 
    7.521377, 6.060873, 4.63544, 4.822312, 6.437052, 5.897691, 5.106303, 
    3.478458,
  2.536837, 2.958106, 4.334505, 9.825414, 11.70893, 10.22899, 13.24324, 
    11.39979, 7.549855, 4.713545, 4.337368, 5.279008, 7.018151, 9.472269, 
    9.110688,
  3.229115, 3.598338, 5.543311, 9.347168, 8.411202, 8.729715, 13.83974, 
    14.43968, 11.86727, 10.85622, 8.453197, 10.08899, 12.92663, 9.077103, 
    8.139907,
  4.057111, 4.604789, 7.34861, 9.231394, 8.07529, 6.820337, 11.07372, 
    15.35523, 16.2486, 15.96297, 15.96411, 16.46889, 14.10901, 11.26587, 
    8.613203,
  4.889728, 5.19251, 6.982358, 8.666441, 10.29051, 7.635639, 5.681685, 
    10.98351, 16.86323, 15.65166, 14.31086, 14.11877, 13.32953, 11.21517, 
    8.115137,
  5.734564, 5.52082, 6.299926, 7.032328, 8.972573, 9.904155, 7.028701, 
    5.327661, 7.248883, 8.35474, 10.46104, 10.58777, 10.40375, 10.22351, 
    8.837163,
  6.8184, 6.286572, 6.621483, 7.042805, 7.57173, 7.785417, 7.521772, 
    4.981303, 2.792164, 3.452803, 4.513565, 7.202951, 7.655639, 7.496092, 
    7.389325,
  7.329075, 7.403028, 7.612999, 7.606234, 7.196562, 6.355442, 4.981586, 
    4.136737, 3.685344, 3.382688, 3.345666, 4.284927, 4.954238, 4.900643, 
    5.132349,
  6.683897, 7.548498, 8.226637, 8.490789, 7.984772, 7.063184, 5.225284, 
    3.615729, 2.915323, 2.117281, 2.170902, 2.665555, 3.056998, 3.500978, 
    3.899722,
  5.809824, 6.717765, 7.467141, 8.34832, 8.727608, 8.294522, 6.685644, 
    3.893833, 3.244611, 3.503972, 3.74928, 3.758724, 3.685271, 3.51516, 
    3.494512,
  4.129466, 5.069407, 6.225089, 7.44302, 9.139974, 10.61569, 9.898829, 
    7.044361, 2.9695, 1.421431, 2.033344, 2.881837, 3.231454, 3.169063, 
    3.064118,
  2.970157, 5.221294, 5.853499, 8.900648, 8.718477, 7.359936, 10.8585, 
    12.64284, 13.04369, 9.837622, 5.904964, 3.931762, 3.623036, 4.55709, 
    4.276134,
  5.15133, 5.40995, 6.540275, 8.229134, 6.661727, 6.478346, 10.01539, 
    11.44299, 12.33919, 12.71007, 9.819398, 4.320601, 3.939177, 3.556392, 
    4.049606,
  6.427784, 6.814312, 7.30449, 7.571208, 6.080245, 5.741426, 9.006838, 
    9.229313, 9.37404, 11.88493, 13.99657, 8.974895, 3.864969, 5.305141, 
    4.96908,
  6.495484, 6.813895, 7.22067, 6.925536, 7.429324, 6.044141, 6.121865, 
    7.86651, 9.985341, 10.48855, 12.73729, 13.71039, 5.59446, 6.285543, 
    6.042218,
  6.154293, 6.505091, 7.011546, 6.204633, 7.556765, 8.111288, 6.76138, 
    5.248099, 6.122297, 6.78222, 9.676294, 11.55824, 9.80412, 6.003584, 
    6.861887,
  5.62944, 6.411924, 7.180392, 7.277688, 8.032253, 8.673295, 8.376656, 
    7.515834, 5.955343, 4.635493, 5.027839, 8.875822, 9.428161, 6.764446, 
    6.939703,
  5.645917, 6.850403, 7.557318, 7.343288, 7.730765, 8.591178, 9.377913, 
    9.209237, 7.160835, 5.044592, 4.840361, 6.573628, 7.729285, 6.839534, 
    6.109477,
  6.65989, 7.709863, 7.695125, 6.881804, 7.189578, 8.283884, 9.183159, 
    8.906203, 6.871612, 4.447245, 3.475779, 4.514612, 5.870365, 6.069664, 
    5.009976,
  8.240059, 8.058333, 6.434917, 5.593608, 6.124615, 7.222778, 9.189708, 
    9.310699, 7.496634, 4.291308, 2.433782, 2.89624, 4.270532, 4.774659, 
    4.343502,
  8.684676, 6.694614, 4.588715, 5.026778, 5.020778, 6.410869, 8.89188, 
    9.454918, 6.872541, 3.188787, 1.442309, 1.670923, 3.032173, 3.743527, 
    3.560758,
  6.173068, 8.79357, 7.616009, 8.803557, 7.916435, 6.851763, 9.055634, 
    8.361834, 7.268116, 6.066, 6.571813, 5.267171, 5.077105, 6.519026, 
    5.646587,
  9.396643, 9.272593, 8.396758, 8.051475, 5.948367, 5.80017, 7.934275, 
    7.105532, 7.054904, 6.604858, 6.535429, 5.593249, 5.162566, 5.511367, 
    5.884459,
  9.301391, 8.736396, 7.901792, 7.400696, 5.44284, 5.181551, 5.818656, 
    5.901892, 5.258086, 6.349253, 7.552786, 5.904832, 4.244686, 6.127415, 
    5.903894,
  8.295926, 7.937299, 8.06512, 7.742296, 8.04239, 4.933505, 3.149324, 
    4.60916, 5.694965, 7.177332, 7.795706, 6.266413, 3.839393, 4.485296, 
    4.575484,
  7.345765, 7.233984, 8.147886, 8.205422, 8.558248, 5.239046, 3.374207, 
    2.480207, 4.113805, 5.425122, 7.320457, 7.012825, 4.12765, 3.217965, 
    2.985607,
  7.594079, 7.174893, 8.195435, 8.777102, 7.870663, 5.077738, 3.82998, 
    2.800831, 4.317341, 4.537219, 4.58999, 7.070213, 5.245402, 4.725518, 
    4.424105,
  7.663872, 7.69953, 8.42201, 7.922668, 5.873648, 4.800638, 3.667835, 
    4.647137, 5.38702, 5.459397, 5.720231, 6.827714, 6.6297, 4.885561, 
    4.794777,
  7.266692, 7.128932, 7.022614, 5.966534, 5.21353, 3.992558, 4.378045, 
    4.775366, 4.664177, 4.396028, 4.841867, 6.396028, 6.80131, 5.594558, 
    4.659537,
  5.835435, 4.894664, 4.317317, 4.069386, 3.76658, 3.720051, 5.888488, 
    6.018336, 4.646605, 3.480286, 4.167299, 6.180474, 6.686422, 5.492376, 
    4.3649,
  3.599001, 2.847361, 3.03203, 2.766639, 2.281169, 3.680812, 6.456867, 
    6.609024, 4.043956, 2.173705, 2.860455, 5.512537, 6.466372, 5.191157, 
    4.188747,
  3.563003, 6.094785, 6.079535, 7.614806, 6.803026, 4.910349, 5.467535, 
    3.63619, 2.995455, 2.16147, 1.957035, 3.973509, 4.665431, 5.032099, 
    5.697142,
  5.401812, 6.192305, 6.491637, 6.5568, 4.610427, 3.905142, 4.872532, 
    3.758277, 3.413956, 1.449859, 2.705306, 5.44357, 6.101377, 4.330386, 
    5.148079,
  5.089451, 5.517632, 6.016797, 5.730915, 4.406908, 3.524543, 4.164386, 
    4.291429, 2.527256, 1.908211, 4.41643, 6.385076, 6.991206, 6.972763, 
    5.503929,
  4.240266, 4.861509, 5.301196, 5.286963, 5.722898, 4.197026, 2.998682, 
    3.620545, 3.499388, 3.282726, 4.62465, 6.775009, 8.157595, 7.769153, 
    5.413695,
  3.685334, 3.800832, 4.332503, 4.270061, 5.265198, 5.792593, 4.049283, 
    2.31338, 3.200153, 3.654185, 5.512053, 7.482768, 8.788976, 8.344231, 
    6.335365,
  3.421201, 3.839141, 4.013798, 3.588358, 4.313582, 5.323528, 5.585064, 
    4.451697, 4.399086, 3.965338, 4.54741, 7.310833, 8.864064, 8.568578, 
    4.921539,
  3.257926, 4.00542, 3.719097, 3.365191, 3.617946, 4.699202, 6.560009, 
    6.674537, 5.875875, 5.377859, 6.271244, 7.415389, 8.665141, 7.29654, 
    3.559526,
  3.036424, 4.083029, 3.698086, 3.349074, 3.246821, 3.92893, 6.734908, 
    6.996368, 6.293121, 5.728782, 6.647537, 7.255539, 7.609257, 5.821623, 
    3.32221,
  3.642215, 4.509266, 4.171875, 3.633387, 2.939147, 3.36152, 6.903512, 
    7.873394, 6.866573, 6.339449, 6.980642, 7.138917, 6.771601, 5.117175, 
    3.891386,
  3.769895, 4.283587, 4.880465, 3.614789, 3.493482, 3.047562, 6.711556, 
    7.816908, 6.349886, 4.593127, 5.222155, 7.092693, 6.649602, 6.013025, 
    5.246552,
  2.371078, 3.733912, 4.346071, 5.979611, 5.337307, 4.309295, 5.382964, 
    5.942914, 5.225554, 3.554037, 3.07011, 3.302032, 3.33289, 3.462025, 
    4.054954,
  3.917878, 4.501789, 5.557296, 6.41396, 4.505875, 3.722063, 5.009765, 
    5.812255, 6.099825, 5.113291, 4.16575, 4.988424, 5.520399, 4.223361, 
    4.967197,
  4.242023, 5.838534, 6.597249, 6.389236, 4.047633, 3.093813, 4.26631, 
    4.965369, 4.955429, 5.49917, 5.700253, 6.180643, 7.262824, 8.366376, 
    7.709289,
  4.545258, 5.907902, 7.204455, 6.739122, 4.945326, 3.443665, 3.109119, 
    5.222024, 6.671719, 6.836798, 6.864665, 6.974563, 7.787764, 8.846927, 
    8.425855,
  4.289573, 5.857435, 7.693781, 7.009717, 5.448933, 3.882871, 2.821952, 
    3.55083, 5.533477, 6.467901, 8.031562, 7.936364, 8.308175, 8.684485, 
    9.080086,
  3.686425, 5.239581, 7.319218, 6.631006, 5.386438, 3.506557, 3.885471, 
    5.77241, 6.341922, 5.97755, 5.901773, 8.259695, 9.08991, 9.288792, 
    9.543114,
  3.030431, 4.75871, 6.603245, 5.492865, 5.258877, 3.381004, 5.39825, 
    7.580389, 7.783244, 7.797855, 8.439961, 9.138906, 9.669049, 9.507186, 
    9.983739,
  2.403503, 4.291116, 6.033339, 4.94511, 5.023834, 4.08532, 5.707613, 
    6.990878, 7.3129, 8.106365, 9.067719, 10.34414, 10.49541, 9.98974, 9.16099,
  2.360564, 3.596058, 4.608272, 4.738157, 5.196245, 4.808421, 6.260164, 
    7.137155, 7.133554, 7.88319, 9.65163, 11.53139, 11.79491, 11.28159, 
    10.22308,
  2.090449, 3.308274, 3.556895, 4.269173, 4.771663, 5.414181, 6.38715, 
    6.674364, 5.79044, 5.315067, 7.449688, 11.95324, 13.40151, 13.76692, 
    12.58605,
  3.025732, 4.388057, 4.43587, 6.158565, 6.068995, 4.720215, 4.802524, 
    4.532814, 5.112736, 4.784064, 5.313695, 5.677998, 4.857633, 3.786477, 
    3.463165,
  4.054319, 4.579547, 4.951855, 5.696508, 4.016025, 3.455048, 4.934821, 
    5.565336, 6.414419, 6.040285, 5.830867, 6.936924, 6.629276, 4.466505, 
    4.107855,
  3.99631, 4.03504, 4.583746, 5.262984, 3.924638, 3.005702, 4.733467, 
    5.968775, 5.798495, 7.031874, 7.954549, 8.154655, 7.660956, 7.082125, 
    5.832409,
  3.661305, 3.742556, 3.936947, 4.838178, 4.750074, 3.335555, 3.275144, 
    5.989672, 8.782182, 9.599318, 9.838425, 9.715942, 9.049025, 8.442188, 
    7.372284,
  2.903829, 3.336305, 2.903111, 3.840565, 4.125857, 4.823015, 3.981586, 
    3.894682, 6.202528, 8.322724, 11.12763, 11.12986, 10.17741, 9.283412, 
    8.885693,
  2.476856, 3.387957, 2.498515, 3.010643, 3.188865, 4.432409, 5.05173, 
    5.183895, 5.384218, 6.671309, 7.959475, 11.70122, 11.19615, 9.183167, 
    8.111078,
  2.800711, 3.902774, 2.481814, 2.693743, 2.802465, 3.996251, 5.169369, 
    7.271048, 9.004292, 10.6216, 12.13321, 12.79301, 11.90475, 9.684036, 
    6.712837,
  3.588108, 4.856163, 2.984513, 2.700518, 2.822259, 3.745628, 4.608013, 
    6.637572, 8.961761, 10.8448, 12.60944, 13.827, 13.20813, 11.39629, 7.36959,
  4.168775, 6.163915, 3.951787, 2.822731, 2.927082, 3.573743, 4.373223, 
    6.526174, 8.928462, 10.49414, 12.39498, 14.24655, 14.25113, 12.59605, 
    8.742614,
  4.523974, 7.502968, 5.530034, 3.4005, 3.168113, 3.824087, 4.088194, 
    5.99678, 6.928421, 6.311909, 8.069599, 13.61909, 14.85162, 13.68565, 
    9.90566,
  2.738188, 3.195323, 2.331898, 2.141834, 2.071858, 2.730647, 3.888318, 
    4.679889, 4.888758, 4.447911, 4.918025, 5.197059, 5.182657, 4.410162, 
    3.612194,
  4.304594, 3.149089, 2.736037, 2.306079, 2.02647, 2.770616, 4.15032, 
    5.094849, 5.765584, 5.457147, 5.227314, 6.845007, 6.220621, 4.234007, 
    4.082566,
  6.127538, 4.767773, 3.867992, 3.143522, 2.51317, 2.602523, 4.20604, 
    4.601324, 4.700732, 5.757039, 6.756876, 7.681459, 7.97559, 7.355861, 
    5.40379,
  6.994355, 6.244806, 4.939726, 4.32364, 3.976697, 3.063454, 3.225912, 
    4.915287, 6.313287, 6.49879, 7.287323, 8.606178, 9.019066, 8.890355, 
    6.45751,
  6.908587, 6.626612, 5.950408, 5.707299, 5.521937, 4.976511, 4.513053, 
    3.766098, 5.466892, 6.490436, 8.257224, 9.559442, 9.756136, 9.6872, 
    8.87927,
  5.915751, 5.97374, 5.949955, 6.388134, 6.758645, 6.782135, 7.02362, 
    7.633542, 7.616799, 7.325448, 6.668839, 9.744223, 10.40841, 10.3769, 
    10.03035,
  5.342714, 5.599019, 5.865134, 6.249621, 7.039826, 7.477186, 8.35737, 
    9.454986, 10.16669, 9.855739, 9.629251, 9.840277, 10.13583, 10.90863, 
    10.48546,
  4.460449, 5.200938, 5.940015, 6.589127, 7.645421, 8.503873, 9.437004, 
    9.72862, 9.990608, 9.831098, 9.603707, 9.250658, 9.825191, 11.19703, 
    10.85965,
  3.786772, 5.119436, 6.315629, 7.29679, 8.493991, 9.194346, 9.826562, 
    9.837547, 9.260954, 8.654163, 8.120065, 8.453798, 9.667005, 10.95417, 
    10.74997,
  3.904502, 5.437088, 7.099237, 8.511621, 9.24276, 9.741487, 9.275127, 
    8.365623, 6.901584, 5.247199, 5.190687, 7.463872, 8.782491, 10.63332, 
    10.37282,
  6.013389, 8.476631, 7.351713, 8.51762, 6.855712, 5.114303, 6.876598, 
    6.935609, 6.517407, 4.859675, 4.435352, 4.0676, 3.253159, 2.73225, 
    2.248256,
  8.568719, 9.08208, 8.472037, 7.805806, 4.487135, 3.876714, 6.387099, 
    7.153781, 7.877005, 6.5421, 5.551101, 5.671068, 5.181068, 3.572262, 
    3.096732,
  7.852459, 7.505268, 7.199591, 6.214971, 4.626069, 3.23074, 5.07914, 
    6.984967, 8.363592, 8.600634, 8.405166, 7.8968, 7.777942, 7.727328, 
    5.552744,
  5.96244, 5.009434, 5.342766, 5.415858, 6.192833, 5.753703, 3.891165, 
    5.152351, 7.305247, 8.017715, 8.602505, 9.020227, 9.16131, 9.501766, 
    8.203864,
  3.876865, 3.456378, 4.320911, 5.027984, 5.84309, 7.285038, 7.286936, 
    5.138441, 5.826635, 5.72197, 8.052115, 9.754173, 10.08442, 10.29293, 
    10.88973,
  3.196308, 3.539397, 4.200294, 5.128266, 6.357978, 7.887444, 9.266786, 
    9.952949, 8.456707, 7.391763, 7.327, 11.00797, 11.57, 11.21959, 11.22333,
  4.225796, 4.666916, 5.160499, 6.192811, 7.671842, 8.869426, 9.181289, 
    9.094543, 9.279971, 9.877098, 10.22251, 10.3864, 10.09944, 9.653162, 
    9.858718,
  5.150714, 5.214503, 6.114443, 7.501764, 9.21305, 9.017083, 8.210098, 
    8.424918, 8.883891, 8.749671, 8.093721, 7.947623, 7.876478, 7.913996, 
    8.179378,
  5.163098, 5.643075, 6.726101, 8.787704, 9.19486, 7.99867, 8.028957, 
    8.364094, 7.886926, 6.864199, 6.963026, 8.432964, 8.74322, 8.49611, 
    8.041276,
  5.039153, 5.961956, 7.953098, 9.680032, 8.387856, 7.625395, 7.243993, 
    7.254753, 6.565723, 5.668063, 7.163712, 9.870276, 8.610125, 7.34805, 
    6.512046,
  3.305653, 5.05236, 4.749658, 5.65913, 4.55979, 2.855164, 3.221373, 
    3.820244, 4.592036, 4.082492, 4.708769, 5.142577, 4.018793, 2.747689, 
    1.807998,
  5.370856, 5.805265, 5.716407, 4.880281, 2.806634, 2.581192, 3.941802, 
    4.850187, 6.1299, 6.362546, 6.244666, 7.18303, 6.952245, 4.258943, 
    3.233962,
  5.647549, 5.66663, 5.803102, 5.134507, 3.800853, 3.322821, 4.679233, 
    5.675139, 7.177587, 8.327398, 8.357808, 8.067593, 7.184076, 6.497176, 
    5.167887,
  5.083356, 5.431839, 6.173975, 6.68945, 6.695181, 5.039047, 4.006532, 
    4.684326, 6.635523, 7.582614, 7.436769, 6.415322, 5.003994, 4.699182, 
    3.708219,
  4.80651, 5.644809, 6.70753, 7.682263, 8.15573, 7.645029, 5.869618, 
    4.376675, 4.826858, 4.615758, 5.474711, 5.071968, 4.83328, 5.198473, 
    5.050274,
  4.839664, 6.023246, 6.896644, 7.765746, 8.088558, 8.147244, 7.48588, 
    5.480357, 3.655433, 3.656464, 3.532534, 4.402289, 4.405489, 4.604714, 
    5.087126,
  4.8221, 6.096343, 6.850808, 7.426653, 7.42874, 7.520417, 7.458199, 7.11461, 
    6.196774, 5.146813, 4.727796, 4.992702, 5.498092, 5.894016, 6.301614,
  4.645754, 5.75221, 6.432049, 6.950935, 7.135554, 7.225884, 7.115294, 
    6.729686, 6.40091, 6.179178, 6.139582, 6.434231, 7.024384, 7.411829, 
    7.509202,
  4.204123, 5.031547, 5.441083, 5.499443, 5.934556, 6.409206, 7.316316, 
    8.281115, 8.026512, 7.776756, 7.298759, 7.522512, 7.727033, 7.697262, 
    7.452783,
  3.708739, 4.266459, 4.275677, 4.348142, 4.803854, 6.135077, 7.940722, 
    8.551419, 7.861922, 6.113187, 6.496526, 8.237024, 7.675691, 7.386023, 
    6.761296,
  4.875767, 6.705606, 6.537482, 7.55252, 6.533724, 6.108841, 8.098567, 
    8.424724, 8.388987, 6.78152, 6.470866, 6.488017, 5.118647, 3.497231, 
    2.079739,
  6.399883, 7.047006, 7.97135, 7.884996, 5.497053, 5.254477, 7.859136, 
    8.599193, 8.935516, 8.340075, 7.392375, 8.327549, 7.177797, 4.139429, 
    3.219544,
  5.467566, 6.085273, 7.439791, 7.546352, 5.718279, 4.397051, 6.344525, 
    6.502168, 6.904, 8.013335, 8.331477, 8.805305, 8.33415, 7.086587, 5.038761,
  4.452192, 5.11412, 5.969694, 6.674297, 6.805243, 4.620148, 4.045507, 
    5.434025, 7.35536, 8.057937, 7.619534, 7.400272, 7.049309, 7.538748, 
    7.064248,
  3.758631, 4.320332, 4.77523, 4.965263, 5.68956, 6.403242, 4.952189, 
    3.693469, 4.965292, 5.747033, 7.083959, 6.831014, 5.671044, 5.122609, 
    5.897942,
  3.615899, 4.018199, 4.114876, 4.358974, 5.254575, 5.418808, 6.127492, 
    5.891308, 5.175908, 4.88869, 4.385783, 6.197071, 5.981263, 4.305419, 
    3.439274,
  3.771403, 4.067837, 3.753364, 3.725339, 4.726554, 4.862643, 6.060981, 
    7.145675, 7.411194, 7.125555, 6.551996, 6.369521, 6.328894, 5.095326, 
    3.143737,
  4.581096, 4.603666, 3.908756, 3.731379, 4.941289, 4.72991, 5.873226, 
    6.527219, 6.892147, 6.764876, 6.553473, 6.676883, 6.616212, 5.718946, 
    4.019164,
  5.490472, 4.828572, 3.811445, 3.949807, 5.051956, 4.468046, 5.750257, 
    6.887949, 7.484652, 7.699315, 7.136168, 7.119806, 6.631167, 5.915597, 
    4.389459,
  5.958161, 4.983526, 4.665157, 4.949707, 5.093077, 4.384046, 5.23619, 
    6.147687, 6.28604, 5.252695, 5.480661, 6.862422, 6.145115, 5.778605, 
    4.578306,
  3.733363, 4.818157, 4.773763, 6.63829, 6.693108, 5.663667, 6.9752, 
    6.861635, 5.952466, 4.597996, 4.801058, 5.300307, 5.261598, 5.284022, 
    5.06571,
  6.08744, 6.563444, 6.861777, 7.862533, 5.887674, 5.116416, 7.163911, 
    7.008981, 6.771699, 5.679075, 4.752075, 5.388735, 5.263871, 4.190175, 
    4.704868,
  6.682047, 7.530148, 8.000917, 8.54917, 6.139652, 4.847384, 6.356835, 
    6.545888, 6.584699, 6.230224, 5.868853, 5.617915, 5.185561, 4.962646, 
    4.579366,
  6.727475, 7.677144, 8.464869, 8.757381, 8.636769, 6.419299, 4.825965, 
    4.793852, 5.972663, 6.573406, 6.139932, 5.564846, 5.178267, 4.966974, 
    3.858509,
  6.786624, 7.345289, 8.593844, 8.773232, 9.256378, 8.872663, 7.155409, 
    4.565448, 4.462164, 4.955766, 5.86217, 5.431387, 5.068362, 5.011137, 
    3.837514,
  6.502294, 7.126547, 7.825589, 8.268197, 9.097902, 9.414172, 9.657617, 
    8.592108, 5.475013, 4.502418, 3.98997, 4.8932, 4.903728, 4.93289, 4.103454,
  6.150062, 6.50293, 6.896884, 7.690698, 8.936546, 8.892022, 9.205179, 
    6.764947, 7.341681, 6.154454, 5.140564, 4.553709, 4.565471, 4.774426, 
    4.313322,
  5.553789, 5.940236, 6.619542, 8.137755, 8.524985, 8.346354, 7.32806, 
    6.48807, 7.43379, 5.543706, 4.356491, 3.935123, 4.090319, 4.676242, 
    4.239934,
  4.696618, 5.410566, 6.786629, 8.151649, 7.950442, 7.73058, 6.89434, 
    6.718284, 5.805406, 3.824841, 2.630821, 3.139716, 3.676525, 4.214162, 
    4.149008,
  4.38447, 5.455795, 7.541557, 8.526927, 8.115942, 6.992361, 6.652779, 
    6.77158, 4.11432, 2.157371, 2.122083, 3.533182, 3.633554, 3.708782, 
    3.747138,
  5.030089, 7.635671, 7.774604, 10.16202, 10.01009, 8.572594, 10.86845, 
    10.97728, 9.396014, 7.053697, 7.363592, 7.344725, 5.811811, 3.813246, 
    2.795027,
  7.179128, 8.078465, 8.931463, 9.841882, 6.359516, 5.585195, 8.913718, 
    9.682654, 8.411827, 6.694199, 6.963369, 8.794448, 8.247634, 4.122684, 
    2.425483,
  6.769485, 7.245292, 8.044274, 7.966333, 5.40472, 4.11964, 6.780901, 
    8.304779, 8.118555, 7.917843, 7.982601, 8.424147, 9.420941, 6.100912, 
    2.553313,
  6.029788, 6.27525, 6.884396, 7.050125, 7.019897, 4.972373, 4.347962, 
    5.977822, 8.107106, 8.682367, 7.693871, 9.538383, 9.383108, 5.823813, 
    2.460596,
  5.614812, 5.643327, 6.310213, 6.823706, 7.658781, 7.600739, 5.617341, 
    4.456107, 5.672052, 5.423202, 8.131817, 10.04403, 8.530675, 5.766497, 
    3.405086,
  5.228539, 5.468494, 5.989915, 6.563969, 7.540301, 8.445187, 8.299379, 
    6.596585, 4.143837, 4.844713, 5.369114, 7.912459, 6.415279, 4.89425, 
    3.782947,
  4.640005, 5.395734, 6.09379, 6.556326, 7.050149, 7.668324, 7.590041, 
    7.990458, 7.497478, 6.609601, 6.041046, 5.059379, 4.339145, 4.120275, 
    3.628431,
  4.345908, 5.788942, 6.424648, 6.901217, 7.124533, 7.08396, 7.113769, 
    7.010029, 6.098073, 5.056329, 3.863583, 2.301799, 2.396056, 3.376446, 
    3.723785,
  5.022658, 6.325091, 6.892479, 7.312233, 7.097653, 6.876248, 6.789196, 
    6.274011, 5.341651, 4.298645, 2.88321, 1.495157, 1.229415, 2.423969, 
    3.933072,
  5.708282, 6.846152, 7.434091, 7.155832, 6.825329, 6.731318, 6.509235, 
    5.873706, 4.755548, 3.118381, 2.399424, 2.0544, 1.678319, 2.092455, 
    3.303101,
  5.130231, 7.97189, 7.380106, 8.137959, 7.02, 7.058786, 9.851826, 10.30065, 
    9.893672, 7.351881, 5.913312, 5.738534, 5.653381, 6.334366, 6.491904,
  6.671037, 8.119482, 9.211805, 8.937675, 5.343812, 5.437273, 9.05003, 
    10.38978, 11.4205, 11.14455, 8.47059, 5.321965, 5.931521, 5.792884, 
    5.864251,
  6.04506, 7.510176, 9.145753, 9.350968, 6.437632, 4.493182, 6.71223, 
    8.250513, 10.11246, 12.84807, 12.35769, 6.914056, 3.972776, 8.457891, 
    7.19174,
  5.623781, 6.838472, 8.212439, 9.230722, 9.02387, 5.906301, 4.191795, 
    6.835984, 11.44586, 13.91238, 13.76886, 10.74642, 7.299641, 8.897576, 
    7.395188,
  5.577715, 6.394, 7.376988, 8.084586, 8.928741, 9.048074, 6.503115, 
    4.732984, 6.546689, 8.491673, 12.19593, 12.8794, 10.93448, 9.594442, 
    8.342923,
  5.586995, 6.118831, 6.90625, 7.619422, 8.20715, 8.478246, 8.57516, 
    7.349016, 4.870141, 4.953914, 6.590765, 10.25544, 10.54532, 10.02623, 
    9.189168,
  5.528462, 6.231934, 6.597878, 7.208973, 7.519813, 8.00359, 7.949673, 
    7.77517, 7.150998, 6.61497, 6.678656, 7.538726, 8.028619, 7.974745, 
    7.636354,
  5.695416, 6.45804, 6.630692, 7.017244, 7.170176, 7.829386, 7.878131, 
    7.148263, 6.340178, 5.477149, 5.013443, 4.689868, 4.811741, 4.91616, 
    5.443671,
  5.851654, 6.319296, 6.284603, 6.393928, 6.793781, 7.454206, 8.002739, 
    7.619155, 6.492896, 5.395409, 4.258661, 3.262049, 2.886217, 2.824627, 
    3.217334,
  5.671166, 5.976677, 6.202265, 6.33356, 6.718823, 7.415916, 8.103863, 
    7.523731, 5.616453, 3.505224, 2.718977, 1.938182, 1.407222, 1.79409, 
    2.236202,
  4.5341, 7.208234, 7.183094, 9.025417, 7.364671, 4.923476, 6.31092, 
    6.987154, 6.652081, 6.365095, 7.472379, 8.156704, 6.66619, 5.30304, 
    4.857944,
  7.90764, 8.444409, 8.224494, 8.366421, 5.391117, 4.624192, 6.623808, 
    7.545889, 7.631449, 7.965908, 8.704692, 9.50306, 8.325081, 5.775013, 
    5.772517,
  8.891034, 9.696839, 9.377176, 7.691337, 5.036367, 4.440203, 6.653004, 
    6.970291, 6.771475, 9.429745, 11.91769, 11.23562, 6.940794, 7.423498, 
    7.194506,
  9.034582, 9.953355, 9.726498, 8.296339, 6.434102, 4.459606, 4.641893, 
    6.052167, 8.274145, 10.52204, 12.74341, 13.47892, 7.947633, 5.122508, 
    7.576662,
  8.988174, 9.687409, 9.697818, 8.563704, 7.294005, 6.249416, 4.8921, 
    3.661159, 5.160456, 7.287263, 10.91483, 13.2899, 12.27116, 6.947807, 
    8.018232,
  8.920984, 9.702572, 9.612028, 8.897494, 7.537151, 6.957684, 6.224391, 
    4.617913, 3.615482, 4.623783, 6.536967, 10.62537, 12.41144, 11.61342, 
    8.599333,
  8.690052, 9.501457, 9.50941, 8.773963, 7.3983, 7.115569, 6.560286, 
    5.827798, 5.552845, 6.787846, 8.301649, 9.181737, 9.785406, 9.806163, 
    8.714789,
  8.508806, 9.449655, 9.370408, 8.584322, 7.44838, 7.079735, 6.463001, 
    5.379172, 4.887107, 6.227301, 7.327082, 8.350623, 8.851926, 8.620948, 
    7.414143,
  7.995178, 8.794388, 8.418941, 7.709094, 7.104321, 6.913029, 6.84712, 
    6.326967, 5.588855, 6.072583, 6.998302, 7.681789, 8.399003, 9.029461, 
    8.241613,
  7.199745, 7.747315, 7.449536, 7.515871, 7.561385, 7.526321, 6.877102, 
    6.530638, 5.282618, 4.018661, 4.443635, 6.715124, 7.926753, 9.002356, 
    9.516198,
  3.730302, 4.757496, 4.283849, 6.54504, 5.674945, 4.359392, 5.461015, 
    5.621859, 4.954644, 4.515191, 5.289076, 5.68545, 6.020315, 6.175553, 
    4.479539,
  5.512421, 4.653363, 4.671892, 5.845747, 4.497976, 4.227147, 6.070745, 
    6.685225, 6.490904, 5.757453, 5.376036, 6.751932, 6.377026, 4.509506, 
    3.988867,
  6.354535, 4.867756, 4.957156, 5.250803, 4.400102, 3.824648, 5.705739, 
    6.244249, 5.780544, 6.374912, 6.847538, 7.216319, 6.259607, 5.17572, 
    4.111101,
  6.371094, 4.969573, 4.821468, 5.219038, 5.473013, 4.045871, 3.852405, 
    6.071121, 8.869392, 9.078269, 8.339254, 7.738572, 6.632608, 4.128643, 
    4.760738,
  6.001711, 4.762549, 4.462961, 4.734615, 5.367531, 6.015384, 4.499115, 
    3.941221, 5.854828, 7.241122, 9.204986, 8.4298, 7.072002, 4.204996, 
    4.176437,
  5.518331, 4.827742, 4.385458, 4.736217, 5.378916, 6.267951, 6.260535, 
    5.754508, 5.353556, 6.244409, 6.979955, 8.99021, 7.252298, 6.168036, 
    3.35749,
  5.123486, 4.898668, 4.323793, 4.507054, 5.123462, 6.104509, 6.70234, 
    7.84323, 8.693141, 10.03622, 11.70744, 11.05829, 7.343699, 6.263604, 
    5.300653,
  5.039083, 4.905472, 4.07759, 4.181283, 4.977445, 6.048189, 6.718656, 
    7.778111, 9.077327, 10.59054, 12.74727, 13.3128, 9.608854, 6.420431, 
    6.477169,
  5.283459, 4.812665, 3.812891, 3.586328, 4.436064, 5.83083, 6.958193, 
    8.574875, 9.92205, 11.28725, 13.38912, 14.8712, 13.44241, 7.139483, 
    6.712635,
  5.649896, 4.695731, 3.456741, 3.153157, 4.240089, 5.701818, 6.992538, 
    8.349966, 8.466695, 7.468859, 9.785301, 14.87202, 15.55883, 12.39998, 
    5.989007,
  5.667792, 9.861054, 5.697868, 3.104542, 2.36109, 3.979468, 6.8244, 
    7.898607, 6.477004, 4.958436, 5.332841, 6.280069, 7.224287, 8.088655, 
    5.932729,
  11.67533, 11.32482, 6.350156, 2.995663, 2.749736, 4.372473, 7.461507, 
    8.766291, 8.179262, 5.785412, 5.17468, 6.527222, 6.717733, 6.270746, 
    6.587019,
  12.53416, 9.883056, 6.434718, 4.091528, 3.587837, 4.055944, 7.573145, 
    8.454372, 7.46233, 6.894836, 6.042554, 5.821153, 5.268262, 6.696894, 
    7.308098,
  10.39168, 7.902397, 5.667711, 4.709157, 5.290252, 4.405002, 5.536764, 
    8.09978, 10.55021, 10.16939, 7.481745, 5.154327, 3.715286, 4.030991, 
    6.641348,
  7.962404, 6.172441, 4.731473, 4.511693, 5.531099, 7.28868, 6.503393, 
    5.396419, 7.16376, 8.446284, 8.985214, 5.200574, 2.89623, 1.86402, 
    5.601025,
  6.151836, 5.152081, 4.385026, 4.685975, 5.993515, 7.656744, 8.803703, 
    8.043556, 6.84602, 7.557886, 6.678556, 5.256769, 2.852347, 3.171849, 
    3.686076,
  5.032794, 4.477167, 4.126705, 4.454681, 5.866613, 7.782741, 9.328668, 
    10.36868, 11.55599, 13.01055, 12.29922, 7.372914, 2.61134, 3.820991, 
    3.589998,
  4.622408, 4.125598, 3.684206, 4.035153, 5.723168, 7.959082, 9.299107, 
    9.952121, 11.34257, 13.21475, 13.5335, 10.11238, 4.013336, 3.812772, 
    3.810479,
  4.447771, 4.030855, 3.008189, 2.989768, 4.814374, 6.957612, 8.948109, 
    10.54067, 11.63918, 12.80642, 13.56216, 12.00141, 6.369207, 2.167198, 
    3.937557,
  4.531761, 3.798745, 2.137663, 2.17039, 3.916909, 5.965846, 8.164853, 
    9.566855, 9.235287, 7.738825, 9.378585, 12.53969, 9.800224, 3.036503, 
    3.279793,
  6.25659, 8.118848, 4.933078, 4.458513, 3.524905, 3.371009, 4.695673, 
    5.515089, 5.627332, 5.105206, 5.537499, 5.675204, 5.384732, 5.535329, 
    6.525201,
  8.9073, 7.533527, 5.791392, 4.925858, 3.780656, 3.760345, 5.394253, 
    6.444239, 7.2481, 5.844193, 5.091877, 5.253482, 4.545837, 3.870698, 
    6.395146,
  7.439638, 6.691087, 6.541468, 6.106449, 4.752018, 3.848323, 6.076629, 
    6.536151, 6.589988, 6.811646, 5.611067, 4.201701, 3.350573, 5.155102, 
    7.427216,
  5.473611, 5.666299, 6.128872, 6.549283, 6.662408, 4.916386, 4.353755, 
    6.406621, 9.172581, 9.305777, 7.055681, 4.628247, 3.990281, 6.183089, 
    7.431144,
  3.967417, 4.657702, 5.67417, 6.537142, 7.159868, 7.44057, 5.472585, 
    4.419492, 6.042244, 7.061566, 7.179514, 5.467759, 4.592757, 6.835124, 
    8.971112,
  2.714394, 3.382589, 4.817349, 6.395445, 7.05924, 7.464474, 7.460787, 
    6.542287, 5.724651, 6.143534, 5.130737, 5.606728, 5.49366, 6.967605, 
    8.911205,
  2.174047, 2.012469, 3.381052, 5.323845, 6.572313, 7.234046, 7.831201, 
    8.232909, 9.292439, 10.16656, 9.026736, 6.331042, 5.422461, 6.734677, 
    8.324047,
  2.434264, 1.52505, 1.735249, 3.649235, 5.648885, 6.837098, 7.522994, 
    7.448736, 8.687477, 10.36223, 10.16249, 7.826664, 5.495412, 6.44179, 
    7.878479,
  3.117228, 2.342123, 1.3238, 1.975197, 3.811753, 5.451927, 7.019375, 
    8.167681, 9.331037, 10.41964, 10.70622, 9.475924, 6.775011, 5.855091, 
    7.072472,
  4.174861, 3.473053, 2.395637, 1.808032, 2.39321, 3.733289, 5.80163, 
    7.382049, 7.61621, 6.626839, 7.347349, 10.03318, 8.213078, 5.677425, 
    5.73209,
  2.125355, 3.230781, 3.920905, 5.232425, 4.216912, 3.0979, 3.911947, 
    4.335047, 4.473898, 4.09817, 4.49556, 4.143344, 3.48183, 3.491853, 
    4.173389,
  2.335519, 2.452754, 4.403342, 5.753551, 3.955862, 3.45841, 4.878748, 
    5.377684, 5.758962, 5.669002, 5.217556, 4.886556, 4.190024, 3.172047, 
    3.635123,
  2.356157, 2.99439, 4.473212, 5.684221, 4.348107, 3.38418, 5.133716, 
    5.227089, 5.205696, 6.563324, 7.117524, 5.765512, 4.698816, 4.968129, 
    5.169871,
  2.311784, 2.447637, 3.878616, 4.957731, 5.363504, 3.886806, 3.659201, 
    4.990788, 7.124381, 8.476176, 8.643362, 7.148588, 5.623805, 5.472908, 
    5.662197,
  2.863462, 1.760832, 3.167349, 4.447094, 5.187026, 5.62389, 4.497539, 
    3.623218, 4.965151, 6.758267, 8.81552, 8.037886, 6.502162, 6.221369, 
    6.695365,
  4.000605, 1.6463, 2.338907, 3.9185, 4.7776, 5.516834, 5.857795, 5.269103, 
    4.904205, 5.527175, 6.218498, 8.096229, 7.38201, 6.978347, 6.62879,
  5.073925, 2.08899, 1.34218, 2.781772, 4.262426, 5.386111, 6.206185, 
    6.637655, 7.279332, 8.699484, 9.734892, 9.334773, 8.16348, 7.712053, 
    5.363132,
  5.895756, 2.894951, 1.439346, 1.639037, 3.82917, 5.263067, 6.245866, 
    6.497888, 7.114894, 8.901579, 10.34737, 10.32066, 9.206928, 8.409966, 
    5.216876,
  6.10259, 3.702544, 3.23012, 1.769029, 2.284001, 4.704071, 6.318354, 
    7.232965, 8.04355, 9.377636, 10.80651, 11.22301, 10.04259, 8.60707, 
    6.182712,
  5.716303, 3.224146, 3.627928, 2.126851, 1.583851, 3.693083, 5.596639, 
    7.133415, 7.203068, 6.342897, 8.138962, 11.47777, 10.6041, 8.655468, 
    6.758204,
  2.32044, 2.451323, 3.148127, 4.333826, 3.655387, 3.040212, 4.079263, 
    4.615154, 4.572065, 4.217107, 5.243555, 6.120952, 5.166992, 3.5121, 
    2.571395,
  3.151183, 1.901879, 3.472002, 4.537079, 3.402725, 3.193837, 4.612344, 
    5.216824, 5.028565, 5.130198, 5.881779, 7.469724, 6.693174, 3.503727, 
    2.907155,
  3.675436, 1.780593, 3.28487, 4.465673, 3.66827, 3.10533, 4.628488, 
    4.628105, 4.028625, 5.563977, 7.486359, 8.418316, 7.667295, 5.834404, 
    3.894398,
  5.085946, 2.241526, 3.227722, 4.174583, 4.66134, 3.694804, 3.50003, 
    4.455936, 5.764039, 7.007546, 8.354527, 9.375966, 8.687266, 6.486197, 
    4.385917,
  5.367703, 2.648633, 2.940411, 3.719416, 4.440848, 5.160017, 4.337641, 
    3.387756, 4.495162, 6.014611, 8.725371, 10.15076, 9.232433, 6.986163, 
    5.489381,
  5.09637, 2.789088, 2.731289, 3.493684, 4.304685, 5.178081, 5.406551, 
    4.95525, 4.549355, 5.261946, 6.561006, 10.25466, 9.183216, 7.057552, 
    5.443787,
  4.28381, 2.80754, 2.385401, 2.875907, 4.108588, 5.205338, 5.837595, 
    6.510145, 7.229435, 8.204713, 9.682145, 10.93926, 9.019213, 7.066102, 
    3.698006,
  3.731261, 2.893796, 2.262275, 2.622382, 4.171014, 5.24008, 5.90797, 
    6.461941, 7.29931, 8.623436, 10.4288, 11.42694, 8.773616, 6.140867, 
    2.673638,
  3.392414, 2.755495, 2.016932, 2.48623, 3.936367, 4.84507, 5.580381, 
    6.904922, 8.177739, 9.327064, 11.1384, 11.53825, 8.334092, 5.03837, 
    3.350187,
  3.09043, 3.409309, 3.313175, 3.564689, 4.057131, 4.115321, 4.480311, 
    6.029708, 6.787979, 6.073861, 8.429012, 10.88835, 7.793093, 4.670509, 
    3.621922,
  1.686502, 2.671853, 3.132903, 4.162825, 3.817627, 3.217187, 4.238862, 
    4.33733, 3.386983, 3.03137, 3.569714, 4.104347, 4.433851, 4.082917, 
    3.649033,
  1.996451, 3.301788, 4.103914, 4.582201, 3.509156, 3.253317, 4.618452, 
    4.633446, 4.223876, 3.96082, 4.044078, 4.991011, 5.639368, 3.676991, 
    3.676436,
  2.430599, 4.335355, 4.833547, 5.03932, 3.833424, 3.497406, 4.59195, 
    4.568292, 4.131503, 4.633475, 5.128411, 6.012105, 6.417562, 5.847018, 
    4.469928,
  3.586803, 5.496468, 6.12054, 6.037518, 5.85377, 4.809917, 4.039382, 
    4.257452, 4.434238, 4.756636, 5.749473, 6.815754, 7.071306, 6.517533, 
    4.832188,
  5.165553, 6.688153, 7.074007, 6.860399, 6.840921, 6.668228, 5.808839, 
    4.17771, 4.141627, 4.528879, 6.388993, 7.523285, 7.654592, 6.815706, 
    5.555126,
  6.512869, 7.781093, 7.483294, 7.00736, 7.112057, 7.374579, 7.552542, 
    7.697651, 6.332778, 5.289978, 5.228106, 7.863252, 7.933676, 6.608442, 
    5.728251,
  7.564444, 8.368467, 8.082239, 7.452971, 7.756711, 7.88951, 8.124894, 
    7.937937, 7.855288, 7.441941, 7.128023, 7.953763, 7.854709, 6.25037, 
    5.379701,
  8.185482, 8.998043, 8.527885, 8.118625, 8.431298, 8.199074, 7.406078, 
    5.947275, 5.047627, 5.693646, 6.563309, 7.862001, 7.692132, 6.17195, 
    4.977793,
  8.660125, 9.116856, 8.293658, 8.12087, 8.589615, 7.915985, 6.262572, 
    3.967452, 3.483189, 4.021519, 6.062839, 7.919308, 7.698816, 5.915386, 
    4.452616,
  8.956388, 8.707696, 8.301989, 8.477445, 8.521746, 7.135811, 4.800728, 
    3.029349, 2.760858, 3.604353, 5.941803, 8.776789, 7.16144, 5.590346, 
    4.369606,
  3.685625, 5.285949, 5.268285, 7.122995, 6.911534, 6.360572, 8.136237, 
    8.160883, 7.560526, 5.268076, 4.257013, 3.57776, 2.411347, 1.571649, 
    1.954484,
  5.569728, 6.97339, 7.682635, 8.502868, 6.249047, 6.38006, 9.557194, 
    9.477779, 9.007659, 7.517758, 5.788081, 5.465451, 4.197347, 1.793829, 
    1.23737,
  6.543299, 8.160968, 8.546268, 8.590949, 5.932563, 5.309897, 7.608562, 
    9.28642, 9.581846, 9.260018, 8.411839, 7.333502, 5.897762, 3.792913, 
    1.632691,
  7.495176, 7.905906, 7.766999, 7.285642, 6.596558, 4.726171, 4.300434, 
    5.447289, 6.958665, 8.800714, 10.04432, 9.011317, 7.168379, 5.153117, 
    2.72073,
  7.696424, 7.338217, 7.35524, 6.887368, 6.314342, 5.466665, 4.490171, 
    3.183173, 3.708358, 4.271169, 7.902797, 10.09885, 8.573471, 6.523205, 
    4.119341,
  7.323919, 7.182924, 7.511789, 7.486452, 7.170782, 6.87372, 6.400703, 
    6.625677, 5.530377, 3.687713, 4.366167, 9.199336, 9.459157, 7.168706, 
    5.008132,
  7.220008, 7.463075, 7.875081, 7.809114, 8.043963, 7.252795, 7.00747, 
    6.74099, 6.129685, 6.177238, 6.46285, 8.662836, 9.570481, 7.690621, 
    5.732122,
  7.581317, 7.802509, 8.038416, 8.383687, 8.983486, 8.033381, 6.173992, 
    5.225332, 3.771315, 4.054854, 6.553249, 8.654038, 9.764725, 8.320726, 
    6.362292,
  7.903901, 7.978513, 8.069279, 8.697926, 9.518082, 8.657922, 6.195903, 
    4.502319, 3.772699, 2.455355, 5.942789, 8.802641, 9.626422, 8.520728, 
    6.353417,
  8.046511, 8.179563, 8.413036, 9.828894, 11.23152, 10.32402, 7.35103, 
    3.710347, 5.140011, 3.669491, 4.991907, 9.299438, 9.560884, 8.4501, 
    6.527164,
  3.096293, 3.590151, 3.20848, 3.2931, 2.716099, 2.312509, 3.460509, 
    4.388363, 5.676505, 4.747056, 4.524399, 4.52176, 3.562664, 2.277769, 
    1.19646,
  4.879488, 4.912076, 5.276945, 5.246616, 3.377175, 2.941529, 3.727559, 
    3.902761, 5.661718, 6.600757, 5.565567, 5.851747, 5.481241, 2.870084, 
    1.184529,
  5.767039, 6.588507, 6.365032, 5.861879, 4.521881, 3.665358, 3.859909, 
    3.185731, 3.970684, 6.675342, 7.669799, 7.203724, 6.552987, 4.928332, 
    1.962119,
  6.844092, 7.309398, 6.975689, 5.261694, 4.955563, 4.602893, 3.209767, 
    2.580037, 2.578793, 4.051567, 7.2169, 8.050968, 7.610229, 5.930317, 
    2.746667,
  7.471982, 7.08797, 5.930838, 3.398798, 3.247629, 4.747588, 5.550014, 
    3.917758, 3.10026, 2.443743, 5.047457, 8.139416, 8.67029, 7.418575, 
    2.78936,
  7.696493, 6.711078, 4.421993, 3.218823, 3.889377, 4.905604, 6.116199, 
    7.890728, 5.814229, 3.229293, 3.1053, 7.705014, 9.637033, 7.887837, 
    3.423576,
  7.674646, 6.446871, 4.397213, 4.019292, 5.431439, 6.307226, 5.577468, 
    6.146436, 7.246934, 6.045132, 4.240312, 7.360747, 10.5637, 8.493814, 
    4.920674,
  7.735454, 6.749447, 5.128788, 5.423997, 6.871085, 6.547233, 4.802649, 
    4.55101, 7.487153, 7.751974, 5.181873, 7.706087, 11.52739, 9.044061, 
    5.910525,
  7.93223, 7.105894, 5.81003, 6.429674, 6.684157, 4.63504, 3.627173, 
    4.213782, 8.4547, 8.226187, 6.007089, 9.377515, 12.30903, 9.170903, 
    5.849138,
  7.884896, 7.527554, 6.61494, 7.021079, 6.534059, 4.568059, 3.853379, 
    6.724612, 8.493989, 5.420573, 5.815576, 11.309, 11.5772, 8.507961, 
    5.001537,
  4.159345, 6.325218, 5.957095, 7.427367, 6.433836, 4.455762, 3.95559, 
    1.892727, 1.578059, 2.837821, 3.648263, 4.268304, 3.978059, 3.201962, 
    2.710592,
  4.730346, 5.545348, 6.039441, 7.055407, 5.572299, 5.549993, 7.172269, 
    4.494085, 2.642428, 3.492016, 4.090087, 5.333202, 5.245983, 3.153945, 
    2.781082,
  4.229478, 4.55782, 4.73049, 5.067556, 4.449118, 4.468998, 6.631915, 
    7.221831, 4.773491, 4.245323, 5.10422, 5.959546, 5.533237, 4.374974, 
    3.470243,
  5.168655, 4.786511, 4.046414, 2.208763, 1.976752, 2.312826, 3.132133, 
    5.205232, 5.353807, 4.888149, 5.529302, 6.095989, 5.870831, 4.660262, 
    3.72726,
  5.668899, 4.279093, 2.807587, 0.9932436, 1.385936, 1.999543, 2.549249, 
    4.445842, 4.15548, 3.837293, 6.033859, 6.366197, 6.087077, 5.493418, 
    3.27793,
  5.828238, 4.028072, 1.778339, 1.964105, 2.331012, 1.218768, 1.845479, 
    5.475215, 5.434137, 4.963375, 5.308749, 7.054428, 6.712421, 5.293649, 
    2.924316,
  5.646012, 4.042382, 2.354627, 1.92731, 3.276054, 1.843713, 1.815829, 
    4.257364, 7.059637, 7.423542, 7.633446, 7.485266, 6.790578, 4.931045, 
    3.256842,
  5.701716, 4.69024, 3.373283, 1.955613, 2.623174, 2.99686, 3.340391, 
    6.462562, 7.77048, 7.906186, 7.778518, 7.685353, 6.451999, 4.632257, 
    3.135002,
  6.205777, 5.720439, 4.044811, 2.775805, 2.649217, 4.218502, 5.455263, 
    7.273319, 8.10288, 8.027838, 7.358194, 7.618468, 6.273396, 4.749903, 
    2.235447,
  6.157211, 6.260479, 5.096251, 4.581851, 4.672826, 5.423843, 6.929907, 
    8.564953, 7.646699, 5.79556, 5.740782, 7.837328, 5.664469, 3.430748, 
    1.640009,
  1.394028, 2.083516, 3.014941, 4.637712, 4.312543, 4.02556, 4.90425, 
    3.837334, 2.406496, 1.918372, 1.299302, 3.113515, 3.828556, 4.516675, 
    5.796059,
  2.608343, 3.842876, 4.401703, 4.575889, 2.827214, 3.162676, 5.147645, 
    4.694308, 2.830601, 2.467092, 1.963205, 3.403646, 4.546727, 3.911058, 
    4.851293,
  3.793535, 4.496412, 4.230668, 3.920918, 2.689933, 2.46387, 4.395526, 
    5.795762, 3.948998, 3.738288, 3.429211, 3.960479, 4.946692, 5.202467, 
    4.916282,
  5.081136, 5.251092, 4.787831, 3.519516, 2.434941, 1.945242, 2.669945, 
    4.166281, 3.952251, 4.304899, 4.634457, 4.347811, 4.648079, 5.082017, 
    5.259093,
  5.654206, 5.278713, 4.037992, 2.720253, 1.819125, 1.674675, 3.118108, 
    3.999199, 3.454686, 3.628148, 5.431635, 4.995209, 4.703285, 5.086613, 
    5.594097,
  5.918975, 4.600214, 2.873176, 1.662995, 3.456665, 2.840858, 1.858785, 
    3.768227, 5.173142, 5.301276, 5.046317, 5.912242, 5.216738, 5.333846, 
    5.630382,
  5.694351, 3.33107, 1.969775, 0.9521869, 3.878565, 3.796572, 1.722267, 
    2.236254, 7.20991, 8.370402, 7.965342, 6.767531, 5.880556, 5.489139, 
    6.127582,
  5.362928, 3.553457, 1.488382, 0.920377, 3.068726, 3.387201, 1.744073, 
    4.705158, 8.399533, 8.766111, 8.083426, 7.107541, 5.391289, 5.198467, 
    5.823062,
  5.801253, 4.994324, 3.111048, 2.920056, 3.867157, 2.804313, 3.014788, 
    6.847915, 9.228541, 8.696585, 8.173409, 6.911164, 5.181894, 5.137623, 
    4.971517,
  6.107138, 6.109696, 5.319133, 4.87165, 4.408502, 4.180257, 6.441334, 
    9.377023, 8.391569, 6.039836, 6.087082, 6.822254, 4.990656, 4.892703, 
    3.631882,
  1.307616, 1.548155, 1.726615, 2.506641, 2.750428, 3.06134, 4.525491, 
    4.85814, 4.541306, 3.441434, 2.57088, 3.212562, 4.333379, 5.54595, 
    6.226547,
  2.254493, 2.856043, 3.735721, 4.055254, 3.031619, 3.551241, 5.437887, 
    4.842277, 4.160699, 2.99284, 2.32666, 3.702293, 5.462535, 5.389098, 
    4.685044,
  2.546785, 3.880473, 4.429324, 4.663224, 3.526691, 3.023165, 3.794998, 
    3.314914, 3.091317, 2.417681, 2.165053, 4.768085, 6.676984, 6.819794, 
    3.704982,
  4.194179, 5.625927, 5.665509, 4.802332, 3.932188, 2.695571, 1.603502, 
    2.080487, 2.688578, 2.204077, 2.571255, 5.237847, 6.557226, 4.718843, 
    4.642734,
  5.732358, 5.635215, 4.572282, 2.48978, 2.403485, 2.523633, 2.525719, 
    2.269091, 2.114722, 1.974374, 3.23862, 5.15098, 4.424369, 4.185804, 
    6.344978,
  5.466173, 4.028532, 1.967994, 1.248399, 1.442161, 1.087922, 2.104369, 
    2.461188, 2.57864, 2.484668, 2.677894, 3.687773, 4.020281, 6.710579, 
    8.427588,
  4.584195, 2.688093, 1.462678, 1.449944, 1.688515, 1.800887, 1.564142, 
    3.800876, 5.021909, 4.333836, 3.923548, 5.108872, 7.895837, 9.602176, 
    10.12197,
  3.537305, 2.535074, 1.658272, 1.768196, 2.381169, 1.923571, 4.005203, 
    6.86781, 6.941155, 5.820214, 6.825029, 8.642351, 10.13863, 10.68263, 
    10.3035,
  3.753837, 3.125594, 2.765312, 3.312557, 3.456764, 3.754842, 6.328453, 
    8.469604, 7.986617, 7.015053, 8.237969, 9.145607, 9.49337, 9.352166, 
    8.398838,
  4.154312, 3.866297, 3.466787, 3.6934, 4.087505, 5.541384, 8.012986, 
    8.980663, 6.881265, 5.212565, 6.233058, 8.3337, 8.284302, 8.039257, 
    7.518186,
  4.139874, 5.313426, 4.647046, 5.20763, 4.424725, 3.470677, 4.597951, 
    5.213777, 5.387692, 3.952996, 3.502793, 3.844421, 3.514037, 3.084018, 
    2.847853,
  6.250857, 4.899128, 3.862625, 3.675088, 2.541308, 3.101267, 5.595132, 
    6.362526, 6.74505, 6.052496, 4.907429, 5.104503, 4.963714, 3.299234, 
    3.164437,
  4.375514, 2.987448, 2.565776, 3.415045, 2.730384, 2.975693, 3.958723, 
    4.960949, 5.418814, 5.012949, 4.875903, 4.908935, 5.017354, 4.881989, 
    4.373243,
  2.659741, 3.499525, 4.454097, 2.997904, 2.183897, 2.244921, 2.474054, 
    2.0145, 3.091057, 4.260273, 4.553153, 4.408583, 4.600162, 5.289343, 
    5.197583,
  3.797436, 4.562211, 3.476512, 1.174137, 1.385342, 3.43711, 3.420933, 
    1.96999, 2.308197, 2.448706, 3.996102, 4.795374, 5.308631, 5.70824, 
    5.640424,
  4.183165, 3.319977, 2.283719, 2.131538, 3.608833, 4.496775, 4.560292, 
    4.32713, 3.049601, 2.042998, 2.675695, 4.80942, 5.253915, 5.150731, 
    5.609466,
  3.348148, 2.370839, 3.007194, 3.647566, 4.464292, 4.219961, 3.186455, 
    2.936748, 3.772895, 4.75186, 4.508108, 4.164834, 4.74053, 5.560352, 
    5.945594,
  2.650772, 3.141231, 3.632376, 3.81172, 3.616614, 2.679405, 2.847957, 
    3.527498, 4.993868, 4.024334, 4.593348, 5.660214, 6.442445, 7.300256, 
    7.418613,
  3.170064, 3.639104, 3.641628, 4.085973, 3.809037, 4.253114, 4.380724, 
    3.900522, 3.277719, 5.63123, 6.939974, 8.103263, 8.69158, 8.426462, 
    7.355602,
  3.619398, 4.320367, 4.635872, 5.80089, 5.964645, 5.202258, 3.618671, 
    4.290895, 5.969665, 5.7955, 7.375075, 9.66654, 9.070355, 8.408607, 
    7.626259,
  6.951286, 8.211737, 5.704196, 6.329492, 5.453324, 3.819982, 4.398412, 
    4.489924, 4.57489, 3.641351, 3.130688, 2.485161, 1.836937, 2.073669, 
    2.240334,
  9.84689, 8.67444, 7.502655, 7.246634, 4.560812, 3.488399, 4.659251, 
    5.029404, 5.674293, 5.254243, 4.317807, 4.328439, 3.293462, 2.145339, 
    1.819131,
  9.877298, 8.865843, 8.163866, 6.943089, 4.383836, 3.100825, 3.368508, 
    3.812658, 4.38136, 4.855301, 4.534564, 4.514787, 4.672301, 3.883861, 
    2.632234,
  10.05776, 9.378069, 7.773365, 5.223779, 3.943919, 3.263061, 2.431302, 
    2.569374, 2.75157, 3.661907, 3.838027, 3.575348, 4.341745, 4.452459, 
    3.388782,
  9.698224, 7.777601, 5.952264, 4.167098, 3.706305, 4.387686, 4.350475, 
    2.595648, 2.623408, 2.43118, 2.96562, 2.897088, 3.640482, 4.52602, 
    4.002055,
  7.342583, 5.56784, 4.465336, 3.929983, 4.612629, 5.775061, 5.832896, 
    5.464408, 3.725378, 1.796152, 1.340501, 2.008973, 2.644294, 4.206679, 
    4.223235,
  5.667292, 4.395339, 4.042178, 4.391224, 5.91449, 6.098384, 5.03345, 
    4.182375, 3.619712, 2.323955, 1.472562, 1.915254, 2.900473, 3.84163, 
    4.180788,
  4.582212, 3.811191, 4.054387, 5.398933, 6.865443, 5.36956, 3.696454, 
    3.063359, 2.872461, 3.015983, 2.291061, 2.253057, 2.87734, 3.293851, 
    3.500862,
  3.35346, 4.195244, 4.747879, 6.680311, 5.686555, 3.580704, 3.776984, 
    3.205806, 3.043994, 3.399115, 3.197488, 2.755806, 2.793803, 3.274516, 
    3.523529,
  3.236859, 5.031218, 5.470143, 5.700101, 3.346754, 2.510483, 3.152459, 
    3.620443, 3.062619, 2.393375, 2.358036, 3.263083, 3.431242, 3.659453, 
    3.557984,
  7.514862, 9.824857, 7.352287, 9.732175, 9.116546, 7.762655, 9.671262, 
    10.36912, 9.989787, 7.091558, 6.575269, 6.608792, 5.796978, 4.293056, 
    3.233154,
  9.408909, 9.960472, 9.423143, 9.617181, 7.241876, 6.088988, 8.511043, 
    8.82201, 8.829655, 7.877429, 6.9923, 7.508587, 6.447099, 3.848763, 
    2.690461,
  9.175187, 9.317482, 9.373819, 9.850688, 7.549833, 5.641829, 5.189419, 
    7.031215, 8.741411, 9.350488, 8.587681, 7.171042, 5.451472, 4.253849, 
    3.031888,
  8.355904, 7.974255, 8.014946, 8.286335, 9.400252, 8.913497, 7.729734, 
    7.637066, 8.524625, 7.705036, 7.217003, 5.587894, 4.475292, 3.906973, 
    2.78859,
  6.810507, 8.006995, 10.30529, 12.19847, 11.84694, 11.31988, 9.359244, 
    6.516198, 5.072853, 4.43798, 5.056102, 4.756609, 4.254679, 3.985486, 
    3.300311,
  13.77484, 15.60547, 15.85187, 14.57053, 12.64516, 9.984213, 8.497131, 
    7.956007, 5.556458, 3.788006, 2.722496, 3.449403, 3.771075, 3.953672, 
    3.57748,
  14.49807, 14.79557, 13.58054, 11.87516, 10.31538, 9.050317, 8.005454, 
    7.198815, 6.200141, 4.624697, 2.533278, 2.155015, 3.55767, 4.362513, 
    3.957042,
  11.67555, 11.45954, 10.25152, 8.806629, 7.972268, 8.21123, 7.752204, 
    7.097328, 5.630671, 4.14741, 2.474146, 3.22913, 4.057134, 4.567956, 
    3.229941,
  8.337463, 8.072527, 7.082008, 6.586489, 6.905415, 6.989456, 6.636785, 
    5.810079, 4.629476, 3.674651, 3.048393, 3.632855, 3.80624, 3.399897, 
    1.6633,
  6.177373, 6.250618, 6.046633, 6.241143, 6.655776, 6.447309, 5.681068, 
    4.462315, 2.982006, 2.160694, 2.430608, 3.292431, 2.970126, 2.146874, 
    1.677321,
  5.72097, 10.89071, 11.26874, 15.27674, 14.31086, 10.81108, 12.19015, 
    12.22087, 11.18716, 7.934265, 7.88931, 8.050259, 7.173957, 6.369071, 
    6.263559,
  9.690592, 13.63069, 15.44635, 15.39377, 9.788487, 7.212472, 9.4973, 
    8.996441, 8.412619, 6.651915, 6.308527, 8.016592, 9.010255, 6.860663, 
    6.852462,
  11.72889, 13.79374, 13.78776, 12.32623, 7.385254, 4.321255, 3.328522, 
    4.447197, 4.643109, 3.702495, 3.36844, 4.757918, 7.612993, 9.871095, 
    8.799854,
  11.15307, 11.80562, 10.63273, 8.633683, 6.392814, 5.980621, 5.864886, 
    8.366776, 12.32363, 10.30205, 8.520135, 7.30755, 7.8245, 9.773837, 
    9.711141,
  9.015068, 9.373736, 9.390231, 11.17124, 12.72466, 11.65646, 8.813233, 
    6.165233, 6.672567, 7.352176, 9.855824, 10.70678, 11.54361, 12.09495, 
    11.35522,
  7.318593, 9.485225, 11.71869, 13.13711, 13.77845, 13.35336, 12.16605, 
    10.63297, 7.024369, 6.347711, 7.383781, 11.59708, 12.29952, 11.98062, 
    10.76521,
  6.090907, 8.251379, 10.12903, 11.19832, 11.50421, 11.21734, 10.77845, 
    10.19812, 9.026281, 8.671287, 8.947016, 9.888791, 10.3839, 10.1306, 
    8.845942,
  5.387882, 7.032693, 8.060462, 9.03459, 9.425648, 9.410253, 8.57325, 
    7.780239, 7.230688, 7.323253, 7.371324, 7.681136, 8.00717, 7.528951, 
    5.876077,
  5.08206, 5.622021, 5.860687, 6.653298, 7.107471, 7.415601, 7.293123, 
    6.954009, 6.455627, 6.122911, 6.412472, 6.67721, 6.553191, 5.346625, 
    3.731801,
  4.942921, 4.468466, 4.352119, 4.788554, 4.988835, 5.088184, 5.412005, 
    5.374502, 4.925735, 4.14259, 4.81939, 6.279142, 5.51935, 4.296762, 
    3.108459,
  5.968748, 7.305185, 6.826405, 8.830269, 7.691085, 4.883582, 5.743217, 
    6.006975, 6.24793, 5.933007, 7.219185, 8.473219, 8.254594, 6.990866, 
    6.003627,
  9.402742, 9.064221, 9.209753, 8.636412, 5.359462, 3.983577, 5.64474, 
    6.29171, 7.039519, 7.25579, 7.834287, 10.1854, 10.5866, 6.911164, 5.732992,
  10.70665, 9.669326, 9.110277, 8.385256, 5.296729, 3.568028, 4.613772, 
    5.229323, 6.62752, 9.007415, 10.79869, 11.32183, 11.12162, 9.845507, 
    6.596533,
  9.420182, 9.450794, 8.943141, 7.784721, 5.971469, 3.897571, 2.976371, 
    3.98045, 6.577118, 9.289709, 11.98551, 12.96907, 11.97711, 8.446168, 
    5.831782,
  11.11313, 9.57101, 8.309858, 6.461749, 4.895535, 4.266561, 3.764251, 
    3.107172, 4.681276, 6.915855, 12.05986, 14.01602, 13.39773, 6.518683, 
    5.243539,
  9.872309, 8.276926, 6.628011, 4.648084, 3.675263, 3.4346, 3.775557, 
    4.275279, 4.494422, 5.552221, 8.226834, 13.42265, 12.94719, 7.978747, 
    6.009706,
  7.097744, 6.102508, 4.480974, 2.928091, 2.659295, 2.921102, 3.707906, 
    4.83317, 5.625301, 7.096753, 9.685291, 11.7921, 10.49352, 9.065828, 
    9.562233,
  4.910827, 4.046904, 2.329307, 1.937584, 2.649029, 3.678136, 4.12321, 
    3.965254, 4.713819, 6.101606, 8.621233, 9.556819, 7.905096, 8.173949, 
    9.130311,
  3.836426, 2.339122, 1.195289, 2.049139, 3.142101, 3.985626, 4.299569, 
    3.845134, 3.968306, 5.002132, 7.044197, 7.642647, 6.123227, 6.386483, 
    7.497486,
  3.710315, 1.460558, 1.313709, 3.113223, 3.675033, 3.635947, 3.577955, 
    3.194839, 2.763613, 2.986612, 4.582068, 5.789166, 5.144267, 6.013829, 
    7.31798,
  9.729269, 13.91445, 12.36124, 15.94815, 13.65107, 9.850479, 11.41197, 
    11.41109, 10.06169, 7.158137, 6.590545, 6.146424, 5.447438, 5.097923, 
    5.27506,
  13.80319, 14.62388, 14.76513, 14.65693, 9.583276, 8.053489, 10.27617, 
    9.722125, 9.830834, 9.041741, 7.202137, 6.99773, 6.579993, 5.197864, 
    5.998962,
  13.14289, 13.64367, 13.33733, 12.95388, 10.20772, 8.623502, 9.552092, 
    11.65163, 11.70341, 9.241956, 7.184424, 6.70882, 7.372483, 9.027465, 
    8.68983,
  11.88571, 12.61122, 12.79486, 14.04561, 14.32402, 11.84466, 9.822556, 
    9.903992, 9.594731, 6.979484, 5.739778, 5.916625, 8.254464, 11.86062, 
    9.865947,
  10.77784, 12.59689, 13.95132, 14.88981, 14.28466, 12.59759, 9.097857, 
    5.987504, 4.590039, 3.60315, 4.351129, 6.276352, 10.08206, 12.2605, 
    7.300433,
  7.859733, 9.739417, 11.01322, 11.57216, 11.11636, 10.14733, 8.01201, 
    6.379817, 4.062398, 3.071515, 3.562857, 7.569849, 10.68195, 8.620585, 
    2.657441,
  5.296824, 6.470161, 7.50641, 7.613502, 7.53929, 7.075568, 5.723751, 
    4.913461, 3.842487, 3.500398, 5.598119, 7.849634, 8.121148, 5.760394, 
    3.970906,
  3.649451, 4.326989, 4.439634, 4.434964, 4.086006, 3.661545, 2.910617, 
    2.284777, 2.316835, 3.836531, 6.596104, 6.424726, 4.818917, 4.816568, 
    5.437138,
  3.214106, 3.241839, 3.014367, 2.848742, 2.256917, 1.6956, 1.901392, 
    1.580946, 2.277437, 4.459561, 6.206844, 4.503366, 3.59966, 4.779689, 
    5.755674,
  3.674176, 3.337338, 4.051155, 4.282445, 2.497905, 0.8963051, 0.9493821, 
    1.247668, 1.602904, 3.057186, 3.586511, 4.014008, 4.618836, 5.860037, 
    6.37162,
  4.566665, 5.73957, 4.776226, 9.004472, 10.62949, 9.920549, 13.0732, 
    13.46873, 11.38326, 7.308867, 5.808895, 8.269007, 10.13635, 9.050732, 
    7.210649,
  5.181449, 4.960437, 5.793924, 8.138896, 7.324691, 8.116054, 12.03615, 
    13.628, 12.8276, 10.70754, 9.945755, 12.19077, 11.72508, 7.203209, 
    5.532135,
  3.687866, 4.302346, 6.281939, 6.758329, 5.990911, 6.174798, 9.586873, 
    12.36067, 13.75897, 14.12669, 12.97893, 11.62341, 9.81438, 7.241813, 
    4.75776,
  3.57527, 4.261025, 6.032994, 5.734393, 6.822223, 5.847518, 5.281719, 
    8.708241, 13.06174, 12.35113, 10.52275, 8.411185, 6.099341, 4.020996, 
    3.45955,
  2.830256, 4.576725, 5.392044, 4.590339, 5.54865, 7.155675, 6.09657, 
    4.756941, 6.205981, 6.726479, 7.294, 5.880918, 3.95004, 2.963044, 3.145937,
  2.647658, 4.473223, 5.388419, 4.654811, 4.684464, 5.487415, 6.417318, 
    6.33904, 5.023706, 5.082079, 4.446656, 5.104445, 4.643462, 4.18486, 
    3.20596,
  2.702453, 4.005078, 5.803762, 5.976366, 5.01317, 4.09611, 4.562609, 
    5.834845, 7.110698, 7.252642, 6.13462, 5.00996, 4.513259, 4.019812, 
    4.551898,
  4.373045, 4.598917, 4.959938, 5.913389, 5.528434, 3.620597, 3.339463, 
    4.213918, 5.734076, 6.256017, 5.872817, 4.907413, 4.321795, 4.137877, 
    4.301745,
  5.0772, 4.412389, 4.051963, 5.335083, 5.539722, 3.9024, 2.606283, 2.986233, 
    4.918272, 5.525475, 5.072638, 4.719071, 4.449382, 4.470676, 4.361481,
  5.004166, 4.227044, 4.08257, 4.879226, 5.53793, 4.053899, 1.745789, 
    2.248958, 3.613988, 3.1782, 3.100884, 4.132089, 4.264055, 4.537349, 
    4.861667,
  2.578507, 3.231148, 2.561214, 4.925063, 5.086739, 2.323211, 4.025913, 
    6.487714, 8.278476, 7.449491, 7.180476, 7.46607, 7.135643, 6.302011, 
    5.44591,
  3.127608, 2.576297, 3.763133, 6.755276, 3.463165, 1.953717, 3.570992, 
    6.327447, 8.233388, 8.446393, 7.191055, 7.810575, 7.725171, 5.5847, 
    4.703831,
  3.768252, 3.876154, 6.302528, 6.109921, 2.517555, 1.693289, 3.756073, 
    5.298323, 6.92299, 8.837653, 8.930089, 7.944199, 7.548165, 7.383819, 
    5.481002,
  4.416405, 3.767884, 6.1043, 5.30712, 2.075357, 1.518629, 2.746898, 4.86742, 
    7.584758, 9.453128, 9.537274, 8.304862, 7.212005, 7.082396, 6.231048,
  4.486826, 3.137636, 4.852022, 4.799227, 3.033293, 1.559057, 2.593517, 
    2.990312, 4.765488, 6.403527, 8.613939, 7.902403, 6.944304, 6.742039, 
    6.546172,
  4.131157, 2.591176, 3.456842, 4.986271, 5.963345, 4.942424, 3.449689, 
    3.960803, 4.743459, 5.43875, 5.696213, 7.005308, 6.51423, 6.393756, 
    6.113472,
  3.390166, 3.603733, 3.839919, 4.936548, 6.081288, 6.192308, 4.423817, 
    3.517274, 6.008022, 7.42472, 7.760346, 7.058645, 6.262535, 6.419023, 
    5.870562,
  4.221092, 4.023413, 3.796343, 4.203461, 4.328714, 4.227703, 3.398725, 
    2.213709, 5.199077, 6.716758, 7.182174, 6.875724, 6.414193, 6.501583, 
    6.018156,
  4.524578, 4.364417, 3.964788, 3.79196, 2.668521, 4.240485, 4.480431, 
    2.290784, 4.747807, 6.01435, 6.493346, 6.50914, 6.365624, 6.673023, 
    6.215126,
  3.918012, 4.401687, 5.248535, 4.708655, 2.918736, 4.881489, 4.38554, 
    2.81492, 4.046171, 3.8797, 4.54807, 5.795297, 6.073484, 6.587388, 6.432084,
  6.084434, 8.068972, 7.148673, 9.391942, 7.63821, 4.500289, 3.958337, 
    3.901067, 4.587611, 5.030398, 6.142195, 6.770978, 5.903592, 4.924731, 
    4.509196,
  8.897402, 9.185845, 8.788509, 7.688766, 4.508142, 3.044667, 3.935743, 
    4.755202, 5.461016, 6.721138, 7.178289, 8.049959, 6.893485, 4.252796, 
    4.222587,
  9.776675, 9.475314, 8.15909, 5.832149, 3.321048, 2.3534, 3.575788, 
    4.193601, 4.412805, 7.137453, 9.176482, 8.838119, 7.165286, 5.842621, 
    4.733214,
  10.20061, 8.993945, 7.06308, 5.003005, 3.287555, 2.532403, 2.743251, 
    4.096309, 6.094682, 8.389143, 9.720734, 9.169725, 7.474607, 5.959756, 
    4.74121,
  9.630903, 7.618942, 5.382354, 3.422093, 2.354905, 3.138715, 3.713633, 
    3.413299, 4.675117, 6.331336, 9.042299, 8.821304, 7.585643, 6.355388, 
    5.603274,
  8.655436, 6.713774, 5.138793, 3.822802, 3.212048, 3.653519, 4.258744, 
    4.908537, 4.583368, 5.405103, 5.854782, 7.807315, 7.466548, 6.513604, 
    5.973603,
  8.139923, 7.02319, 6.195512, 5.8312, 5.426626, 5.067983, 5.010443, 
    5.900962, 6.118107, 7.22398, 7.674193, 7.48475, 7.054881, 6.797509, 
    6.750087,
  7.877615, 6.70252, 5.81726, 5.806335, 6.25481, 6.54376, 6.484674, 6.28363, 
    6.482932, 6.614762, 7.081485, 7.113154, 6.778552, 7.166646, 7.507485,
  7.425463, 6.194591, 5.142911, 5.270324, 6.013222, 6.565032, 6.526864, 
    6.728936, 6.841133, 6.61425, 6.861776, 6.88857, 6.504981, 7.3982, 7.377754,
  6.940652, 5.653308, 4.70545, 4.932364, 5.783169, 6.461397, 6.947235, 
    6.901775, 5.91229, 4.4483, 5.134927, 6.628623, 6.37788, 7.082258, 7.506353,
  7.443436, 8.830438, 5.396954, 4.750201, 3.270135, 2.818722, 3.909804, 
    4.881592, 5.520867, 5.115001, 5.798831, 6.164289, 5.122076, 3.939429, 
    3.399234,
  9.663918, 8.03284, 5.744534, 4.088457, 2.95023, 3.086249, 4.765794, 
    6.275388, 6.886387, 6.683034, 6.503424, 7.234287, 6.170165, 3.923161, 
    3.877316,
  8.937181, 6.808421, 5.370986, 4.837787, 3.702304, 3.262977, 5.176557, 
    5.564097, 5.552172, 6.78358, 8.149739, 7.822779, 6.793291, 6.016077, 
    5.126537,
  8.163181, 5.841264, 4.579003, 4.999186, 5.202277, 4.297071, 4.106473, 
    5.341384, 6.452888, 7.322016, 8.555694, 8.318347, 7.280718, 6.941268, 
    5.870325,
  7.479594, 4.904557, 3.850221, 4.556492, 5.276158, 6.032076, 5.238713, 
    3.868681, 4.857858, 6.067864, 8.293118, 8.437496, 7.780133, 7.704091, 
    7.375225,
  6.823903, 4.489832, 3.903683, 4.835734, 5.756822, 6.461123, 6.268765, 
    5.607107, 5.317203, 5.453798, 5.896907, 8.065314, 8.13402, 8.008396, 
    7.517764,
  6.649617, 4.540398, 3.912299, 4.838732, 6.160708, 6.957278, 7.027182, 
    7.011385, 7.186962, 7.482113, 8.161801, 8.538381, 8.160316, 7.997959, 
    7.327442,
  6.393133, 4.094501, 3.748367, 5.254678, 6.565691, 7.298712, 7.04408, 
    6.821303, 7.046202, 7.482174, 8.351067, 8.612493, 8.2096, 8.078849, 
    7.500876,
  5.885612, 3.516909, 3.436052, 5.16285, 6.680999, 7.516103, 7.304945, 
    7.294888, 7.433271, 7.648993, 8.230218, 8.667066, 8.335119, 8.150845, 
    7.238098,
  5.108588, 3.051543, 3.693625, 5.343654, 7.063961, 7.827036, 7.559279, 
    7.18174, 6.177115, 5.010316, 5.803638, 8.050215, 8.089046, 8.082212, 
    7.257362,
  4.652858, 5.687837, 3.892633, 4.096245, 3.675138, 3.24162, 4.678705, 
    5.744971, 5.276903, 4.323086, 4.893898, 5.643377, 5.921574, 5.314015, 
    4.437138,
  6.011617, 5.013546, 4.544637, 4.702092, 3.766623, 3.673494, 5.227595, 
    6.01695, 5.768956, 5.090009, 5.547692, 7.361078, 7.274546, 4.791304, 
    4.430137,
  5.446683, 4.104946, 4.402699, 5.234233, 4.175748, 3.863304, 5.813213, 
    5.324454, 4.412287, 5.4448, 7.457614, 8.258209, 7.389779, 6.097433, 
    4.668443,
  4.457997, 3.34329, 4.170568, 5.36531, 5.64071, 4.757866, 4.328369, 
    4.986431, 5.348096, 6.41604, 8.25492, 8.641547, 7.259491, 5.765297, 
    3.846611,
  3.530918, 2.958135, 4.400486, 5.608913, 6.418237, 6.280226, 5.076686, 
    3.546366, 4.447924, 5.863933, 8.596588, 8.541612, 6.638381, 5.41921, 
    4.349879,
  2.787829, 2.984489, 4.745108, 5.926569, 6.918806, 7.172493, 6.188945, 
    5.642689, 5.606257, 5.836391, 6.104379, 7.430709, 6.224082, 5.600541, 
    4.826008,
  2.327468, 3.119877, 4.951993, 6.005224, 7.194591, 7.651114, 7.514721, 
    7.446488, 7.367102, 7.451462, 7.540776, 6.785213, 5.937396, 6.010017, 
    5.424652,
  2.182599, 3.577334, 5.192337, 6.309313, 7.555552, 8.149636, 8.00158, 
    7.446622, 7.209827, 7.236029, 6.870722, 6.257405, 6.022545, 6.182257, 
    5.924354,
  2.468798, 4.096445, 5.090364, 6.066605, 7.470377, 8.350773, 8.612132, 
    8.162002, 7.480428, 6.857183, 6.294489, 5.977381, 5.75667, 6.037643, 
    5.84421,
  3.022678, 4.767258, 5.239201, 6.251131, 7.942361, 9.236679, 9.010199, 
    8.126148, 6.243183, 4.582788, 4.488494, 5.363643, 4.94983, 5.093126, 
    5.081191,
  3.510148, 3.568302, 2.806002, 4.886309, 5.043803, 4.324579, 5.466763, 
    6.211999, 5.265723, 3.81323, 3.734246, 3.765343, 3.623667, 3.105183, 
    2.425612,
  3.904027, 2.215195, 3.969098, 5.617564, 4.754234, 4.642085, 6.253866, 
    6.969957, 6.709616, 5.323512, 4.465867, 5.032444, 4.597116, 2.766902, 
    2.213319,
  2.657267, 2.096815, 4.741139, 6.218047, 4.965067, 4.791895, 7.098656, 
    6.999095, 6.56335, 6.15366, 5.988784, 6.003641, 5.31697, 4.338974, 
    2.918247,
  1.773443, 3.034988, 5.810017, 7.084332, 6.979499, 5.810116, 5.895841, 
    6.718745, 6.409164, 5.609342, 6.29279, 6.615903, 5.940412, 5.032027, 
    3.600158,
  1.667097, 4.263512, 6.921751, 7.377625, 7.999217, 8.027457, 6.860871, 
    5.492474, 5.540708, 5.209855, 6.528203, 7.233687, 6.519502, 5.743093, 
    4.945245,
  2.289981, 5.625086, 7.433821, 7.515643, 8.547606, 9.227502, 8.853489, 
    8.215578, 7.09355, 5.932242, 5.237381, 7.287799, 6.775018, 6.200098, 
    5.735801,
  3.296724, 6.371831, 7.230726, 7.425498, 8.513923, 9.400626, 9.962536, 
    9.552691, 8.247339, 7.005391, 6.31759, 6.48488, 6.379492, 6.306053, 
    6.155266,
  4.285204, 6.680775, 6.899928, 7.274683, 8.444448, 9.577949, 9.683411, 
    8.892779, 7.758016, 6.5441, 5.460681, 4.642043, 5.152205, 5.817284, 
    5.711402,
  5.298802, 6.598237, 5.905826, 6.692853, 8.098804, 9.300637, 9.475121, 
    9.125298, 7.778394, 6.037069, 4.555848, 3.276026, 3.289892, 4.267163, 
    4.80992,
  5.998925, 6.348254, 5.722981, 6.502735, 8.331654, 9.399215, 9.178941, 
    8.398985, 6.491601, 4.378747, 3.75394, 3.484225, 2.570668, 3.409486, 
    4.56056,
  3.961302, 3.938841, 1.829641, 4.699436, 5.891311, 5.200517, 6.694751, 
    7.049599, 6.163695, 4.568396, 4.229771, 4.079998, 3.293356, 2.255652, 
    1.060518,
  4.229977, 1.618651, 3.739586, 5.982693, 4.848755, 4.617608, 6.582582, 
    7.193106, 6.483713, 5.011147, 4.416325, 5.23716, 5.153856, 2.976444, 
    1.465423,
  2.775343, 2.231209, 5.220922, 5.918705, 4.368438, 4.428874, 6.048573, 
    6.471203, 5.894968, 4.564513, 4.280564, 5.206669, 6.387516, 5.509103, 
    2.988375,
  1.580218, 3.912913, 5.778943, 5.992256, 5.935798, 4.810228, 4.883358, 
    5.141255, 4.69748, 3.433193, 3.453153, 4.411375, 6.200716, 6.391632, 
    4.521099,
  1.811112, 4.622564, 5.565541, 5.945582, 7.150774, 6.784921, 5.486651, 
    4.167355, 3.729585, 2.996564, 3.397436, 4.070026, 6.063494, 7.200484, 
    6.282054,
  2.713555, 4.369704, 5.260134, 6.656686, 8.15206, 8.389306, 7.372664, 
    6.355908, 4.89603, 3.593253, 2.724032, 3.681464, 5.650462, 7.344178, 
    6.978189,
  3.133896, 4.079565, 5.329723, 7.428953, 8.923047, 8.948499, 8.393973, 
    7.00301, 5.895844, 4.757103, 3.384584, 3.168375, 5.46642, 7.440119, 
    7.587461,
  3.533773, 4.252082, 5.793657, 8.117177, 9.650985, 9.636585, 8.652927, 
    6.373183, 5.77106, 4.928487, 3.313741, 3.154536, 5.261129, 7.28497, 
    7.668458,
  3.573808, 3.954098, 5.501093, 8.180192, 9.947165, 10.16742, 9.327611, 
    7.2477, 5.756925, 5.121824, 3.532803, 3.54726, 5.374897, 7.187072, 
    7.789378,
  3.998962, 3.810606, 5.52222, 8.659118, 10.82462, 11.13792, 10.27442, 
    8.24513, 5.253314, 4.084838, 3.766505, 4.627475, 6.010468, 7.320277, 
    7.452598,
  4.593127, 5.074707, 2.829183, 3.132869, 3.529236, 3.273968, 4.066905, 
    3.635206, 3.582778, 3.031706, 3.436708, 3.918738, 3.376921, 2.220147, 
    1.807525,
  4.498754, 3.221072, 3.589457, 4.204761, 3.767017, 3.6548, 4.80493, 
    3.969554, 3.450287, 3.345849, 3.471351, 5.06222, 5.182308, 2.747345, 
    2.018504,
  3.032837, 3.294162, 4.384931, 5.314302, 4.478287, 4.144092, 4.083385, 
    3.87234, 3.631629, 3.751463, 4.271932, 5.895147, 6.059231, 4.322983, 
    2.739554,
  2.558171, 4.093118, 5.507698, 6.825188, 6.984971, 4.779856, 2.739717, 
    2.454788, 3.162791, 3.513704, 4.749067, 6.236986, 6.512786, 5.009397, 
    3.172538,
  2.782366, 4.510483, 6.428663, 7.508706, 8.055825, 5.857471, 3.00889, 
    2.584203, 2.635954, 2.77189, 5.345867, 6.559332, 7.024455, 5.780061, 
    4.02284,
  2.910197, 4.855429, 6.905313, 7.832013, 8.01616, 6.834067, 3.534248, 
    4.073774, 4.432196, 4.521874, 4.601462, 6.743392, 7.141952, 6.117825, 
    4.666445,
  3.274265, 5.305025, 6.869614, 7.855854, 7.984631, 7.089448, 5.770415, 
    4.831483, 6.657166, 6.610988, 6.302245, 7.137002, 7.444102, 6.716065, 
    5.443997,
  3.94106, 5.793549, 6.707504, 7.750443, 8.13084, 7.847519, 6.955901, 
    6.612029, 6.856847, 6.315151, 6.494046, 7.421209, 7.583839, 7.03123, 
    5.85858,
  4.553251, 5.828889, 6.401479, 7.339746, 7.756388, 7.778035, 7.255027, 
    6.620713, 6.167236, 5.627468, 6.346132, 7.734414, 7.794248, 7.138212, 
    5.852251,
  4.873408, 5.644233, 6.600768, 7.687816, 7.825012, 7.374688, 6.755183, 
    5.911225, 4.62433, 4.15536, 5.422693, 8.122777, 7.692417, 6.969933, 
    5.612424,
  2.112349, 1.938897, 1.765726, 3.007736, 3.607843, 3.383726, 3.611677, 
    3.124149, 2.323736, 2.529611, 3.153374, 2.56186, 1.154825, 1.660343, 
    3.134291,
  2.431624, 2.215174, 2.644233, 3.530991, 3.187398, 2.594927, 3.118295, 
    2.937578, 3.073661, 3.252403, 3.464662, 3.323867, 1.620951, 1.718469, 
    3.213398,
  2.929339, 2.28373, 2.808897, 3.442934, 2.92259, 2.292918, 1.253935, 
    2.495476, 3.680459, 4.25955, 4.613438, 3.831308, 2.004441, 2.945107, 
    3.559594,
  2.716973, 2.317202, 3.038785, 3.718026, 3.317595, 1.421009, 1.214193, 
    3.20164, 3.645521, 4.195246, 5.136121, 3.951216, 2.658972, 3.700219, 
    3.581654,
  3.203964, 3.193929, 3.749726, 4.000719, 3.304827, 1.494517, 2.019152, 
    2.985132, 2.949565, 3.444325, 4.869134, 3.51046, 3.16042, 3.6133, 3.604018,
  4.215957, 4.178389, 4.380737, 4.73728, 4.605488, 3.905914, 3.469256, 
    4.518987, 4.673696, 4.869235, 3.699721, 4.00953, 3.691201, 3.976868, 
    5.136459,
  5.293286, 5.105473, 4.723985, 5.308014, 5.684165, 6.054245, 6.177609, 
    6.432252, 7.134417, 6.768421, 5.680859, 5.13605, 5.160396, 6.101845, 
    7.085255,
  6.180939, 5.533978, 4.757706, 5.41505, 5.864539, 6.366319, 6.953441, 
    7.460179, 7.660124, 7.539793, 7.157724, 6.987378, 7.139089, 7.300676, 
    7.262776,
  6.645617, 5.55127, 4.867862, 5.394397, 6.046981, 6.633699, 7.160275, 
    7.644794, 7.972369, 7.876359, 7.823992, 7.867248, 7.747328, 7.659399, 
    6.848152,
  6.783386, 5.864025, 5.347458, 5.271443, 5.666945, 6.363478, 7.155316, 
    7.350777, 6.694509, 5.625304, 6.275286, 8.093423, 8.02153, 8.098676, 
    7.518355,
  5.323083, 6.547487, 5.45559, 5.773393, 4.494079, 3.247134, 3.727078, 
    3.38602, 1.75193, 0.4886339, 2.01238, 2.210936, 1.030248, 2.52713, 
    4.144566,
  8.345502, 7.513963, 5.910537, 4.555771, 2.687877, 2.226647, 3.644198, 
    3.457841, 2.489383, 1.120707, 1.519376, 1.480535, 1.29069, 2.536952, 
    4.44015,
  9.225501, 7.107168, 5.01255, 3.309081, 2.239658, 1.339236, 1.905803, 
    3.369461, 3.041189, 2.290324, 2.03644, 1.76213, 1.869601, 4.149532, 
    5.430993,
  8.716697, 6.133072, 3.624037, 2.211602, 2.323681, 1.456449, 0.9135218, 
    2.475263, 2.673128, 2.495208, 2.69638, 2.222168, 3.483416, 5.957811, 
    5.33309,
  7.802373, 5.197698, 2.733415, 1.621115, 1.725087, 2.182214, 1.578119, 
    1.877507, 2.085502, 1.929093, 2.625328, 2.593348, 4.748963, 6.040844, 
    4.535234,
  7.083781, 4.963465, 3.171259, 2.200475, 1.734929, 1.778754, 1.953367, 
    2.165243, 2.282483, 2.014568, 1.345366, 2.905423, 4.803412, 4.01893, 
    2.503887,
  6.672111, 5.107272, 3.578007, 2.925256, 2.974498, 3.277131, 3.269618, 
    2.453985, 1.912932, 2.082134, 2.76304, 3.444835, 3.222574, 2.305282, 
    3.39055,
  6.313592, 5.131826, 3.769, 3.315205, 3.236792, 3.044706, 2.912228, 
    2.444618, 2.155585, 2.42624, 2.993462, 3.111759, 2.5107, 3.674245, 
    5.255366,
  6.613481, 5.810369, 4.977878, 4.545085, 4.115565, 3.528343, 3.35208, 
    3.157401, 3.158082, 3.301092, 3.54069, 3.554394, 4.45442, 5.541081, 
    5.997453,
  7.168694, 6.748442, 6.243951, 5.765567, 5.314854, 4.573498, 4.395575, 
    3.969903, 3.410305, 2.950871, 3.758171, 5.870842, 6.393638, 6.925784, 
    7.378078,
  4.492879, 6.433449, 7.76363, 11.72882, 11.37677, 8.596026, 9.78044, 
    8.486322, 5.825492, 3.542471, 2.935062, 2.703412, 2.132231, 2.76632, 
    3.964048,
  7.25491, 9.197427, 10.8113, 13.05062, 9.334537, 7.148826, 8.657099, 
    7.445328, 4.729696, 2.768892, 1.851113, 1.929201, 2.750225, 3.308379, 
    5.005332,
  9.133286, 10.37429, 11.49125, 11.67111, 8.263697, 6.10818, 6.297534, 
    5.880544, 4.005445, 2.244102, 1.028944, 2.146568, 3.810201, 6.089744, 
    6.558998,
  10.80422, 10.92151, 10.69419, 9.583282, 8.033422, 6.225557, 4.681412, 
    3.753198, 2.82775, 2.396253, 2.491693, 3.454337, 5.575734, 8.039979, 
    6.239913,
  10.9298, 9.879169, 8.806252, 7.58128, 6.060916, 5.558741, 5.312748, 
    3.451055, 2.170838, 2.142968, 2.676457, 4.133526, 6.447542, 8.393238, 
    5.89833,
  9.60912, 8.315928, 6.860953, 5.413033, 5.005381, 4.45375, 4.302803, 
    3.793687, 2.180811, 1.483281, 1.451653, 4.567258, 7.31517, 6.585628, 
    3.365438,
  7.406801, 6.300727, 4.731768, 3.215047, 3.587983, 4.155447, 3.711793, 
    2.847689, 2.703008, 1.982354, 2.494646, 5.964189, 6.285355, 3.166959, 
    3.56909,
  4.813438, 3.777536, 2.545421, 2.09554, 2.730744, 3.716673, 4.465297, 
    4.513498, 3.074902, 1.642556, 4.473336, 5.8209, 3.281438, 3.014512, 
    5.099977,
  3.12783, 2.373512, 2.308245, 2.251225, 2.797329, 3.538068, 4.328125, 
    4.173468, 2.396126, 3.037446, 4.732606, 3.090226, 2.614494, 4.889056, 
    6.427299,
  2.844944, 2.6435, 2.811254, 2.899779, 3.174659, 3.664759, 4.474132, 
    3.830334, 2.577326, 2.490495, 2.144869, 2.316149, 4.677498, 6.607718, 
    8.245794,
  3.350342, 5.208306, 6.038963, 8.616463, 8.686428, 8.7562, 12.02026, 
    11.78938, 10.21155, 7.068875, 5.923479, 4.519629, 2.785463, 1.654064, 
    1.48364,
  5.3555, 7.510163, 9.335673, 11.29968, 9.899303, 9.979164, 12.57156, 
    11.65946, 9.93343, 7.819829, 5.194863, 3.840545, 2.149468, 1.291052, 
    2.044202,
  6.043754, 8.786137, 11.02838, 13.63931, 11.7241, 10.39064, 10.38643, 
    10.4472, 9.45225, 6.848524, 3.904366, 2.180785, 2.402987, 4.099425, 
    3.779627,
  7.582534, 10.77722, 12.95332, 13.91485, 13.88465, 11.52383, 8.989481, 
    7.405899, 5.563577, 2.973212, 1.481692, 2.611008, 4.956118, 6.281328, 
    4.583825,
  9.399341, 11.84604, 13.312, 13.48678, 12.35805, 11.5807, 9.717013, 
    5.986004, 2.646849, 1.27721, 1.314972, 4.460739, 6.437719, 6.547581, 
    4.211971,
  10.85648, 12.65913, 13.33466, 13.27221, 12.25133, 9.212277, 6.898428, 
    6.391608, 3.825391, 2.255361, 2.226424, 6.236782, 6.470547, 4.483719, 
    1.901668,
  11.71817, 13.01267, 13.22054, 12.7942, 11.27023, 9.183258, 7.193345, 
    6.416307, 5.320942, 3.260052, 4.776575, 6.157645, 4.704956, 2.911617, 
    3.046642,
  11.7401, 12.48563, 12.17059, 11.39424, 10.24799, 9.05962, 8.061252, 6.9768, 
    4.076562, 3.067142, 5.769854, 5.26148, 3.317932, 3.028853, 3.943807,
  10.64422, 11.24398, 10.80005, 10.00642, 9.313128, 8.498592, 7.070443, 
    4.675784, 2.478216, 4.377243, 5.805562, 4.131948, 2.710633, 3.102617, 
    4.122482,
  9.296144, 9.909732, 9.565985, 8.769542, 8.302839, 7.68655, 5.994524, 
    3.138779, 2.053572, 3.458204, 3.645, 2.623274, 3.120944, 4.449511, 
    6.079962,
  5.307834, 7.689221, 7.622944, 9.7141, 8.68327, 7.380922, 9.327675, 
    10.15812, 9.891477, 8.08188, 7.439319, 6.788157, 5.105536, 3.205649, 
    1.69473,
  5.611659, 7.56321, 9.22979, 10.10778, 8.226689, 7.674519, 9.963756, 
    10.82749, 10.81592, 9.580626, 7.658125, 7.511306, 5.391117, 2.318782, 
    1.142509,
  5.429908, 7.922499, 9.628836, 11.59921, 9.594709, 9.251943, 9.762693, 
    11.10141, 11.57088, 10.15805, 8.61991, 6.21192, 3.881357, 2.844165, 
    2.097631,
  7.768142, 9.288099, 9.966231, 11.23137, 11.35087, 11.46286, 10.1517, 
    9.455685, 8.641166, 6.929673, 5.737508, 4.211576, 3.863485, 4.763323, 
    4.456717,
  8.752702, 9.784859, 10.36541, 11.71821, 12.05754, 11.72865, 10.18772, 
    7.656278, 4.667713, 3.585036, 4.174286, 4.538383, 5.643821, 6.604434, 
    6.9301,
  9.59452, 10.52079, 10.773, 12.48745, 12.13482, 9.108303, 7.285314, 
    8.210038, 6.301459, 3.836416, 2.390356, 4.6243, 5.885256, 4.945672, 
    4.600136,
  10.02547, 11.35627, 12.34851, 12.92678, 12.12183, 10.40443, 9.057784, 
    8.124415, 6.617699, 3.035604, 2.574009, 3.151957, 2.805465, 1.854979, 
    2.43291,
  11.29556, 12.68254, 12.9415, 12.74332, 11.71804, 10.57476, 9.650527, 
    7.645362, 4.509909, 2.370878, 1.807746, 1.807232, 1.990548, 2.168762, 
    2.539461,
  12.91545, 13.71483, 13.38867, 12.56792, 11.47421, 9.834125, 7.635831, 
    5.533505, 4.10456, 3.548961, 3.344698, 2.853104, 2.432015, 2.437912, 
    2.866537,
  13.95029, 14.13318, 13.29822, 12.03456, 10.32614, 8.354545, 6.305112, 
    4.951518, 3.538447, 2.610122, 2.714729, 3.32082, 3.021569, 3.684152, 
    4.939462,
  7.526241, 7.237547, 4.913599, 3.717779, 4.881094, 4.999369, 5.297647, 
    4.777257, 5.927516, 6.466885, 7.492273, 8.225288, 7.706977, 5.316778, 
    3.641923,
  10.49711, 9.152086, 7.659022, 5.21232, 3.660429, 3.583177, 4.731077, 
    5.248475, 5.314406, 6.421004, 7.767774, 9.471597, 9.949802, 5.421128, 
    3.854753,
  8.408777, 8.981205, 8.058387, 6.840285, 4.497072, 2.910816, 2.926933, 
    4.303191, 5.419873, 7.577154, 9.452744, 9.979228, 9.779704, 7.319693, 
    5.187578,
  8.334959, 8.723668, 8.020819, 7.08527, 5.888256, 4.187221, 2.952271, 
    4.458419, 5.933664, 5.969016, 9.507608, 10.72703, 9.22171, 7.135568, 
    5.136609,
  9.621422, 8.907662, 8.206658, 7.200862, 6.004178, 5.434869, 5.187474, 
    4.377917, 3.655417, 4.096328, 8.672186, 10.30171, 8.913139, 7.125668, 
    5.653861,
  11.07155, 9.748174, 8.56524, 7.343872, 6.000964, 5.070413, 5.016436, 
    6.618071, 6.239886, 6.766042, 6.933266, 9.174501, 7.758317, 6.386684, 
    5.192681,
  11.42555, 10.55178, 9.491512, 8.499122, 7.986619, 7.880147, 8.305653, 
    9.156181, 10.26504, 9.869476, 8.982243, 7.327109, 5.544071, 4.290128, 
    3.710449,
  11.92553, 11.81993, 11.26685, 11.04438, 11.1989, 11.55454, 11.74076, 
    11.36943, 10.16096, 8.390798, 6.462622, 4.369446, 3.246639, 2.380667, 
    2.091633,
  11.96248, 12.18665, 12.01363, 11.97761, 11.73215, 11.22076, 10.24617, 
    9.023, 7.407491, 5.753458, 4.044907, 3.276837, 2.917262, 1.851512, 
    1.195624,
  11.50305, 11.76998, 11.78285, 11.25272, 10.46975, 9.729711, 8.643811, 
    7.310935, 5.198575, 3.480392, 3.444107, 4.661504, 4.302035, 3.258085, 
    2.805991,
  2.775185, 2.917824, 1.746094, 2.980581, 5.625031, 5.513534, 7.09855, 
    7.635716, 7.122707, 5.290862, 5.582362, 5.909791, 6.439266, 5.463192, 
    3.993279,
  5.283486, 3.888653, 2.087459, 3.269582, 4.289331, 5.305911, 7.657098, 
    7.789406, 7.909644, 7.392296, 6.806741, 7.574872, 8.478504, 5.611314, 
    5.121096,
  5.553885, 4.30358, 3.835726, 5.100145, 4.684995, 5.183946, 6.594779, 
    7.320766, 8.085533, 8.609184, 8.70574, 8.567899, 8.700787, 8.671327, 
    6.94019,
  5.488324, 4.842212, 4.946596, 5.928045, 6.545852, 5.510627, 5.21764, 
    5.897007, 6.834455, 7.679961, 9.209903, 9.566014, 9.291985, 9.03583, 
    7.329372,
  5.362506, 4.960872, 5.028304, 5.274485, 5.544338, 7.001375, 5.900908, 
    5.005644, 4.132093, 4.765216, 8.547848, 10.16649, 10.53114, 9.630301, 
    7.731281,
  5.255696, 5.200638, 5.220131, 5.081663, 4.868718, 5.731453, 6.00887, 
    4.752025, 4.232653, 5.604672, 7.213036, 10.74067, 10.57784, 9.220948, 
    7.041637,
  5.762497, 6.125134, 6.05367, 6.334447, 6.536511, 6.609125, 6.704527, 
    6.584285, 7.490578, 9.144408, 10.31174, 11.23734, 10.50544, 8.979618, 
    7.222423,
  7.868483, 8.690602, 8.761815, 9.624242, 10.41031, 10.4961, 10.42792, 
    10.56252, 10.68561, 10.94197, 10.95002, 10.67942, 9.49915, 8.061516, 
    6.639201,
  10.26575, 10.68256, 11.03351, 11.87033, 12.45729, 12.77293, 12.67363, 
    12.1485, 11.56225, 10.61618, 9.979596, 9.405378, 8.292573, 6.856054, 
    5.544287,
  10.56089, 10.61128, 10.98563, 11.06623, 11.25851, 11.35075, 11.32848, 
    10.91902, 8.958592, 6.682334, 6.698585, 7.867575, 6.573941, 5.267165, 
    4.123254,
  3.474753, 4.03143, 3.61297, 4.792715, 4.522716, 3.701345, 4.296802, 
    5.308021, 5.976187, 3.147759, 1.533848, 2.516747, 4.161571, 4.225686, 
    3.292921,
  6.068634, 6.142813, 5.692944, 5.527792, 3.549018, 3.501865, 4.929893, 
    5.438673, 6.058026, 4.142796, 1.442838, 2.664692, 5.2005, 4.064755, 
    3.833578,
  7.607922, 7.637062, 7.458606, 7.411335, 5.559192, 4.101174, 4.206063, 
    5.633392, 6.764155, 5.194894, 2.338679, 2.716835, 4.377849, 5.963567, 
    5.901174,
  8.81743, 8.713732, 8.180127, 8.840391, 10.11609, 7.330832, 4.866857, 
    4.457161, 5.576282, 4.670491, 3.037865, 2.787762, 4.038094, 6.049178, 
    6.69073,
  10.35898, 9.84794, 8.794621, 7.714772, 10.6164, 11.21926, 9.345628, 
    6.765659, 4.485798, 3.19539, 3.672823, 3.478301, 4.557477, 7.062501, 
    9.156579,
  11.62296, 11.15017, 9.368301, 4.892226, 9.188533, 12.13107, 11.08555, 
    9.318898, 6.086436, 4.301757, 3.350479, 4.44818, 5.385212, 7.165557, 
    8.21145,
  12.52827, 12.45267, 9.601436, 5.149517, 8.509732, 11.91973, 10.20848, 
    7.908988, 7.060442, 6.351167, 5.486054, 5.70435, 6.413223, 7.563715, 
    8.043307,
  12.96172, 13.46305, 11.47878, 8.597486, 10.17907, 11.18448, 9.688319, 
    8.886436, 7.793475, 6.538233, 5.887767, 6.460299, 7.090076, 8.111259, 
    8.338476,
  12.59676, 13.68254, 12.92204, 11.73626, 11.65816, 11.19165, 9.675533, 
    8.464055, 7.507902, 6.600886, 6.50205, 7.328193, 8.064488, 8.816447, 
    8.544014,
  11.35092, 13.34006, 14.06527, 13.11353, 11.84958, 10.89121, 9.806964, 
    8.713435, 6.831774, 5.023928, 5.552676, 8.229177, 8.6334, 8.820601, 
    7.682074,
  3.401387, 4.799524, 4.998209, 6.078526, 5.66992, 4.647433, 5.394286, 
    5.041995, 4.496493, 3.719604, 2.720994, 2.499259, 2.566438, 2.869145, 
    3.320728,
  6.023068, 7.245213, 7.604006, 7.687506, 4.74919, 4.038935, 5.459596, 
    4.806417, 4.821895, 4.230046, 2.23188, 2.709743, 3.970801, 3.321084, 
    3.973204,
  7.291216, 8.892542, 8.967738, 8.243851, 5.659421, 4.175705, 3.968385, 
    3.966854, 4.185298, 4.115258, 2.124917, 2.641604, 4.525533, 5.477861, 
    6.610081,
  8.944961, 9.966869, 9.834556, 8.9939, 8.546962, 6.012475, 3.395938, 
    1.705111, 2.641578, 2.639133, 1.630827, 2.882981, 4.676459, 6.273156, 
    7.536399,
  10.50753, 10.64167, 10.37319, 9.196906, 8.716568, 8.842624, 6.916265, 
    3.754986, 2.162327, 1.709227, 1.882211, 3.263948, 5.726909, 7.984727, 
    9.745482,
  10.94326, 10.70656, 9.610979, 8.509042, 8.210636, 8.889717, 8.902181, 
    6.590706, 3.745441, 2.553494, 1.751889, 4.125323, 7.079236, 8.360414, 
    8.421423,
  10.9354, 10.42124, 7.964578, 6.266479, 7.181136, 8.60927, 8.203122, 
    5.25493, 4.187626, 3.781818, 3.039828, 5.865248, 7.525175, 8.315766, 
    8.487534,
  10.57152, 9.63395, 5.814607, 2.792288, 6.995783, 9.056296, 8.712554, 
    6.754275, 5.431685, 4.096931, 4.446428, 6.635538, 7.53808, 8.418462, 
    8.991082,
  10.25154, 9.54628, 6.980147, 6.535919, 9.024757, 9.564078, 8.338859, 
    6.484004, 5.737754, 4.848068, 5.348483, 6.889003, 7.924553, 9.142179, 
    9.436306,
  9.27603, 9.409713, 9.300041, 9.21309, 9.251458, 8.930807, 7.924055, 
    7.139286, 5.321671, 3.727863, 4.328834, 6.857671, 8.261016, 9.399374, 
    8.371819,
  3.006135, 4.124927, 3.927167, 5.014788, 4.867869, 4.740211, 6.50417, 
    6.965465, 6.875519, 5.337157, 5.605123, 5.746657, 4.917598, 4.230541, 
    3.955782,
  3.519307, 4.0101, 4.527236, 5.289698, 3.879048, 4.286747, 7.163624, 
    7.425045, 7.560474, 6.754385, 6.128335, 6.518106, 5.7101, 3.889907, 
    3.899985,
  2.880117, 3.733949, 5.278544, 6.434294, 5.325291, 4.597637, 5.824998, 
    7.099271, 7.338202, 6.970058, 6.856325, 6.515921, 5.860122, 5.290824, 
    4.135547,
  4.955483, 7.262222, 8.642375, 9.233256, 9.509992, 7.329875, 4.692343, 
    3.856311, 5.313264, 5.996239, 5.702863, 5.185871, 4.759024, 4.388706, 
    4.027902,
  8.882757, 9.896937, 10.36273, 10.24376, 10.17361, 10.00041, 7.982892, 
    4.641161, 3.179333, 2.839556, 3.228874, 3.740078, 3.482846, 4.308908, 
    5.62497,
  10.05221, 10.00775, 9.586461, 9.440598, 9.446986, 9.484324, 9.901513, 
    8.893309, 4.272437, 2.597857, 2.84728, 4.253334, 4.096179, 5.899557, 
    6.333845,
  9.309406, 8.486599, 7.797218, 7.053235, 7.272843, 7.616357, 7.826637, 
    7.328125, 5.71084, 5.384355, 5.826317, 4.815242, 6.363375, 7.066927, 
    8.355978,
  7.70793, 7.470363, 5.633401, 3.642552, 3.818337, 5.482789, 6.309928, 
    6.140309, 5.447157, 5.578964, 4.697579, 6.202789, 7.736673, 8.950753, 
    10.57773,
  7.013495, 6.398411, 5.26811, 4.039137, 4.213778, 5.327099, 5.640692, 
    4.369602, 3.605803, 3.595146, 5.538477, 8.392316, 9.809714, 11.18912, 
    10.84591,
  6.065263, 6.260602, 6.054527, 5.466807, 4.979349, 4.873323, 4.182468, 
    3.052818, 2.438024, 3.288848, 6.758769, 10.36036, 10.71399, 10.83041, 
    9.498553,
  4.771297, 5.949106, 5.023509, 6.229692, 5.449824, 4.035744, 5.012703, 
    4.628866, 3.813023, 2.893858, 2.82701, 2.773844, 3.60579, 5.645966, 
    7.049871,
  6.757607, 6.791123, 6.209363, 6.189419, 4.560802, 3.596622, 4.863028, 
    4.686846, 4.255019, 3.765617, 2.78407, 3.077784, 5.096293, 5.588117, 
    7.706246,
  7.650397, 7.089321, 5.870754, 5.525173, 4.86857, 3.644294, 3.756277, 
    5.081248, 5.348271, 4.457025, 3.44089, 4.22905, 6.102228, 7.587686, 
    8.150611,
  7.952559, 6.06117, 5.626781, 5.469392, 5.68918, 5.008163, 3.657321, 
    3.124814, 4.282526, 4.57151, 4.282172, 3.970725, 4.565882, 6.756877, 
    6.686429,
  5.407135, 5.529634, 5.854462, 5.981646, 6.046612, 6.716352, 6.582891, 
    4.765185, 3.114243, 2.752347, 3.145581, 1.897676, 2.411053, 5.718931, 
    5.903516,
  4.664464, 4.8297, 5.366481, 5.856351, 6.425826, 6.927681, 8.215537, 
    8.86484, 5.270947, 3.002533, 2.44902, 2.46829, 2.399898, 4.939703, 
    4.703473,
  5.351723, 4.886478, 5.206175, 5.956482, 6.73502, 7.082877, 7.439281, 
    7.771141, 6.7937, 5.499582, 4.87675, 3.715677, 1.741023, 3.540948, 
    5.372167,
  5.445718, 5.405824, 5.626616, 6.256125, 6.592615, 6.874523, 7.275496, 
    8.053418, 8.352966, 6.994541, 5.895192, 4.14114, 1.775428, 3.206836, 
    6.805009,
  6.080042, 6.42066, 6.407734, 6.309405, 5.47905, 5.430425, 6.60751, 
    7.614252, 8.203394, 7.689709, 6.755205, 4.499308, 2.806082, 5.298325, 
    7.330272,
  6.889575, 7.500194, 6.26756, 4.844078, 3.857524, 4.526871, 6.228007, 
    7.719975, 7.361559, 5.608391, 5.159583, 4.906621, 4.632962, 7.199097, 
    8.112029,
  8.764199, 7.877611, 3.822595, 6.283848, 6.7219, 7.304638, 11.16217, 
    10.94514, 9.575599, 8.034684, 7.199025, 5.285167, 3.382046, 3.426749, 
    3.535747,
  11.09461, 7.344759, 5.278272, 7.617711, 6.763711, 7.394744, 10.34596, 
    10.68228, 10.42392, 9.744804, 7.116471, 5.4765, 4.108067, 2.740862, 
    3.131847,
  11.55522, 7.387227, 5.737859, 8.224138, 7.91221, 7.439523, 7.953716, 
    9.52312, 10.98675, 9.61219, 6.706225, 4.53324, 3.87944, 3.923696, 3.331713,
  13.95558, 8.540824, 5.74445, 8.3228, 9.248665, 8.835874, 8.230157, 
    8.266933, 8.645768, 6.557708, 5.270415, 3.559714, 3.500555, 4.19592, 
    3.542605,
  13.78609, 11.08038, 5.937087, 8.553916, 8.92709, 9.68792, 10.15031, 
    8.102933, 4.677975, 3.215854, 4.056982, 3.150974, 3.295597, 4.016831, 
    4.453091,
  10.70099, 11.17075, 7.400594, 8.373795, 8.566898, 8.252116, 8.334518, 
    8.139454, 5.852145, 4.594676, 3.669826, 3.87785, 3.53408, 4.359591, 
    5.513425,
  6.511325, 8.523251, 7.165061, 7.074338, 7.486809, 7.515647, 6.658889, 
    6.399565, 7.071671, 6.789527, 5.755173, 4.300159, 4.09647, 5.549392, 
    6.638815,
  3.05358, 5.153729, 5.663061, 5.855079, 6.63325, 7.132846, 7.279863, 
    7.49727, 7.583908, 6.752384, 5.65288, 4.425648, 4.613679, 5.595643, 
    5.959683,
  2.464071, 3.039056, 4.455592, 5.464352, 6.191049, 6.844649, 6.970182, 
    6.994821, 7.271744, 6.26518, 5.340816, 4.75932, 4.806981, 4.995825, 
    4.843226,
  3.597784, 3.944723, 4.817676, 5.82425, 6.345942, 6.919253, 7.383012, 
    7.608333, 6.376141, 4.334155, 4.166292, 5.222756, 4.974719, 5.256585, 
    5.723138,
  6.341107, 10.83976, 8.823115, 8.45902, 6.418128, 5.029895, 8.196727, 
    10.25821, 10.51389, 8.505161, 8.62526, 8.035576, 6.744782, 5.339475, 
    3.804637,
  8.181557, 10.53881, 9.140781, 7.629435, 7.155796, 7.540196, 10.86221, 
    10.97253, 10.91008, 9.448105, 8.784444, 8.567597, 7.219652, 3.960924, 
    2.651301,
  7.495365, 10.00955, 7.287779, 6.17613, 6.74229, 6.471496, 9.245654, 
    10.93628, 11.83895, 10.6849, 9.28597, 8.008835, 6.425981, 4.450497, 
    3.078124,
  7.042449, 9.210582, 5.427816, 5.182, 7.255434, 6.085771, 6.787819, 
    9.385942, 10.59398, 8.583773, 8.145993, 7.170505, 6.341466, 5.249379, 
    4.17452,
  6.544911, 7.827337, 3.895379, 4.754435, 6.48583, 6.094203, 5.155256, 
    5.562873, 4.656131, 4.46014, 6.416672, 6.716185, 6.606447, 6.119861, 
    5.711893,
  6.064644, 6.82529, 3.312964, 4.356499, 5.873203, 4.8548, 4.45834, 6.34875, 
    6.056769, 4.926392, 4.923239, 6.847845, 6.498847, 6.422534, 6.095851,
  5.48048, 6.190969, 3.048249, 4.740534, 6.230367, 5.760315, 6.464291, 
    7.865478, 7.731878, 7.204741, 7.013679, 6.785767, 6.148965, 5.487364, 
    5.142855,
  4.501649, 5.534325, 3.030907, 5.187149, 7.428945, 7.269705, 8.378889, 
    9.425632, 8.847477, 7.961762, 6.956933, 6.220843, 5.152202, 4.328479, 
    3.843132,
  3.320643, 4.420231, 3.143526, 5.021569, 8.350395, 8.55103, 9.314709, 
    9.098018, 8.541685, 7.377637, 6.201391, 5.211763, 4.265819, 3.73057, 
    3.515331,
  2.11459, 3.172889, 3.814344, 4.669136, 8.963868, 9.932427, 10.45922, 
    9.417968, 7.040546, 4.769721, 4.464002, 4.746527, 4.236407, 4.254245, 
    4.433413,
  4.895441, 5.457362, 4.031568, 4.493909, 3.857341, 3.617407, 5.290527, 
    5.984023, 6.37107, 5.144282, 5.409388, 5.639904, 5.631036, 5.592321, 
    5.372873,
  8.102873, 7.298892, 5.954859, 5.377881, 4.063879, 4.190941, 6.227142, 
    6.444605, 6.539688, 5.88177, 6.027861, 6.581379, 6.318485, 4.006005, 
    3.662915,
  9.121426, 8.567737, 7.455547, 6.736969, 5.518513, 4.586431, 5.630278, 
    6.667044, 6.962353, 6.561688, 6.562931, 6.822064, 6.514612, 5.091942, 
    3.339982,
  10.98028, 10.25864, 8.935369, 8.235326, 7.877962, 6.551228, 5.26802, 
    5.207098, 5.47281, 5.237845, 6.260062, 6.594309, 6.208323, 5.437226, 
    4.132678,
  12.33615, 11.14355, 10.11714, 9.42401, 8.550694, 8.181841, 6.777822, 
    4.605456, 3.437151, 3.667571, 5.783823, 6.136298, 5.606153, 5.140803, 
    4.397835,
  12.36541, 11.39334, 10.79798, 10.13558, 9.339741, 7.896911, 6.313283, 
    5.731121, 5.243187, 5.344291, 4.600097, 5.599951, 4.403528, 3.585338, 
    2.895682,
  11.13799, 10.48782, 10.51179, 10.64107, 9.75931, 8.128725, 6.452934, 
    5.876254, 7.308482, 7.705529, 6.22604, 4.935259, 3.044804, 2.082412, 
    2.440267,
  10.26757, 9.168105, 8.163693, 9.404113, 9.871246, 8.931346, 8.622907, 
    8.781632, 8.913465, 8.094223, 6.12072, 4.054743, 2.287678, 1.963428, 
    2.455557,
  8.219985, 7.811659, 6.362936, 7.928233, 10.07164, 9.425247, 9.13597, 
    9.001863, 9.037432, 7.344121, 5.119528, 3.284714, 2.222678, 2.597287, 
    2.76496,
  5.468838, 6.100594, 4.881977, 7.096457, 9.525796, 9.74007, 9.873559, 
    9.686917, 7.647559, 4.871364, 3.827992, 3.247207, 2.481851, 3.314687, 
    3.656773,
  4.856919, 5.958483, 5.300701, 5.3798, 3.783406, 2.76229, 3.330795, 
    3.144691, 3.382277, 2.92728, 3.252316, 3.177695, 2.984639, 2.936482, 
    3.097259,
  6.451963, 5.960823, 5.993693, 5.053934, 3.156441, 2.644112, 3.909877, 
    4.016714, 4.257825, 3.954369, 4.310053, 4.560706, 4.006134, 2.129683, 
    1.725881,
  5.880063, 5.197948, 4.845639, 4.381755, 3.0066, 2.523216, 3.56987, 
    4.446575, 5.119485, 5.123972, 5.747009, 5.815612, 4.426738, 3.252071, 
    2.241172,
  4.473745, 4.154109, 4.345843, 4.675807, 4.20635, 3.647499, 3.448128, 
    3.735668, 4.478722, 5.01586, 5.904694, 6.210719, 5.162748, 4.021371, 
    3.07535,
  3.681, 4.737454, 6.289669, 6.7519, 6.910068, 6.755624, 6.123393, 4.313725, 
    3.988552, 3.810951, 6.034224, 6.642538, 6.113847, 5.009855, 3.736877,
  5.908927, 7.572368, 8.816413, 9.374795, 9.498336, 9.725106, 9.605769, 
    9.472946, 6.600896, 5.38523, 5.160168, 7.16326, 6.667161, 5.208774, 
    2.838696,
  8.179172, 9.731719, 10.82516, 11.30585, 11.5391, 10.96843, 11.1731, 
    9.927972, 9.069762, 9.173327, 8.463593, 7.938223, 6.968513, 4.792111, 
    2.549035,
  9.874085, 11.24985, 12.29174, 12.82271, 12.90779, 12.52697, 12.52957, 
    11.13676, 10.71719, 10.27648, 9.23417, 8.477435, 6.964707, 4.462785, 
    2.284553,
  10.45598, 12.26689, 12.51635, 13.77858, 13.29644, 13.64802, 13.08269, 
    11.76047, 11.20545, 10.47052, 9.786209, 8.750044, 6.731177, 4.37383, 
    2.644032,
  9.567395, 11.08139, 12.63369, 11.75156, 10.70997, 10.87275, 12.05752, 
    12.47425, 10.39009, 8.150321, 8.087931, 8.692059, 6.059055, 4.573244, 
    3.363755,
  5.095816, 6.669696, 5.48365, 6.68114, 5.581913, 4.654222, 5.635038, 
    3.970187, 2.822906, 2.001362, 2.228679, 3.22207, 4.087158, 3.421025, 
    1.853695,
  8.901944, 9.727968, 9.809859, 9.247342, 7.05416, 6.200647, 7.113941, 
    5.616723, 4.290644, 3.560037, 3.459509, 3.277899, 4.367136, 3.672973, 
    2.651763,
  11.78589, 11.55759, 10.52633, 8.44801, 5.23056, 3.177397, 3.389716, 
    2.685423, 2.528389, 3.13956, 3.811212, 4.419418, 4.641477, 5.053554, 
    3.96506,
  10.46747, 9.758495, 8.286391, 6.506525, 4.470928, 2.521685, 1.607154, 
    2.395563, 1.769274, 2.3436, 3.154191, 4.202782, 5.124385, 5.318207, 
    4.902085,
  6.842549, 5.531592, 4.41431, 3.797505, 3.521644, 3.275235, 3.379689, 
    2.056691, 1.650301, 1.720141, 2.980837, 3.81841, 5.237499, 5.746255, 
    6.176231,
  3.300912, 3.601396, 3.945282, 4.438937, 5.157836, 6.108057, 7.313029, 
    8.219937, 5.837998, 3.944988, 3.160258, 3.476887, 4.337955, 4.928586, 
    5.687095,
  3.242043, 4.048459, 4.761926, 5.840171, 7.247582, 8.481062, 9.871485, 
    10.74615, 9.831508, 8.355762, 6.278503, 3.880922, 3.668633, 4.827628, 
    6.072401,
  3.911315, 5.446394, 6.135077, 7.336526, 8.893971, 10.16903, 11.4873, 
    11.54181, 11.05684, 9.739491, 7.462476, 4.661253, 4.179734, 5.949833, 
    6.592796,
  5.195327, 6.331345, 6.641488, 7.809633, 9.533514, 9.836067, 9.924506, 
    8.603547, 8.11933, 8.395448, 7.311809, 5.270021, 5.671714, 7.478117, 
    6.129735,
  6.311141, 6.944431, 5.892725, 7.344551, 8.087946, 6.213342, 4.960057, 
    5.310446, 5.996823, 5.383107, 5.033202, 6.466913, 7.701811, 7.604761, 
    5.347944,
  7.028694, 10.64195, 10.9291, 13.6614, 12.8978, 10.70429, 12.70907, 
    12.19083, 10.7371, 7.842993, 6.593657, 5.661095, 5.091051, 5.297849, 
    5.72447,
  8.438213, 9.715081, 11.39983, 12.54454, 9.745272, 9.310986, 11.43436, 
    11.52899, 11.41173, 9.789445, 8.594566, 7.940831, 6.157727, 4.074429, 
    4.760899,
  9.922235, 10.57897, 10.56689, 10.66299, 9.072794, 7.591312, 8.048326, 
    8.605666, 9.230232, 9.94186, 9.779834, 8.507111, 6.609456, 4.493724, 
    4.9933,
  10.27023, 12.52916, 13.92043, 13.91512, 11.66969, 8.380016, 6.751686, 
    7.427485, 8.613161, 7.274038, 7.999055, 7.497152, 6.626199, 4.741838, 
    5.314224,
  8.085166, 9.484995, 11.09851, 11.95785, 11.88345, 10.24445, 6.833245, 
    5.152062, 5.458782, 5.811602, 7.727582, 7.004285, 6.429543, 5.479308, 
    5.140218,
  6.490534, 7.455637, 8.094666, 8.434374, 8.293175, 8.207557, 6.920693, 
    5.35784, 5.165458, 5.099389, 5.2632, 6.002999, 5.170694, 5.234885, 
    3.917954,
  5.395487, 5.991727, 6.291533, 6.897727, 6.625959, 5.662983, 5.361573, 
    5.884772, 5.825631, 6.869003, 6.617472, 5.23145, 3.809045, 4.177136, 
    4.775024,
  4.411446, 4.622979, 5.089219, 6.005301, 6.175967, 5.611557, 4.310242, 
    3.889102, 4.910666, 6.230625, 6.164032, 4.668979, 3.36277, 4.515412, 
    7.741251,
  3.661052, 3.461867, 4.132383, 5.367166, 6.022191, 6.083495, 5.300116, 
    4.208152, 3.47782, 4.474551, 5.445365, 4.920897, 4.594382, 6.796452, 
    7.656184,
  2.901376, 3.045726, 3.959919, 5.247986, 6.168332, 6.725642, 6.698537, 
    6.159797, 5.082872, 4.436319, 4.938486, 5.820471, 6.154412, 6.999577, 
    6.457168,
  7.213525, 8.368214, 6.207285, 6.471536, 5.5265, 4.581683, 6.073585, 
    7.916316, 8.55278, 8.180918, 9.709243, 11.18131, 11.15084, 10.22952, 
    9.208579,
  7.307653, 6.52938, 5.935091, 5.336448, 4.287819, 4.468304, 6.595137, 
    9.020411, 9.658677, 8.901062, 10.11771, 13.23498, 13.93829, 9.81917, 
    8.734571,
  4.684958, 4.507169, 4.727111, 4.960705, 4.333033, 4.535334, 7.3329, 
    7.996437, 7.485653, 8.423338, 11.0934, 13.37947, 12.56797, 11.07544, 
    7.594855,
  2.932611, 3.030916, 3.380894, 4.791726, 4.949446, 4.889506, 5.850035, 
    6.493715, 7.623352, 9.80025, 11.23213, 11.24865, 9.681664, 7.990447, 
    5.289001,
  2.690071, 2.496079, 3.280641, 4.539895, 5.309381, 5.712247, 5.144096, 
    4.00531, 5.819771, 8.496035, 11.65303, 10.00358, 7.316319, 6.457363, 
    6.53884,
  3.156308, 2.413141, 2.971916, 4.058523, 5.391058, 5.619038, 4.602715, 
    4.415654, 5.303369, 6.669967, 6.907678, 8.885803, 9.823861, 9.852771, 
    9.708825,
  2.921088, 1.852051, 2.363204, 4.268739, 5.102563, 4.28224, 3.598276, 
    4.626799, 6.172086, 7.391205, 6.815008, 7.633138, 9.537362, 10.88069, 
    11.48498,
  1.54109, 1.457306, 2.604942, 4.058218, 4.219053, 3.476736, 2.761937, 
    3.501129, 5.00721, 5.951344, 5.783169, 6.582488, 8.441476, 9.743121, 
    10.08804,
  1.882925, 1.757863, 2.513991, 3.426818, 3.472221, 3.193777, 2.985902, 
    3.457291, 4.342843, 5.15292, 5.270474, 5.882341, 7.142393, 7.977903, 
    8.18788,
  3.150651, 2.271961, 2.949041, 3.585849, 3.778373, 3.69475, 3.436255, 
    3.128183, 3.178876, 3.022184, 3.502244, 5.391356, 6.07242, 7.026118, 
    7.804147,
  4.849519, 6.697682, 6.247329, 7.844195, 6.757779, 7.331517, 9.636107, 
    9.473237, 7.62007, 5.230213, 4.574164, 4.151122, 4.067165, 4.657979, 
    5.489256,
  12.03947, 7.935115, 9.070918, 8.839728, 6.868136, 6.909606, 8.512488, 
    8.693694, 7.63705, 6.16502, 5.101448, 5.163026, 4.885547, 4.304946, 
    5.594584,
  14.53053, 12.98183, 10.20273, 9.444815, 7.832664, 7.142177, 7.293772, 
    7.86096, 7.616495, 6.173853, 5.316803, 4.740098, 4.764718, 5.787791, 
    5.796064,
  12.29752, 13.03901, 12.15689, 10.06677, 8.650727, 7.275253, 6.502321, 
    6.204388, 5.800838, 4.506689, 4.690324, 4.136286, 5.081362, 6.041972, 
    4.721054,
  9.298114, 10.3285, 10.64142, 9.63623, 7.985795, 6.528892, 6.297173, 
    4.724793, 3.268876, 3.17347, 3.890576, 3.406426, 4.683069, 5.669099, 
    5.173812,
  6.72336, 7.784155, 7.937356, 7.329429, 6.82881, 6.000018, 4.71829, 
    4.506767, 3.74256, 3.263551, 2.363359, 2.445959, 3.971004, 4.437923, 
    4.595152,
  5.255044, 6.349622, 5.882463, 5.37505, 5.283039, 5.14339, 4.823349, 
    4.542672, 4.195524, 3.793675, 2.53326, 1.956472, 2.882977, 3.28725, 
    3.975866,
  4.721154, 4.806427, 3.912508, 3.955722, 3.989755, 4.011432, 3.786649, 
    3.39777, 3.173409, 3.367092, 2.346022, 2.070395, 2.601384, 2.541119, 
    3.085972,
  4.264127, 3.196545, 2.383366, 2.449608, 2.538494, 2.868284, 2.68791, 
    2.142464, 2.258997, 2.740186, 2.425166, 2.078836, 2.275029, 2.387333, 
    2.83533,
  2.689933, 1.713213, 1.657744, 1.532416, 1.649835, 1.847466, 1.9799, 
    1.759528, 1.355135, 1.077939, 1.166522, 1.705947, 2.335178, 3.272196, 
    4.617418,
  5.446392, 5.238118, 4.416406, 3.869411, 2.867603, 2.750278, 4.995563, 
    7.253987, 7.080687, 5.707461, 6.019893, 6.922927, 6.521385, 4.517231, 
    2.42585,
  8.829627, 6.592779, 5.556293, 4.693962, 2.401077, 1.823459, 3.460289, 
    5.753863, 6.991104, 6.460632, 6.761354, 8.549068, 8.443936, 4.585291, 
    2.597812,
  9.535536, 8.930303, 5.797768, 4.726174, 3.317416, 2.805788, 1.857745, 
    3.369798, 6.886041, 8.264245, 8.651887, 9.490877, 8.820193, 5.758525, 
    3.37664,
  9.73194, 10.08341, 8.793593, 4.719197, 4.636816, 4.817885, 3.926577, 
    3.613769, 3.868354, 6.807208, 8.917513, 9.317327, 8.037491, 5.502522, 
    3.351651,
  9.491121, 10.43446, 10.52185, 8.492375, 4.807645, 5.720863, 7.133018, 
    6.056583, 4.13975, 4.658035, 8.554315, 9.571018, 8.278092, 5.993183, 
    3.86116,
  8.807062, 9.713847, 10.75879, 10.16564, 7.986231, 4.80788, 6.920769, 
    9.270761, 7.414253, 7.182706, 7.321981, 9.657363, 8.283387, 6.187466, 
    4.500975,
  7.775854, 8.743905, 9.739348, 10.18149, 9.5331, 7.578257, 5.524167, 
    7.100517, 9.44803, 10.21691, 10.17731, 9.770988, 8.110232, 6.351974, 
    5.027245,
  6.24199, 7.432822, 8.577971, 9.462882, 9.655067, 8.552699, 7.395772, 
    9.170116, 10.94244, 10.94289, 10.52888, 9.482881, 7.523209, 6.123614, 
    4.842787,
  4.160594, 5.611945, 6.947287, 8.292248, 9.189067, 9.034992, 8.640772, 
    9.760755, 10.94089, 10.72233, 9.881694, 8.29712, 6.532421, 5.407978, 
    4.359436,
  1.912566, 3.561745, 5.399423, 6.883632, 8.22743, 8.955896, 9.462241, 
    9.786531, 8.645732, 6.79964, 6.434638, 6.793284, 5.560605, 4.897193, 
    4.556606,
  6.894981, 8.477451, 7.408788, 7.191946, 5.275501, 2.574337, 4.469018, 
    5.878564, 5.647833, 4.325972, 4.390372, 4.272595, 4.502282, 4.380605, 
    4.487089,
  8.951414, 9.161383, 9.77741, 8.445866, 5.092245, 3.742932, 3.769081, 
    3.734448, 4.863478, 4.206432, 4.356809, 5.540048, 6.025453, 4.739902, 
    4.915941,
  8.198508, 8.672601, 9.080655, 8.928103, 6.283056, 3.591544, 3.952872, 
    2.739358, 3.864243, 4.376059, 4.41196, 5.341108, 6.678141, 6.772247, 
    6.353806,
  7.292546, 7.775356, 8.177082, 8.49297, 7.509329, 4.384715, 2.931775, 
    4.090069, 4.119691, 2.66319, 3.831117, 4.485607, 5.563385, 6.456314, 
    6.880931,
  5.668055, 6.55447, 7.273026, 7.498227, 6.913019, 5.644059, 3.719604, 
    2.202728, 2.70635, 2.020335, 3.007312, 3.784902, 5.012343, 6.931277, 
    8.580631,
  4.166437, 5.169961, 6.304863, 6.972683, 6.809396, 5.933918, 5.161427, 
    5.305657, 3.904666, 2.427546, 2.062012, 2.934891, 4.165476, 6.710786, 
    8.372405,
  4.273325, 4.379354, 5.402464, 6.57966, 7.024457, 6.448889, 6.382019, 
    6.453076, 5.943045, 5.575696, 4.61981, 3.646059, 4.691202, 6.697053, 
    8.548772,
  4.769485, 4.067357, 5.178155, 6.496868, 6.996431, 6.849244, 6.663252, 
    7.170614, 7.788753, 7.571014, 6.569674, 6.292196, 6.946683, 7.959548, 
    9.354668,
  3.942078, 3.425509, 4.633104, 5.811302, 6.56644, 6.897014, 7.2482, 
    6.673256, 6.983768, 7.253531, 8.14058, 8.952731, 9.252007, 9.921359, 
    9.98681,
  3.08034, 2.620667, 4.021649, 5.393831, 6.443192, 7.305288, 8.045398, 
    7.11769, 5.854347, 5.303143, 6.875795, 10.10259, 10.491, 11.10038, 
    10.08122,
  13.13416, 13.22418, 8.946644, 8.746314, 7.269735, 6.040694, 7.814629, 
    8.381728, 7.554328, 5.681574, 5.028837, 4.255634, 4.155594, 3.3015, 
    3.68283,
  17.06646, 16.42697, 13.03458, 9.449042, 6.431849, 5.799402, 7.160745, 
    7.291222, 6.429863, 4.964789, 4.733939, 5.222225, 5.205321, 3.457781, 
    3.556006,
  15.16313, 16.4949, 15.82368, 12.00936, 7.808858, 5.422373, 5.7002, 
    7.435496, 8.045794, 6.637553, 5.095074, 4.613773, 5.013182, 4.290956, 
    4.055051,
  12.62999, 14.17358, 15.19056, 14.49618, 10.79091, 6.275465, 5.194381, 
    7.217674, 9.435438, 7.306308, 6.129875, 4.278567, 3.264741, 3.17085, 
    4.112574,
  9.07763, 10.81748, 12.49263, 13.32673, 12.32681, 9.335169, 6.825334, 
    5.803777, 3.969116, 3.984956, 5.954625, 5.091694, 3.623789, 3.022007, 
    4.492898,
  5.695218, 6.761245, 8.778517, 10.42833, 11.20617, 10.84186, 9.18921, 
    7.177787, 4.582901, 3.814633, 3.96455, 5.47993, 4.307748, 3.224613, 
    3.437693,
  4.233797, 3.418757, 4.253102, 6.537618, 8.188684, 9.083473, 9.186789, 
    8.605873, 7.502001, 6.084728, 5.307794, 4.825275, 4.152715, 3.609135, 
    3.285234,
  4.88066, 2.951183, 2.628366, 3.154004, 4.689366, 5.853837, 6.445164, 
    6.653204, 6.393076, 5.941787, 5.628731, 5.035728, 4.167665, 3.665191, 
    3.608237,
  5.391673, 3.975232, 3.108789, 2.872565, 2.53288, 3.500651, 4.462963, 
    5.415377, 5.759231, 5.317258, 4.875828, 4.777114, 4.748961, 4.404317, 
    3.842753,
  4.690629, 4.181886, 4.049606, 4.03226, 3.596185, 2.926877, 3.215047, 
    3.884419, 3.974143, 3.313015, 3.89499, 5.284369, 5.465339, 5.464512, 
    5.110958,
  8.82373, 4.502766, 6.782233, 7.112494, 4.024956, 3.360124, 6.900246, 
    8.948024, 8.700441, 7.721816, 7.282036, 6.5457, 6.164057, 4.63747, 
    3.912602,
  15.23502, 5.500703, 6.366843, 6.857337, 3.796307, 2.920209, 6.036795, 
    8.295141, 8.429219, 7.26784, 7.253067, 7.649803, 7.455578, 4.67877, 
    3.934631,
  17.06556, 10.31511, 4.947399, 4.952072, 3.62499, 3.715375, 3.805992, 
    6.266484, 8.585501, 8.499972, 8.299003, 8.466105, 7.914664, 6.51083, 
    4.687759,
  16.74542, 14.73749, 7.795951, 3.981294, 3.782686, 4.936934, 5.463252, 
    5.080249, 4.954477, 5.776124, 7.665699, 7.893254, 7.179914, 5.941054, 
    4.688737,
  15.22263, 15.94014, 13.20772, 7.4376, 3.575706, 5.870448, 8.185777, 
    7.784316, 3.846896, 2.754889, 6.243372, 7.437523, 6.921732, 6.024578, 
    5.585401,
  12.38815, 14.60624, 15.24258, 12.35792, 6.899786, 4.784735, 7.511741, 
    8.843608, 6.395909, 4.797386, 5.127626, 7.436916, 7.252568, 6.175236, 
    4.974196,
  10.33969, 12.0183, 13.62376, 14.20562, 11.84437, 6.987851, 5.783485, 
    6.272863, 6.939361, 7.615171, 7.968435, 8.116656, 7.739203, 6.944548, 
    5.695306,
  8.484245, 9.190569, 10.72125, 12.69333, 13.43422, 10.8542, 7.366512, 
    7.937701, 8.285395, 8.400275, 8.533827, 8.449413, 8.012759, 7.424284, 
    6.345759,
  6.744414, 6.040021, 6.832954, 9.098031, 11.69339, 12.2778, 10.0245, 
    8.269794, 8.296827, 8.26159, 8.525517, 8.526464, 8.006399, 7.475688, 
    6.250872,
  5.048091, 3.947186, 3.939659, 5.257596, 8.014087, 10.16755, 10.64253, 
    9.12299, 6.915665, 5.478219, 6.151503, 7.790438, 7.134297, 6.560935, 
    5.363628,
  9.155606, 7.062159, 5.457249, 7.744963, 5.40996, 2.902866, 1.851812, 
    5.693299, 3.32926, 5.293374, 7.38138, 7.128666, 6.889565, 5.653759, 
    5.612637,
  13.03429, 7.447168, 3.962338, 7.71385, 5.565305, 3.138498, 2.749649, 
    4.599032, 4.087406, 3.999299, 7.799711, 8.344926, 7.814964, 5.378044, 
    4.849393,
  13.07407, 9.109155, 2.23417, 6.885345, 5.854567, 3.074416, 2.148866, 
    3.134564, 3.072026, 6.52974, 9.236265, 9.166161, 8.133965, 6.434314, 
    4.341554,
  13.07491, 10.90151, 3.298849, 5.430676, 6.086651, 4.751099, 2.359554, 
    1.86496, 3.972288, 5.366837, 8.86335, 8.893727, 7.961802, 6.30617, 
    4.412956,
  12.67781, 12.26396, 7.638721, 2.591517, 5.584771, 5.358903, 4.740006, 
    3.669361, 2.703204, 2.950822, 7.690864, 8.546163, 7.9704, 6.484456, 
    4.951147,
  10.64942, 12.47238, 10.56213, 4.754796, 3.966083, 5.873827, 6.291904, 
    6.330359, 3.907019, 3.620124, 5.26643, 8.39141, 8.022913, 6.668335, 
    5.052404,
  9.561071, 11.68722, 11.50898, 9.213329, 3.578922, 5.842888, 6.918415, 
    5.754853, 4.870613, 5.390426, 7.137321, 8.603675, 8.377584, 7.2376, 
    5.702349,
  8.024294, 10.24938, 11.02248, 11.18165, 8.934473, 3.878348, 7.542635, 
    8.161186, 7.438506, 6.466627, 6.645336, 8.093866, 8.356019, 7.591771, 
    6.252765,
  5.91396, 7.799906, 9.296934, 11.01853, 11.6371, 7.518558, 5.612966, 
    8.278048, 7.853463, 6.636777, 6.402252, 7.395855, 7.998558, 7.718518, 
    6.586434,
  3.881672, 5.077774, 6.857814, 9.522912, 12.1377, 12.05439, 6.258943, 
    7.195383, 7.176999, 5.268175, 5.142565, 7.10473, 7.443623, 7.689149, 
    6.916959,
  5.164035, 7.932854, 7.006207, 8.409231, 7.152252, 5.168714, 5.020635, 
    5.35068, 6.304421, 4.922925, 4.765639, 4.675841, 4.71022, 4.507028, 
    4.885571,
  7.776678, 8.927336, 8.155127, 7.927776, 5.564947, 4.229182, 4.897328, 
    5.435915, 6.352144, 4.989834, 5.147924, 5.281723, 5.367083, 4.179287, 
    4.340236,
  8.571608, 9.326718, 7.55374, 6.754242, 5.206567, 3.384226, 3.497126, 
    5.409825, 5.170029, 5.708859, 5.629691, 5.936276, 5.705239, 4.802189, 
    3.657056,
  8.823874, 9.159299, 6.795011, 5.529991, 5.270615, 4.367245, 2.356508, 
    2.350541, 3.333331, 5.068872, 6.133062, 6.08517, 5.315892, 4.894925, 
    3.829165,
  8.437321, 9.221612, 6.923173, 4.229639, 4.059733, 3.644211, 2.933925, 
    2.674262, 2.552289, 2.792619, 6.577591, 6.069457, 5.118259, 5.074435, 
    5.048997,
  7.080398, 9.091602, 7.683642, 3.61771, 3.455913, 3.167454, 3.29459, 
    4.122608, 3.784014, 4.34095, 5.018593, 6.277502, 5.246156, 4.99191, 
    5.416875,
  5.808038, 8.713177, 8.437987, 4.253547, 2.306669, 2.497292, 2.786858, 
    4.236498, 4.92165, 7.300268, 7.761946, 7.090953, 5.784944, 5.254837, 
    5.260636,
  4.88026, 7.984374, 9.057528, 6.440904, 2.577509, 2.415875, 2.920164, 
    3.402395, 5.11643, 7.312286, 7.804193, 7.256716, 6.224021, 5.397762, 
    4.714524,
  3.89826, 6.296294, 8.597513, 8.642954, 5.016088, 2.770928, 2.33588, 
    3.408221, 4.326931, 6.477668, 7.031742, 6.982741, 6.405489, 5.611956, 
    4.480409,
  3.120549, 4.259376, 6.966366, 9.706118, 9.299993, 5.747087, 2.859148, 
    3.084452, 4.410027, 4.308087, 4.893874, 6.457248, 6.123126, 5.773396, 
    4.826194,
  2.208369, 2.613814, 2.531166, 4.468501, 4.687168, 3.841121, 4.91228, 
    5.891494, 5.7616, 5.317498, 6.396518, 4.635158, 2.873797, 4.465592, 
    4.835207,
  3.746592, 3.840329, 3.223744, 4.283708, 3.905568, 3.565547, 4.974542, 
    5.810862, 6.101556, 5.582231, 6.118119, 4.286261, 3.770484, 4.392477, 
    5.000389,
  3.966678, 4.02202, 3.943467, 4.148715, 3.560373, 3.311895, 4.269326, 
    4.49086, 4.682515, 5.364942, 5.755418, 2.915123, 4.348617, 5.820222, 
    5.246014,
  3.812805, 4.048143, 4.121704, 4.560594, 4.725406, 4.577282, 3.679518, 
    4.197295, 4.546856, 4.970923, 4.395502, 2.046375, 4.533478, 6.275774, 
    5.53631,
  4.013972, 3.946543, 4.581974, 5.698781, 6.118657, 6.278297, 5.629612, 
    3.14497, 3.163141, 3.515553, 3.876245, 2.137939, 4.31838, 6.830602, 
    6.860566,
  4.001795, 4.091582, 5.840725, 6.979544, 7.348427, 7.345922, 7.053062, 
    6.793381, 4.295692, 3.021831, 2.906549, 2.07416, 3.906929, 6.809902, 
    6.972611,
  4.537658, 5.682896, 7.09245, 7.692375, 7.907038, 7.528639, 7.368187, 
    6.341737, 5.178372, 4.03298, 3.751572, 2.150457, 4.360098, 6.866338, 
    7.226377,
  6.041417, 6.974679, 7.594732, 7.581002, 7.406912, 7.457977, 7.441743, 
    7.487858, 6.753515, 4.76974, 3.651074, 2.538024, 4.978662, 7.195449, 
    7.078366,
  7.029872, 6.689198, 6.543024, 7.349446, 6.455606, 7.249287, 7.837016, 
    7.502401, 6.709147, 5.019769, 4.214327, 3.253537, 5.622864, 7.59697, 
    6.878005,
  7.22835, 5.732898, 5.366126, 7.89891, 7.251448, 6.150222, 7.93618, 
    8.183071, 6.432843, 3.863955, 3.405776, 3.814185, 5.949995, 7.700608, 
    6.633212,
  3.734597, 4.571475, 4.052641, 5.193661, 5.197143, 5.556209, 7.808095, 
    8.620811, 8.43556, 6.726915, 6.296112, 5.254887, 4.780618, 5.002146, 
    5.651872,
  4.773776, 4.326461, 2.80522, 3.256109, 3.237171, 3.805671, 6.005261, 
    7.783999, 8.994744, 8.812435, 7.419776, 5.718769, 5.408138, 4.003829, 
    4.605845,
  4.735138, 5.110541, 3.013344, 1.461923, 2.162066, 2.409953, 4.075742, 
    4.804381, 6.760654, 9.581813, 10.13194, 6.908973, 5.488644, 4.635751, 
    3.546661,
  3.161077, 4.528432, 4.38562, 2.988048, 1.416, 1.669374, 2.087781, 3.86212, 
    5.859931, 8.663264, 10.37311, 7.881028, 5.01109, 4.720503, 3.563085,
  1.534946, 2.26097, 4.231514, 4.618116, 3.898331, 2.89699, 2.562579, 
    1.816852, 3.071601, 5.058673, 8.538294, 8.901331, 5.068403, 4.608878, 
    4.495711,
  2.704643, 3.461367, 4.519759, 5.448011, 5.959195, 6.087643, 5.295117, 
    4.124422, 2.869802, 2.790856, 4.802467, 8.296811, 5.190074, 4.481622, 
    4.464855,
  5.111732, 5.028253, 5.612343, 6.238102, 7.012059, 7.582553, 7.46891, 
    6.496912, 4.838844, 3.617757, 4.266809, 6.367482, 5.143775, 4.17275, 
    4.392303,
  5.141289, 5.237875, 6.022956, 6.950103, 7.65423, 8.150665, 8.349325, 
    8.408996, 7.504627, 5.810707, 4.23905, 4.395581, 4.349041, 3.846516, 
    4.210544,
  5.45635, 6.064852, 6.604811, 7.450222, 7.991413, 8.314653, 8.670855, 
    8.763239, 8.277762, 7.202728, 5.659241, 3.967233, 3.373574, 3.738333, 
    4.005767,
  6.41678, 7.372137, 7.649807, 7.935794, 7.995557, 8.299212, 8.868142, 
    9.012712, 7.858825, 5.936742, 5.02608, 4.676367, 3.10219, 3.878608, 
    3.998158 ;

 sftlf =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.141347, 0.07456003, 0.2762221, 0, 0.2154952, 0.5089986, 0.007178012, 0, 
    0.1467785, 25.31165, 20.60715, 2.120196, 15.979, 48.81725, 63.64272,
  0.001503375, 0, 0, 0, 0.8848332, 11.68672, 0, 0, 0, 0.4694104, 0.9680001, 
    0.09868675, 1.334438, 150.908, 101.0153,
  0, 0, 0, 0, 8.803595, 280.9762, 7.478715, 0, 0, 0, 0.0046135, 0, 
    0.00845787, 0.9458157, 6.678408,
  0, 0, 0, 0, 0, 12.95772, 307.1121, 15.76765, 0, 0, 0, 0, 0.001950179, 
    0.08926713, 2.882818,
  0, 0, 0, 0, 0, 0, 9.245329, 485.3841, 540.1508, 15.00115, 0.01623012, 0, 0, 
    0.06344586, 0.01027276,
  0, 0, 0, 0, 0, 0, 0, 1.278773, 12.13823, 0.8518202, 0.2699268, 0, 0, 
    0.01012854, 0.01599434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05785002, 0, 0, 0, 0, 0.2725836,
  0, 0, 0, 0, 0, 0, 0, 0.3482242, 1.154397, 3.605569, 0.8750445, 0, 0.158783, 
    0.02233585, 0.6264485 ;
}
