netcdf \20030101.atmos_static_cmip.tile1 {
dimensions:
	grid_xt = 96 ;
	grid_yt = 96 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:associated_files = "area: 20030101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 time = 0 ;

 orog =
  8.54475, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  110.6839, 9.015973, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  118.8102, 18.13202, 0.007421071, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  130.705, 39.06387, 3.106806, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  141.0809, 84.24564, 11.19796, 0.4508977, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.9822, 184.6116, 106.8482, 7.492514, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.08320683, 3.271346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  180.4211, 249.8835, 220.8967, 76.21671, 1.021369, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21.94272, 34.81591, 74.42256, 66.43814, 11.87937, 0, 0, 0, 0, 0, 0, 0, 0,
  149.0657, 196.1795, 177.1756, 126.4176, 11.39334, 0.5445582, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.201014, 10.06274, 
    26.85098, 48.46229, 196.196, 446.1897, 398.605, 448.8601, 587.3398, 
    619.0617, 478.8845, 191.0291, 9.431361, 0, 0, 0, 0, 0, 0,
  247.4764, 260.0786, 196.9956, 132.1378, 48.361, 5.852092, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.821061, 227.5061, 
    341.0564, 416.8428, 546.1491, 760.7002, 800.6117, 811.9203, 918.2296, 
    1199.078, 1194.457, 1065.196, 779.4019, 539.7784, 68.59048, 0, 0, 0, 0, 0,
  254.4188, 378.3603, 367.6226, 301.4343, 162.2049, 108.9995, 0.9085217, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.392265, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    84.11958, 610.6379, 784.4166, 873.3272, 803.2366, 954.6566, 1133.667, 
    1193.683, 1333.627, 1518.089, 1657.062, 1719.367, 1548.189, 1097.09, 
    488.3766, 19.6729, 0, 0, 0, 0,
  282.803, 388.1694, 501.5489, 557.1978, 613.9719, 624.3671, 154.6011, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.850073, 136.7001, 
    621.1481, 1059.969, 1205.403, 1271.604, 1289.321, 1373.992, 1468.906, 
    1399.973, 1501.777, 1674.687, 2147.529, 2156.621, 1497.179, 907.9773, 
    341.0655, 33.16307, 0, 0, 0,
  281.039, 423.6907, 485.7559, 651.8676, 783.3052, 889.3768, 610.0162, 
    16.97377, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    129.3114, 660.4066, 997.0892, 1271.035, 1259.05, 1269.307, 1282.922, 
    1357.486, 1418.984, 1464.053, 1694.626, 2161.078, 2172.453, 1467.212, 
    1030.81, 612.332, 164.4304, 1.996331, 0, 0,
  322.6488, 427.8226, 549.0103, 681.7765, 829.639, 1022.879, 837.8648, 
    305.3638, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.138049, 280.6169, 659.5826, 1002.684, 1031.975, 1099.151, 1099.102, 
    1133.435, 1221.698, 1317.967, 1415.099, 1513.935, 1787.441, 1850.336, 
    1464.755, 1240.903, 696.9532, 172.8423, 13.54243, 0, 0,
  246.0376, 453.1236, 631.008, 871.3788, 1047.864, 932.1511, 816.0308, 
    317.9274, 6.631444, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    150.0291, 674.2753, 908.9203, 930.3144, 938.6702, 1006.137, 1124.25, 
    1170.841, 1154.932, 1264.449, 1330.767, 1451.47, 1585.219, 1689.979, 
    1656.847, 1377.684, 685.7067, 148.093, 7.893209, 0, 0,
  302.9081, 427.2077, 600.2842, 822.6921, 987.5324, 917.3104, 668.1157, 
    303.2888, 0.4759156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05529097, 404.3319, 849.9101, 942.0059, 899.2049, 892.3331, 1045.702, 
    1259.788, 1338.622, 1238.361, 1260.895, 1324.21, 1411.141, 1544.977, 
    1598.17, 1706.571, 1414.926, 652.4966, 175.4458, 20.1155, 25.00171, 
    36.41872,
  304.3976, 367.4553, 507.5162, 723.1177, 889.1189, 890.2856, 860.1849, 
    487.2796, 0.9306844, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    48.47385, 456.4773, 788.9446, 784.0788, 797.9801, 888.491, 1040.636, 
    1257.102, 1379.351, 1308.995, 1358.369, 1450.252, 1468.341, 1489.487, 
    1519.486, 1585.82, 1321.473, 545.1862, 138.8361, 40.63335, 49.9632, 
    84.77402,
  357.9227, 326.5664, 409.4615, 533.1976, 722.5844, 805.3265, 892.149, 
    651.6109, 85.95663, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.497938, 272.2702, 615.2929, 908.9059, 917.061, 841.0509, 900.0991, 
    989.4551, 1097.285, 1229.295, 1245.714, 1381.851, 1374.066, 1291.548, 
    1248.401, 1166.31, 1273.148, 967.5308, 443.7959, 159.7697, 64.36124, 
    74.43269, 110.2169,
  374.3119, 313.8954, 345.6318, 445.4458, 583.0211, 721.8264, 795.6353, 
    683.6541, 309.0318, 22.92986, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 217.3822, 804.5779, 921.5053, 1073.372, 1032.455, 914.3887, 915.9861, 
    975.9174, 1025.77, 1091.464, 1183.756, 1203.829, 1146.519, 1118.986, 
    1206.85, 1186.365, 1061.127, 699.5498, 315.4096, 174.5182, 91.69196, 
    117.5326, 129.1317,
  384.2018, 316.835, 329.2943, 348.3972, 449.1535, 490.7008, 580.1392, 
    682.83, 561.0168, 450.0525, 74.4604, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.625334, 529.3156, 1179.003, 1083.251, 1046.369, 1010.433, 952.2749, 
    974.9957, 1008.044, 1025.375, 1088.216, 1136.371, 1137.306, 977.9841, 
    966.8591, 1095.862, 1080.748, 967.8829, 583.6017, 349.6461, 208.4064, 
    122.2884, 137.5921, 124.6154,
  425.9325, 402.693, 356.9512, 342.1429, 387.3358, 451.6554, 543.8193, 
    598.1646, 671.4254, 663.9327, 658.8842, 342.5872, 1.323529, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 55.75727, 723.3252, 1345.097, 1208.163, 1096.152, 
    1057.105, 1042.026, 1052.195, 1075.99, 1085.4, 1083.792, 1107.45, 
    1089.932, 1003.74, 908.7562, 881.2886, 806.4973, 725.7192, 521.3715, 
    374.6654, 268.3831, 172.0694, 131.0901, 57.53464,
  461.6035, 467.3536, 394.1595, 343.5833, 356.553, 412.9582, 456.8489, 
    546.8406, 586.7995, 714.7881, 969.0544, 855.0431, 500.8872, 32.52318, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 123.6441, 855.6476, 1413.006, 1269.892, 
    1172.559, 1156.56, 1149.75, 1151.305, 1144.381, 1103.469, 1061.514, 
    1045.96, 1102.312, 1112.108, 971.346, 808.2177, 695.4062, 630.5798, 
    525.356, 437.357, 384.1834, 350.2086, 123.1665, 31.22814,
  464.4684, 508.0797, 455.048, 373.7856, 366.4037, 387.9864, 443.3236, 
    495.3125, 589.3275, 739.6755, 988.6879, 1060.314, 904.9486, 528.0706, 
    225.8937, 27.69355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 174.664, 879.7312, 1444.223, 
    1357.686, 1256.545, 1275.17, 1242.061, 1206.494, 1137.42, 1064.367, 
    1009.382, 1009.102, 1074.426, 1101.382, 1013.848, 935.0889, 872.3643, 
    823.5287, 742.5305, 702.767, 638.2717, 610.8529, 236.0903, 19.05215,
  377.5986, 476.2537, 554.4959, 498.4242, 421.1341, 410.7194, 460.7333, 
    508.1182, 604.0519, 780.8995, 940.6996, 912.0196, 1031.078, 860.0245, 
    593.0319, 288.8579, 12.86605, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 211.1246, 927.424, 
    1489.004, 1561.025, 1444.746, 1376.06, 1280.973, 1179.52, 1098.244, 
    1019.69, 975.9384, 963.2079, 978.0944, 1029.098, 1103.491, 1163.96, 
    1175.215, 1136.579, 1103.248, 1014.715, 943.465, 803.7495, 369.8148, 
    113.7734,
  332.751, 472.4073, 685.3926, 635.038, 517.4619, 464.7151, 489.6293, 
    589.0376, 704.1102, 888.3381, 946.3566, 843.2612, 937.7106, 952.2573, 
    593.1406, 408.6372, 87.12373, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 274.805, 948.42, 
    1506.014, 1601.052, 1578.846, 1456.921, 1284.965, 1163.84, 1079.576, 
    1015.096, 961.92, 924.3301, 919.1673, 969.1686, 1080.93, 1206.276, 
    1290.624, 1303.251, 1316.85, 1354.376, 1136.7, 970.1143, 487.621, 182.6047,
  386.6328, 599.5612, 743.3576, 737.4709, 670.9242, 536.273, 553.6517, 
    674.8468, 801.8613, 965.2466, 953.0202, 781.4857, 825.5333, 884.1866, 
    743.7918, 650.3617, 509.5243, 47.25615, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34.19665, 536.6432, 
    1112.04, 1443.481, 1515.864, 1440.972, 1356.049, 1192.005, 1062.608, 
    976.4597, 953.9917, 942.6937, 942.3792, 969.4203, 966.9082, 1031.604, 
    1100.836, 1155.753, 1179.703, 1365.894, 1379.681, 1287.486, 922.5301, 
    544.6479, 214.8122,
  407.2789, 556.476, 691.2809, 737.9501, 749.3389, 662.7368, 563.8776, 
    667.7236, 775.2804, 860.3702, 857.4185, 735.3098, 719.4968, 858.9086, 
    655.9019, 560.5863, 441.2978, 138.1514, 0.004807308, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 245.0765, 
    740.5414, 1216.22, 1399.232, 1428.595, 1324.44, 1244.887, 1171.623, 
    1058.757, 978.5461, 948.2759, 945.5349, 979.3757, 1012.527, 980.8537, 
    912.5103, 983.9648, 1005.987, 1126.251, 1280.425, 1263.255, 944.915, 
    620.7706, 330.2798, 198.4007,
  485.9347, 536.7831, 520.842, 574.1156, 628.2961, 593.3192, 671.6805, 
    760.3802, 792.5333, 809.5409, 713.7068, 694.2451, 762.8157, 893.8396, 
    750.4239, 489.7271, 319.0528, 122.3887, 1.660121, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1749505, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36.20846, 
    639.6878, 1064.495, 1200.584, 1345.762, 1339.131, 1276.558, 1206.219, 
    1145.992, 1077.639, 997.5162, 966.3801, 956.3568, 970.2714, 1008.335, 
    951.059, 828.9758, 706.606, 863.0428, 1080.806, 1123.896, 920.291, 
    656.9827, 373.7796, 334.5416, 526.0103,
  571.2805, 576.3853, 467.4599, 411.0854, 392.3285, 505.7308, 722.9926, 
    869.4109, 931.8525, 811.3553, 662.9765, 604.0966, 688.219, 858.3245, 
    825.9299, 572.1747, 408.3769, 146.4941, 9.387668, 0.001074584, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    273.4626, 965.0869, 1142.758, 1166.024, 1121.857, 1187.254, 1166.343, 
    1151.341, 1121.571, 1066.005, 1020.396, 995.9119, 976.3922, 999.8099, 
    1080.855, 1153.143, 949.2833, 796.8798, 704.9807, 751.8674, 635.2756, 
    537.6038, 460.5406, 432.7109, 753.7834, 783.1511,
  541.8253, 527.6813, 442.9381, 349.75, 282.5704, 372.3629, 647.7617, 
    839.8668, 941.1125, 907.2533, 705.0693, 633.6419, 637.7145, 768.287, 
    809.7827, 674.5598, 493.8878, 279.3312, 44.60109, 0.003030813, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59.35226, 753.0102, 1128.37, 1213.516, 1102.814, 1106.985, 1138.11, 
    1148.302, 1144.664, 1119.719, 1075.693, 1028.648, 1007.681, 1040.419, 
    1070.42, 1085.326, 1113.797, 1101.634, 964.3666, 826.3594, 688.6269, 
    581.0179, 749.9571, 747.4507, 813.9899, 1027.863, 909.4127,
  451.7546, 465.3449, 395.6716, 335.8462, 247.0956, 298.3383, 466.0626, 
    661.6984, 813.6958, 827.1074, 757.3602, 671.0699, 631.3232, 636.7422, 
    748.9434, 753.5067, 653.6973, 358.9735, 111.3765, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 237.6711, 881.6313, 
    1209.199, 1111.17, 1116.662, 1148.323, 1170.288, 1177.596, 1179.032, 
    1162.061, 1096.823, 1040.075, 1027.026, 1072.69, 1144.079, 1132.332, 
    1099.773, 1094.171, 1114.551, 970.8142, 812.7686, 713.1152, 878.1364, 
    977.2021, 1026.251, 1069.996, 736.0057,
  391.2837, 370.3196, 366.6443, 340.5762, 263.041, 234.9373, 359.7917, 
    485.6016, 684.4538, 736.9855, 740.4536, 781.7585, 658.1667, 565.2335, 
    713.5017, 808.0051, 692.545, 472.7854, 120.2969, 0.03788849, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 152.0637, 
    745.3533, 1129.647, 1190.232, 1165.257, 1217.449, 1233.613, 1242.039, 
    1225.1, 1190.186, 1129.522, 1051.2, 1039.217, 1088.383, 1158.137, 
    1160.562, 1157.639, 1146.778, 1176.388, 1196.262, 1103.755, 939.6448, 
    773.607, 786.1696, 1066.588, 999.4681, 658.9298,
  343.9839, 329.1209, 326.8227, 338.2211, 268.4422, 231.5902, 273.1661, 
    411.1793, 556.3333, 647.4001, 724.2601, 776.667, 679.067, 508.2994, 
    620.4402, 716.1536, 666.8013, 484.4005, 195.8266, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49.35054, 549.8828, 
    1179.242, 1286.947, 1285.081, 1347.293, 1373.125, 1342.854, 1282.255, 
    1234.189, 1156.042, 1075.134, 1044.677, 1093.778, 1146.635, 1190.949, 
    1194.665, 1203.338, 1225.234, 1270.81, 1379.499, 1236.873, 994.0289, 
    744.1392, 1000.295, 1032.345, 591.7537,
  341.9223, 323.5297, 312.363, 327.7422, 256.121, 211.4899, 232.2774, 
    293.0904, 373.0227, 483.3326, 649.4127, 771.75, 673.2164, 571.9428, 
    626.7587, 791.145, 642.7789, 521.3182, 201.4202, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.703202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.91209, 
    566.6647, 1165.319, 1443.802, 1442.337, 1513.629, 1471.694, 1443.57, 
    1354.923, 1276.675, 1185.226, 1087.362, 1080.905, 1145.881, 1175.568, 
    1221.021, 1282.013, 1268.265, 1230.614, 1228.024, 1211.29, 1307.737, 
    1161.229, 873.0657, 933.2297, 1159.808, 670.6091,
  346.7993, 338.6057, 314.9171, 289.7007, 236.9087, 190.2888, 202.9013, 
    268.8091, 310.8858, 411.589, 656.1295, 740.801, 656.6727, 541.4875, 
    678.8455, 853.9406, 730.4851, 459.3751, 220.1203, 13.96118, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    413.7036, 981.3401, 1411.613, 1624.979, 1620.908, 1479.521, 1444.335, 
    1392.403, 1297.059, 1161.221, 1098.89, 1153.009, 1254.525, 1302.453, 
    1335.512, 1364.571, 1280.526, 1204.677, 1180.655, 1170.281, 1240.504, 
    1336.752, 1084.095, 1070.497, 1113.52, 930.3657,
  373.4141, 339.6274, 318.1039, 291.9559, 260.7186, 191.6193, 197.949, 
    276.8808, 356.4713, 444.8528, 671.9672, 707.4572, 541.8743, 515.196, 
    593.6595, 844.5728, 740.3514, 450.5794, 236.8895, 126.5775, 12.02609, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    74.79279, 582.2818, 1387.929, 1653.479, 1656.323, 1452.037, 1384.894, 
    1380.74, 1263.157, 1129.277, 1087.819, 1140.283, 1291.528, 1349.267, 
    1427.148, 1380.747, 1211.18, 1182.415, 1173.129, 1242.567, 1253.907, 
    1328.973, 1235.93, 1102.579, 1212.149, 1188.651,
  411.907, 359.5694, 312.9021, 316.0843, 319.7564, 228.2056, 193.8342, 
    296.6815, 321.6121, 390.0383, 586.1972, 616.8071, 522.6686, 497.1555, 
    514.1055, 625.6185, 709.9496, 500.6991, 322.1615, 233.313, 73.02024, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 251.8302, 1240.724, 1602.32, 1519.831, 1331.846, 1307.905, 1319.815, 
    1247.846, 1123.754, 1088.791, 1091.119, 1166.166, 1236.438, 1262.825, 
    1296.363, 1122.022, 1172.453, 1197.705, 1311.24, 1400.86, 1405.443, 
    1374.509, 1337.278, 1486.886, 1500.223,
  361.1769, 319.2283, 308.7516, 344.1496, 351.8325, 252.6501, 205.3004, 
    264.0542, 284.5062, 319.0981, 459.6907, 492.8576, 454.6547, 494.1764, 
    467.236, 499.1732, 633.0408, 550.3798, 449.2036, 364.1278, 174.6403, 
    28.89057, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 104.2696, 1010.841, 1362.054, 1315.101, 1130.426, 1149.357, 
    1245.088, 1169.575, 1095.747, 1041.157, 1027.792, 1023.939, 991.415, 
    1043.899, 1006.476, 1261.374, 1189.962, 1103.186, 1205.096, 1273.994, 
    1571.499, 1265.122, 1354.616, 1342.277, 1499.963,
  288.3837, 296.7624, 328.1481, 349.2853, 354.0044, 300.8336, 209.8271, 
    242.339, 257.6059, 315.6365, 438.6422, 454.057, 469.7331, 499.5292, 
    472.8086, 418.0537, 492.4049, 451.988, 414.6512, 387.9483, 298.7437, 
    224.9868, 30.84828, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.8451669, 71.35338, 642.9059, 1073.645, 1063.941, 
    943.9172, 1026.204, 1114.221, 1073.748, 1012.559, 1027.82, 1014.382, 
    1057.285, 1027.442, 823.2462, 941.8942, 1091.702, 1226.689, 1104.525, 
    1242.194, 1126.849, 1339.002, 1262.845, 1232.307, 1363.345, 1223.546,
  260.1389, 284.7289, 287.6657, 321.2379, 323.3841, 321.9951, 239.3829, 
    211.8097, 231.2988, 276.1485, 389.8618, 400.1599, 419.2465, 413.5182, 
    379.3967, 365.7533, 402.7262, 476.0164, 436.6118, 442.7455, 523.3729, 
    513.603, 263.7818, 2.99741, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 6.84726, 127.0682, 564.7839, 1027.651, 923.8217, 
    809.4365, 946.3239, 1098.568, 971.295, 901.8392, 924.174, 968.075, 
    986.755, 1009.199, 898.538, 673.96, 868.1624, 893.8102, 1322.028, 
    1317.703, 1118.277, 1254.662, 1102.685, 1225.965, 1365.095, 1100.581,
  256.0101, 258.5121, 265.4595, 271.6456, 281.9239, 339.2019, 239.4398, 
    201.6286, 231.9184, 272.3331, 346.6201, 365.2863, 335.9691, 301.0338, 
    258.306, 271.6318, 450.0833, 557.5646, 531.2784, 522.4316, 549.2473, 
    622.1465, 329.0093, 25.54767, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.427928, 262.789, 692.8567, 1032.231, 824.3097, 
    711.4518, 954.0336, 994.9745, 852.847, 765.702, 840.2001, 873.9611, 
    851.5475, 920.1156, 891.8646, 743.049, 630.5678, 807.291, 1051.364, 
    1174.423, 1034.36, 1105.102, 1130.744, 1221.451, 1312.698, 1236.457,
  244.8726, 235.7898, 238.6499, 250.9584, 264.177, 304.3681, 231.7038, 
    171.5492, 194.0964, 237.4297, 322.8626, 324.8877, 315.0707, 258.6005, 
    236.6363, 277.2534, 457.8071, 528.7694, 405.2236, 342.8656, 385.32, 
    442.8686, 295.1935, 24.17916, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.293201, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52.95097, 347.3517, 720.2449, 929.5432, 
    735.391, 780.5626, 910.9541, 885.9318, 687.3369, 662.2593, 723.8735, 
    755.4806, 723.0743, 769.8126, 788.1163, 702.8589, 630.3057, 768.6213, 
    1059.849, 972.3868, 1188.259, 1177.481, 1121.192, 1184.726, 1279.616, 
    1302.242,
  235.042, 217.7554, 200.0201, 218.5201, 210.6107, 214.8637, 159.0711, 
    132.8887, 194.6062, 222.7486, 255.3079, 243.1668, 189.8971, 189.5496, 
    151.8132, 254.9043, 441.0879, 450.9707, 312.1183, 209.6811, 199.2862, 
    258.3366, 160.7645, 4.592148, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1700515, 92.22056, 366.6779, 594.3502, 777.5218, 
    693.3395, 719.6742, 801.9887, 715.3484, 599.9813, 555.8511, 606.0909, 
    628.077, 622.9703, 659.368, 666.463, 613.6947, 660.4321, 819.1418, 
    1024.8, 1005.07, 1167.154, 1107.55, 1131.997, 1173.377, 1208.152, 1350.651,
  196.7365, 204.5998, 198.4898, 193.5049, 169.7109, 154.1599, 121.315, 
    140.5267, 197.9303, 241.7397, 228.9246, 149.1499, 105.5863, 101.0614, 
    123.9294, 166.2768, 433.4229, 365.3992, 271.7154, 133.414, 51.558, 
    55.21501, 35.0076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13.58836, 185.3467, 334.9186, 518.5123, 624.0504, 611.5664, 
    573.1268, 551.8474, 545.7886, 508.7069, 509.3336, 518.7409, 552.8677, 
    565.2957, 587.2665, 552.8708, 585.5536, 619.3701, 901.4293, 1212.324, 
    1221.37, 1192.156, 1120.597, 1169.473, 1176.514, 1126.01, 1376.636,
  146.6925, 179.7951, 169.8683, 144.5109, 115.9851, 100.912, 77.22723, 
    96.99864, 139.7948, 160.3108, 134.8792, 69.91695, 26.29307, 64.91444, 
    76.29048, 164.2859, 290.0237, 281.2162, 184.3736, 70.43913, 2.701435, 0, 
    0, 0, 0, 0.09234287, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.41791, 93.65132, 238.9857, 412.0441, 452.2166, 553.3406, 506.5167, 
    421.6122, 392.6665, 425.7772, 440.7444, 462.4359, 492.6555, 517.598, 
    531.2183, 527.7665, 529.114, 571.4398, 752.8386, 1117.882, 1654.942, 
    1618.519, 1398.75, 1202.588, 1191.508, 1195.801, 1221.172, 1415.927,
  69.31319, 104.212, 110.316, 83.84324, 63.33185, 52.58361, 41.60804, 
    45.76586, 76.87368, 101.9827, 93.67348, 33.04323, 20.12624, 46.1826, 
    54.88905, 34.84738, 115.9459, 49.21751, 40.83882, 0.5943004, 0, 0, 0, 0, 
    0, 0.0057942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.398386, 
    119.9112, 199.3601, 411.994, 476.3767, 578.0508, 529.0004, 436.2539, 
    335.8598, 335.8933, 358.957, 401.7341, 439.7245, 481.3549, 499.7074, 
    519.8088, 515.3641, 502.7769, 560.4839, 723.5606, 1163.4, 1705.951, 
    1771.096, 1455.29, 1286.019, 1198.102, 1179.159, 1260.96, 1461.374,
  79.25274, 98.79363, 46.67113, 25.34361, 28.43618, 24.51583, 16.18622, 
    19.50146, 37.39209, 67.61229, 56.61288, 32.74178, 14.21986, 3.174914, 
    2.647948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01747818, 46.90157, 207.9118, 460.4455, 514.9199, 
    602.9887, 590.7431, 513.9005, 364.6547, 319.0529, 315.5271, 335.9451, 
    373.1736, 425.5178, 449.45, 464.8029, 490.2738, 503.6892, 494.0532, 
    586.5953, 751.3316, 1115.167, 1723.364, 1792.263, 1481.577, 1256.694, 
    1160.092, 1138.162, 1189.935, 1531.006,
  304.3052, 225.9071, 146.4976, 49.22798, 14.06787, 15.70426, 14.31254, 
    10.55259, 21.65571, 34.42345, 26.47721, 10.16362, 1.715719, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3261773, 0, 0, 5.140869, 66.8336, 316.336, 486.2376, 557.2535, 
    481.0815, 482.611, 398.9484, 317.3685, 310.7681, 323.2128, 329.6191, 
    362.9882, 389.781, 416.3743, 421.8354, 456.8871, 480.976, 483.8488, 
    540.1299, 714.4539, 990.8341, 1670.664, 1620.258, 1494.627, 1232.962, 
    1134.55, 1134, 1203.068, 1431.174,
  377.3476, 300.3462, 179.3239, 123.5264, 29.18042, 8.49296, 10.41877, 
    2.594529, 2.675612, 3.391332, 0.1138654, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007269558, 0, 
    7.853471, 62.3085, 274.8862, 413.5488, 423.2161, 435.7926, 444.4748, 
    361.6428, 308.9561, 319.7975, 321.1809, 340.5662, 354.3437, 378.4564, 
    404.6211, 438.1272, 444.1309, 457.4094, 472.3898, 582.7078, 713.5034, 
    965.1596, 1325.418, 1513.297, 1287.996, 1268.213, 1155.886, 1135.109, 
    1137.983, 1441.737,
  397.6618, 290.1455, 262.0854, 164.1737, 72.91979, 9.641136, 3.297817, 
    0.002408294, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24.52353, 0, 1.134986, 131.7988, 
    413.9996, 487.4259, 485.74, 514.1754, 483.7487, 398.7583, 334.6064, 
    318.3876, 329.1971, 343.4026, 364.3184, 386.8412, 433.8055, 462.0353, 
    443.1543, 453.2259, 475.2897, 560.871, 675.3644, 778.7476, 1195.336, 
    1219.456, 1293.797, 1255.619, 1167.165, 1128.763, 1127.737, 1605.608,
  359.7442, 322.1634, 256.7101, 190.8573, 99.29717, 20.20619, 2.261762, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.042433, 1.061284, 0.06026918, 221.4693, 588.1027, 
    609.5046, 567.6266, 539.7374, 519.683, 443.9848, 375.9164, 330.9009, 
    328.2888, 345.5885, 367.2719, 396.1122, 425.6252, 436.9988, 445.1413, 
    455.4268, 478.2379, 538.37, 618.6725, 704.752, 879.9337, 1044.206, 
    1143.218, 1000.543, 1114.351, 1055.759, 1244.916, 1644.584,
  339.5918, 283.2596, 244.217, 182.1556, 115.8238, 16.9204, 1.281723, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 118.1892, 542.7286, 664.8825, 616.7386, 
    595.4612, 551.9771, 495.2496, 416.2375, 373.1087, 345.3355, 352.5166, 
    377.2891, 390.3913, 413.6357, 444.6428, 442.3636, 488.6983, 526.4742, 
    581.7993, 665.6102, 783.5282, 909.798, 1160.341, 1189.347, 1036.943, 
    1004.612, 1053.218, 1059.908, 1416.363,
  279.6242, 227.4193, 199.1174, 149.1774, 83.37285, 3.592551, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 101.2812, 60.90662, 478.8484, 643.0255, 690.905, 
    652.9017, 619.0784, 549.6542, 517.7484, 445.3293, 372.7345, 391.3872, 
    396.3501, 434.3335, 453.7928, 469.5943, 484.0396, 513.5276, 579.3093, 
    651.2834, 708.0594, 776.8271, 870.302, 1036.794, 1245.989, 901.5364, 
    940.5923, 1070.94, 1195.01, 1146.841,
  196.4323, 187.7343, 179.3497, 120.5639, 39.21375, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.005413, 45.81821, 62.24737, 21.02495, 
    3.207724, 0.02404907, 1.234567, 12.24459, 1.728072, 0, 0, 0, 0, 0, 0, 
    3.453561, 7.352701, 19.79626, 158.7443, 296.7885, 521.1622, 627.5361, 
    662.5475, 682.7275, 655.5103, 590.583, 580.2885, 526.9755, 427.6072, 
    407.3717, 430.1629, 446.7533, 474.6825, 500.0133, 519.8837, 559.5943, 
    617.9446, 655.3353, 686.9636, 713.472, 753.1322, 906.1678, 1018.012, 
    815.1847, 882.2279, 1056.679, 1259.787, 1045.098,
  141.7976, 159.4438, 144.7507, 76.36758, 7.418705, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.733681, 94.68479, 175.18, 187.5313, 
    155.0462, 110.0206, 72.29835, 93.21919, 121.2557, 115.5466, 66.30669, 
    6.150113, 0, 0, 0, 3.670892, 28.15756, 46.06707, 79.14339, 305.7281, 
    712.5394, 940.3807, 751.7666, 698.2665, 746.433, 768.7173, 723.7104, 
    672.3049, 616.0403, 509.8206, 453.0623, 453.5248, 504.1813, 528.5236, 
    544.4155, 565.7984, 598.8699, 625.6595, 655.5828, 686.7064, 683.7915, 
    732.2036, 789.5637, 840.5327, 723.5177, 745.4189, 965.6844, 1038.274, 
    796.5178,
  95.12392, 103.6217, 82.47251, 13.03405, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.002540734, 15.74638, 122.9433, 222.9018, 302.6361, 
    279.6983, 224.5893, 190.8986, 149.559, 188.5142, 236.7475, 212.6731, 
    150.321, 153.6949, 48.69242, 25.20141, 29.67488, 91.25098, 132.1451, 
    112.2913, 103.7838, 263.8452, 764.3199, 1062.096, 1009.38, 884.1952, 
    931.0499, 977.1282, 882.8214, 713.9742, 616.5552, 536.9384, 509.7403, 
    500.2069, 555.3665, 585.5272, 600.3098, 607.6362, 615.286, 634.0374, 
    661.1276, 645.6732, 626.6214, 638.4325, 669.1021, 625.0273, 530.0295, 
    528.0609, 601.1044, 644.5855, 548.4876,
  30.5022, 27.99392, 7.313161, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.7658302, 12.3739, 142.0602, 300.8344, 465.4789, 498.4969, 
    391.7122, 316.7618, 249.2353, 219.1284, 259.9997, 244.4664, 174.3858, 
    179.9653, 249.7257, 193.2922, 150.1301, 234.5797, 302.7541, 285.0494, 
    207.801, 158.7262, 115.508, 347.3649, 690.9739, 928.4409, 982.3543, 
    1030.41, 1034.681, 877.8196, 652.1367, 503.6282, 493.2419, 491.9219, 
    520.8734, 593.4538, 643.876, 652.7304, 662.8006, 652.0361, 676.1411, 
    653.5867, 602.203, 551.5805, 537.899, 522.2339, 492.5406, 445.3781, 
    430.9313, 431.1991, 487.3873, 602.6268,
  0.766829, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.8648, 
    83.18796, 276.2613, 500.1916, 600.5903, 597.6884, 475.5048, 352.7767, 
    314.1613, 281.9288, 287.8528, 237.377, 131.9863, 144.99, 306.4143, 
    294.3946, 305.1169, 332.2526, 310.4181, 229.8286, 185.2745, 224.0371, 
    255.049, 135.4041, 273.2138, 527.6912, 587.1231, 611.7789, 642.2618, 
    595.1403, 463.5603, 424.1609, 415.3838, 429.1796, 490.9037, 608.7256, 
    694.1671, 728.9787, 711.6575, 716.4285, 701.124, 642.769, 552.2159, 
    495.597, 465.6459, 440.4718, 429.3813, 424.0435, 422.3978, 418.5041, 
    446.8545, 718.7314,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.295444, 78.97375, 
    275.3757, 455.0948, 458.2011, 506.2027, 494.194, 412.8863, 375.2495, 
    355.046, 307.8675, 307.6067, 255.4145, 162.655, 174.7049, 269.6479, 
    362.2924, 358.3284, 318.2245, 211.9518, 198.9956, 327.952, 577.7234, 
    678.533, 449.4442, 258.9631, 309.9615, 318.2204, 354.7622, 372.4727, 
    407.3471, 409.3253, 394.0547, 388.1353, 397.6263, 455.2305, 588.9576, 
    706.325, 787.8987, 810.1958, 757.8834, 690.1829, 588.7928, 504.9205, 
    456.3733, 419.4193, 401.9965, 409.1686, 411.8871, 415.8695, 412.8529, 
    415.983, 653.3243,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04495476, 1.543852, 
    40.60966, 249.5493, 570.8077, 624.9529, 503.8392, 404.5659, 388.5279, 
    371.8024, 372.5071, 373.0171, 344.5746, 314.8991, 279.2988, 232.3392, 
    204.3131, 251.619, 321.1378, 336.9094, 265.9687, 241.0423, 314.6817, 
    503.8398, 693.5359, 810.1852, 579.9879, 386.7859, 384.9114, 418.0108, 
    446.1444, 373.0016, 350.7278, 352.2296, 366.1898, 378.6504, 386.957, 
    403.5961, 448.4445, 545.6042, 676.7407, 741.8482, 705.261, 612.5644, 
    508.2358, 457.7974, 419.8724, 397.5679, 394.2395, 399.4266, 405.9669, 
    407.882, 402.7976, 410.4689, 789.8555,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7914926, 10.71653, 
    37.00443, 201.4314, 448.087, 531.7697, 431.7727, 398.7067, 393.9764, 
    349.5272, 333.6953, 360.2705, 337.4265, 298.6373, 309.2917, 282.9134, 
    270.9925, 231.9091, 272.6257, 235.9534, 234.1443, 273.3409, 414.232, 
    561.9924, 633.738, 604.2332, 478.0908, 428.5763, 404.8661, 464.5562, 
    464.1216, 373.5608, 319.6164, 329.3439, 353.2355, 408.3477, 412.724, 
    410.5272, 419.3637, 448.9814, 538.6779, 576.0292, 562.1622, 501.3907, 
    457.8747, 424.4431, 405.648, 395.4491, 393.9858, 397.7108, 400.8848, 
    400.0156, 396.7203, 474.1039, 980.1252,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.459178, 23.89642, 
    39.5673, 52.56926, 168.347, 227.195, 285.7491, 353.7228, 381.3757, 
    362.791, 311.1005, 312.541, 320.0593, 289.4526, 308.0459, 311.635, 
    295.6172, 265.5541, 242.1341, 228.7672, 222.6893, 264.653, 356.3772, 
    481.8984, 514.7236, 444.572, 376.3537, 375.8529, 367.9664, 341.9634, 
    351.7896, 291.5329, 307.0333, 322.6101, 365.6251, 444.1953, 465.1169, 
    441.8697, 452.7754, 478.7091, 527.0575, 540.0756, 491.8977, 461.4532, 
    433.0887, 417.837, 414.4355, 413.9627, 410.6415, 421.8182, 400.1716, 
    394.3721, 399.2646, 611.9307, 1308.194,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.790205, 27.87427, 
    37.87522, 49.99376, 77.3848, 129.5688, 225.8023, 291.5181, 345.4376, 
    327.5065, 299.076, 285.3165, 292.4263, 320.6955, 306.0085, 310.2983, 
    291.4063, 262.9675, 246.8307, 238.5132, 249.1621, 271.4966, 326.77, 
    393.712, 450.9673, 416.2671, 374.2629, 344.2727, 333.5673, 305.9854, 
    280.9805, 285.871, 292.4921, 298.5072, 329.7079, 419.0633, 450.0066, 
    465.448, 502.8485, 574.8007, 637.0599, 703.0728, 587.3303, 483.8123, 
    452.7943, 442.7585, 455.8902, 478.3641, 513.434, 528.1032, 446.6922, 
    395.0017, 396.0436, 580.3947, 1096.152,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7.539374, 13.82793, 0, 0, 0, 0, 0, 0.3629586, 
    22.22618, 38.05198, 50.36842, 51.9423, 55.76481, 123.9351, 200.9567, 
    248.0657, 288.369, 296.5797, 284.997, 272.4008, 306.0285, 313.191, 
    326.7126, 292.9926, 277.2778, 264.6691, 265.5726, 260.786, 272.6996, 
    322.4322, 380.3541, 402.2595, 439.8839, 455.1393, 427.6396, 381.3865, 
    336.1739, 308.6934, 286.1038, 296.1768, 298.6016, 292.2509, 297.8213, 
    348.2343, 392.0045, 441.4889, 561.517, 686.3062, 815.3308, 935.5671, 
    875.5865, 574.7263, 510.7076, 481.0591, 505.4455, 569.8447, 637.2155, 
    645.5725, 578.0183, 406.8309, 416.0845, 555.6661, 828.242,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.968982, 31.56356, 1.362759, 0, 0, 0, 0, 0, 
    9.483889, 33.60556, 38.53296, 50.37358, 74.38406, 139.3567, 205.6824, 
    215.1312, 223.8199, 264.2617, 295.2328, 280.9891, 269.5547, 301.0195, 
    283.1612, 300.8699, 290.1711, 288.1376, 298.2253, 296.4409, 301.7662, 
    372.0651, 450.2336, 467.1264, 467.0771, 487.0597, 462.8398, 408.4555, 
    374.192, 332.696, 321.5491, 328.5142, 322.4901, 299.8736, 293.3217, 
    324.0511, 366.8441, 447.5163, 626.8708, 836.7401, 890.7211, 1096.81, 
    1047.843, 760.592, 575.9907, 540.1681, 540.2332, 595.8331, 628.45, 
    649.7249, 568.4493, 455.0399, 431.6068, 517.0565, 601.8608,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.797053, 7.747849, 3.450143, 0, 0, 0, 0, 0, 
    0.9109401, 18.42504, 39.59516, 52.26551, 97.90691, 235.892, 219.3992, 
    208.2924, 216.5296, 262.5898, 292.2108, 286.3712, 274.5794, 269.5547, 
    279.5371, 287.6822, 293.7041, 308.5545, 345.3323, 335.1651, 328.9469, 
    369.3367, 444.4053, 470.777, 502.3892, 510.839, 472.6234, 420.1351, 
    393.2463, 375.5051, 344.6975, 341.879, 320.9992, 295.3217, 288.8875, 
    310.2828, 356.9085, 436.3004, 643.2478, 908.5942, 908.9702, 1001.605, 
    1072.39, 855.878, 706.8087, 615.7324, 594.7244, 607.8818, 589.8001, 
    519.1802, 495.0875, 398.2069, 416.0681, 481.5428, 468.7679,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 45.77684, 0, 0, 0, 0, 0, 0, 0, 0, 19.37672, 
    35.37803, 69.18604, 153.2726, 288.3199, 317.8352, 244.572, 258.4949, 
    287.7384, 311.5768, 297.4268, 289.1551, 278.5264, 276.3994, 304.6932, 
    323.0869, 346.2746, 396.4057, 380.4884, 341.7323, 349.6577, 376.4726, 
    426.947, 504.5984, 651.9197, 501.9165, 434.0541, 415.7284, 411.0024, 
    387.9035, 340.0662, 290.0233, 265.8179, 252.4831, 284.6985, 349.8331, 
    406.4402, 572.5109, 805.2451, 886.5491, 902.3984, 984.8835, 957.6617, 
    842.1849, 709.3141, 604.957, 577.4132, 542.0748, 476.5501, 421.5896, 
    398.5287, 416.1053, 436.3309, 444.6508,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2233779, 7.883308, 
    46.45991, 63.79469, 184.3558, 336.8821, 374.0247, 374.8209, 335.6512, 
    339.178, 324.0201, 312.332, 293.5074, 275.675, 291.9893, 330.8283, 
    374.3214, 414.9174, 493.441, 464.5028, 388.4646, 358.354, 358.3539, 
    399.2584, 604.8146, 824.4387, 636.0546, 425.0211, 422.0507, 444.4562, 
    444.8008, 388.2694, 300.7451, 240.5886, 216.5688, 229.7297, 312.2461, 
    400.7599, 488.0696, 759.7354, 869.7776, 810.3863, 836.918, 927.7097, 
    906.3384, 778.0356, 610.2334, 542.7169, 508.4426, 490.6646, 424.6607, 
    396.6208, 405.9286, 424.3958, 467.8904,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.524688, 44.15213, 
    88.41959, 159.127, 276.4428, 370.4227, 392.6274, 382.1442, 366.4334, 
    336.8749, 317.2722, 299.4598, 286.5885, 283.6873, 292.2945, 335.28, 
    393.107, 469.711, 592.4265, 585.6436, 482.2569, 415.559, 389.8748, 
    408.3621, 619.8497, 895.7261, 639.1478, 447.5954, 410.7881, 450.1098, 
    465.333, 443.5472, 380.2547, 332.284, 295.5856, 256.3805, 299.0791, 
    379.3657, 547.1831, 780.5206, 955.9313, 825.8504, 679.0082, 745.6443, 
    771.3798, 700.3216, 547.1471, 488.1773, 493.5975, 534.8677, 465.9749, 
    408.6629, 406.9938, 428.9316, 486.2154,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.648079, 90.31952, 
    139.5776, 213.0849, 372.9224, 415.0632, 410.2803, 377.4778, 360.1422, 
    341.8087, 303.7456, 280.1181, 284.2162, 290.7113, 310.3253, 325.1641, 
    379.646, 458.2865, 595.5748, 642.431, 599.8919, 527.5738, 473.18, 
    483.1668, 614.2881, 799.8925, 603.7574, 431.5247, 413.0665, 434.388, 
    454.1592, 461.4271, 468.4397, 452.5511, 440.9289, 400.6418, 349.5063, 
    404.0337, 485.1346, 668.6317, 844.2675, 779.2899, 658.3606, 603.169, 
    619.9202, 579.0063, 475.0612, 424.7502, 455.7198, 513.4985, 468.9218, 
    415.5838, 421.0052, 460.8036, 482.3849,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.58741, 141.5162, 
    204.9548, 236.1427, 343.1058, 379.2624, 360.7214, 335.7108, 336.3476, 
    332.6995, 308.2321, 285.1463, 271.4974, 292.8643, 320.6105, 328.3786, 
    355.2569, 397.3354, 482.0117, 568.8033, 603.5388, 619.1583, 583.2557, 
    547.499, 603.738, 696.2391, 558.0874, 454.7069, 434.771, 488.2554, 
    465.5451, 480.1592, 528.2115, 662.0346, 767.2975, 774.6315, 505.6811, 
    453.9677, 500.7877, 584.0219, 721.4752, 757.2107, 622.8404, 564.5931, 
    553.7775, 544.0915, 438.6134, 401.1854, 402.1854, 448.803, 413.0183, 
    422.9466, 438.3102, 442.5483, 441.3457,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.301848, 158.3098, 
    258.9337, 303.8173, 299.6194, 299.056, 279.9115, 262.4927, 294.193, 
    317.6132, 308.028, 282.2506, 265.0864, 268.781, 299.4977, 330.493, 
    349.1855, 376.8177, 421.5884, 502.247, 599.8027, 734.8414, 890.7762, 
    678.5621, 700.035, 677.1342, 600.2327, 509.2974, 559.8538, 608.821, 
    538.714, 488.7658, 668.5876, 1060.59, 1373.92, 1418.137, 819.2729, 
    541.28, 535.3813, 612.2632, 721.4976, 746.7157, 652.4662, 555.7067, 
    576.511, 582.4625, 469.2462, 383.6081, 342.5653, 332.923, 354.656, 
    407.8102, 443.4485, 401.7837, 378.6187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 86.89892, 228.9686, 
    307.1906, 284.381, 247.07, 238.9294, 245.0831, 292.1502, 321.7906, 
    317.2473, 299.972, 288.464, 279.9789, 285.0193, 296.3184, 328.2048, 
    358.1512, 417.3985, 513.0966, 649.8973, 1018.273, 1282.382, 1139.754, 
    900.5889, 797.8112, 659.6571, 681.5824, 716.9097, 741.9376, 622.0638, 
    551.46, 815.8694, 1147.539, 1486.932, 1523.49, 1029.805, 601.8781, 
    552.1006, 578.9692, 660.6729, 721.0251, 691.4706, 615.808, 579.7531, 
    580.8895, 447.5938, 336.6733, 275.8545, 256.4472, 302.6965, 384.8403, 
    451.3116, 391.0798, 372.3258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.010157, 137.2761, 
    246.5296, 275.4832, 286.3332, 281.9478, 285.9474, 335.5515, 358.7326, 
    329.0612, 289.5595, 278.5055, 274.489, 270.4537, 278.7563, 306.5069, 
    345.374, 407.7699, 519.6101, 695.6252, 1020.536, 1431.428, 1296.497, 
    1159.715, 894.8511, 889.3289, 837.659, 898.1722, 824.8221, 688.373, 
    685.1447, 783.9781, 882.051, 899.179, 1132.87, 975.0953, 703.803, 
    579.3523, 556.1559, 602.6837, 672.3351, 701.9514, 668.7778, 612.2599, 
    538.6722, 430.2552, 334.1217, 260.4696, 247.4416, 300.6423, 367.5648, 
    419.1653, 385.3712, 385.5648,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57.55773, 181.7126, 
    294.1019, 358.642, 376.2969, 381.9689, 378.035, 391.0516, 372.8776, 
    348.465, 324.6873, 307.1947, 273.0872, 273.6699, 274.8869, 275.7082, 
    315.3789, 463.814, 693.0596, 959.1632, 1143.813, 1204.84, 1186.019, 
    1113.179, 1009.146, 981.3286, 895.3462, 765.3611, 644.151, 603.1124, 
    711.8834, 624.4473, 590.9575, 727.5765, 872.574, 675.1846, 577.9081, 
    544.3901, 554.0104, 578.1396, 636.2142, 666.0281, 591.5745, 499.7725, 
    416.1812, 362.9875, 301.6709, 266.8849, 341.4141, 365.0664, 373.7022, 
    355.0049, 393.6327,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.672453, 76.61076, 
    200.5678, 304.525, 397.0667, 442.379, 428.145, 388.1142, 388.5081, 
    408.9069, 422.5594, 380.0047, 325.1395, 271.7728, 229.48, 221.3898, 
    214.3802, 330.7382, 597.4027, 826.9779, 1010.901, 1106.384, 1267.898, 
    1164.386, 1014.269, 812.2874, 856.5626, 721.2389, 588.0623, 545.859, 
    605.4478, 543.02, 491.1708, 537.3549, 686.0102, 599.1124, 549.1641, 
    530.5813, 510.3197, 549.0093, 608.9304, 682.692, 603.2574, 419.0844, 
    360.2815, 332.0342, 312.2987, 297.1729, 354.3885, 423.995, 364.6626, 
    357.3581, 429.184,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.492652, 0, 5.913332, 0, 
    9.827749, 122.8932, 239.9646, 413.3958, 469.7688, 442.4698, 411.2574, 
    384.8907, 404.1997, 419.0803, 395.6619, 331.3684, 275.5099, 249.502, 
    270.0858, 300.564, 302.8828, 432.2428, 627.8237, 685.1678, 758.2089, 
    829.3271, 816.4886, 691.1724, 675.4188, 734.3888, 674.1106, 540.9742, 
    509.9907, 540.2866, 512.6861, 438.8988, 428.1956, 510.8031, 492.1108, 
    477.0582, 467.651, 481.3288, 477.3205, 570.1652, 742.3004, 660.6039, 
    434.6603, 307.3639, 286.5654, 295.7912, 296.1364, 355.3662, 457.1753, 
    393.4307, 396.5924, 493.4605,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.18091, 177.9759, 
    78.61066, 5.231147, 20.97725, 4.670784, 80.24761, 276.9565, 515.89, 
    480.1449, 420.3515, 475.0774, 450.7651, 429.4347, 397.8179, 353.9267, 
    293.7534, 272.3435, 388.218, 463.1545, 491.6412, 475.5977, 481.5441, 
    496.2309, 455.1932, 510.3101, 537.7867, 541.0651, 539.1157, 607.288, 
    534.366, 475.9772, 458.8337, 508.1748, 500.2999, 470.7975, 373.0616, 
    372.9929, 372.6212, 339.7219, 379.8255, 402.0655, 426.9336, 542.4205, 
    772.5742, 775.2917, 518.3701, 319.2849, 250.5893, 235.3483, 234.3458, 
    282.5884, 389.9496, 389.2494, 430.362, 541.4569,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42.64318, 0, 0, 0, 14.13362, 
    0, 0, 97.32533, 567.0143, 755.1489, 660.1171, 552.6977, 559.0915, 
    519.6163, 501.7351, 442.0413, 369.866, 317.342, 371.9945, 499.4051, 
    535.2877, 491.8406, 421.9243, 376.5453, 400.5975, 453.606, 510.7452, 
    552.5534, 541.176, 503.5962, 466.0743, 452.3511, 428.7473, 469.4224, 
    558.7114, 555.1274, 362.4989, 286.6256, 277.3649, 257.8876, 279.6031, 
    357.494, 406.6543, 470.3801, 647.2722, 685.0935, 537.283, 372.8993, 
    288.5817, 221.9755, 181.4825, 209.1741, 291.7701, 287.4789, 395.4302, 
    561.2106,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01953389, 0, 0, 0, 
    0, 0, 455.7978, 1051.609, 1211.341, 1040.144, 739.9411, 620.1765, 
    620.5828, 543.5131, 502.523, 425.7497, 412.7139, 442.9023, 449.829, 
    379.7539, 314.4379, 297.9188, 320.5314, 397.3131, 505.9446, 602.7551, 
    619.6101, 569.6279, 539.3142, 520.7625, 497.6906, 523.4991, 613.6224, 
    612.6038, 400.595, 262.5043, 224.5589, 204.1281, 205.329, 279.9945, 
    355.9917, 390.6264, 461.2118, 514.0649, 484.4973, 380.1658, 331.9442, 
    259.4583, 192.7791, 282.2837, 280.4692, 273.8584, 398.2701, 491.5527,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    524.9088, 1227.854, 1514.503, 1593.471, 1283.125, 835.2573, 726.7971, 
    681.4029, 629.7035, 589.2842, 510.3927, 473.1457, 430.4084, 306.1007, 
    237.6619, 228.5278, 244.4046, 284.5834, 374.7751, 497.4753, 605.6686, 
    636.1135, 616.2618, 595.865, 525.5728, 477.7885, 496.7985, 413.9014, 
    286.8343, 221.6673, 207.5997, 165.5916, 149.3675, 196.3652, 251.1849, 
    278.328, 301.5162, 361.5432, 350.5833, 304.2287, 281.5658, 276.7146, 
    189.8026, 362.6567, 363.6728, 247.8723, 372.7149, 441.053,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    109.9336, 398.2949, 940.3243, 1436.861, 1731.173, 1299.493, 1035.062, 
    902.295, 892.6244, 738.1326, 628.37, 557.6457, 490.0444, 346.9488, 
    207.4061, 175.4873, 181.6765, 210.3732, 258.1815, 368.8855, 533.0062, 
    620.7709, 626.9582, 508.8629, 400.888, 363.2095, 333.2734, 270.4286, 
    219.8917, 179.2967, 159.2247, 142.6616, 109.0908, 142.8433, 178.4309, 
    190.0326, 221.8169, 245.1929, 268.4247, 231.8128, 307.9815, 330.6054, 
    275.8257, 397.8697, 359.8254, 219.364, 334.6523, 463.7612,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06423091, 57.11491, 0, 0, 
    0, 0, 0, 0, 7.836217, 136.0153, 314.1614, 994.2757, 1493.946, 1517.679, 
    1301.398, 1272.304, 1158.99, 1018.497, 845.142, 688.6971, 603.6498, 
    439.0118, 236.4267, 146.054, 144.4927, 163.0123, 225.2119, 349.3079, 
    489.0631, 592.2128, 608.7792, 410.0895, 244.743, 193.4141, 256.4616, 
    227.5397, 197.2503, 107.2875, 83.52959, 68.98138, 80.46129, 115.9747, 
    132.9302, 145.9669, 152.7381, 174.7173, 173.7455, 175.6978, 235.3297, 
    318.201, 276.576, 340.2295, 316.9229, 225.2303, 420.5147, 420.0156,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.182514, 89.51676, 343.4627, 955.3691, 1260.624, 1151.738, 1138.569, 
    1236.952, 1157.061, 1085.779, 1005.899, 794.526, 562.4872, 299.4979, 
    123.4399, 98.68906, 119.4459, 185.4302, 329.3733, 361.4457, 432.3123, 
    502.7655, 379.1094, 146.3032, 62.53582, 92.53636, 99.53645, 60.84525, 
    11.73829, 14.53334, 21.45396, 50.65263, 84.13147, 89.0048, 93.22248, 
    110.0247, 112.9956, 145.8865, 186.0687, 228.4272, 220.4345, 204.2188, 
    252.7047, 291.9086, 311.514, 407.4745, 196.5356,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 37.47989, 422.1205, 709.343, 683.818, 813.1848, 1012.258, 1090.199, 
    1166.657, 1117.992, 963.0756, 744.8711, 327.3204, 67.59232, 51.20574, 
    51.10489, 136.7648, 215.8003, 145.3761, 67.80409, 186.2934, 218.4242, 
    88.11556, 0.4354767, 0, 0, 0, 0, 34.36349, 48.50853, 69.10825, 73.94706, 
    66.00063, 75.26979, 83.438, 52.38344, 29.00477, 151.119, 204.1204, 
    143.2567, 130.4681, 270.9427, 483.1219, 465.0688, 362.5184, 4.126702,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.66449, 261.7532, 151.233, 91.45276, 90.23305, 372.949, 595.9958, 
    811.2404, 1056.335, 1019.892, 820.1436, 449.4274, 159.2536, 109.9366, 
    231.9172, 190.1881, 121.1451, 13.04661, 0.002457884, 0.07684267, 
    1.469449, 0.02487941, 0, 0, 0, 0, 0, 69.92484, 163.3495, 125.5531, 
    119.3953, 127.3019, 150.9474, 169.9525, 115.3876, -54.83441, 78.6655, 
    169.3711, 172.5084, 110.4562, 298.2401, 618.7454, 450.6016, 111.6259, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18.18774, 198.2974, 24.82351, 0.01659623, 0, 9.641451, 62.01321, 
    362.3916, 663.819, 745.0246, 764.4761, 729.5575, 860.1415, 989.5406, 
    901.2372, 633.0322, 214.5284, 22.94515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    71.94882, 276.9225, 273.4788, 160.4362, 155.9303, 183.5391, 191.451, 
    188.135, 115.3398, 35.40816, 124.8625, 162.5711, 94.14777, 280.8703, 
    519.7524, 233.8496, 268.5618, 36.8153,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1127852, 103.1683, 83.84983, 125.6781, 310.4157, 588.7912, 843.4153, 
    526.3326, 1.147217, 0, 31.65186, 188.915, 342.4284, 556.4823, 714.2188, 
    878.2565, 858.4985, 833.0258, 646.3763, 302.5152, 38.86568, 0, 
    0.01003916, 0, 0, 0, 0, 0, 0, 0, 0, 50.22194, 269.6366, 109.4844, 
    37.02338, 59.75043, 26.35164, 79.59688, 104.9516, 76.24226, 67.52459, 
    111.2902, 103.7956, 226.3943, 374.5558, 285.326, 834.7192, 451.0992,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.3265, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.225108, 103.0244, 258.1696, 347.2978, 418.1593, 560.3155, 894.6843, 
    791.2195, 306.0076, 0.8998873, 0, 0, 0, 14.49841, 35.44591, 118.7575, 
    200.4224, 258.1529, 344.5415, 204.937, 28.87837, 0, 0.1383204, 0, 
    2.479101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01911015, 
    8.849098, 12.94733, 55.8584, 180.516, 374.3842, 761.2708, 606.065,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15.89997, 14.70358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37.67767, 140.6756, 246.9203, 375.567, 456.3772, 603.2179, 
    768.8178, 926.5468, 582.7935, 196.5176, 0, 0.4811277, 0, 0, 0, 0, 0, 0, 
    24.83666, 45.255, 12.15549, 2.415782, 0, 0.09825284, 1.407857, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6392468, 2.363386, 28.96285, 
    234.0622, 386.0693, 563.9972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17.55955, 29.1074, 15.34933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10.62364, 190.7695, 391.3156, 404.325, 600.9966, 680.045, 
    704.8675, 862.8046, 749.6393, 130.0502, 3.100419, 5.116066, 6.17757, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4328433, 76.46776, 242.6619, 291.0963, 5.134037, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8376673, 0, 0, 0, 0, 0, 0, 0, 0, 0.008186113, 
    0.07604827, 15.87589, 119.0556, 379.1627,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.163343, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 255.9357, 568.2272, 791.1302, 892.6254, 903.9981, 891.0063, 
    1059.328, 1098.428, 617.2275, 6.932829, 0.3629374, 65.03675, 7.93887, 0, 
    0, 0, 0.8275996, 112.0045, 17.52323, 0, 0, 57.19586, 246.4086, 451.7093, 
    100.6016, 0.06041526, 0, 0, 0, 0, 0, 0, 0.5732526, 182.9803, 198.6564, 
    161.3975, 11.53954, 0, 0, 0, 0, 0, 0, 0, 0, 0.992954, 173.7827,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.585627, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 257.8992, 621.7795, 752.3851, 846.557, 900.2053, 1019.242, 1113.99, 
    880.9015, 529.3146, 159.8383, 6.419941, 0, 0, 0, 0, 0, 0.03464887, 
    317.7343, 145.3232, 0, 0, 0.1035934, 0, 5.595896, 134.9415, 159.4373, 0, 
    0, 0, 0, 0.5597559, 213.3741, 71.13373, 0, 0, 10.51704, 18.63104, 
    3.763446, 0, 0, 0, 0, 0, 0, 0, 0, 34.35713,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.43994, 381.3143, 748.3234, 941.8181, 893.6531, 933.1523, 1035.22, 
    860.355, 610.6863, 554.7979, 525.4812, 498.002, 75.12685, 0, 0, 0, 0, 
    11.73125, 325.2318, 124.1923, 0, 0, 0, 0, 0, 42.32673, 450.324, 9.972672, 
    0, 0, 34.3005, 62.80934, 603.7728, 328.5521, 8.121914, 9.169447, 
    6.230115, 1.321965, 11.59744, 3.048517, 0, 0, 0, 0, 0, 0, 0, 6.704556,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30.85074, 297.304, 660.8721, 966.9948, 998.4858, 885.1306, 751.5646, 
    655.1858, 732.1314, 1084.44, 1349.639, 1119.806, 408.8793, 0, 0, 0, 0, 0, 
    140.0299, 7.918328, 0, 0, 0.1702392, 1.991248, 53.83979, 472.2008, 
    346.2012, 2.112901, 0.005206824, 0, 24.37175, 219.4124, 598.756, 
    329.5864, 98.26838, 18.94595, 28.95024, 2.492014, 22.5628, 50.42095, 0, 
    0, 0, 0, 22.81216, 24.65398, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26.93062, 106.7775, 98.48605, 75.9237, 51.93491, 62.07972, 66.57274, 
    176.725, 422.3495, 479.3473, 519.7673, 215.12, 2.231832, 0.004072465, 
    1.405816, 0.08232938, 0, 495.7819, 40.24272, 0, 7.263184, 112.9553, 
    325.7667, 421.6084, 533.7393, 301.4734, 91.60561, 24.09392, 33.98492, 
    380.9341, 705.0402, 632.1104, 263.1127, 138.8074, 37.80578, 1.129739, 
    35.61073, 95.76726, 325.1597, 511.9413, 832.47, 77.51266, 0, 41.77975, 
    292.1154, 30.66951, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 23.8246, 73.93395, 126.2193, 321.1346, 494.5471, 
    282.6015, 106.8233, 331.644, 202.062, 0, 24.80076, 24.1915, 49.88836, 
    269.6974, 671.1443, 778.3289, 494.5531, 183.3987, 40.72751, 10.41955, 0, 
    92.49084, 767.71, 1000.381, 579.1232, 178.2135, 9.95975, 6.408473, 
    10.95331, 70.58002, 197.3521, 552.4769, 928.8527, 1256.867, 539.4283, 
    47.92098, 154.266, 98.49847, 27.90792, 1.357446 ;
}
