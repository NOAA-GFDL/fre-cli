netcdf atmos.1980-1981.alb_sfc.04 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:17 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.04.nc reduced/atmos.1980-1981.alb_sfc.04.nc\n",
			"Mon Aug 25 14:40:04 2025: cdo -O -s -select,month=4 merged_output.nc monthly_nc_files/all_years.4.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  10.17506, 10.34687, 10.39664, 10.04403, 10.37535, 10.30696, 10.37304, 
    10.49578, 10.32739, 10.31409, 10.77876, 10.35706, 10.36029, 10.56685, 
    10.57548, 10.62285, 10.55661, 10.49646, 10.1098, 10.07648, 10.09658, 
    10.23055, 9.94339, 10.11824, 10.08967, 10.60355, 10.58841, 10.59269, 
    10.33088,
  19.00928, 21.95174, 17.02231, 23.46513, 27.66054, 27.62418, 30.24759, 
    27.77559, 27.74319, 27.85352, 27.51577, 27.36524, 27.67224, 16.6535, 
    8.171993, 6.117301, 6.300015, 3.363888, 3.108542, 3.818256, 14.28573, 
    13.49114, 25.43802, 28.50901, 30.97534, 27.81471, 15.67716, 5.820986, 
    19.04185,
  3.649509, 3.711534, 4.148434, 3.80628, 3.921348, 3.752871, 3.739745, 
    3.816878, 3.658071, 3.685964, 3.914557, 3.421335, 3.186375, 3.552358, 
    3.920477, 3.793256, 3.521006, 3.37693, 3.52585, 3.617719, 3.616264, 
    3.437983, 3.344326, 3.670508, 3.279581, 3.391854, 3.247155, 3.612114, 
    3.698802,
  3.425123, 3.543334, 3.489604, 3.717349, 3.711251, 3.504045, 3.72509, 
    3.743647, 3.803928, 3.674218, 3.586309, 3.644969, 3.641523, 3.735444, 
    3.785143, 3.782576, 3.773204, 3.728181, 3.596585, 3.635291, 3.423252, 
    3.461358, 3.685841, 6.673156, 3.952131, 3.838429, 3.802125, 3.692227, 
    3.546192,
  3.667484, 3.592069, 3.817947, 3.774054, 3.641324, 3.743829, 3.767117, 
    3.684308, 3.637321, 3.696648, 3.631402, 3.714461, 4.182073, 4.02251, 
    8.091396, 3.782749, 3.77611, 3.544719, 3.764357, 3.64257, 3.671102, 
    3.736082, 3.760887, 7.992327, 4.095751, 3.889305, 3.829881, 3.838686, 
    3.544152,
  3.922848, 3.875879, 11.30232, 3.76468, 3.828202, 3.812728, 3.628883, 
    3.863199, 3.539303, 4.024624, 8.984606, 13.47036, 9.536808, 3.973724, 
    3.845654, 3.665733, 3.732253, 3.570317, 3.68306, 3.562364, 3.570363, 
    3.902476, 3.863683, 4.29673, 8.449537, 3.823218, 3.546736, 3.841413, 
    3.71239,
  3.604418, 9.474848, 9.74848, 3.650055, 3.528545, 3.534727, 3.436677, 
    3.69836, 3.447464, 3.844562, 12.0921, 11.43484, 3.671887, 3.650176, 
    3.471658, 3.447522, 3.550918, 3.464666, 3.74015, 3.726095, 3.876029, 
    3.730717, 3.457626, 3.440653, 8.686346, 8.855945, 3.666655, 3.85588, 
    3.67703,
  3.312147, 6.464054, 8.699188, 8.565091, 3.410318, 3.340126, 3.213651, 
    3.433171, 3.248914, 3.334031, 4.521204, 3.440553, 4.099717, 3.317961, 
    3.429661, 3.200667, 3.404907, 3.61327, 3.509827, 3.638924, 3.694595, 
    3.453199, 3.229338, 8.627817, 8.159281, 8.787914, 3.738759, 3.444099, 
    3.491243,
  3.085088, 8.404028, 8.187752, 9.708523, 3.483654, 3.530845, 3.508086, 
    3.38312, 8.610996, 8.175154, 3.281808, 3.305061, 3.157861, 3.422521, 
    3.363621, 3.46149, 3.458388, 3.527724, 3.47356, 3.451664, 3.458107, 
    3.421351, 3.261666, 8.20139, 8.325867, 3.323549, 3.199236, 3.243976, 
    3.09024,
  10.12701, 10.45427, 10.47324, 9.854937, 15.00554, 3.250327, 5.317032, 
    3.361509, 3.609287, 3.387492, 4.487518, 3.294055, 3.414907, 3.276591, 
    3.220608, 3.359467, 3.271201, 3.311265, 3.333187, 3.377179, 3.222859, 
    3.434927, 8.879153, 7.552234, 3.525756, 3.281205, 3.129554, 3.212574, 
    8.847616,
  18.17624, 20.83453, 22.87333, 3.566541, 22.7756, 3.525362, 10.93584, 
    3.464999, 9.91872, 3.274202, 3.605289, 3.609395, 3.761668, 3.801834, 
    3.754453, 3.877979, 3.59555, 3.801422, 3.355684, 3.554606, 3.63324, 
    6.545098, 3.729053, 4.371435, 3.862963, 3.501264, 3.593875, 3.442076, 
    23.69124,
  24.06986, 20.33024, 21.01896, 19.51342, 12.65938, 14.35067, 12.61054, 
    18.56179, 8.785735, 10.16657, 3.466849, 3.470922, 3.41175, 3.495042, 
    3.63209, 3.563735, 3.526203, 3.815447, 3.490995, 3.928687, 10.50747, 
    11.85238, 9.369282, 3.581663, 3.803839, 3.596276, 3.771416, 3.655037, 
    11.41738,
  7.765381, 4.086432, 6.013519, 10.90557, 2.09387, 15.4515, 17.82203, 
    15.4425, 13.44672, 10.99661, 8.152763, 3.811582, 3.750215, 3.789702, 
    3.712769, 3.683611, 3.693204, 3.805667, 3.627367, 12.20406, 11.70161, 
    14.42378, 13.58505, 4.551152, 3.780712, 3.791294, 3.778115, 3.772772, 
    5.300657,
  6.06729, 12.56274, 15.14699, 16.13959, 13.54663, 18.02957, 9.101006, 
    37.50301, 11.27762, 8.376409, 8.203783, 19.17479, 11.18044, 4.101985, 
    4.11036, 4.222049, 4.093166, 4.031904, 4.210052, 21.27369, 11.73486, 
    15.35893, 21.06082, 32.20111, 10.18414, 3.802861, 4.014256, 4.359132, 
    4.244776,
  4.73652, 13.7879, 16.50302, 18.34985, 21.65412, 18.8244, 27.42126, 
    34.27948, 28.79816, 30.23542, 26.37563, 45.13363, 46.19276, 40.32684, 
    11.79234, 30.68948, 35.72057, 18.39208, 41.09412, 14.49545, 18.53337, 
    44.19654, 53.46863, 46.30341, 4.543104, 11.67899, 5.190823, 4.885833, 
    4.767662,
  5.22267, 5.87256, 32.10634, 5.723254, 45.7923, 55.96578, 51.44799, 
    52.06663, 52.08028, 51.43078, 37.40095, 32.54665, 51.7729, 61.06168, 
    60.62331, 61.73666, 54.94989, 54.04713, 59.06818, 58.58297, 51.47298, 
    57.09022, 53.18268, 52.66552, 60.6999, 52.58768, 52.42189, 57.15929, 
    5.598478,
  77.02435, 73.35914, 74.04105, 77.1144, 76.28472, 77.30383, 80.36185, 
    81.08687, 81.46243, 82.12009, 82.125, 82.15228, 81.97961, 81.79935, 
    81.9388, 82.09886, 82.0745, 81.82104, 81.69016, 81.78006, 81.72695, 
    77.22157, 71.78038, 72.82487, 69.39729, 68.93155, 69.23479, 70.63942, 
    80.96623 ;

 average_DT = 730 ;

 average_T1 = 106 ;

 average_T2 = 836 ;

 climatology_bounds =
  106, 836 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
