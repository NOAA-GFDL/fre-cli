netcdf atmos_month.198001-198012.aliq {
dimensions:
	time = UNLIMITED ; // (12 currently)
	pfull = 65 ;
	lat = 2 ;
	lon = 2 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:cell_methods = "time: mean" ;
		aliq:interp_method = "conserve_order2" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:10 2025" ;
		:hostname = "pp033" ;
		:history = "Tue Sep 23 14:27:36 2025: ncks -d lon,0,1 atmos_month.198001-198012.aliq.nc_lat01 atmos_month.198001-198012.aliq.nc_lat01_lon01\n",
			"Tue Sep 23 14:26:17 2025: ncks -d lat,0,1 atmos_month.198001-198012.aliq.nc atmos_month.198001-198012.aliq.nc_lat01\n",
			"Mon Aug 11 16:16:54 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198001-198012.aliq.nc reduced/atmos_month.198001-198012.aliq.nc\n",
			"Mon Aug 11 20:02:14 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.3.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -1.903176e-05, 0,
  0, 0,
  0.0121547, 0.008161363,
  0, 0,
  0.06501345, 0.02135089,
  8.785783e-09, 5.590953e-09,
  0.1428165, 0.08510327,
  0.002939393, 0.001987103,
  0.2557682, 0.1874608,
  0.05468941, 0.05095281,
  0.2539347, 0.2629735,
  0.07082365, 0.06972443,
  0.2560496, 0.269366,
  0.07199486, 0.06983482,
  0.228195, 0.2628424,
  0.09812149, 0.09578804,
  0.2298899, 0.2502919,
  0.1267387, 0.1250323,
  0.2373341, 0.2178164,
  0.1310529, 0.1308487,
  0.2460021, 0.2085861,
  0.1995048, 0.2002687,
  0.2216481, 0.2018702,
  0.2625196, 0.2618038,
  0.2523988, 0.2091967,
  0.255346, 0.2593552,
  0.2741496, 0.2189191,
  0.2551941, 0.2605655,
  0.2815016, 0.2265071,
  0.2703033, 0.2749571,
  0.229144, 0.2730744,
  0.2689278, 0.2741974,
  0.1832122, 0.2486309,
  0.2748757, 0.2809682,
  0.1385254, 0.198225,
  0.216422, 0.2239572,
  0.1053532, 0.1415415,
  0.1407903, 0.1463517,
  0.07865272, 0.1105382,
  0.09309179, 0.09744438,
  0.0689756, 0.1030117,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, -1.757755e-08,
  1.550498e-05, 5.04163e-06,
  -0.0008809567, -4.098656e-05,
  0.007066551, 0.006271057,
  0.006030335, 1.379079e-05,
  0.03892121, 0.03680561,
  0.08309711, 0.01622687,
  0.07216924, 0.06890453,
  0.08641893, 0.06942788,
  0.09311233, 0.0903368,
  0.07210723, 0.06494962,
  0.08248186, 0.08157716,
  0.0509961, 0.0549494,
  0.08843844, 0.08719351,
  0.04479598, 0.04906452,
  0.09118559, 0.08987503,
  0.04027409, 0.04334169,
  0.100023, 0.09964643,
  0.04200535, 0.04575753,
  0.1149001, 0.1144186,
  0.04214699, 0.04915907,
  0.1242735, 0.1244703,
  0.03330694, 0.05728827,
  0.1733709, 0.1712074,
  0.0263656, 0.05740754,
  0.2691303, 0.2681251,
  0.02007959, 0.0535381,
  0.3860271, 0.3870821,
  0.02894714, 0.0717443,
  0.4845036, 0.4915984,
  0.03050267, 0.08193073,
  0.5371985, 0.5458538,
  0.04646148, 0.09572122,
  0.5117947, 0.5172998,
  0.06510687, 0.08072527,
  0.386596, 0.3897896,
  0.07288758, 0.06823067,
  0.2883959, 0.2918073,
  0.08649805, 0.07038835,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.001269084, 0,
  0, 0,
  0.003174752, -0.0001079531,
  0, 0,
  0.0223729, 0.004021255,
  0, 0,
  0.06323196, 0.03809451,
  0.002499975, 0.001813969,
  0.1488183, 0.03445232,
  0.03642909, 0.03419077,
  0.3008322, 0.05210298,
  0.07355022, 0.06964004,
  0.3423942, 0.1291718,
  0.1716236, 0.1668534,
  0.3654023, 0.2743756,
  0.2285265, 0.2252701,
  0.3632489, 0.3423707,
  0.3042807, 0.3001232,
  0.342408, 0.3600067,
  0.3715583, 0.3692498,
  0.3142951, 0.3875316,
  0.4237208, 0.4234163,
  0.2903997, 0.4068105,
  0.4688378, 0.469766,
  0.3047067, 0.4441353,
  0.4858305, 0.4872543,
  0.322566, 0.5097123,
  0.4968948, 0.4935788,
  0.3785984, 0.5892029,
  0.3602235, 0.3580395,
  0.4308827, 0.5595596,
  0.2271547, 0.227679,
  0.4199008, 0.4808587,
  0.07568359, 0.07368695,
  0.395285, 0.4188643,
  0.04348774, 0.04363547,
  0.4133147, 0.325191,
  0.03229425, 0.0320038,
  0.3281704, 0.2329517,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0006693949, -7.566133e-06,
  4.385775e-05, 4.385775e-05,
  0.0004087718, -4.93201e-05,
  0.0001984276, 0.0001812432,
  0.01354727, -0.000234678,
  0.01256921, 0.01144051,
  0.03691494, 0.007345036,
  0.02753257, 0.0255592,
  0.06373479, 0.03909881,
  0.07186773, 0.06564563,
  0.08012234, 0.04464604,
  0.1588344, 0.1500731,
  0.1115285, 0.07558514,
  0.2562161, 0.2474208,
  0.1241159, 0.09782873,
  0.3003374, 0.2942557,
  0.1187288, 0.1074577,
  0.3328915, 0.3284591,
  0.1172309, 0.1252135,
  0.3681359, 0.3673311,
  0.1230053, 0.1438777,
  0.400963, 0.403028,
  0.1305353, 0.1695595,
  0.4257114, 0.4279828,
  0.1477159, 0.1868984,
  0.4513431, 0.4535102,
  0.1757396, 0.2471377,
  0.4753781, 0.4742626,
  0.2376152, 0.3482167,
  0.3653514, 0.3618405,
  0.2853765, 0.3674977,
  0.2737293, 0.2692288,
  0.312907, 0.3103174,
  0.1920229, 0.1834596,
  0.3483743, 0.2742096,
  0.1678627, 0.1660403,
  0.3435206, 0.2074582,
  0.1657239, 0.1641073,
  0.2655927, 0.1419661,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  4.244298e-05, 4.244298e-05,
  -2.760227e-05, 0,
  0.002817712, 0.002147224,
  -9.475026e-05, 0,
  0.06244681, 0.05529452,
  -0.001292572, -2.575446e-05,
  0.1596455, 0.1557184,
  0.01434967, -0.0008734533,
  0.2365951, 0.235928,
  0.0607516, 0.002980232,
  0.2527589, 0.2539192,
  0.1002498, 0.03602106,
  0.3013707, 0.3044307,
  0.1283372, 0.1003454,
  0.3261281, 0.3284515,
  0.1389281, 0.1957614,
  0.3658895, 0.3689875,
  0.1516593, 0.2509073,
  0.4102564, 0.4145253,
  0.1815312, 0.3070099,
  0.4384012, 0.4430297,
  0.2070991, 0.3335978,
  0.4339935, 0.4381829,
  0.2452309, 0.3665509,
  0.3853813, 0.3901182,
  0.2860303, 0.365562,
  0.2851419, 0.2876454,
  0.3023286, 0.3388455,
  0.2236998, 0.2233455,
  0.3218701, 0.2817795,
  0.1599583, 0.156792,
  0.3757266, 0.2360641,
  0.1298458, 0.1275699,
  0.4501016, 0.1901356,
  0.1142291, 0.1111387,
  0.3889688, 0.1094372,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.002399456, 0,
  1.073616e-06, 3.451996e-07,
  -0.001885479, 0,
  0.001102697, 0.0006314904,
  0.02886408, -0.00110208,
  0.02229615, 0.01872572,
  0.06581829, 0.005058833,
  0.07222524, 0.06773897,
  0.1017247, 0.04196965,
  0.1152714, 0.1120449,
  0.1259371, 0.1177407,
  0.1255099, 0.1244332,
  0.1567555, 0.1483307,
  0.1449172, 0.1426661,
  0.1848758, 0.1825048,
  0.1756151, 0.1719283,
  0.2189726, 0.1882457,
  0.2020522, 0.1982561,
  0.227085, 0.1913392,
  0.2222029, 0.2180355,
  0.2318976, 0.20593,
  0.1960303, 0.1936831,
  0.2712145, 0.2228032,
  0.1526051, 0.1496233,
  0.2593804, 0.2424669,
  0.03631271, 0.03447295,
  0.2502342, 0.1715394,
  0.01062638, 0.01064972,
  0.2399901, 0.1106699,
  0.004458392, 0.004630582,
  0.1668659, 0.076603,
  0.003017554, 0.003269679,
  0.1405581, 0.02841221,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -9.909024e-05, -4.007819e-06,
  1.341797e-05, 3.779102e-06,
  -0.002178703, -0.0002003084,
  6.10212e-05, 5.603315e-05,
  -0.005564602, -0.0008649079,
  0.0004863774, 0.0004109764,
  0.03698276, 0.007683921,
  0.009834158, 0.009580641,
  0.08800703, 0.01513108,
  0.02420903, 0.02415885,
  0.1042449, 0.04537813,
  0.04153079, 0.04124913,
  0.1175527, 0.09448731,
  0.0599519, 0.0574755,
  0.1174143, 0.1103957,
  0.08444641, 0.07964391,
  0.09850796, 0.1200001,
  0.1390322, 0.1334855,
  0.0782954, 0.1083198,
  0.1642184, 0.159615,
  0.07852578, 0.1151201,
  0.2157677, 0.2129067,
  0.08349716, 0.1126601,
  0.2232485, 0.2196473,
  0.08397945, 0.09468019,
  0.1200811, 0.1160422,
  0.08360814, 0.05772583,
  0.03526216, 0.03352587,
  0.06743748, 0.05211816,
  0.01526833, 0.01406171,
  0.06677447, 0.06787933,
  0.007301806, 0.006589465,
  0.05158073, 0.04500922,
  0.006030517, 0.005746993,
  0.01315673, 0.01630084,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0001481954, 9.430615e-05,
  -0.003089417, 0,
  0.01355244, 0.01171181,
  0.02348906, -4.27804e-05,
  0.02967546, 0.02777132,
  0.122583, -0.005069637,
  0.05576523, 0.051435,
  0.1631925, 0.01606301,
  0.1170336, 0.1128706,
  0.2129585, 0.05194824,
  0.1466008, 0.1404632,
  0.2292565, 0.1133222,
  0.2039614, 0.1972816,
  0.2318809, 0.1477728,
  0.2218536, 0.2178232,
  0.2319861, 0.1528771,
  0.2261455, 0.2239303,
  0.2264886, 0.1551652,
  0.2194332, 0.218079,
  0.2210793, 0.1512545,
  0.1769586, 0.1744665,
  0.2225234, 0.1258079,
  0.09321445, 0.09017443,
  0.2157615, 0.1073802,
  0.02515564, 0.02247247,
  0.1819369, 0.09167586,
  0.01440501, 0.01380268,
  0.1586076, 0.06623261,
  0.003076577, 0.003191179,
  0.06755415, 0.03215805,
  0.00251772, 0.002610245,
  0.02413257, 0.01362237,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0005570832, 0,
  0, 0,
  0.002879241, -0.0003239195,
  0, 0,
  0.01253692, 0.00167431,
  1.881689e-05, 1.200311e-05,
  0.06458889, 0.006456007,
  0.003274292, 0.002119844,
  0.09254536, 0.02910665,
  0.04760399, 0.0384461,
  0.1480272, 0.06183461,
  0.168439, 0.1551169,
  0.1690663, 0.07180968,
  0.2528341, 0.2436806,
  0.1832339, 0.08408518,
  0.286597, 0.2815888,
  0.1986619, 0.09331097,
  0.3021533, 0.2996509,
  0.2091256, 0.106077,
  0.2722183, 0.2704413,
  0.2283738, 0.1207343,
  0.2331161, 0.2317068,
  0.2175328, 0.1341003,
  0.1082781, 0.1056106,
  0.2153779, 0.1122836,
  0.005673736, 0.005389275,
  0.2400678, 0.08253906,
  0.003098136, 0.003332698,
  0.2325847, 0.07793682,
  0.002048941, 0.002089897,
  0.1668127, 0.07191476,
  0.001871879, 0.001887264,
  0.1019444, 0.04080886,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -1.821549e-05, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.005257796, 0,
  0, 0,
  0.01892745, -0.0002736447,
  0.0003883444, 0.0002716848,
  0.1073103, -0.002577145,
  0.008033142, 0.005041669,
  0.2343454, 0.003473091,
  0.07106643, 0.06676165,
  0.2541608, 0.07001664,
  0.09580622, 0.08998394,
  0.2487421, 0.1963657,
  0.1480571, 0.1438056,
  0.2455886, 0.2686774,
  0.1537506, 0.1504861,
  0.2547307, 0.2704693,
  0.1418939, 0.1407577,
  0.2596151, 0.275584,
  0.1262513, 0.1254863,
  0.281264, 0.2809329,
  0.1132192, 0.1117519,
  0.3080943, 0.2932978,
  0.09338196, 0.09071989,
  0.3187168, 0.2886704,
  0.05107618, 0.04976555,
  0.3126582, 0.2743697,
  0.02197386, 0.01974013,
  0.2898149, 0.2412924,
  0.004051184, 0.003536265,
  0.2746014, 0.2083342,
  0.001986551, 0.001687597,
  0.2511431, 0.09400836,
  0.001809807, 0.001398553,
  0.2245727, 0.04111981,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.005807792, 0,
  0, 0,
  0.04682167, -0.001002102,
  0.002258079, 0.001228736,
  0.1150018, 0.01118559,
  0.08450992, 0.07685507,
  0.1499721, 0.04051647,
  0.1784922, 0.1723485,
  0.1824355, 0.07230795,
  0.238776, 0.2337206,
  0.216827, 0.1110514,
  0.2799259, 0.2782658,
  0.2196311, 0.1588986,
  0.3002201, 0.297475,
  0.2242833, 0.1812991,
  0.3265011, 0.3241398,
  0.2296282, 0.2018863,
  0.3487751, 0.3470336,
  0.2373523, 0.2307075,
  0.3528084, 0.3508893,
  0.241697, 0.2572981,
  0.3925946, 0.3916629,
  0.2417884, 0.2529759,
  0.4333732, 0.435076,
  0.2514358, 0.2597913,
  0.42853, 0.4325115,
  0.2448828, 0.2613389,
  0.4127883, 0.414814,
  0.2140058, 0.246437,
  0.3317362, 0.3338371,
  0.1811901, 0.2120274,
  0.2489596, 0.2506604,
  0.1539144, 0.1544172,
  0.1813499, 0.1831295,
  0.1586418, 0.1348162,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.003990239, 0.002360163,
  -0.001139022, -2.046406e-05,
  0.06727315, 0.06590822,
  0.03966309, -0.001063082,
  0.08475678, 0.08434079,
  0.1126059, 0.01425214,
  0.1425587, 0.1371274,
  0.1224593, 0.1008512,
  0.2133387, 0.2105108,
  0.1348311, 0.1685959,
  0.2245434, 0.2263062,
  0.1282396, 0.1872784,
  0.2106881, 0.2120548,
  0.1223254, 0.180681,
  0.1849882, 0.1856724,
  0.1176915, 0.1657309,
  0.1654041, 0.1652822,
  0.1161799, 0.1485025,
  0.1573271, 0.1572207,
  0.1193676, 0.1459998,
  0.1429823, 0.1426574,
  0.1207952, 0.1669818,
  0.139992, 0.1406398,
  0.1649158, 0.192272,
  0.2284337, 0.2263003,
  0.1803104, 0.2126425,
  0.3125763, 0.3141736,
  0.2280552, 0.2292765,
  0.3295633, 0.3325611,
  0.2022519, 0.2286711,
  0.2736285, 0.2775607,
  0.1516945, 0.1765874,
  0.2197597, 0.2236073,
  0.1146186, 0.1284907,
  0.1388423, 0.1424826,
  0.08461437, 0.09215746,
  0.1068983, 0.1095244,
  0.06781885, 0.06706832,
  0.07674241, 0.07860156,
  0.06298608, 0.05691301 ;

 lat = -89.5, -79.5 ;

 lat_bnds =
  -90, -89,
  -80, -79 ;

 lon = 0.625, 13.125 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 380.5, 410.5, 440.5, 471, 501.5, 532, 562.5, 593.5, 624, 654.5, 685, 
    715.5 ;

 time_bnds =
  365, 396,
  396, 425,
  425, 456,
  456, 486,
  486, 517,
  517, 547,
  547, 578,
  578, 609,
  609, 639,
  639, 670,
  670, 700,
  700, 731 ;
}
