netcdf \00010101.huss.atmos_daily.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float huss(time, grid_yt, grid_xt) ;
		huss:_FillValue = 1.e+20f ;
		huss:missing_value = 1.e+20f ;
		huss:units = "1.0" ;
		huss:long_name = "Near-Surface Specific Humidity" ;
		huss:cell_methods = "time: mean" ;
		huss:cell_measures = "area: area" ;
		huss:coordinates = "height2m" ;
		huss:time_avg_info = "average_T1,average_T2,average_DT" ;
		huss:standard_name = "specific_humidity" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:_FillValue = NaN ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 huss =
  0.0007530822, 0.0008768799, 0.0009092166, 0.0009961284, 0.0008377059, 
    0.0006539731, 0.0006554869, 0.0006321146, 0.0006374769, 0.0003675956, 
    0.0003955099, 0.0004174119, 0.0002630356, 0.0002883163, 0.0001339794,
  0.0009561618, 0.0009128363, 0.0008647798, 0.0009378794, 0.0007641964, 
    0.000571433, 0.0005947688, 0.0005371174, 0.0005777993, 0.0005743248, 
    0.000425976, 0.0005255786, 0.0005168005, 0.0002419239, 0.0001384041,
  0.0009307395, 0.0008935601, 0.0008646884, 0.0008629375, 0.0007758569, 
    0.000447036, 0.0005087287, 0.0005155887, 0.0005337982, 0.0005408757, 
    0.0005119591, 0.0005206638, 0.0005404028, 0.0005288417, 0.0003520976,
  0.00113384, 0.0008631091, 0.0007961398, 0.000777832, 0.0007899554, 
    0.0006982922, 0.0002854749, 0.0004015622, 0.0005369425, 0.0004798827, 
    0.0004437493, 0.0004648793, 0.0004996103, 0.0005274226, 0.0004602039,
  0.001308236, 0.0009967769, 0.0007881733, 0.0007331111, 0.0007056717, 
    0.0007090645, 0.0006824931, 0.0002410056, 0.0002850571, 0.000307249, 
    0.0003930083, 0.0004322271, 0.0004758358, 0.0005212312, 0.0005475282,
  0.001277564, 0.001101121, 0.0008742156, 0.0007632893, 0.0007157979, 
    0.0006666422, 0.0006203346, 0.000634043, 0.0004587235, 0.0003683333, 
    0.0003368547, 0.0004292976, 0.000463269, 0.0005085627, 0.0005444105,
  0.001292239, 0.001102979, 0.0009468182, 0.0008127367, 0.0007604, 
    0.000716044, 0.0006858966, 0.0006329794, 0.0005738842, 0.0005391051, 
    0.0005011102, 0.0004579447, 0.0004766339, 0.0004995739, 0.0005359706,
  0.001269325, 0.001140613, 0.0009690849, 0.0008696977, 0.0007979057, 
    0.0007449095, 0.0007039802, 0.0006580271, 0.0006178524, 0.000594656, 
    0.0005557326, 0.000506365, 0.000502655, 0.0005263335, 0.0005416659,
  0.001244844, 0.001108353, 0.0009590478, 0.00087578, 0.0008185451, 
    0.0007577097, 0.0007120819, 0.0006731761, 0.0006527828, 0.0006173366, 
    0.0005922007, 0.0005354744, 0.0005365719, 0.0005552122, 0.0005691127,
  0.00120875, 0.001076314, 0.0009777534, 0.0009040253, 0.0008143926, 
    0.0007660507, 0.000730239, 0.0006923698, 0.0006145052, 0.0004795597, 
    0.0005147595, 0.0005403934, 0.0005401413, 0.000535469, 0.0005393531,
  0.0008980546, 0.001073442, 0.0007530436, 0.0007996496, 0.0007115795, 
    0.0006337609, 0.0006757569, 0.000664669, 0.0005938851, 0.000487438, 
    0.0006053591, 0.0006448331, 0.0005523701, 0.0005115941, 0.0003655333,
  0.0009984722, 0.0009372503, 0.0009599963, 0.0008575451, 0.0006437195, 
    0.0006573037, 0.000687752, 0.0006974107, 0.0006615157, 0.0005874933, 
    0.0006035316, 0.0006897251, 0.0006359905, 0.0004011344, 0.0003123115,
  0.001074921, 0.0009965914, 0.000949616, 0.0009052905, 0.0007076812, 
    0.0004398235, 0.0006716397, 0.0006833635, 0.0007061739, 0.000649713, 
    0.0006716747, 0.0006925944, 0.000664248, 0.0006261519, 0.0004388681,
  0.001036437, 0.0009981121, 0.0009270424, 0.0008431557, 0.0007757313, 
    0.0006916833, 0.0003898216, 0.0005880829, 0.0006791412, 0.0006300923, 
    0.0006466847, 0.0006645711, 0.000654576, 0.0006103413, 0.0004900293,
  0.0009850053, 0.0009462467, 0.0008758054, 0.0008179686, 0.0007526397, 
    0.0007389758, 0.0007264304, 0.0004323155, 0.0004583884, 0.0005554088, 
    0.0005839331, 0.0006172941, 0.0006310287, 0.0006179803, 0.0005850727,
  0.00100065, 0.0009398441, 0.0008752222, 0.0008142266, 0.0007571048, 
    0.0007260385, 0.0007007107, 0.0006955507, 0.0005986123, 0.0005738524, 
    0.0005592173, 0.0005869356, 0.0006149106, 0.0006228877, 0.0006070727,
  0.001049451, 0.0009741975, 0.0008805915, 0.0008200234, 0.000767327, 
    0.0007287167, 0.0007060217, 0.0006818941, 0.0006670841, 0.0007052703, 
    0.0006286543, 0.0005583372, 0.0005866491, 0.0006084851, 0.000592471,
  0.001070552, 0.001012136, 0.0009234792, 0.0008583146, 0.0008035842, 
    0.000737306, 0.0006885672, 0.0006683614, 0.0006711602, 0.000704921, 
    0.0006311021, 0.0005381237, 0.0005557536, 0.0005766152, 0.0005672105,
  0.001083633, 0.001032597, 0.0009645977, 0.0009015722, 0.0008255244, 
    0.0007754309, 0.000734996, 0.0007179205, 0.0007071889, 0.0006815303, 
    0.0006291486, 0.0005264693, 0.0005363925, 0.0005512457, 0.0005467192,
  0.001096405, 0.001044034, 0.0009823715, 0.0009309803, 0.0008686552, 
    0.000819184, 0.0007656894, 0.0007355547, 0.0006617467, 0.0005681547, 
    0.0005667752, 0.0005314429, 0.0005299909, 0.0005417115, 0.0005458943,
  0.00135655, 0.000957029, 0.0009171431, 0.0007683452, 0.0007847981, 
    0.0008719563, 0.0008990131, 0.0008399659, 0.0007519785, 0.0005911266, 
    0.0005688903, 0.0005197859, 0.0004917724, 0.0005261312, 0.000397647,
  0.00105266, 0.0009244414, 0.0008820223, 0.0008166908, 0.0008227486, 
    0.0008938395, 0.0008435775, 0.0007689197, 0.0007478251, 0.0007469565, 
    0.0006169259, 0.0006135405, 0.0006456155, 0.0004667959, 0.0003591249,
  0.001022252, 0.0009121695, 0.0008965994, 0.0008758614, 0.0007884059, 
    0.0005282015, 0.0008091156, 0.0007307418, 0.0008211561, 0.0007840539, 
    0.0007080858, 0.000688506, 0.0007019042, 0.0007336077, 0.0005690817,
  0.001037595, 0.000917552, 0.0009029151, 0.0009244372, 0.0009551837, 
    0.0008529504, 0.0004783327, 0.0007189242, 0.000844559, 0.0007809772, 
    0.0007529865, 0.000746544, 0.0007570798, 0.0007377694, 0.0006500371,
  0.001061363, 0.0009329103, 0.0009097412, 0.0009228921, 0.000979447, 
    0.0009935297, 0.0009780178, 0.0005340397, 0.0005798342, 0.0007495183, 
    0.000801663, 0.0008105797, 0.0007985095, 0.0007743195, 0.0007421008,
  0.001092793, 0.000962796, 0.0009194835, 0.0009393317, 0.000981658, 
    0.001031706, 0.001059151, 0.001062984, 0.0009285291, 0.000889072, 
    0.0008250752, 0.0008427274, 0.0008258965, 0.0008209722, 0.0007943487,
  0.001142343, 0.001037194, 0.0009523911, 0.0009400369, 0.0009724433, 
    0.001024681, 0.001104523, 0.001156345, 0.00117752, 0.001154777, 
    0.0009591159, 0.0008804561, 0.0008590887, 0.0008834685, 0.0008635087,
  0.001166665, 0.001084921, 0.001017527, 0.0009777739, 0.00098604, 
    0.00101646, 0.001080766, 0.001176205, 0.00124537, 0.001251715, 
    0.001027212, 0.0009111268, 0.0009123381, 0.0009668338, 0.0008624067,
  0.00117681, 0.001115904, 0.001056893, 0.001002287, 0.0009845035, 
    0.001015987, 0.00106609, 0.001157736, 0.001246354, 0.001265802, 
    0.001057588, 0.0009349418, 0.0009632639, 0.0009499122, 0.0007702274,
  0.001193253, 0.001137045, 0.001062313, 0.001022832, 0.001004515, 
    0.001004244, 0.001034052, 0.001115969, 0.001112094, 0.001008649, 
    0.0009774503, 0.0009476212, 0.0009797541, 0.0008969891, 0.0008073791,
  0.001627185, 0.001509548, 0.001357412, 0.001181064, 0.001317018, 
    0.001360065, 0.001155056, 0.0008835946, 0.0007219403, 0.0003829865, 
    0.0004272309, 0.0003292248, 0.0002595325, 0.0003015403, 0.0001728117,
  0.001619205, 0.00134769, 0.001134195, 0.001035277, 0.000908931, 
    0.001100016, 0.001314754, 0.001084897, 0.0008672302, 0.0006225342, 
    0.0004528249, 0.0004215558, 0.0004344355, 0.0002632265, 0.0001726813,
  0.001543007, 0.001241649, 0.001038922, 0.00100364, 0.001034016, 
    0.0006833803, 0.00130439, 0.001133973, 0.000982509, 0.0007315299, 
    0.0005624832, 0.0004503138, 0.0004284699, 0.000503736, 0.0003884511,
  0.001403165, 0.001116892, 0.001022387, 0.001012057, 0.00102764, 
    0.001341936, 0.0007136638, 0.001069162, 0.0009523394, 0.0006865243, 
    0.0005382542, 0.0004492979, 0.0004391255, 0.0004859319, 0.0004871878,
  0.001259651, 0.001033163, 0.001014809, 0.001016426, 0.001020862, 
    0.001243402, 0.001435786, 0.0006782218, 0.0005928428, 0.0005330672, 
    0.0005076898, 0.0004604468, 0.000481087, 0.0005415746, 0.0005476545,
  0.001170587, 0.001023674, 0.001020593, 0.001016725, 0.001017304, 
    0.001225119, 0.001474348, 0.001267614, 0.0008449564, 0.000723758, 
    0.000517319, 0.0005026202, 0.0005421782, 0.0005924528, 0.0005231393,
  0.001108071, 0.001009802, 0.001025058, 0.001023635, 0.001069359, 
    0.001267876, 0.001416581, 0.001269477, 0.001146613, 0.001043686, 
    0.000680681, 0.0005857383, 0.0006191225, 0.0006142892, 0.0005862893,
  0.001047952, 0.001011261, 0.001055091, 0.001086339, 0.001177726, 
    0.001345669, 0.001377834, 0.001321993, 0.001225931, 0.001125887, 
    0.0007595569, 0.0006781573, 0.0006688548, 0.0006475661, 0.0006368958,
  0.001017296, 0.001026587, 0.001121003, 0.001198748, 0.001313804, 
    0.001407519, 0.001367448, 0.001349563, 0.001296851, 0.001184901, 
    0.0008603281, 0.0007526244, 0.0007148192, 0.0007080482, 0.0006962098,
  0.0009922312, 0.001070923, 0.001206234, 0.001319489, 0.001392032, 
    0.001417328, 0.001398169, 0.001380107, 0.001271977, 0.0009811533, 
    0.0008374979, 0.0007975359, 0.0007816156, 0.000742277, 0.0007940147,
  0.001244931, 0.001500216, 0.001518027, 0.001651438, 0.001625377, 
    0.001482349, 0.001083796, 0.0005888687, 0.0004478158, 0.0002904466, 
    0.0002569427, 0.0002614844, 0.0002300165, 0.0002828164, 9.693115e-05,
  0.001584934, 0.001652695, 0.001691091, 0.001635522, 0.001549146, 
    0.001266933, 0.0008635756, 0.0006096173, 0.0004933051, 0.0003930131, 
    0.0002985082, 0.0003892836, 0.0004560337, 0.0002105278, 8.913482e-05,
  0.001648976, 0.001702621, 0.001676034, 0.001637538, 0.001684307, 
    0.0007899839, 0.000874568, 0.0006835842, 0.0005567619, 0.0004712873, 
    0.0004627351, 0.0004345903, 0.0004524546, 0.0005335872, 0.000291738,
  0.001720609, 0.001707252, 0.001646413, 0.001639671, 0.001775707, 
    0.00139257, 0.0006251337, 0.0006531405, 0.0005855231, 0.0005366409, 
    0.0004771214, 0.0004510333, 0.0004884864, 0.000519788, 0.0003997945,
  0.001762109, 0.001710972, 0.00161092, 0.001591451, 0.001693794, 
    0.001697783, 0.001229759, 0.0005217785, 0.0004206049, 0.0004834959, 
    0.0004714851, 0.000477387, 0.0005233486, 0.0005751593, 0.0006096233,
  0.001765804, 0.001701539, 0.001576418, 0.001536617, 0.001578487, 
    0.001684929, 0.001532269, 0.001232063, 0.0007983778, 0.00065925, 
    0.000499821, 0.0005090066, 0.0005520935, 0.0006098123, 0.0006266892,
  0.001803496, 0.001676399, 0.001534792, 0.001493325, 0.001488797, 
    0.001624539, 0.001570885, 0.001323628, 0.001168588, 0.001017788, 
    0.0006608014, 0.0005387455, 0.0005938174, 0.0006497502, 0.0006695391,
  0.001819151, 0.001646176, 0.0014741, 0.001451923, 0.001467006, 0.001626738, 
    0.001548359, 0.001329417, 0.001240335, 0.001076151, 0.0006604787, 
    0.0005730179, 0.0006407145, 0.0006896465, 0.0007292586,
  0.001788189, 0.001579517, 0.001432194, 0.001430467, 0.001530756, 
    0.001678904, 0.00149353, 0.001309232, 0.001239069, 0.001096383, 
    0.0007117121, 0.0006164405, 0.0006933659, 0.0007289145, 0.0007595762,
  0.001690051, 0.001488864, 0.001415162, 0.001478484, 0.001611821, 
    0.001688063, 0.001448498, 0.001311227, 0.001169003, 0.0008710331, 
    0.0006851083, 0.0006731757, 0.0007302076, 0.0007467864, 0.0009168799,
  0.00088528, 0.001201036, 0.001079171, 0.00125862, 0.001014239, 0.001034869, 
    0.0009659665, 0.0006281153, 0.0004475539, 0.0002527351, 0.0002212355, 
    0.000376318, 0.000362545, 0.0003735471, 0.0001366704,
  0.001296363, 0.001383019, 0.001416203, 0.00146578, 0.001206658, 
    0.001146873, 0.000894357, 0.0005875426, 0.0004556496, 0.0003573807, 
    0.0002785535, 0.000474667, 0.000610749, 0.0003192766, 0.000151656,
  0.001364552, 0.001452958, 0.001496675, 0.001574523, 0.001456165, 
    0.0009470491, 0.0008003141, 0.0005728637, 0.0004803931, 0.0004580799, 
    0.0004601229, 0.000506894, 0.0006509511, 0.0006714613, 0.000356046,
  0.001441461, 0.001504462, 0.001556391, 0.001672607, 0.001727208, 
    0.001317889, 0.000594279, 0.0005274338, 0.0004936859, 0.0004924979, 
    0.0004695536, 0.00052552, 0.0006918043, 0.0006787174, 0.0004769487,
  0.001558232, 0.00156873, 0.001619871, 0.001735362, 0.001832251, 
    0.001683983, 0.001125137, 0.0004301983, 0.0003278341, 0.0004281811, 
    0.0004725989, 0.0005441894, 0.0007414487, 0.0007703389, 0.0007549651,
  0.001662471, 0.001665466, 0.001681468, 0.001796095, 0.001886602, 
    0.00177396, 0.001537758, 0.001216602, 0.0008166729, 0.0006324744, 
    0.0005109624, 0.0006097996, 0.0007381557, 0.0007931156, 0.0008247024,
  0.001735576, 0.001728542, 0.001744724, 0.001861559, 0.001903245, 
    0.00177547, 0.001584364, 0.001368414, 0.001118225, 0.0009636085, 
    0.0007170626, 0.0006543247, 0.000766579, 0.0008115225, 0.0008470005,
  0.001842155, 0.001794712, 0.001820874, 0.001917504, 0.001934704, 
    0.001770031, 0.001569013, 0.001341478, 0.001213365, 0.001072069, 
    0.0007431243, 0.0006946061, 0.0008016748, 0.0008381997, 0.0009229468,
  0.001903303, 0.001878514, 0.001899447, 0.001982551, 0.001950409, 
    0.001769725, 0.001554188, 0.001342279, 0.001222701, 0.00110814, 
    0.0007905091, 0.0007411053, 0.0007933188, 0.0008469958, 0.0009073482,
  0.001927466, 0.001914913, 0.001925961, 0.002005461, 0.001962456, 
    0.001789356, 0.001523918, 0.001323816, 0.001178437, 0.0009667049, 
    0.0007902536, 0.0007792472, 0.0008167436, 0.0008544762, 0.0009759422,
  0.000772438, 0.001163808, 0.0010059, 0.001219889, 0.0006638478, 
    0.0005627173, 0.0006315805, 0.0005536226, 0.0005698404, 0.0004648798, 
    0.0004917078, 0.0006475924, 0.000390827, 0.0002845594, 0.0001847626,
  0.00133039, 0.001358878, 0.001353296, 0.001324019, 0.0007065058, 
    0.0006569041, 0.0006965324, 0.0005668725, 0.0005829588, 0.0006339918, 
    0.0006075518, 0.0007922468, 0.0007004802, 0.0002596571, 0.0001687422,
  0.001467045, 0.001414186, 0.001396409, 0.001387421, 0.0009642097, 
    0.0006303654, 0.0006942466, 0.000579554, 0.0005710205, 0.0006404648, 
    0.0007308832, 0.0008222234, 0.0007878378, 0.0006394278, 0.0003634478,
  0.001588381, 0.001502888, 0.001453981, 0.001459778, 0.00140206, 
    0.001051989, 0.0006071811, 0.0005456786, 0.000593778, 0.0006425751, 
    0.0007123311, 0.0008540399, 0.0008345716, 0.0006993202, 0.000474708,
  0.001676755, 0.001584322, 0.001518958, 0.00153641, 0.001477903, 
    0.001331103, 0.001025055, 0.0003863266, 0.0003047553, 0.0004963411, 
    0.0006873384, 0.0008411941, 0.0008748884, 0.00080411, 0.0007477585,
  0.00174588, 0.001662803, 0.001574419, 0.001575332, 0.001535129, 0.00145588, 
    0.001288368, 0.001224113, 0.0008843751, 0.0008195325, 0.0006759848, 
    0.0008405477, 0.0008459722, 0.0008404177, 0.0007752199,
  0.001857922, 0.001750271, 0.001636379, 0.001625334, 0.001595527, 
    0.001502593, 0.001352495, 0.001204588, 0.001052843, 0.001021997, 
    0.0008472624, 0.0008264109, 0.0008687042, 0.0008616764, 0.0008023459,
  0.001958499, 0.001826381, 0.001703547, 0.001656095, 0.001649977, 
    0.001531689, 0.001452415, 0.001382723, 0.001226002, 0.001084211, 
    0.0008751647, 0.0008399083, 0.0008875154, 0.0009009796, 0.000876707,
  0.002021183, 0.001890926, 0.00178963, 0.001697908, 0.00167827, 0.001593973, 
    0.001539589, 0.001564428, 0.001370621, 0.00113467, 0.0009251445, 
    0.0008383736, 0.0008766534, 0.00092754, 0.0009199308,
  0.002033893, 0.001893284, 0.001803636, 0.001733431, 0.001705684, 
    0.001635366, 0.001647215, 0.001738247, 0.001509409, 0.001231084, 
    0.0009567636, 0.0008677692, 0.000840957, 0.0009351274, 0.0009560644,
  0.0008458176, 0.001190368, 0.0008845752, 0.001084112, 0.0006570603, 
    0.0005646124, 0.0006926673, 0.0007068245, 0.0006670813, 0.0004240672, 
    0.0003271729, 0.0003047152, 0.0002451753, 0.000259932, 0.0001568898,
  0.001496093, 0.001510897, 0.001399384, 0.001277391, 0.0006873483, 
    0.0005112923, 0.000702277, 0.0007348695, 0.0007319978, 0.0006415503, 
    0.0004539293, 0.0004806627, 0.000463364, 0.0002150851, 0.0001551139,
  0.001680422, 0.001684084, 0.001515253, 0.001398753, 0.0009546456, 
    0.0004645502, 0.000714039, 0.0007344856, 0.0007861954, 0.000744412, 
    0.0006692006, 0.0006173963, 0.000581963, 0.0005312226, 0.0003779555,
  0.001756507, 0.001748445, 0.001622341, 0.00150387, 0.001328078, 
    0.001041593, 0.0003740854, 0.0007271524, 0.0008317417, 0.0008160004, 
    0.000748889, 0.0006856118, 0.0006400816, 0.0005952384, 0.0004971575,
  0.001724403, 0.001799866, 0.001673218, 0.001536297, 0.001412271, 
    0.001253327, 0.001062977, 0.0003586949, 0.0004535542, 0.0007161964, 
    0.0008431548, 0.0007507892, 0.0007203926, 0.0006607264, 0.0006330814,
  0.001756601, 0.001826778, 0.001701048, 0.001573465, 0.001473585, 
    0.001294467, 0.001117284, 0.00111505, 0.0009746728, 0.0008537669, 
    0.0008141619, 0.0007889356, 0.000736739, 0.0007158141, 0.0006783006,
  0.001839038, 0.001846468, 0.001727474, 0.00162604, 0.001505711, 
    0.001366977, 0.001152952, 0.001121571, 0.001153011, 0.001043601, 
    0.0008733693, 0.0008198628, 0.0007661768, 0.0007316038, 0.0007075011,
  0.001937845, 0.001903498, 0.001797273, 0.00168416, 0.001550114, 
    0.001467586, 0.00123796, 0.001159139, 0.001213907, 0.001135179, 
    0.0008790755, 0.0008391079, 0.0008001305, 0.0007523518, 0.0007066864,
  0.002128603, 0.001998359, 0.001866944, 0.001771548, 0.00163725, 
    0.001559009, 0.001366663, 0.001207929, 0.001248538, 0.001188893, 
    0.0008963486, 0.0008594687, 0.0008102524, 0.0007735668, 0.0007376147,
  0.00240006, 0.002104545, 0.001973284, 0.00186841, 0.001720868, 0.001640318, 
    0.001467237, 0.001302073, 0.001296729, 0.001149365, 0.0008986455, 
    0.0008806097, 0.0008392516, 0.0008358302, 0.0008460688,
  0.0009499397, 0.001149502, 0.0007682691, 0.0009003985, 0.0005971981, 
    0.000568375, 0.00050288, 0.0004347326, 0.0004046461, 0.0002776233, 
    0.0002694313, 0.0003518319, 0.0002644564, 0.0002780122, 0.0001469581,
  0.001342832, 0.001474158, 0.001364417, 0.00119469, 0.0006357197, 
    0.0005701555, 0.0005671176, 0.0004952668, 0.0004546067, 0.0004283974, 
    0.0003414695, 0.0004923914, 0.0005315549, 0.0002249122, 0.0001758391,
  0.001423813, 0.001612327, 0.001540148, 0.001368562, 0.0008749946, 
    0.0004309369, 0.0006135506, 0.0005655137, 0.0005074158, 0.0004902874, 
    0.0004987904, 0.000530626, 0.000566921, 0.0005664405, 0.0004686276,
  0.001488455, 0.001662728, 0.001623156, 0.001500361, 0.001250613, 
    0.0009569713, 0.0004500638, 0.0006042387, 0.000532969, 0.0004999242, 
    0.0004968515, 0.0005274737, 0.000598839, 0.0006075615, 0.0005892752,
  0.00159126, 0.001716183, 0.001638218, 0.001518766, 0.00137599, 0.001248318, 
    0.001010921, 0.0004574817, 0.0003843172, 0.0004663018, 0.0005309322, 
    0.0005534811, 0.0006127105, 0.0006598222, 0.0006762806,
  0.001679538, 0.001758969, 0.001666014, 0.001550281, 0.001415143, 
    0.001316036, 0.001245789, 0.001186371, 0.0008895199, 0.0007372125, 
    0.0006253528, 0.000607106, 0.0006345148, 0.0006927265, 0.0007001914,
  0.001762336, 0.001824967, 0.001684023, 0.001551474, 0.001418927, 
    0.001337155, 0.001294001, 0.001299163, 0.001194505, 0.0009966001, 
    0.0007740417, 0.0006804593, 0.0006741179, 0.0007082425, 0.0007342691,
  0.001853498, 0.001842372, 0.001702707, 0.001551111, 0.001408467, 
    0.001363692, 0.001323492, 0.001366799, 0.00132725, 0.00120011, 
    0.0008475368, 0.0007592109, 0.0007294266, 0.0007415477, 0.0007675747,
  0.001802848, 0.001869602, 0.001728557, 0.001585005, 0.001447891, 
    0.001399313, 0.00134403, 0.001365151, 0.001402971, 0.001252707, 
    0.0009403671, 0.0008329428, 0.0007623697, 0.0007690038, 0.0007539341,
  0.001868906, 0.001863841, 0.001764924, 0.001634837, 0.001485711, 
    0.001445699, 0.001384234, 0.001382799, 0.001437627, 0.001259611, 
    0.0009653283, 0.0008624629, 0.0007916858, 0.0007723793, 0.0007599458,
  0.0006798884, 0.0009273534, 0.0005796482, 0.0006608103, 0.0004814486, 
    0.0004714799, 0.0005278075, 0.0005502158, 0.0005886609, 0.00045812, 
    0.0004042562, 0.0005589795, 0.0004087429, 0.0003560864, 0.0001946153,
  0.001176487, 0.001217431, 0.001106654, 0.00098748, 0.0004817574, 
    0.0004257961, 0.000531052, 0.0005457469, 0.0005764399, 0.0006147923, 
    0.0004663036, 0.0007179814, 0.0007537344, 0.0003987499, 0.0003305572,
  0.00138231, 0.001364927, 0.001269183, 0.001169216, 0.0007256914, 
    0.000329046, 0.000513851, 0.0005435139, 0.000555283, 0.0005686608, 
    0.0006163557, 0.0007253342, 0.0008122339, 0.0008388328, 0.0006753516,
  0.001476959, 0.001448341, 0.001373286, 0.001281204, 0.001096852, 
    0.0008199436, 0.0003577206, 0.0004773551, 0.0005557741, 0.000553521, 
    0.0005882949, 0.0006964356, 0.0008280664, 0.0009100551, 0.0008928301,
  0.001586157, 0.001521092, 0.001416144, 0.001337198, 0.001202348, 
    0.00111714, 0.0009070458, 0.0002796284, 0.0003022251, 0.0004461132, 
    0.0006012633, 0.0006826049, 0.0008393758, 0.0009476088, 0.001038018,
  0.0016845, 0.001584252, 0.001488847, 0.001426884, 0.001287733, 0.001214396, 
    0.001114098, 0.001043793, 0.0008507161, 0.0007033524, 0.0005808385, 
    0.000685019, 0.0008334256, 0.0009559054, 0.001054576,
  0.001782312, 0.001677385, 0.001535428, 0.001463733, 0.001377879, 
    0.001301077, 0.001213597, 0.001089582, 0.0009625062, 0.0008288816, 
    0.0006907607, 0.0007047806, 0.000842174, 0.000958983, 0.001076277,
  0.001884768, 0.001778794, 0.001622893, 0.001542567, 0.001431314, 
    0.001381897, 0.001327644, 0.001175244, 0.001110879, 0.001021823, 
    0.0007425516, 0.0007307242, 0.0008326205, 0.0009313844, 0.001029254,
  0.001969611, 0.001953857, 0.001751087, 0.001625228, 0.001518527, 
    0.001469287, 0.001410406, 0.001342807, 0.001226469, 0.001122528, 
    0.0008596066, 0.0007590873, 0.0008196975, 0.000912409, 0.0009862127,
  0.002047504, 0.00199633, 0.001895577, 0.001766649, 0.001590899, 
    0.001525608, 0.001485578, 0.001443221, 0.001365813, 0.001296134, 
    0.0009303325, 0.0007913189, 0.0008148858, 0.0009087075, 0.0009863926,
  0.0005373147, 0.0007805214, 0.0005494839, 0.000688454, 0.0006035151, 
    0.0005343809, 0.000637004, 0.0006768154, 0.000782443, 0.0006551942, 
    0.0006120364, 0.0007427997, 0.0004999139, 0.0004425556, 0.0002340348,
  0.001027295, 0.001005504, 0.0009166581, 0.0008526498, 0.0005107899, 
    0.0004301495, 0.0006526909, 0.0006751962, 0.0007709893, 0.0009061305, 
    0.0007893663, 0.0009951666, 0.000932599, 0.0004062481, 0.0003589842,
  0.001194022, 0.001099992, 0.001016954, 0.0009169065, 0.000756191, 
    0.0003515301, 0.0005720931, 0.0006900679, 0.0007957664, 0.0009209301, 
    0.0010626, 0.001146029, 0.001105798, 0.001030551, 0.0008822888,
  0.001263715, 0.001164421, 0.001088056, 0.001011363, 0.0009564605, 
    0.0008251561, 0.0003314013, 0.0005498652, 0.0007373804, 0.0008821575, 
    0.001074097, 0.001199308, 0.001253918, 0.001227383, 0.001170399,
  0.001384472, 0.00128414, 0.001205278, 0.0011191, 0.00106159, 0.0009778483, 
    0.00100376, 0.0003562877, 0.0004935193, 0.0007496522, 0.00105561, 
    0.001203255, 0.001278205, 0.001284672, 0.001289382,
  0.001573931, 0.00149022, 0.001390371, 0.001291875, 0.001173697, 
    0.001082886, 0.001017811, 0.001078487, 0.0008554214, 0.0008177335, 
    0.0009578709, 0.00114646, 0.001208172, 0.001255337, 0.001285275,
  0.001847709, 0.001745894, 0.001634079, 0.001521914, 0.001432419, 
    0.001259308, 0.001100925, 0.001113743, 0.0009630601, 0.0008648491, 
    0.0009729539, 0.001030203, 0.001079856, 0.001157657, 0.001176759,
  0.002167573, 0.002016585, 0.001866266, 0.001725203, 0.001628359, 
    0.001502276, 0.001414135, 0.001286658, 0.001152089, 0.0009404718, 
    0.0009455087, 0.0009860464, 0.001018292, 0.00106275, 0.001061653,
  0.002766941, 0.002561068, 0.002344088, 0.002050011, 0.001799255, 
    0.001653079, 0.001551699, 0.001477036, 0.001362495, 0.001017129, 
    0.0009170455, 0.000954263, 0.001006527, 0.001003009, 0.001081152,
  0.003370462, 0.003073762, 0.002814954, 0.002461525, 0.002052115, 
    0.001787674, 0.00163222, 0.001580021, 0.001502705, 0.001090751, 
    0.0009016439, 0.0009133887, 0.0009744045, 0.0009527082, 0.000928279,
  0.0005341409, 0.0008826249, 0.0009600315, 0.001047156, 0.0007562609, 
    0.000584148, 0.0008892031, 0.001049999, 0.001167649, 0.0008060374, 
    0.0007696306, 0.0009845537, 0.0008126931, 0.0007442924, 0.0005443592,
  0.001040602, 0.001075951, 0.0009898562, 0.0009579254, 0.0006458763, 
    0.0004938116, 0.0008551904, 0.001015583, 0.001103399, 0.001110524, 
    0.0009045989, 0.00116826, 0.001149286, 0.0006721864, 0.0006703583,
  0.00121307, 0.001147719, 0.001091314, 0.001044464, 0.00117624, 
    0.0004658278, 0.0006519388, 0.001005674, 0.001107991, 0.001102994, 
    0.001084485, 0.001137539, 0.001129116, 0.001069996, 0.001038198,
  0.001355185, 0.001272149, 0.001253757, 0.001222565, 0.001185567, 
    0.001282745, 0.000334508, 0.0006546882, 0.0009608683, 0.001023664, 
    0.001028946, 0.001054963, 0.001086033, 0.001063013, 0.001050826,
  0.001524473, 0.001497808, 0.001458212, 0.001387928, 0.001265825, 
    0.001212428, 0.001366718, 0.000367339, 0.0006267116, 0.0007608711, 
    0.0009521634, 0.0009843967, 0.001014404, 0.001011328, 0.0009952179,
  0.001735846, 0.001725, 0.001662737, 0.001593734, 0.001512472, 0.001266592, 
    0.001425831, 0.001206863, 0.0008933156, 0.0008955363, 0.0009561845, 
    0.0009532101, 0.0009628076, 0.0009675283, 0.0009682935,
  0.002045075, 0.001932436, 0.001862278, 0.001777547, 0.001738863, 
    0.001592762, 0.001503929, 0.00119044, 0.0009233949, 0.0008149219, 
    0.001059868, 0.000981533, 0.0009577794, 0.0009486928, 0.0009455047,
  0.002888527, 0.002589704, 0.002339725, 0.002073884, 0.001902553, 
    0.00176095, 0.001644253, 0.00154557, 0.001174547, 0.0008917419, 
    0.0009982439, 0.0009940504, 0.0009661579, 0.0009524039, 0.0009235491,
  0.002989678, 0.002987709, 0.002969476, 0.002798998, 0.002446956, 
    0.002086795, 0.001808255, 0.001745381, 0.00160857, 0.001083056, 
    0.001033956, 0.0009709422, 0.0009494151, 0.0009543331, 0.0009152948,
  0.002413466, 0.002476096, 0.002556591, 0.002960916, 0.00289151, 0.00256091, 
    0.00209713, 0.001861234, 0.001759731, 0.001230514, 0.001099309, 
    0.0009974861, 0.0009327075, 0.0009302826, 0.0008835403,
  0.000552893, 0.0008929609, 0.0009882366, 0.001260897, 0.001088799, 
    0.0006892661, 0.0008799786, 0.0009201678, 0.000943662, 0.0006675241, 
    0.000623949, 0.0008122245, 0.0007855237, 0.000775423, 0.0005889317,
  0.001104261, 0.001247855, 0.001326396, 0.00132429, 0.0009368055, 
    0.0005478994, 0.0007878274, 0.0008937292, 0.0008923783, 0.0008558935, 
    0.0007508846, 0.0008794786, 0.0009293854, 0.000703922, 0.0006539749,
  0.00128977, 0.001258296, 0.001239815, 0.001366237, 0.00152618, 
    0.0005731707, 0.0006570735, 0.0008422083, 0.0008530967, 0.0008403381, 
    0.000812908, 0.0008768275, 0.0009082113, 0.001000202, 0.0009943329,
  0.001365829, 0.001331817, 0.001278924, 0.001369915, 0.00145947, 
    0.001603981, 0.0005563722, 0.00061446, 0.0007305252, 0.0008060838, 
    0.0007800685, 0.0008539949, 0.0008914869, 0.0009640569, 0.001054368,
  0.00150186, 0.001454037, 0.001417143, 0.001442067, 0.001486795, 
    0.001723685, 0.00165601, 0.000374269, 0.0004001498, 0.0007283142, 
    0.0008174353, 0.0008468534, 0.0008667379, 0.0009219896, 0.001056243,
  0.001631551, 0.001597764, 0.0015486, 0.001528376, 0.001584384, 0.001627145, 
    0.001767067, 0.001675269, 0.00107615, 0.0009142941, 0.0008415225, 
    0.0009039906, 0.0008648193, 0.000872373, 0.0009711111,
  0.001846651, 0.001746741, 0.001689313, 0.001628597, 0.001652272, 
    0.001671363, 0.001750827, 0.001635544, 0.001357218, 0.001064977, 
    0.001070352, 0.001038734, 0.0009333307, 0.0008568658, 0.0009155434,
  0.002201915, 0.001986342, 0.001871417, 0.001804298, 0.001773144, 
    0.001768922, 0.001833677, 0.001769201, 0.001685568, 0.001431528, 
    0.001293811, 0.001198343, 0.001039515, 0.0009004368, 0.0008854038,
  0.002394401, 0.00226598, 0.002208276, 0.002136066, 0.0020488, 0.001976997, 
    0.001990201, 0.001976351, 0.001903861, 0.001815302, 0.001586839, 
    0.001381361, 0.001176397, 0.0009948596, 0.0009237388,
  0.002370987, 0.002291222, 0.002254694, 0.00230897, 0.002306225, 
    0.002317201, 0.002299361, 0.002301476, 0.002202974, 0.002048776, 
    0.001860846, 0.001585289, 0.001319788, 0.001102283, 0.0009940605,
  0.0006755121, 0.0008474457, 0.0007146689, 0.0007368508, 0.0007282908, 
    0.0006791523, 0.0007444739, 0.000720392, 0.0007642721, 0.0005719279, 
    0.000597754, 0.0007150251, 0.0007185221, 0.0007549985, 0.0005324639,
  0.001217584, 0.00133114, 0.001353839, 0.00122484, 0.0007395571, 
    0.0005881015, 0.0007312061, 0.0007829908, 0.0007713556, 0.0007045662, 
    0.000622788, 0.0008922705, 0.001015559, 0.0006633607, 0.0006205223,
  0.001406589, 0.001410181, 0.001433711, 0.001394995, 0.001291472, 
    0.0004760293, 0.0009073554, 0.0007851818, 0.0007767596, 0.0007278598, 
    0.0007847825, 0.001002138, 0.001101404, 0.001108407, 0.001020487,
  0.001421558, 0.001400608, 0.001430688, 0.001473772, 0.001503381, 
    0.001603098, 0.0008177204, 0.000769066, 0.0008854743, 0.0007979902, 
    0.0008216473, 0.001067279, 0.001138487, 0.001173758, 0.001087694,
  0.001408303, 0.00139127, 0.001350541, 0.001391966, 0.001502815, 0.00165702, 
    0.001787057, 0.001076275, 0.0008854249, 0.0009459851, 0.0009442134, 
    0.00119766, 0.001256358, 0.001258711, 0.001157919,
  0.001430536, 0.001409882, 0.001378882, 0.001382363, 0.001447495, 
    0.001482901, 0.001665601, 0.001998274, 0.001661808, 0.001411274, 
    0.001191822, 0.001383294, 0.00148565, 0.001424069, 0.001313887,
  0.001480456, 0.001453133, 0.001419892, 0.0014122, 0.001440885, 0.001491514, 
    0.001549642, 0.001680142, 0.002047418, 0.002005052, 0.001753208, 
    0.001749158, 0.001767343, 0.001652846, 0.001449171,
  0.001571106, 0.001532083, 0.001499469, 0.001484787, 0.00151539, 
    0.001577635, 0.00166841, 0.001745716, 0.001855526, 0.002109743, 
    0.002073617, 0.00202966, 0.001987494, 0.001834719, 0.001657312,
  0.001699813, 0.00167232, 0.001652212, 0.001652831, 0.00169244, 0.001748815, 
    0.00181815, 0.001890395, 0.001991543, 0.002105271, 0.002076475, 
    0.00207196, 0.002090856, 0.001962824, 0.001834271,
  0.001893193, 0.001808029, 0.001801415, 0.001833273, 0.001892647, 
    0.001963301, 0.002027125, 0.002119849, 0.002241175, 0.002143055, 
    0.002193006, 0.002110961, 0.002078997, 0.002020758, 0.001927831,
  0.0007152242, 0.0008318364, 0.0007638162, 0.000768077, 0.0006625067, 
    0.0005937974, 0.0006507834, 0.0006394563, 0.0006145029, 0.0005030361, 
    0.0005064808, 0.0006863811, 0.0007530211, 0.000934726, 0.0005782566,
  0.001162282, 0.001304111, 0.001308041, 0.001043943, 0.0006541855, 
    0.0005863697, 0.0006901795, 0.0006818559, 0.0006953478, 0.0007521355, 
    0.0006846727, 0.0009078538, 0.00123332, 0.001182003, 0.0006318286,
  0.001452836, 0.001534318, 0.001554312, 0.001393188, 0.0009059472, 
    0.0004818485, 0.0007574465, 0.0007563143, 0.0008719402, 0.0009974671, 
    0.00106104, 0.001312933, 0.001499479, 0.001589967, 0.000926148,
  0.001567465, 0.001638812, 0.00163147, 0.001535972, 0.001372576, 
    0.001092238, 0.0005287361, 0.000713298, 0.001277442, 0.001381364, 
    0.001348761, 0.001560515, 0.001753439, 0.001708115, 0.001072198,
  0.001603156, 0.001650623, 0.001642448, 0.00156528, 0.00146826, 0.001394933, 
    0.001367623, 0.000795011, 0.001049342, 0.001560173, 0.001673619, 
    0.001752669, 0.001880362, 0.001918858, 0.001279709,
  0.001640499, 0.001643406, 0.001599604, 0.00153851, 0.001483597, 
    0.001462336, 0.001448104, 0.001540226, 0.001508851, 0.001811892, 
    0.001760342, 0.001868297, 0.001952122, 0.002015541, 0.001586202,
  0.0016725, 0.001653704, 0.001604979, 0.001545453, 0.001521908, 0.001507511, 
    0.001514627, 0.001533778, 0.001724925, 0.002049942, 0.002002914, 
    0.001970698, 0.001978321, 0.002027512, 0.00176195,
  0.001669067, 0.001641816, 0.001597452, 0.001556685, 0.0015306, 0.001538252, 
    0.001547033, 0.001594135, 0.001704924, 0.001891246, 0.001866029, 
    0.001897239, 0.001969662, 0.002071979, 0.001978893,
  0.0016385, 0.001613835, 0.001578916, 0.00154789, 0.001527505, 0.001538938, 
    0.001579936, 0.001669915, 0.001755652, 0.001968544, 0.001931839, 
    0.001993196, 0.002019028, 0.002111709, 0.002200688,
  0.001577043, 0.001546877, 0.001538685, 0.001554168, 0.001572407, 
    0.001609553, 0.001671082, 0.001746873, 0.001944382, 0.0019266, 
    0.002081373, 0.002223962, 0.002272513, 0.002332616, 0.00238812,
  0.0006399217, 0.0007436967, 0.0006720006, 0.0007074457, 0.0006096797, 
    0.0005158479, 0.0005751852, 0.0006405133, 0.0008366935, 0.0009964192, 
    0.0009304913, 0.000911308, 0.000577361, 0.0003797749, 0.0002072982,
  0.001212562, 0.001250322, 0.001212675, 0.0008779019, 0.0005933613, 
    0.0004913741, 0.0006522388, 0.0006690617, 0.0009278533, 0.001243974, 
    0.00131382, 0.001371565, 0.001120669, 0.0005583861, 0.0003896057,
  0.001550528, 0.001509903, 0.001452224, 0.001303954, 0.0008521124, 
    0.0003978443, 0.000665337, 0.0007179885, 0.00103521, 0.001465134, 
    0.001696442, 0.001825414, 0.001609524, 0.0012815, 0.0008210012,
  0.001694216, 0.001629946, 0.001562512, 0.001503406, 0.001360213, 
    0.001063915, 0.0004733276, 0.0006757177, 0.001136875, 0.001697748, 
    0.001699669, 0.001802116, 0.001926178, 0.001642767, 0.001176294,
  0.001728136, 0.001661641, 0.001615873, 0.001592689, 0.001493573, 
    0.001398712, 0.001245145, 0.000520603, 0.0007356763, 0.001518421, 
    0.001733886, 0.001761356, 0.001873448, 0.001794476, 0.001499333,
  0.001747927, 0.001700606, 0.001665378, 0.001631599, 0.001583634, 
    0.001487135, 0.001402169, 0.001510815, 0.001242288, 0.001534973, 
    0.001713628, 0.001786427, 0.001799054, 0.001708836, 0.001791314,
  0.001785782, 0.001766114, 0.001728073, 0.001671967, 0.001590073, 
    0.001495953, 0.001460526, 0.001398789, 0.001346234, 0.001541825, 
    0.001839971, 0.001883263, 0.001745622, 0.001796509, 0.00195506,
  0.001793228, 0.001810102, 0.001814131, 0.001764478, 0.001661437, 
    0.001551032, 0.001510049, 0.001462653, 0.001389684, 0.001605127, 
    0.001763706, 0.001813625, 0.001869358, 0.001976732, 0.002115096,
  0.00179936, 0.001839361, 0.001862653, 0.00181951, 0.001746863, 0.001644525, 
    0.001546473, 0.001501706, 0.001479853, 0.001645314, 0.001588511, 
    0.001616553, 0.00195056, 0.002013252, 0.00216947,
  0.001804967, 0.001830861, 0.001829621, 0.001810204, 0.001771326, 
    0.001708287, 0.001631921, 0.001554876, 0.001569871, 0.001531968, 
    0.001772571, 0.001790676, 0.001791875, 0.002029203, 0.002202246,
  0.0005546997, 0.0006438819, 0.0005687734, 0.0006905457, 0.0006276005, 
    0.0005129021, 0.0007762783, 0.001018135, 0.001252765, 0.001243826, 
    0.00125186, 0.001450251, 0.00140048, 0.001222659, 0.0006667318,
  0.001077508, 0.001087011, 0.00108648, 0.0008024375, 0.0004941471, 
    0.0003988909, 0.0006993039, 0.000849886, 0.001128399, 0.001354674, 
    0.001327486, 0.001553943, 0.001682579, 0.00134884, 0.0008224295,
  0.001359686, 0.001340087, 0.001318234, 0.001223641, 0.000842914, 
    0.0002809544, 0.000627997, 0.0007396014, 0.00101136, 0.001333233, 
    0.001394806, 0.001542983, 0.001696993, 0.00154061, 0.001029769,
  0.001518312, 0.00146591, 0.001446389, 0.001408556, 0.001365549, 
    0.001190589, 0.0004497012, 0.0006766762, 0.0008755163, 0.001263477, 
    0.001350476, 0.001479164, 0.001658964, 0.001567368, 0.001132106,
  0.001596008, 0.0015498, 0.001499734, 0.001476685, 0.00145451, 0.001421796, 
    0.001418607, 0.0005866642, 0.0005048659, 0.0009783038, 0.00132427, 
    0.001408002, 0.00162087, 0.001605785, 0.001304505,
  0.001662869, 0.001644569, 0.001593091, 0.001559491, 0.001551103, 
    0.001517796, 0.001491101, 0.001577457, 0.00134732, 0.0012027, 
    0.001195421, 0.001430198, 0.001561503, 0.001617254, 0.00137821,
  0.001760017, 0.001744019, 0.001660342, 0.001606949, 0.001589101, 
    0.001580857, 0.001556474, 0.001564142, 0.001609548, 0.001534907, 
    0.001401651, 0.001428962, 0.00154877, 0.001656213, 0.001514172,
  0.001833746, 0.001758732, 0.001715945, 0.001690237, 0.001673387, 
    0.001666671, 0.00166148, 0.001636303, 0.001630707, 0.001677382, 
    0.001461319, 0.001418725, 0.00147637, 0.001606505, 0.00162753,
  0.001893629, 0.001875348, 0.001867759, 0.001857447, 0.001862801, 
    0.001864135, 0.001841903, 0.001818325, 0.001756637, 0.001740225, 
    0.001538153, 0.001433396, 0.0013849, 0.001397194, 0.001767821,
  0.00189059, 0.001956306, 0.002013876, 0.00205155, 0.002083672, 0.002117622, 
    0.002107689, 0.002072674, 0.002003253, 0.001772325, 0.001753278, 
    0.001581199, 0.001366842, 0.00132212, 0.001744313,
  0.0007241182, 0.0009032185, 0.000885118, 0.0009491201, 0.0007176324, 
    0.0005786545, 0.0007864104, 0.0008492902, 0.0008903458, 0.0005727883, 
    0.0005645187, 0.0005719436, 0.000259701, 0.0001440574, 8.19065e-05,
  0.001215434, 0.00118177, 0.00119123, 0.001013099, 0.0005383793, 
    0.0004769819, 0.0008191947, 0.0009546555, 0.0009949026, 0.0007990211, 
    0.000608502, 0.0006609882, 0.0003760233, 0.0001216634, 8.008149e-05,
  0.001327455, 0.001251052, 0.001190657, 0.001122814, 0.00096764, 
    0.0004069997, 0.0008184594, 0.00104674, 0.001142321, 0.0009812211, 
    0.0008674367, 0.0006841945, 0.0004265632, 0.0002747808, 0.0001684489,
  0.001405973, 0.0013454, 0.001305404, 0.001295012, 0.001313527, 0.001295781, 
    0.0008498309, 0.001120001, 0.001260284, 0.001075744, 0.0009242778, 
    0.0007748912, 0.0004679832, 0.0002964043, 0.0002333029,
  0.001480902, 0.001384801, 0.001327737, 0.001354692, 0.001428958, 
    0.001539308, 0.001575427, 0.001046569, 0.001124756, 0.001074435, 
    0.0009886094, 0.000830099, 0.0005806389, 0.0003588048, 0.0003164147,
  0.001500556, 0.001502338, 0.001495241, 0.001531269, 0.001619591, 
    0.00167521, 0.001721934, 0.001916439, 0.001747145, 0.001488174, 
    0.001012802, 0.0009333655, 0.0007152631, 0.0004361532, 0.0003739221,
  0.001585115, 0.001632098, 0.001662944, 0.001707396, 0.00176867, 
    0.001826991, 0.001861096, 0.001877925, 0.002009093, 0.001870518, 
    0.001353983, 0.001082057, 0.0009234918, 0.0005546029, 0.0004393814,
  0.001683079, 0.001685944, 0.001723017, 0.001775006, 0.001843165, 
    0.001893738, 0.001919581, 0.001894396, 0.001995322, 0.001996093, 
    0.001509255, 0.001237752, 0.001160859, 0.0007596762, 0.0005350077,
  0.00176689, 0.001757296, 0.001798232, 0.001848219, 0.00195022, 0.001973364, 
    0.002002429, 0.002096235, 0.002027673, 0.002069849, 0.00162487, 
    0.00138307, 0.001191263, 0.001068881, 0.0006670808,
  0.001888414, 0.001894016, 0.001959585, 0.00205647, 0.002093467, 
    0.002137283, 0.002273837, 0.002335529, 0.002370083, 0.001991491, 
    0.001911539, 0.001530083, 0.001273909, 0.001111755, 0.001158145,
  0.001011945, 0.001070649, 0.000900061, 0.001097145, 0.000978273, 
    0.0008341064, 0.001062182, 0.000929612, 0.0005320949, 0.000215528, 
    0.0001686452, 0.000196181, 0.0001625248, 0.0001944151, 0.0001696597,
  0.001118703, 0.001040105, 0.001119513, 0.001246139, 0.0009754961, 
    0.0008650382, 0.001250837, 0.00128711, 0.0007884277, 0.0004153641, 
    0.000258016, 0.0003062661, 0.000330714, 0.000183368, 0.0001826304,
  0.001184081, 0.001079991, 0.001055778, 0.001246713, 0.001468002, 
    0.0008529571, 0.001348443, 0.001518704, 0.001161882, 0.0006689625, 
    0.0004543115, 0.0003825845, 0.0003567094, 0.0003711366, 0.0003498574,
  0.001275005, 0.00117553, 0.001188951, 0.00138506, 0.001647404, 0.001863416, 
    0.001400426, 0.001549657, 0.00131492, 0.0008610422, 0.0005577827, 
    0.0004335799, 0.0003901842, 0.0003883474, 0.0004105546,
  0.001370085, 0.001309964, 0.001336675, 0.001532742, 0.001762114, 
    0.001972416, 0.002198869, 0.001540276, 0.001289247, 0.0009402534, 
    0.0006789364, 0.000523798, 0.0004232656, 0.0004274448, 0.0004520239,
  0.001483923, 0.001474753, 0.001495246, 0.00168535, 0.001845235, 0.00201331, 
    0.002106791, 0.002286825, 0.001686163, 0.001228366, 0.0007581012, 
    0.000608984, 0.0004962829, 0.000455825, 0.0004795869,
  0.001578284, 0.001586504, 0.001654015, 0.001738999, 0.001859031, 
    0.002035678, 0.002112809, 0.002069438, 0.002082617, 0.001568908, 
    0.001070801, 0.000765688, 0.0005828826, 0.0005112399, 0.0005214442,
  0.001681235, 0.001666268, 0.001696638, 0.001743512, 0.001891154, 
    0.002048455, 0.002090076, 0.002044824, 0.002148803, 0.001801384, 
    0.001206083, 0.0009024697, 0.0007288269, 0.00056999, 0.0005611127,
  0.001733423, 0.0017363, 0.001750985, 0.001798249, 0.001965513, 0.002032434, 
    0.002068631, 0.002153226, 0.001981073, 0.001985841, 0.00161863, 
    0.001285802, 0.0009926077, 0.0007077972, 0.0005921789,
  0.001783836, 0.001763607, 0.001779322, 0.001851615, 0.001964916, 
    0.001974782, 0.002094628, 0.002018015, 0.002007436, 0.001783119, 
    0.001840524, 0.001569021, 0.001245699, 0.0009175009, 0.0006752075,
  0.0006891138, 0.0009053152, 0.0009228467, 0.001148973, 0.001127763, 
    0.00115084, 0.001438358, 0.001423014, 0.001045001, 0.000871529, 
    0.0006844496, 0.0005937198, 0.000340051, 0.0003368688, 0.0002758084,
  0.001167, 0.001198509, 0.001297872, 0.001403518, 0.001098799, 0.001144961, 
    0.001524102, 0.001474195, 0.001231443, 0.001210722, 0.0008774535, 
    0.0008145621, 0.0005669123, 0.0003110611, 0.0002946844,
  0.001283128, 0.001259918, 0.001289319, 0.001348023, 0.001557069, 
    0.001194655, 0.001548743, 0.001518868, 0.001367108, 0.001217326, 
    0.001175581, 0.0009446606, 0.0006095088, 0.0005738156, 0.0005165777,
  0.001388078, 0.00136364, 0.001368269, 0.001438028, 0.001642602, 
    0.001916641, 0.001252117, 0.001415641, 0.001403864, 0.001323674, 
    0.001225082, 0.0009907987, 0.0006596657, 0.0006051211, 0.0005786285,
  0.001414535, 0.001426133, 0.001449454, 0.00153648, 0.001729385, 
    0.001853705, 0.002119693, 0.001551975, 0.001540363, 0.001302743, 
    0.001248281, 0.001010937, 0.0007269967, 0.0006369418, 0.0006451333,
  0.001419205, 0.001445715, 0.001496307, 0.001606587, 0.001751732, 
    0.001848792, 0.001946479, 0.002195363, 0.00185003, 0.001790744, 
    0.001399592, 0.001158239, 0.0008108285, 0.0006622463, 0.0006483495,
  0.001525165, 0.001537761, 0.001581834, 0.001662928, 0.001754125, 
    0.001827131, 0.001914349, 0.001979847, 0.002194604, 0.002003897, 
    0.001750783, 0.001296222, 0.0009588992, 0.0006782047, 0.0006592525,
  0.001622043, 0.001633731, 0.001644926, 0.001688099, 0.001750435, 
    0.001812569, 0.001881293, 0.001946454, 0.00214736, 0.001987186, 
    0.001720892, 0.001404346, 0.001098212, 0.0007497136, 0.0006495544,
  0.001706886, 0.001728236, 0.001745677, 0.001739178, 0.001771189, 
    0.001821802, 0.001869722, 0.002097195, 0.002059748, 0.001912389, 
    0.001650961, 0.001471064, 0.001241744, 0.0008969016, 0.0006326871,
  0.00179405, 0.00177456, 0.001767276, 0.001778896, 0.001802006, 0.00187317, 
    0.00211003, 0.002152956, 0.00215794, 0.001713887, 0.001594709, 
    0.001505308, 0.001361685, 0.001179339, 0.0006925558,
  0.000728547, 0.0008389141, 0.000802741, 0.0008535275, 0.0008588271, 
    0.0008752742, 0.0009984776, 0.001106636, 0.001154936, 0.001116903, 
    0.001047013, 0.001017584, 0.0008721931, 0.0006121976, 0.0002900136,
  0.001116366, 0.001150287, 0.001200538, 0.001118788, 0.0008724961, 
    0.0009117621, 0.001162086, 0.001244093, 0.001301431, 0.0012832, 
    0.001176197, 0.001230998, 0.001137654, 0.0005714473, 0.0002376136,
  0.001312441, 0.00134687, 0.001403043, 0.001394891, 0.001400566, 
    0.0009298103, 0.001299199, 0.001387226, 0.0014125, 0.001384244, 
    0.001394528, 0.001376385, 0.001226173, 0.0008873023, 0.0003446112,
  0.001321249, 0.001401057, 0.00146473, 0.001512083, 0.001539555, 
    0.001605565, 0.001002569, 0.001313777, 0.001464233, 0.001473395, 
    0.001469263, 0.001463591, 0.001330688, 0.0009449971, 0.0004005529,
  0.001389205, 0.001480517, 0.001522401, 0.00157069, 0.001640705, 
    0.001695211, 0.001807211, 0.001321521, 0.001406153, 0.001379345, 
    0.001523979, 0.001498216, 0.00132436, 0.0009915003, 0.0005099634,
  0.001503768, 0.001564141, 0.001622208, 0.001698762, 0.001771902, 
    0.001831229, 0.001875574, 0.001966004, 0.001779384, 0.001613056, 
    0.001549704, 0.001594511, 0.001403314, 0.001040868, 0.0005861561,
  0.001835385, 0.001881036, 0.001928149, 0.001969447, 0.002025402, 
    0.002080848, 0.002142184, 0.002152846, 0.002167171, 0.0020616, 
    0.001903404, 0.001776811, 0.001502109, 0.001031725, 0.0005960962,
  0.002269211, 0.002287496, 0.002308153, 0.002341062, 0.002367453, 
    0.002402682, 0.00238511, 0.002312532, 0.002258292, 0.002176277, 
    0.002004016, 0.001854323, 0.001592517, 0.001026506, 0.0005701969,
  0.002573137, 0.002552042, 0.002537875, 0.002568557, 0.00260155, 
    0.002596208, 0.002452173, 0.002267361, 0.002217629, 0.002190038, 
    0.002091617, 0.00201002, 0.001658197, 0.0009972638, 0.000545404,
  0.002650793, 0.002676548, 0.002703668, 0.002744016, 0.002733956, 
    0.00263714, 0.002328216, 0.002176527, 0.002150555, 0.002064756, 
    0.002153034, 0.002130338, 0.001722128, 0.001005196, 0.0005359699,
  0.000699554, 0.0008198161, 0.0008361782, 0.0008853439, 0.0008195323, 
    0.0008181051, 0.000883347, 0.0008547409, 0.0008305495, 0.0007374068, 
    0.0007580665, 0.0007650347, 0.000775832, 0.0008242911, 0.0005635891,
  0.001103955, 0.00116016, 0.001256764, 0.001118203, 0.0007946377, 
    0.000854279, 0.001019641, 0.000992397, 0.0009725541, 0.0009312031, 
    0.001030779, 0.001165821, 0.001213479, 0.0009968622, 0.0005728762,
  0.001478889, 0.001482619, 0.001514723, 0.001481982, 0.001361945, 
    0.001039262, 0.00120927, 0.001243707, 0.001250267, 0.001301238, 
    0.001429166, 0.001602229, 0.001565523, 0.001393116, 0.0006128948,
  0.00171345, 0.001668374, 0.001635794, 0.001658227, 0.001664144, 0.00157775, 
    0.0009832403, 0.001361276, 0.001631058, 0.001746622, 0.002015434, 
    0.002009296, 0.001853636, 0.001549823, 0.000540811,
  0.001994272, 0.001881796, 0.001812508, 0.001811242, 0.001836097, 
    0.001862434, 0.001961708, 0.00164447, 0.001737116, 0.002137845, 
    0.002390249, 0.002101635, 0.001945733, 0.001563852, 0.0005319812,
  0.002434041, 0.002215894, 0.002054477, 0.002009465, 0.002029703, 
    0.002105238, 0.002232598, 0.002381328, 0.002502173, 0.002582751, 
    0.002313078, 0.001903123, 0.001899005, 0.001529317, 0.0004932131,
  0.002907392, 0.002677176, 0.002422991, 0.002299126, 0.002297581, 
    0.002359516, 0.002482549, 0.002639697, 0.002756238, 0.002486657, 
    0.001970892, 0.001824371, 0.001895514, 0.001292284, 0.0004454981,
  0.003234242, 0.003057419, 0.002830182, 0.00264621, 0.002558755, 
    0.002564156, 0.002623181, 0.002708294, 0.002448575, 0.002137295, 
    0.001718504, 0.001788519, 0.001869629, 0.001053781, 0.0003830277,
  0.003356381, 0.003252131, 0.003094602, 0.002881117, 0.00269839, 
    0.002633526, 0.002683086, 0.002623501, 0.002344706, 0.002133796, 
    0.001705492, 0.001815623, 0.001631507, 0.0007619575, 0.0002886952,
  0.003487154, 0.003374263, 0.00320562, 0.003026349, 0.002852073, 
    0.002759614, 0.002686532, 0.002489035, 0.002242773, 0.001851196, 
    0.001875475, 0.00182678, 0.001329434, 0.0005718228, 0.0003013432,
  0.0005653467, 0.0006503145, 0.0005754103, 0.0005638853, 0.0004959096, 
    0.0005122497, 0.0005771958, 0.0005580473, 0.0005469393, 0.0004914161, 
    0.0005083476, 0.0005760791, 0.0006128071, 0.0007766383, 0.000987743,
  0.001030076, 0.001044545, 0.001059994, 0.0008369387, 0.0004932333, 
    0.0005926592, 0.0007051868, 0.0006460512, 0.0006164488, 0.0005918749, 
    0.0005968311, 0.0007296065, 0.0008902244, 0.001141711, 0.001135792,
  0.001998008, 0.001745371, 0.001678479, 0.001545426, 0.0009355238, 
    0.000542226, 0.0007909504, 0.0007964802, 0.0007483989, 0.000725998, 
    0.0007637213, 0.0009157605, 0.001201304, 0.00142039, 0.0007627523,
  0.002638689, 0.002391872, 0.002125182, 0.001960309, 0.001757931, 
    0.001212068, 0.0006723693, 0.0008147266, 0.0009070331, 0.0009265517, 
    0.0009868335, 0.001205382, 0.00139437, 0.001380577, 0.0005289999,
  0.003200987, 0.003043976, 0.00279311, 0.002489886, 0.002220431, 0.00192935, 
    0.001514868, 0.0008159127, 0.000802559, 0.0009957084, 0.001191048, 
    0.001418144, 0.001523184, 0.001340613, 0.0005363777,
  0.003429885, 0.003359039, 0.003257617, 0.003058162, 0.002816097, 
    0.002500387, 0.00214814, 0.0016953, 0.001145376, 0.001081984, 
    0.001227081, 0.001507372, 0.001608677, 0.00110805, 0.0004609544,
  0.003293086, 0.003307332, 0.003352431, 0.003295023, 0.003244393, 
    0.003045368, 0.002770844, 0.002371054, 0.001928779, 0.001441952, 
    0.001407541, 0.001577815, 0.001502238, 0.0008322605, 0.0004164633,
  0.003235451, 0.00316531, 0.003233959, 0.00328374, 0.003319487, 0.003235711, 
    0.003075318, 0.002828456, 0.002510644, 0.001888882, 0.001626289, 
    0.001666274, 0.00141767, 0.0006550042, 0.0003647048,
  0.002666799, 0.002672524, 0.002842701, 0.003022116, 0.003131397, 
    0.003161776, 0.003022793, 0.002877151, 0.002733193, 0.002229221, 
    0.001816058, 0.001750398, 0.001275474, 0.0005207355, 0.0002949758,
  0.002536069, 0.002536399, 0.002712088, 0.002916442, 0.003100101, 
    0.003193051, 0.003148705, 0.003011506, 0.002843312, 0.002465795, 
    0.002073945, 0.00179914, 0.001098369, 0.0004498032, 0.0003100481,
  0.0006801357, 0.000764827, 0.0005610632, 0.0005722246, 0.0004503362, 
    0.0004434017, 0.000516502, 0.0004648652, 0.0004188386, 0.0002663599, 
    0.0002680117, 0.0003179486, 0.0002580939, 0.0002807371, 0.0002758795,
  0.001049558, 0.001086708, 0.000945367, 0.000705266, 0.0004249398, 
    0.0005290616, 0.0006166216, 0.0005080157, 0.0004598014, 0.0003707023, 
    0.0003250674, 0.000412379, 0.0004102991, 0.0003074974, 0.0002285541,
  0.001850608, 0.001618847, 0.001565045, 0.00130702, 0.0006143142, 
    0.0004399866, 0.0007271691, 0.0006192874, 0.0005144798, 0.0004357111, 
    0.0004421151, 0.0004252936, 0.0004359834, 0.0004674838, 0.0003640762,
  0.002718682, 0.002060678, 0.001886634, 0.001752448, 0.001386986, 
    0.0008578105, 0.0005414248, 0.000676735, 0.0006611613, 0.0005672392, 
    0.0005167002, 0.0004708103, 0.0004728396, 0.0005408352, 0.0004600755,
  0.00333237, 0.002616994, 0.002153359, 0.00199256, 0.001728831, 0.001521341, 
    0.001164922, 0.0005888499, 0.0005898732, 0.0006959871, 0.0007058849, 
    0.0006350819, 0.0005539877, 0.0006149995, 0.0005679997,
  0.002877526, 0.002867276, 0.002380818, 0.002195499, 0.001975042, 
    0.001809442, 0.001658665, 0.001435444, 0.0009012813, 0.0007790829, 
    0.0007850325, 0.0007761691, 0.0006728346, 0.0006900053, 0.0005980527,
  0.002721866, 0.002625021, 0.002409217, 0.00230155, 0.002126652, 
    0.001988027, 0.001866289, 0.001770607, 0.001625708, 0.001210466, 
    0.0009925193, 0.0008704768, 0.0007629557, 0.0007669591, 0.000578968,
  0.002678064, 0.00272123, 0.002629659, 0.002528702, 0.002390665, 
    0.002308975, 0.002190161, 0.002102792, 0.001967083, 0.001609177, 
    0.001257107, 0.001019281, 0.0008545594, 0.0007943923, 0.0005433467,
  0.002208588, 0.002297543, 0.002408716, 0.00240745, 0.002344756, 
    0.002351286, 0.002465079, 0.002457506, 0.002364893, 0.002077708, 
    0.001589581, 0.001188856, 0.0009318095, 0.0008058015, 0.0004308886,
  0.001902439, 0.001891904, 0.001857515, 0.001862941, 0.001937144, 
    0.001984441, 0.002150239, 0.002356383, 0.002594274, 0.002475013, 
    0.001991077, 0.00141547, 0.001035514, 0.0007986691, 0.0004506409,
  0.0007295397, 0.0008324006, 0.0007061284, 0.0007345272, 0.0006288448, 
    0.0006408401, 0.0007649553, 0.0005519106, 0.0004788841, 0.0003008391, 
    0.0002717559, 0.0002970071, 0.0001777537, 0.0001662506, 9.81405e-05,
  0.0009889022, 0.001068711, 0.0009282262, 0.0007779954, 0.0005619676, 
    0.0007151836, 0.0007954491, 0.000574571, 0.000529778, 0.0004376115, 
    0.0003476395, 0.0004578891, 0.0004044951, 0.0001562303, 9.111016e-05,
  0.001559616, 0.001463871, 0.001380804, 0.001093641, 0.0007463832, 
    0.000564754, 0.0008020338, 0.0006118673, 0.0005529851, 0.0004999259, 
    0.0005360996, 0.0004666483, 0.0003984795, 0.0003146709, 0.0001519918,
  0.001850971, 0.001748496, 0.001657002, 0.001524613, 0.001275157, 
    0.0009494949, 0.0005738006, 0.0006191641, 0.0006027998, 0.0005305011, 
    0.0005232096, 0.000480603, 0.0004106072, 0.0003658515, 0.0002325363,
  0.002078286, 0.001903944, 0.001784254, 0.001702762, 0.001551712, 
    0.001443962, 0.001193492, 0.0005305298, 0.0004884254, 0.0005503827, 
    0.0005935581, 0.0005669403, 0.0004569535, 0.0004641544, 0.0003687094,
  0.002264915, 0.002052471, 0.001909533, 0.00182865, 0.001700823, 
    0.001627614, 0.00158425, 0.001329946, 0.0008181965, 0.0006770099, 
    0.0006700777, 0.0006690326, 0.0005338861, 0.0005071366, 0.0004356909,
  0.002311235, 0.002207427, 0.002020054, 0.001895097, 0.001786723, 
    0.001713606, 0.001657722, 0.001586745, 0.001425917, 0.0009973689, 
    0.0008172445, 0.0007382343, 0.0006130614, 0.0005416268, 0.000475291,
  0.002318952, 0.002239102, 0.002081084, 0.001986654, 0.001852466, 
    0.001778331, 0.001692434, 0.001647165, 0.001563011, 0.001206807, 
    0.0008886121, 0.0007708575, 0.0006733821, 0.0005550971, 0.0004640881,
  0.002308368, 0.002263878, 0.002165323, 0.00205551, 0.001927608, 
    0.001836539, 0.001736998, 0.00167619, 0.001546799, 0.001331366, 
    0.001003389, 0.0008694191, 0.0007358936, 0.0005753356, 0.0004258345,
  0.002041172, 0.00209274, 0.002067862, 0.002034053, 0.001957567, 
    0.001890552, 0.001809561, 0.001762569, 0.001619371, 0.001375315, 
    0.001225714, 0.0009864488, 0.0008175382, 0.0006413048, 0.0004758633,
  0.0006924176, 0.000785089, 0.0007415057, 0.0007232876, 0.0005653313, 
    0.000544225, 0.0005748299, 0.0003997071, 0.0003769669, 0.0002224255, 
    0.0001756261, 0.0002068886, 0.0001607106, 0.0001554543, 0.0001161939,
  0.0009938903, 0.001042548, 0.001007521, 0.0007563527, 0.0005404075, 
    0.0005860864, 0.0005418597, 0.0004260966, 0.0004065919, 0.0003578054, 
    0.0002842385, 0.0003627777, 0.000338151, 0.0001402639, 0.0001053811,
  0.001461687, 0.001361495, 0.001335145, 0.0009544346, 0.0007474078, 
    0.0004153663, 0.0005218023, 0.0004619775, 0.0004611704, 0.0004571723, 
    0.0004602894, 0.0003616413, 0.0003451021, 0.0003112165, 0.0001754105,
  0.001705227, 0.001631223, 0.001575283, 0.00144781, 0.001225383, 
    0.0008673404, 0.0003997506, 0.0004810041, 0.0004874336, 0.0004389953, 
    0.0004248263, 0.0003546767, 0.0003300109, 0.0003195394, 0.000300882,
  0.001829736, 0.00174327, 0.001665047, 0.001607806, 0.00150465, 0.00133652, 
    0.001044295, 0.0004342902, 0.0003684447, 0.0003980269, 0.0004751119, 
    0.000428449, 0.0003760955, 0.0003906198, 0.0003893851,
  0.001921491, 0.001818144, 0.001728896, 0.001645071, 0.001591721, 
    0.001505118, 0.001427005, 0.001197398, 0.0008058314, 0.0006718881, 
    0.0006067447, 0.0005806125, 0.0004580909, 0.000429121, 0.0003854443,
  0.002043021, 0.001928245, 0.001794532, 0.001698048, 0.001603407, 
    0.001559556, 0.001450502, 0.001351744, 0.001238666, 0.00098761, 
    0.0008171339, 0.0006992315, 0.0005495303, 0.0004834245, 0.0004098232,
  0.002148894, 0.002017749, 0.001860049, 0.001753366, 0.001650754, 
    0.001586144, 0.001504414, 0.001453628, 0.001350679, 0.001071228, 
    0.0008455387, 0.0006986639, 0.0005965147, 0.0004848515, 0.000404595,
  0.002197345, 0.00209347, 0.001970924, 0.001814062, 0.001699995, 
    0.001603049, 0.001558949, 0.001488519, 0.001359148, 0.0011325, 
    0.0008524375, 0.0007399777, 0.0006477156, 0.0005126146, 0.0004200353,
  0.002225563, 0.002109728, 0.001968168, 0.001863603, 0.001750124, 
    0.001653766, 0.001564936, 0.001485748, 0.00142708, 0.001069214, 
    0.001067875, 0.0008652624, 0.0007183675, 0.0006029613, 0.0004960757,
  0.0005856088, 0.0006542181, 0.0006054405, 0.0005714492, 0.0004502237, 
    0.0004115941, 0.000448596, 0.0004011734, 0.0004419372, 0.0003177136, 
    0.0002583889, 0.0003183697, 0.0002269185, 0.0001838898, 0.0001324752,
  0.0009595355, 0.0009130124, 0.0008729884, 0.0005684305, 0.0004269073, 
    0.000376967, 0.0004147608, 0.0004094234, 0.0004410677, 0.0004655865, 
    0.0003472005, 0.0004403875, 0.0004347783, 0.0002007242, 0.0001454669,
  0.001318085, 0.001170483, 0.001103017, 0.0006910622, 0.0005854084, 
    0.0002807908, 0.0004097836, 0.0004373883, 0.0004547601, 0.0004669891, 
    0.0004639566, 0.0004352486, 0.0004535422, 0.0004228121, 0.0002457704,
  0.00151722, 0.001440006, 0.001360184, 0.00113792, 0.001020543, 
    0.0006556257, 0.0003290131, 0.0004038284, 0.000432577, 0.0004195703, 
    0.000416479, 0.000413151, 0.0004371831, 0.000462166, 0.0004259939,
  0.001592805, 0.0014896, 0.001413063, 0.001321107, 0.00120365, 0.001066488, 
    0.0009455788, 0.0003461261, 0.0002796785, 0.0003870326, 0.000476735, 
    0.0004918539, 0.0004637253, 0.0004987291, 0.0005519452,
  0.001597805, 0.001503231, 0.001439677, 0.001360388, 0.001291887, 
    0.001209173, 0.001138792, 0.0009952913, 0.0007396303, 0.0006839994, 
    0.0005417907, 0.0005729682, 0.0005075648, 0.0004952345, 0.0005332779,
  0.001600043, 0.001516102, 0.001451074, 0.001377596, 0.001347307, 
    0.001291168, 0.001223658, 0.001111259, 0.001048288, 0.0008592383, 
    0.0007015942, 0.0006278704, 0.000564535, 0.0005177733, 0.0005041157,
  0.001620217, 0.001538604, 0.00146637, 0.001409505, 0.001375973, 
    0.001349368, 0.001287955, 0.001247152, 0.001074428, 0.0008601648, 
    0.0007181838, 0.000652898, 0.0006163655, 0.0005208545, 0.0005463911,
  0.001653038, 0.001571015, 0.001527611, 0.001445692, 0.001391886, 
    0.001369118, 0.001304432, 0.001250981, 0.001105719, 0.0008392819, 
    0.0007528021, 0.0007381953, 0.000696536, 0.0005850735, 0.0005862475,
  0.001663509, 0.001562643, 0.001510915, 0.001450657, 0.001397134, 
    0.00134126, 0.001270592, 0.001206954, 0.001079183, 0.000700467, 
    0.0008202506, 0.0008618213, 0.0007969311, 0.0006861088, 0.0006486044,
  0.0005718856, 0.0006575185, 0.000581726, 0.0005798685, 0.0004978992, 
    0.0004434825, 0.0004855823, 0.000452778, 0.0004439391, 0.000286967, 
    0.0002118449, 0.0002300698, 0.0002009032, 0.0002044125, 0.0001564908,
  0.000962219, 0.0008876296, 0.0007969941, 0.000594289, 0.0004487896, 
    0.0003780686, 0.0004909456, 0.0004998168, 0.0005144307, 0.0005024357, 
    0.0004056095, 0.0004557274, 0.0004740272, 0.0002956806, 0.0002305706,
  0.001332828, 0.001097304, 0.001045105, 0.0007215677, 0.0006638818, 
    0.0002905615, 0.000471285, 0.0005333505, 0.0005577914, 0.0005630927, 
    0.0005647501, 0.0005649414, 0.0005839382, 0.0005873004, 0.0004456201,
  0.001554049, 0.001409102, 0.001295386, 0.001108189, 0.001060434, 
    0.0007900883, 0.0003398995, 0.0005312208, 0.0006076843, 0.0005964773, 
    0.0005905885, 0.000625112, 0.0006765665, 0.0007384684, 0.0007092804,
  0.001653976, 0.001513857, 0.00140855, 0.001341148, 0.001234739, 
    0.001146543, 0.001217879, 0.0004293392, 0.000455818, 0.0006248479, 
    0.0006669543, 0.0007317648, 0.0007570075, 0.0008416215, 0.0008694509,
  0.001713462, 0.001582627, 0.001495232, 0.001422251, 0.001368435, 
    0.001339724, 0.001257881, 0.001132843, 0.0009529184, 0.0008073782, 
    0.0006767202, 0.0007712537, 0.0008301546, 0.0008903242, 0.0009823235,
  0.0017863, 0.001686725, 0.00155625, 0.001473905, 0.001424833, 0.001406805, 
    0.001379112, 0.001320676, 0.001168384, 0.0009218896, 0.000796016, 
    0.0007762514, 0.0008206377, 0.0008830959, 0.0009879469,
  0.001832729, 0.001716812, 0.001611666, 0.001521661, 0.001443346, 
    0.001420659, 0.00138205, 0.001347773, 0.001167099, 0.0009128304, 
    0.0008228784, 0.0007666813, 0.0007644899, 0.0008074811, 0.0009338213,
  0.001819699, 0.00174293, 0.001659033, 0.001552702, 0.001464309, 
    0.001408877, 0.001362894, 0.001293366, 0.001258953, 0.001017803, 
    0.0009370961, 0.0008281206, 0.0007402391, 0.0007579487, 0.0008346671,
  0.001780895, 0.001698511, 0.001640098, 0.001540311, 0.0014702, 0.001361023, 
    0.001278393, 0.001257438, 0.001207715, 0.000980781, 0.001076019, 
    0.0008929817, 0.0007392342, 0.0006933187, 0.000774834,
  0.0006187005, 0.0006576809, 0.0005988256, 0.0005145984, 0.000441419, 
    0.0003932725, 0.0003685628, 0.0003525113, 0.0003623695, 0.0002307781, 
    0.000202856, 0.0002700946, 0.0002514528, 0.0002700058, 0.0002093802,
  0.0008827003, 0.0007882376, 0.0007035334, 0.0005636833, 0.0004722332, 
    0.0003722064, 0.000455437, 0.0004257986, 0.0004215823, 0.0003921341, 
    0.0003131181, 0.0004162567, 0.0004505159, 0.0002473947, 0.0001795486,
  0.001139758, 0.0009596285, 0.0009475602, 0.0006904483, 0.000642782, 
    0.0002975216, 0.0005415981, 0.0005700586, 0.0005587896, 0.0005276586, 
    0.0005005422, 0.0005260546, 0.0005367108, 0.0005166429, 0.0003029112,
  0.001339609, 0.001263264, 0.001228132, 0.001083822, 0.001057791, 
    0.000837152, 0.0004386109, 0.0006647559, 0.0006985556, 0.0006202398, 
    0.000564122, 0.0005747019, 0.000580575, 0.0005753569, 0.0004347412,
  0.001440472, 0.001402037, 0.001425468, 0.001488343, 0.001399742, 
    0.001306242, 0.001198223, 0.000573448, 0.0005647462, 0.0006407632, 
    0.0007083645, 0.000676349, 0.0006772261, 0.0006839155, 0.0005588837,
  0.001574434, 0.001537906, 0.001545052, 0.001602249, 0.001653891, 
    0.001552669, 0.001421333, 0.001230917, 0.001044134, 0.0009565089, 
    0.0007746632, 0.0008407736, 0.000780293, 0.0007134754, 0.0006710378,
  0.001686243, 0.001661366, 0.001655966, 0.00168232, 0.001670577, 
    0.001708584, 0.001633301, 0.001464978, 0.001214125, 0.001075625, 
    0.001020806, 0.0009364937, 0.0008480718, 0.0007394461, 0.0007220028,
  0.001800049, 0.001739491, 0.00169577, 0.001690458, 0.001682626, 
    0.001676549, 0.001598556, 0.001466744, 0.001161866, 0.001073006, 
    0.001060551, 0.001043072, 0.001016147, 0.001044748, 0.001099097,
  0.001862204, 0.001783245, 0.001724745, 0.001685196, 0.001646061, 
    0.001629141, 0.001573864, 0.001428878, 0.001214002, 0.001070262, 
    0.001049793, 0.001041796, 0.001012451, 0.0009542105, 0.0009074672,
  0.001878266, 0.001775865, 0.001701103, 0.00163127, 0.001547736, 
    0.001516532, 0.001455474, 0.001383164, 0.001124563, 0.001004735, 
    0.0009698153, 0.0008945802, 0.0008738083, 0.0008339591, 0.0008403087,
  0.0005247268, 0.0005166846, 0.0004362356, 0.0004599867, 0.0004034601, 
    0.0004306459, 0.000509102, 0.0005583526, 0.0005952805, 0.0005120296, 
    0.0004786394, 0.0004708976, 0.000365667, 0.0003343772, 0.0002320368,
  0.0007512511, 0.00067175, 0.0005970386, 0.0005017136, 0.0004091033, 
    0.0003795661, 0.0005355185, 0.0005893821, 0.0006297979, 0.0006534199, 
    0.0005711545, 0.0006045422, 0.0005594786, 0.0003176811, 0.0002414889,
  0.001058288, 0.0008611314, 0.0008543879, 0.0005987749, 0.0005371646, 
    0.0002926128, 0.0005163579, 0.0005851996, 0.0006259656, 0.0006505011, 
    0.0006494515, 0.0006293396, 0.0006058646, 0.0004891727, 0.0003546571,
  0.001322816, 0.00120849, 0.00115602, 0.000923404, 0.0008615024, 
    0.0006656286, 0.0003646857, 0.0005181297, 0.000591674, 0.0005979706, 
    0.0006160634, 0.0006066205, 0.0005863518, 0.0005067084, 0.0004394632,
  0.001463922, 0.001421149, 0.001356309, 0.001262846, 0.001175242, 
    0.00105552, 0.001032866, 0.0004134533, 0.000372236, 0.000530567, 
    0.0006512934, 0.000672565, 0.0006680376, 0.000623363, 0.0005709312,
  0.001622652, 0.001604425, 0.001556579, 0.001479653, 0.001417674, 
    0.001280261, 0.001152468, 0.001089926, 0.0008878991, 0.0007254849, 
    0.0006813114, 0.0007465268, 0.0007227878, 0.0006958267, 0.0006727126,
  0.001783108, 0.001805619, 0.001741442, 0.001637089, 0.001563679, 
    0.001494439, 0.001358996, 0.001239676, 0.001082664, 0.0008601652, 
    0.0008037882, 0.0007434867, 0.000721026, 0.0006649557, 0.0006572898,
  0.001906366, 0.001897818, 0.001862454, 0.001761604, 0.001685654, 
    0.001573412, 0.00148202, 0.00142743, 0.001065721, 0.0008834114, 
    0.0008306673, 0.000792676, 0.0008215234, 0.0007718826, 0.000690217,
  0.001970042, 0.001888875, 0.001849998, 0.001803312, 0.00174351, 
    0.001640602, 0.001540977, 0.001437642, 0.001093965, 0.0009749447, 
    0.0009575898, 0.0009466455, 0.0008583429, 0.0007019087, 0.000591682,
  0.001969372, 0.001864054, 0.001827213, 0.001762563, 0.001694011, 
    0.001614165, 0.001536811, 0.001412467, 0.001089657, 0.001010443, 
    0.001014651, 0.0009541269, 0.0007618876, 0.0006473941, 0.0006275031,
  0.0004073874, 0.0005107169, 0.0004740721, 0.0005027748, 0.0004340613, 
    0.0005044807, 0.0006188334, 0.000599008, 0.0005433502, 0.0004235375, 
    0.0003992458, 0.0003560575, 0.0002565107, 0.0002085072, 0.000147591,
  0.0006541832, 0.0006702241, 0.0006318553, 0.0005459759, 0.000418003, 
    0.0004876664, 0.0006866258, 0.0006453819, 0.0006266379, 0.0005779359, 
    0.0004003131, 0.0004101819, 0.0003623016, 0.0002020372, 0.0001893421,
  0.0009999098, 0.0008748423, 0.0008717897, 0.0007165194, 0.0006760177, 
    0.0005079159, 0.0007202918, 0.000715833, 0.0006756208, 0.0005862821, 
    0.000501714, 0.0004573408, 0.0004207325, 0.0003758379, 0.0002813645,
  0.001226679, 0.001141382, 0.001111684, 0.001004678, 0.0009535495, 
    0.0008199952, 0.0005356367, 0.0006528233, 0.000603213, 0.0005578814, 
    0.0004979548, 0.0004475554, 0.0004138827, 0.0003930281, 0.0003847441,
  0.001315163, 0.001253072, 0.001234828, 0.001303126, 0.001311996, 
    0.001156464, 0.001065033, 0.0004814526, 0.0004228103, 0.0004726764, 
    0.0004907349, 0.0004482598, 0.0004385923, 0.000454229, 0.00045684,
  0.001427961, 0.001336003, 0.001347264, 0.001442376, 0.001484175, 
    0.001405685, 0.001287055, 0.001101972, 0.0008650123, 0.000652621, 
    0.0005190957, 0.0004920925, 0.0004804502, 0.0004933071, 0.0005077912,
  0.001579026, 0.001494256, 0.001479561, 0.001540067, 0.001588886, 
    0.001515774, 0.001426502, 0.001269408, 0.001033285, 0.0007253136, 
    0.0006055257, 0.0005441133, 0.000517192, 0.000497528, 0.0005207729,
  0.001731668, 0.001623924, 0.001585322, 0.001601228, 0.001616978, 
    0.001555127, 0.00153636, 0.00144524, 0.001002362, 0.0007510739, 
    0.0006286799, 0.0005876807, 0.0005415299, 0.0005082281, 0.0005263515,
  0.001903144, 0.001801499, 0.001742473, 0.001677367, 0.00165415, 0.00158608, 
    0.00155488, 0.001377153, 0.0009638484, 0.0007640557, 0.0006607713, 
    0.0006202154, 0.0005427513, 0.000517075, 0.0005337641,
  0.002030627, 0.001907552, 0.001804237, 0.001701253, 0.001654983, 
    0.00159922, 0.001496471, 0.001310767, 0.0008989641, 0.0007840237, 
    0.0007173171, 0.0006520152, 0.0005693614, 0.0005567972, 0.0005688053,
  0.0004303547, 0.0005326619, 0.0005326574, 0.0005586045, 0.0005672906, 
    0.0006011114, 0.0006316047, 0.000548024, 0.0004873729, 0.0003341761, 
    0.0002858212, 0.0002826518, 0.0002444095, 0.0002090949, 0.0001454625,
  0.0006786347, 0.0006983176, 0.0006924506, 0.0006323516, 0.0004721299, 
    0.0004894248, 0.0005655062, 0.0005047912, 0.0004580795, 0.0004165851, 
    0.0003427831, 0.0003741953, 0.00037416, 0.0001973809, 0.0001571866,
  0.001063292, 0.001005129, 0.0009631138, 0.0008463382, 0.0006772261, 
    0.0003279746, 0.00054142, 0.0004864706, 0.0004690681, 0.0004782249, 
    0.0004672509, 0.0004189939, 0.0004115146, 0.0003756038, 0.0002558292,
  0.001251503, 0.001249624, 0.001214031, 0.001114155, 0.001078113, 
    0.0008249928, 0.0003696456, 0.0004372478, 0.000457124, 0.0004684186, 
    0.0004530007, 0.0003985562, 0.0003967448, 0.0003607258, 0.0003565148,
  0.001354336, 0.001341466, 0.001349892, 0.001325526, 0.001329054, 
    0.001243493, 0.001000724, 0.0003344009, 0.0003012358, 0.0003811678, 
    0.0004263748, 0.0003920261, 0.0003969672, 0.0004059383, 0.0004262927,
  0.001458962, 0.001432228, 0.001424491, 0.001417033, 0.001395479, 
    0.00142582, 0.00119264, 0.0009944973, 0.0006853417, 0.0005314907, 
    0.0004457197, 0.0004134396, 0.000414441, 0.0004358093, 0.0004709706,
  0.001589975, 0.001554282, 0.001538829, 0.001518989, 0.001514671, 
    0.001499439, 0.001361248, 0.001151722, 0.000828848, 0.0005807749, 
    0.0005001341, 0.0004523921, 0.0004405593, 0.0004462778, 0.0004856369,
  0.001688718, 0.001659646, 0.001642105, 0.001627009, 0.001600607, 
    0.001539336, 0.001491547, 0.001342492, 0.0008895045, 0.0005810359, 
    0.000515798, 0.0004751439, 0.0004581274, 0.0004433861, 0.0004803547,
  0.00176017, 0.001748205, 0.001764371, 0.001727974, 0.001716216, 
    0.001592448, 0.001551704, 0.001441663, 0.000929083, 0.0005750755, 
    0.0005085748, 0.0004911426, 0.0004653758, 0.0004494547, 0.0004877269,
  0.001817578, 0.001813841, 0.001819916, 0.00175543, 0.001726169, 
    0.001603694, 0.001581057, 0.001558635, 0.000935591, 0.0006089162, 
    0.0005748129, 0.0005330728, 0.0004934762, 0.000498339, 0.0005160999,
  0.0005127306, 0.0005749416, 0.0006136285, 0.0006841084, 0.0006089194, 
    0.0005742068, 0.000535237, 0.000429338, 0.0003139288, 0.0001737405, 
    0.0001842047, 0.0002430909, 0.000240153, 0.0001845627, 0.0001208891,
  0.0006810588, 0.0007002176, 0.0007640107, 0.0008527758, 0.0005465564, 
    0.0004139814, 0.0005164683, 0.0004617228, 0.0003609374, 0.0003059128, 
    0.0002270492, 0.0003333046, 0.0004009366, 0.000175794, 0.0001179894,
  0.00115758, 0.001082612, 0.001010269, 0.001020879, 0.0008706738, 
    0.0003541229, 0.000433091, 0.0004750963, 0.0004071372, 0.0003671065, 
    0.0003308249, 0.000375557, 0.0004471321, 0.0003772949, 0.0002302658,
  0.001465496, 0.001395941, 0.001340597, 0.001261311, 0.001427426, 
    0.001050678, 0.0003086906, 0.0004182582, 0.0004326778, 0.0004176333, 
    0.0003659884, 0.0003633382, 0.0004275634, 0.0004008291, 0.0003045686,
  0.001580023, 0.001502439, 0.001463306, 0.001417994, 0.001453734, 
    0.001773983, 0.001152365, 0.0003285585, 0.0002882202, 0.000403541, 
    0.0003805824, 0.0003656714, 0.0004032585, 0.0004141425, 0.000374797,
  0.001705385, 0.001609118, 0.00153036, 0.00148323, 0.001472427, 0.001625243, 
    0.001664533, 0.001060917, 0.0006880607, 0.0006165573, 0.0004834192, 
    0.0004020072, 0.0003989803, 0.0003986054, 0.0003937005,
  0.001827581, 0.00171268, 0.001600359, 0.001549551, 0.001520419, 
    0.001551976, 0.001729217, 0.001586599, 0.001066657, 0.0007054508, 
    0.0005610836, 0.0004352505, 0.0004108092, 0.0003919176, 0.0003984916,
  0.001859566, 0.001733822, 0.001650438, 0.001605535, 0.001589191, 
    0.001584646, 0.001668806, 0.001726685, 0.001258229, 0.0007848954, 
    0.0005856288, 0.0004649977, 0.0004180476, 0.0003858688, 0.0003910066,
  0.0018702, 0.001752419, 0.001700523, 0.001668845, 0.001665621, 0.001667712, 
    0.0017311, 0.001796085, 0.001286869, 0.0007665904, 0.0005920796, 
    0.0004998082, 0.0004353566, 0.0003918699, 0.0003999998,
  0.001831736, 0.00172062, 0.001704715, 0.001718669, 0.001755595, 
    0.001824973, 0.001995602, 0.001977602, 0.001243934, 0.0008305419, 
    0.0007094428, 0.0005371905, 0.0004656737, 0.0004307771, 0.0004202875,
  0.0006322965, 0.0006231727, 0.0005519156, 0.0005999494, 0.0005706662, 
    0.0004112769, 0.0003251959, 0.0003335803, 0.0002884123, 0.0001565802, 
    0.0001812143, 0.0002466754, 0.0001911947, 0.0001567366, 9.944328e-05,
  0.0008096626, 0.0007615653, 0.0006914344, 0.0006693723, 0.0005338459, 
    0.0003507842, 0.0003428124, 0.0003357922, 0.0002942935, 0.0002578018, 
    0.0002560167, 0.0003415314, 0.0003455105, 0.0001487824, 9.119018e-05,
  0.001291418, 0.001138995, 0.0009557988, 0.0007771789, 0.0006309345, 
    0.0002707906, 0.0003394031, 0.0003394329, 0.0003040755, 0.0003157899, 
    0.0003358297, 0.0004445845, 0.0005018587, 0.0003350989, 0.0002077825,
  0.001808081, 0.001590736, 0.001435761, 0.001171531, 0.0009440146, 
    0.0005944336, 0.0002716359, 0.0003085485, 0.0003197436, 0.0003315659, 
    0.0003390249, 0.0004176011, 0.0005239177, 0.0004106844, 0.0002713884,
  0.001980488, 0.00182539, 0.001650825, 0.001490263, 0.001364868, 
    0.001173966, 0.0008764457, 0.0002887363, 0.0002322767, 0.0002995268, 
    0.0003464627, 0.0003860197, 0.0004957968, 0.0005034846, 0.0003391684,
  0.002058572, 0.001973154, 0.001786517, 0.001625386, 0.001506016, 
    0.001420674, 0.001297388, 0.0009788538, 0.0006643861, 0.0006118299, 
    0.000446722, 0.0004008396, 0.0004311253, 0.0004661773, 0.0004105966,
  0.002124534, 0.002082193, 0.001904556, 0.001739875, 0.001599889, 
    0.001513185, 0.001496438, 0.001420739, 0.00116432, 0.0008327502, 
    0.0005829454, 0.000435194, 0.0004209805, 0.0004322569, 0.0004081672,
  0.002159232, 0.002125997, 0.001952673, 0.001785281, 0.001656811, 
    0.001563771, 0.001516516, 0.001584591, 0.001513697, 0.001162049, 
    0.0007101358, 0.0004787908, 0.0004234045, 0.0003936396, 0.0003809863,
  0.002135344, 0.002128656, 0.002010815, 0.001823467, 0.001676293, 
    0.001587593, 0.001541808, 0.001581278, 0.001535262, 0.001362893, 
    0.001040132, 0.0006484551, 0.0004637388, 0.000386225, 0.000361999,
  0.002085827, 0.002098765, 0.002005548, 0.00183694, 0.001691083, 
    0.001606739, 0.001596637, 0.001723992, 0.001463401, 0.001317217, 
    0.001294283, 0.0009749298, 0.0006592514, 0.0004801042, 0.0003849557,
  0.00158845, 0.001377933, 0.0008541885, 0.0005373025, 0.0003824715, 
    0.0003146108, 0.000323176, 0.0003459796, 0.0003158007, 0.0001713678, 
    0.0001737625, 0.0001631344, 0.0001296445, 0.0001329196, 8.302342e-05,
  0.001874593, 0.001561322, 0.001051528, 0.0005817279, 0.0003722941, 
    0.000292436, 0.000326121, 0.0003456204, 0.0003299418, 0.0002641934, 
    0.0002339711, 0.0002589065, 0.0002442328, 0.0001212231, 8.409774e-05,
  0.002289322, 0.001972532, 0.001249155, 0.0006778628, 0.0004822811, 
    0.0002439988, 0.0003054616, 0.0003338121, 0.0003301409, 0.0003204297, 
    0.0003237636, 0.0003348644, 0.0003096777, 0.0002637092, 0.000178404,
  0.002478483, 0.002337811, 0.001775541, 0.001073807, 0.0007646697, 
    0.0005092127, 0.0002547379, 0.0002794756, 0.0003154978, 0.0003198836, 
    0.0003426086, 0.0003833497, 0.0003672465, 0.0003049737, 0.0002309412,
  0.002532377, 0.002489975, 0.002056215, 0.001545686, 0.001256097, 
    0.0009891891, 0.0007780224, 0.0002787478, 0.0002253275, 0.0002819333, 
    0.0003473227, 0.0004030042, 0.0004073649, 0.0003649933, 0.0002928606,
  0.002513417, 0.002525598, 0.002257532, 0.001726128, 0.001483816, 
    0.001301132, 0.001114577, 0.0008278551, 0.0005746404, 0.0005336804, 
    0.0004156426, 0.0004116021, 0.0004277247, 0.0003994276, 0.0003226194,
  0.002493319, 0.002495968, 0.00239591, 0.001847126, 0.001592779, 
    0.001435368, 0.001294059, 0.00103447, 0.0008246849, 0.0006852256, 
    0.0005418635, 0.0004400201, 0.000437693, 0.0004056235, 0.0003548785,
  0.002387463, 0.002432771, 0.002477369, 0.001989007, 0.001637984, 
    0.001528635, 0.001367236, 0.001255106, 0.0009848808, 0.0007482301, 
    0.000577055, 0.0004630541, 0.0004403637, 0.000393348, 0.0003616354,
  0.002228634, 0.002322911, 0.002481524, 0.002101625, 0.001716024, 
    0.001515864, 0.001419264, 0.001272161, 0.00101058, 0.000766686, 
    0.0006381872, 0.0005033936, 0.000449755, 0.0003854001, 0.0003442006,
  0.002056411, 0.002239886, 0.002405729, 0.002149654, 0.001777704, 
    0.001503761, 0.00135573, 0.001270329, 0.000978082, 0.0008158032, 
    0.0008165108, 0.0006756607, 0.0005218682, 0.0004325178, 0.0003647451,
  0.001788514, 0.002083512, 0.002064215, 0.001379205, 0.0007337383, 
    0.0004241287, 0.0003917962, 0.0003739761, 0.0002841234, 0.0001324584, 
    0.0001323175, 0.0001258613, 0.0001005381, 0.0001086667, 7.77211e-05,
  0.002280897, 0.002479991, 0.002305895, 0.001269693, 0.0005013824, 
    0.0003713685, 0.000363158, 0.0003495768, 0.0002770648, 0.0002186525, 
    0.0001616173, 0.0002000587, 0.0001900841, 9.789969e-05, 7.170482e-05,
  0.002570158, 0.002651348, 0.002378656, 0.001230249, 0.0005892372, 
    0.0002734232, 0.0003186292, 0.0003312869, 0.0002818084, 0.0002602013, 
    0.0002336933, 0.0002266548, 0.0002197879, 0.0001936639, 0.0001392066,
  0.002665909, 0.002745451, 0.00266172, 0.001554082, 0.0008924948, 
    0.0005761168, 0.0002488112, 0.0002677501, 0.0002747794, 0.0002601634, 
    0.0002407563, 0.0002396113, 0.0002294277, 0.0002101772, 0.0001883238,
  0.002612764, 0.002666098, 0.002758419, 0.002087655, 0.001323277, 0.0010004, 
    0.0007515568, 0.0002527315, 0.0001886493, 0.0002334275, 0.0002595131, 
    0.0002587342, 0.0002538525, 0.0002410527, 0.000231522,
  0.002556524, 0.002516488, 0.002750165, 0.002343241, 0.00167217, 
    0.001360676, 0.001068804, 0.0007332303, 0.0005039957, 0.0004524034, 
    0.000326003, 0.0002969279, 0.0002762744, 0.0002647685, 0.000242752,
  0.002448656, 0.002356928, 0.002635016, 0.002495634, 0.001820792, 
    0.001482749, 0.001214966, 0.0008595723, 0.000639924, 0.0005562777, 
    0.0004265732, 0.0003328327, 0.0003031396, 0.0002864437, 0.0002645411,
  0.002124674, 0.002171137, 0.002506094, 0.002552831, 0.001887156, 
    0.001531169, 0.001311573, 0.001111578, 0.0007839386, 0.0005395281, 
    0.000424881, 0.0003544182, 0.0003295632, 0.0003079343, 0.0002874906,
  0.001988614, 0.002119085, 0.002436906, 0.002571176, 0.001944025, 
    0.001515406, 0.001328809, 0.001195157, 0.0007543462, 0.0005386302, 
    0.0004450878, 0.0003857067, 0.0003606166, 0.0003277659, 0.0002993692,
  0.002107645, 0.002393509, 0.002553513, 0.002536366, 0.001902389, 
    0.00149546, 0.001263589, 0.001117065, 0.0006825865, 0.0005573121, 
    0.0005249615, 0.0004236083, 0.0003964195, 0.0003599145, 0.0003182816,
  0.0014721, 0.001507686, 0.001520399, 0.00162025, 0.001435081, 0.001073944, 
    0.0008217612, 0.000576797, 0.000339223, 0.0001588538, 0.0001528539, 
    0.0001399442, 0.0001159103, 0.0001203024, 8.000408e-05,
  0.001723359, 0.001677391, 0.001634382, 0.001678849, 0.00130113, 
    0.0008496913, 0.0006383686, 0.0004696124, 0.0003164354, 0.0002457236, 
    0.000181658, 0.0002154088, 0.000202649, 9.648546e-05, 6.521778e-05,
  0.00212047, 0.002068869, 0.001939861, 0.001813709, 0.001339113, 
    0.0005349072, 0.000442088, 0.000397558, 0.0002948052, 0.0002730586, 
    0.0002536751, 0.000245971, 0.000225632, 0.0001933391, 0.0001351125,
  0.002290971, 0.002257395, 0.002217982, 0.002115353, 0.00160935, 
    0.0008707701, 0.0003268787, 0.0002781323, 0.0002712007, 0.0002524453, 
    0.0002597742, 0.0002414861, 0.0002187049, 0.0001935934, 0.0001713781,
  0.002467302, 0.002431209, 0.002383968, 0.002365045, 0.001913374, 
    0.001271744, 0.0009206377, 0.0002718186, 0.0001918067, 0.0002185572, 
    0.0002555993, 0.0002451218, 0.0002220033, 0.0002071245, 0.0001972469,
  0.002457139, 0.002559354, 0.002547817, 0.002506684, 0.002215912, 
    0.001740774, 0.001341747, 0.0008794629, 0.0005413385, 0.0004347629, 
    0.0003212593, 0.0002675259, 0.0002322971, 0.0002060173, 0.000194373,
  0.002319959, 0.002519393, 0.002600126, 0.002592246, 0.002249224, 
    0.001799351, 0.001423892, 0.000940942, 0.0006402343, 0.0005589069, 
    0.0004159654, 0.0002851874, 0.0002408873, 0.000211045, 0.0001996041,
  0.002377447, 0.002466627, 0.002580328, 0.002604974, 0.002209782, 
    0.00178451, 0.001441664, 0.001114036, 0.0006937112, 0.000467519, 
    0.0003599089, 0.0002804305, 0.000241019, 0.0002142884, 0.0002098369,
  0.002183978, 0.002340618, 0.002465471, 0.002518597, 0.002118156, 
    0.00171053, 0.001404293, 0.001152458, 0.0005977495, 0.0003998225, 
    0.0003272045, 0.0002698214, 0.0002464637, 0.0002255907, 0.0002242257,
  0.002214205, 0.00232341, 0.002432878, 0.002434932, 0.001969228, 
    0.001570355, 0.001264045, 0.000937485, 0.000461581, 0.0004038838, 
    0.0003686268, 0.0002850552, 0.0002696054, 0.0002491255, 0.0002445522,
  0.001682732, 0.001637013, 0.001573536, 0.001514004, 0.001418405, 
    0.00132385, 0.001309588, 0.001134887, 0.0008546943, 0.0004394516, 
    0.000278323, 0.0002176622, 0.0001344137, 0.0001279439, 0.0001078438,
  0.002065493, 0.001952807, 0.001778976, 0.001628828, 0.001458698, 
    0.001328439, 0.00124336, 0.00103556, 0.0007671715, 0.0004976078, 
    0.0003122342, 0.0002924677, 0.0002446827, 0.0001138705, 8.886679e-05,
  0.002302187, 0.002275081, 0.002113603, 0.001784727, 0.001531687, 
    0.001039922, 0.001002856, 0.0008729914, 0.0006316206, 0.0004742864, 
    0.0003656188, 0.000334881, 0.0002887954, 0.0002416324, 0.0001799217,
  0.002351838, 0.0023164, 0.002280603, 0.002052877, 0.001708228, 0.00136983, 
    0.0005739869, 0.0004935617, 0.0004410739, 0.0003989936, 0.0003544728, 
    0.0003166939, 0.0002965113, 0.0002570392, 0.0002218883,
  0.002554665, 0.002550329, 0.002433244, 0.002210638, 0.001813459, 
    0.001562095, 0.001154278, 0.000371131, 0.0002830619, 0.0003026123, 
    0.000324561, 0.0003164102, 0.000295331, 0.0002671587, 0.0002432657,
  0.00239094, 0.002536242, 0.002603415, 0.002311832, 0.001904651, 
    0.001631405, 0.001461031, 0.0010268, 0.0007010218, 0.0005014083, 
    0.0003955241, 0.0003357001, 0.0002919812, 0.0002534097, 0.0002264192,
  0.002303933, 0.002341088, 0.002667683, 0.002386919, 0.001910156, 
    0.001659612, 0.001420807, 0.001166737, 0.0009215279, 0.0006842738, 
    0.0005194001, 0.0003404091, 0.0002818911, 0.0002345094, 0.0002211235,
  0.002495742, 0.002556324, 0.002700903, 0.002289371, 0.001924546, 
    0.001653782, 0.001481798, 0.00128762, 0.0008795908, 0.000556442, 
    0.0004503621, 0.0003206656, 0.0002716365, 0.0002224706, 0.0002203884,
  0.002694115, 0.002674519, 0.002573563, 0.002195125, 0.001862943, 
    0.001652143, 0.001574004, 0.001293028, 0.0006846573, 0.0004367235, 
    0.0003694253, 0.0002932709, 0.0002459498, 0.0002160875, 0.0002356524,
  0.002487849, 0.002401477, 0.002247307, 0.002023692, 0.001785313, 
    0.001646662, 0.001480209, 0.000820075, 0.0004333786, 0.0004049456, 
    0.0003876448, 0.0002880701, 0.0002561111, 0.0002353433, 0.0002663662,
  0.001388963, 0.001414516, 0.001342994, 0.001289736, 0.001190149, 
    0.001072975, 0.001081156, 0.001052365, 0.001031396, 0.000716695, 
    0.0006263231, 0.0005870977, 0.0004108562, 0.0003447016, 0.0002773058,
  0.002048249, 0.001826081, 0.001620185, 0.001446345, 0.001274716, 
    0.001188412, 0.001183155, 0.001098835, 0.001045177, 0.0009851148, 
    0.0007819667, 0.0007620232, 0.0005785798, 0.0002788048, 0.0002087615,
  0.002513092, 0.002522325, 0.002356638, 0.001954539, 0.001550898, 
    0.00111032, 0.001131791, 0.001079289, 0.0009477386, 0.0009374568, 
    0.000874248, 0.00075061, 0.0005664859, 0.0003852696, 0.0002522979,
  0.002599277, 0.002691265, 0.002756071, 0.002728193, 0.002217709, 
    0.00159661, 0.000864241, 0.0008034654, 0.0007419052, 0.0007506339, 
    0.0007370946, 0.0006392387, 0.0004887801, 0.0003422306, 0.0002578513,
  0.002463548, 0.002659298, 0.002767337, 0.002869544, 0.002749179, 
    0.002231137, 0.001593711, 0.0007453364, 0.0006505611, 0.000547498, 
    0.0006003301, 0.0005571686, 0.0004147899, 0.0003216909, 0.0002623099,
  0.002280655, 0.002509686, 0.002639315, 0.00287073, 0.002828708, 
    0.002301225, 0.001780605, 0.001347582, 0.001011422, 0.0008194334, 
    0.0006303372, 0.0004930773, 0.0003726489, 0.000288576, 0.0002420636,
  0.002170723, 0.002357901, 0.002712758, 0.0028019, 0.002517783, 0.001959955, 
    0.001531567, 0.001195132, 0.001011854, 0.0008831205, 0.0006940941, 
    0.0004496667, 0.0003369999, 0.0002671945, 0.0002289221,
  0.002009826, 0.002025074, 0.002054397, 0.002053303, 0.00181563, 
    0.001550847, 0.00138301, 0.001203043, 0.0008626697, 0.0007165617, 
    0.0005538819, 0.0003811897, 0.0003201945, 0.0002447026, 0.0002342846,
  0.001869195, 0.001780119, 0.001711967, 0.001627842, 0.001562279, 
    0.001442541, 0.001376767, 0.001145918, 0.0006703355, 0.000503657, 
    0.0004071661, 0.0003461873, 0.0002808864, 0.0002415118, 0.0002566103,
  0.001913085, 0.001798001, 0.001708533, 0.0016132, 0.001543768, 0.001483711, 
    0.001329945, 0.0007947728, 0.0004568266, 0.0004297218, 0.0004081008, 
    0.0003184665, 0.0002905878, 0.000278559, 0.0003277237,
  0.001633178, 0.001703297, 0.001558274, 0.00136955, 0.00113656, 
    0.0008154227, 0.0008043157, 0.0007251547, 0.0006392506, 0.0003546642, 
    0.000365503, 0.0004341379, 0.0003590252, 0.0003477817, 0.0002994717,
  0.002244129, 0.00222266, 0.002122467, 0.001873206, 0.001436732, 0.00115347, 
    0.000957703, 0.0007739895, 0.0006820089, 0.0005765987, 0.0004918765, 
    0.0005844228, 0.0005560868, 0.0003416044, 0.0002857016,
  0.002144144, 0.002421296, 0.002421959, 0.002247388, 0.001831129, 
    0.001230372, 0.001139484, 0.0009830699, 0.0007980962, 0.0007052155, 
    0.0006716324, 0.0006828617, 0.0006632307, 0.0005828509, 0.0003830774,
  0.001943731, 0.002149047, 0.00230976, 0.002511868, 0.002349092, 
    0.001725907, 0.001069632, 0.0008949384, 0.0008159694, 0.0007942463, 
    0.0007459503, 0.0007254554, 0.0006944022, 0.000618932, 0.0004291098,
  0.001848371, 0.002057046, 0.002173472, 0.002482216, 0.002503837, 
    0.002387535, 0.001598026, 0.0008226589, 0.0006935589, 0.0007783909, 
    0.0007712726, 0.0007682319, 0.0007167393, 0.0006255656, 0.0004646794,
  0.001714302, 0.001866553, 0.002034185, 0.002253935, 0.0024585, 0.002316548, 
    0.001831174, 0.001589166, 0.001343168, 0.001185896, 0.0009105777, 
    0.0008272383, 0.0007501284, 0.0005578988, 0.0004093362,
  0.001600531, 0.001647695, 0.001741822, 0.001798156, 0.00186022, 
    0.001854109, 0.001645617, 0.001490348, 0.001390704, 0.00133748, 
    0.001055671, 0.0008423261, 0.0006832257, 0.0004739259, 0.0003618706,
  0.001529175, 0.001509314, 0.001507278, 0.001496326, 0.001496301, 
    0.001478788, 0.001392712, 0.001294081, 0.001143751, 0.001110466, 
    0.0009168214, 0.0007406309, 0.0005734049, 0.0003956051, 0.0003145515,
  0.00157983, 0.001494688, 0.001463959, 0.001407707, 0.001388267, 
    0.001296814, 0.001217577, 0.001110805, 0.000714245, 0.0007108227, 
    0.0006824336, 0.0005868374, 0.0004192384, 0.0003079838, 0.0002490108,
  0.001640507, 0.001521979, 0.001446019, 0.001367549, 0.001317969, 
    0.001201844, 0.001035223, 0.000739312, 0.0005262051, 0.0004864633, 
    0.0005240488, 0.0004313963, 0.0003525126, 0.0002930302, 0.0002637699,
  0.001825624, 0.001970233, 0.001884324, 0.001883718, 0.001799833, 
    0.001628638, 0.00154712, 0.001303071, 0.0009683384, 0.0004642591, 
    0.0004352594, 0.0005026374, 0.0004316548, 0.0004116788, 0.0003708834,
  0.001862601, 0.001846504, 0.001741439, 0.001823272, 0.001762599, 
    0.001770384, 0.001655081, 0.001407683, 0.001170302, 0.0007039827, 
    0.0005388567, 0.0005775466, 0.0005175869, 0.0003317908, 0.0003114476,
  0.001569981, 0.001648873, 0.001843566, 0.001655465, 0.001671096, 
    0.001560741, 0.001531624, 0.001438145, 0.001275145, 0.001042104, 
    0.0007752518, 0.0006508117, 0.0005420355, 0.0004558194, 0.0003487959,
  0.001585949, 0.001493275, 0.001521697, 0.001620218, 0.001705728, 
    0.001673565, 0.001160805, 0.001027762, 0.0009809176, 0.0009608493, 
    0.0008045253, 0.0006467485, 0.000580003, 0.0004864785, 0.0003846252,
  0.001615025, 0.001448388, 0.001490684, 0.001525764, 0.001568582, 
    0.001572844, 0.001464087, 0.0006163863, 0.0008258751, 0.0008915081, 
    0.0008943029, 0.0007287987, 0.0006072329, 0.0005186225, 0.0004325546,
  0.001625673, 0.001465708, 0.00150165, 0.00155891, 0.001550337, 0.001482842, 
    0.001335792, 0.001178118, 0.001200199, 0.00129249, 0.001030901, 
    0.0008076152, 0.0006385343, 0.0005469909, 0.0004388696,
  0.001673672, 0.001549075, 0.001592668, 0.001642852, 0.001616161, 
    0.001522337, 0.001357075, 0.001080942, 0.001087925, 0.001296415, 
    0.001111949, 0.0007922358, 0.0006378445, 0.0005505322, 0.0004352457,
  0.00174568, 0.001653248, 0.001759408, 0.001776222, 0.001688324, 
    0.001573767, 0.001372368, 0.00110641, 0.0008940429, 0.001032962, 
    0.0009663888, 0.0007516131, 0.0006340744, 0.0005254907, 0.0004074726,
  0.00181253, 0.001810196, 0.001914657, 0.001905376, 0.001734367, 
    0.001552145, 0.001368537, 0.001050294, 0.0007910948, 0.0007781612, 
    0.0008525105, 0.0007092295, 0.0006165666, 0.0004448923, 0.000311205,
  0.001944996, 0.002070736, 0.002139593, 0.001941261, 0.00174155, 
    0.001548182, 0.001317045, 0.0009662181, 0.0006686266, 0.000520319, 
    0.0007445154, 0.0006573119, 0.0005431154, 0.0003804537, 0.0003145558,
  0.001472957, 0.001779011, 0.001209052, 0.001567627, 0.00131058, 
    0.001256714, 0.001427995, 0.001428504, 0.001394361, 0.0009766886, 
    0.0008474697, 0.0008306035, 0.0006451422, 0.0005696235, 0.0004716694,
  0.001714603, 0.001538663, 0.001405471, 0.00142028, 0.00117447, 0.001272243, 
    0.001426357, 0.001392908, 0.001403623, 0.001212161, 0.000984703, 
    0.0009689364, 0.0009061706, 0.0005844765, 0.0004516602,
  0.001694748, 0.001642511, 0.001836904, 0.001699717, 0.001483096, 
    0.001280977, 0.001463323, 0.001486243, 0.001409121, 0.001193517, 
    0.001064176, 0.001016967, 0.0008955913, 0.000755146, 0.0005445628,
  0.001824847, 0.001774293, 0.001883162, 0.002106875, 0.002219745, 
    0.002168302, 0.001829291, 0.001490546, 0.001317801, 0.001102575, 
    0.0008655043, 0.000812522, 0.0008006607, 0.0007157011, 0.0005687225,
  0.001981687, 0.002015285, 0.002148349, 0.002316578, 0.00250235, 
    0.002611069, 0.002487366, 0.001655164, 0.001166081, 0.0008692613, 
    0.0008170411, 0.0008128854, 0.0007812965, 0.0007417861, 0.0005695479,
  0.00199848, 0.002141278, 0.002343389, 0.002506057, 0.002595386, 
    0.002605857, 0.002483992, 0.002151479, 0.001492013, 0.001099722, 
    0.0008084027, 0.000821439, 0.000761422, 0.000676713, 0.0005264259,
  0.002158254, 0.002429411, 0.002552011, 0.002552578, 0.002568208, 
    0.002433668, 0.002140808, 0.001910331, 0.001545016, 0.001156262, 
    0.0008802086, 0.0006608785, 0.0006879788, 0.000635652, 0.0004923887,
  0.00242378, 0.002620025, 0.002661285, 0.002520511, 0.002448329, 
    0.002188114, 0.001748542, 0.001730407, 0.001422103, 0.0009764711, 
    0.0006948558, 0.0005453053, 0.0006412159, 0.0005553052, 0.0004550355,
  0.002689573, 0.002851184, 0.0027288, 0.002422562, 0.002320482, 0.00188613, 
    0.001523463, 0.001584294, 0.001231129, 0.0007952666, 0.0005794992, 
    0.0005495823, 0.0005819856, 0.0004701304, 0.0003760798,
  0.002989514, 0.003058385, 0.002739742, 0.00231746, 0.002188134, 
    0.001689314, 0.001355228, 0.001429447, 0.0009914414, 0.0005740112, 
    0.0005143, 0.000551186, 0.000520608, 0.0004038553, 0.000340298,
  0.001095661, 0.001275994, 0.001086177, 0.001304415, 0.00129309, 
    0.001303964, 0.001418369, 0.001392831, 0.001387196, 0.001288983, 
    0.001352431, 0.00144989, 0.001342688, 0.001191725, 0.0008221027,
  0.00149339, 0.001679571, 0.001594108, 0.001545159, 0.001437129, 
    0.001500426, 0.001513561, 0.001452901, 0.001369227, 0.001314632, 
    0.001408381, 0.001568717, 0.001475506, 0.0009608893, 0.0007112641,
  0.00199002, 0.002274055, 0.002318193, 0.002098051, 0.001785951, 
    0.001448883, 0.001534747, 0.001478943, 0.001344881, 0.001236083, 
    0.001353433, 0.00133978, 0.001146383, 0.000928239, 0.0006901833,
  0.002323939, 0.002566692, 0.002462053, 0.002235777, 0.002033039, 
    0.001546749, 0.001154212, 0.001201505, 0.001140958, 0.0009854981, 
    0.001000212, 0.0009821854, 0.0009080904, 0.0008624945, 0.0007501879,
  0.002603782, 0.002746935, 0.002461037, 0.002156901, 0.001865491, 
    0.001560786, 0.001392209, 0.0009408469, 0.0009155572, 0.0007535369, 
    0.000726137, 0.0007509474, 0.0007700869, 0.0008265372, 0.0008195732,
  0.002849808, 0.002852487, 0.00253362, 0.002180214, 0.001905473, 
    0.001544772, 0.001336011, 0.001278039, 0.0009975265, 0.0007634833, 
    0.0006175489, 0.0006762415, 0.0007756341, 0.0008630602, 0.0006907039,
  0.002947164, 0.002823755, 0.002581405, 0.002379274, 0.00205864, 
    0.001685799, 0.001426873, 0.001251774, 0.0009956722, 0.0007804204, 
    0.0006382219, 0.0005983187, 0.0006997176, 0.0006943263, 0.000525489,
  0.002922795, 0.002836222, 0.002638303, 0.002541164, 0.002209932, 
    0.001881453, 0.001572386, 0.00134701, 0.0009631332, 0.0007196489, 
    0.0005980846, 0.0005663016, 0.0005894932, 0.0004576457, 0.000424851,
  0.002874884, 0.002878371, 0.002680537, 0.002615247, 0.002356303, 
    0.001996623, 0.001741403, 0.001497311, 0.001052957, 0.0007103377, 
    0.0005609513, 0.0005030886, 0.0004708965, 0.0004122336, 0.000400987,
  0.002907881, 0.003164535, 0.002899154, 0.002707722, 0.002438292, 
    0.002133173, 0.001835675, 0.001613146, 0.001156596, 0.0006502434, 
    0.0004948576, 0.0004822298, 0.0004419921, 0.0003982688, 0.0003824709,
  0.001197677, 0.001367203, 0.001032372, 0.001107849, 0.0009416444, 
    0.0009975081, 0.001224684, 0.001134236, 0.000875624, 0.000538616, 
    0.0006449121, 0.0007816917, 0.0006717227, 0.0006297696, 0.0004957234,
  0.001721779, 0.001514848, 0.001166724, 0.001181929, 0.001033346, 
    0.001287794, 0.001371668, 0.001326521, 0.001028751, 0.0006690388, 
    0.0006384757, 0.0007671493, 0.0006882318, 0.0004462106, 0.0003786619,
  0.001921709, 0.001803494, 0.001793389, 0.001777189, 0.001513432, 
    0.001324677, 0.001639054, 0.001570825, 0.001293765, 0.0007197195, 
    0.0007008008, 0.0007671792, 0.0007075938, 0.000555385, 0.0004338996,
  0.002067305, 0.002056846, 0.002095214, 0.002265992, 0.002199524, 
    0.001982795, 0.001725738, 0.00160148, 0.001517973, 0.000904951, 
    0.000686351, 0.0007691569, 0.0007701837, 0.0005859516, 0.0004596287,
  0.002171226, 0.002197966, 0.002299535, 0.002366993, 0.002374392, 
    0.002600872, 0.002409377, 0.001816165, 0.001620059, 0.001292799, 
    0.0007036676, 0.0007206504, 0.000754267, 0.0006556228, 0.0006397484,
  0.002456779, 0.002649279, 0.002607343, 0.002472697, 0.002441725, 
    0.002634505, 0.002662151, 0.002481996, 0.002265503, 0.001836764, 
    0.0007642262, 0.0007389336, 0.000697626, 0.0005669484, 0.0004830077,
  0.002513648, 0.0025047, 0.002700668, 0.002863623, 0.002417533, 0.002569324, 
    0.002571733, 0.002655427, 0.002439778, 0.002148153, 0.001169086, 
    0.0007178773, 0.0006995433, 0.0004814119, 0.0003938702,
  0.002556482, 0.00255252, 0.00252687, 0.002731379, 0.002422567, 0.002511101, 
    0.002516737, 0.002663131, 0.00254026, 0.002317568, 0.001612485, 
    0.0008649575, 0.0006861278, 0.0004957649, 0.0003497594,
  0.00256506, 0.002492955, 0.002419111, 0.002630481, 0.002548064, 
    0.002670312, 0.002533951, 0.002581162, 0.002553971, 0.002404191, 
    0.001824761, 0.001113932, 0.0007553747, 0.0004515079, 0.0003721931,
  0.00251692, 0.002563526, 0.002627002, 0.002635289, 0.002672142, 
    0.002579404, 0.0025868, 0.002540952, 0.002559327, 0.002475011, 
    0.002007403, 0.001320984, 0.0008820249, 0.0005468515, 0.0004242188,
  0.001197214, 0.001355147, 0.001491584, 0.001934114, 0.00198742, 
    0.002089821, 0.002211505, 0.001881576, 0.0009305906, 0.0004042655, 
    0.0004558269, 0.0005422513, 0.0003705064, 0.0002797733, 0.0002449645,
  0.001444982, 0.001636731, 0.001857911, 0.002040151, 0.001918783, 
    0.002017945, 0.002123126, 0.001945465, 0.001542759, 0.0006650097, 
    0.0004300236, 0.0005784177, 0.0004907231, 0.0002291245, 0.0001887532,
  0.001857781, 0.001854562, 0.002111173, 0.002233587, 0.001925885, 
    0.001724076, 0.002024422, 0.002051316, 0.002117196, 0.001286299, 
    0.0007464121, 0.0006227792, 0.000531142, 0.0004808127, 0.0003642019,
  0.002008668, 0.002079617, 0.002058479, 0.002017011, 0.002141117, 
    0.002001902, 0.001789706, 0.001606881, 0.002180826, 0.002011778, 
    0.001197272, 0.0007688208, 0.0005788789, 0.000478075, 0.0004719683,
  0.002113499, 0.002106259, 0.002080799, 0.002016276, 0.001996096, 
    0.002094585, 0.002271587, 0.001854136, 0.002010396, 0.00224562, 
    0.001676544, 0.001250702, 0.0007151208, 0.000534448, 0.0005765051,
  0.002174111, 0.002215918, 0.002083083, 0.002018709, 0.002023786, 
    0.002086422, 0.002247155, 0.002355668, 0.002258444, 0.002310661, 
    0.002037317, 0.001702153, 0.001181243, 0.0006958183, 0.0005215818,
  0.002173523, 0.002286852, 0.002102131, 0.002114714, 0.002091902, 
    0.002164953, 0.002190666, 0.002324168, 0.002300048, 0.002278452, 
    0.002258629, 0.001897046, 0.001505223, 0.0009811496, 0.0005974316,
  0.002292191, 0.002376874, 0.002315252, 0.002320912, 0.002274765, 
    0.002327535, 0.002358803, 0.002377757, 0.002336503, 0.002260418, 
    0.00226263, 0.001998618, 0.001713606, 0.001254491, 0.0007880938,
  0.002539722, 0.002599395, 0.002612405, 0.002613745, 0.002680936, 
    0.002548986, 0.002605425, 0.00253823, 0.002409807, 0.002368011, 
    0.002316309, 0.002058317, 0.001847517, 0.001474163, 0.000988109,
  0.002650151, 0.002751037, 0.002951506, 0.002653825, 0.002591166, 
    0.002533094, 0.002527143, 0.002402727, 0.002417913, 0.002294425, 
    0.002311699, 0.002207031, 0.001895325, 0.001588009, 0.001171254,
  0.001593446, 0.001691067, 0.001627348, 0.001743715, 0.001767036, 
    0.001825449, 0.001870709, 0.001614079, 0.001296843, 0.0006878494, 
    0.000442366, 0.0004626252, 0.0002522281, 0.0002510417, 0.000220084,
  0.001818534, 0.00173924, 0.001774961, 0.001735633, 0.001558744, 
    0.001641261, 0.001563285, 0.001719643, 0.001690448, 0.001411006, 
    0.0008157885, 0.0007273052, 0.0005934549, 0.0003671588, 0.0002654229,
  0.001879734, 0.001810619, 0.001841015, 0.001796501, 0.001617912, 
    0.001274542, 0.001647446, 0.001722952, 0.001776667, 0.001719582, 
    0.001455952, 0.001190694, 0.0009654665, 0.0008246428, 0.0005868103,
  0.001908798, 0.00185153, 0.001802443, 0.001708305, 0.001816148, 
    0.001722345, 0.001529552, 0.001390313, 0.001492729, 0.001570522, 
    0.001605996, 0.001513018, 0.001336847, 0.001154325, 0.0009832438,
  0.001929536, 0.001846179, 0.001827133, 0.001834507, 0.001879059, 
    0.001934477, 0.002040659, 0.001764804, 0.001732081, 0.001675839, 
    0.001821429, 0.001863404, 0.001739217, 0.001472497, 0.001237363,
  0.001968476, 0.001928445, 0.001980172, 0.002009985, 0.002073796, 
    0.002162913, 0.002205192, 0.002342806, 0.002311826, 0.002250276, 
    0.002230828, 0.002067134, 0.002044392, 0.001881009, 0.001584682,
  0.002182157, 0.002203045, 0.002241403, 0.002288234, 0.002347143, 0.0023923, 
    0.00244018, 0.002537569, 0.002573333, 0.002493907, 0.002400056, 
    0.002230647, 0.002167428, 0.002080029, 0.001906935,
  0.0023926, 0.002449053, 0.002486793, 0.00260009, 0.002634332, 0.002669673, 
    0.002718527, 0.00282168, 0.002843264, 0.002788336, 0.002733844, 
    0.002505794, 0.002389273, 0.00227824, 0.002068375,
  0.002577102, 0.002662159, 0.002796532, 0.002858835, 0.00295013, 
    0.002887518, 0.002928641, 0.002991127, 0.003020156, 0.002986613, 
    0.00291494, 0.002767504, 0.002632319, 0.002370545, 0.002136943,
  0.002814104, 0.002919601, 0.003020798, 0.003077378, 0.00307386, 
    0.003098425, 0.003105165, 0.003088806, 0.003116458, 0.003083678, 
    0.003030586, 0.002930662, 0.002808811, 0.002522489, 0.002062878,
  0.001772866, 0.001402606, 0.001040889, 0.0009296859, 0.0007640691, 
    0.0007911069, 0.0009378688, 0.00104194, 0.001157236, 0.001084746, 
    0.001168077, 0.001255522, 0.00121886, 0.001192004, 0.00137395,
  0.001736543, 0.001541859, 0.001228013, 0.001035672, 0.0007643104, 
    0.0008898039, 0.001179414, 0.001225636, 0.001265939, 0.001255768, 
    0.001289026, 0.001513288, 0.001686879, 0.001609037, 0.001550981,
  0.001869081, 0.001685846, 0.001511011, 0.001246269, 0.0009318269, 
    0.0006911602, 0.00110331, 0.001242955, 0.001455963, 0.001579626, 
    0.001742211, 0.001980284, 0.002140824, 0.002143161, 0.002074207,
  0.002147491, 0.002056505, 0.001972743, 0.001874454, 0.001651724, 
    0.001234772, 0.001225879, 0.00149709, 0.001910407, 0.002133588, 
    0.002346538, 0.002487891, 0.00241279, 0.002305752, 0.002216694,
  0.002233656, 0.002138877, 0.002086326, 0.002061168, 0.002076982, 
    0.002139559, 0.002174383, 0.002019189, 0.002153972, 0.002416911, 
    0.002718423, 0.002677288, 0.002523999, 0.002411791, 0.002313168,
  0.002246875, 0.002210691, 0.002178535, 0.002190467, 0.002251314, 
    0.002329287, 0.00244531, 0.002550458, 0.002771603, 0.002989307, 
    0.002934063, 0.002619227, 0.002489393, 0.002391609, 0.00224623,
  0.002278314, 0.002305115, 0.002326653, 0.00233893, 0.002483877, 
    0.002593469, 0.002734248, 0.002928646, 0.003165699, 0.00309193, 
    0.002637065, 0.002453575, 0.002350894, 0.002242552, 0.002160781,
  0.002406995, 0.002447285, 0.00250544, 0.002600465, 0.00272791, 0.002855574, 
    0.003012174, 0.003180551, 0.0031747, 0.002580883, 0.002361587, 
    0.002230428, 0.002139952, 0.002049289, 0.002010199,
  0.002467615, 0.002598133, 0.002694768, 0.002779745, 0.002903272, 
    0.003030662, 0.003233615, 0.003239531, 0.002593408, 0.002190389, 
    0.002061267, 0.001945863, 0.001852684, 0.001822913, 0.001830328,
  0.002666582, 0.00277438, 0.002893725, 0.003008143, 0.00313591, 0.003286332, 
    0.00330771, 0.002538147, 0.002054518, 0.001770506, 0.001785299, 
    0.001709125, 0.001665755, 0.00166437, 0.001619376,
  0.001750855, 0.001598393, 0.001276566, 0.0010787, 0.0008386324, 
    0.0006914485, 0.000743359, 0.0006351423, 0.0005809816, 0.0005116706, 
    0.0006020249, 0.0008594726, 0.00114534, 0.001327774, 0.00105734,
  0.001935506, 0.001870246, 0.001501591, 0.001191292, 0.000827459, 
    0.0007384188, 0.0008289882, 0.0007131753, 0.0006897079, 0.0006646268, 
    0.0007517918, 0.001192625, 0.0014953, 0.001152159, 0.0008672056,
  0.002008689, 0.001959585, 0.001848724, 0.001527324, 0.0009636477, 
    0.000724673, 0.0009610312, 0.0009907881, 0.000952001, 0.0009066963, 
    0.001081674, 0.001458096, 0.001435402, 0.001134346, 0.00085743,
  0.00214138, 0.002200679, 0.00218685, 0.002100584, 0.001696112, 0.001036651, 
    0.0008593376, 0.0009763405, 0.001167889, 0.001210758, 0.001509643, 
    0.001658004, 0.001371972, 0.001209727, 0.0009835846,
  0.002221899, 0.002201303, 0.002205901, 0.002198073, 0.00219429, 
    0.002138321, 0.001683887, 0.001172503, 0.00112381, 0.001525934, 
    0.001929331, 0.001758089, 0.001523187, 0.001386886, 0.001219137,
  0.002220121, 0.002233843, 0.002252691, 0.002292186, 0.002302935, 
    0.002297713, 0.002277185, 0.002068288, 0.001869838, 0.002050433, 
    0.002138217, 0.001881287, 0.001712807, 0.001516737, 0.001267293,
  0.002249029, 0.002289985, 0.002272281, 0.002264506, 0.00227442, 
    0.002276799, 0.00230639, 0.002360515, 0.002369057, 0.002398715, 
    0.002223886, 0.001959434, 0.001762885, 0.001528219, 0.001278595,
  0.002232117, 0.002268502, 0.002265068, 0.002267782, 0.002305454, 
    0.002320343, 0.002362769, 0.002472159, 0.002454048, 0.00239874, 
    0.002203712, 0.001948179, 0.001721602, 0.001470249, 0.001251808,
  0.002293395, 0.002256599, 0.002267646, 0.002310849, 0.002351591, 
    0.002442947, 0.002492506, 0.002531758, 0.002554247, 0.002427534, 
    0.002221591, 0.001932882, 0.00170089, 0.001430484, 0.001234371,
  0.002376693, 0.002321689, 0.002294132, 0.002330602, 0.002461746, 
    0.002545764, 0.002508414, 0.00254305, 0.002509065, 0.002256683, 
    0.002154258, 0.001881943, 0.001610451, 0.001354296, 0.001160674,
  0.001960485, 0.001944831, 0.001922286, 0.001962247, 0.001853736, 
    0.001700818, 0.001652761, 0.001358963, 0.001062729, 0.0006040452, 
    0.0004800328, 0.0005064311, 0.0004173317, 0.0003749656, 0.0003461389,
  0.002023904, 0.002065046, 0.00205142, 0.002074284, 0.001913461, 
    0.001730885, 0.001712736, 0.001403375, 0.001077349, 0.0008645827, 
    0.0007105546, 0.0007028715, 0.0006466308, 0.0004630618, 0.0004558688,
  0.002089819, 0.002147558, 0.002239011, 0.002253696, 0.002099026, 
    0.001667182, 0.001758157, 0.001607037, 0.001173684, 0.001072775, 
    0.001042602, 0.001005401, 0.0009466298, 0.0009817573, 0.0009528702,
  0.002258996, 0.002286192, 0.002377956, 0.002457297, 0.002500994, 
    0.002067391, 0.001671364, 0.001525894, 0.001414592, 0.001376944, 
    0.001361405, 0.001335749, 0.001397205, 0.001263701, 0.001017184,
  0.002395622, 0.002437117, 0.002530087, 0.002629683, 0.002657337, 
    0.002711355, 0.002365196, 0.001574322, 0.001532683, 0.00166854, 
    0.001913792, 0.001804035, 0.001565951, 0.001140918, 0.001008547,
  0.00267457, 0.002722523, 0.002775104, 0.002765519, 0.002702647, 
    0.002599235, 0.002657761, 0.002396017, 0.002174356, 0.002099049, 
    0.002228572, 0.001974961, 0.001402621, 0.001120014, 0.00103162,
  0.003043597, 0.003010023, 0.002921917, 0.002782535, 0.00268445, 
    0.002531709, 0.002439101, 0.002552352, 0.002283718, 0.002372294, 
    0.002075938, 0.001508039, 0.001124136, 0.0009631194, 0.000906623,
  0.003321502, 0.003216061, 0.003025287, 0.002769663, 0.002695115, 
    0.002425398, 0.002442812, 0.002523849, 0.0025434, 0.002180337, 
    0.001476662, 0.001073287, 0.000883735, 0.0007847676, 0.0007593411,
  0.003524161, 0.003257733, 0.00304096, 0.002846039, 0.002643629, 
    0.002516338, 0.00241677, 0.002591808, 0.002289978, 0.001768746, 
    0.001326027, 0.0008870054, 0.0007161392, 0.0006264119, 0.0006236268,
  0.00342256, 0.003314827, 0.003068473, 0.002751345, 0.002627253, 
    0.002377786, 0.002450461, 0.002154013, 0.001714137, 0.001257628, 
    0.001129085, 0.0008380304, 0.0006295195, 0.0005318927, 0.0005016471,
  0.001588472, 0.001774826, 0.001774676, 0.002098376, 0.002137193, 
    0.002313338, 0.002519681, 0.002559268, 0.002417641, 0.001973553, 
    0.001568504, 0.001355379, 0.0009493666, 0.0007248968, 0.0005014867,
  0.001993761, 0.002074482, 0.002314406, 0.002575756, 0.002544312, 
    0.002740597, 0.00286771, 0.002747931, 0.002487748, 0.00196996, 
    0.001706284, 0.00154847, 0.001298228, 0.0008348296, 0.0006535889,
  0.002533752, 0.002765682, 0.002863808, 0.003004603, 0.003048887, 
    0.002982263, 0.002962776, 0.002834182, 0.002492107, 0.002057717, 
    0.001883059, 0.001708569, 0.001540821, 0.001362951, 0.00107536,
  0.002824835, 0.003230144, 0.003255719, 0.003272318, 0.003347853, 
    0.003313923, 0.00302131, 0.002759036, 0.002418464, 0.002150357, 
    0.001940264, 0.001800891, 0.001734328, 0.00160203, 0.001418969,
  0.003305302, 0.003396617, 0.003404716, 0.003481546, 0.003465274, 
    0.003399444, 0.003279729, 0.002640268, 0.002428049, 0.00219665, 
    0.00223483, 0.002159958, 0.001997365, 0.001790676, 0.001569078,
  0.003579899, 0.003648521, 0.003665603, 0.003607717, 0.003556737, 
    0.003409417, 0.003229641, 0.00297577, 0.002773766, 0.00254808, 
    0.002369616, 0.002268093, 0.002122728, 0.001876879, 0.001468046,
  0.003941685, 0.003963031, 0.003864956, 0.003663966, 0.003556926, 
    0.003322246, 0.003119535, 0.002961068, 0.002649402, 0.002420326, 
    0.002252298, 0.002257218, 0.002034086, 0.001622718, 0.001104079,
  0.004009501, 0.004026616, 0.003927781, 0.00367785, 0.003495376, 
    0.003248008, 0.003031377, 0.00288851, 0.002682655, 0.002529255, 
    0.002433971, 0.002202735, 0.001754963, 0.00111715, 0.0007829082,
  0.004198727, 0.004144677, 0.003959814, 0.003629117, 0.003351001, 
    0.003184733, 0.003032312, 0.002815964, 0.002619787, 0.002578524, 
    0.002474533, 0.001795717, 0.001100163, 0.0007645632, 0.0006283305,
  0.004123782, 0.003941381, 0.003715003, 0.003438132, 0.003262762, 
    0.003083427, 0.002856343, 0.002720001, 0.002718594, 0.002464062, 
    0.001949873, 0.001120284, 0.0007661739, 0.0005443532, 0.000448117,
  0.001047509, 0.001288099, 0.001364413, 0.001621857, 0.001772813, 
    0.002087987, 0.002313684, 0.002383074, 0.002251777, 0.002039941, 
    0.001972315, 0.002053547, 0.001888582, 0.001966638, 0.001907242,
  0.00155277, 0.001677634, 0.00176118, 0.001797771, 0.001927296, 0.002352315, 
    0.002433396, 0.002341313, 0.002240142, 0.002073635, 0.002005829, 
    0.002063125, 0.002170867, 0.0022024, 0.002143758,
  0.001928178, 0.002157965, 0.002280511, 0.002163662, 0.002415063, 
    0.002338186, 0.00255738, 0.002413387, 0.002272636, 0.002170541, 
    0.002256514, 0.002391959, 0.002598554, 0.002618704, 0.002463378,
  0.002178746, 0.002400769, 0.002566375, 0.002735169, 0.00270949, 
    0.002763308, 0.002640874, 0.002546361, 0.002448086, 0.002411182, 
    0.002545675, 0.002715121, 0.002784051, 0.002753249, 0.002246657,
  0.00243137, 0.002550601, 0.00269103, 0.002815981, 0.002905346, 0.002942261, 
    0.002964036, 0.002597491, 0.002552524, 0.002652856, 0.002830755, 
    0.002871684, 0.002896295, 0.002763978, 0.002056276,
  0.002632642, 0.002747111, 0.002889529, 0.002976718, 0.003079781, 
    0.003098352, 0.003105533, 0.00304594, 0.002954113, 0.002966054, 
    0.002915557, 0.002891133, 0.002915306, 0.002615465, 0.001741265,
  0.002952303, 0.003038112, 0.003118195, 0.00315968, 0.003171318, 
    0.003195748, 0.003171562, 0.00311522, 0.003036616, 0.00290769, 
    0.002825963, 0.002857188, 0.002886249, 0.002184664, 0.001261524,
  0.00314072, 0.003173252, 0.003248189, 0.003274191, 0.003294231, 
    0.003272262, 0.003188645, 0.003145796, 0.003039936, 0.002919001, 
    0.002837927, 0.002955772, 0.002657921, 0.00144657, 0.0007337006,
  0.003322209, 0.003405735, 0.003460829, 0.003450434, 0.003370269, 
    0.003281274, 0.003248629, 0.003158733, 0.003044214, 0.002947619, 
    0.002994221, 0.0029268, 0.001880427, 0.0007447009, 0.0004806179,
  0.003526863, 0.003518667, 0.003521134, 0.003416957, 0.003350389, 
    0.003273872, 0.003158616, 0.002982339, 0.002939658, 0.002894537, 
    0.003000979, 0.002452421, 0.000940351, 0.0004665662, 0.0003691338,
  0.0008801502, 0.001001508, 0.001005879, 0.001090868, 0.0009811004, 
    0.000972425, 0.001227312, 0.001324864, 0.001516275, 0.00166931, 
    0.001788269, 0.00193053, 0.001944254, 0.002003195, 0.002062151,
  0.001376716, 0.001422939, 0.001326226, 0.001211518, 0.001093285, 
    0.001433928, 0.001748564, 0.001787885, 0.001949251, 0.002034108, 
    0.002081443, 0.002112863, 0.002041577, 0.00202607, 0.002239654,
  0.001864826, 0.001947779, 0.002004821, 0.001951326, 0.002033918, 
    0.001938231, 0.00213525, 0.002188836, 0.002163102, 0.002110056, 
    0.00203874, 0.002074662, 0.002242444, 0.002565322, 0.0028116,
  0.00205062, 0.002190684, 0.00228543, 0.002327912, 0.002315867, 0.002290588, 
    0.002235152, 0.00231006, 0.002246781, 0.002025803, 0.002142826, 
    0.00236432, 0.002674421, 0.002882431, 0.002894473,
  0.002244209, 0.002288918, 0.002353252, 0.002387139, 0.002422053, 
    0.002492019, 0.002545631, 0.002298847, 0.00223646, 0.002386164, 
    0.002690165, 0.002816898, 0.002932451, 0.002972029, 0.002881972,
  0.002382588, 0.002430358, 0.002448343, 0.002458596, 0.002532599, 
    0.00264489, 0.002728842, 0.002765644, 0.002772581, 0.002846011, 
    0.002940095, 0.002998096, 0.003011358, 0.003007712, 0.002717651,
  0.002593942, 0.002608728, 0.002605445, 0.002655468, 0.002749395, 
    0.002823302, 0.002888463, 0.002967464, 0.003020797, 0.003051804, 
    0.003072675, 0.003072312, 0.003051559, 0.002990696, 0.00232737,
  0.002772795, 0.002772296, 0.002810969, 0.002909334, 0.003014968, 
    0.003078501, 0.003121079, 0.00316237, 0.003179231, 0.003173402, 
    0.003151679, 0.003124431, 0.003108229, 0.002801764, 0.002010711,
  0.003011542, 0.003040434, 0.003121624, 0.003163913, 0.003181742, 
    0.003197023, 0.003217041, 0.003232011, 0.003248667, 0.003251657, 
    0.003241901, 0.003186053, 0.003092036, 0.002529621, 0.001733446,
  0.003368257, 0.003356701, 0.003371887, 0.003319924, 0.00327297, 
    0.003251001, 0.003243379, 0.003238443, 0.003269994, 0.003296311, 
    0.00326756, 0.003222377, 0.002904851, 0.002252904, 0.001523831,
  0.0008100203, 0.0008952832, 0.0009323322, 0.0009914668, 0.000906995, 
    0.0009080417, 0.001018886, 0.0009500477, 0.0009801154, 0.001035106, 
    0.001167748, 0.001277723, 0.001377032, 0.001504743, 0.001611394,
  0.001318794, 0.001185859, 0.001060734, 0.001000163, 0.0008580679, 
    0.001087316, 0.001245199, 0.001292281, 0.001341114, 0.00141453, 
    0.001519589, 0.001638304, 0.001749614, 0.001778337, 0.001875827,
  0.001822979, 0.00195242, 0.001913018, 0.001717122, 0.001301007, 0.00127345, 
    0.001652239, 0.00174339, 0.001764977, 0.001760116, 0.001777395, 
    0.001863443, 0.001962574, 0.002045486, 0.002153202,
  0.001962075, 0.002059679, 0.002108631, 0.002171325, 0.002126143, 
    0.001797347, 0.00169773, 0.00191704, 0.001994479, 0.002028047, 
    0.002002182, 0.001957507, 0.002055024, 0.002139177, 0.002250352,
  0.002171496, 0.002181932, 0.002216537, 0.002272906, 0.002268782, 
    0.002350881, 0.002304538, 0.001991747, 0.001933358, 0.00204678, 
    0.0022561, 0.002128389, 0.002156018, 0.002294016, 0.002295026,
  0.002329641, 0.002347745, 0.002342887, 0.002312512, 0.002310451, 
    0.002319652, 0.002393399, 0.002430407, 0.002275598, 0.002286099, 
    0.00233805, 0.002286935, 0.002309131, 0.00241286, 0.002507863,
  0.002494061, 0.002489203, 0.002481912, 0.002431952, 0.002423706, 
    0.002406357, 0.002424648, 0.002516962, 0.002557571, 0.002490954, 
    0.002443166, 0.002411402, 0.00247475, 0.002541267, 0.002629094,
  0.002472667, 0.002486888, 0.002470376, 0.002502193, 0.002547694, 
    0.002547806, 0.002555714, 0.002581456, 0.002625669, 0.002591572, 
    0.002536954, 0.002517168, 0.002531239, 0.002561337, 0.002665637,
  0.002394536, 0.002415875, 0.002458399, 0.002570771, 0.00270569, 0.00277769, 
    0.002794588, 0.002780998, 0.002733167, 0.002723972, 0.002725287, 
    0.002636716, 0.002655662, 0.002669635, 0.002716418,
  0.002070188, 0.002079196, 0.002145875, 0.002305816, 0.002471309, 
    0.002668273, 0.002820028, 0.002950295, 0.002997495, 0.002950223, 
    0.002946792, 0.002926121, 0.002892, 0.002861783, 0.002836911,
  0.0008246755, 0.0008893264, 0.0009353479, 0.0009928164, 0.000849131, 
    0.0007936718, 0.0008583909, 0.0007366468, 0.0006071838, 0.000566079, 
    0.0005892422, 0.0006184601, 0.0005825044, 0.0005804308, 0.0005868389,
  0.00115782, 0.0009875314, 0.0009330808, 0.0008850403, 0.0007544952, 
    0.0009574367, 0.001034153, 0.0009207142, 0.0007377438, 0.0006556678, 
    0.000680143, 0.0007400432, 0.0007384444, 0.0006670719, 0.0007107087,
  0.001750788, 0.001715117, 0.001567614, 0.00129312, 0.0008112721, 
    0.0007363309, 0.001214637, 0.001237728, 0.001069593, 0.0008299568, 
    0.0008559303, 0.0008756873, 0.0008593259, 0.0008701875, 0.0009202625,
  0.00204233, 0.002035413, 0.002008862, 0.002005013, 0.001857375, 
    0.001129926, 0.001002416, 0.001371403, 0.001525366, 0.00139511, 
    0.00125346, 0.001249254, 0.001270684, 0.00133849, 0.001366016,
  0.00210382, 0.002213388, 0.002242836, 0.002225348, 0.002178255, 
    0.002170708, 0.001757788, 0.001321546, 0.001351233, 0.001554393, 
    0.001762245, 0.001768813, 0.001770743, 0.00180062, 0.001786079,
  0.001828849, 0.001962623, 0.002151127, 0.002257589, 0.002308823, 
    0.002370862, 0.002430414, 0.002232893, 0.001781031, 0.001753898, 
    0.001806478, 0.00195483, 0.002003382, 0.002033291, 0.002040034,
  0.001535335, 0.001520672, 0.001516003, 0.001539525, 0.001635645, 
    0.001750484, 0.001887824, 0.002078247, 0.002196247, 0.002089617, 
    0.002171755, 0.002207063, 0.002241612, 0.00223625, 0.002180899,
  0.00141805, 0.001344841, 0.001306063, 0.001294556, 0.001356332, 
    0.001485929, 0.001649091, 0.001846832, 0.002008264, 0.002018386, 
    0.002159987, 0.002205206, 0.002268927, 0.002299136, 0.002277666,
  0.001366389, 0.001264412, 0.001173152, 0.001096256, 0.001092338, 
    0.00118924, 0.0014406, 0.001733526, 0.001926292, 0.002048135, 
    0.002196193, 0.002223044, 0.002236057, 0.002224038, 0.002214779,
  0.001321925, 0.001205912, 0.001120222, 0.001042289, 0.000976963, 
    0.0009573312, 0.001009081, 0.001107625, 0.001583638, 0.001864772, 
    0.002168621, 0.002300651, 0.002141848, 0.002223133, 0.002283322,
  0.0009777204, 0.0009922357, 0.0010096, 0.001068382, 0.001030131, 
    0.001039245, 0.001094834, 0.0009636332, 0.0008454649, 0.0007253094, 
    0.000675974, 0.0007171768, 0.0006091589, 0.0005621969, 0.0004727418,
  0.001381529, 0.001135869, 0.001037232, 0.0009962376, 0.00089325, 
    0.001083333, 0.001125187, 0.001050117, 0.0008904628, 0.0008022611, 
    0.0007942883, 0.0008191938, 0.0007305196, 0.0005501655, 0.0004726195,
  0.002116481, 0.002057527, 0.00184094, 0.001445352, 0.001013503, 
    0.0008742471, 0.001190825, 0.001174345, 0.001066863, 0.0008577434, 
    0.0009086686, 0.0008512791, 0.0007646254, 0.0006441908, 0.0005369551,
  0.001828266, 0.001939877, 0.002087782, 0.002243678, 0.002014847, 
    0.001179744, 0.0009624924, 0.001248945, 0.00127586, 0.001171617, 
    0.001045071, 0.0009954328, 0.0008682815, 0.0008051965, 0.0006746216,
  0.001505742, 0.001551537, 0.001715002, 0.001870686, 0.002099599, 
    0.002181376, 0.001514756, 0.001036088, 0.0009970228, 0.001227543, 
    0.001413033, 0.001274461, 0.001064967, 0.0008964101, 0.0007596684,
  0.001454884, 0.00136734, 0.001414689, 0.001627589, 0.001786879, 
    0.001902737, 0.002055048, 0.001804877, 0.001410361, 0.001249282, 
    0.001383301, 0.001498165, 0.001537835, 0.00149346, 0.001397758,
  0.001455379, 0.001354475, 0.001291382, 0.0012865, 0.001313004, 0.001368963, 
    0.001548057, 0.001668056, 0.00177021, 0.001702451, 0.001732766, 
    0.001686848, 0.001707501, 0.001742187, 0.001761489,
  0.001525907, 0.001383812, 0.001265232, 0.001229882, 0.00118503, 
    0.001212742, 0.001176248, 0.001146552, 0.00117367, 0.001080053, 
    0.001017958, 0.0009365601, 0.000913711, 0.0009225557, 0.0009751134,
  0.00156496, 0.001426305, 0.001292589, 0.001183335, 0.001127522, 
    0.001079778, 0.001086587, 0.001059863, 0.000954217, 0.0008592362, 
    0.0009622464, 0.0008682274, 0.0008229208, 0.000777343, 0.0008224346,
  0.001553982, 0.00141275, 0.001270753, 0.001162036, 0.001080406, 
    0.0009893312, 0.0007876516, 0.0006332809, 0.0006365567, 0.0006158061, 
    0.0007633237, 0.0007142038, 0.000719753, 0.0007774472, 0.0009182403,
  0.001031637, 0.001078921, 0.001053107, 0.001071543, 0.0010248, 0.001063435, 
    0.00109149, 0.0010663, 0.0009849933, 0.0008165739, 0.0007795118, 
    0.0008028967, 0.0007651369, 0.0007258549, 0.0007035244,
  0.001647054, 0.001459637, 0.001228868, 0.001101321, 0.0009372259, 
    0.001095976, 0.001144442, 0.001108415, 0.001043928, 0.0009636599, 
    0.0009318426, 0.0008996411, 0.0008398609, 0.0007163387, 0.0006910202,
  0.002163815, 0.002196257, 0.002064571, 0.001769975, 0.001147023, 
    0.0009718311, 0.001240498, 0.00122292, 0.00117427, 0.001062473, 
    0.001067672, 0.0009926135, 0.0009017125, 0.0008322666, 0.0007494094,
  0.00211809, 0.001969862, 0.001934448, 0.002023401, 0.002041718, 
    0.001328098, 0.001071227, 0.001354568, 0.001380673, 0.00129725, 
    0.001250321, 0.001154025, 0.001035107, 0.0009432147, 0.0008435753,
  0.001977896, 0.001828498, 0.001735397, 0.001612781, 0.001658326, 
    0.002049331, 0.001693933, 0.001211065, 0.001186787, 0.001300899, 
    0.001458611, 0.001359443, 0.001238257, 0.001092543, 0.0009915996,
  0.001832272, 0.001710116, 0.001634319, 0.001548423, 0.001420212, 
    0.001420081, 0.001608435, 0.001719164, 0.00154898, 0.001276452, 
    0.001286283, 0.001311247, 0.001257947, 0.001224568, 0.001171076,
  0.001691649, 0.001628057, 0.001557416, 0.001407107, 0.001329884, 
    0.001324632, 0.001302527, 0.001317781, 0.00135855, 0.001418766, 
    0.001439241, 0.00143674, 0.001434823, 0.001353435, 0.001163656,
  0.001606051, 0.001522141, 0.001402568, 0.001309756, 0.001204515, 
    0.001178665, 0.001118663, 0.001075575, 0.000999607, 0.0008793192, 
    0.0009347954, 0.0008883191, 0.0008943662, 0.000872609, 0.0008111453,
  0.001498174, 0.001397945, 0.001290293, 0.001151064, 0.001021745, 
    0.0009367861, 0.0008688696, 0.000786986, 0.0006844208, 0.0006530259, 
    0.00070133, 0.0006297463, 0.0006832753, 0.000627748, 0.0005855297,
  0.001364119, 0.001203044, 0.001104122, 0.0009486931, 0.0007883804, 
    0.0006518768, 0.0005320814, 0.0004878597, 0.000485826, 0.00046201, 
    0.0005057855, 0.0004639231, 0.0004536689, 0.000435992, 0.0005245095,
  0.001124005, 0.001184177, 0.001127027, 0.001099218, 0.001008004, 
    0.0009615598, 0.001018064, 0.0009604082, 0.0008896826, 0.0006474645, 
    0.0007011953, 0.0007173775, 0.0006238603, 0.0005524, 0.0005091423,
  0.001798441, 0.001595143, 0.001356591, 0.001152974, 0.001026137, 
    0.001073494, 0.001093523, 0.0009982253, 0.0008828876, 0.0007495491, 
    0.0007935766, 0.0008337779, 0.0007726974, 0.0005935198, 0.0005811156,
  0.001956433, 0.002040443, 0.00205877, 0.001752255, 0.001196175, 
    0.0009549785, 0.001224809, 0.001162212, 0.001020735, 0.0007820245, 
    0.0008836493, 0.0008749249, 0.0008097648, 0.000742314, 0.0006470495,
  0.001730715, 0.001766109, 0.001990241, 0.002212265, 0.002112199, 
    0.001267125, 0.001042771, 0.001296148, 0.001288361, 0.001080241, 
    0.0009892273, 0.0009379369, 0.0008491293, 0.0008393113, 0.0007632701,
  0.001538926, 0.001616457, 0.001701765, 0.001854641, 0.002046308, 
    0.002057023, 0.00146854, 0.001117792, 0.001075643, 0.001204158, 
    0.001235842, 0.001106623, 0.0009858847, 0.0009102043, 0.000831659,
  0.001530808, 0.00147338, 0.001381856, 0.001428318, 0.001584399, 
    0.001710104, 0.001750985, 0.001626036, 0.001379075, 0.001274117, 
    0.001270792, 0.001224259, 0.001116193, 0.001019192, 0.0009187168,
  0.001501546, 0.001317317, 0.001125773, 0.001086937, 0.001156996, 
    0.001268087, 0.001361523, 0.001413152, 0.001329862, 0.001311294, 
    0.001302114, 0.00124221, 0.001215045, 0.001134148, 0.0010527,
  0.001435433, 0.001199428, 0.0009967335, 0.0008954843, 0.0008624331, 
    0.0008739527, 0.0008782568, 0.000867256, 0.0007282804, 0.0007116045, 
    0.0009463611, 0.0009955278, 0.001029279, 0.001011559, 0.0009894335,
  0.001438805, 0.001149261, 0.0009552732, 0.0008380873, 0.0007513899, 
    0.0006829017, 0.0006340738, 0.0005548009, 0.0004903829, 0.0004995267, 
    0.0006013149, 0.000595572, 0.0006433064, 0.0006683168, 0.0007205412,
  0.001531761, 0.001145021, 0.0009218964, 0.0007552583, 0.0006606437, 
    0.0005409879, 0.0004384156, 0.000381423, 0.0003593895, 0.0003951254, 
    0.0003990389, 0.0003586819, 0.0003600371, 0.0004120469, 0.0004813702,
  0.001513367, 0.001459134, 0.001321708, 0.001280318, 0.001092225, 
    0.001004572, 0.001009953, 0.0009071754, 0.0008565169, 0.0006424931, 
    0.000631003, 0.000641009, 0.000464669, 0.0004050213, 0.0003295533,
  0.00184346, 0.001682404, 0.001508933, 0.001379783, 0.001112532, 
    0.001211294, 0.001195704, 0.00102517, 0.0008816154, 0.0008020084, 
    0.0007408521, 0.0007720058, 0.0006690788, 0.0004420313, 0.0003696006,
  0.002231688, 0.002012162, 0.001893591, 0.001679561, 0.001362755, 
    0.00110365, 0.001323289, 0.00127458, 0.001066745, 0.0008352044, 
    0.0008961793, 0.0008616488, 0.0007546059, 0.0006460577, 0.0004815561,
  0.00235878, 0.002035244, 0.001769686, 0.001699915, 0.001886989, 0.00150206, 
    0.001164514, 0.001338573, 0.001321245, 0.001085547, 0.0009549256, 
    0.0009181504, 0.0008431481, 0.0007503408, 0.0006149282,
  0.002360238, 0.001982094, 0.001588808, 0.001271087, 0.001328758, 
    0.001743409, 0.001572792, 0.001162534, 0.0009261962, 0.001155164, 
    0.001207597, 0.001045168, 0.0009525534, 0.0008577945, 0.0006955179,
  0.002257422, 0.001884489, 0.0013773, 0.001096306, 0.001197373, 0.001302951, 
    0.001443614, 0.001361617, 0.001040083, 0.000919417, 0.001030425, 
    0.001110933, 0.001003543, 0.0009166485, 0.0007584455,
  0.002107692, 0.00179764, 0.001327329, 0.001035088, 0.0009496295, 
    0.00100475, 0.001079648, 0.001062638, 0.0008388747, 0.0007567674, 
    0.0009059209, 0.0009928219, 0.0009949782, 0.0009189517, 0.0008316161,
  0.00205895, 0.001690806, 0.001252141, 0.001083073, 0.00101323, 
    0.0009905124, 0.0009115019, 0.0007814025, 0.0005954111, 0.0005841488, 
    0.0006417083, 0.000780144, 0.0009804411, 0.0009222892, 0.0008476617,
  0.001925496, 0.001561921, 0.001248531, 0.001094768, 0.001076856, 
    0.0009720977, 0.0008009498, 0.000630435, 0.0004906472, 0.0004369125, 
    0.0005006593, 0.0005011008, 0.0007617266, 0.0009096746, 0.0008466841,
  0.00141365, 0.001240138, 0.001056993, 0.0008851796, 0.0007644636, 
    0.0005669782, 0.000440639, 0.0003769642, 0.0003227428, 0.0003183137, 
    0.0003547644, 0.0003599271, 0.000550886, 0.000844863, 0.0008592446,
  0.001826258, 0.001908918, 0.001801293, 0.001656003, 0.001351493, 
    0.001118346, 0.001133909, 0.0009926257, 0.001005993, 0.0007707268, 
    0.0007834131, 0.0007594606, 0.0005511739, 0.0004351646, 0.000330007,
  0.001831241, 0.001899765, 0.001835895, 0.0016522, 0.001323154, 0.001271521, 
    0.001218525, 0.001086951, 0.001018705, 0.0009946499, 0.000893696, 
    0.0008952506, 0.0007479794, 0.0004916351, 0.0003735546,
  0.001959231, 0.001951278, 0.001868728, 0.001707142, 0.001342921, 
    0.001090411, 0.001257786, 0.001206289, 0.001077756, 0.0009362994, 
    0.001065933, 0.001020845, 0.0008768063, 0.0006939523, 0.0005042367,
  0.002095855, 0.002053602, 0.001948363, 0.001851084, 0.001512274, 
    0.001158463, 0.0009941767, 0.001235649, 0.001234307, 0.001039193, 
    0.001008579, 0.0009948205, 0.000952181, 0.0008437853, 0.0006535426,
  0.00221815, 0.002055366, 0.001895056, 0.001797731, 0.001692708, 
    0.001500816, 0.001266031, 0.00104029, 0.001025851, 0.001119205, 
    0.00115601, 0.001026615, 0.0009408502, 0.0009249815, 0.0008114635,
  0.002214983, 0.001989402, 0.001826739, 0.001625427, 0.001446402, 
    0.00145774, 0.001582167, 0.001422358, 0.001080628, 0.001026541, 
    0.001020906, 0.001094446, 0.0009931289, 0.000890463, 0.0008166145,
  0.002127401, 0.001930876, 0.001717948, 0.001486867, 0.00134603, 
    0.001245398, 0.001351469, 0.001521529, 0.00133741, 0.001065181, 
    0.000839002, 0.0007307331, 0.0007865172, 0.000787377, 0.00077521,
  0.002140985, 0.001913104, 0.001673541, 0.001426211, 0.001292589, 
    0.001238636, 0.001274567, 0.001351313, 0.001227911, 0.0009232637, 
    0.0006937421, 0.000593739, 0.000509167, 0.0004786184, 0.0005389614,
  0.001889191, 0.001632558, 0.00135387, 0.001097598, 0.0009838481, 
    0.0009865612, 0.001214505, 0.001329983, 0.001135379, 0.0008360263, 
    0.0006330571, 0.0004894103, 0.0004011955, 0.0003563526, 0.0003892047,
  0.001378313, 0.001195898, 0.0009695489, 0.0006921684, 0.0005644907, 
    0.0005150688, 0.0006496388, 0.000821265, 0.0007343219, 0.0005881364, 
    0.0004411548, 0.0003468173, 0.0003225182, 0.0003300517, 0.0003895741,
  0.001292302, 0.001674844, 0.001760545, 0.001864769, 0.001851336, 
    0.001771941, 0.001709454, 0.001415967, 0.001171751, 0.0008575801, 
    0.0007151788, 0.0005971566, 0.0004186329, 0.0003904151, 0.0004069933,
  0.001495096, 0.00164677, 0.001740364, 0.001748915, 0.001642878, 
    0.001861636, 0.001857576, 0.001505168, 0.00121476, 0.0009464971, 
    0.0008044792, 0.0007752152, 0.0006304414, 0.0003608857, 0.0003829453,
  0.001506374, 0.001656317, 0.001759402, 0.001757629, 0.001671323, 
    0.001616084, 0.001808665, 0.001565497, 0.00125305, 0.001004395, 
    0.0009918716, 0.0008743986, 0.0006534662, 0.0005727668, 0.0004452399,
  0.001586739, 0.001683358, 0.001738191, 0.001831083, 0.001791379, 
    0.001600683, 0.001474559, 0.001463711, 0.001233546, 0.0009728086, 
    0.0009344465, 0.0009057774, 0.0007408706, 0.0006242748, 0.0005510382,
  0.001820665, 0.001793177, 0.001731958, 0.001686045, 0.001676727, 
    0.001639361, 0.001436773, 0.001014333, 0.0009021251, 0.0009252696, 
    0.0009088656, 0.0008924567, 0.0008347257, 0.0007513419, 0.0005824679,
  0.001868581, 0.001748483, 0.001644042, 0.001577846, 0.001538776, 
    0.001481712, 0.001503974, 0.001298713, 0.001031422, 0.0009400339, 
    0.0008850959, 0.0009160078, 0.0009309995, 0.0009047482, 0.0006672354,
  0.001826811, 0.001756098, 0.001660988, 0.001556777, 0.001482955, 
    0.001392601, 0.001290938, 0.001259773, 0.001290046, 0.001128579, 
    0.0009504523, 0.0008907028, 0.0009150573, 0.0009512226, 0.0008482409,
  0.001555766, 0.001455278, 0.001342344, 0.001222341, 0.001140481, 
    0.001073289, 0.0009678273, 0.0009189001, 0.0009963405, 0.001096747, 
    0.001072254, 0.0009330246, 0.0009029701, 0.0009092559, 0.0008916768,
  0.001230985, 0.001137925, 0.001050741, 0.0009538901, 0.0007975296, 
    0.000678191, 0.0006628201, 0.0006356242, 0.0006328046, 0.0007910933, 
    0.001128029, 0.001018218, 0.0008941265, 0.0008379885, 0.000791706,
  0.001015483, 0.0009309087, 0.0008533891, 0.0006196437, 0.0004752462, 
    0.0004227841, 0.0004245772, 0.0004585165, 0.0004925792, 0.0006832032, 
    0.0009711073, 0.0009782707, 0.0008450185, 0.0007891406, 0.0007794151,
  0.001150681, 0.001341942, 0.001240159, 0.001419108, 0.0014117, 0.001440032, 
    0.001415104, 0.00127047, 0.001008799, 0.0009408019, 0.0009089399, 
    0.0009184623, 0.0008894747, 0.0008656664, 0.0008116303,
  0.001499546, 0.001438049, 0.001419224, 0.001366088, 0.001332549, 
    0.001449706, 0.001522888, 0.001430257, 0.001171878, 0.001087105, 
    0.001055166, 0.001084587, 0.001007182, 0.0007892211, 0.0007543621,
  0.001695996, 0.001653507, 0.001591359, 0.001484925, 0.001290843, 
    0.001196956, 0.001530209, 0.001583139, 0.001454949, 0.001222012, 
    0.001247386, 0.001170377, 0.001028615, 0.0008971345, 0.0007342766,
  0.001668001, 0.001591536, 0.001675123, 0.001729849, 0.001624509, 
    0.001439832, 0.001301631, 0.001623763, 0.001590664, 0.001333484, 
    0.001264901, 0.001209983, 0.001036713, 0.0009083073, 0.0007545594,
  0.001611639, 0.001622773, 0.001646683, 0.001625759, 0.001762557, 
    0.001669168, 0.001596174, 0.001379015, 0.001307685, 0.001283005, 
    0.001295012, 0.001171659, 0.0009765766, 0.0008525467, 0.0007074815,
  0.001399476, 0.001421683, 0.001565447, 0.001646494, 0.001655513, 
    0.001664536, 0.001723068, 0.001685989, 0.001440208, 0.001388846, 
    0.001328265, 0.001200182, 0.0009653148, 0.000782607, 0.0006378187,
  0.001200629, 0.001197516, 0.001255539, 0.001378756, 0.001520584, 0.0015982, 
    0.001594886, 0.001611922, 0.001631897, 0.001480967, 0.001365649, 
    0.001142305, 0.0009006484, 0.0007061965, 0.0005402166,
  0.001033226, 0.0009861306, 0.0009910939, 0.00102877, 0.001051722, 
    0.001147547, 0.001155248, 0.001315465, 0.001344574, 0.001410181, 
    0.001280237, 0.001079084, 0.0008412617, 0.0006467658, 0.0005107562,
  0.0009988053, 0.0009430912, 0.0009157675, 0.0008742134, 0.0007801328, 
    0.0006949915, 0.0006758279, 0.0007053092, 0.0009440535, 0.001156201, 
    0.001190425, 0.001000415, 0.0007296153, 0.0005845652, 0.0004911806,
  0.001060416, 0.0009115685, 0.0007951865, 0.0006109793, 0.0004547451, 
    0.0004073704, 0.0004225858, 0.0004906275, 0.0005496104, 0.0007348044, 
    0.0009404558, 0.0008246137, 0.0006738613, 0.0005778368, 0.0005490076,
  0.001119773, 0.00128926, 0.001030732, 0.001262456, 0.001286535, 
    0.001131106, 0.001039471, 0.0009123924, 0.000877483, 0.0008126728, 
    0.0008937704, 0.001019348, 0.001029456, 0.00101287, 0.0009098376,
  0.001400711, 0.001303919, 0.001099588, 0.001206899, 0.00119159, 
    0.001155154, 0.001066447, 0.0009368692, 0.0008875334, 0.000936691, 
    0.0009815148, 0.0011007, 0.001118415, 0.0008747082, 0.0008054513,
  0.001574736, 0.001702324, 0.001398978, 0.001131198, 0.001115057, 
    0.0008297915, 0.001105841, 0.001016027, 0.0009898745, 0.001010576, 
    0.001094818, 0.001085572, 0.001012951, 0.0009580094, 0.0008269169,
  0.001435889, 0.001594324, 0.001677983, 0.001404153, 0.001230065, 
    0.001073101, 0.0009301979, 0.001075642, 0.001075601, 0.001067232, 
    0.001087592, 0.001060006, 0.0009408618, 0.0008917514, 0.0008690783,
  0.001242705, 0.001452039, 0.001626634, 0.001620628, 0.001431133, 
    0.001342693, 0.001136413, 0.0007777347, 0.0008333444, 0.001024515, 
    0.001086193, 0.001033342, 0.0009361758, 0.0009050407, 0.0008856294,
  0.001108668, 0.001192032, 0.001573083, 0.001618918, 0.001556608, 
    0.001523654, 0.001402457, 0.001218118, 0.001081964, 0.001093328, 
    0.001131675, 0.001069601, 0.000966835, 0.000882122, 0.0008418383,
  0.001019022, 0.001037708, 0.0012392, 0.001538923, 0.001567035, 0.001522479, 
    0.001487682, 0.001467257, 0.001292082, 0.001241763, 0.001187002, 
    0.001065181, 0.0009442242, 0.000880995, 0.0008755149,
  0.001007357, 0.0009726716, 0.0010228, 0.001189188, 0.001390634, 
    0.001456569, 0.001467454, 0.001509698, 0.001375524, 0.001226951, 
    0.001096468, 0.001076898, 0.0009834528, 0.0008982152, 0.0008868988,
  0.001030023, 0.0009459839, 0.0009376146, 0.0009452218, 0.0008595409, 
    0.0009716028, 0.001090004, 0.001211915, 0.001319275, 0.00122786, 
    0.001095039, 0.001102741, 0.001015364, 0.0009195401, 0.0008030375,
  0.000986967, 0.0008421813, 0.0007705322, 0.000612502, 0.0004821771, 
    0.0004673317, 0.0006431363, 0.0009510267, 0.001015336, 0.00103561, 
    0.001118207, 0.00114023, 0.001039776, 0.0009410867, 0.0007534442,
  0.001390358, 0.001501217, 0.001360177, 0.001506426, 0.001402244, 
    0.001268526, 0.001167357, 0.001135221, 0.001144363, 0.0008614194, 
    0.0008554411, 0.0009237347, 0.0007736135, 0.0007445771, 0.0006839352,
  0.00153096, 0.001608503, 0.001523456, 0.001525211, 0.001343394, 
    0.001114401, 0.001039788, 0.001096658, 0.001040366, 0.0009873824, 
    0.0009089131, 0.001029598, 0.001045702, 0.0006964196, 0.0006415643,
  0.00143486, 0.001581999, 0.001617108, 0.001519794, 0.001174232, 
    0.0007870342, 0.0009702298, 0.0009846864, 0.0009632005, 0.0009741849, 
    0.001019013, 0.001018731, 0.00103605, 0.0009902403, 0.0007427314,
  0.001385329, 0.00161932, 0.001600858, 0.00145138, 0.00119254, 0.0009016466, 
    0.000649146, 0.0008575417, 0.0009165077, 0.0009507945, 0.0009826575, 
    0.001002816, 0.0009911139, 0.0009734341, 0.0008818741,
  0.001348334, 0.001595224, 0.001614161, 0.001502928, 0.001326791, 
    0.001036794, 0.0009078312, 0.0006249087, 0.0006813305, 0.0008497216, 
    0.0009429863, 0.001001495, 0.0009790096, 0.0009767106, 0.000912035,
  0.001345119, 0.001570269, 0.001637695, 0.001569414, 0.001460156, 
    0.001303009, 0.001099016, 0.001000907, 0.0009805887, 0.001065807, 
    0.001093274, 0.001053602, 0.0009727369, 0.0008596587, 0.0007715569,
  0.001313738, 0.001499627, 0.001660436, 0.001638668, 0.001528327, 
    0.001462122, 0.001319026, 0.001203848, 0.001134988, 0.001169805, 
    0.00115477, 0.001039399, 0.0009007553, 0.0007504934, 0.0005929264,
  0.001299482, 0.001425258, 0.001570457, 0.001626245, 0.001605097, 
    0.001523312, 0.001401877, 0.001310519, 0.001206591, 0.001168063, 
    0.001036574, 0.0009278462, 0.0007435338, 0.000558676, 0.0004619062,
  0.001256595, 0.001359156, 0.001447721, 0.001400771, 0.001307296, 
    0.00134775, 0.001290299, 0.001230645, 0.001156735, 0.001012138, 
    0.0008621163, 0.0007444351, 0.0005938276, 0.0005261329, 0.0004999809,
  0.001119404, 0.001143706, 0.001122587, 0.0008847295, 0.0008840785, 
    0.001050537, 0.001113143, 0.001064424, 0.0008956454, 0.0008246301, 
    0.0007268554, 0.0006527665, 0.0005986193, 0.0005511029, 0.0005639835,
  0.001537543, 0.001781634, 0.001712083, 0.001485812, 0.001380445, 
    0.001505521, 0.001270214, 0.001034894, 0.000922363, 0.0007998899, 
    0.0008822234, 0.0008983836, 0.0008228428, 0.0007125082, 0.0006141741,
  0.001755777, 0.0016646, 0.001365983, 0.00102194, 0.0009412126, 0.00134763, 
    0.001316636, 0.001069582, 0.0009438088, 0.0008903826, 0.0008855583, 
    0.0009559113, 0.0009431236, 0.000622668, 0.0005298762,
  0.001606998, 0.001516556, 0.001259597, 0.0009446089, 0.0009351025, 
    0.001035538, 0.001247774, 0.001058327, 0.0009822886, 0.0009340504, 
    0.0009317723, 0.0009346124, 0.0008980136, 0.0007940062, 0.0005961107,
  0.001614352, 0.001496084, 0.001342597, 0.001179588, 0.001088682, 
    0.00112906, 0.0008962839, 0.0009748939, 0.0009580398, 0.0009144518, 
    0.0009011399, 0.000871475, 0.0008256586, 0.0008815777, 0.0007721047,
  0.001655116, 0.001531504, 0.001423516, 0.001307878, 0.001208792, 
    0.001106133, 0.001057327, 0.0006940116, 0.0007096997, 0.0007165204, 
    0.000808617, 0.0008057086, 0.0007784809, 0.0008635067, 0.0008621356,
  0.001689485, 0.001577926, 0.001469902, 0.001378843, 0.001342507, 
    0.001275105, 0.00108802, 0.0009859108, 0.0009370252, 0.0009286536, 
    0.0008012537, 0.000785849, 0.000773399, 0.0008149383, 0.0008128066,
  0.001708281, 0.001631232, 0.001525066, 0.001422549, 0.001367313, 
    0.001317637, 0.001252927, 0.001122727, 0.001047528, 0.00103461, 
    0.0009299916, 0.0007679053, 0.000758754, 0.0007558947, 0.0007222137,
  0.001777689, 0.001691832, 0.001573371, 0.001475324, 0.001418723, 
    0.001338933, 0.001277991, 0.001189306, 0.001024618, 0.0008902259, 
    0.000798544, 0.0007448134, 0.0006921132, 0.0006414647, 0.000548194,
  0.001776966, 0.001688705, 0.001588099, 0.001452916, 0.001319234, 
    0.001259846, 0.001198359, 0.001089327, 0.0008890619, 0.0006962285, 
    0.0006380381, 0.0007008233, 0.000600689, 0.0005166248, 0.0004567807,
  0.001476107, 0.001389846, 0.001333849, 0.001143689, 0.00109328, 
    0.001037735, 0.0009991238, 0.0009235775, 0.0007016764, 0.0005786828, 
    0.0005304811, 0.0005711301, 0.0004982231, 0.0004502238, 0.0004489468,
  0.001248508, 0.001219567, 0.001018534, 0.001063043, 0.0009009029, 
    0.0008609207, 0.0009629054, 0.0009775952, 0.000890159, 0.0005626698, 
    0.0005986087, 0.0009018746, 0.0008886118, 0.000869943, 0.001181401,
  0.001276013, 0.001156347, 0.001102016, 0.00103509, 0.0009484941, 
    0.001047879, 0.001070993, 0.0009831832, 0.0007605267, 0.0008688467, 
    0.0008284794, 0.001057971, 0.001026643, 0.0008056707, 0.0008668484,
  0.00144209, 0.001287118, 0.001178664, 0.001148325, 0.001101614, 
    0.0008984886, 0.000923562, 0.0008384815, 0.0008186367, 0.0008825391, 
    0.0009155108, 0.0009571592, 0.001012868, 0.0009609894, 0.0008584068,
  0.001504205, 0.001490825, 0.001438543, 0.001277312, 0.001044591, 
    0.0009328554, 0.0006600128, 0.000641721, 0.0007434404, 0.0008000587, 
    0.0008356635, 0.0008847598, 0.0009559576, 0.0009710098, 0.0009067976,
  0.001416616, 0.001413205, 0.001397824, 0.001341615, 0.001123613, 
    0.0009974929, 0.0009350016, 0.0004632602, 0.0005804804, 0.000729915, 
    0.0007897485, 0.0008372758, 0.0008989378, 0.0009967422, 0.0009386044,
  0.001412176, 0.001350625, 0.001327268, 0.001291696, 0.001238101, 0.0010943, 
    0.0009198358, 0.0008785078, 0.0007590157, 0.0007609452, 0.0007656016, 
    0.0008043321, 0.0009064105, 0.0009068316, 0.0008448118,
  0.001429282, 0.001338733, 0.001255423, 0.001221641, 0.001181421, 
    0.00113667, 0.001090998, 0.0008761383, 0.000806116, 0.0008023941, 
    0.0007466408, 0.0007374029, 0.0007877438, 0.0007925822, 0.0007420597,
  0.001444662, 0.001373963, 0.001288622, 0.001233073, 0.001194222, 
    0.001166324, 0.001109412, 0.0009326158, 0.00074176, 0.0007048444, 
    0.0006513527, 0.0006607374, 0.000645643, 0.0006259012, 0.000553315,
  0.001551493, 0.001456493, 0.001381139, 0.001231877, 0.00110937, 
    0.001038847, 0.0009803852, 0.0008420358, 0.0007138521, 0.0005641287, 
    0.0005079288, 0.0005359222, 0.0005119178, 0.000514988, 0.0005453617,
  0.001470941, 0.001356772, 0.001259541, 0.000975835, 0.0008783055, 
    0.000809159, 0.0007700078, 0.0007634776, 0.0006384858, 0.0004771789, 
    0.0004815481, 0.0005396588, 0.0005536377, 0.0005171645, 0.0005813757,
  0.0009020907, 0.0009367033, 0.0007864323, 0.0007844973, 0.0006257721, 
    0.0006359988, 0.0007526646, 0.0007982185, 0.0008329937, 0.0007845858, 
    0.0008583507, 0.001159275, 0.001146059, 0.00106756, 0.0009847258,
  0.00109148, 0.0009597733, 0.0008664211, 0.0007580524, 0.0006444335, 
    0.0006415929, 0.0007760911, 0.0007434114, 0.0007335758, 0.0008258015, 
    0.0008170918, 0.001074609, 0.001172077, 0.0009512314, 0.0008620259,
  0.001340134, 0.001089289, 0.0009617395, 0.0009064375, 0.0008163765, 
    0.0005018722, 0.0006779765, 0.0007119311, 0.0007446186, 0.0007236237, 
    0.0007885942, 0.0009177874, 0.001059646, 0.00109889, 0.0009738854,
  0.00129569, 0.001317026, 0.001237516, 0.001036373, 0.0008842243, 
    0.0008061365, 0.0004367381, 0.0004653325, 0.0005744679, 0.0006223764, 
    0.0006268548, 0.0008216393, 0.0008825937, 0.001001969, 0.0009947278,
  0.001213163, 0.001167675, 0.001162717, 0.001112162, 0.0009054122, 
    0.0008411473, 0.0008291461, 0.00049883, 0.0005684985, 0.0005813292, 
    0.000589602, 0.0006780695, 0.0007446253, 0.0009460734, 0.001022927,
  0.001216124, 0.001149347, 0.001080457, 0.001058564, 0.001011955, 
    0.000916763, 0.0007905338, 0.0007755546, 0.0007527891, 0.000700965, 
    0.0005732503, 0.0007366954, 0.0007586654, 0.0008949809, 0.0009322634,
  0.001322972, 0.001211502, 0.001095704, 0.001048618, 0.0009985243, 
    0.0009940432, 0.0009231191, 0.0007608363, 0.0007237767, 0.0006627347, 
    0.0005685399, 0.0007130982, 0.0008224678, 0.0009211147, 0.0008739953,
  0.001396201, 0.001290898, 0.001179021, 0.001156181, 0.001077399, 
    0.0009749516, 0.0009191326, 0.000785764, 0.0005980327, 0.0005093881, 
    0.0004861858, 0.0006567746, 0.0008561123, 0.000889616, 0.0007377327,
  0.001565599, 0.001426304, 0.001222224, 0.001077731, 0.001023428, 
    0.0009181585, 0.0008217912, 0.0006855927, 0.0005345994, 0.0004657251, 
    0.0004266863, 0.0004812531, 0.0006968397, 0.0007659394, 0.0006879277,
  0.001462692, 0.001322732, 0.001260882, 0.0008872684, 0.0008260815, 
    0.000692594, 0.0006969623, 0.0006902147, 0.0004732784, 0.0004029291, 
    0.0003456725, 0.0004263966, 0.0004722591, 0.0006204438, 0.0006346827,
  0.0007959139, 0.0008278707, 0.0007499365, 0.0008087077, 0.0007697158, 
    0.0007045017, 0.0007251283, 0.000719674, 0.0007588518, 0.0008469204, 
    0.0009707537, 0.001006758, 0.0007920092, 0.0007294178, 0.0008298266,
  0.001019865, 0.0009008486, 0.000867166, 0.0008536577, 0.0008304002, 
    0.0006156023, 0.0007322711, 0.0006980602, 0.0007650138, 0.0008728279, 
    0.00105334, 0.001124637, 0.0009396084, 0.000678622, 0.000672542,
  0.001108987, 0.001020433, 0.0009670351, 0.0009344861, 0.0008749817, 
    0.0005959937, 0.0007353437, 0.0006735315, 0.0007271938, 0.0008895612, 
    0.00110218, 0.001166774, 0.0009660999, 0.0008522857, 0.0007606078,
  0.001156829, 0.001033769, 0.0009930191, 0.0009436014, 0.0009389207, 
    0.0009092838, 0.0006815242, 0.0005678691, 0.0006552087, 0.0008530015, 
    0.001020845, 0.001088827, 0.0009468314, 0.0008677288, 0.0008657616,
  0.001294718, 0.001139726, 0.001068497, 0.0009931142, 0.0009351152, 
    0.0009662934, 0.0008807979, 0.0005339693, 0.0005495992, 0.0007475789, 
    0.0008886897, 0.0009350759, 0.0009002652, 0.0008902009, 0.0009098123,
  0.001664636, 0.001521832, 0.001350242, 0.001151961, 0.001043172, 
    0.001023424, 0.0008728153, 0.0007534691, 0.0006560004, 0.0007309137, 
    0.0007879969, 0.0008476507, 0.0008297626, 0.0008299477, 0.0008649663,
  0.00196688, 0.001875558, 0.001750451, 0.001579372, 0.001333742, 
    0.001054357, 0.001026757, 0.0008147209, 0.0006909305, 0.0006675959, 
    0.0007507769, 0.0007929906, 0.0007659638, 0.0007652989, 0.0007820574,
  0.002033851, 0.001903482, 0.00180613, 0.001597762, 0.00146523, 0.001169314, 
    0.001019777, 0.0008430178, 0.0005880365, 0.0005881807, 0.0006179316, 
    0.0007356987, 0.0007373016, 0.0007039838, 0.0006787834,
  0.002176214, 0.001990064, 0.001797579, 0.001517567, 0.001388821, 
    0.001248256, 0.000981768, 0.0006948082, 0.0005318859, 0.0005070095, 
    0.0004886934, 0.0005432263, 0.0006858638, 0.0006642923, 0.0007055941,
  0.002452204, 0.00215318, 0.001909796, 0.001540056, 0.00119771, 0.001021066, 
    0.0008995443, 0.00074064, 0.0004908129, 0.0004451608, 0.0003590433, 
    0.0004321272, 0.0004754027, 0.0005832507, 0.0006880375,
  0.0007588147, 0.0008599744, 0.0009153812, 0.0009825152, 0.0009743248, 
    0.0009341948, 0.0009665536, 0.0009263335, 0.0008902802, 0.0007467238, 
    0.0006180495, 0.0005993113, 0.0006273686, 0.0007752799, 0.0008247537,
  0.001170023, 0.001038611, 0.001030799, 0.001027169, 0.00102939, 
    0.000887874, 0.001020923, 0.0009510684, 0.0008668701, 0.0008306029, 
    0.0007226936, 0.0007580962, 0.0008195339, 0.0007403792, 0.0007499843,
  0.001599644, 0.00144435, 0.001420125, 0.001312734, 0.001314663, 
    0.001056704, 0.001152501, 0.0009158971, 0.0008385842, 0.0008452622, 
    0.0008039051, 0.0007802176, 0.0008150977, 0.0009494136, 0.0008775015,
  0.001605705, 0.001514139, 0.001452599, 0.001495652, 0.001630029, 
    0.001534781, 0.0007992656, 0.0007691326, 0.0008008351, 0.0008991141, 
    0.0008718648, 0.0008259561, 0.0007970626, 0.0009156633, 0.0009302878,
  0.001620389, 0.001496979, 0.001543731, 0.001669464, 0.001611421, 
    0.001165749, 0.0008206983, 0.0005320663, 0.000567553, 0.0008700428, 
    0.0008676708, 0.0007851627, 0.0007907608, 0.0009279551, 0.0009589278,
  0.001721564, 0.001602951, 0.001730446, 0.001757091, 0.001518904, 
    0.001055573, 0.0008334413, 0.0007648517, 0.0007979857, 0.0009213449, 
    0.0008018901, 0.0007448637, 0.0007786644, 0.0009485499, 0.0009361622,
  0.001856573, 0.001722543, 0.001802282, 0.001718343, 0.001468105, 
    0.001143911, 0.001009479, 0.0008754724, 0.0008864444, 0.0008598427, 
    0.0007790743, 0.0007230468, 0.0007791852, 0.0008982635, 0.0008860402,
  0.001927777, 0.001804153, 0.001836304, 0.001640692, 0.001406946, 
    0.001191608, 0.001056149, 0.0008846395, 0.0008137409, 0.0007560281, 
    0.0006822525, 0.0006692402, 0.0008116559, 0.0008379252, 0.0007384133,
  0.002011182, 0.001963532, 0.001854514, 0.001500266, 0.001122338, 
    0.0009425132, 0.0008255097, 0.0007279345, 0.0007024345, 0.0006578375, 
    0.000632196, 0.0006742512, 0.0007358841, 0.0007321155, 0.0006290278,
  0.002094554, 0.001970285, 0.001629522, 0.001011808, 0.0008029936, 
    0.0006903734, 0.0006445073, 0.0006284373, 0.0005459277, 0.0004922534, 
    0.0004782732, 0.000578059, 0.0006080359, 0.0005631063, 0.0005513872,
  0.0009770471, 0.0009416079, 0.0008803158, 0.0008095417, 0.000739452, 
    0.0007092837, 0.0007609021, 0.000721974, 0.0007295062, 0.0006894237, 
    0.0006736764, 0.0007354516, 0.0007318081, 0.0007144432, 0.0005979612,
  0.001136523, 0.00101087, 0.0009412069, 0.0008759109, 0.0007772172, 
    0.0007860491, 0.0008659492, 0.0008541182, 0.0008565372, 0.0009195675, 
    0.0008583619, 0.0008947222, 0.0009647377, 0.0006853217, 0.0005105183,
  0.00118615, 0.001045692, 0.0009819301, 0.0009352486, 0.000884773, 
    0.0007318124, 0.0009078397, 0.0009769684, 0.000992212, 0.001070524, 
    0.0009901325, 0.0008903714, 0.0009599624, 0.0009724534, 0.0006924202,
  0.001385666, 0.001342375, 0.001370026, 0.001324651, 0.001169282, 
    0.00113187, 0.0008429622, 0.0009306949, 0.001017711, 0.0009232527, 
    0.000813438, 0.0007213739, 0.0008798402, 0.0008302261, 0.0007167552,
  0.001475243, 0.001537002, 0.00149413, 0.001506527, 0.001168921, 
    0.001035124, 0.001163141, 0.0006825135, 0.0006036005, 0.0005564322, 
    0.0005758435, 0.0007593962, 0.0008461857, 0.0007757562, 0.0007063359,
  0.001467673, 0.001398994, 0.001333002, 0.001335834, 0.001240121, 
    0.001065572, 0.001089792, 0.0009486999, 0.0007982657, 0.0007901291, 
    0.0006633208, 0.0008233491, 0.0008097116, 0.0007510225, 0.0006585752,
  0.001473303, 0.001383792, 0.00132886, 0.001245368, 0.001186118, 
    0.001155298, 0.001090661, 0.000899142, 0.0008577092, 0.0008090224, 
    0.0007438433, 0.0006966428, 0.0006425941, 0.0005498342, 0.0005320327,
  0.001507652, 0.001442932, 0.001344395, 0.001267771, 0.001236169, 
    0.001204753, 0.001155397, 0.0009043369, 0.0007821356, 0.0006885321, 
    0.0006566272, 0.0006163934, 0.0005521618, 0.0004797131, 0.0004415567,
  0.001559165, 0.001501144, 0.001412512, 0.00125007, 0.001127878, 
    0.001052068, 0.0009325749, 0.0007929422, 0.0007068668, 0.000636872, 
    0.0006294586, 0.000614602, 0.0005650042, 0.0005200089, 0.0005318986,
  0.001531289, 0.001420555, 0.001222484, 0.0008489952, 0.0008306061, 
    0.0007823551, 0.0007337054, 0.0007172926, 0.0006539724, 0.0005890488, 
    0.0005795005, 0.0005953415, 0.0005903534, 0.0005207544, 0.0005596928,
  0.001082741, 0.001017632, 0.0009538549, 0.0009537684, 0.0008034174, 
    0.0006818417, 0.0007428267, 0.0006363709, 0.0005430976, 0.0003142463, 
    0.0003337042, 0.0003908947, 0.0003298467, 0.0003509618, 0.0003466005,
  0.001202655, 0.001102809, 0.001045433, 0.0009925644, 0.0008266486, 
    0.0007759575, 0.0007854326, 0.0006679785, 0.0006047484, 0.0005253815, 
    0.0004834991, 0.0005788236, 0.0006175407, 0.0004823738, 0.0004438057,
  0.001216008, 0.001036034, 0.001030205, 0.001039163, 0.0008889139, 
    0.0006899404, 0.0007766615, 0.0006904908, 0.0006022807, 0.0006372326, 
    0.0006664629, 0.0007261792, 0.0008174467, 0.0008677837, 0.0008499991,
  0.001083204, 0.001102029, 0.001199441, 0.00114102, 0.0009237305, 
    0.0008895134, 0.0006205906, 0.0006062184, 0.0006039311, 0.0006448353, 
    0.0007716069, 0.0008264898, 0.0009062712, 0.0009435913, 0.0009452845,
  0.001217311, 0.001163461, 0.001208748, 0.001251096, 0.0009820515, 
    0.0009455259, 0.0009622163, 0.0004876812, 0.0004338718, 0.0004734774, 
    0.0005156694, 0.0006989641, 0.0007567276, 0.0007440575, 0.0007652062,
  0.001372469, 0.001285243, 0.001259756, 0.001236421, 0.00117867, 
    0.001096402, 0.001019776, 0.001017253, 0.0008550216, 0.0007577292, 
    0.0005133243, 0.0005870583, 0.0005561797, 0.0005747034, 0.0006091971,
  0.001430465, 0.001364741, 0.00130962, 0.001244702, 0.001230041, 
    0.001237276, 0.001074743, 0.0009016237, 0.0007429132, 0.0005895031, 
    0.0005095061, 0.0004888137, 0.0004641767, 0.0004436454, 0.0004900029,
  0.001485167, 0.001427555, 0.001321736, 0.001311987, 0.001305645, 
    0.001270823, 0.001139719, 0.0007706865, 0.0005877159, 0.0004792941, 
    0.0004248209, 0.0004068023, 0.000400431, 0.0003930209, 0.0004096263,
  0.001538244, 0.001476913, 0.001448564, 0.001351246, 0.001216254, 
    0.001083665, 0.0008600367, 0.0006064564, 0.0005310505, 0.0004150589, 
    0.0003634578, 0.0003655943, 0.0003752216, 0.000410642, 0.0004092008,
  0.001618857, 0.00152617, 0.001345477, 0.0009557265, 0.0008689412, 
    0.0007321787, 0.0006708898, 0.0006108917, 0.0004751649, 0.0003268232, 
    0.000276361, 0.0003574005, 0.0003873791, 0.0004015279, 0.000415713,
  0.001108572, 0.001206161, 0.001151764, 0.001157695, 0.0009627831, 
    0.0008086499, 0.0008404998, 0.0006808156, 0.0005009954, 0.0003054441, 
    0.0003081355, 0.0003638522, 0.0002774343, 0.0002964442, 0.0002500317,
  0.001297451, 0.001216393, 0.001129071, 0.001103696, 0.0008106588, 
    0.0007984095, 0.0008067867, 0.0006142588, 0.0004882666, 0.0004169063, 
    0.0003683562, 0.0004880503, 0.0005215287, 0.0003720983, 0.0003482983,
  0.001613224, 0.001217965, 0.001026756, 0.0009905687, 0.0008506567, 
    0.0006382747, 0.0006728002, 0.0005373836, 0.0004592803, 0.0005136082, 
    0.0005481804, 0.0005794271, 0.0006374783, 0.000700767, 0.0006847883,
  0.001431559, 0.001287804, 0.001203846, 0.001102875, 0.0009409455, 
    0.0008602662, 0.0004501653, 0.0004555745, 0.0004254622, 0.0004744226, 
    0.000572951, 0.0006224292, 0.0006997235, 0.0007443849, 0.000736053,
  0.001365144, 0.001304393, 0.001286544, 0.001333799, 0.0009981568, 
    0.0009641431, 0.0009071147, 0.000413028, 0.0003268056, 0.0004445652, 
    0.0004723718, 0.000568315, 0.0006556978, 0.0006492913, 0.0006090511,
  0.001405829, 0.00137713, 0.001343892, 0.001337221, 0.001248411, 
    0.001100484, 0.0009327309, 0.0009318975, 0.0007495832, 0.000670723, 
    0.0003862058, 0.0005370085, 0.0005335225, 0.0005069676, 0.0005487896,
  0.00146952, 0.001431105, 0.001392801, 0.001332032, 0.001327052, 
    0.001267995, 0.001073542, 0.0009684042, 0.0006927985, 0.0005534294, 
    0.0004600151, 0.0004290574, 0.0004322092, 0.0004279163, 0.0004862879,
  0.001475846, 0.001400495, 0.001321806, 0.001278269, 0.001253751, 
    0.001235431, 0.001154643, 0.0008657611, 0.000561304, 0.0004563914, 
    0.0003993834, 0.0003911187, 0.0004075095, 0.0004322006, 0.0004858337,
  0.001494146, 0.00140213, 0.001327673, 0.001260075, 0.001178488, 
    0.001118155, 0.0009783359, 0.0006411453, 0.0004826605, 0.0003936906, 
    0.0003588674, 0.0003631783, 0.0003953537, 0.0004523667, 0.0004620464,
  0.001583705, 0.001524605, 0.001449187, 0.001179557, 0.00100865, 
    0.000818508, 0.0007614465, 0.000615009, 0.0004282775, 0.0002851952, 
    0.0002356774, 0.0003297899, 0.0003728092, 0.0003935049, 0.0004010651,
  0.0009781726, 0.0009871953, 0.0009741007, 0.0009885472, 0.0009328161, 
    0.0007728367, 0.0009857015, 0.0008271234, 0.0006940152, 0.0005813903, 
    0.0005122109, 0.0004757582, 0.0003551274, 0.0003149803, 0.0002367092,
  0.0011337, 0.001013778, 0.001084197, 0.001071126, 0.0007018996, 
    0.0007146806, 0.0007421414, 0.0006985838, 0.0006449798, 0.0006134629, 
    0.0005107575, 0.0005144039, 0.0004538537, 0.0002643706, 0.0002744727,
  0.001574817, 0.001272418, 0.001107973, 0.001038138, 0.0007760378, 
    0.0005157415, 0.0006120368, 0.0006092804, 0.0006051542, 0.0005924946, 
    0.0005404379, 0.0004972406, 0.0005236655, 0.000535211, 0.000543373,
  0.001320522, 0.001230282, 0.001185554, 0.0009885393, 0.0008099469, 
    0.0007366975, 0.0004061735, 0.0004657768, 0.0004685052, 0.0004304144, 
    0.0005213706, 0.0005473381, 0.0006112816, 0.0006176644, 0.0006248661,
  0.001371433, 0.001281428, 0.001283129, 0.001184952, 0.0008470022, 
    0.0008374313, 0.0008009743, 0.0003667693, 0.0002913841, 0.0003327101, 
    0.0003958281, 0.0005005851, 0.0005950238, 0.000593011, 0.0006290062,
  0.001389331, 0.001346341, 0.001324628, 0.001237403, 0.001074142, 
    0.000891683, 0.0008244085, 0.0008369664, 0.0007058925, 0.000535327, 
    0.0004000901, 0.0004806364, 0.0005379428, 0.0005779134, 0.0006177929,
  0.001356518, 0.001335276, 0.001289749, 0.001227701, 0.001208313, 
    0.001154217, 0.0009425708, 0.0007866902, 0.0006129178, 0.0005375383, 
    0.0004760008, 0.0004401173, 0.0004371923, 0.0004732376, 0.0005696358,
  0.001366192, 0.0013105, 0.001249379, 0.001184404, 0.001161985, 0.001163382, 
    0.001116904, 0.000689049, 0.0005126707, 0.0004457936, 0.0003918787, 
    0.000389392, 0.0003902134, 0.000439586, 0.0004879393,
  0.001468599, 0.001372139, 0.001275579, 0.001205577, 0.001183776, 
    0.001119274, 0.0009031068, 0.0005565797, 0.0004714675, 0.0003975846, 
    0.0003735356, 0.0003882587, 0.0004198042, 0.0004462633, 0.0004313198,
  0.00161566, 0.001517367, 0.001462267, 0.00134992, 0.001041695, 
    0.0008801417, 0.0007012562, 0.0005022381, 0.0004112757, 0.0003038025, 
    0.0003022074, 0.0003789594, 0.000395592, 0.000389771, 0.0004037582,
  0.001006736, 0.0009823011, 0.0008874878, 0.0007315426, 0.0006184022, 
    0.0005356625, 0.0006942084, 0.0007402005, 0.0007676345, 0.0005720399, 
    0.0004743141, 0.0005136624, 0.0004298514, 0.0003250871, 0.0002397101,
  0.001084617, 0.0009902683, 0.000792174, 0.0006713173, 0.0005153423, 
    0.0004821184, 0.0005546432, 0.0005939304, 0.0006490304, 0.0006551039, 
    0.000511672, 0.0005348908, 0.0005101548, 0.0002350139, 0.0001595515,
  0.001346509, 0.001011347, 0.0008044319, 0.0007302599, 0.0006105584, 
    0.0003623689, 0.0004475604, 0.0004969691, 0.0005599964, 0.0006301169, 
    0.0006274083, 0.0006034864, 0.0006189318, 0.0005587117, 0.000395723,
  0.001409433, 0.001261334, 0.001114473, 0.0008423994, 0.0007391425, 
    0.0007316986, 0.0002917075, 0.0003919668, 0.0004616416, 0.0005081396, 
    0.0006030259, 0.0006131324, 0.0006191154, 0.0005881498, 0.0005118567,
  0.001428873, 0.001249513, 0.001200358, 0.001065016, 0.0008064589, 
    0.000821251, 0.000804072, 0.0003258072, 0.0003164207, 0.0004214085, 
    0.0004891125, 0.0005445878, 0.0005570347, 0.0005311203, 0.0004789382,
  0.001461449, 0.001303449, 0.001175147, 0.00109004, 0.0009566693, 
    0.000853584, 0.0007723112, 0.0007406707, 0.00052466, 0.0004963193, 
    0.000429213, 0.0004876847, 0.0005102656, 0.0005055268, 0.0004747191,
  0.001488205, 0.001360382, 0.001208093, 0.001093737, 0.001074931, 
    0.001093902, 0.0007228786, 0.0005476631, 0.0004962853, 0.0004538521, 
    0.0004214401, 0.000414136, 0.0004379236, 0.0004425447, 0.0004849657,
  0.001488189, 0.001316328, 0.001189709, 0.001154589, 0.001176598, 
    0.00114725, 0.0009248391, 0.0005429522, 0.0004543608, 0.0004062059, 
    0.0003761995, 0.0003745249, 0.000388433, 0.0004217351, 0.0004576464,
  0.00149041, 0.001349246, 0.001286127, 0.001242493, 0.001162141, 
    0.0009549573, 0.0006337868, 0.000492281, 0.000416848, 0.0003772881, 
    0.0003509984, 0.0003622883, 0.0003787088, 0.0003953232, 0.0003987014,
  0.001554734, 0.001479088, 0.001403205, 0.0009271907, 0.0006806531, 
    0.00057799, 0.0005329731, 0.0004764055, 0.000387404, 0.0003026479, 
    0.0002889397, 0.0003605629, 0.0003604764, 0.0003598072, 0.0003797565,
  0.000815442, 0.0008080525, 0.0006601411, 0.000636693, 0.0005149605, 
    0.0004168105, 0.0005043528, 0.0005206161, 0.0006009801, 0.0004032758, 
    0.0003365766, 0.0004151254, 0.0003796435, 0.0002847764, 0.0002212644,
  0.0008552846, 0.0007416122, 0.000664587, 0.0005755597, 0.0004232028, 
    0.0003113548, 0.0003888155, 0.0004232192, 0.000487779, 0.0005130972, 
    0.0003851796, 0.0004726382, 0.0004767054, 0.0002448696, 0.0001634662,
  0.001111611, 0.0008411235, 0.0007828386, 0.000714715, 0.0006317958, 
    0.0002609754, 0.0003100012, 0.0003747315, 0.0004006842, 0.0004363623, 
    0.0004620081, 0.0004645016, 0.0004491427, 0.0004111839, 0.0002606832,
  0.001243675, 0.001139069, 0.001008268, 0.0008580562, 0.0008009616, 
    0.0008128871, 0.0002245405, 0.0003228473, 0.0003934147, 0.0003885679, 
    0.0004234854, 0.0004482013, 0.0004376528, 0.0003917114, 0.0002969306,
  0.001276826, 0.00107942, 0.001048217, 0.001051699, 0.0008740925, 
    0.0008180593, 0.0008010201, 0.0002483797, 0.0002801519, 0.0003567876, 
    0.0003935566, 0.0004182245, 0.0004451402, 0.0004251336, 0.0003956697,
  0.001334028, 0.001146922, 0.001086416, 0.001056286, 0.0009366604, 
    0.0007247217, 0.0006704648, 0.0006089559, 0.0004677011, 0.0004440974, 
    0.0003781649, 0.0004056222, 0.0004416755, 0.0004432807, 0.0004351067,
  0.00142139, 0.001198665, 0.001119733, 0.001088442, 0.00108936, 
    0.0009682815, 0.0006481112, 0.0005300141, 0.0004742463, 0.000441247, 
    0.0004113343, 0.0003885933, 0.0003852471, 0.0003939106, 0.0004372668,
  0.001459663, 0.001232189, 0.001173544, 0.00114831, 0.001126496, 
    0.001050126, 0.0008333417, 0.0005256619, 0.0004536333, 0.0004058556, 
    0.0003658168, 0.0003590616, 0.0003500679, 0.0003790727, 0.0004372428,
  0.001448672, 0.001326327, 0.001302855, 0.001226004, 0.001102891, 
    0.0008888337, 0.0006121858, 0.0005023406, 0.0004277102, 0.0003614656, 
    0.0003190647, 0.0003191986, 0.0003351055, 0.0003597747, 0.0003562193,
  0.001556367, 0.001537045, 0.001357904, 0.0007817216, 0.0005891986, 
    0.00054078, 0.000529752, 0.0004976285, 0.0003941773, 0.0002695176, 
    0.0002157287, 0.0002925751, 0.0002863934, 0.0002967532, 0.0003225438,
  0.0007792658, 0.0007978053, 0.0007073295, 0.0007094082, 0.000636753, 
    0.0005756925, 0.0005650753, 0.0005490176, 0.0005503531, 0.0003770168, 
    0.0003126809, 0.0003245716, 0.0002564679, 0.0002492509, 0.0001738773,
  0.0008090225, 0.0007351886, 0.0006696404, 0.0005967765, 0.0005022148, 
    0.0003653282, 0.000454962, 0.0004856481, 0.0005110267, 0.00046742, 
    0.0003157099, 0.0003949489, 0.0004236759, 0.0002442692, 0.0001749141,
  0.001073201, 0.0007696434, 0.0006821746, 0.0006013443, 0.0005177924, 
    0.0002720373, 0.0003255642, 0.0004010783, 0.0004283263, 0.0004460037, 
    0.0004023466, 0.0003995444, 0.0004349974, 0.0004628592, 0.0003387882,
  0.001197906, 0.001149292, 0.0009933759, 0.0007340589, 0.0006279324, 
    0.0006192905, 0.0002411612, 0.0003176743, 0.0003689053, 0.0003628729, 
    0.0003843466, 0.0004166499, 0.0004505158, 0.000436639, 0.0003410149,
  0.001170214, 0.001143075, 0.001138757, 0.0009882255, 0.0008004906, 
    0.0006707669, 0.000696309, 0.0002390708, 0.0001933152, 0.0002623137, 
    0.0003519757, 0.000413559, 0.0004425879, 0.0004078885, 0.0003754014,
  0.001182909, 0.001156283, 0.001119742, 0.001041204, 0.0008563318, 
    0.0007277254, 0.0006864177, 0.0007128517, 0.0005415883, 0.0004026037, 
    0.0003115328, 0.0003784746, 0.0004505824, 0.000457018, 0.0004158358,
  0.001260074, 0.001243743, 0.001153838, 0.001070734, 0.001044183, 
    0.0009278925, 0.0006774574, 0.0005910512, 0.000476715, 0.0004087875, 
    0.0003561393, 0.0003338977, 0.0003360062, 0.0003666945, 0.0004005918,
  0.001356293, 0.001291406, 0.001218307, 0.00112661, 0.001078342, 
    0.001038931, 0.0008073382, 0.0005442577, 0.0004388015, 0.0003415903, 
    0.0002945777, 0.0002942128, 0.0002814742, 0.0003114296, 0.0003682152,
  0.001354429, 0.001332435, 0.001322847, 0.00115425, 0.001069125, 
    0.0009779597, 0.0007031334, 0.0005195667, 0.0004197154, 0.0003004325, 
    0.0002761423, 0.0002737108, 0.0002754579, 0.0003154317, 0.0003794183,
  0.001580715, 0.001527839, 0.001355515, 0.0009719137, 0.0008251839, 
    0.0007299088, 0.0006067126, 0.0005202705, 0.0003737676, 0.0002331646, 
    0.0002078555, 0.000273221, 0.0002860063, 0.0003247862, 0.0003819149,
  0.0008180825, 0.0008213343, 0.0007751962, 0.0007903856, 0.0008291377, 
    0.0008151812, 0.0008514627, 0.0008601123, 0.0008762326, 0.0007276786, 
    0.0006566011, 0.0006460142, 0.0005502373, 0.0004983796, 0.0003677678,
  0.0009366769, 0.0008485586, 0.0008162688, 0.000793685, 0.0006996822, 
    0.0005886605, 0.0006674854, 0.0006924053, 0.0007161078, 0.0006950386, 
    0.0005686797, 0.0005924291, 0.0005461558, 0.0003245826, 0.0002489909,
  0.001164395, 0.0009264625, 0.0008505213, 0.000808205, 0.0006749147, 
    0.000406754, 0.0004565342, 0.0005121627, 0.0005425741, 0.0005671016, 
    0.0005365878, 0.0005070189, 0.0005008792, 0.0004533154, 0.0003218246,
  0.001198572, 0.00119472, 0.001064908, 0.0008273622, 0.0007266935, 
    0.000631541, 0.0003330561, 0.0003784074, 0.000395071, 0.0004136067, 
    0.0004671064, 0.0004721211, 0.0004826011, 0.0004665899, 0.0003946336,
  0.001200792, 0.001163553, 0.001136943, 0.0009499963, 0.000733779, 
    0.0006506806, 0.0006730625, 0.0002666424, 0.000220073, 0.000285416, 
    0.0003601979, 0.0004320757, 0.0004626038, 0.0004566531, 0.0004713353,
  0.001251942, 0.001156304, 0.001119548, 0.0009943915, 0.0008264941, 
    0.0007298416, 0.0006671858, 0.0006951952, 0.0005121151, 0.0003590183, 
    0.0002814598, 0.0003342451, 0.0003926606, 0.0004175387, 0.0004162028,
  0.001462818, 0.001269485, 0.001137362, 0.001028404, 0.0009576251, 
    0.0008611985, 0.0006506376, 0.0005510626, 0.0003953394, 0.0003511984, 
    0.0003249434, 0.0003123973, 0.0003218288, 0.0003276466, 0.0003687723,
  0.001876618, 0.001662223, 0.001450573, 0.001295374, 0.001043134, 
    0.0008977501, 0.0007296606, 0.0005402687, 0.0004402356, 0.0003847159, 
    0.0003290576, 0.0003028122, 0.0002724215, 0.0002769205, 0.0003626503,
  0.001949548, 0.001811755, 0.001703357, 0.001527064, 0.001233842, 
    0.0009458121, 0.0007186661, 0.0005766231, 0.0005220349, 0.0004635092, 
    0.0004247548, 0.0003900007, 0.0003554054, 0.000360786, 0.0003669768,
  0.001860698, 0.001750619, 0.001734375, 0.00140869, 0.0009594513, 
    0.0007563318, 0.0006289817, 0.0006048528, 0.0005704242, 0.000492131, 
    0.0005070035, 0.0005196314, 0.0004695216, 0.0004468874, 0.000422948,
  0.001022461, 0.001055812, 0.001008657, 0.0009472386, 0.0009328287, 
    0.0009613413, 0.001277146, 0.001404269, 0.001498591, 0.001368197, 
    0.001435451, 0.001616472, 0.001395327, 0.001219752, 0.0009888337,
  0.00110504, 0.001113675, 0.001073979, 0.00106408, 0.0008817837, 
    0.0007114915, 0.0008472382, 0.001154588, 0.001338743, 0.001418217, 
    0.00128914, 0.001455789, 0.001329706, 0.0009081534, 0.0007349025,
  0.001239235, 0.001174762, 0.00109946, 0.001085667, 0.0009388826, 
    0.0006094952, 0.0006124187, 0.0006991014, 0.0009170517, 0.001129563, 
    0.001199781, 0.00121155, 0.001157614, 0.001004344, 0.0007138519,
  0.001340996, 0.001311515, 0.001238323, 0.001050586, 0.000969241, 
    0.0008893372, 0.000495255, 0.000505869, 0.000508078, 0.000659899, 
    0.0008349406, 0.0008639639, 0.0008434071, 0.0007500855, 0.0006112217,
  0.001438931, 0.001341152, 0.001333925, 0.001261031, 0.0009565796, 
    0.0009311294, 0.0008971266, 0.0003418934, 0.0003007912, 0.0004172217, 
    0.0005303318, 0.0006390263, 0.0006798876, 0.0006322861, 0.0005788276,
  0.001635883, 0.0014833, 0.001381793, 0.001331848, 0.0009982716, 
    0.0009118152, 0.0008388027, 0.0007318854, 0.0005020377, 0.0004169452, 
    0.0003578543, 0.0004500708, 0.0005413783, 0.0005662742, 0.000534322,
  0.002009894, 0.001796728, 0.001517194, 0.001418977, 0.001260445, 
    0.001173802, 0.0008831957, 0.0006882718, 0.0005175858, 0.0004247949, 
    0.0003669481, 0.0003767691, 0.0003857167, 0.0004313163, 0.0004788921,
  0.002176474, 0.002055305, 0.001847862, 0.001553003, 0.00139848, 
    0.001310176, 0.00112329, 0.0008826027, 0.0007945755, 0.0005625237, 
    0.0004105573, 0.0003504374, 0.0003051471, 0.0003191053, 0.0004446536,
  0.00207685, 0.002019979, 0.001951881, 0.001626408, 0.001410067, 
    0.001189279, 0.0009790377, 0.0008279905, 0.0007807678, 0.0007368695, 
    0.0006128406, 0.0004476574, 0.000359972, 0.0003541067, 0.0003755324,
  0.001977966, 0.001852736, 0.001539825, 0.001182421, 0.001088137, 
    0.0009953824, 0.0009157652, 0.0007543843, 0.0006202045, 0.000533309, 
    0.0006683358, 0.0006616216, 0.000493212, 0.0004190254, 0.0004032513,
  0.001286084, 0.001614162, 0.001300476, 0.00119115, 0.001125455, 
    0.0008979059, 0.001075814, 0.001410669, 0.001510187, 0.001208218, 
    0.001257478, 0.001696936, 0.001385937, 0.001433805, 0.001144207,
  0.001436912, 0.001627913, 0.001444422, 0.001276987, 0.001117425, 
    0.0007853275, 0.0007973178, 0.001104362, 0.001594331, 0.001658259, 
    0.001425001, 0.00183953, 0.001721996, 0.001353106, 0.001095958,
  0.001789608, 0.001824406, 0.001632646, 0.001323527, 0.001188561, 
    0.0007457069, 0.0006830815, 0.0007222001, 0.0008871002, 0.001260499, 
    0.001613675, 0.001698183, 0.001726988, 0.001609374, 0.001218934,
  0.001780994, 0.001895779, 0.00203895, 0.00147329, 0.001272692, 0.001211383, 
    0.0005274396, 0.0005904481, 0.0006052454, 0.0006579369, 0.0009841735, 
    0.001285238, 0.001435885, 0.001409409, 0.001257179,
  0.001896313, 0.002024675, 0.002011105, 0.001940933, 0.001361128, 
    0.001324634, 0.001081175, 0.0003504598, 0.0003711884, 0.0004753399, 
    0.0005453885, 0.0008332562, 0.001000856, 0.001145516, 0.001189137,
  0.002045468, 0.002070188, 0.001978762, 0.001857229, 0.001647211, 
    0.001427625, 0.001109903, 0.0008346786, 0.0005664157, 0.0004654386, 
    0.0003862766, 0.0004899714, 0.0006719359, 0.0008301081, 0.0009206258,
  0.002051182, 0.002023276, 0.001942984, 0.001740955, 0.001499936, 
    0.001483921, 0.001127254, 0.0008872725, 0.0007053936, 0.0005298725, 
    0.0004319856, 0.0003685596, 0.0004056394, 0.0005284895, 0.0006829827,
  0.001903577, 0.002036653, 0.001995364, 0.001567888, 0.001498111, 
    0.001394181, 0.001038688, 0.0007584877, 0.0007179833, 0.00063156, 
    0.0005291625, 0.0003450981, 0.0003067057, 0.0003530065, 0.0004634905,
  0.0018204, 0.001920704, 0.001912998, 0.00167236, 0.001365858, 0.001036216, 
    0.0007739161, 0.0006583245, 0.0005352875, 0.0004803124, 0.0004638143, 
    0.0004256152, 0.0003602535, 0.0003309302, 0.0003372074,
  0.001750177, 0.001819137, 0.001766281, 0.00133048, 0.001010331, 
    0.0007093762, 0.0006283787, 0.0006157032, 0.0004578153, 0.0003560875, 
    0.0004798109, 0.000459754, 0.000366375, 0.0003243907, 0.0003251439,
  0.00111781, 0.001255709, 0.001310091, 0.001158166, 0.0009967927, 
    0.0005496881, 0.0006264641, 0.0008827169, 0.00124621, 0.001112587, 
    0.0008985429, 0.001151221, 0.001217854, 0.0009927083, 0.0009104236,
  0.001317111, 0.001280582, 0.001311975, 0.001492234, 0.001223312, 
    0.0004590916, 0.0005358015, 0.0006158284, 0.0008930475, 0.001106367, 
    0.001213307, 0.001570572, 0.001578072, 0.001069962, 0.0008973698,
  0.001808091, 0.001528183, 0.001474429, 0.00162762, 0.001521996, 
    0.0006892555, 0.0004818226, 0.0005052597, 0.000579291, 0.0006709707, 
    0.0009520277, 0.001223143, 0.001436836, 0.001500944, 0.001301369,
  0.001983375, 0.001920858, 0.001806155, 0.001759692, 0.001729712, 
    0.001575775, 0.0005603743, 0.0004814407, 0.0005244231, 0.0005031041, 
    0.0005537754, 0.0008224495, 0.001040511, 0.001168082, 0.001122892,
  0.002024458, 0.001961735, 0.001883381, 0.001951863, 0.00176889, 
    0.001781991, 0.001497917, 0.0004587717, 0.0003173932, 0.0004150133, 
    0.000439359, 0.0005118366, 0.000696922, 0.0008662255, 0.001015644,
  0.002050909, 0.002017063, 0.001936559, 0.001972088, 0.002017697, 
    0.001750838, 0.001455763, 0.001192424, 0.0007396257, 0.0004971298, 
    0.000365536, 0.0004159934, 0.0004626866, 0.0005900572, 0.0007303155,
  0.002051453, 0.002048595, 0.001997766, 0.001920981, 0.001986589, 
    0.002014553, 0.001298648, 0.0009712565, 0.0007182927, 0.0006042273, 
    0.0004644264, 0.0003679558, 0.0003688473, 0.0004279824, 0.0005311299,
  0.002054484, 0.002063713, 0.002048116, 0.001945387, 0.001860833, 
    0.001858885, 0.001281658, 0.0008693836, 0.0006644891, 0.0006125896, 
    0.0005108429, 0.0003622507, 0.0003126371, 0.0003577459, 0.0004305893,
  0.002080595, 0.002103183, 0.002099436, 0.001993829, 0.001820431, 
    0.001705031, 0.001130497, 0.0007735031, 0.0005926779, 0.0005121005, 
    0.0004482247, 0.0003780789, 0.0003141874, 0.0003206725, 0.0003692629,
  0.002109462, 0.002135679, 0.002159531, 0.0019408, 0.001462594, 0.001261047, 
    0.0009249378, 0.0007551391, 0.0005181837, 0.0004485158, 0.0005280533, 
    0.000374547, 0.0003052806, 0.0002922487, 0.0003265309,
  0.001230475, 0.001203414, 0.001203597, 0.001264527, 0.001138255, 
    0.0006815317, 0.0005595648, 0.0006225819, 0.0009751492, 0.001187163, 
    0.001226355, 0.001338986, 0.001215216, 0.0007791803, 0.0007118567,
  0.00172923, 0.001272071, 0.001296159, 0.001363962, 0.001158862, 
    0.0005959668, 0.0005420545, 0.0005585329, 0.0006650078, 0.000893132, 
    0.001174107, 0.001396803, 0.001308426, 0.001117904, 0.0008857357,
  0.002119131, 0.001560262, 0.00134131, 0.001463989, 0.001316777, 
    0.0007599687, 0.000545878, 0.0004885035, 0.000529058, 0.0005966622, 
    0.0006988025, 0.0008423495, 0.0009332428, 0.0009482253, 0.0009212002,
  0.002135239, 0.002122917, 0.001785622, 0.00157733, 0.001509647, 
    0.001305247, 0.0007575731, 0.0005131818, 0.0005149741, 0.0004827103, 
    0.0005809863, 0.000630582, 0.0006406901, 0.0006386392, 0.0006250623,
  0.002243398, 0.002183509, 0.002007984, 0.001743691, 0.001599617, 
    0.001564817, 0.001420164, 0.0008547282, 0.0007477304, 0.000446454, 
    0.0004692003, 0.000520591, 0.0005618276, 0.0005566038, 0.0005661027,
  0.002356319, 0.002285663, 0.002187089, 0.00190301, 0.001722428, 
    0.001678037, 0.001672695, 0.001589797, 0.00107523, 0.0006749837, 
    0.0004264342, 0.0004313, 0.0004313913, 0.0004861394, 0.000526095,
  0.002443274, 0.002382699, 0.002331797, 0.002124125, 0.001893936, 
    0.00183077, 0.001711191, 0.001414555, 0.0009811968, 0.0006341342, 
    0.0004842067, 0.0004209684, 0.0003721169, 0.0004108412, 0.0004974366,
  0.002401232, 0.002409314, 0.002395139, 0.002282013, 0.002017599, 
    0.001860389, 0.001853379, 0.001239212, 0.0007419903, 0.0005785726, 
    0.0004488661, 0.0003899981, 0.000304478, 0.0003652088, 0.0004813352,
  0.002277443, 0.002353478, 0.002395521, 0.00234675, 0.002126766, 
    0.002021969, 0.001728747, 0.001044531, 0.000639692, 0.0005380626, 
    0.0004149127, 0.0003802309, 0.0002787624, 0.0003315173, 0.0004453424,
  0.002226796, 0.002323685, 0.002464361, 0.002342869, 0.002042459, 
    0.001930092, 0.001481556, 0.0008215974, 0.0005509335, 0.000463242, 
    0.000421913, 0.0003388217, 0.0002657373, 0.0002849407, 0.0003868696,
  0.002017991, 0.001870029, 0.001459422, 0.001225164, 0.0009337231, 
    0.0008392639, 0.0009618272, 0.001132891, 0.00124507, 0.001200785, 
    0.001184019, 0.001172165, 0.001089993, 0.0008049131, 0.0006287515,
  0.002215037, 0.001957225, 0.001448684, 0.001100042, 0.0007706279, 
    0.0006684245, 0.0008785174, 0.001061039, 0.001204199, 0.001288189, 
    0.001302832, 0.001300818, 0.001191158, 0.0006028782, 0.0006041392,
  0.002451937, 0.002137207, 0.001484349, 0.001181403, 0.0009129557, 
    0.000537499, 0.0006738589, 0.0008412594, 0.001040383, 0.00111911, 
    0.001161401, 0.001086162, 0.0009086547, 0.000767834, 0.000504423,
  0.002389753, 0.002379254, 0.001712484, 0.001274924, 0.001081256, 
    0.0009357628, 0.0005663992, 0.0006828886, 0.0007594756, 0.0008349826, 
    0.0008698109, 0.0007485589, 0.000696534, 0.0006407787, 0.0005229144,
  0.002295776, 0.002362304, 0.001839933, 0.001492798, 0.001146557, 
    0.00110511, 0.0009668241, 0.0005538448, 0.0005624032, 0.000571379, 
    0.000651039, 0.00066213, 0.0006462955, 0.0005988895, 0.0005458863,
  0.002239395, 0.00241837, 0.001915001, 0.001572488, 0.001312818, 
    0.001174659, 0.001103383, 0.001094191, 0.001009285, 0.0007001462, 
    0.0005604736, 0.000558293, 0.0005330345, 0.0005016355, 0.000522305,
  0.002270832, 0.002441358, 0.002066532, 0.001667642, 0.001580383, 
    0.001426633, 0.001279454, 0.001342387, 0.0009961835, 0.0006920836, 
    0.0005915611, 0.0005065778, 0.0004314363, 0.0004327528, 0.000511064,
  0.002298185, 0.002455521, 0.002154669, 0.001787172, 0.001631165, 
    0.001562684, 0.001468127, 0.00119555, 0.0008151279, 0.0006054206, 
    0.0004917046, 0.000403042, 0.0003251312, 0.0004113762, 0.0005133692,
  0.002362747, 0.002491688, 0.00225159, 0.001885046, 0.001716661, 
    0.001643978, 0.001552633, 0.001084001, 0.0006744064, 0.00051825, 
    0.0004050641, 0.0003257227, 0.0002758867, 0.0003681307, 0.0004773526,
  0.002498278, 0.002592649, 0.002464388, 0.002132835, 0.001734303, 
    0.001724698, 0.001472503, 0.0008466794, 0.0005312057, 0.000430539, 
    0.0003587687, 0.0002921286, 0.0002525074, 0.0003073652, 0.000427264,
  0.001951266, 0.002049258, 0.002012427, 0.001709447, 0.001087262, 
    0.0005869581, 0.0007672379, 0.0009931793, 0.001049459, 0.0008875585, 
    0.0008304305, 0.0007771081, 0.000721704, 0.0006445663, 0.0004865573,
  0.002213022, 0.0021945, 0.002088708, 0.001529562, 0.0008752351, 
    0.0004941225, 0.0006847664, 0.0009513267, 0.001112066, 0.001086662, 
    0.0009876962, 0.000941917, 0.0008608068, 0.0005629021, 0.0005015853,
  0.002326432, 0.00234272, 0.002025749, 0.001452598, 0.001004952, 
    0.0004918188, 0.0006125927, 0.0008932625, 0.001121092, 0.001214008, 
    0.001147341, 0.001030609, 0.0009225996, 0.0008401438, 0.0006355738,
  0.002392712, 0.002424931, 0.002203015, 0.001382795, 0.001126124, 
    0.001007062, 0.0005398131, 0.0008093247, 0.000960212, 0.001083471, 
    0.001039768, 0.0009073435, 0.0008340388, 0.000742292, 0.0005687833,
  0.002443549, 0.002424401, 0.002117525, 0.001462073, 0.001061822, 
    0.001086317, 0.00104511, 0.0005522514, 0.0005423598, 0.0007527765, 
    0.0008072983, 0.0007446968, 0.0007241724, 0.0006678167, 0.0006081357,
  0.00252843, 0.002438741, 0.001968428, 0.001441915, 0.001175751, 
    0.0009787232, 0.00107133, 0.001119119, 0.0008668688, 0.0007195615, 
    0.0006515793, 0.0006446354, 0.0006379443, 0.0006329961, 0.0006086548,
  0.002525654, 0.002341371, 0.001819815, 0.001456494, 0.001354163, 
    0.001234253, 0.001099505, 0.0009648922, 0.0007830376, 0.0006865684, 
    0.0005988221, 0.0005603948, 0.0005646744, 0.0005776195, 0.0005698181,
  0.002428381, 0.002218348, 0.001717926, 0.001487015, 0.00142532, 
    0.001400517, 0.001013978, 0.0008348034, 0.000667141, 0.0005907334, 
    0.0005009044, 0.0004710081, 0.0004400183, 0.0004990011, 0.0005431903,
  0.002318941, 0.002055935, 0.001683423, 0.001539757, 0.001515653, 
    0.001321558, 0.0008717534, 0.0007335859, 0.0005550496, 0.0004630602, 
    0.000398468, 0.0003746646, 0.0003469823, 0.0004458477, 0.0004792541,
  0.002244136, 0.002017824, 0.001753278, 0.001680854, 0.001202228, 
    0.001052038, 0.0007566992, 0.0006142239, 0.0004645511, 0.0003726457, 
    0.0003263428, 0.0003224973, 0.0002952228, 0.0003689563, 0.0004286015,
  0.002377272, 0.002460612, 0.002472619, 0.002422248, 0.002331149, 
    0.002034876, 0.001662813, 0.0014164, 0.001189913, 0.0008449402, 
    0.0007990356, 0.0007953385, 0.000721753, 0.0007075733, 0.0005932546,
  0.00264369, 0.002610534, 0.002499936, 0.002345009, 0.002022746, 0.00122084, 
    0.001068612, 0.000937066, 0.0009074023, 0.0008866591, 0.0008570227, 
    0.0008983294, 0.0008618737, 0.0006291463, 0.0005290802,
  0.002607807, 0.002490164, 0.002268687, 0.002018384, 0.001470515, 
    0.0008402144, 0.0008859165, 0.0009341282, 0.0008918006, 0.000920364, 
    0.000924224, 0.0009298891, 0.0009353556, 0.0009276645, 0.0007182309,
  0.002322913, 0.002186685, 0.001980103, 0.001656647, 0.001332643, 
    0.001016366, 0.0006535868, 0.000754795, 0.0007146394, 0.0007841114, 
    0.0008163132, 0.000882169, 0.0009519254, 0.0009444479, 0.0007577699,
  0.002050645, 0.00194738, 0.001823999, 0.001512928, 0.001202449, 0.00113792, 
    0.001055053, 0.0005494541, 0.0004064198, 0.000667811, 0.0007843638, 
    0.0008619613, 0.0009360203, 0.0009128299, 0.0007732642,
  0.001916088, 0.001740558, 0.001580448, 0.001380378, 0.001188335, 
    0.00108881, 0.001058543, 0.001014496, 0.0008737723, 0.0007329892, 
    0.0007466403, 0.000839707, 0.0008792908, 0.0008330938, 0.0007409381,
  0.001782773, 0.001624968, 0.001480635, 0.001336702, 0.001231214, 
    0.001085834, 0.0009620049, 0.0008906795, 0.0007808362, 0.0007552212, 
    0.0007684331, 0.000794357, 0.0007925308, 0.0007422456, 0.0006938882,
  0.001695895, 0.001586156, 0.001453183, 0.00134903, 0.001291174, 
    0.001154706, 0.0008386388, 0.0007542982, 0.0006996089, 0.0006959334, 
    0.000699502, 0.0007135955, 0.0006946589, 0.0006822253, 0.0006386921,
  0.00171947, 0.001614927, 0.001488826, 0.001345778, 0.001213772, 
    0.0009532992, 0.0007005081, 0.000633059, 0.0005949749, 0.0005966555, 
    0.0006010482, 0.0006041003, 0.0005842394, 0.0005696241, 0.0004761631,
  0.001759125, 0.001642888, 0.001468306, 0.0009917313, 0.0007952874, 
    0.0007179255, 0.0006230433, 0.0005543083, 0.0004933972, 0.0004714997, 
    0.0004788772, 0.0004989338, 0.0004637418, 0.0004401315, 0.0004080656,
  0.00161198, 0.00152262, 0.001312623, 0.001191315, 0.001208979, 0.001007911, 
    0.0008731415, 0.0008795007, 0.0009421796, 0.0009443749, 0.0009305333, 
    0.0009375758, 0.001014129, 0.001152883, 0.001108293,
  0.001719968, 0.001512815, 0.001289079, 0.001114953, 0.001024709, 
    0.0008692474, 0.0007634101, 0.0006631343, 0.0007696607, 0.0008354838, 
    0.0007905397, 0.0008675578, 0.0008311736, 0.0006534219, 0.0008228389,
  0.001879052, 0.001518154, 0.001252199, 0.001141159, 0.001006713, 
    0.0007384457, 0.000714926, 0.0006778566, 0.0007440093, 0.0008285051, 
    0.0008880025, 0.0008919197, 0.0008549558, 0.0008880214, 0.0008760106,
  0.001841984, 0.001591951, 0.001338691, 0.001172734, 0.001005043, 
    0.000895082, 0.000588421, 0.0005787453, 0.000651709, 0.0007975307, 
    0.0009094933, 0.0009642822, 0.0008858835, 0.0008855279, 0.0008636959,
  0.001867131, 0.001589751, 0.001395866, 0.001178148, 0.001015249, 
    0.0008894111, 0.0008551871, 0.0004309434, 0.0004687386, 0.0007242825, 
    0.0008770856, 0.0009336999, 0.0009453263, 0.0009137665, 0.0008566302,
  0.001891735, 0.001617021, 0.001401353, 0.001199572, 0.001019216, 
    0.0008485071, 0.0007976954, 0.0007501081, 0.0007347471, 0.0008630308, 
    0.0008613874, 0.0009531502, 0.0009742467, 0.000910331, 0.0008197959,
  0.001909434, 0.001666584, 0.001457695, 0.001249832, 0.001150178, 
    0.0009284234, 0.0007180147, 0.0007119391, 0.0007676648, 0.0009099395, 
    0.0009631139, 0.0009573855, 0.0009430978, 0.0008706667, 0.0008028957,
  0.001943578, 0.001732538, 0.001491085, 0.001276562, 0.001196458, 
    0.001003821, 0.0006711011, 0.0006492372, 0.0006523965, 0.000766155, 
    0.0008761779, 0.0009087939, 0.0008714325, 0.0007931128, 0.0007439881,
  0.002009646, 0.001747329, 0.001510915, 0.001228465, 0.00104588, 
    0.0007776379, 0.0006319786, 0.0006154765, 0.0005992246, 0.0006091037, 
    0.0006712403, 0.0006949503, 0.0006713447, 0.0006250993, 0.0005346395,
  0.002078133, 0.001829791, 0.001477004, 0.0008949405, 0.0006769074, 
    0.0006157926, 0.000596309, 0.0005928189, 0.0005406184, 0.0005000343, 
    0.0005078209, 0.0005506317, 0.0005387895, 0.0005141385, 0.0004752348,
  0.001904575, 0.001700556, 0.001287191, 0.00108416, 0.0009447274, 
    0.0006763662, 0.0006448628, 0.0006191005, 0.0007220629, 0.0007156762, 
    0.0007778588, 0.0008913815, 0.0008847368, 0.0008311799, 0.0008909944,
  0.002344269, 0.001828219, 0.001437836, 0.001108119, 0.0008851351, 
    0.00058777, 0.0006379056, 0.0006104137, 0.0007178515, 0.0008459137, 
    0.0008527303, 0.001007385, 0.0009855507, 0.0006878111, 0.0008527417,
  0.00256523, 0.001918092, 0.001502559, 0.001128744, 0.0009282115, 
    0.0005211084, 0.0006008879, 0.0006799973, 0.000802343, 0.0009250853, 
    0.0009933783, 0.001020287, 0.001005198, 0.00102627, 0.001095871,
  0.002667002, 0.002239703, 0.001679251, 0.001221667, 0.001002215, 
    0.0007709306, 0.0004845785, 0.0005627354, 0.0007387408, 0.0009341124, 
    0.001016791, 0.001027416, 0.001022507, 0.001039054, 0.000974199,
  0.002917876, 0.002465901, 0.001899651, 0.001327826, 0.0009981729, 
    0.0007837531, 0.0007315332, 0.0003949188, 0.0005626506, 0.0008525462, 
    0.0009708612, 0.0009968219, 0.001001771, 0.0009830057, 0.00095339,
  0.003147508, 0.002784358, 0.002142752, 0.001516102, 0.001118258, 
    0.0007729478, 0.0006979538, 0.0006550129, 0.0007342866, 0.0008608249, 
    0.0008497908, 0.0009412091, 0.0009659376, 0.0009298858, 0.0008830112,
  0.003385325, 0.003097618, 0.002529769, 0.001737368, 0.001316929, 
    0.000951752, 0.0006597834, 0.0006422239, 0.0006759538, 0.0007763018, 
    0.000789923, 0.0008324093, 0.0008548695, 0.0008367079, 0.0007972993,
  0.003596723, 0.00335516, 0.002905269, 0.002036594, 0.00145263, 0.001060254, 
    0.0006450261, 0.0006031657, 0.0005746305, 0.0006202371, 0.0006498238, 
    0.0006853257, 0.0006827031, 0.0006819282, 0.000654544,
  0.003766105, 0.003558737, 0.003205968, 0.002463904, 0.001605036, 
    0.000929892, 0.0006382565, 0.000588619, 0.0005281198, 0.0004803443, 
    0.0004983115, 0.000524291, 0.00054322, 0.0005428261, 0.0005006506,
  0.00382983, 0.003648069, 0.003301458, 0.002690512, 0.001616765, 
    0.0008104254, 0.0006350463, 0.0005950925, 0.0004701588, 0.000362481, 
    0.0003663411, 0.0004523518, 0.0004681914, 0.000500483, 0.0005369979,
  0.003589258, 0.003069437, 0.002029315, 0.001210774, 0.0007384885, 
    0.0005005234, 0.0004490084, 0.0005136208, 0.0008047348, 0.0007747687, 
    0.000839164, 0.0008885839, 0.0007288604, 0.0006563858, 0.000500523,
  0.003625028, 0.002969195, 0.00191801, 0.001053109, 0.000651792, 
    0.0004477979, 0.0004870332, 0.00054799, 0.0007652032, 0.0008776246, 
    0.0008716864, 0.00103134, 0.0009579335, 0.0005902865, 0.0004078005,
  0.003570673, 0.002922822, 0.001850368, 0.001109867, 0.0008131618, 
    0.0004212557, 0.0004882502, 0.0006148732, 0.0008229468, 0.0009352501, 
    0.0009844017, 0.0009857184, 0.0009332309, 0.0008288722, 0.000736375,
  0.003720038, 0.003166733, 0.002159022, 0.001264341, 0.0009979189, 
    0.0008042902, 0.0003991735, 0.0005547234, 0.000694942, 0.000880677, 
    0.0009906451, 0.0009842854, 0.0009531521, 0.0009088552, 0.0008709874,
  0.003822675, 0.003216115, 0.00245388, 0.00147421, 0.001023002, 
    0.0009139127, 0.0008544769, 0.0004120239, 0.0005758793, 0.0007091288, 
    0.0008699928, 0.0009327912, 0.0009279074, 0.0008776907, 0.0008289074,
  0.003676945, 0.00330786, 0.002504741, 0.00162269, 0.001065352, 0.000874456, 
    0.0008162895, 0.000740419, 0.0006554796, 0.0007345562, 0.0007138686, 
    0.0008219648, 0.0008333994, 0.0008074583, 0.0007896387,
  0.003508082, 0.003200477, 0.002615046, 0.001760387, 0.001340842, 
    0.0009664918, 0.0007317612, 0.0006362522, 0.0006000409, 0.0006258981, 
    0.0006418684, 0.0007248248, 0.0007551207, 0.000767266, 0.0007697839,
  0.003315809, 0.003048013, 0.002655256, 0.001879591, 0.001520713, 
    0.001157071, 0.0006955708, 0.0006118018, 0.0005282519, 0.0004954804, 
    0.0005113464, 0.000575135, 0.0006151578, 0.0006743719, 0.0006763285,
  0.003145999, 0.002927236, 0.002667387, 0.001962037, 0.001554668, 
    0.001011364, 0.0006577063, 0.0005855576, 0.0004999475, 0.000443556, 
    0.0004513534, 0.0005097114, 0.000556592, 0.0006258979, 0.000646026,
  0.002995629, 0.002824452, 0.002532064, 0.00184049, 0.001230859, 
    0.0008026839, 0.0006711447, 0.0006146083, 0.0005056271, 0.0004044014, 
    0.0004185672, 0.0005290192, 0.0005805603, 0.0006428482, 0.0006841128,
  0.001255018, 0.0009093675, 0.0007445657, 0.0006883454, 0.0006342211, 
    0.0005935621, 0.0006615885, 0.0005099822, 0.0006022456, 0.000483344, 
    0.0005514912, 0.0006168347, 0.0005494026, 0.0004742463, 0.0004158733,
  0.001248007, 0.0009356985, 0.0008560162, 0.0007714835, 0.000677385, 
    0.000583168, 0.0006787112, 0.0005917646, 0.0006511435, 0.0006116066, 
    0.0005973116, 0.0007013446, 0.0006462407, 0.0003732153, 0.0003301636,
  0.001388733, 0.001021122, 0.0009411006, 0.0009312864, 0.0008539097, 
    0.0004942897, 0.0006235373, 0.0006826836, 0.0008045384, 0.00076551, 
    0.0007886252, 0.0007603976, 0.000675754, 0.0005783097, 0.0004708465,
  0.001570508, 0.001420249, 0.001180646, 0.001009395, 0.0009780327, 
    0.0008895074, 0.000571051, 0.0006410636, 0.0007263173, 0.0008260168, 
    0.0008818401, 0.0008681336, 0.0007855933, 0.0007050644, 0.0006010926,
  0.001646094, 0.001515618, 0.001424808, 0.001113197, 0.00100811, 
    0.0009694459, 0.0009238906, 0.000473456, 0.0005685543, 0.0007456848, 
    0.0008294933, 0.0008772094, 0.0008875646, 0.0008214274, 0.0007281164,
  0.001694029, 0.001557105, 0.001426508, 0.001228462, 0.001036852, 
    0.0008974667, 0.0008602149, 0.0007865605, 0.0007412031, 0.0007979457, 
    0.0007704106, 0.0008046225, 0.0008427865, 0.000857919, 0.0007976487,
  0.00173406, 0.001633845, 0.001526002, 0.001390398, 0.001313244, 
    0.0009627344, 0.0008235078, 0.0007834432, 0.0007741686, 0.0008062471, 
    0.0008518521, 0.0008414565, 0.0008217331, 0.0008414877, 0.0008434146,
  0.00176361, 0.001690138, 0.001590522, 0.001485878, 0.001413299, 
    0.001102946, 0.0008423148, 0.000801545, 0.0007563161, 0.0007653222, 
    0.0008421252, 0.0009205008, 0.0008941888, 0.0008680509, 0.0008665102,
  0.001789516, 0.001713494, 0.001583008, 0.001444705, 0.001281998, 
    0.0009890303, 0.0008792453, 0.0008440876, 0.0007770695, 0.0007419059, 
    0.00075232, 0.0009055078, 0.000966591, 0.0009598053, 0.0009460416,
  0.001761584, 0.001639823, 0.001425969, 0.001126218, 0.0009487774, 
    0.0009372723, 0.0009029029, 0.0008675854, 0.0007636906, 0.0006830014, 
    0.0006785047, 0.0007725714, 0.0009372034, 0.001019817, 0.001004726,
  0.00105142, 0.001036399, 0.0009677032, 0.0009397966, 0.0008138882, 
    0.000596525, 0.0005749064, 0.0005388296, 0.0005682071, 0.0003881711, 
    0.0004031649, 0.0005273013, 0.0005557218, 0.0005850081, 0.0006507518,
  0.001268767, 0.001119935, 0.001024377, 0.0009547278, 0.000810696, 
    0.0005867769, 0.0006269817, 0.0005881778, 0.0006586338, 0.0005254174, 
    0.0004205755, 0.0005650694, 0.0006580129, 0.000425585, 0.0004741231,
  0.001425364, 0.001313517, 0.001123072, 0.0009607191, 0.0008870423, 
    0.0005390471, 0.0006079383, 0.000643442, 0.0006980151, 0.0006979576, 
    0.0006112571, 0.0005737077, 0.0006347052, 0.0006614095, 0.0006142684,
  0.001515536, 0.001461024, 0.001314152, 0.001009537, 0.0009176117, 
    0.0007990326, 0.0005342376, 0.0005604847, 0.0006848972, 0.0007065622, 
    0.00073349, 0.0006226744, 0.0006106888, 0.0006532872, 0.0006028943,
  0.001596784, 0.001534377, 0.001437653, 0.001121622, 0.0009268043, 
    0.0008234644, 0.0007550019, 0.0004222323, 0.0005040216, 0.0006843514, 
    0.0006794287, 0.0006940038, 0.0006253918, 0.0006314315, 0.0006325062,
  0.001640476, 0.001574459, 0.001440885, 0.00121165, 0.001025685, 
    0.0007941153, 0.0007278734, 0.0006424772, 0.0006453866, 0.0008102487, 
    0.0006088343, 0.0007462534, 0.000691171, 0.000630661, 0.0006041096,
  0.001671516, 0.001602279, 0.001496779, 0.001292141, 0.00118244, 
    0.0008373785, 0.0007167908, 0.0006447837, 0.0006449363, 0.0008030799, 
    0.0007929649, 0.0007522337, 0.0007310984, 0.0006750022, 0.0006006518,
  0.001652518, 0.001576993, 0.001456988, 0.00133398, 0.001199241, 
    0.0008802766, 0.0007178247, 0.0006323771, 0.0005646136, 0.0006271283, 
    0.0008480641, 0.0008376854, 0.0007273451, 0.0007312993, 0.0006529929,
  0.001596109, 0.001504444, 0.001349463, 0.001167079, 0.000931591, 
    0.0007139514, 0.0007034824, 0.0006648615, 0.0005592393, 0.0005570815, 
    0.0006404204, 0.0009047274, 0.0008828918, 0.0008025714, 0.0007480159,
  0.001467225, 0.001331734, 0.001125628, 0.0007582949, 0.0006021328, 
    0.0006007156, 0.0006111335, 0.0006904941, 0.000551102, 0.0004845251, 
    0.0005119936, 0.0006951869, 0.0009361113, 0.0009386976, 0.0008438092,
  0.0009472769, 0.0009058112, 0.0008424453, 0.0008046235, 0.0006714729, 
    0.0004789553, 0.0004532833, 0.0004814663, 0.0005243015, 0.0004612073, 
    0.0004474945, 0.0004602661, 0.000416672, 0.0004531701, 0.0004300257,
  0.00112471, 0.0009686805, 0.0008872023, 0.0008194909, 0.0007276097, 
    0.0004358596, 0.0004582766, 0.0004797229, 0.0005439153, 0.0005509281, 
    0.0004791189, 0.0005384573, 0.0006020165, 0.0004414637, 0.0003884858,
  0.00140199, 0.00109804, 0.0009082519, 0.000804381, 0.0007485097, 
    0.0004695918, 0.0004710156, 0.0005055488, 0.0005579318, 0.0005857142, 
    0.0006084812, 0.000600192, 0.0006162696, 0.0006550269, 0.000628482,
  0.00132285, 0.001197729, 0.001000918, 0.0008055926, 0.0007281876, 
    0.0006571552, 0.0004065652, 0.0004602324, 0.0005362362, 0.000676411, 
    0.0006951056, 0.0006681572, 0.0006391446, 0.0006660682, 0.0006511753,
  0.001353053, 0.001233696, 0.001083071, 0.0008270033, 0.0007284746, 
    0.0006391299, 0.0005751328, 0.000309832, 0.0003766604, 0.0006317717, 
    0.0007270314, 0.0006767458, 0.0006201423, 0.0006552034, 0.0007209104,
  0.001360598, 0.001263699, 0.001091609, 0.0008984182, 0.0007661585, 
    0.0006157244, 0.0005821352, 0.0005096999, 0.0005301441, 0.0006710888, 
    0.0006482523, 0.0006057793, 0.0005827729, 0.0006467005, 0.0006788574,
  0.001359199, 0.001277826, 0.001165542, 0.001010634, 0.0009232913, 
    0.0006304019, 0.0005787765, 0.0005414042, 0.0005737385, 0.0007257247, 
    0.0007235698, 0.0005722637, 0.0005432994, 0.0005882472, 0.0006154954,
  0.00132912, 0.001263879, 0.001194058, 0.001113118, 0.0009737053, 
    0.0006447543, 0.0005652161, 0.0005435412, 0.0005463476, 0.0006801374, 
    0.0007100469, 0.0006055965, 0.0005138205, 0.0005269899, 0.0005548963,
  0.001300915, 0.00123129, 0.001137088, 0.0009781546, 0.0007016059, 
    0.0005299671, 0.0005474304, 0.0005598607, 0.0005416375, 0.000625092, 
    0.0007151364, 0.0006809713, 0.0005238838, 0.0005280161, 0.0005096583,
  0.001287223, 0.001142804, 0.0009277884, 0.0005823972, 0.0004725026, 
    0.0004545295, 0.0004774937, 0.0006295143, 0.000553059, 0.0005149716, 
    0.0006038379, 0.0007391288, 0.0006383123, 0.000526719, 0.0005142727,
  0.0007476927, 0.0007859663, 0.0007243161, 0.0006722991, 0.0005794151, 
    0.0004700169, 0.0004394657, 0.0003957782, 0.0004030085, 0.0003610807, 
    0.0004430497, 0.0004599231, 0.0003918952, 0.0003850904, 0.000369333,
  0.0008772985, 0.0007997387, 0.0007759221, 0.0007044197, 0.0005811552, 
    0.000392423, 0.0004231266, 0.0004138559, 0.0004204716, 0.0004597994, 
    0.000481745, 0.0004958143, 0.0004923136, 0.0004165353, 0.0003264058,
  0.001055908, 0.0008112363, 0.0007659335, 0.0007607116, 0.0006635159, 
    0.0003706959, 0.000429914, 0.000436849, 0.0004318441, 0.0005013405, 
    0.000580008, 0.0005806905, 0.0005503968, 0.0005022069, 0.0004237457,
  0.001133015, 0.00100067, 0.0008926823, 0.00073253, 0.0006857108, 
    0.0006099236, 0.0003562837, 0.0004682188, 0.0005028166, 0.0005793279, 
    0.0006636269, 0.0006931036, 0.0006602438, 0.0006173151, 0.000546707,
  0.001124468, 0.001067062, 0.0009670703, 0.0007803343, 0.0007031055, 
    0.0006193497, 0.0005807237, 0.0002927426, 0.0003763178, 0.0006228992, 
    0.0007076288, 0.0007009389, 0.0006982088, 0.0006936839, 0.0006728509,
  0.001132765, 0.001065169, 0.0009743075, 0.0008376734, 0.0007573247, 
    0.0006230649, 0.0005956122, 0.0005531119, 0.0005376263, 0.0006107982, 
    0.0006058226, 0.0006587427, 0.0006804266, 0.0006646266, 0.0006625896,
  0.00112009, 0.001097358, 0.001020247, 0.000943715, 0.0008894454, 
    0.0006396307, 0.0005764881, 0.0005511024, 0.0005448625, 0.0006082985, 
    0.0006070001, 0.0005457225, 0.0005634956, 0.0006059438, 0.0006135138,
  0.001155886, 0.001103839, 0.001071601, 0.001032795, 0.0009487614, 
    0.0006710792, 0.0005725309, 0.0005485864, 0.0005099563, 0.0005177518, 
    0.0005154228, 0.0005217538, 0.0005580965, 0.0006185339, 0.0006138132,
  0.001193975, 0.001103297, 0.001085614, 0.0009997139, 0.0007915088, 
    0.0006350927, 0.0005763255, 0.0005804567, 0.0005315288, 0.0004975469, 
    0.0004650951, 0.0005158656, 0.0005255165, 0.0006032545, 0.0005852731,
  0.00118562, 0.00112228, 0.001046482, 0.0008395472, 0.0007333658, 
    0.0006575939, 0.0005942706, 0.0007116654, 0.0005852801, 0.0004201838, 
    0.000348485, 0.000433802, 0.0004956418, 0.0005744825, 0.0005707838,
  0.0007127001, 0.0006903253, 0.0006112379, 0.0005912379, 0.0004889209, 
    0.000364624, 0.0003956069, 0.0004099735, 0.0004389174, 0.000367658, 
    0.0004260733, 0.0004977189, 0.0004751761, 0.0005105597, 0.0005422946,
  0.0007820532, 0.0007415753, 0.0007228855, 0.0007143551, 0.0006069371, 
    0.0004485995, 0.0004584765, 0.0004583816, 0.0004758557, 0.0004419604, 
    0.0004372821, 0.0004773112, 0.0005041888, 0.0004258989, 0.0004209753,
  0.001174847, 0.0009620452, 0.0008692938, 0.0008848684, 0.0008246343, 
    0.0004927136, 0.0005040477, 0.0005278556, 0.0004917044, 0.000513681, 
    0.0005369427, 0.0005216391, 0.0005084919, 0.000495391, 0.0004467555,
  0.001450406, 0.001485385, 0.001509691, 0.00125653, 0.001163609, 
    0.0009840134, 0.0006179939, 0.0006023913, 0.0005800461, 0.0006076497, 
    0.0006214461, 0.0006288015, 0.0006050807, 0.0005796887, 0.0005021132,
  0.001503986, 0.001583698, 0.001663161, 0.001616116, 0.001532139, 
    0.001361678, 0.001141666, 0.0006468134, 0.0005346916, 0.0006526398, 
    0.0006986875, 0.0006778962, 0.0006618379, 0.0006534968, 0.000624544,
  0.001710644, 0.001825034, 0.001816887, 0.001795855, 0.001715303, 
    0.001472826, 0.001245672, 0.00101565, 0.0008045602, 0.0006928645, 
    0.0006843804, 0.000677089, 0.0006554977, 0.0006639578, 0.0006567809,
  0.001976311, 0.001994282, 0.001877939, 0.001729865, 0.001582378, 
    0.001356972, 0.001128341, 0.0009661631, 0.0007745828, 0.0006677688, 
    0.0006008255, 0.0005979902, 0.0006128644, 0.000633633, 0.0006460434,
  0.002149164, 0.002027142, 0.001780328, 0.001625856, 0.001470273, 
    0.001204902, 0.0009845544, 0.0008297953, 0.0006940794, 0.0006096539, 
    0.0005598153, 0.0005239526, 0.000520355, 0.0005645634, 0.0005991564,
  0.002159569, 0.001916633, 0.001725595, 0.001535237, 0.001263131, 
    0.001022503, 0.0008232666, 0.0007380693, 0.0006503778, 0.0005685089, 
    0.0005113709, 0.0004831067, 0.0004801393, 0.0005155943, 0.0005538065,
  0.002066573, 0.001864755, 0.001642146, 0.001338032, 0.001067784, 
    0.0008521616, 0.0006818335, 0.000676254, 0.0006028894, 0.000503752, 
    0.0004498713, 0.0004416149, 0.000431073, 0.0004580593, 0.0004945492,
  0.001185783, 0.001180058, 0.001209894, 0.001183774, 0.0009628521, 
    0.0006526145, 0.000574505, 0.0005062557, 0.0004780627, 0.0003626005, 
    0.0003912115, 0.00043643, 0.0003744526, 0.0003965333, 0.0003531089,
  0.001402697, 0.001342749, 0.001352541, 0.001418527, 0.001174317, 
    0.001014004, 0.000931195, 0.0008380773, 0.0006875253, 0.0006052094, 
    0.000582164, 0.0005881114, 0.0005515824, 0.000430297, 0.00038688,
  0.00177664, 0.001674295, 0.001778335, 0.002042238, 0.001785716, 
    0.001571573, 0.001224819, 0.0009615127, 0.0008598232, 0.0007974796, 
    0.0007187006, 0.0007229695, 0.0006510311, 0.0005742349, 0.0004950191,
  0.001748419, 0.00205356, 0.002476169, 0.002496722, 0.002303728, 
    0.001834846, 0.00107548, 0.0009316236, 0.0008767149, 0.000810112, 
    0.0007984892, 0.0007530668, 0.0007014382, 0.0007134379, 0.0006523159,
  0.002035195, 0.00238526, 0.002642585, 0.00254891, 0.002024498, 0.001560354, 
    0.001178064, 0.0006472599, 0.0006172406, 0.0007296733, 0.0007707749, 
    0.0007395913, 0.0007070366, 0.0007044058, 0.0006922607,
  0.002473089, 0.002631937, 0.002649725, 0.002246372, 0.001830969, 
    0.001433512, 0.00124088, 0.0009586959, 0.0007108211, 0.0005440969, 
    0.0005843801, 0.000580802, 0.0005765079, 0.0005975054, 0.0006343157,
  0.002657731, 0.002543022, 0.002204242, 0.001830234, 0.001616372, 
    0.001307917, 0.0009939063, 0.0007434878, 0.0005823079, 0.0004802371, 
    0.0004625547, 0.000476183, 0.0004807632, 0.0004888787, 0.0005265286,
  0.002530755, 0.002232945, 0.001933358, 0.001634933, 0.001377143, 
    0.0008507821, 0.0005911979, 0.0005086185, 0.0004810452, 0.0004544097, 
    0.0004534351, 0.0004607714, 0.0004623398, 0.0004484611, 0.000472496,
  0.002265769, 0.002036655, 0.001718097, 0.00135856, 0.0009106269, 
    0.000589897, 0.0004814447, 0.0004895604, 0.000510965, 0.0004844301, 
    0.0004653594, 0.0004433124, 0.000430438, 0.0004112076, 0.0004181283,
  0.002097805, 0.001785024, 0.001443688, 0.0009189653, 0.0006385842, 
    0.0004615872, 0.0004153854, 0.0005207103, 0.0005031731, 0.0004320835, 
    0.0004422799, 0.0004319599, 0.0003824356, 0.000358322, 0.000374336,
  0.001134202, 0.001088975, 0.001119272, 0.001158469, 0.001435994, 
    0.001574167, 0.001944311, 0.001628883, 0.001299222, 0.0009334955, 
    0.0008560192, 0.0007961497, 0.0005869456, 0.0005205133, 0.0004621269,
  0.001195608, 0.001185746, 0.001190973, 0.001342269, 0.001567886, 
    0.001613091, 0.001946123, 0.00149253, 0.001341195, 0.001125935, 
    0.001008449, 0.001006146, 0.0009199283, 0.0007543216, 0.0006903257,
  0.001385427, 0.001440848, 0.001573476, 0.001976928, 0.002204719, 
    0.001924371, 0.001431606, 0.001213441, 0.001038908, 0.0009102431, 
    0.0008385472, 0.0009021432, 0.0008654587, 0.0008353696, 0.0007485675,
  0.001611964, 0.001851562, 0.002312985, 0.00248649, 0.002124323, 
    0.001317915, 0.0008679762, 0.0008255879, 0.000777462, 0.0007167021, 
    0.0007187008, 0.0007303948, 0.0007364224, 0.0007664124, 0.0007809128,
  0.001870797, 0.002306619, 0.002595197, 0.001964329, 0.001104985, 
    0.0008807656, 0.0008309454, 0.0005485353, 0.0005534069, 0.000632481, 
    0.0007003968, 0.0007033886, 0.0006830906, 0.0007017827, 0.0007510424,
  0.002454967, 0.002708749, 0.002411936, 0.001424142, 0.0009844011, 
    0.0006473728, 0.0005706962, 0.0005276168, 0.000485547, 0.0004189049, 
    0.0004908352, 0.0005646378, 0.0005660814, 0.0005964296, 0.0006276412,
  0.002750733, 0.002540268, 0.001782308, 0.001109686, 0.0009213192, 
    0.0006178207, 0.0005086307, 0.0004676901, 0.0004372009, 0.0004105709, 
    0.0004093241, 0.0004176408, 0.0004361186, 0.0004419606, 0.0004499367,
  0.002573509, 0.001784062, 0.001201117, 0.0009803547, 0.0008843828, 
    0.0005893902, 0.0005084023, 0.0004925668, 0.0004770661, 0.0004552006, 
    0.0004416632, 0.0004353325, 0.0004289931, 0.0004248405, 0.0004270697,
  0.002079122, 0.001363251, 0.001070751, 0.0008714659, 0.0005976395, 
    0.0005311367, 0.0005177338, 0.000535309, 0.0005259035, 0.0004993952, 
    0.0004663066, 0.0004379739, 0.0004510054, 0.0004660822, 0.0004449423,
  0.001651964, 0.0010983, 0.0008748528, 0.0005978745, 0.0005703925, 
    0.000545315, 0.0005473082, 0.0005794812, 0.0005394064, 0.0004486525, 
    0.0004245633, 0.0004255733, 0.0004677036, 0.0005030665, 0.0004380641,
  0.001173823, 0.00119557, 0.001140871, 0.001101278, 0.001034363, 
    0.001032407, 0.001252667, 0.001407561, 0.001259979, 0.0009098929, 
    0.000678023, 0.0005410404, 0.0004641312, 0.0004747481, 0.0004611165,
  0.001358565, 0.001282357, 0.00121462, 0.00116216, 0.001031109, 0.001060379, 
    0.001302572, 0.001103654, 0.0007865817, 0.0006507816, 0.0005122678, 
    0.0004980351, 0.0004827795, 0.0004167954, 0.0004369623,
  0.001852906, 0.001570006, 0.001385774, 0.001357027, 0.001393193, 
    0.00130767, 0.001150428, 0.0009021197, 0.0006937459, 0.0005906138, 
    0.0005338745, 0.0005098424, 0.0004948027, 0.0004710268, 0.0004486278,
  0.001886868, 0.0019993, 0.001970454, 0.001953598, 0.001875336, 0.001663873, 
    0.000938239, 0.0007219878, 0.0006154592, 0.0005836037, 0.0005657987, 
    0.0005317205, 0.0005004573, 0.0004792694, 0.000447111,
  0.001827663, 0.001915903, 0.00207039, 0.002097425, 0.001762756, 
    0.001509792, 0.00111828, 0.000559333, 0.0004620798, 0.0005507903, 
    0.0005734633, 0.0005242006, 0.0004832358, 0.0004661984, 0.0004536381,
  0.001850314, 0.001999489, 0.002165223, 0.002130813, 0.001827117, 
    0.001407937, 0.001132915, 0.0007287192, 0.0005377593, 0.0004077468, 
    0.0004047026, 0.0004706768, 0.0004666906, 0.0004511181, 0.0004350398,
  0.002068688, 0.002250417, 0.002287293, 0.002014319, 0.001774267, 
    0.001321366, 0.0007893017, 0.0005428245, 0.0004780211, 0.0004504058, 
    0.000485172, 0.0004775341, 0.0004621043, 0.0004287164, 0.0004137484,
  0.002532829, 0.002514478, 0.002244606, 0.001922373, 0.001662571, 
    0.0008440498, 0.0005806817, 0.000521721, 0.0005342234, 0.000523204, 
    0.0005145639, 0.0004725125, 0.0004233554, 0.0004003675, 0.0004215407,
  0.002985447, 0.002732621, 0.002267346, 0.001689137, 0.001011543, 
    0.000666698, 0.000572257, 0.0005824763, 0.000588234, 0.000569593, 
    0.0004777662, 0.0004020531, 0.0003873868, 0.0004070091, 0.0004294726,
  0.002764169, 0.002568285, 0.001867664, 0.001055234, 0.0006958539, 
    0.0006063593, 0.0005423889, 0.0005784211, 0.000569283, 0.0004351789, 
    0.0003553139, 0.0003244683, 0.0003446025, 0.0004239017, 0.0004339685,
  0.001618509, 0.001604786, 0.001487517, 0.001415475, 0.001253158, 
    0.001193861, 0.001180086, 0.001100894, 0.001047695, 0.001023205, 
    0.001083143, 0.001128339, 0.001056614, 0.001012707, 0.0008568307,
  0.001658055, 0.00160139, 0.001509568, 0.001333365, 0.001175835, 
    0.001166566, 0.001216133, 0.001123305, 0.001081953, 0.001085454, 
    0.001007585, 0.0009468025, 0.0008918149, 0.0008002875, 0.0007032616,
  0.001838436, 0.00165808, 0.001497888, 0.00136668, 0.00124948, 0.001016094, 
    0.001167057, 0.001202184, 0.001123833, 0.001110341, 0.001035319, 
    0.0009434809, 0.0008657224, 0.00078679, 0.0007147373,
  0.001929171, 0.00204947, 0.001957939, 0.001631191, 0.001352071, 
    0.001311686, 0.0009577252, 0.001144065, 0.001214845, 0.00118412, 
    0.001111364, 0.001011891, 0.0008989797, 0.0007875301, 0.0006976629,
  0.001883972, 0.002029584, 0.002137972, 0.001921485, 0.001491762, 
    0.001446876, 0.001302398, 0.0009985052, 0.001013209, 0.001137557, 
    0.001205806, 0.001084109, 0.0009207477, 0.00079284, 0.0006902132,
  0.001836425, 0.001944036, 0.002086684, 0.002086374, 0.001818502, 
    0.001552898, 0.001466429, 0.001277108, 0.001162065, 0.0009539077, 
    0.0008674543, 0.0008892867, 0.0007827507, 0.0006787395, 0.0005834097,
  0.00185273, 0.00186792, 0.002016623, 0.002134689, 0.002111814, 0.001834795, 
    0.00162038, 0.00138005, 0.001124318, 0.0008811448, 0.0007811615, 
    0.0007001345, 0.0006341015, 0.0005194715, 0.0004560074,
  0.001867293, 0.001860435, 0.001973574, 0.002110713, 0.002160166, 
    0.002017752, 0.001716639, 0.001392132, 0.001084377, 0.0007876011, 
    0.0006733639, 0.0005670505, 0.0004722803, 0.0004192212, 0.000396189,
  0.001987596, 0.001994076, 0.002039595, 0.002124196, 0.002283034, 
    0.001992721, 0.001683063, 0.001230333, 0.0009435075, 0.0007232427, 
    0.0005411694, 0.0004322024, 0.0003754695, 0.0003438595, 0.0003502296,
  0.002253911, 0.0025854, 0.002681162, 0.002279871, 0.00198514, 0.001536062, 
    0.001170157, 0.0008811866, 0.000652167, 0.0004423143, 0.0003101931, 
    0.0002860843, 0.0002848745, 0.0003115495, 0.0003538645,
  0.001562689, 0.001701102, 0.001711679, 0.001679516, 0.001616721, 
    0.001551795, 0.001514963, 0.00150219, 0.001364917, 0.001112548, 
    0.001078314, 0.001055852, 0.000893097, 0.0008973491, 0.0008493119,
  0.001910079, 0.001933343, 0.001885808, 0.001760861, 0.001601021, 
    0.001536433, 0.001480716, 0.001419628, 0.001345228, 0.001220963, 
    0.001145974, 0.001132723, 0.001015381, 0.0008630692, 0.0008304362,
  0.002113204, 0.002000569, 0.001886614, 0.001832683, 0.001710236, 
    0.001391507, 0.001455267, 0.001383555, 0.001345525, 0.001227694, 
    0.001164962, 0.001114347, 0.001024917, 0.000934526, 0.0009010791,
  0.002049562, 0.001899793, 0.001958428, 0.001913768, 0.001770066, 
    0.001598771, 0.001158437, 0.001262758, 0.001256026, 0.001195564, 
    0.001156474, 0.001116408, 0.001053469, 0.0009584053, 0.0009443772,
  0.00188011, 0.001815823, 0.001924326, 0.001831242, 0.001647601, 
    0.001638331, 0.001377166, 0.001007052, 0.0009724052, 0.001101474, 
    0.00122572, 0.001183374, 0.001087241, 0.00100804, 0.0009942539,
  0.001857204, 0.001764979, 0.001880895, 0.001844025, 0.00158372, 0.0015457, 
    0.001440487, 0.001201064, 0.001044267, 0.0009477453, 0.001025646, 
    0.001101812, 0.001051643, 0.001037343, 0.001018805,
  0.001867739, 0.001859515, 0.001885935, 0.001879117, 0.001700384, 
    0.001467458, 0.001325895, 0.001155028, 0.001017319, 0.0009706746, 
    0.0009599163, 0.0009267731, 0.0009541257, 0.0009285128, 0.0009106674,
  0.001993923, 0.001945191, 0.001960201, 0.00193593, 0.001816634, 
    0.001421507, 0.001283425, 0.001136089, 0.001005227, 0.0009202053, 
    0.0008913222, 0.00091406, 0.0008220714, 0.0006740401, 0.0006283196,
  0.002167981, 0.002081863, 0.002021398, 0.001902972, 0.001726331, 
    0.001442484, 0.001301582, 0.001134009, 0.0009526518, 0.0007472433, 
    0.000549793, 0.000482239, 0.0004282456, 0.0003659039, 0.0003244541,
  0.002150861, 0.002127594, 0.001842553, 0.001456689, 0.00125909, 
    0.001055366, 0.0009048677, 0.0007629891, 0.0005504694, 0.0003646627, 
    0.0002880031, 0.0002554972, 0.0002509417, 0.0002574939, 0.0002877158,
  0.00200915, 0.002070203, 0.002150425, 0.002089427, 0.001948756, 
    0.001850852, 0.001864424, 0.001853494, 0.001773389, 0.001570214, 
    0.001448747, 0.001437854, 0.00130942, 0.001205854, 0.001151374,
  0.002211966, 0.002221346, 0.002164452, 0.001979098, 0.001861907, 
    0.001836016, 0.001822261, 0.001730084, 0.001804243, 0.001692819, 
    0.001548458, 0.001499953, 0.001413906, 0.001172013, 0.001023164,
  0.002122905, 0.002030504, 0.001885233, 0.001771245, 0.001733249, 
    0.001589667, 0.001722582, 0.001711139, 0.001657532, 0.001636984, 
    0.001503404, 0.001373847, 0.001295426, 0.001195336, 0.001088483,
  0.001862706, 0.001811649, 0.001753754, 0.001624199, 0.001613721, 
    0.001679997, 0.001356046, 0.001519093, 0.001440101, 0.001403628, 
    0.001317985, 0.001260525, 0.001210046, 0.001217222, 0.001110154,
  0.001803054, 0.001732609, 0.001671449, 0.001462049, 0.001388535, 
    0.001492345, 0.001503535, 0.001047958, 0.00107993, 0.001254798, 
    0.001281883, 0.001238718, 0.001170778, 0.001131919, 0.001099919,
  0.001744068, 0.001654921, 0.001550041, 0.001376143, 0.001193166, 
    0.001142047, 0.001243343, 0.001241482, 0.001181405, 0.001176075, 
    0.001182992, 0.001195337, 0.001133702, 0.001098558, 0.001026196,
  0.001689053, 0.001594314, 0.00149514, 0.00134683, 0.001172892, 
    0.0008746026, 0.0008825044, 0.0009400795, 0.0009772929, 0.001000851, 
    0.0009982605, 0.0009904896, 0.0009789701, 0.0009451128, 0.0009304158,
  0.00162223, 0.001518408, 0.001405494, 0.00132454, 0.001168985, 
    0.0007509262, 0.0007113471, 0.0006682614, 0.000665142, 0.0006477133, 
    0.0006426886, 0.0006454756, 0.0006361104, 0.0006383155, 0.0006425383,
  0.001589321, 0.001482243, 0.001303271, 0.001035923, 0.0006988005, 
    0.0006260394, 0.0005932684, 0.0005505145, 0.0004738886, 0.0004054906, 
    0.0003617326, 0.0003778269, 0.0003850802, 0.0003815368, 0.0003646968,
  0.001595886, 0.001442637, 0.001147851, 0.000664936, 0.0005134764, 
    0.000492795, 0.0005416108, 0.0005757877, 0.0004383535, 0.0003248964, 
    0.0002894695, 0.0003040963, 0.0003132532, 0.0003236656, 0.0003222699,
  0.001616202, 0.001571653, 0.001619623, 0.001453465, 0.001207544, 
    0.001113968, 0.001163232, 0.00115739, 0.001227333, 0.001307968, 
    0.001411922, 0.001513218, 0.001547079, 0.001528378, 0.001483219,
  0.001755969, 0.001667908, 0.001590975, 0.001414354, 0.001082351, 
    0.001014156, 0.001015925, 0.0009976722, 0.001069352, 0.001204596, 
    0.001378511, 0.001514595, 0.001574023, 0.001446622, 0.001397114,
  0.001838899, 0.001789445, 0.001588689, 0.001377493, 0.001049414, 
    0.0007766407, 0.0008550165, 0.0008791732, 0.0009590176, 0.001091756, 
    0.001252769, 0.001328092, 0.001386823, 0.00140453, 0.001344504,
  0.001710678, 0.001682668, 0.001695778, 0.001531525, 0.001145949, 
    0.0008886408, 0.0005974848, 0.0006934214, 0.0007763283, 0.0008788479, 
    0.0009959341, 0.001064723, 0.001136139, 0.001191114, 0.001243792,
  0.001849945, 0.001753894, 0.001701026, 0.001557517, 0.001170053, 
    0.0008696842, 0.000776166, 0.0004406858, 0.0005404717, 0.0007295326, 
    0.0008143427, 0.0008397487, 0.0008318122, 0.0008763185, 0.0009823535,
  0.00214639, 0.001985301, 0.001853147, 0.001644715, 0.001147585, 
    0.0007461557, 0.0006716647, 0.0006025126, 0.0005841639, 0.0005911464, 
    0.0005930309, 0.0006472765, 0.0006659396, 0.0007031218, 0.0007563367,
  0.002425057, 0.002294166, 0.002100929, 0.001808033, 0.00108677, 
    0.0006513441, 0.0005588297, 0.0005388401, 0.0005294294, 0.0005174655, 
    0.0004967056, 0.0004974261, 0.0005094977, 0.0005453097, 0.0006028753,
  0.002513856, 0.002479003, 0.002397169, 0.001732689, 0.001018104, 
    0.0006072327, 0.000506134, 0.0004758833, 0.0004722553, 0.0004442276, 
    0.0004180599, 0.0004391308, 0.000413207, 0.0004423693, 0.0004680846,
  0.002530378, 0.002445946, 0.002273294, 0.001485265, 0.0007753439, 
    0.0005946782, 0.0005316663, 0.0005233305, 0.0004660634, 0.0004085689, 
    0.0003758151, 0.0003838979, 0.0003614342, 0.0003768636, 0.0004076173,
  0.002389014, 0.002236757, 0.001928914, 0.001066398, 0.0006185776, 
    0.0005253216, 0.0005125692, 0.0005347712, 0.0004479248, 0.0003669451, 
    0.0003318708, 0.0003337054, 0.0003159243, 0.0003321831, 0.000355861,
  0.001855302, 0.001854481, 0.001732974, 0.001718594, 0.001550595, 
    0.001544665, 0.001665865, 0.001427633, 0.001231246, 0.001069057, 
    0.0009526201, 0.0008787776, 0.0007493514, 0.00068748, 0.0006553045,
  0.001680919, 0.001697893, 0.00171695, 0.001649395, 0.001526028, 
    0.001550788, 0.001486561, 0.001331054, 0.001183697, 0.001013698, 
    0.0009222465, 0.0008972461, 0.000776857, 0.0006229254, 0.0005537752,
  0.002134283, 0.001950938, 0.001649024, 0.00158552, 0.001386198, 0.00119833, 
    0.001303293, 0.001223762, 0.001060871, 0.001060044, 0.001036161, 
    0.0009214581, 0.0008296453, 0.0006990618, 0.000590514,
  0.001999314, 0.002090076, 0.002220287, 0.001948074, 0.00152587, 
    0.001427013, 0.001168743, 0.001202725, 0.001173876, 0.001005336, 
    0.0008652417, 0.0007437536, 0.0006798116, 0.0006172088, 0.000535182,
  0.002092271, 0.002035652, 0.002049127, 0.002060506, 0.001799362, 
    0.001873001, 0.001717727, 0.0008550609, 0.0005249445, 0.0006026519, 
    0.0006053452, 0.0005514427, 0.000525881, 0.0005036715, 0.0004909175,
  0.002475859, 0.002306752, 0.002081894, 0.001734473, 0.001422671, 
    0.001189084, 0.0008856113, 0.0006751373, 0.0005182089, 0.0004201543, 
    0.0003918975, 0.0004201351, 0.0004173164, 0.0004109128, 0.0004063049,
  0.002285682, 0.002094972, 0.001733978, 0.00126984, 0.0008836339, 
    0.000627514, 0.0005665803, 0.0004909714, 0.0004201322, 0.0003943295, 
    0.0003796548, 0.0003665536, 0.0003602002, 0.0003387986, 0.000337124,
  0.001937518, 0.001729091, 0.001492241, 0.001198793, 0.0008635374, 
    0.0005275501, 0.0004606892, 0.0004047815, 0.0003865637, 0.0003692772, 
    0.0003374303, 0.0003282063, 0.0002980219, 0.0003010376, 0.0003213861,
  0.001614163, 0.001448871, 0.001235784, 0.0009362221, 0.0005476989, 
    0.0004611766, 0.0004209042, 0.0004021406, 0.0003789979, 0.0003470253, 
    0.0003092822, 0.0002832384, 0.0002698074, 0.0002629448, 0.0002885758,
  0.0013947, 0.001227537, 0.0009444089, 0.0005306888, 0.0004514824, 
    0.0004293965, 0.0004155081, 0.0004220959, 0.0003815812, 0.0003086889, 
    0.0002878938, 0.0002783665, 0.0002583197, 0.0002496631, 0.0002646917,
  0.001932382, 0.001915655, 0.001834995, 0.001847892, 0.002122976, 
    0.002407313, 0.002506752, 0.002281505, 0.002095731, 0.001996711, 
    0.001885997, 0.001774678, 0.001625026, 0.001501591, 0.001325781,
  0.001972555, 0.001860923, 0.001787912, 0.001757113, 0.001711429, 
    0.001791282, 0.001958616, 0.001970024, 0.001920601, 0.00186793, 
    0.001735943, 0.001734376, 0.001588343, 0.001367504, 0.001228755,
  0.002096205, 0.001878737, 0.001733198, 0.001629255, 0.00148463, 
    0.001296064, 0.00140976, 0.00148897, 0.00156546, 0.001683839, 
    0.001693445, 0.001593295, 0.001486867, 0.001398088, 0.001254077,
  0.001972758, 0.002007284, 0.001944187, 0.001707951, 0.001427422, 
    0.001351848, 0.001211518, 0.001234843, 0.001243384, 0.00124668, 
    0.001196343, 0.001064278, 0.001009215, 0.0009128819, 0.0007688146,
  0.001983418, 0.001955418, 0.001917113, 0.001703513, 0.001395912, 
    0.001475684, 0.001358256, 0.0008129185, 0.0006479567, 0.0007083039, 
    0.0007568595, 0.0006577411, 0.0006191734, 0.0005738689, 0.0005244827,
  0.001796468, 0.001647751, 0.001485174, 0.001049733, 0.0008957943, 
    0.0008718789, 0.001000045, 0.0008812759, 0.0005933025, 0.0004803043, 
    0.0004456273, 0.0004759349, 0.0004415752, 0.000419398, 0.0003889808,
  0.001394043, 0.001294516, 0.001181058, 0.000770357, 0.0006970257, 
    0.0006086418, 0.0005941417, 0.0005484516, 0.000464637, 0.0004569755, 
    0.0004226055, 0.0003888772, 0.0003883868, 0.0003793274, 0.0003650816,
  0.001297012, 0.001205849, 0.001111315, 0.001003079, 0.0007982653, 
    0.0005397465, 0.000466812, 0.0004588169, 0.0004628115, 0.0004417224, 
    0.0004107972, 0.0003958303, 0.0003823647, 0.0003800735, 0.0003799452,
  0.001452232, 0.0013247, 0.001215851, 0.001061784, 0.0008992367, 
    0.0007304939, 0.0006251661, 0.0005717028, 0.0005406583, 0.0005349024, 
    0.0005256911, 0.0004878241, 0.0004654549, 0.0004462535, 0.0004191874,
  0.001676923, 0.001581049, 0.001422356, 0.001179871, 0.0009518731, 
    0.0008107287, 0.0006846017, 0.0006490113, 0.000647894, 0.0006303781, 
    0.0006723742, 0.0006308866, 0.0005710219, 0.0005657126, 0.0005358551,
  0.001501272, 0.001468065, 0.001520379, 0.001691663, 0.002348869, 
    0.002632697, 0.002823007, 0.002610797, 0.002766546, 0.002586555, 
    0.002484446, 0.002471447, 0.002397998, 0.002252834, 0.002188146,
  0.001610277, 0.001484912, 0.001498085, 0.001559053, 0.001798494, 
    0.002387932, 0.002719926, 0.002715463, 0.002756947, 0.002603479, 
    0.002496376, 0.002448273, 0.002334193, 0.002038314, 0.001953908,
  0.001628826, 0.001561156, 0.001528754, 0.001493815, 0.00155266, 
    0.001672618, 0.002357549, 0.002665851, 0.002711715, 0.002609442, 
    0.002509073, 0.002381782, 0.002248758, 0.002077942, 0.001798557,
  0.001620253, 0.001639907, 0.001669426, 0.001395267, 0.001434594, 
    0.001675793, 0.001785884, 0.002200027, 0.002413416, 0.002448658, 
    0.002420413, 0.002274133, 0.002150404, 0.001940036, 0.001641816,
  0.001577991, 0.001549921, 0.001644168, 0.001265737, 0.001207611, 
    0.001411592, 0.001707601, 0.001525521, 0.001486324, 0.002063721, 
    0.002193887, 0.002038965, 0.001937664, 0.001776971, 0.001555255,
  0.001584949, 0.001503318, 0.001545821, 0.001149422, 0.001055737, 
    0.001099864, 0.001273808, 0.00150531, 0.001536054, 0.001706961, 
    0.001772494, 0.001725873, 0.001670488, 0.00152999, 0.001320002,
  0.00171584, 0.001664452, 0.001577746, 0.001229304, 0.001013318, 
    0.0009102435, 0.0009763828, 0.001087834, 0.001312922, 0.001421757, 
    0.001406677, 0.001399077, 0.001368997, 0.001250788, 0.001046517,
  0.002048686, 0.001994323, 0.001941269, 0.001900124, 0.001264256, 
    0.000736066, 0.0007457, 0.0007848819, 0.000863355, 0.001040953, 
    0.001127656, 0.001114106, 0.001076723, 0.0009844197, 0.0008363031,
  0.002484252, 0.002380886, 0.002300918, 0.002208272, 0.001711428, 
    0.00092887, 0.0006938152, 0.0006595371, 0.0006984565, 0.000762736, 
    0.0008478194, 0.0008732556, 0.0008206152, 0.0007236667, 0.000622944,
  0.002909424, 0.002874445, 0.002817933, 0.002566969, 0.002232545, 
    0.001281854, 0.0007318272, 0.0006059899, 0.0005954569, 0.0005959725, 
    0.000701244, 0.00068583, 0.0006568912, 0.0006265602, 0.0005880228,
  0.001289906, 0.001255658, 0.001251492, 0.001595095, 0.001830421, 
    0.001962928, 0.00189761, 0.001626033, 0.001552858, 0.00182938, 
    0.001697461, 0.001985888, 0.002057586, 0.002054602, 0.001951292,
  0.001573623, 0.001485245, 0.001520146, 0.001813475, 0.001818821, 
    0.001914305, 0.001909669, 0.001558476, 0.001956345, 0.001884834, 
    0.001907609, 0.00216096, 0.002321516, 0.002235024, 0.001930478,
  0.002224303, 0.002054595, 0.001912797, 0.001919986, 0.001746428, 
    0.001944972, 0.002199905, 0.00181204, 0.002386512, 0.00240952, 
    0.002330519, 0.002296508, 0.002452688, 0.002387648, 0.002031932,
  0.00237501, 0.002272707, 0.002068495, 0.002058427, 0.001771274, 
    0.002045379, 0.001994814, 0.002091449, 0.002491836, 0.002538375, 
    0.002483061, 0.002347054, 0.002342816, 0.002126389, 0.001769356,
  0.002543003, 0.002380069, 0.002156141, 0.001943914, 0.001697778, 
    0.00190243, 0.00252789, 0.002225748, 0.002199574, 0.00245976, 
    0.002503055, 0.002265293, 0.002194421, 0.001873813, 0.001688511,
  0.002477386, 0.002349134, 0.002226893, 0.002000301, 0.001750335, 
    0.001695185, 0.002058839, 0.00231239, 0.002321468, 0.002363299, 
    0.002329949, 0.002278249, 0.001987127, 0.00160413, 0.00145682,
  0.002356744, 0.002303641, 0.002230599, 0.002212103, 0.001938253, 
    0.001559828, 0.001893553, 0.002145078, 0.002315389, 0.002380318, 
    0.002246492, 0.002182683, 0.001860562, 0.001547213, 0.001259693,
  0.002225541, 0.002213982, 0.002226747, 0.002294888, 0.002231118, 
    0.001370148, 0.001464265, 0.001736484, 0.002081525, 0.002231043, 
    0.002163038, 0.002115139, 0.001811119, 0.001433294, 0.001074302,
  0.001953676, 0.002037951, 0.002178127, 0.002396503, 0.002405486, 
    0.001702303, 0.001251206, 0.001596122, 0.001731258, 0.001955174, 
    0.002131807, 0.002056559, 0.001739202, 0.001269499, 0.0009575327,
  0.001474228, 0.001493304, 0.001566984, 0.001827142, 0.002434531, 
    0.001940074, 0.001269059, 0.001266229, 0.001484436, 0.001684483, 
    0.001950309, 0.001974977, 0.001644497, 0.001182686, 0.0009947596,
  0.001469133, 0.00147512, 0.001416744, 0.001427157, 0.001574161, 
    0.001395431, 0.001538369, 0.00154228, 0.00150291, 0.001449893, 
    0.001345726, 0.001523169, 0.001608673, 0.001590411, 0.00145265,
  0.001737019, 0.001648888, 0.00157771, 0.001523532, 0.001622669, 
    0.001335237, 0.001444849, 0.001431347, 0.001479243, 0.001247412, 
    0.001311454, 0.001571891, 0.001640227, 0.001597754, 0.00123431,
  0.001651511, 0.001746121, 0.001593882, 0.001557365, 0.001598157, 
    0.001386722, 0.001254685, 0.001159653, 0.00153002, 0.001463314, 
    0.001668728, 0.001792178, 0.001797274, 0.001743416, 0.001592195,
  0.001483597, 0.001595821, 0.001776655, 0.001796652, 0.001746238, 
    0.001743673, 0.001405112, 0.001314959, 0.001763823, 0.001821912, 
    0.001514651, 0.001637785, 0.001737708, 0.00186529, 0.001767373,
  0.001383469, 0.001404441, 0.0015902, 0.001640895, 0.001706095, 0.001877217, 
    0.001988612, 0.001676593, 0.00135326, 0.001593197, 0.001695068, 
    0.001778644, 0.001812488, 0.001854177, 0.00184993,
  0.00133017, 0.001272746, 0.001364724, 0.001528029, 0.00167064, 0.001887232, 
    0.002006815, 0.001887602, 0.001788595, 0.001911115, 0.00158323, 
    0.00171256, 0.001845838, 0.001920575, 0.001669098,
  0.001278256, 0.001210683, 0.001270369, 0.001393377, 0.001627917, 
    0.001757209, 0.001942873, 0.001589509, 0.001938684, 0.002037727, 
    0.00177111, 0.001751644, 0.001881697, 0.001673229, 0.001047367,
  0.001220783, 0.001194826, 0.00126751, 0.001423284, 0.001809582, 
    0.001630377, 0.001490707, 0.001752826, 0.001852543, 0.001961508, 
    0.001700129, 0.001747459, 0.001567974, 0.0009734753, 0.0005819513,
  0.001164704, 0.001189338, 0.001258757, 0.001214982, 0.001780295, 
    0.001894406, 0.001532192, 0.001649875, 0.001898079, 0.001810114, 
    0.001654196, 0.001548006, 0.0009925236, 0.0006347705, 0.0005317213,
  0.001054384, 0.001050233, 0.0009150985, 0.0008040927, 0.001570102, 
    0.001965982, 0.001687334, 0.001863836, 0.001671803, 0.001646563, 
    0.001486935, 0.001140509, 0.0007454238, 0.000621621, 0.0005720523,
  0.001366898, 0.001223002, 0.001072734, 0.001069749, 0.001285273, 
    0.001426008, 0.001262013, 0.001337208, 0.001395087, 0.001368782, 
    0.001421681, 0.001706009, 0.001556527, 0.001432359, 0.001362663,
  0.001595916, 0.001284278, 0.001158499, 0.001111875, 0.001235791, 
    0.001340474, 0.001408947, 0.001340795, 0.00145978, 0.001396867, 
    0.001316084, 0.001501994, 0.001506061, 0.001265824, 0.00110189,
  0.001622151, 0.001497368, 0.001295491, 0.00118165, 0.001141067, 
    0.001326708, 0.001299751, 0.001233293, 0.00119718, 0.001267695, 
    0.001364939, 0.001420215, 0.001397821, 0.001305944, 0.0009463158,
  0.001662177, 0.001620048, 0.001495635, 0.001367477, 0.001299495, 
    0.001485891, 0.001333454, 0.00117502, 0.001324963, 0.001441567, 
    0.001357645, 0.00134548, 0.00129403, 0.001137329, 0.0009040036,
  0.001690353, 0.001667194, 0.00164192, 0.001589173, 0.001509267, 
    0.001596516, 0.001742253, 0.0009969342, 0.001100532, 0.001243537, 
    0.001374345, 0.001339017, 0.001205726, 0.001057466, 0.0008863715,
  0.001683862, 0.001705018, 0.00173247, 0.001793041, 0.001778983, 
    0.001688812, 0.001776498, 0.00169512, 0.001418158, 0.00138699, 
    0.00127061, 0.001241017, 0.001105423, 0.0009175675, 0.000765547,
  0.001684148, 0.001730607, 0.001805892, 0.001872835, 0.001930677, 
    0.001609289, 0.001618392, 0.001517586, 0.001456057, 0.001366385, 
    0.001269602, 0.001139453, 0.0009057822, 0.0006810474, 0.0005831618,
  0.001641391, 0.001715352, 0.001798058, 0.00189769, 0.001983923, 
    0.001586007, 0.001417987, 0.001424843, 0.00129125, 0.001278426, 
    0.001102422, 0.0008350561, 0.0006123064, 0.000511993, 0.0004757053,
  0.001477172, 0.001518802, 0.001542234, 0.001442519, 0.00161681, 
    0.001629639, 0.001340487, 0.001321671, 0.001339649, 0.001062094, 
    0.0007937021, 0.0005978481, 0.0005054623, 0.0004879786, 0.0004895558,
  0.001250486, 0.001173395, 0.001036173, 0.000968173, 0.001238186, 
    0.001424755, 0.001389673, 0.001278979, 0.001158521, 0.0008588617, 
    0.0006194782, 0.0005086628, 0.0004917104, 0.0004990507, 0.0005351671,
  0.001701227, 0.001480503, 0.001329678, 0.001411367, 0.001322328, 
    0.001113446, 0.001037366, 0.001101859, 0.001194715, 0.00113643, 
    0.001078901, 0.001145563, 0.00105594, 0.0009325731, 0.0008364317,
  0.001997185, 0.001620613, 0.001509209, 0.001443892, 0.00125568, 
    0.0009745678, 0.0009884943, 0.001025568, 0.001021317, 0.001057311, 
    0.0009923457, 0.001086506, 0.001068076, 0.0008772452, 0.0008228284,
  0.00204276, 0.001916123, 0.0015966, 0.00151104, 0.001190495, 0.0009941995, 
    0.0008588873, 0.0009291168, 0.0008892458, 0.0009184621, 0.0009088746, 
    0.0009862023, 0.001042324, 0.00101074, 0.00087924,
  0.002000821, 0.0018915, 0.001728661, 0.001494418, 0.001281166, 0.001138585, 
    0.000737514, 0.0007679374, 0.0008050974, 0.0007943293, 0.000768607, 
    0.0008122115, 0.0009104088, 0.0009581269, 0.0009229483,
  0.001992926, 0.001838807, 0.001725049, 0.001454243, 0.001245386, 0.0011631, 
    0.001055663, 0.0006469615, 0.0006471236, 0.0007046797, 0.0006871711, 
    0.0006813119, 0.0007382489, 0.0007943358, 0.000855657,
  0.001967907, 0.001848037, 0.001706345, 0.001602102, 0.001354051, 
    0.001057793, 0.0009927112, 0.000916268, 0.0007500554, 0.0007131583, 
    0.00061602, 0.0006269886, 0.0006174822, 0.0006515139, 0.000725576,
  0.002030521, 0.001836901, 0.00178049, 0.001705862, 0.001479307, 
    0.0009688846, 0.0008003513, 0.0007472837, 0.0007008163, 0.000643192, 
    0.0005874408, 0.0005699864, 0.0005660331, 0.0005612036, 0.0005916686,
  0.002086368, 0.001845943, 0.001771703, 0.001796788, 0.001657562, 
    0.001041603, 0.0007386934, 0.0006247454, 0.0005628231, 0.000529632, 
    0.0004976849, 0.000514213, 0.0005204238, 0.0005310808, 0.000532061,
  0.002171193, 0.001870255, 0.001712812, 0.00144756, 0.001458305, 
    0.001363915, 0.0007914605, 0.0006184523, 0.000510825, 0.0004583677, 
    0.0004469074, 0.000468133, 0.0004757746, 0.0005093632, 0.0005419841,
  0.002306292, 0.001893607, 0.001544019, 0.001262419, 0.001212088, 
    0.001178715, 0.0008875637, 0.0006788526, 0.0005187768, 0.0004200174, 
    0.0004202041, 0.0004328925, 0.0004356935, 0.0004724289, 0.0005291961,
  0.002426483, 0.002184019, 0.001840585, 0.001756373, 0.001506625, 
    0.001160634, 0.0009979656, 0.0008786447, 0.0008275257, 0.0007846206, 
    0.0007819207, 0.0008875486, 0.0008174957, 0.0008072017, 0.0008634331,
  0.002813528, 0.00258749, 0.002201971, 0.001951502, 0.001679039, 
    0.001338503, 0.001141654, 0.0009908675, 0.0008975088, 0.0008664833, 
    0.0007694621, 0.0008644203, 0.0009052259, 0.0007156596, 0.0006721846,
  0.003087261, 0.002948059, 0.002559418, 0.002134769, 0.001702018, 
    0.001277189, 0.001145488, 0.0009845475, 0.0009060364, 0.000853295, 
    0.0007971501, 0.000812948, 0.0008956388, 0.000891675, 0.0007106186,
  0.003352122, 0.002988839, 0.002734477, 0.002282422, 0.001837267, 
    0.001469068, 0.001054167, 0.0009299014, 0.0008752279, 0.0008241546, 
    0.0007822719, 0.0007442016, 0.0008018165, 0.0008566714, 0.0008019963,
  0.003559967, 0.003024275, 0.002677623, 0.002268113, 0.001841787, 
    0.001476103, 0.001246002, 0.0007968053, 0.0006848703, 0.0007767662, 
    0.0007526199, 0.0007288347, 0.0007075435, 0.0007615671, 0.0008236152,
  0.003593361, 0.003052925, 0.002561921, 0.002210115, 0.001837872, 
    0.001475038, 0.001230718, 0.001133239, 0.001016297, 0.0009534345, 
    0.0007805986, 0.0007404403, 0.0006667647, 0.000667126, 0.0007245081,
  0.003528399, 0.002996152, 0.00245715, 0.00207941, 0.001748664, 0.001429942, 
    0.001218504, 0.001126906, 0.001056712, 0.0009651357, 0.0008343706, 
    0.0007577246, 0.0006647861, 0.0006149907, 0.0006559378,
  0.003272598, 0.002787567, 0.002292146, 0.001950787, 0.001652138, 
    0.001376276, 0.001195378, 0.001150362, 0.00108424, 0.001009643, 
    0.0009241706, 0.0007962871, 0.0006532774, 0.0005717099, 0.0005731959,
  0.002961244, 0.002499798, 0.002091164, 0.001669614, 0.001366597, 
    0.001194276, 0.00115329, 0.001192812, 0.001145913, 0.001069315, 
    0.0009738471, 0.0008267818, 0.0006480992, 0.0005664915, 0.0005642948,
  0.002588017, 0.002118487, 0.001656611, 0.001331012, 0.001109571, 
    0.0009948834, 0.001041744, 0.001200572, 0.001209131, 0.001088001, 
    0.0009785679, 0.0007978298, 0.0006202321, 0.0005579722, 0.0005643357,
  0.002381458, 0.002311113, 0.002025817, 0.001674186, 0.001397396, 
    0.001198036, 0.00115109, 0.001075659, 0.001022958, 0.0009479533, 
    0.0009206752, 0.0008544806, 0.0008302217, 0.00088703, 0.0008796356,
  0.002433849, 0.002189519, 0.001837226, 0.001427702, 0.001179524, 
    0.00099627, 0.0009881257, 0.0009592862, 0.000939671, 0.0009577281, 
    0.0008294196, 0.0008315044, 0.0008625963, 0.0008168729, 0.0008040164,
  0.002313565, 0.002049342, 0.001751827, 0.001308597, 0.001079469, 
    0.000906371, 0.0009240297, 0.0009409822, 0.0009138558, 0.0008542598, 
    0.0008321815, 0.0008246762, 0.0008501893, 0.0009144586, 0.0009322269,
  0.002148106, 0.001978993, 0.001720666, 0.001290945, 0.001063624, 
    0.0009434544, 0.0008390659, 0.0008963691, 0.00091502, 0.0009201762, 
    0.0008315232, 0.0008668842, 0.0008710459, 0.0009895741, 0.0009926412,
  0.002053336, 0.001878101, 0.00161551, 0.00120264, 0.0010418, 0.0009806207, 
    0.0009732083, 0.0008019479, 0.0008001304, 0.0009300669, 0.0008523688, 
    0.0008771872, 0.0009845401, 0.001010324, 0.0009846435,
  0.001998852, 0.001739231, 0.001483983, 0.001159166, 0.001031733, 
    0.0009993664, 0.001030801, 0.00105012, 0.001035453, 0.0009594786, 
    0.0007946916, 0.0008706744, 0.0009701864, 0.000985979, 0.0009612843,
  0.00202366, 0.001652123, 0.001475791, 0.001251077, 0.00103534, 
    0.0009450775, 0.001015663, 0.001057079, 0.001056952, 0.0009917065, 
    0.000864203, 0.0008662505, 0.0008943175, 0.0008750522, 0.0008353967,
  0.002187214, 0.001670753, 0.001465037, 0.001296831, 0.001067375, 
    0.0008850504, 0.0009409111, 0.0009973509, 0.0009886189, 0.0009664124, 
    0.0008463783, 0.0008507207, 0.0008097368, 0.000754579, 0.0007192733,
  0.002395898, 0.00178818, 0.001490186, 0.001040103, 0.0008926989, 
    0.0008304134, 0.0008794756, 0.000939025, 0.0009271708, 0.0008862674, 
    0.0008310952, 0.0007873147, 0.0007157063, 0.0006340183, 0.000580975,
  0.002500471, 0.00176265, 0.001303878, 0.0009665323, 0.0008685227, 
    0.0008005587, 0.0008029251, 0.0008999658, 0.0008502303, 0.0007340249, 
    0.0006664183, 0.0006656045, 0.0006041757, 0.0005829994, 0.0005629144,
  0.001807843, 0.00171226, 0.001494837, 0.00131263, 0.001256056, 0.001031374, 
    0.0009519373, 0.0009292764, 0.0008751422, 0.0008195394, 0.0009075223, 
    0.0007721221, 0.0006467634, 0.0006735134, 0.0006650802,
  0.002266464, 0.002076031, 0.001838311, 0.001542399, 0.001384671, 
    0.001122819, 0.001080238, 0.001004251, 0.0009311665, 0.0008983368, 
    0.0007891905, 0.000929145, 0.0009195214, 0.0007498228, 0.0006368427,
  0.002646487, 0.002457574, 0.002283731, 0.00193512, 0.001565538, 
    0.001179065, 0.001156416, 0.001080988, 0.0009843427, 0.0008943279, 
    0.0008632608, 0.000912889, 0.000951436, 0.0009559045, 0.0008162921,
  0.002966271, 0.002775615, 0.002631192, 0.002332673, 0.001972545, 
    0.001528078, 0.001147976, 0.001062424, 0.001039017, 0.0009403707, 
    0.0008446135, 0.0009097848, 0.0009357763, 0.0009585242, 0.0008994003,
  0.003336979, 0.003064611, 0.00292443, 0.00262837, 0.002311978, 0.001906152, 
    0.001435492, 0.000948988, 0.0008718135, 0.0009436118, 0.0008349803, 
    0.0007965808, 0.0008562281, 0.000895219, 0.0009248104,
  0.003730808, 0.003463379, 0.003164757, 0.002909397, 0.002619534, 
    0.002283076, 0.001838535, 0.001392983, 0.001148205, 0.0009625413, 
    0.0007863138, 0.0007294673, 0.0007140276, 0.0007539876, 0.000816178,
  0.004050678, 0.003808398, 0.003456576, 0.003122356, 0.002848433, 
    0.002519388, 0.002163731, 0.001785705, 0.001430624, 0.001099593, 
    0.0008437177, 0.0007288761, 0.0006585187, 0.000638188, 0.0006701946,
  0.004109637, 0.003937975, 0.003633127, 0.003314558, 0.003084707, 
    0.002762973, 0.002388754, 0.002066372, 0.001716985, 0.001327983, 
    0.0009201385, 0.0007219902, 0.0006357325, 0.0005859432, 0.0005937112,
  0.003981696, 0.003823163, 0.003696515, 0.003472788, 0.003238712, 
    0.002934335, 0.002611575, 0.00230042, 0.001965035, 0.00152579, 
    0.001046378, 0.0007485606, 0.0006158624, 0.0005499253, 0.0005613679,
  0.00373886, 0.003627535, 0.00357647, 0.003513188, 0.003306511, 0.003061768, 
    0.002747466, 0.002453114, 0.002139477, 0.001551147, 0.001037008, 
    0.0007409096, 0.0005788876, 0.0005012218, 0.0005484797,
  0.003039782, 0.003143935, 0.003230782, 0.003309397, 0.00327543, 
    0.003125571, 0.002939464, 0.002630468, 0.00216753, 0.00155164, 
    0.001417281, 0.001234595, 0.0009784758, 0.000855198, 0.0007424272,
  0.003199445, 0.003243058, 0.003364628, 0.003496706, 0.003502046, 
    0.003356119, 0.003183174, 0.002976918, 0.002661617, 0.002031914, 
    0.001602686, 0.001399206, 0.001213913, 0.0009695702, 0.0007992818,
  0.003257701, 0.003198595, 0.003293161, 0.003496765, 0.003602256, 
    0.003354675, 0.003255255, 0.003190382, 0.002935613, 0.00259175, 
    0.002086842, 0.001681851, 0.00138562, 0.001176427, 0.001007372,
  0.003284625, 0.003211682, 0.003208604, 0.00333975, 0.003510488, 0.00353364, 
    0.003245892, 0.003091688, 0.002897322, 0.002686673, 0.002308662, 
    0.001939571, 0.001573287, 0.001301151, 0.001116066,
  0.003280476, 0.003079166, 0.003084642, 0.00318459, 0.003296315, 
    0.003347311, 0.003354593, 0.002884774, 0.002728093, 0.002815018, 
    0.002707321, 0.002301766, 0.001824667, 0.001418756, 0.001165836,
  0.003224189, 0.002988904, 0.002904675, 0.002986986, 0.003034901, 
    0.003034179, 0.003086317, 0.003079589, 0.00305838, 0.002994138, 
    0.00281614, 0.002515943, 0.002038478, 0.001539976, 0.001182709,
  0.003184866, 0.002908331, 0.002784241, 0.002733841, 0.002744976, 
    0.002731574, 0.002756186, 0.002798702, 0.002829911, 0.002843668, 
    0.002700465, 0.002428773, 0.001904947, 0.001424226, 0.001104573,
  0.003145357, 0.002866529, 0.002666241, 0.00250769, 0.002436653, 
    0.002424855, 0.002459604, 0.002478877, 0.002462708, 0.002542973, 
    0.002495658, 0.002133447, 0.001532157, 0.001140925, 0.000974283,
  0.003120731, 0.002827301, 0.00254629, 0.002205284, 0.002078995, 
    0.002129753, 0.002142668, 0.002157434, 0.002135629, 0.002123259, 
    0.00197217, 0.001494478, 0.001095014, 0.0008993087, 0.0007654267,
  0.003034913, 0.002717449, 0.002294231, 0.001986517, 0.00179137, 
    0.001768697, 0.001754026, 0.001794661, 0.001733598, 0.001529932, 
    0.001308289, 0.0009828423, 0.0008018341, 0.00069244, 0.0006107542,
  0.003290345, 0.003113189, 0.002970607, 0.002680254, 0.002324362, 
    0.002101452, 0.002057592, 0.002221119, 0.002630728, 0.002663226, 
    0.0026674, 0.002463366, 0.00178674, 0.001335128, 0.001063517,
  0.00348314, 0.003247089, 0.003012241, 0.002675972, 0.002159468, 
    0.001780881, 0.001753255, 0.001835693, 0.00203182, 0.002244659, 
    0.002351667, 0.002432908, 0.002122417, 0.001490719, 0.001174407,
  0.003554555, 0.003258161, 0.0030493, 0.002755369, 0.002150547, 0.001515765, 
    0.001560203, 0.001507989, 0.001597456, 0.001907233, 0.002127567, 
    0.002353149, 0.002378064, 0.001982576, 0.001447893,
  0.003837175, 0.003533461, 0.003242569, 0.002858867, 0.002281076, 
    0.001654004, 0.001205862, 0.001309693, 0.001308664, 0.00147665, 
    0.001775212, 0.002155951, 0.002375337, 0.002331305, 0.001771063,
  0.004085165, 0.003684605, 0.003392687, 0.002988678, 0.002413993, 
    0.001702443, 0.001332475, 0.0009503568, 0.001049253, 0.001258852, 
    0.001558299, 0.001944292, 0.002279773, 0.002432766, 0.002214478,
  0.004314541, 0.00391165, 0.003466369, 0.003095657, 0.002642644, 
    0.001973698, 0.001406595, 0.001148761, 0.001002583, 0.001098995, 
    0.001348876, 0.00177244, 0.002132548, 0.002412803, 0.002237656,
  0.004481693, 0.00413052, 0.003690057, 0.003237618, 0.00282846, 0.00226195, 
    0.00165627, 0.00122131, 0.001009272, 0.0009745385, 0.001126235, 
    0.001485941, 0.001860042, 0.001929643, 0.001649989,
  0.00451214, 0.004207946, 0.003817244, 0.003381487, 0.002995802, 
    0.002482658, 0.001906655, 0.001367443, 0.001021784, 0.0008540834, 
    0.0009394719, 0.0009755394, 0.001082, 0.001121029, 0.001046193,
  0.004439234, 0.004174737, 0.003850784, 0.003441398, 0.003039799, 
    0.002575943, 0.002085807, 0.001572386, 0.001140725, 0.000876486, 
    0.0007988815, 0.0008655968, 0.0008007089, 0.0007620329, 0.000704928,
  0.004150582, 0.003930656, 0.003640061, 0.00329745, 0.002966932, 
    0.002620379, 0.002231156, 0.001803442, 0.00135993, 0.0009393427, 
    0.0007237231, 0.000689726, 0.0006633883, 0.000625178, 0.0006256519,
  0.003876847, 0.003589261, 0.003548523, 0.003654256, 0.003546953, 
    0.002952364, 0.002587354, 0.001988325, 0.001467971, 0.001409209, 
    0.001162834, 0.001463207, 0.001815837, 0.00188757, 0.001741795,
  0.003775412, 0.00349999, 0.003435762, 0.003525936, 0.003549115, 
    0.003065452, 0.002652216, 0.00205089, 0.001472416, 0.001357997, 
    0.001365385, 0.001511023, 0.001616865, 0.001712518, 0.001586549,
  0.003796358, 0.003374635, 0.003292936, 0.003362597, 0.003551943, 
    0.003054237, 0.002658116, 0.002200262, 0.001650481, 0.001464233, 
    0.001334151, 0.001474194, 0.001574416, 0.001846434, 0.001853191,
  0.003973646, 0.003560633, 0.003314929, 0.003221027, 0.003414456, 
    0.003455916, 0.002721781, 0.002139705, 0.001785131, 0.001582342, 
    0.001406944, 0.001324306, 0.001471221, 0.001711217, 0.001998225,
  0.004050054, 0.003580577, 0.003247915, 0.003088603, 0.003182963, 
    0.003373086, 0.003158822, 0.002146025, 0.00176124, 0.001858051, 
    0.001647323, 0.001386287, 0.001481641, 0.001601248, 0.001900605,
  0.004105685, 0.003687938, 0.003112264, 0.002900378, 0.002952159, 
    0.003093388, 0.003128912, 0.002869149, 0.002427235, 0.001950287, 
    0.00162577, 0.00143305, 0.001332489, 0.001517763, 0.001801864,
  0.004103205, 0.003741449, 0.003104147, 0.002703728, 0.002669055, 
    0.002743158, 0.002857841, 0.00284454, 0.00260294, 0.002149198, 
    0.001717938, 0.001419231, 0.001260192, 0.001339593, 0.001578777,
  0.004091356, 0.003697101, 0.003051713, 0.002552861, 0.00231704, 
    0.002374944, 0.002520517, 0.002616245, 0.00253084, 0.002148377, 
    0.00176327, 0.001461944, 0.001219653, 0.001061479, 0.001307776,
  0.00399728, 0.003615759, 0.002982126, 0.002287228, 0.002024538, 
    0.002016578, 0.002147352, 0.002244485, 0.002250283, 0.001979951, 
    0.001672085, 0.001458371, 0.001295087, 0.001069159, 0.0009389014,
  0.00381568, 0.003384754, 0.002768342, 0.002089716, 0.00172478, 0.001626145, 
    0.001764938, 0.001835079, 0.00186376, 0.001679825, 0.001474185, 
    0.001372483, 0.001262294, 0.001130617, 0.0009346181,
  0.003571734, 0.003316985, 0.00314422, 0.002750717, 0.00240088, 0.002484387, 
    0.00270734, 0.003053278, 0.00279535, 0.002232094, 0.001565275, 
    0.001385791, 0.001120465, 0.001470955, 0.001870107,
  0.003558639, 0.003361169, 0.00308127, 0.002541964, 0.002003448, 
    0.002047195, 0.002390611, 0.002772039, 0.002827407, 0.002438905, 
    0.001972489, 0.001659344, 0.001272951, 0.001198198, 0.001645613,
  0.003500998, 0.003272867, 0.002978675, 0.002412696, 0.001814874, 
    0.001791365, 0.002091391, 0.002425956, 0.002535632, 0.002385169, 
    0.002150039, 0.001967701, 0.001579317, 0.00133208, 0.001443357,
  0.003487808, 0.003274466, 0.002943645, 0.002264089, 0.001665194, 
    0.001655894, 0.001782764, 0.001915025, 0.002023682, 0.00209598, 
    0.00206391, 0.002062382, 0.001933185, 0.001580617, 0.001480198,
  0.003380563, 0.003123377, 0.002861609, 0.002125512, 0.001519271, 
    0.001419189, 0.001602834, 0.001476387, 0.001483834, 0.001807519, 
    0.001984891, 0.002017051, 0.002081044, 0.001911102, 0.001629503,
  0.003248968, 0.002982107, 0.002673606, 0.001985599, 0.001375065, 
    0.001163693, 0.00127083, 0.00132979, 0.001388074, 0.001449729, 
    0.001542696, 0.001664996, 0.001785393, 0.001901915, 0.001796752,
  0.003141603, 0.002835838, 0.002516739, 0.001839317, 0.001220549, 
    0.001006886, 0.0009940437, 0.0009951729, 0.001003334, 0.001023751, 
    0.001057374, 0.00119328, 0.001383047, 0.001545751, 0.00172424,
  0.003012037, 0.002633022, 0.002313109, 0.001605442, 0.00109624, 
    0.0008812035, 0.0008397801, 0.0007931886, 0.0007617666, 0.0007417716, 
    0.0007438876, 0.0008345159, 0.001024061, 0.001279636, 0.001487123,
  0.002820328, 0.002491243, 0.00207251, 0.001253147, 0.0009064778, 
    0.0008184955, 0.000775018, 0.0007334251, 0.0006794692, 0.0006521214, 
    0.0006132985, 0.0006418448, 0.0007421927, 0.001016258, 0.001231109,
  0.002544786, 0.002249935, 0.001694813, 0.001083715, 0.000853806, 
    0.0007574818, 0.0007248382, 0.0006756171, 0.0006131597, 0.0005458441, 
    0.0005124791, 0.0005417839, 0.0005891242, 0.0007818033, 0.001002458,
  0.001644808, 0.001305958, 0.001049229, 0.0009811468, 0.0009680468, 
    0.0009295014, 0.0008908338, 0.0009862294, 0.001120047, 0.001221972, 
    0.001373493, 0.001599346, 0.00167826, 0.001538307, 0.001363247,
  0.001841619, 0.001411724, 0.00105779, 0.0009232163, 0.0008502901, 
    0.0007121126, 0.0007502104, 0.0007685352, 0.0008001725, 0.000857058, 
    0.001018541, 0.001369725, 0.001472905, 0.001400027, 0.001312193,
  0.001800334, 0.001524498, 0.001303046, 0.0009317927, 0.0008141127, 
    0.0006227801, 0.0006685999, 0.0006436678, 0.00062056, 0.0006385393, 
    0.0006935248, 0.000972163, 0.00126503, 0.00138174, 0.001493831,
  0.001802726, 0.001524164, 0.001354987, 0.0009829275, 0.0008546578, 
    0.0007056865, 0.0005346184, 0.0005747867, 0.0005842895, 0.0005790457, 
    0.0005712454, 0.0006793141, 0.0009595053, 0.001234657, 0.001452172,
  0.001807857, 0.00152158, 0.001335564, 0.001026935, 0.0009307024, 
    0.0007196388, 0.0006386363, 0.000424308, 0.0004499831, 0.0005486591, 
    0.0005403392, 0.0005510286, 0.0006529355, 0.0009565349, 0.001330714,
  0.001815931, 0.001545394, 0.0013288, 0.001110489, 0.0009698277, 
    0.000755766, 0.0006586661, 0.0005790835, 0.0005028787, 0.000439567, 
    0.0004216223, 0.0004717033, 0.0005347132, 0.0006636381, 0.001063469,
  0.001811165, 0.001566654, 0.001351053, 0.001149694, 0.000968953, 
    0.0007781312, 0.0007025022, 0.0006317506, 0.000569412, 0.0004916659, 
    0.0004369909, 0.000434387, 0.0004872418, 0.0005428554, 0.0007575863,
  0.001797881, 0.001596456, 0.001371787, 0.001149502, 0.0009710077, 
    0.0008304517, 0.0007454034, 0.0006598338, 0.0005873609, 0.0005290566, 
    0.0004592189, 0.0004250442, 0.0004371836, 0.0004814427, 0.0006604188,
  0.001757639, 0.001600139, 0.001357507, 0.001112767, 0.0009663706, 
    0.0008443494, 0.0007258898, 0.000624066, 0.0005710716, 0.000516897, 
    0.000461027, 0.000412797, 0.0003962998, 0.0004478593, 0.0005854227,
  0.001699945, 0.00149644, 0.001247903, 0.001113616, 0.0009640587, 
    0.0008285373, 0.000695843, 0.0005904722, 0.0005358367, 0.0004473961, 
    0.0004146062, 0.0003999943, 0.0003701199, 0.0004180591, 0.0005290944,
  0.00190767, 0.00182861, 0.001697497, 0.001632659, 0.001613826, 0.001337132, 
    0.0009230187, 0.0006232899, 0.0005525102, 0.0004767743, 0.0004410334, 
    0.000535895, 0.0007844092, 0.001143021, 0.001534709,
  0.002257218, 0.00204217, 0.001819479, 0.001750365, 0.001661486, 
    0.001310462, 0.0008945783, 0.0006593763, 0.000596532, 0.0005623176, 
    0.0004302333, 0.0005033229, 0.0006014645, 0.0007145106, 0.001103414,
  0.002048596, 0.001879252, 0.001837254, 0.001800752, 0.001719477, 
    0.001125013, 0.0009817644, 0.0007794544, 0.0006875502, 0.0006003589, 
    0.0005360468, 0.0004748456, 0.0005619074, 0.0006809899, 0.0009284851,
  0.001913762, 0.001773174, 0.001695133, 0.001647163, 0.00167526, 
    0.001267494, 0.0008982548, 0.0008489216, 0.0007748932, 0.0007301033, 
    0.0006304782, 0.0004984356, 0.0004919597, 0.0005727548, 0.0007571938,
  0.001789882, 0.001638667, 0.001573689, 0.001518887, 0.001509258, 
    0.001413622, 0.001059746, 0.000735841, 0.0006216324, 0.0007595575, 
    0.0007268983, 0.0005726449, 0.0004562205, 0.0005060395, 0.0006219874,
  0.00168202, 0.0015039, 0.001397583, 0.001282385, 0.001236769, 0.001187584, 
    0.001133742, 0.0009214043, 0.0007659352, 0.0006488687, 0.0006246876, 
    0.0005681597, 0.0004708053, 0.000460681, 0.0005708817,
  0.001571119, 0.001411784, 0.001252448, 0.001091423, 0.000943481, 
    0.0009023575, 0.0009240006, 0.00080673, 0.0007262913, 0.000653553, 
    0.0006427145, 0.0005694383, 0.000488464, 0.0004363049, 0.0005362103,
  0.00150006, 0.001318227, 0.001131161, 0.0009193073, 0.0008082752, 
    0.0007301595, 0.0006835712, 0.0006710234, 0.0006208202, 0.0006082536, 
    0.0006097342, 0.0005626608, 0.0004918571, 0.0004310742, 0.0005238682,
  0.001423039, 0.001232773, 0.0009885681, 0.0007758633, 0.0007462507, 
    0.0006527046, 0.0006168975, 0.0005998996, 0.0005671842, 0.0005405249, 
    0.0005749537, 0.0005392884, 0.0004757093, 0.0004322263, 0.0004894037,
  0.001272057, 0.001023981, 0.0008254665, 0.0007081704, 0.0006733424, 
    0.0006270459, 0.0005900778, 0.0005750564, 0.0005391904, 0.0005120735, 
    0.0005369482, 0.0005064388, 0.0004410576, 0.0004097887, 0.000451037,
  0.001400018, 0.00139149, 0.001259903, 0.001213929, 0.001277425, 
    0.001494759, 0.001556923, 0.001348207, 0.001112914, 0.0008542673, 
    0.0007070147, 0.0005589618, 0.0006642734, 0.001032161, 0.001647825,
  0.00152797, 0.0013999, 0.001281855, 0.001181653, 0.001338838, 0.001490079, 
    0.001372477, 0.001164063, 0.0009669877, 0.0007418655, 0.000593851, 
    0.0005700403, 0.00073637, 0.001018405, 0.00151486,
  0.00134989, 0.001195028, 0.001122857, 0.001158699, 0.001357898, 
    0.001157956, 0.001141974, 0.0009173836, 0.0007485735, 0.0006342258, 
    0.0005890948, 0.0005704362, 0.0007377066, 0.001130308, 0.001601721,
  0.001274819, 0.001128968, 0.001047278, 0.001025297, 0.001128588, 
    0.001077511, 0.0007702378, 0.0007286791, 0.0006255739, 0.0005892835, 
    0.0005521876, 0.0005855267, 0.0007680571, 0.001100852, 0.001468016,
  0.001203559, 0.001042816, 0.0009380149, 0.0008270773, 0.0009391172, 
    0.0009655415, 0.0008659541, 0.0005795921, 0.0004815386, 0.0005954275, 
    0.0005803498, 0.0005697064, 0.0007155468, 0.00104457, 0.001367149,
  0.00118802, 0.00102883, 0.0008982109, 0.0007144334, 0.0007308106, 
    0.0008996845, 0.0009670362, 0.0008156862, 0.0006702113, 0.0006415723, 
    0.0005505196, 0.0005701453, 0.000675539, 0.0009978685, 0.001292989,
  0.001158669, 0.001060347, 0.0009726989, 0.0008350351, 0.0008264756, 
    0.0009409014, 0.001018211, 0.0008912592, 0.0007624577, 0.0006778945, 
    0.00063133, 0.0005899985, 0.0007143412, 0.001012572, 0.001299137,
  0.001151163, 0.001079287, 0.001006391, 0.0009089863, 0.0009404841, 
    0.0009768406, 0.0009571888, 0.0008404463, 0.0007062397, 0.0006545089, 
    0.0006007717, 0.0005957836, 0.0007421511, 0.001000811, 0.001255763,
  0.001106896, 0.001022819, 0.0008690823, 0.0007824085, 0.0009055233, 
    0.0009260441, 0.0008737325, 0.000745683, 0.0006563104, 0.0005941071, 
    0.0005493627, 0.0005736793, 0.0006984943, 0.0009704908, 0.001165337,
  0.0009945076, 0.000804599, 0.0007192523, 0.0006957232, 0.0007768238, 
    0.0008263242, 0.0007776055, 0.0007237532, 0.0006055292, 0.0005074374, 
    0.0005002827, 0.0005376404, 0.0006321866, 0.0009065329, 0.00118516,
  0.001034401, 0.001055592, 0.0009596502, 0.0008412446, 0.0008794856, 
    0.0008796429, 0.0008714689, 0.0008637072, 0.001063479, 0.001409666, 
    0.00161258, 0.001377993, 0.001169014, 0.00101096, 0.0008229619,
  0.001238875, 0.001148734, 0.001027727, 0.0008702846, 0.0009099949, 
    0.0009227512, 0.001038971, 0.001016089, 0.001188695, 0.001441363, 
    0.001502745, 0.001299668, 0.001139406, 0.0008379028, 0.0007645772,
  0.001237273, 0.001167428, 0.001089737, 0.0009076091, 0.0008843861, 
    0.0008201971, 0.001070736, 0.001119587, 0.001236216, 0.001423151, 
    0.001366949, 0.001199162, 0.001091724, 0.0009122733, 0.0008714764,
  0.001238869, 0.001194188, 0.00113326, 0.0009157935, 0.000881592, 
    0.0008376971, 0.0007500318, 0.0009447588, 0.00110769, 0.001233355, 
    0.001120166, 0.001054821, 0.00104808, 0.0009882838, 0.001009783,
  0.001240056, 0.001184394, 0.001120812, 0.0008967721, 0.0008516276, 
    0.0008370466, 0.0008078321, 0.0005567301, 0.0005761823, 0.0008904942, 
    0.0009217422, 0.0007665027, 0.0009419784, 0.001132901, 0.001153922,
  0.001249354, 0.00121533, 0.001122808, 0.0009330978, 0.0008497242, 
    0.0007687519, 0.0007451077, 0.0007404902, 0.0006085008, 0.0005823851, 
    0.0005713984, 0.0007236112, 0.001097428, 0.001278338, 0.001282173,
  0.001243348, 0.001221582, 0.001177367, 0.0009829332, 0.0008517843, 
    0.0007261246, 0.0006715029, 0.0006438607, 0.0006137009, 0.0005444862, 
    0.00063122, 0.0009619766, 0.001353006, 0.001495736, 0.001453166,
  0.001245347, 0.001239428, 0.00115243, 0.0009566618, 0.0007977359, 
    0.0007069603, 0.0006484597, 0.0006223857, 0.0005948172, 0.000679738, 
    0.0008896512, 0.001326223, 0.001555436, 0.001592943, 0.001588374,
  0.001155579, 0.001115378, 0.0009710206, 0.0008263192, 0.0007573419, 
    0.0006772476, 0.0006834587, 0.0006920794, 0.0007251316, 0.0008472528, 
    0.001162155, 0.001522094, 0.001595051, 0.001532747, 0.001486298,
  0.00102505, 0.0008584465, 0.0007708358, 0.0007497828, 0.0007291737, 
    0.0006973778, 0.0007198097, 0.0008167292, 0.0009016356, 0.0009919099, 
    0.001165804, 0.001385948, 0.001425983, 0.001464705, 0.001525458,
  0.001400537, 0.001130762, 0.0009126462, 0.0008348114, 0.0009494098, 
    0.001112406, 0.001350562, 0.001403357, 0.001378253, 0.001329444, 
    0.001313142, 0.001440554, 0.001617566, 0.001584261, 0.00156544,
  0.001621519, 0.00126982, 0.001001821, 0.0008828363, 0.0009582398, 
    0.001092337, 0.001360674, 0.001452238, 0.00151263, 0.001578733, 
    0.001763652, 0.001925451, 0.001841345, 0.001632531, 0.001652476,
  0.001491602, 0.001257436, 0.001105424, 0.0009100071, 0.0009303685, 
    0.0009886986, 0.001224161, 0.001340848, 0.001418798, 0.00145748, 
    0.001495443, 0.001601002, 0.001680644, 0.001696824, 0.001641309,
  0.001385191, 0.001206329, 0.001114854, 0.0009130169, 0.0009319472, 
    0.001028884, 0.00110198, 0.001180638, 0.001192288, 0.001239553, 
    0.001236226, 0.001272394, 0.00137108, 0.001460005, 0.001510655,
  0.00126401, 0.001171602, 0.001082409, 0.000899911, 0.0009131963, 
    0.0009641332, 0.001118504, 0.0009058382, 0.0009178494, 0.001122701, 
    0.001092402, 0.001029341, 0.001073889, 0.001175911, 0.001313361,
  0.001259493, 0.001176664, 0.001053731, 0.00093238, 0.0009225672, 
    0.0009143528, 0.0009626435, 0.0009458924, 0.0007828056, 0.0008486368, 
    0.0008829923, 0.0009648051, 0.0009874178, 0.0009996864, 0.001088727,
  0.00127878, 0.001200202, 0.001104464, 0.0009737898, 0.0009097174, 
    0.0009265571, 0.000941578, 0.0008734871, 0.0008049695, 0.000764017, 
    0.0007736592, 0.0008832732, 0.0009526635, 0.0009604666, 0.00104769,
  0.00125759, 0.001199468, 0.001107566, 0.0009508182, 0.0009088139, 
    0.000959714, 0.00105661, 0.001090862, 0.0009989265, 0.0008281903, 
    0.0008092371, 0.0007924899, 0.0008673089, 0.001006345, 0.001068001,
  0.001232714, 0.001152436, 0.0009533829, 0.0008569018, 0.0008802523, 
    0.0009283614, 0.001099031, 0.001191192, 0.001180597, 0.001084005, 
    0.001125232, 0.001110449, 0.001126133, 0.001085576, 0.001206647,
  0.001126584, 0.0009195128, 0.0008619379, 0.0008160305, 0.0008216816, 
    0.0008552846, 0.001074977, 0.001334811, 0.001416734, 0.001443293, 
    0.001496613, 0.001435477, 0.001423885, 0.001310806, 0.001331111,
  0.001249313, 0.001257483, 0.001153896, 0.001125771, 0.001229582, 
    0.001076905, 0.0009795481, 0.0009682788, 0.001126018, 0.001328143, 
    0.001338999, 0.001034625, 0.0007495118, 0.0008262652, 0.0008276614,
  0.001555387, 0.001476521, 0.001291156, 0.001159214, 0.001177554, 
    0.001018545, 0.0009814291, 0.0009433152, 0.0009921457, 0.001205993, 
    0.001328904, 0.001306093, 0.0008819611, 0.000720128, 0.0007491629,
  0.001521306, 0.001500939, 0.001444671, 0.001176944, 0.001051857, 
    0.000925357, 0.0009678291, 0.0009421946, 0.0009627182, 0.001014917, 
    0.001137851, 0.001443507, 0.00119267, 0.0009241049, 0.0008173009,
  0.001570038, 0.001527684, 0.001453408, 0.001209515, 0.001090627, 
    0.0009901354, 0.0008898249, 0.0008974616, 0.000956822, 0.001004654, 
    0.000961808, 0.001260574, 0.001544482, 0.001243409, 0.000996485,
  0.001599668, 0.001532565, 0.001433837, 0.001226271, 0.001126588, 
    0.001019011, 0.001019011, 0.0008436634, 0.0008880103, 0.001056124, 
    0.0009472661, 0.001056706, 0.00139599, 0.001429227, 0.001292743,
  0.001625134, 0.001555111, 0.001475515, 0.00131612, 0.00115666, 0.00103363, 
    0.001023357, 0.001102204, 0.001203041, 0.001106169, 0.0009101456, 
    0.0009771342, 0.001224922, 0.001480924, 0.001437394,
  0.00167946, 0.001651968, 0.001586126, 0.00140906, 0.001171784, 0.00104822, 
    0.001026136, 0.001141989, 0.001351707, 0.001223688, 0.0009932544, 
    0.0009561126, 0.001151123, 0.001406565, 0.001535985,
  0.001865505, 0.001846657, 0.0017643, 0.001478177, 0.001236918, 0.001036793, 
    0.000983173, 0.001160284, 0.001448185, 0.001375754, 0.001088568, 
    0.001000722, 0.001096562, 0.001326061, 0.001473071,
  0.002302455, 0.002209106, 0.001967799, 0.001582551, 0.001253256, 
    0.0009929057, 0.0009362854, 0.001159316, 0.001455396, 0.001514607, 
    0.001276609, 0.001103299, 0.001152156, 0.001291686, 0.001316047,
  0.00270017, 0.002395989, 0.002078322, 0.001639964, 0.001352292, 
    0.0009300431, 0.0008748749, 0.001138592, 0.001448575, 0.001617, 
    0.00144046, 0.001218242, 0.00128827, 0.001338915, 0.001346911,
  0.001284378, 0.001568092, 0.001744971, 0.001742869, 0.001675705, 
    0.001632506, 0.001539956, 0.001308693, 0.001065109, 0.001212723, 
    0.001116331, 0.001016268, 0.0009282693, 0.0009883634, 0.001035925,
  0.002169358, 0.002270683, 0.002164775, 0.002067037, 0.001998119, 
    0.001837339, 0.001720852, 0.001342084, 0.001003664, 0.001235298, 
    0.001161457, 0.001084816, 0.001016676, 0.0009105866, 0.0009474595,
  0.002510078, 0.002663171, 0.002654094, 0.002335898, 0.002089278, 
    0.001967084, 0.001874831, 0.001379339, 0.0009784348, 0.00129457, 
    0.001180998, 0.001187587, 0.001076083, 0.001099208, 0.0009871003,
  0.002914312, 0.002881221, 0.002760867, 0.002537093, 0.002432807, 
    0.002310597, 0.001834066, 0.00113217, 0.000911614, 0.001226493, 
    0.001217834, 0.001237748, 0.001159939, 0.001073361, 0.0009541531,
  0.003185764, 0.003051563, 0.002860496, 0.002693129, 0.002567156, 
    0.00223355, 0.001681461, 0.0007767713, 0.0007946956, 0.001172188, 
    0.001265256, 0.001291576, 0.001324086, 0.001106598, 0.001043228,
  0.003177981, 0.003085364, 0.002897626, 0.002744904, 0.00247161, 
    0.001958281, 0.001223891, 0.0009135256, 0.000949936, 0.001212212, 
    0.001246706, 0.001304081, 0.001479472, 0.001406849, 0.001211838,
  0.003175076, 0.003138476, 0.002974945, 0.002640017, 0.002175937, 
    0.001486321, 0.001061235, 0.001006868, 0.001082231, 0.001373188, 
    0.001260724, 0.001312767, 0.001483083, 0.001581136, 0.001535005,
  0.003296023, 0.003160228, 0.002917278, 0.002300079, 0.001725942, 
    0.001151911, 0.001015059, 0.001028723, 0.00112753, 0.001441296, 
    0.001271372, 0.001287644, 0.001403664, 0.001508903, 0.001612737,
  0.003352856, 0.00296998, 0.002641053, 0.00183779, 0.001370882, 0.001033843, 
    0.0009707122, 0.001079646, 0.001232314, 0.001425296, 0.001293534, 
    0.00130927, 0.001368242, 0.001467972, 0.001485913,
  0.003374136, 0.002752101, 0.002322861, 0.001759847, 0.001412822, 
    0.000924892, 0.0009329832, 0.001141986, 0.00128556, 0.001375769, 
    0.001295805, 0.001340687, 0.001432607, 0.001563936, 0.001447234,
  0.001998475, 0.002314961, 0.002556758, 0.002540882, 0.00248721, 
    0.002484994, 0.002559658, 0.002477501, 0.002158856, 0.001381967, 
    0.001031212, 0.001232639, 0.001222166, 0.00118544, 0.001146239,
  0.002932234, 0.002871537, 0.002628975, 0.002382956, 0.002099084, 
    0.002165242, 0.002333462, 0.002183055, 0.001719001, 0.001131991, 
    0.00103071, 0.001287189, 0.001280928, 0.00115736, 0.001136445,
  0.003112193, 0.002818367, 0.002496885, 0.002024746, 0.00182134, 
    0.001691838, 0.001802474, 0.001574978, 0.001135978, 0.001030647, 
    0.001191919, 0.001284089, 0.001329351, 0.001354576, 0.001331224,
  0.003061235, 0.002572264, 0.002249012, 0.001717596, 0.001502747, 
    0.001396901, 0.00116488, 0.001126714, 0.00091627, 0.001012909, 
    0.001116561, 0.001276416, 0.001322556, 0.001414155, 0.00136852,
  0.002956212, 0.002375514, 0.0019967, 0.001432494, 0.001271739, 0.001048106, 
    0.001029161, 0.0007515305, 0.0007205075, 0.001005924, 0.001163737, 
    0.001290554, 0.00134895, 0.001430978, 0.001529053,
  0.003035051, 0.00233738, 0.001893496, 0.001526291, 0.001334551, 
    0.001067003, 0.0009300863, 0.0009627963, 0.0009962447, 0.001044413, 
    0.001198598, 0.001274217, 0.001407, 0.001518862, 0.001538701,
  0.003229211, 0.002582107, 0.002152237, 0.001684969, 0.001435791, 
    0.001101285, 0.0009430086, 0.001002117, 0.001177998, 0.001253902, 
    0.00128788, 0.001391993, 0.001543464, 0.001614135, 0.001461962,
  0.003423722, 0.002751032, 0.002464822, 0.001970819, 0.00162273, 
    0.001136543, 0.000932932, 0.0010661, 0.001332735, 0.001374673, 
    0.001451472, 0.001552107, 0.001697867, 0.001671358, 0.001444669,
  0.003541504, 0.003165876, 0.002806206, 0.002298226, 0.001828848, 
    0.001207936, 0.0009220462, 0.001123178, 0.001398083, 0.001536121, 
    0.001584042, 0.001709006, 0.00174799, 0.001649103, 0.001539108,
  0.003675838, 0.003341851, 0.002839515, 0.002638722, 0.001956707, 
    0.001084597, 0.0008805208, 0.001212411, 0.00148187, 0.001571179, 
    0.00172617, 0.001812155, 0.001750797, 0.001606184, 0.001576289,
  0.002023255, 0.00156714, 0.001505291, 0.001352354, 0.001212348, 
    0.001175889, 0.001057032, 0.001149139, 0.001233234, 0.001295885, 
    0.001247931, 0.001269383, 0.001249059, 0.001192911, 0.001185439,
  0.002459365, 0.001984647, 0.001887767, 0.001723398, 0.00150707, 
    0.001182432, 0.00107554, 0.0009526468, 0.001046175, 0.001152562, 
    0.001197117, 0.001203155, 0.001149873, 0.001022776, 0.001053969,
  0.002725532, 0.002460827, 0.002437987, 0.002139937, 0.001836214, 
    0.001334287, 0.001050396, 0.0009954441, 0.001102077, 0.001209085, 
    0.001307325, 0.001334185, 0.001291022, 0.001265074, 0.001252035,
  0.003143962, 0.002956377, 0.002786584, 0.002444387, 0.002226264, 
    0.001725416, 0.001125923, 0.0009390645, 0.001147905, 0.001367634, 
    0.001456737, 0.001482422, 0.00145214, 0.001534939, 0.001603282,
  0.003673364, 0.003373599, 0.002933776, 0.002718107, 0.002455305, 
    0.001948854, 0.001156953, 0.0009456789, 0.001074393, 0.001503126, 
    0.001534402, 0.001531995, 0.001476295, 0.001517579, 0.001545466,
  0.004035862, 0.003568753, 0.002902469, 0.00292909, 0.002426534, 
    0.001874286, 0.001237738, 0.001325985, 0.001506072, 0.001610407, 
    0.001528266, 0.001486505, 0.001486655, 0.001431756, 0.001444416,
  0.004063688, 0.003353891, 0.002742673, 0.002918403, 0.002221111, 
    0.001583233, 0.001232001, 0.00144507, 0.001660802, 0.001579242, 
    0.001482416, 0.001480072, 0.001450513, 0.001487756, 0.001552948,
  0.003867687, 0.003105125, 0.002503014, 0.002644158, 0.001937414, 
    0.001351057, 0.001304501, 0.001587403, 0.001600618, 0.001474668, 
    0.001387623, 0.001412118, 0.001467121, 0.0015969, 0.001701906,
  0.003683982, 0.002988225, 0.002309989, 0.002213222, 0.001489916, 
    0.001156166, 0.001381414, 0.001621702, 0.001552125, 0.00137987, 
    0.00130355, 0.001348019, 0.001455705, 0.00161325, 0.001738066,
  0.003833327, 0.002932535, 0.002094037, 0.00186018, 0.001163545, 
    0.001145064, 0.001441595, 0.001645076, 0.001507482, 0.00127444, 
    0.001209779, 0.001285896, 0.001388901, 0.001533413, 0.001673669,
  0.002391356, 0.002624394, 0.00267193, 0.002402879, 0.002146144, 
    0.001896047, 0.001395901, 0.001289257, 0.001259055, 0.001331127, 
    0.001332062, 0.001379311, 0.001395414, 0.001206638, 0.0010891,
  0.002976497, 0.002997434, 0.002595461, 0.00224038, 0.002055267, 
    0.001598444, 0.001415577, 0.001157205, 0.001183074, 0.00122419, 
    0.001340362, 0.001384927, 0.001421232, 0.00131442, 0.001213562,
  0.003265969, 0.002817159, 0.002324073, 0.002158189, 0.001817216, 
    0.00148409, 0.001306112, 0.001220545, 0.001254023, 0.001304184, 
    0.001319208, 0.001352084, 0.001378661, 0.001328887, 0.001304108,
  0.003424564, 0.002719976, 0.002071502, 0.00202805, 0.001645992, 
    0.001400016, 0.001135199, 0.001199209, 0.001260131, 0.001307525, 
    0.001296729, 0.001348895, 0.001372512, 0.001373015, 0.001344785,
  0.003422529, 0.002532559, 0.00196223, 0.001897656, 0.001484763, 
    0.001357727, 0.001300355, 0.001006838, 0.001052418, 0.001268604, 
    0.001326761, 0.00138725, 0.001473137, 0.001530742, 0.001443243,
  0.003550394, 0.002436428, 0.001834546, 0.001836773, 0.001450569, 
    0.001321492, 0.001340733, 0.001250569, 0.001167518, 0.001204263, 
    0.001278947, 0.00142815, 0.001578106, 0.001612906, 0.001625269,
  0.003586102, 0.002437671, 0.001702973, 0.001775732, 0.001427899, 0.0013506, 
    0.001326216, 0.001240181, 0.00120937, 0.00123474, 0.00127775, 
    0.001414539, 0.00153822, 0.001657763, 0.001656834,
  0.003577456, 0.002505054, 0.001728736, 0.001582648, 0.001389392, 
    0.001471937, 0.00129899, 0.001226468, 0.001249312, 0.00126383, 
    0.001253236, 0.001349048, 0.001463529, 0.001602181, 0.001576254,
  0.003693986, 0.002737247, 0.001799097, 0.001424386, 0.001327593, 
    0.001415759, 0.001286364, 0.001265121, 0.001303656, 0.001293631, 
    0.001212656, 0.001263138, 0.001381033, 0.001551295, 0.001549174,
  0.003939443, 0.002864618, 0.001907922, 0.001514651, 0.00131124, 
    0.001414165, 0.001335373, 0.001339029, 0.001304406, 0.001148264, 
    0.001116435, 0.001206294, 0.001315865, 0.001509126, 0.001598881,
  0.001813841, 0.001673155, 0.001604198, 0.001214347, 0.001062315, 
    0.001014812, 0.000942568, 0.000973176, 0.001030535, 0.001106765, 
    0.001099233, 0.001076101, 0.001233467, 0.001212606, 0.00114514,
  0.002261061, 0.001868877, 0.001728663, 0.001337949, 0.001171186, 
    0.001054152, 0.001018593, 0.001038519, 0.001082849, 0.001086776, 
    0.001054364, 0.001089493, 0.001141719, 0.001165287, 0.001128158,
  0.002754187, 0.002226085, 0.001964876, 0.00146257, 0.001284166, 
    0.001095751, 0.001107941, 0.001098263, 0.001105138, 0.001164208, 
    0.001129727, 0.001107378, 0.001178474, 0.00119412, 0.001222799,
  0.003170833, 0.002677941, 0.002246505, 0.001790871, 0.001519443, 
    0.001332292, 0.001107432, 0.001148975, 0.001170891, 0.001204519, 
    0.001183136, 0.001123667, 0.001169567, 0.001186846, 0.00120774,
  0.003508218, 0.003108826, 0.002622003, 0.002193057, 0.001833153, 
    0.001528028, 0.001423411, 0.001042557, 0.001007011, 0.001242013, 
    0.001248181, 0.001173039, 0.001161256, 0.001147202, 0.001245497,
  0.003804522, 0.003453966, 0.002826938, 0.002506927, 0.002165718, 
    0.001839248, 0.001545916, 0.001399336, 0.001289748, 0.001259781, 
    0.001226734, 0.001190279, 0.001186192, 0.001145842, 0.001257964,
  0.004207509, 0.003882814, 0.003139538, 0.002741941, 0.002389005, 
    0.002017962, 0.001724042, 0.001583946, 0.001472315, 0.001426453, 
    0.001361657, 0.001251329, 0.001168959, 0.001167283, 0.001276913,
  0.004265041, 0.00397795, 0.003340093, 0.002900003, 0.002581197, 0.00231364, 
    0.002084364, 0.00188994, 0.001804825, 0.001705278, 0.001527816, 
    0.001307214, 0.001160203, 0.001194785, 0.00126086,
  0.004111379, 0.003888241, 0.003414546, 0.00307112, 0.002807352, 
    0.002594536, 0.002377647, 0.002238694, 0.002107314, 0.001925709, 
    0.001654679, 0.001341003, 0.00120226, 0.001179926, 0.001251903,
  0.00383683, 0.003575038, 0.003516774, 0.003360188, 0.003051528, 
    0.002866803, 0.002643678, 0.002534908, 0.002286805, 0.001978721, 
    0.001592398, 0.001275414, 0.001110811, 0.001144366, 0.001234491,
  0.002527491, 0.002457368, 0.002415891, 0.002236841, 0.002068738, 
    0.001718172, 0.001472396, 0.001307873, 0.00133375, 0.001294091, 
    0.001278337, 0.001088368, 0.001047212, 0.0009443313, 0.000808906,
  0.003113473, 0.002953666, 0.002709788, 0.002389435, 0.002058698, 
    0.001936346, 0.001572671, 0.001537516, 0.001578349, 0.00145545, 
    0.001443601, 0.001278873, 0.001182455, 0.00103791, 0.0009440678,
  0.003493187, 0.003356352, 0.003132513, 0.002586344, 0.002417365, 
    0.00202123, 0.002035638, 0.001995678, 0.001948176, 0.001891423, 
    0.001816872, 0.001664548, 0.001512131, 0.001296396, 0.001171717,
  0.003798401, 0.003701091, 0.003487866, 0.003041219, 0.002837692, 
    0.002314449, 0.002163875, 0.002252431, 0.002208471, 0.002179102, 
    0.002054609, 0.001876672, 0.001730429, 0.001617936, 0.00140694,
  0.004125405, 0.003773956, 0.003542385, 0.003285918, 0.003214238, 
    0.003114416, 0.002935791, 0.002444467, 0.002374289, 0.002576141, 
    0.002599271, 0.002495531, 0.002299577, 0.002087654, 0.001788216,
  0.004191882, 0.00394336, 0.003491971, 0.003292907, 0.003310276, 
    0.003387864, 0.003379035, 0.003309284, 0.003214867, 0.003098657, 
    0.00290982, 0.002730318, 0.002597849, 0.002469605, 0.002294212,
  0.004246153, 0.004002531, 0.003601486, 0.003366591, 0.0033944, 0.003457692, 
    0.003477975, 0.003348493, 0.00303218, 0.002771251, 0.002645263, 
    0.002575063, 0.002534931, 0.002462453, 0.002373618,
  0.004430218, 0.00411248, 0.003638614, 0.00348252, 0.003513137, 0.003480121, 
    0.003217819, 0.00275185, 0.002516235, 0.002449537, 0.002400849, 
    0.002306992, 0.002159549, 0.002078023, 0.002037905,
  0.004511569, 0.004070032, 0.003529842, 0.003503077, 0.003345692, 
    0.003002811, 0.002494274, 0.002230708, 0.00215098, 0.002033212, 
    0.001736051, 0.00167223, 0.001706582, 0.001701029, 0.001703236,
  0.004190269, 0.00358775, 0.003459896, 0.003268478, 0.002888601, 
    0.002246081, 0.0019602, 0.001837028, 0.001639183, 0.001321082, 
    0.001331301, 0.001449348, 0.001547823, 0.001552124, 0.001553173,
  0.003089791, 0.003062344, 0.003291399, 0.003169173, 0.003069167, 
    0.003006847, 0.002741517, 0.002364795, 0.002158037, 0.001968549, 
    0.002007035, 0.002125217, 0.00208184, 0.002038803, 0.001833428,
  0.003450035, 0.003378873, 0.003332552, 0.003238891, 0.003172205, 
    0.003122513, 0.002826588, 0.002516588, 0.002275845, 0.002162606, 
    0.002219636, 0.002317388, 0.002344375, 0.002130825, 0.001925909,
  0.003725162, 0.003534386, 0.003425117, 0.003197744, 0.00322898, 
    0.002824391, 0.002756483, 0.002602887, 0.002377816, 0.002374464, 
    0.00246907, 0.00265409, 0.002744669, 0.002712364, 0.002369458,
  0.00390259, 0.003661952, 0.003392256, 0.003103507, 0.003027616, 
    0.002712601, 0.002317614, 0.002245307, 0.002251758, 0.002324692, 
    0.002372374, 0.002527531, 0.002574861, 0.002560711, 0.002456039,
  0.004016749, 0.003503195, 0.003148127, 0.00279655, 0.002615192, 
    0.002442608, 0.002301953, 0.00188818, 0.001857546, 0.001965235, 
    0.001876703, 0.001788289, 0.00162483, 0.001576677, 0.001706136,
  0.00393835, 0.003396646, 0.002804197, 0.002457205, 0.002247379, 
    0.002019321, 0.001912359, 0.001870909, 0.001732385, 0.001330995, 
    0.001146833, 0.001079162, 0.001067226, 0.001057085, 0.001141633,
  0.003751064, 0.003147446, 0.002579495, 0.002073105, 0.001793469, 
    0.001542619, 0.001371736, 0.001290779, 0.00119742, 0.001121669, 
    0.001074792, 0.001019074, 0.001083054, 0.001049364, 0.001055211,
  0.003417548, 0.002800073, 0.002154458, 0.001631673, 0.00136346, 
    0.001187696, 0.001112101, 0.001116036, 0.001114423, 0.001076048, 
    0.001072708, 0.001097995, 0.001113584, 0.001098184, 0.001069541,
  0.002994095, 0.002392636, 0.001656274, 0.001237887, 0.001169352, 
    0.001108531, 0.001085862, 0.001148131, 0.001130524, 0.001082655, 
    0.001145249, 0.00114136, 0.001170747, 0.001146762, 0.001145797,
  0.002573732, 0.001962332, 0.001372958, 0.001161373, 0.001116759, 
    0.001088269, 0.001081124, 0.001169185, 0.001155029, 0.001119566, 
    0.001208185, 0.00119579, 0.001176507, 0.001136245, 0.001086292,
  0.002275156, 0.002163805, 0.002072692, 0.001930306, 0.001897784, 
    0.00172484, 0.001523917, 0.001434153, 0.001385237, 0.001442881, 
    0.001517997, 0.00163543, 0.001798438, 0.002037131, 0.002349679,
  0.002257053, 0.001985563, 0.001712458, 0.001604098, 0.001581147, 
    0.001364836, 0.001232469, 0.001180308, 0.001161088, 0.001195427, 
    0.001355339, 0.001474365, 0.001637766, 0.001778407, 0.002064809,
  0.00217343, 0.001935809, 0.001646587, 0.001280974, 0.001203475, 
    0.001046083, 0.001041243, 0.001068503, 0.001069015, 0.001079721, 
    0.001115754, 0.001195414, 0.00131184, 0.001525972, 0.001954511,
  0.002130368, 0.001886377, 0.001676706, 0.0012813, 0.00115919, 0.001034708, 
    0.0009119933, 0.0009372996, 0.001015363, 0.001088291, 0.001100053, 
    0.001080107, 0.001073384, 0.001185127, 0.001446238,
  0.002236358, 0.001940224, 0.001735382, 0.001363812, 0.001177444, 
    0.001098984, 0.000992923, 0.0008111458, 0.0009034763, 0.001099267, 
    0.001131737, 0.001060188, 0.001053995, 0.001036095, 0.001074252,
  0.002385544, 0.002146279, 0.001849164, 0.001481424, 0.001237177, 
    0.001117657, 0.001052883, 0.001087539, 0.001155409, 0.00108946, 
    0.00108897, 0.001033923, 0.001079639, 0.001039648, 0.00102211,
  0.002602299, 0.002354901, 0.001999134, 0.001580847, 0.001273019, 
    0.001128834, 0.001028907, 0.001113956, 0.001192561, 0.001176762, 
    0.001172967, 0.001097999, 0.001140206, 0.001154881, 0.001175266,
  0.002969422, 0.002685553, 0.002151284, 0.001665771, 0.001368999, 
    0.001237982, 0.001027783, 0.001101449, 0.001226221, 0.001217516, 
    0.001223686, 0.001137151, 0.001206649, 0.001267463, 0.001192394,
  0.003328756, 0.002960913, 0.002257935, 0.001838244, 0.0015319, 0.001331775, 
    0.001107182, 0.001170467, 0.00122252, 0.001216979, 0.001188269, 
    0.001146398, 0.001195814, 0.001228653, 0.001279751,
  0.003535126, 0.003018563, 0.002497492, 0.002189647, 0.001825214, 
    0.001499765, 0.001151378, 0.001192042, 0.001244309, 0.001197562, 
    0.001118049, 0.001105091, 0.001153351, 0.001246107, 0.001325401,
  0.002088611, 0.001889082, 0.001732109, 0.001644355, 0.001601057, 
    0.001556586, 0.001331683, 0.001146242, 0.001105627, 0.001146978, 
    0.001184955, 0.001039756, 0.001086657, 0.001209996, 0.001446452,
  0.002635509, 0.002422628, 0.002214942, 0.002055699, 0.001990179, 
    0.001794801, 0.001585154, 0.001357618, 0.001187353, 0.001122458, 
    0.00108771, 0.000972158, 0.001001475, 0.001179717, 0.001160617,
  0.002997889, 0.002778581, 0.002697467, 0.002478009, 0.002347904, 
    0.001993436, 0.001751881, 0.001527469, 0.001311625, 0.001172619, 
    0.001072314, 0.001018955, 0.00104181, 0.001192926, 0.001161464,
  0.003353157, 0.00317244, 0.00309931, 0.002962675, 0.002768512, 0.002437456, 
    0.001863447, 0.001494503, 0.001285308, 0.001194485, 0.001097431, 
    0.001005544, 0.001051017, 0.001186185, 0.001138107,
  0.003713883, 0.003501497, 0.003433964, 0.003285828, 0.003084493, 
    0.002767953, 0.002292796, 0.001506111, 0.001170783, 0.001205656, 
    0.001106254, 0.001006045, 0.00104705, 0.001198999, 0.001196657,
  0.003985651, 0.003818033, 0.003565831, 0.003447981, 0.003334455, 
    0.003042431, 0.00262265, 0.002106308, 0.001552897, 0.00123728, 
    0.001040177, 0.0009825873, 0.001019721, 0.001114572, 0.001262554,
  0.004215085, 0.004162035, 0.003857358, 0.0035711, 0.00347675, 0.003122103, 
    0.002724112, 0.002226562, 0.001532929, 0.001235048, 0.001067032, 
    0.00104947, 0.001025755, 0.001139157, 0.00125129,
  0.004340478, 0.004115218, 0.003866612, 0.003662394, 0.003514477, 
    0.003112758, 0.002672875, 0.002120843, 0.001526172, 0.001310537, 
    0.001142135, 0.00108764, 0.001073934, 0.001148304, 0.001183939,
  0.004394445, 0.00411048, 0.00365996, 0.003685364, 0.003416157, 0.002955082, 
    0.002643596, 0.002031868, 0.00154368, 0.001287581, 0.001110445, 
    0.001034306, 0.001042477, 0.001102298, 0.001123183,
  0.004054082, 0.003720462, 0.003642159, 0.003508436, 0.003146996, 
    0.002825821, 0.002478607, 0.001907096, 0.00142915, 0.00117037, 
    0.000943625, 0.0009712526, 0.0009741951, 0.001053143, 0.001098591,
  0.003316605, 0.003242862, 0.003205954, 0.003043729, 0.002915078, 
    0.002825421, 0.002774165, 0.002818791, 0.002687682, 0.002362258, 
    0.002162179, 0.001789002, 0.001409121, 0.001078899, 0.0009332568,
  0.003614429, 0.003479273, 0.003411839, 0.003311128, 0.003211683, 
    0.003067709, 0.002855476, 0.002840157, 0.002802695, 0.002527319, 
    0.002296814, 0.001915542, 0.001401177, 0.00105512, 0.0009192184,
  0.003872746, 0.003616328, 0.003453614, 0.003324543, 0.003169668, 
    0.002959545, 0.002909113, 0.002807936, 0.002643291, 0.002284567, 
    0.002053266, 0.001829657, 0.001336475, 0.001080282, 0.001033758,
  0.00409523, 0.003711479, 0.003480831, 0.003182641, 0.002928709, 
    0.002906713, 0.002595793, 0.002399398, 0.002145684, 0.001977051, 
    0.001836924, 0.001518738, 0.001198971, 0.001054074, 0.0009883011,
  0.004252407, 0.003624606, 0.003314298, 0.002907768, 0.002718565, 
    0.002646763, 0.002402562, 0.001819829, 0.001658491, 0.001680228, 
    0.001483047, 0.001285812, 0.001149878, 0.001024709, 0.0009891465,
  0.004174334, 0.003541705, 0.002991602, 0.002634201, 0.002441998, 
    0.002255805, 0.0020203, 0.001848633, 0.001532855, 0.001356212, 
    0.001292134, 0.001162513, 0.001113636, 0.001030223, 0.000981398,
  0.003996512, 0.003326204, 0.002831928, 0.002431377, 0.002215598, 
    0.001862157, 0.001671637, 0.001439824, 0.001296197, 0.001139879, 
    0.001102191, 0.001133841, 0.001098921, 0.001047604, 0.001035315,
  0.003794323, 0.003106876, 0.002609574, 0.002228387, 0.001859457, 
    0.001619915, 0.00148291, 0.001286793, 0.00121256, 0.001163115, 
    0.001094166, 0.001092502, 0.001131661, 0.001126762, 0.001066606,
  0.003512857, 0.00296363, 0.002248737, 0.001808619, 0.001562875, 
    0.001437893, 0.001346778, 0.001243431, 0.001198044, 0.001146145, 
    0.001066206, 0.001027543, 0.0009846304, 0.001036402, 0.001006943,
  0.003086281, 0.002482834, 0.001855139, 0.00151699, 0.001303939, 
    0.001168165, 0.001133308, 0.001167298, 0.001122908, 0.001009758, 
    0.0008898739, 0.0008993532, 0.0008513692, 0.0008725924, 0.0009107482,
  0.002112158, 0.002025351, 0.00199209, 0.001991922, 0.001804552, 
    0.001442884, 0.001308641, 0.001364847, 0.001515829, 0.00169786, 
    0.001927882, 0.002162898, 0.002252889, 0.002202434, 0.001924394,
  0.002213786, 0.0019155, 0.001719664, 0.001642483, 0.001626287, 0.001207977, 
    0.00111091, 0.001126486, 0.001202984, 0.001417874, 0.001751764, 
    0.002395248, 0.002420152, 0.002107078, 0.001833839,
  0.002215345, 0.001879044, 0.001662513, 0.001416462, 0.00133742, 
    0.001123555, 0.001045272, 0.00104386, 0.001100293, 0.001296857, 
    0.001605791, 0.002153061, 0.002511815, 0.002099404, 0.001725631,
  0.00220403, 0.001852011, 0.001641401, 0.001305677, 0.001199859, 
    0.001125003, 0.0009302668, 0.0009520866, 0.001012139, 0.001175334, 
    0.001445466, 0.001869816, 0.002021194, 0.001811325, 0.001604962,
  0.002195518, 0.001814386, 0.001627241, 0.001276664, 0.001183686, 
    0.001147424, 0.001128625, 0.0008704488, 0.0008685838, 0.001098815, 
    0.001248664, 0.001505821, 0.001652768, 0.001676182, 0.001662399,
  0.002249534, 0.001842345, 0.0015711, 0.001330138, 0.001167903, 0.001122033, 
    0.001107283, 0.001087512, 0.001010937, 0.001083683, 0.001144234, 
    0.001294004, 0.001443268, 0.00146719, 0.001419132,
  0.002188366, 0.001881118, 0.001562556, 0.001330525, 0.001143112, 
    0.001108559, 0.001115392, 0.001101837, 0.001117151, 0.001082114, 
    0.001101523, 0.001144501, 0.001167317, 0.001217375, 0.00120898,
  0.002055878, 0.001850958, 0.001509493, 0.00121781, 0.001123229, 
    0.001090585, 0.001096406, 0.001103805, 0.001100294, 0.00111279, 
    0.001063702, 0.001122186, 0.001111585, 0.001074134, 0.001054958,
  0.001914492, 0.001801158, 0.001368627, 0.001208049, 0.001117554, 
    0.001079565, 0.001107253, 0.001142058, 0.001161555, 0.001156429, 
    0.001104349, 0.001077056, 0.00104664, 0.001085487, 0.001012648,
  0.001732987, 0.001588756, 0.001414314, 0.001285519, 0.001146353, 
    0.001074743, 0.001089128, 0.001145332, 0.001150055, 0.001119274, 
    0.001059913, 0.0009797105, 0.0009745049, 0.000983621, 0.001023851,
  0.001679172, 0.001780919, 0.001763241, 0.001655435, 0.001516254, 
    0.001180697, 0.001038385, 0.0009391616, 0.000961786, 0.00109271, 
    0.001217247, 0.001498506, 0.001682949, 0.001789105, 0.001850318,
  0.002017917, 0.002043611, 0.001892881, 0.00172742, 0.001492274, 
    0.001144601, 0.001061305, 0.001008771, 0.0009871792, 0.001045103, 
    0.001256008, 0.001611962, 0.00187217, 0.001882194, 0.001808438,
  0.002122894, 0.002101155, 0.001964199, 0.001712205, 0.001417849, 
    0.001161212, 0.001033959, 0.001060092, 0.001008907, 0.001103056, 
    0.001267507, 0.001683382, 0.002063753, 0.002030218, 0.001998395,
  0.002184621, 0.00213365, 0.00195426, 0.00171077, 0.001432589, 0.001168063, 
    0.000929179, 0.0009950628, 0.001030483, 0.00113587, 0.00122307, 
    0.001587643, 0.002156883, 0.002257828, 0.002139231,
  0.002266129, 0.002145958, 0.001927171, 0.00163654, 0.001415567, 
    0.001178297, 0.001060827, 0.0008596627, 0.0008810684, 0.001106195, 
    0.001170049, 0.001375842, 0.00180469, 0.002196679, 0.002196921,
  0.002304009, 0.002159676, 0.001874744, 0.001611467, 0.001410088, 
    0.001219795, 0.001078297, 0.001086531, 0.001045468, 0.001074033, 
    0.001111134, 0.001198873, 0.001367457, 0.001647701, 0.001842292,
  0.002344368, 0.002175437, 0.001861978, 0.001561204, 0.001385767, 
    0.001213452, 0.001093246, 0.001103285, 0.001083104, 0.001059547, 
    0.001095768, 0.001149626, 0.001215679, 0.001272944, 0.001358372,
  0.002356185, 0.002184846, 0.001814315, 0.001528045, 0.001364583, 
    0.001202239, 0.001135946, 0.001121759, 0.001111621, 0.001062975, 
    0.001044737, 0.001077571, 0.001170244, 0.001216416, 0.001261017,
  0.00241369, 0.002146902, 0.001740605, 0.001495152, 0.00134824, 0.001193293, 
    0.001147731, 0.00111769, 0.001124391, 0.001089169, 0.001040789, 
    0.001032359, 0.001100803, 0.001188036, 0.001279438,
  0.002387988, 0.00207011, 0.001720521, 0.00144877, 0.00130935, 0.001179261, 
    0.0011719, 0.001135518, 0.001150108, 0.001122801, 0.001071163, 
    0.001040273, 0.001051586, 0.001140214, 0.001292879,
  0.002513873, 0.002019904, 0.001494236, 0.001362816, 0.001316584, 
    0.001178481, 0.0009689892, 0.0009492526, 0.0009257091, 0.001059558, 
    0.001111491, 0.001171298, 0.001325354, 0.001638255, 0.002319196,
  0.002856578, 0.001966121, 0.001483622, 0.001284458, 0.001248119, 
    0.001061839, 0.0009741609, 0.0009923939, 0.0009856843, 0.000969036, 
    0.00108708, 0.001226756, 0.001390542, 0.001480873, 0.001764344,
  0.002788247, 0.001847394, 0.001480999, 0.001232771, 0.001143947, 
    0.001031945, 0.000983858, 0.001048906, 0.00107165, 0.001095958, 
    0.001111416, 0.001320398, 0.001447933, 0.001529124, 0.001588603,
  0.002675972, 0.001800342, 0.001454622, 0.001183063, 0.001163282, 
    0.001010616, 0.000910688, 0.001015262, 0.00108037, 0.00118359, 
    0.001228863, 0.001297792, 0.001474046, 0.001692746, 0.001610446,
  0.002535899, 0.001703167, 0.001414929, 0.001171876, 0.001131305, 
    0.001104724, 0.001016128, 0.0008869951, 0.0009368843, 0.00119089, 
    0.001295642, 0.001367456, 0.001442706, 0.001692899, 0.001899888,
  0.002380907, 0.001736355, 0.001368934, 0.001192774, 0.001088912, 
    0.001140061, 0.001125127, 0.001139718, 0.001185254, 0.001239235, 
    0.001323538, 0.001486391, 0.001489011, 0.001454965, 0.001827017,
  0.002317294, 0.001776998, 0.001397994, 0.001096426, 0.001064089, 
    0.001130338, 0.00116449, 0.001179067, 0.001237883, 0.001278466, 
    0.001361794, 0.001553543, 0.001735025, 0.001528315, 0.001472588,
  0.002315565, 0.00174034, 0.001285327, 0.001065308, 0.001059695, 
    0.001120517, 0.001207852, 0.001217677, 0.001246427, 0.001283475, 
    0.001362625, 0.001595727, 0.001881753, 0.001928199, 0.00164336,
  0.002376448, 0.00168685, 0.001190006, 0.001060377, 0.001074791, 
    0.001129219, 0.001239163, 0.001249817, 0.001272326, 0.001283139, 
    0.001365865, 0.001581501, 0.00192424, 0.002221371, 0.00198861,
  0.002341127, 0.001643556, 0.00122997, 0.001058908, 0.001073046, 
    0.001170115, 0.00124712, 0.001280236, 0.001300511, 0.001281986, 
    0.001352875, 0.001532073, 0.001831562, 0.002246997, 0.002473737,
  0.002545594, 0.001973592, 0.001334874, 0.001106348, 0.0009596135, 
    0.001036458, 0.001144084, 0.001283406, 0.001305224, 0.001349244, 
    0.001346905, 0.001307174, 0.001403751, 0.001767377, 0.00254773,
  0.002521872, 0.001706239, 0.001282613, 0.001104207, 0.001080704, 
    0.001041221, 0.001252958, 0.00131847, 0.001339242, 0.001195192, 
    0.001314774, 0.001434882, 0.001405521, 0.001607577, 0.002257475,
  0.00234039, 0.001745107, 0.001370355, 0.001193699, 0.001092609, 
    0.001042142, 0.001263085, 0.001406889, 0.001427427, 0.001443578, 
    0.00137303, 0.001548441, 0.001482924, 0.001582883, 0.002204563,
  0.002127491, 0.001648354, 0.00139211, 0.001151705, 0.001156335, 0.00117889, 
    0.001207837, 0.001328975, 0.001382257, 0.001556683, 0.001640862, 
    0.001681907, 0.001580736, 0.001412424, 0.001985078,
  0.001940224, 0.001533414, 0.001345312, 0.00115997, 0.001183195, 
    0.001256459, 0.001330745, 0.001152625, 0.001189043, 0.001593252, 
    0.001855679, 0.001941612, 0.001713806, 0.001305563, 0.001809848,
  0.001823569, 0.001523036, 0.001283528, 0.001161015, 0.001172055, 
    0.001256349, 0.001312617, 0.001367062, 0.001432377, 0.001661927, 
    0.001957875, 0.002090184, 0.001829187, 0.00151951, 0.001664354,
  0.001823901, 0.001522593, 0.001304742, 0.001102851, 0.001173982, 
    0.001239272, 0.001283118, 0.001363279, 0.001451257, 0.001686074, 
    0.002000308, 0.002205826, 0.00194824, 0.001593145, 0.001535404,
  0.001830714, 0.001499363, 0.001235619, 0.001067548, 0.00117606, 
    0.001255796, 0.001265635, 0.001279355, 0.001356204, 0.001580551, 
    0.001920978, 0.00218701, 0.002130589, 0.00170481, 0.001561729,
  0.00188642, 0.001538226, 0.001102449, 0.001057876, 0.001158063, 
    0.001260272, 0.001258052, 0.00126495, 0.001334358, 0.001523204, 
    0.00177858, 0.002085257, 0.002321579, 0.00198175, 0.001505485,
  0.001867031, 0.001427026, 0.001100454, 0.001054694, 0.001147041, 
    0.00124091, 0.001215285, 0.00122684, 0.001260031, 0.001378825, 
    0.001633417, 0.00188525, 0.002225895, 0.002452051, 0.001735073,
  0.001754438, 0.001623175, 0.001374, 0.001190187, 0.001184169, 0.001096533, 
    0.001207395, 0.001313829, 0.001511873, 0.001683138, 0.001825141, 
    0.001850044, 0.001801091, 0.001786592, 0.001792526,
  0.001694921, 0.001495331, 0.00134004, 0.001272886, 0.001247138, 
    0.001175779, 0.001333977, 0.001505283, 0.001662763, 0.001616128, 
    0.001916132, 0.001946086, 0.00187844, 0.001652287, 0.001774404,
  0.001689009, 0.001566485, 0.001423216, 0.001360094, 0.001255261, 
    0.001147688, 0.00137181, 0.001526546, 0.001699106, 0.001925117, 
    0.002028772, 0.001911236, 0.00178589, 0.001695176, 0.002031141,
  0.00159135, 0.001566428, 0.001473104, 0.001354554, 0.001262813, 0.00123712, 
    0.001245872, 0.001403145, 0.00162145, 0.001952306, 0.002063203, 
    0.001781819, 0.001632783, 0.001708499, 0.002409449,
  0.001539334, 0.001518982, 0.001439188, 0.001339688, 0.001266435, 
    0.001251617, 0.001307539, 0.001280674, 0.001405679, 0.001924203, 
    0.002076892, 0.001742901, 0.001667241, 0.001789544, 0.002547764,
  0.001522279, 0.001460436, 0.001336548, 0.001300726, 0.00124962, 
    0.001192917, 0.001320469, 0.001440622, 0.001657228, 0.00189388, 
    0.002067877, 0.001875038, 0.001703861, 0.001768082, 0.002391333,
  0.001514845, 0.001408388, 0.001270613, 0.001238305, 0.001272904, 
    0.001155816, 0.001268135, 0.001455491, 0.001651444, 0.001862697, 
    0.002068417, 0.002176638, 0.00177064, 0.001743314, 0.002168298,
  0.001621736, 0.00143907, 0.001226724, 0.001135665, 0.001281627, 
    0.001139787, 0.001208672, 0.001367887, 0.001490148, 0.001711667, 
    0.00192962, 0.002223822, 0.002102086, 0.001771787, 0.001960519,
  0.001831956, 0.001643232, 0.001225927, 0.001060708, 0.001249847, 
    0.001167831, 0.00115615, 0.001334402, 0.001440742, 0.00163609, 
    0.001743845, 0.002167606, 0.002304062, 0.00195307, 0.001836708,
  0.002013956, 0.001812481, 0.001352715, 0.001098165, 0.001264888, 
    0.001161796, 0.001113571, 0.001299222, 0.001389716, 0.00150288, 
    0.001551488, 0.001868941, 0.002340611, 0.002298365, 0.001861758,
  0.001388551, 0.001505456, 0.001276594, 0.001291201, 0.001247565, 
    0.001217105, 0.001310702, 0.001539989, 0.001687688, 0.001824756, 
    0.002046461, 0.002094951, 0.002059091, 0.002028173, 0.002021491,
  0.001596097, 0.001471848, 0.001383978, 0.001309269, 0.001321911, 
    0.001174316, 0.001272956, 0.001566103, 0.001715528, 0.001962889, 
    0.002194639, 0.002150392, 0.002032161, 0.001755002, 0.00173863,
  0.00150469, 0.001578144, 0.001476404, 0.001295032, 0.001236967, 
    0.001159251, 0.001253647, 0.001435236, 0.001731603, 0.002027756, 
    0.002213765, 0.002221867, 0.00212472, 0.001938474, 0.001890858,
  0.001507211, 0.001557362, 0.001477515, 0.001268299, 0.00122821, 
    0.001128274, 0.00120426, 0.001318271, 0.001575727, 0.001934717, 
    0.002197785, 0.002367454, 0.002209906, 0.002210809, 0.002288174,
  0.001555467, 0.001453196, 0.001427962, 0.001258241, 0.0012242, 0.00120807, 
    0.001356148, 0.001251403, 0.001347575, 0.001865428, 0.002166291, 
    0.002421328, 0.002296819, 0.00233169, 0.002445943,
  0.00169005, 0.00143273, 0.001366832, 0.001274916, 0.001240156, 0.001215507, 
    0.001344181, 0.001482294, 0.001605364, 0.001866956, 0.002108982, 
    0.002429314, 0.002385304, 0.002392491, 0.002523474,
  0.001872012, 0.001511327, 0.001384919, 0.001291914, 0.001274547, 
    0.001233188, 0.001323784, 0.001392436, 0.001539914, 0.001787303, 
    0.0020108, 0.002386874, 0.002442475, 0.002428113, 0.002523311,
  0.002002601, 0.001647045, 0.001549969, 0.001233745, 0.001322917, 
    0.001240794, 0.001328988, 0.001358104, 0.001400416, 0.001604478, 
    0.001830293, 0.002286974, 0.002445864, 0.002440813, 0.002487547,
  0.002184042, 0.002035712, 0.001815891, 0.001270673, 0.001308924, 
    0.001243393, 0.001331362, 0.001332028, 0.001354833, 0.001499181, 
    0.00164946, 0.002106472, 0.002456869, 0.002457601, 0.002443557,
  0.002231391, 0.002170874, 0.00197717, 0.001343492, 0.001321885, 
    0.001233349, 0.001287897, 0.001325112, 0.001351401, 0.001403854, 
    0.001500691, 0.001857982, 0.002420267, 0.002487344, 0.002386904,
  0.001440078, 0.001404061, 0.00132272, 0.001260634, 0.001254234, 0.0012669, 
    0.001396281, 0.001473744, 0.001613952, 0.001790549, 0.001903077, 
    0.002172774, 0.002293942, 0.002268721, 0.002154613,
  0.001697205, 0.001548634, 0.001386146, 0.001249958, 0.001267781, 
    0.001282144, 0.001331414, 0.001351487, 0.001428477, 0.001680937, 
    0.001830138, 0.002077535, 0.002271851, 0.002251128, 0.002278413,
  0.001794402, 0.001552887, 0.001447256, 0.00125272, 0.001243006, 
    0.001193852, 0.001235941, 0.00123386, 0.001411545, 0.001568971, 
    0.001683352, 0.001991133, 0.002264789, 0.002396884, 0.002480916,
  0.001892911, 0.001501484, 0.001449506, 0.001259722, 0.001293118, 
    0.001273225, 0.001214721, 0.001169018, 0.00127399, 0.001449022, 0.001558, 
    0.001880322, 0.002242765, 0.002347331, 0.002425221,
  0.001909934, 0.001525729, 0.001511657, 0.001280192, 0.001308055, 
    0.001269035, 0.001332774, 0.001118805, 0.001134627, 0.001355854, 
    0.001479291, 0.001842478, 0.002253419, 0.002349209, 0.002455231,
  0.001887224, 0.001624256, 0.001572895, 0.001306962, 0.001333907, 
    0.001295337, 0.001310291, 0.001299758, 0.00129189, 0.001305247, 
    0.001435683, 0.001854372, 0.002299951, 0.00243024, 0.002547793,
  0.001829054, 0.001742486, 0.001771572, 0.001351198, 0.001308715, 
    0.001297232, 0.00130253, 0.001300444, 0.001288966, 0.001272883, 
    0.001460197, 0.001879651, 0.002309193, 0.00242779, 0.002384828,
  0.001878253, 0.00181284, 0.001871888, 0.001328798, 0.001287618, 
    0.001361217, 0.001316514, 0.001286053, 0.001285427, 0.001255677, 
    0.001451292, 0.00189804, 0.002278408, 0.002284669, 0.002328118,
  0.00202726, 0.002050986, 0.00202924, 0.001516111, 0.001418155, 0.001350267, 
    0.00133455, 0.001285236, 0.001268694, 0.001288836, 0.001420157, 
    0.001906476, 0.002193102, 0.002066734, 0.002079407,
  0.002125619, 0.002503971, 0.002385214, 0.00198944, 0.001784726, 
    0.001514317, 0.001335777, 0.001305886, 0.001270279, 0.001292226, 
    0.001377489, 0.001901194, 0.002093125, 0.002010829, 0.001936219,
  0.001311359, 0.001511692, 0.001458227, 0.001362395, 0.001336358, 
    0.001272215, 0.001288709, 0.001338776, 0.001264551, 0.001307256, 
    0.001261907, 0.001281035, 0.00147457, 0.001752198, 0.001861808,
  0.001525287, 0.001687084, 0.001611582, 0.001506172, 0.001449068, 
    0.00134374, 0.001293219, 0.001159259, 0.001130683, 0.001189915, 
    0.001233333, 0.001284029, 0.00145974, 0.001762803, 0.001782924,
  0.001702139, 0.001836882, 0.001829605, 0.001704393, 0.001566153, 
    0.001367825, 0.001280494, 0.001276766, 0.00119272, 0.001251529, 
    0.001166938, 0.001315132, 0.001562402, 0.00182436, 0.00188755,
  0.001879156, 0.00199826, 0.0020591, 0.001927633, 0.001900622, 0.001681905, 
    0.00135252, 0.001254537, 0.001219188, 0.001239058, 0.001261161, 
    0.001329522, 0.001571877, 0.001776458, 0.001906984,
  0.002103442, 0.002225493, 0.002384912, 0.002246974, 0.002175655, 
    0.002002321, 0.001713762, 0.001281398, 0.001110848, 0.001232014, 
    0.001251241, 0.001335897, 0.001565512, 0.001773419, 0.001841143,
  0.002293093, 0.002460646, 0.002631168, 0.002509723, 0.002307774, 
    0.002114308, 0.001951856, 0.001749182, 0.001487324, 0.001328981, 
    0.001298853, 0.001387539, 0.001620369, 0.001758499, 0.001828743,
  0.002498336, 0.002635718, 0.002724601, 0.002524015, 0.002224687, 
    0.002027552, 0.002040465, 0.001968179, 0.001739032, 0.001448232, 
    0.00136885, 0.001425295, 0.001683308, 0.001806112, 0.001814256,
  0.002600493, 0.002636755, 0.002660742, 0.002458276, 0.002124839, 
    0.001987939, 0.002037103, 0.002149695, 0.001861939, 0.001529641, 
    0.001367889, 0.001486962, 0.00171596, 0.001838392, 0.001862557,
  0.002581225, 0.002552029, 0.002511112, 0.002334769, 0.002147647, 
    0.001981076, 0.001955638, 0.001931446, 0.001591842, 0.001290013, 
    0.001326679, 0.00154049, 0.001817088, 0.001887657, 0.001942235,
  0.002543729, 0.002509487, 0.002312508, 0.002138451, 0.001979929, 
    0.001777528, 0.001660947, 0.00162785, 0.001370388, 0.001394057, 
    0.001391683, 0.001725423, 0.001962541, 0.001993269, 0.001890307,
  0.001906782, 0.001830231, 0.001864227, 0.001825281, 0.001853968, 
    0.001865446, 0.001810727, 0.001764514, 0.001741763, 0.001664461, 
    0.001522696, 0.001316569, 0.001217773, 0.001273726, 0.001507055,
  0.002470227, 0.002236012, 0.002274169, 0.002246827, 0.002221713, 
    0.002199733, 0.002090932, 0.001999959, 0.001852515, 0.001728073, 
    0.00159012, 0.001371225, 0.001124321, 0.00121067, 0.001311725,
  0.002550818, 0.002525014, 0.002485837, 0.002451391, 0.002498969, 
    0.002390408, 0.002490086, 0.002448282, 0.002278842, 0.002040741, 
    0.001723368, 0.001508642, 0.001181121, 0.001235579, 0.001304064,
  0.002543184, 0.002455402, 0.002355102, 0.002255727, 0.002208402, 
    0.002259207, 0.002158771, 0.002309873, 0.002315689, 0.002342709, 
    0.002132752, 0.001761269, 0.001300844, 0.001233181, 0.001256708,
  0.002404244, 0.002287747, 0.002097333, 0.001916755, 0.00183701, 
    0.001804136, 0.001835205, 0.001680505, 0.001635747, 0.002111934, 
    0.002208162, 0.001945984, 0.001398198, 0.001219218, 0.001165676,
  0.002211533, 0.002022807, 0.001806864, 0.001686313, 0.001641887, 
    0.001574242, 0.001566156, 0.001674359, 0.001682647, 0.001717551, 
    0.002005524, 0.001981422, 0.001568055, 0.001251668, 0.001207848,
  0.002044145, 0.001853331, 0.001681904, 0.001667564, 0.001673401, 
    0.001668886, 0.001635688, 0.001769842, 0.001850759, 0.001860693, 
    0.001943173, 0.001928721, 0.001606075, 0.001352899, 0.001358152,
  0.001989601, 0.001854166, 0.001696965, 0.00168173, 0.001719844, 
    0.001809451, 0.001838609, 0.001839659, 0.001848031, 0.002045308, 
    0.001977653, 0.001873197, 0.001622894, 0.001456255, 0.001369423,
  0.0020127, 0.001874682, 0.001680608, 0.001711951, 0.001804484, 0.001952731, 
    0.00203989, 0.001860971, 0.001699882, 0.001805551, 0.00199973, 
    0.001812335, 0.001614138, 0.001455109, 0.001461051,
  0.002031485, 0.001808722, 0.001707896, 0.001744129, 0.001855318, 
    0.002058005, 0.002190574, 0.002103554, 0.001763923, 0.001667017, 
    0.001870482, 0.001765646, 0.001592329, 0.0014772, 0.001516607,
  0.00200172, 0.001953771, 0.002029005, 0.001767777, 0.001626447, 
    0.001569257, 0.00166801, 0.00184507, 0.00172704, 0.00158777, 0.001632718, 
    0.001591914, 0.001370718, 0.001223088, 0.001308082,
  0.002237373, 0.002233316, 0.002124147, 0.002004982, 0.001938686, 
    0.001873392, 0.001861463, 0.001948738, 0.001933177, 0.001720536, 
    0.001686775, 0.001716178, 0.001519041, 0.001256585, 0.001249344,
  0.00249395, 0.002510954, 0.002467394, 0.002262686, 0.00208086, 0.001809851, 
    0.001650498, 0.001693147, 0.001919956, 0.002002852, 0.001830022, 
    0.001827996, 0.001643469, 0.00139585, 0.001295497,
  0.002576485, 0.002561276, 0.002532324, 0.002420996, 0.002253534, 
    0.002041241, 0.001546665, 0.00141987, 0.001381034, 0.001875237, 
    0.001996502, 0.002001997, 0.001825994, 0.001533563, 0.001322734,
  0.002618742, 0.002530977, 0.002380219, 0.002344699, 0.002099684, 
    0.002044635, 0.001855113, 0.001413723, 0.001158478, 0.001331658, 
    0.002030829, 0.002160708, 0.001930147, 0.001662611, 0.001179442,
  0.002561791, 0.002356553, 0.002160701, 0.00188873, 0.001792006, 
    0.001787652, 0.001947663, 0.001840536, 0.001488342, 0.001346414, 
    0.001920773, 0.002274311, 0.002061842, 0.001543, 0.001366846,
  0.002395535, 0.002200241, 0.001908767, 0.001806692, 0.001813824, 
    0.001975658, 0.002109727, 0.002149805, 0.001909147, 0.001458367, 
    0.001723835, 0.00228295, 0.002047526, 0.001544554, 0.001597816,
  0.002284847, 0.002074895, 0.001840017, 0.001883482, 0.002047171, 
    0.002165333, 0.002147694, 0.00211743, 0.001960456, 0.001732269, 
    0.001704475, 0.002269149, 0.0019473, 0.001542883, 0.001551463,
  0.002186301, 0.002025059, 0.001935925, 0.001992344, 0.002137063, 
    0.002115067, 0.002242164, 0.002164955, 0.001975255, 0.001697372, 
    0.00176974, 0.002200078, 0.001770945, 0.001545463, 0.001493711,
  0.002126352, 0.001963023, 0.002002775, 0.002116185, 0.002233787, 
    0.002306802, 0.002250907, 0.002147868, 0.001765297, 0.001695851, 
    0.001965204, 0.002092794, 0.001618871, 0.001515768, 0.001480387,
  0.002731265, 0.002619199, 0.00263968, 0.002519478, 0.002236102, 0.00195299, 
    0.001874754, 0.001849145, 0.001893126, 0.00202457, 0.001927974, 
    0.001666776, 0.001539113, 0.001456468, 0.001644586,
  0.002960655, 0.00272424, 0.002610682, 0.002662415, 0.002593947, 
    0.002490932, 0.002214093, 0.001901004, 0.001886526, 0.00208364, 
    0.002048323, 0.001818138, 0.001510742, 0.001267347, 0.001452964,
  0.003198608, 0.003175918, 0.003037738, 0.002987043, 0.002917289, 
    0.002624895, 0.002518019, 0.00225779, 0.001911123, 0.002103854, 
    0.002028234, 0.001878573, 0.001642326, 0.001347431, 0.001410164,
  0.002946944, 0.002825385, 0.002719252, 0.00272666, 0.002665004, 0.00278169, 
    0.002454627, 0.002354852, 0.001893426, 0.001930105, 0.001973178, 
    0.001850693, 0.001662808, 0.00138484, 0.001279752,
  0.002617569, 0.002386675, 0.002201091, 0.002305317, 0.001915307, 
    0.002107133, 0.002107263, 0.002053159, 0.001642778, 0.001794343, 
    0.001996579, 0.001837902, 0.001653077, 0.00143253, 0.001312066,
  0.002319793, 0.002195982, 0.002099389, 0.002054803, 0.001840425, 
    0.001515008, 0.002044375, 0.002101025, 0.001778027, 0.001713395, 
    0.001830231, 0.001825617, 0.001701485, 0.001427539, 0.00134647,
  0.002157904, 0.002089851, 0.001952455, 0.002117065, 0.001922829, 
    0.001631423, 0.001943081, 0.002041942, 0.001814238, 0.001739082, 
    0.001830707, 0.0018107, 0.001676798, 0.001491188, 0.001694851,
  0.002028905, 0.001978681, 0.001971716, 0.002020248, 0.002012055, 
    0.00194497, 0.001873905, 0.002039815, 0.001792559, 0.001751006, 
    0.001808643, 0.001819496, 0.001677641, 0.00161861, 0.001677964,
  0.00195167, 0.001961101, 0.001946871, 0.001892772, 0.002080162, 
    0.001929267, 0.002037975, 0.001975434, 0.001852239, 0.001742325, 
    0.001807627, 0.001842809, 0.001647659, 0.001604913, 0.001611027,
  0.00191601, 0.001951924, 0.001999406, 0.00198842, 0.001963122, 0.001998028, 
    0.001992024, 0.001959434, 0.001821324, 0.001747878, 0.001881635, 
    0.001848942, 0.001635688, 0.001574872, 0.001605632,
  0.002824596, 0.002573733, 0.002592213, 0.002692037, 0.002734389, 
    0.002520383, 0.002259867, 0.002266794, 0.00218491, 0.002190778, 
    0.001882776, 0.001689413, 0.00200946, 0.002151057, 0.002507075,
  0.003199606, 0.002936634, 0.002756564, 0.002942208, 0.002861652, 
    0.002558805, 0.002414187, 0.002236443, 0.001975478, 0.00187499, 
    0.002048989, 0.001773953, 0.001938576, 0.002001511, 0.002398997,
  0.003441923, 0.003343159, 0.003145196, 0.002723549, 0.002625641, 
    0.002444801, 0.002471843, 0.002277846, 0.002046126, 0.002051213, 
    0.002029652, 0.001759975, 0.001947656, 0.00198182, 0.002221292,
  0.002610645, 0.002536662, 0.002436037, 0.002446767, 0.00243902, 
    0.002585121, 0.002511439, 0.00247233, 0.002091985, 0.002147483, 
    0.001972159, 0.001719445, 0.00180455, 0.001891874, 0.002044271,
  0.002351731, 0.002292547, 0.002247797, 0.002473661, 0.002399371, 
    0.002445709, 0.002693755, 0.002238276, 0.001999887, 0.002083178, 
    0.001908812, 0.001780669, 0.001791784, 0.001859206, 0.002003899,
  0.002046726, 0.001985728, 0.001976926, 0.002180671, 0.002174712, 
    0.00183328, 0.002291204, 0.002545824, 0.002166771, 0.00209962, 
    0.001930225, 0.001727331, 0.00176472, 0.001803013, 0.002003407,
  0.001920014, 0.001820943, 0.001740584, 0.001892946, 0.002086407, 
    0.00183547, 0.00178869, 0.002454577, 0.002281629, 0.002067549, 
    0.001903546, 0.001711991, 0.001707649, 0.001881421, 0.001961573,
  0.001823191, 0.001740749, 0.001642041, 0.001795958, 0.002035643, 
    0.001828307, 0.001761536, 0.002321171, 0.002210373, 0.001957784, 
    0.001808365, 0.001665178, 0.001736474, 0.001848949, 0.001890999,
  0.001829254, 0.001859679, 0.001954539, 0.001948118, 0.001984794, 
    0.001853217, 0.002106452, 0.002318311, 0.002187463, 0.001864065, 
    0.001697455, 0.001633953, 0.001699718, 0.001756869, 0.001755886,
  0.0018634, 0.001913692, 0.00201083, 0.00201487, 0.002019849, 0.002095333, 
    0.002229255, 0.002247765, 0.002009658, 0.001758338, 0.001578032, 
    0.001581961, 0.001652751, 0.001621688, 0.001636288,
  0.002734944, 0.002676569, 0.002596698, 0.002664851, 0.002596716, 
    0.00242672, 0.002423208, 0.002638163, 0.002704879, 0.002600323, 
    0.002204874, 0.002097062, 0.002040705, 0.002049474, 0.002427476,
  0.003204499, 0.003033279, 0.002763306, 0.002761211, 0.002848053, 
    0.002602069, 0.002586406, 0.002654612, 0.002547096, 0.002381089, 
    0.002174214, 0.002051754, 0.002043383, 0.002191209, 0.002630858,
  0.003504223, 0.003432278, 0.003231781, 0.002699608, 0.002846774, 
    0.002297511, 0.002281255, 0.002369333, 0.002331894, 0.002227363, 
    0.001920792, 0.001919304, 0.002035157, 0.002383599, 0.002859922,
  0.002526416, 0.00254034, 0.002560595, 0.002528345, 0.002278156, 
    0.002301725, 0.002295151, 0.002161909, 0.00224657, 0.001979527, 
    0.001743094, 0.001795896, 0.002215204, 0.00260838, 0.002941728,
  0.002311178, 0.002279616, 0.002205046, 0.002421451, 0.00218344, 
    0.002299107, 0.002477921, 0.001890256, 0.001664512, 0.002033034, 
    0.0018176, 0.00209548, 0.002455124, 0.002789532, 0.002835104,
  0.002096906, 0.001969527, 0.0019408, 0.002130298, 0.002099616, 0.002099564, 
    0.002310376, 0.00207697, 0.001923933, 0.001880943, 0.001938638, 
    0.002358107, 0.002685306, 0.002781934, 0.002691064,
  0.001948626, 0.001812294, 0.001730975, 0.001905898, 0.002002438, 
    0.002043153, 0.002466943, 0.002230457, 0.002043319, 0.002079967, 
    0.002304673, 0.002584951, 0.002683759, 0.00268583, 0.002586325,
  0.001826928, 0.001719858, 0.001598315, 0.0017712, 0.002019831, 0.002132558, 
    0.002406639, 0.002317656, 0.002065063, 0.002195147, 0.002353643, 
    0.002508462, 0.002531963, 0.002454016, 0.002382868,
  0.001769534, 0.001841331, 0.00192443, 0.001909037, 0.002004003, 
    0.002179477, 0.002392738, 0.002226323, 0.002050382, 0.002107662, 
    0.002217878, 0.002355136, 0.002332712, 0.002291068, 0.002237295,
  0.001806281, 0.00189857, 0.00200195, 0.00201909, 0.002199989, 0.002293164, 
    0.002284325, 0.00208571, 0.001955686, 0.001967445, 0.002048206, 
    0.002114446, 0.002144661, 0.002136238, 0.002143058,
  0.003391913, 0.003078708, 0.002851414, 0.002973518, 0.002713574, 
    0.002793904, 0.002875512, 0.002813631, 0.002607765, 0.002508506, 
    0.002440069, 0.002498238, 0.002491093, 0.00233314, 0.002199048,
  0.003254837, 0.002871041, 0.002800258, 0.00278551, 0.00293335, 0.002925461, 
    0.002913898, 0.00281304, 0.002640944, 0.002614526, 0.002482193, 
    0.002566846, 0.002550289, 0.002263231, 0.002165418,
  0.003332175, 0.003168056, 0.003175384, 0.002829632, 0.002795817, 
    0.002171393, 0.00221543, 0.002330012, 0.002378163, 0.002346016, 
    0.00232464, 0.002469276, 0.002385431, 0.002179815, 0.002065124,
  0.002678859, 0.0025674, 0.00262425, 0.00278924, 0.002198262, 0.00217991, 
    0.001940771, 0.00193085, 0.002115678, 0.002310389, 0.002289619, 
    0.002322193, 0.002192558, 0.002157916, 0.002268657,
  0.002474341, 0.002504354, 0.002360073, 0.002253168, 0.001842857, 
    0.001903843, 0.001974195, 0.001725778, 0.001586954, 0.001836259, 
    0.002135439, 0.002137106, 0.002117351, 0.002162529, 0.002445225,
  0.002437293, 0.002178502, 0.002020857, 0.001985265, 0.001779541, 
    0.001866331, 0.001947757, 0.001875028, 0.002005376, 0.001845015, 
    0.001909974, 0.002120088, 0.00223856, 0.002499665, 0.002472577,
  0.002090647, 0.001977775, 0.001675646, 0.001896504, 0.001903741, 
    0.001984758, 0.002083124, 0.001972543, 0.002132751, 0.002194581, 
    0.002311186, 0.002438062, 0.002546408, 0.002511389, 0.002398413,
  0.001922684, 0.001837944, 0.001723551, 0.001956762, 0.0020645, 0.002232926, 
    0.002142491, 0.00207448, 0.00215654, 0.002394115, 0.002545159, 
    0.002590794, 0.002514793, 0.002323573, 0.002214138,
  0.001837051, 0.001915672, 0.001953477, 0.002033751, 0.002123364, 
    0.002181084, 0.002186187, 0.002231851, 0.002372328, 0.002615398, 
    0.002626361, 0.002504725, 0.002357894, 0.00225863, 0.002295586,
  0.001874138, 0.001962027, 0.002091979, 0.002137359, 0.002175625, 
    0.002231944, 0.002264365, 0.002425315, 0.002594329, 0.002543672, 
    0.002432246, 0.002340466, 0.002284741, 0.00234398, 0.002435311,
  0.003531136, 0.00321705, 0.002984217, 0.002831341, 0.002750177, 
    0.002730081, 0.002613311, 0.002532524, 0.002407073, 0.002394612, 
    0.002480321, 0.002156527, 0.002218322, 0.002181174, 0.002158443,
  0.003360159, 0.003104165, 0.002977428, 0.00283891, 0.002771107, 
    0.002787609, 0.002598628, 0.002481026, 0.002362166, 0.002408199, 
    0.002516364, 0.002394935, 0.002227834, 0.002196421, 0.001966532,
  0.003553107, 0.003385102, 0.003206841, 0.003007474, 0.00278242, 
    0.002285813, 0.002143886, 0.002020833, 0.002059803, 0.002159778, 
    0.002282287, 0.002493079, 0.002429808, 0.002138785, 0.002095814,
  0.003550994, 0.00317796, 0.003068236, 0.002906023, 0.0025497, 0.002181162, 
    0.001662799, 0.001637521, 0.001664653, 0.00178161, 0.002109147, 
    0.002427822, 0.002527791, 0.002402748, 0.002245904,
  0.00335608, 0.003198749, 0.00301792, 0.002616455, 0.002098302, 0.001961374, 
    0.001830122, 0.001664311, 0.001333841, 0.001652872, 0.001940208, 
    0.002248809, 0.002506145, 0.002306556, 0.002161145,
  0.003063365, 0.002721605, 0.0024776, 0.002286443, 0.00198719, 0.002007678, 
    0.002042573, 0.001966382, 0.001834775, 0.001649729, 0.001788494, 
    0.001939687, 0.002203152, 0.002276729, 0.002267129,
  0.00251198, 0.002247629, 0.002165582, 0.002006088, 0.001952784, 
    0.002063211, 0.002083174, 0.002031934, 0.00210335, 0.001886, 0.00193038, 
    0.002125052, 0.002260752, 0.002180371, 0.002157247,
  0.002116586, 0.001947662, 0.001997052, 0.001977195, 0.002086469, 
    0.002110714, 0.001993877, 0.002037999, 0.001881658, 0.0017839, 
    0.00192912, 0.002085232, 0.002123077, 0.002074165, 0.002084632,
  0.001886245, 0.001963888, 0.002051824, 0.002098551, 0.002221064, 
    0.001984169, 0.001990326, 0.001963626, 0.002050078, 0.001989295, 
    0.001836957, 0.002067347, 0.002088835, 0.00204747, 0.002061815,
  0.001918517, 0.002051726, 0.002057036, 0.002246133, 0.002160162, 
    0.002384724, 0.002247503, 0.002289043, 0.002216695, 0.002085817, 
    0.002010845, 0.002072966, 0.002067962, 0.002051473, 0.002100481,
  0.004959674, 0.004561756, 0.004189422, 0.004137703, 0.004001113, 
    0.003866927, 0.003680406, 0.003508057, 0.003311618, 0.003124717, 
    0.002957867, 0.002721703, 0.002585319, 0.002464193, 0.002292778,
  0.004237161, 0.004242615, 0.004126579, 0.00405054, 0.004093833, 
    0.003778156, 0.003614246, 0.003414956, 0.003186044, 0.002910224, 
    0.002728421, 0.002462743, 0.002416602, 0.002259146, 0.002062888,
  0.004337595, 0.004214833, 0.004119747, 0.004017307, 0.003793592, 
    0.003493165, 0.003140354, 0.002962394, 0.002782914, 0.002538878, 
    0.002375202, 0.002242532, 0.002309451, 0.00221965, 0.002219553,
  0.004433058, 0.004305761, 0.004050106, 0.003764012, 0.003527277, 
    0.003134392, 0.002476783, 0.002490696, 0.002390817, 0.00224439, 
    0.002192059, 0.002059411, 0.002052349, 0.002250432, 0.002200806,
  0.004334421, 0.003946872, 0.003673169, 0.003257334, 0.002891787, 
    0.002546321, 0.002234375, 0.001970866, 0.001769884, 0.002033701, 
    0.001840028, 0.00179151, 0.001894787, 0.002179377, 0.002258763,
  0.003533775, 0.003359257, 0.003072273, 0.002752913, 0.002418095, 
    0.002213818, 0.002049811, 0.002019951, 0.001990389, 0.001909556, 
    0.001789449, 0.001875394, 0.002012091, 0.002199575, 0.00229976,
  0.003082713, 0.002918495, 0.002754851, 0.002329799, 0.0021746, 0.002101423, 
    0.002006616, 0.001969388, 0.001926296, 0.001860251, 0.001696602, 
    0.001800261, 0.002198636, 0.002299677, 0.002319966,
  0.002660815, 0.002557287, 0.002472941, 0.002170375, 0.002073016, 
    0.002170706, 0.001989474, 0.001949895, 0.001861398, 0.001881193, 
    0.001828525, 0.00205768, 0.0022797, 0.002340186, 0.002196321,
  0.002420616, 0.002308698, 0.002328857, 0.002152261, 0.002246598, 
    0.002064756, 0.00196754, 0.001893784, 0.001817596, 0.001789706, 
    0.001911324, 0.002001267, 0.002080275, 0.001970814, 0.001833236,
  0.002284222, 0.002225419, 0.002261413, 0.002304624, 0.002110266, 
    0.002056317, 0.001963242, 0.001883958, 0.001791237, 0.00179798, 
    0.001834584, 0.001825008, 0.00186587, 0.001889344, 0.001791963,
  0.002871404, 0.003009218, 0.003090433, 0.003195695, 0.003332098, 
    0.003444728, 0.003515763, 0.003617904, 0.003697127, 0.003737071, 
    0.003788857, 0.003794538, 0.003834636, 0.003718592, 0.00360619,
  0.00308782, 0.002999297, 0.003050629, 0.003257009, 0.003457591, 
    0.003547277, 0.003631682, 0.00369851, 0.00374244, 0.003788386, 
    0.003825273, 0.003834197, 0.003769991, 0.003595484, 0.003449925,
  0.002912948, 0.002911244, 0.00309582, 0.003355165, 0.003550736, 
    0.003594583, 0.003602111, 0.00322915, 0.003286134, 0.003388281, 
    0.00347593, 0.00354103, 0.003513319, 0.00341593, 0.003268068,
  0.002764647, 0.002927485, 0.003128518, 0.003285419, 0.003378775, 
    0.003302019, 0.002635228, 0.002609214, 0.002673659, 0.002902573, 
    0.002978899, 0.003106391, 0.003187902, 0.003112479, 0.002937182,
  0.002662622, 0.002784583, 0.002840529, 0.002755682, 0.002656622, 
    0.002576087, 0.002343288, 0.00213813, 0.002084834, 0.002573227, 
    0.002685253, 0.002748575, 0.002810586, 0.002775377, 0.002643337,
  0.00246574, 0.002451628, 0.0024006, 0.002279837, 0.002180122, 0.002133803, 
    0.002128458, 0.002221185, 0.002296062, 0.002362117, 0.002437869, 
    0.002473982, 0.002491581, 0.002477647, 0.00241156,
  0.00228001, 0.00228056, 0.002107463, 0.00202306, 0.001984037, 0.00195409, 
    0.001930489, 0.001957913, 0.002041458, 0.002185332, 0.002247502, 
    0.002252835, 0.00227235, 0.002267234, 0.002230168,
  0.002188874, 0.002122457, 0.001945798, 0.001944703, 0.001920967, 0.0019863, 
    0.001975819, 0.001975637, 0.001966314, 0.001997265, 0.002151529, 
    0.002156111, 0.002181153, 0.002160901, 0.002044022,
  0.002097467, 0.002008321, 0.001796096, 0.001774511, 0.001771384, 
    0.001827012, 0.001905724, 0.001993373, 0.002046649, 0.002113397, 
    0.002142394, 0.002196164, 0.002133088, 0.002079467, 0.00199634,
  0.002014015, 0.001896868, 0.001793839, 0.001752328, 0.001723169, 
    0.001721659, 0.001765844, 0.001886143, 0.001937422, 0.002063683, 
    0.002133004, 0.002170175, 0.002046812, 0.002064807, 0.002240119,
  0.003036485, 0.002960595, 0.002712046, 0.002496848, 0.002596266, 
    0.002620983, 0.00255431, 0.002288973, 0.00225708, 0.002417391, 
    0.002624766, 0.002790074, 0.002955321, 0.003088265, 0.003267163,
  0.003236259, 0.002882221, 0.002590109, 0.002446299, 0.002524889, 
    0.002384384, 0.002314241, 0.002133378, 0.002094308, 0.002228135, 
    0.00247005, 0.002738438, 0.002959603, 0.00312862, 0.003358426,
  0.00321478, 0.002833379, 0.00252995, 0.002381035, 0.002360302, 0.002130867, 
    0.002139947, 0.001995057, 0.001950353, 0.002065517, 0.002227075, 
    0.002567488, 0.002913305, 0.003271034, 0.003488355,
  0.003232092, 0.002788051, 0.002456238, 0.002385881, 0.002212103, 
    0.002140306, 0.001871932, 0.001834277, 0.001868541, 0.002013305, 
    0.002111823, 0.002433856, 0.002904205, 0.003367217, 0.003574556,
  0.002936405, 0.00248336, 0.002305601, 0.002280927, 0.002071444, 
    0.001961399, 0.001996963, 0.001830009, 0.001762119, 0.001982777, 
    0.002022027, 0.002321729, 0.002859123, 0.003384472, 0.003613438,
  0.002505494, 0.002197164, 0.002048425, 0.002121851, 0.001935948, 
    0.001907858, 0.002075926, 0.002191115, 0.002198694, 0.002089853, 
    0.001952639, 0.002298989, 0.002760999, 0.003120102, 0.003407759,
  0.002242049, 0.002027906, 0.001795915, 0.001826082, 0.001791091, 
    0.001826857, 0.001838898, 0.002094347, 0.002117237, 0.002084207, 
    0.001934915, 0.002318327, 0.002731356, 0.002907516, 0.003032737,
  0.002135522, 0.001941503, 0.001647382, 0.001565415, 0.001602057, 
    0.001674689, 0.001756949, 0.00194282, 0.002041024, 0.001906729, 
    0.001917337, 0.002363391, 0.002728704, 0.002764583, 0.002736981,
  0.002167732, 0.001820542, 0.001523432, 0.001562913, 0.001624264, 
    0.001691911, 0.001773907, 0.001910418, 0.001927584, 0.001872828, 
    0.001905477, 0.00237626, 0.00270361, 0.002766082, 0.002663642,
  0.00209949, 0.001694227, 0.001560377, 0.001682605, 0.001787669, 
    0.001755042, 0.001756955, 0.001868758, 0.001807456, 0.001773068, 
    0.00196746, 0.002460742, 0.002651273, 0.00278475, 0.002697166,
  0.002573714, 0.00284328, 0.003044419, 0.003178172, 0.00329392, 0.003357753, 
    0.003310783, 0.003101841, 0.002825846, 0.002613286, 0.002343944, 
    0.002158509, 0.002037704, 0.001875845, 0.001874504,
  0.002836562, 0.002865471, 0.003032455, 0.003197944, 0.003354081, 
    0.003352409, 0.003270859, 0.002934209, 0.002639829, 0.002365935, 
    0.002229192, 0.002105698, 0.0018637, 0.001796615, 0.00191041,
  0.002812607, 0.002856326, 0.002989712, 0.003106394, 0.003230453, 
    0.003024355, 0.002908268, 0.002595616, 0.002378886, 0.002186799, 
    0.002101387, 0.002008836, 0.001823678, 0.001907076, 0.002312079,
  0.002739505, 0.002712792, 0.002826351, 0.002874346, 0.002854664, 
    0.002635809, 0.002296978, 0.002336806, 0.002176974, 0.002065359, 
    0.001941077, 0.00181975, 0.00185153, 0.002305985, 0.002839345,
  0.002534883, 0.002404668, 0.002466304, 0.002401675, 0.002450099, 
    0.002380461, 0.002203726, 0.001807877, 0.001693291, 0.001907015, 
    0.001789239, 0.001758428, 0.002147626, 0.002803797, 0.003399314,
  0.002420977, 0.002165508, 0.002091216, 0.002021186, 0.002082887, 
    0.002121782, 0.002101845, 0.002005251, 0.001898291, 0.001852338, 
    0.001841392, 0.002056704, 0.002575017, 0.003225514, 0.003623799,
  0.002320967, 0.001949372, 0.001794892, 0.001808851, 0.00177855, 
    0.001763941, 0.001805944, 0.001809184, 0.001755951, 0.001810857, 
    0.001873021, 0.002425211, 0.002817526, 0.003344471, 0.003621182,
  0.002235171, 0.001861281, 0.001613803, 0.001645465, 0.001613996, 
    0.001594708, 0.001655069, 0.001735177, 0.001794049, 0.001816614, 
    0.002150044, 0.00265568, 0.002889959, 0.003079507, 0.003232169,
  0.002290579, 0.001949125, 0.001708159, 0.001730622, 0.001745449, 
    0.001772116, 0.001744097, 0.001721105, 0.001810631, 0.001989743, 
    0.002442425, 0.002900854, 0.002877439, 0.002907173, 0.002880882,
  0.002360272, 0.00214057, 0.002051874, 0.002088235, 0.002063059, 
    0.001723967, 0.001780219, 0.001865612, 0.001789729, 0.002072513, 
    0.002658308, 0.002786209, 0.002667798, 0.002578195, 0.002496309,
  0.002418474, 0.002757654, 0.002750803, 0.002235527, 0.002049491, 
    0.002140473, 0.002310459, 0.002623141, 0.002933291, 0.003144855, 
    0.00321737, 0.002943604, 0.002757254, 0.002550314, 0.002466793,
  0.003080705, 0.002978142, 0.002645446, 0.00203655, 0.001942358, 
    0.002022705, 0.002150564, 0.002420021, 0.002707676, 0.002838474, 
    0.002781389, 0.002645891, 0.002469671, 0.002290667, 0.002194968,
  0.003361106, 0.003079877, 0.002504826, 0.001926088, 0.001834176, 
    0.001947145, 0.001986661, 0.002159609, 0.002349169, 0.002486279, 
    0.002431355, 0.002345336, 0.002219306, 0.00215918, 0.00221612,
  0.003657049, 0.003192865, 0.002416593, 0.001834276, 0.001778582, 
    0.001977774, 0.001885387, 0.001953651, 0.002105386, 0.002361627, 
    0.002420821, 0.002350674, 0.002262287, 0.002275012, 0.002460032,
  0.003821093, 0.003131284, 0.002374048, 0.001762521, 0.001751461, 
    0.001885568, 0.001952163, 0.001751638, 0.001800817, 0.002375476, 
    0.002500708, 0.002603076, 0.002744845, 0.003007339, 0.003346464,
  0.003646143, 0.003158202, 0.002442162, 0.001949837, 0.00181507, 
    0.001802343, 0.001877745, 0.001971564, 0.002069298, 0.00239092, 
    0.002557351, 0.002750125, 0.003096333, 0.003473622, 0.003522421,
  0.003090973, 0.002944192, 0.002694549, 0.002313792, 0.002012052, 
    0.001863096, 0.001807908, 0.001914411, 0.002039065, 0.002442828, 
    0.002703075, 0.002868321, 0.00326316, 0.003552625, 0.003593133,
  0.003007893, 0.002940309, 0.002903856, 0.00263641, 0.002335757, 
    0.001980274, 0.001823903, 0.00192589, 0.002023546, 0.002339556, 
    0.002677063, 0.002881281, 0.003236926, 0.003509584, 0.003474351,
  0.002703535, 0.002703639, 0.00283423, 0.002780547, 0.002589434, 
    0.002152262, 0.001899893, 0.002034523, 0.002058484, 0.002330167, 
    0.002656244, 0.002821025, 0.003009475, 0.003103015, 0.003070511,
  0.002554796, 0.002575903, 0.002547175, 0.00258774, 0.002670499, 0.00233974, 
    0.002075366, 0.002036885, 0.002035749, 0.002340244, 0.002556516, 
    0.002499107, 0.002538446, 0.002674597, 0.002661488,
  0.002710751, 0.002951732, 0.003104002, 0.002889334, 0.002125857, 
    0.001695266, 0.001580208, 0.001885345, 0.002300781, 0.002803326, 
    0.003083937, 0.003109811, 0.003032975, 0.002937348, 0.002943339,
  0.003253463, 0.003268241, 0.003180719, 0.002629034, 0.002033367, 
    0.001657507, 0.00155013, 0.001842325, 0.002157208, 0.002874146, 
    0.003180349, 0.003208359, 0.003104038, 0.002968894, 0.003044778,
  0.003570339, 0.003360891, 0.002972529, 0.002367876, 0.001858263, 
    0.001656684, 0.001621183, 0.001766025, 0.002097559, 0.00277953, 
    0.003129342, 0.003330385, 0.003252276, 0.003214041, 0.003203623,
  0.003941755, 0.003504055, 0.002898637, 0.002275631, 0.001674337, 
    0.00168706, 0.001686209, 0.001730392, 0.001944963, 0.002532874, 
    0.003006456, 0.003356806, 0.003351429, 0.003287336, 0.003224224,
  0.003779327, 0.003562752, 0.003133258, 0.002353411, 0.001907647, 
    0.001866546, 0.001882688, 0.001720623, 0.0017521, 0.002376553, 
    0.002883156, 0.003292551, 0.003299107, 0.003178626, 0.00308579,
  0.003124209, 0.003199336, 0.003373412, 0.002887908, 0.002432037, 
    0.002148918, 0.002068734, 0.002088851, 0.002015017, 0.00238474, 
    0.002821827, 0.003186997, 0.003188532, 0.003002964, 0.00291268,
  0.002688199, 0.002604238, 0.003074434, 0.003054723, 0.002930712, 
    0.00276664, 0.002600995, 0.002246226, 0.001972966, 0.002338246, 
    0.002759867, 0.003029335, 0.003037256, 0.002880418, 0.002814291,
  0.002780729, 0.002772294, 0.002673182, 0.002715526, 0.002736546, 
    0.003059311, 0.0028724, 0.002119358, 0.001990968, 0.002265603, 
    0.002657857, 0.002851111, 0.002861559, 0.002784917, 0.002804552,
  0.002494816, 0.00227766, 0.002418784, 0.002559683, 0.002678508, 0.00297775, 
    0.002576107, 0.002093187, 0.001998374, 0.002172098, 0.002643651, 
    0.002737991, 0.002757816, 0.002769265, 0.00286738,
  0.00239171, 0.002197917, 0.002373899, 0.002556996, 0.002608607, 
    0.002673414, 0.002284388, 0.002001127, 0.001976922, 0.002175828, 
    0.002589823, 0.002659172, 0.002750507, 0.002824224, 0.002918272,
  0.003265034, 0.002980269, 0.002780332, 0.002376633, 0.002042274, 
    0.00185576, 0.001690286, 0.00166534, 0.00194005, 0.002469371, 
    0.002816829, 0.002988331, 0.00296519, 0.00287344, 0.002909556,
  0.003112296, 0.002873871, 0.002583227, 0.002273401, 0.002058994, 
    0.001848033, 0.001720753, 0.001717787, 0.001782079, 0.002372779, 
    0.002758482, 0.002941702, 0.002966673, 0.002768767, 0.002767349,
  0.003069937, 0.002822377, 0.002583559, 0.002327859, 0.002089329, 
    0.001909353, 0.001892041, 0.001971241, 0.001844812, 0.002325921, 
    0.00273264, 0.002936862, 0.003004249, 0.002892104, 0.002854384,
  0.003051797, 0.0027369, 0.002512722, 0.002338189, 0.002021871, 0.002092227, 
    0.002034748, 0.001991373, 0.001949682, 0.002321465, 0.002730877, 
    0.002948167, 0.003065316, 0.003030465, 0.002959403,
  0.002891892, 0.002565102, 0.002456974, 0.002587033, 0.002146845, 
    0.002252596, 0.002338309, 0.001952935, 0.001860259, 0.002298156, 
    0.002740274, 0.00294346, 0.003125679, 0.003175161, 0.003163982,
  0.002851636, 0.002790059, 0.002731506, 0.00284178, 0.00280624, 0.002545942, 
    0.002388739, 0.002328486, 0.002306153, 0.002469436, 0.002759886, 
    0.002971173, 0.003187539, 0.003311363, 0.00337779,
  0.002676947, 0.002541467, 0.002447708, 0.002486606, 0.002532179, 
    0.002520903, 0.002439327, 0.002277919, 0.002335442, 0.002521435, 
    0.002693038, 0.002939893, 0.003230914, 0.003388482, 0.003454695,
  0.002615896, 0.002452395, 0.00229231, 0.002336269, 0.002263836, 
    0.002300979, 0.00227474, 0.002392534, 0.00246663, 0.002468599, 
    0.002707275, 0.003024542, 0.003292036, 0.003389986, 0.003426751,
  0.002530542, 0.002384949, 0.002293798, 0.00226228, 0.002216947, 
    0.002167653, 0.002254795, 0.002383888, 0.002503956, 0.002493916, 
    0.002708562, 0.003092132, 0.003347592, 0.003364993, 0.003369103,
  0.002487239, 0.002289496, 0.002170341, 0.002113475, 0.002103643, 
    0.002147322, 0.002249257, 0.002353961, 0.002407038, 0.002499379, 
    0.002719104, 0.003153334, 0.003385012, 0.003413421, 0.003369755,
  0.002207838, 0.002449317, 0.002341141, 0.002248066, 0.002181201, 
    0.002024016, 0.001978991, 0.002070284, 0.002298067, 0.002508626, 
    0.002763843, 0.002998057, 0.003151234, 0.003039989, 0.003076684,
  0.002515745, 0.002513797, 0.002376181, 0.00230853, 0.00220692, 0.002132029, 
    0.002091375, 0.002207581, 0.002290531, 0.002528305, 0.002798982, 
    0.003089727, 0.003149147, 0.002998833, 0.003064496,
  0.00262854, 0.002543915, 0.002362828, 0.002211583, 0.002112074, 
    0.002048803, 0.002137614, 0.002312502, 0.00241608, 0.002528176, 
    0.002774062, 0.003058744, 0.003114375, 0.003187139, 0.003201746,
  0.002700802, 0.002638995, 0.002368008, 0.002174154, 0.002083241, 
    0.002124572, 0.002134447, 0.002200717, 0.002380768, 0.002473041, 
    0.002731812, 0.003024821, 0.0030786, 0.003164216, 0.003215525,
  0.002709616, 0.002415138, 0.002201826, 0.00219722, 0.002116809, 
    0.002146652, 0.002243345, 0.002099082, 0.002105422, 0.002430572, 
    0.00277636, 0.002969438, 0.003108478, 0.003199837, 0.003259045,
  0.002612262, 0.002292328, 0.002103707, 0.002079365, 0.002092649, 
    0.002220256, 0.00229593, 0.00238302, 0.002502695, 0.002632244, 
    0.002838423, 0.002977364, 0.003158116, 0.003259907, 0.00334271,
  0.002589083, 0.002215137, 0.002011084, 0.002030775, 0.002096066, 
    0.002240649, 0.002287489, 0.00233144, 0.0025481, 0.002698909, 
    0.002811162, 0.003069288, 0.003253155, 0.003316981, 0.003404229,
  0.002485674, 0.002079157, 0.00197617, 0.002045644, 0.002145236, 0.00224253, 
    0.002223239, 0.002254459, 0.002531571, 0.002668697, 0.002815099, 
    0.003128214, 0.003284708, 0.003343535, 0.003391952,
  0.002325961, 0.001974074, 0.001995035, 0.002051635, 0.002200408, 
    0.002218626, 0.002136875, 0.002190439, 0.002465502, 0.00260693, 
    0.002808558, 0.003140115, 0.003307843, 0.003363174, 0.003372821,
  0.002185455, 0.001971949, 0.002033713, 0.002057929, 0.002204464, 
    0.002160463, 0.002058756, 0.002104485, 0.002381139, 0.002524486, 
    0.002815001, 0.003107992, 0.003298836, 0.003413716, 0.003412788,
  0.002306184, 0.002450043, 0.00222531, 0.00214091, 0.002132559, 0.002177465, 
    0.002159858, 0.002322519, 0.002423563, 0.002567429, 0.002635158, 
    0.00273052, 0.002879266, 0.002935005, 0.003011807,
  0.00245036, 0.002282623, 0.002114893, 0.002057691, 0.002153145, 
    0.002173588, 0.002178412, 0.002390604, 0.002481546, 0.002586848, 
    0.002681387, 0.002827789, 0.003032672, 0.003024529, 0.003101076,
  0.002476807, 0.002200748, 0.002120845, 0.002082671, 0.002169388, 
    0.002039466, 0.002116248, 0.002344007, 0.002461678, 0.00257708, 
    0.002700248, 0.003005545, 0.003145144, 0.00325433, 0.003338289,
  0.002428544, 0.002250782, 0.00216592, 0.002143171, 0.002169506, 
    0.002136183, 0.002068453, 0.002189402, 0.002339698, 0.002541919, 
    0.002760936, 0.003168309, 0.00325609, 0.003263393, 0.003420681,
  0.002358465, 0.002073506, 0.002182458, 0.002127144, 0.002152526, 
    0.002141628, 0.002135094, 0.001968577, 0.002056734, 0.002520142, 
    0.00289506, 0.003304311, 0.003304879, 0.003275581, 0.003396024,
  0.002216307, 0.002071857, 0.002133016, 0.002139475, 0.002166017, 
    0.002121464, 0.00218267, 0.002365491, 0.002579915, 0.002715833, 
    0.003124714, 0.003462652, 0.00331511, 0.003181322, 0.003256258,
  0.002181379, 0.002122381, 0.002146587, 0.002179489, 0.00218548, 
    0.002088232, 0.002158837, 0.002443011, 0.002672874, 0.002896452, 
    0.003297279, 0.003525177, 0.003354644, 0.003175974, 0.00316891,
  0.002181367, 0.002176163, 0.002200021, 0.002178806, 0.002172481, 
    0.00210845, 0.002239757, 0.002522555, 0.00275897, 0.003019642, 
    0.003382039, 0.003537731, 0.003439214, 0.00332735, 0.003128359,
  0.002172557, 0.00226441, 0.002317, 0.002210936, 0.002154676, 0.002135995, 
    0.002329239, 0.002639425, 0.002855468, 0.003137419, 0.003423454, 
    0.003522333, 0.003470945, 0.003385975, 0.003224138,
  0.002286327, 0.002423199, 0.002432583, 0.002224104, 0.002207943, 
    0.002184815, 0.002442233, 0.002719256, 0.002975466, 0.003288507, 
    0.003441965, 0.003498978, 0.003464213, 0.003437372, 0.003287548,
  0.002256578, 0.002276199, 0.002310039, 0.002221901, 0.002207727, 
    0.00224553, 0.002285959, 0.002399335, 0.002513106, 0.002654342, 
    0.002760304, 0.002993797, 0.003061201, 0.003045981, 0.003267521,
  0.002317671, 0.00226842, 0.002284801, 0.002285579, 0.002309972, 
    0.002249344, 0.002317439, 0.002340667, 0.002467022, 0.002611269, 
    0.002756803, 0.002893408, 0.002957143, 0.002949665, 0.003137326,
  0.002333709, 0.002273941, 0.002397284, 0.002374233, 0.002367689, 
    0.002255487, 0.002333226, 0.002439442, 0.002552477, 0.002590253, 
    0.002675464, 0.002777805, 0.002852679, 0.002913189, 0.003102561,
  0.002258245, 0.002368552, 0.002464043, 0.002464668, 0.00247525, 
    0.002504532, 0.002407587, 0.002543673, 0.002546377, 0.002549987, 
    0.002652354, 0.00276347, 0.002916429, 0.002979347, 0.003081287,
  0.002322477, 0.002360505, 0.002561784, 0.002631168, 0.002593806, 
    0.00268841, 0.002786976, 0.002368473, 0.002323807, 0.002602609, 
    0.002700266, 0.002800357, 0.003018673, 0.003075256, 0.003139021,
  0.002348225, 0.002584861, 0.002680226, 0.002765071, 0.002663542, 
    0.002818871, 0.00296681, 0.003017218, 0.002982841, 0.002939556, 
    0.002914529, 0.00289246, 0.003030347, 0.003125956, 0.003118671,
  0.002526627, 0.002775792, 0.002812827, 0.002757396, 0.002768843, 
    0.002983663, 0.003070636, 0.003102719, 0.003083334, 0.003075292, 
    0.003042683, 0.003024307, 0.003102005, 0.003041231, 0.003041961,
  0.002798613, 0.002942185, 0.002805126, 0.002736501, 0.00286277, 
    0.003079234, 0.003129396, 0.003149221, 0.003136446, 0.003116847, 
    0.003093333, 0.003160833, 0.003173101, 0.003108122, 0.003157013,
  0.002938342, 0.002895312, 0.002843451, 0.002787946, 0.002937333, 
    0.003151576, 0.003173678, 0.00320752, 0.003215858, 0.003213862, 
    0.003280644, 0.003322072, 0.003147613, 0.003216104, 0.003299203,
  0.002968598, 0.002959898, 0.002849669, 0.002922276, 0.003003101, 
    0.003195047, 0.003210735, 0.003244349, 0.003277004, 0.003322544, 
    0.003361032, 0.003383445, 0.003291557, 0.00332915, 0.003309417,
  0.002471925, 0.002394755, 0.002398608, 0.0025822, 0.00278426, 0.002829636, 
    0.002897623, 0.002999858, 0.00303608, 0.003065129, 0.003025466, 
    0.00288775, 0.002886131, 0.002640844, 0.002858354,
  0.00237379, 0.002253649, 0.0025139, 0.002917731, 0.002925445, 0.002937276, 
    0.003002374, 0.003083153, 0.0031592, 0.003174939, 0.003171207, 
    0.003009113, 0.002899311, 0.002747128, 0.002865823,
  0.002448348, 0.002497849, 0.002756667, 0.002976901, 0.003000017, 
    0.002858121, 0.003048546, 0.003122517, 0.003237084, 0.003246392, 
    0.003212977, 0.003118714, 0.002943912, 0.002895291, 0.002880416,
  0.002487587, 0.002782538, 0.00285017, 0.003003567, 0.003066036, 
    0.003212094, 0.002944679, 0.003020072, 0.003151698, 0.003237488, 
    0.003239935, 0.003154795, 0.002943554, 0.002911857, 0.002943591,
  0.002708793, 0.002938158, 0.002823213, 0.003013257, 0.003118876, 
    0.003281735, 0.003255186, 0.002796243, 0.002761941, 0.003212223, 
    0.003350019, 0.003236092, 0.003007597, 0.002926809, 0.002962194,
  0.00306221, 0.00301807, 0.002829915, 0.003027122, 0.003165883, 0.003315033, 
    0.003330175, 0.003349105, 0.003340118, 0.003402288, 0.003452537, 
    0.003318397, 0.003073576, 0.002933806, 0.002972787,
  0.003158541, 0.002977568, 0.002817749, 0.003093679, 0.003251469, 
    0.003367853, 0.003367646, 0.003380367, 0.003385243, 0.003406608, 
    0.003504227, 0.003362258, 0.003098388, 0.002894572, 0.002911668,
  0.003078138, 0.002878987, 0.002745174, 0.00315866, 0.003322063, 
    0.003401094, 0.003424625, 0.003413325, 0.003373453, 0.003391496, 
    0.00353637, 0.003472543, 0.003179577, 0.002882414, 0.002856987,
  0.002983755, 0.002839809, 0.002814402, 0.00319732, 0.003353338, 
    0.003431705, 0.003464672, 0.003434168, 0.003371078, 0.003366271, 
    0.003448798, 0.003561868, 0.003161101, 0.00286325, 0.002826223,
  0.003100547, 0.002984029, 0.002912493, 0.003195547, 0.003337994, 
    0.003416346, 0.003474729, 0.00345392, 0.003419936, 0.003363149, 
    0.003429078, 0.003538172, 0.003253599, 0.002877578, 0.00281063,
  0.002562635, 0.00266767, 0.002656814, 0.002740099, 0.002912275, 
    0.002956842, 0.002991586, 0.003033574, 0.003093434, 0.00317306, 
    0.003195219, 0.003076688, 0.00289202, 0.002646262, 0.002749063,
  0.00272404, 0.002674916, 0.0026936, 0.00294565, 0.003076816, 0.003085479, 
    0.003095877, 0.003064551, 0.003059247, 0.003210894, 0.003233102, 
    0.003044782, 0.002871585, 0.002715693, 0.002730932,
  0.002894665, 0.002788013, 0.002716824, 0.00306354, 0.003273907, 
    0.003022113, 0.003168069, 0.003157785, 0.003073054, 0.003160451, 
    0.003224621, 0.003262652, 0.002937808, 0.002887073, 0.003008947,
  0.00301369, 0.002818561, 0.002859307, 0.003187122, 0.003355525, 
    0.003434861, 0.003119157, 0.003192475, 0.003045876, 0.003175055, 
    0.003323434, 0.003333531, 0.00297599, 0.002913565, 0.002903228,
  0.003066532, 0.002869869, 0.002966693, 0.003245753, 0.003416622, 
    0.003539702, 0.003545298, 0.002968313, 0.002646232, 0.003226569, 
    0.003395263, 0.003330254, 0.003005598, 0.002925144, 0.002880287,
  0.003078318, 0.002987675, 0.00303598, 0.003319098, 0.003463228, 
    0.003568849, 0.003613455, 0.003349121, 0.00312424, 0.00336322, 
    0.003429473, 0.003290659, 0.003048141, 0.003025674, 0.00299172,
  0.003061262, 0.003044043, 0.003150855, 0.003353181, 0.003447382, 
    0.003546298, 0.003512667, 0.003357921, 0.003334677, 0.00343368, 
    0.003416036, 0.003284299, 0.003126091, 0.003109096, 0.003044132,
  0.003068221, 0.00303397, 0.003238934, 0.003355484, 0.0034005, 0.003437988, 
    0.00337626, 0.003315104, 0.003428521, 0.003452137, 0.003426154, 
    0.003259432, 0.003152597, 0.00314718, 0.003105293,
  0.003038942, 0.003052511, 0.003257606, 0.003335504, 0.003391002, 
    0.003398198, 0.003385744, 0.003353491, 0.003383136, 0.003459902, 
    0.003408845, 0.003232385, 0.003181284, 0.003159871, 0.003134084,
  0.003080571, 0.003143964, 0.003294265, 0.003362272, 0.003418553, 
    0.003434316, 0.00344401, 0.003383345, 0.003409063, 0.003432621, 
    0.003382582, 0.003219596, 0.003174707, 0.003137086, 0.003112121,
  0.002573937, 0.002620959, 0.002766988, 0.002873074, 0.003034233, 
    0.003124151, 0.003311723, 0.003273132, 0.003006808, 0.00295158, 
    0.002815667, 0.002700639, 0.002820674, 0.002679696, 0.00304904,
  0.002708938, 0.002938489, 0.002855056, 0.00288427, 0.003071458, 
    0.003339879, 0.003440145, 0.003444245, 0.003185993, 0.003041744, 
    0.002916954, 0.002707161, 0.00246824, 0.002616462, 0.003162451,
  0.002928107, 0.002841309, 0.002694135, 0.002813021, 0.003179424, 
    0.00321055, 0.003439014, 0.003474508, 0.003207321, 0.003118633, 
    0.002950542, 0.002805679, 0.002369002, 0.002677703, 0.003344872,
  0.002883743, 0.002746144, 0.00269283, 0.002987617, 0.003430422, 
    0.003510182, 0.003155324, 0.003372889, 0.003146295, 0.003096231, 
    0.002980058, 0.002850358, 0.002682089, 0.003019463, 0.003380679,
  0.002869524, 0.002722902, 0.002773697, 0.003248412, 0.003542124, 
    0.00344644, 0.003360078, 0.002711192, 0.002530564, 0.003050954, 
    0.003003963, 0.00296358, 0.0030052, 0.003178566, 0.003396162,
  0.002908185, 0.002782287, 0.002954452, 0.003358629, 0.003371029, 
    0.003436256, 0.003320026, 0.002952382, 0.002917374, 0.003009137, 
    0.003082597, 0.003115235, 0.003244602, 0.003300887, 0.003459573,
  0.002911642, 0.002817493, 0.003071112, 0.003329798, 0.003167813, 
    0.003061612, 0.002969672, 0.00292931, 0.003058899, 0.003159964, 
    0.003231383, 0.00329451, 0.003342067, 0.003382889, 0.00345165,
  0.002909183, 0.002842889, 0.003266771, 0.003304482, 0.003315463, 
    0.003262473, 0.003236176, 0.003217062, 0.003223481, 0.003269083, 
    0.003269595, 0.003301692, 0.003328663, 0.003333068, 0.003388734,
  0.002958573, 0.00308905, 0.003346157, 0.003324444, 0.003318371, 0.00331779, 
    0.003287435, 0.003289168, 0.003286386, 0.003256264, 0.003268282, 
    0.00328681, 0.003302473, 0.003330722, 0.003354979,
  0.002975588, 0.003270624, 0.003401895, 0.003415711, 0.00340182, 
    0.003364217, 0.003340338, 0.003276268, 0.00322324, 0.003205603, 
    0.003246147, 0.003266623, 0.003269901, 0.003284988, 0.003311233,
  0.003506077, 0.003263942, 0.003216129, 0.002974885, 0.002796155, 
    0.002744895, 0.002838403, 0.003131792, 0.003159787, 0.002694519, 
    0.003141455, 0.002746979, 0.002513786, 0.002657252, 0.003059604,
  0.003316854, 0.003197215, 0.003008078, 0.002728265, 0.002658505, 
    0.002908026, 0.003046867, 0.00314237, 0.00316704, 0.003085011, 
    0.00305424, 0.002560437, 0.002344328, 0.002700398, 0.003050724,
  0.003347398, 0.003085616, 0.002725889, 0.002575105, 0.002688332, 
    0.002776424, 0.003333796, 0.003385308, 0.003318135, 0.002999924, 
    0.002926561, 0.002706191, 0.002325919, 0.002595474, 0.003248278,
  0.003285831, 0.002906822, 0.002562158, 0.002495905, 0.002798946, 
    0.003135808, 0.002836044, 0.003399677, 0.003312672, 0.003068683, 
    0.002972432, 0.002751399, 0.002477792, 0.002789515, 0.003473098,
  0.003050679, 0.002674889, 0.00250277, 0.002642256, 0.002989069, 0.00333089, 
    0.003370112, 0.00278021, 0.002542247, 0.002833385, 0.002873232, 
    0.002559915, 0.002682985, 0.003268594, 0.003669228,
  0.002885628, 0.002641088, 0.002565376, 0.002875376, 0.003062733, 
    0.003226082, 0.003261471, 0.002882983, 0.002744124, 0.002710552, 
    0.00260341, 0.002707534, 0.003203498, 0.003632962, 0.003704047,
  0.002814965, 0.002654382, 0.002650853, 0.002864578, 0.0030422, 0.003090674, 
    0.003018314, 0.002861387, 0.002723453, 0.00271292, 0.002946013, 
    0.003161405, 0.003527372, 0.003685059, 0.00369938,
  0.002813979, 0.002771555, 0.003040542, 0.002840183, 0.002975409, 
    0.00301172, 0.003027136, 0.003040458, 0.003087596, 0.003220626, 
    0.003257994, 0.003492128, 0.00364154, 0.003660254, 0.003638204,
  0.002910682, 0.003069099, 0.003158536, 0.003090671, 0.003077411, 
    0.003141308, 0.003227646, 0.003295814, 0.003339075, 0.003366187, 
    0.00352392, 0.003623334, 0.003634743, 0.003617229, 0.00358338,
  0.00301599, 0.003124356, 0.003204226, 0.003117073, 0.00314893, 0.00318242, 
    0.003153742, 0.003225541, 0.003384922, 0.003515659, 0.003607733, 
    0.003619674, 0.003598568, 0.003564528, 0.003518612,
  0.005352847, 0.004075862, 0.004393763, 0.003480387, 0.003288331, 
    0.003106636, 0.002867039, 0.002814926, 0.00282716, 0.002945787, 
    0.002825507, 0.002619939, 0.002510667, 0.002720712, 0.002973268,
  0.003962945, 0.003780751, 0.003606422, 0.003291894, 0.003206281, 
    0.002982687, 0.002851569, 0.002808731, 0.002899359, 0.002875023, 
    0.002699086, 0.0022876, 0.002471191, 0.002671859, 0.002997274,
  0.0039211, 0.003697131, 0.003449706, 0.003193506, 0.003068339, 0.002806898, 
    0.002776313, 0.002754319, 0.002853138, 0.002664399, 0.002560091, 
    0.002474276, 0.002702703, 0.002801397, 0.003307965,
  0.003879969, 0.003600946, 0.003338838, 0.00313195, 0.002951382, 
    0.002817354, 0.002627777, 0.002828929, 0.002946039, 0.002710918, 
    0.002669649, 0.002742057, 0.002740853, 0.003001237, 0.003530554,
  0.00364225, 0.003341876, 0.003137452, 0.002931045, 0.002820287, 
    0.002823041, 0.002844522, 0.002594255, 0.002435644, 0.002605187, 
    0.002621052, 0.002644266, 0.0027878, 0.003353381, 0.003659302,
  0.003155299, 0.002981215, 0.002823217, 0.002739453, 0.002745362, 
    0.002888557, 0.002964922, 0.002791998, 0.002626257, 0.002588474, 
    0.002654796, 0.002708867, 0.003126743, 0.003599838, 0.003685518,
  0.002736859, 0.002629075, 0.002520424, 0.002775156, 0.002925149, 
    0.003016158, 0.003100445, 0.002876563, 0.00263626, 0.002692142, 
    0.002642434, 0.002912019, 0.003512057, 0.003661284, 0.003682178,
  0.002519367, 0.002428485, 0.002926224, 0.002714227, 0.002943009, 
    0.00309017, 0.003181738, 0.00291268, 0.00271803, 0.002642236, 
    0.002808661, 0.003391061, 0.003631738, 0.003653685, 0.003686272,
  0.002627661, 0.002717112, 0.002988507, 0.002990994, 0.003033933, 
    0.003073001, 0.003195641, 0.003064016, 0.002623232, 0.002728348, 
    0.003169744, 0.003616043, 0.003633587, 0.003634277, 0.003634014,
  0.002770915, 0.002878002, 0.003050266, 0.002930796, 0.003049689, 
    0.003120498, 0.003080896, 0.002901271, 0.002873187, 0.003186044, 
    0.003627679, 0.003640628, 0.003610621, 0.003596763, 0.003568919,
  0.006419483, 0.004975914, 0.00557236, 0.004152661, 0.003862522, 
    0.003630489, 0.003425476, 0.003266354, 0.003134561, 0.003107334, 
    0.003025692, 0.002871685, 0.002757013, 0.00261023, 0.00273182,
  0.004763334, 0.004494915, 0.004173465, 0.003743554, 0.003688925, 
    0.003527537, 0.00334156, 0.003123543, 0.002973644, 0.002925095, 
    0.002805662, 0.002614876, 0.002493304, 0.002543924, 0.002727112,
  0.004530817, 0.004267276, 0.003838796, 0.003574731, 0.003468917, 
    0.003293794, 0.0031068, 0.002928806, 0.002758063, 0.002601657, 
    0.002507356, 0.002511796, 0.002597889, 0.002697997, 0.003146299,
  0.004519406, 0.004163117, 0.003752665, 0.00353491, 0.003323048, 0.00305448, 
    0.002786336, 0.002806717, 0.002625797, 0.002440088, 0.002382611, 
    0.002565253, 0.002739976, 0.003135547, 0.003533738,
  0.004444832, 0.003989377, 0.003708069, 0.00343275, 0.003236209, 
    0.002918397, 0.002710371, 0.002376672, 0.002211547, 0.002332663, 
    0.002444687, 0.002839654, 0.00330354, 0.003596833, 0.003699113,
  0.00431719, 0.003878986, 0.003527679, 0.003273792, 0.00311576, 0.002839869, 
    0.002698651, 0.002572581, 0.002601813, 0.002634944, 0.002731732, 
    0.00323301, 0.003591022, 0.003683442, 0.003698276,
  0.004091286, 0.003775207, 0.003380009, 0.003166693, 0.003006664, 
    0.002841146, 0.002752896, 0.002615723, 0.002589101, 0.002671598, 
    0.002997923, 0.003518516, 0.003652902, 0.003679711, 0.003712332,
  0.003760995, 0.003527789, 0.003173695, 0.003033383, 0.002884412, 
    0.002792062, 0.002778868, 0.002623249, 0.00249427, 0.002560846, 
    0.003251465, 0.0035879, 0.003635475, 0.003685565, 0.003715061,
  0.003452953, 0.003233477, 0.003005784, 0.002946465, 0.002828314, 
    0.002777227, 0.002795215, 0.002517379, 0.002339333, 0.002843722, 
    0.003440412, 0.003619384, 0.003631884, 0.003653977, 0.003672163,
  0.003231653, 0.003094976, 0.002966075, 0.002899292, 0.002823171, 
    0.002784317, 0.002829885, 0.002833377, 0.002778661, 0.00315398, 
    0.003566989, 0.003638133, 0.003612374, 0.003593338, 0.00356362,
  0.005527923, 0.004640535, 0.005188029, 0.004399619, 0.004319856, 
    0.004320093, 0.004106665, 0.003828174, 0.003626247, 0.003615435, 
    0.003528295, 0.003165987, 0.002933834, 0.00277885, 0.002630771,
  0.004241121, 0.004172189, 0.004173533, 0.004071536, 0.004233961, 
    0.003904311, 0.003854664, 0.003697007, 0.00358587, 0.003480091, 
    0.003269344, 0.002950547, 0.002661899, 0.002714539, 0.002879363,
  0.004378444, 0.004238581, 0.004065173, 0.004065818, 0.003809539, 
    0.003845559, 0.003687249, 0.00359451, 0.003430421, 0.003184247, 
    0.002964657, 0.00269079, 0.002502498, 0.002518424, 0.002961508,
  0.004461398, 0.004205644, 0.003983141, 0.003875128, 0.003669377, 
    0.003567413, 0.003306711, 0.003233282, 0.003111482, 0.00294083, 
    0.002671855, 0.002504635, 0.002764026, 0.002988273, 0.003224314,
  0.00451884, 0.004111383, 0.003951444, 0.003764544, 0.003649911, 
    0.003403071, 0.003194683, 0.002914199, 0.002517659, 0.002671448, 
    0.002608275, 0.002815411, 0.003106195, 0.003391636, 0.003543759,
  0.004533597, 0.004092967, 0.003774056, 0.003635007, 0.003494804, 
    0.003227867, 0.003047894, 0.002928255, 0.002732686, 0.002703584, 
    0.00271521, 0.00315049, 0.003473347, 0.003637982, 0.003678482,
  0.00447678, 0.004072579, 0.003636207, 0.003379453, 0.003070842, 
    0.002806175, 0.002754973, 0.002714337, 0.002701702, 0.002941674, 
    0.00334742, 0.003595961, 0.003661358, 0.003650697, 0.003616828,
  0.004434214, 0.003952415, 0.003397162, 0.00305709, 0.002833228, 
    0.002778169, 0.002855222, 0.002967367, 0.003122425, 0.003497354, 
    0.003641023, 0.003650772, 0.003638328, 0.003637788, 0.003624247,
  0.004150697, 0.003593055, 0.003073267, 0.002859626, 0.002828127, 0.0028384, 
    0.002917382, 0.003073447, 0.003344213, 0.003608086, 0.003654805, 
    0.003649087, 0.003644496, 0.003640056, 0.003637178,
  0.00381239, 0.00330701, 0.002997048, 0.002861677, 0.002869977, 0.002899863, 
    0.002983541, 0.003188381, 0.003400497, 0.0036125, 0.00364365, 0.00363095, 
    0.003606032, 0.003588875, 0.003554419,
  0.004095216, 0.00370648, 0.004172163, 0.003919837, 0.00399834, 0.003978968, 
    0.003916197, 0.003938984, 0.004082974, 0.003974371, 0.003811656, 
    0.003595053, 0.003444513, 0.003634907, 0.003718552,
  0.004113457, 0.003790418, 0.00379076, 0.003745425, 0.003914812, 
    0.003802566, 0.00381149, 0.003931057, 0.003974709, 0.00391496, 
    0.003725973, 0.00353297, 0.003415331, 0.003437587, 0.003453018,
  0.004362618, 0.004089459, 0.003870755, 0.003725586, 0.003780709, 
    0.003865069, 0.00374342, 0.003848863, 0.003922985, 0.003902039, 
    0.003706367, 0.003531266, 0.003361706, 0.003302443, 0.003255328,
  0.004440519, 0.004211539, 0.003953911, 0.003826609, 0.003730212, 
    0.003731019, 0.003965269, 0.003843471, 0.003875703, 0.003790623, 
    0.003686828, 0.003486321, 0.003408711, 0.003265161, 0.003107914,
  0.004458425, 0.004143961, 0.003999481, 0.003847419, 0.003807564, 
    0.003597839, 0.003644582, 0.003910865, 0.003706448, 0.003704183, 
    0.003625032, 0.003502016, 0.003294843, 0.003140175, 0.003101652,
  0.004383679, 0.004135876, 0.003897518, 0.003823935, 0.003810931, 
    0.003834722, 0.003783426, 0.003654449, 0.003527049, 0.003497506, 
    0.003445115, 0.003338378, 0.003208036, 0.003158984, 0.003235784,
  0.004245054, 0.004045694, 0.003750835, 0.003691411, 0.003663405, 
    0.003603609, 0.003538864, 0.003419689, 0.003319774, 0.003287817, 
    0.00326634, 0.003246904, 0.003276592, 0.003365579, 0.003422188,
  0.004020405, 0.003813236, 0.003484487, 0.003410263, 0.00339789, 
    0.003357713, 0.003281318, 0.003258784, 0.003236843, 0.003295586, 
    0.003366045, 0.003409427, 0.003485244, 0.003539931, 0.003546404,
  0.003703748, 0.003476171, 0.003277384, 0.003303793, 0.00333729, 
    0.003360178, 0.003384158, 0.003439849, 0.003544512, 0.00357496, 
    0.003566786, 0.003591212, 0.003612407, 0.003600611, 0.003584682,
  0.003561139, 0.003400465, 0.003296678, 0.003349188, 0.003482438, 
    0.003578622, 0.003639172, 0.00362954, 0.003668967, 0.003671747, 
    0.003669213, 0.003615381, 0.003479292, 0.00327793, 0.00340197,
  0.004577772, 0.004018121, 0.004355425, 0.003972348, 0.003875495, 
    0.003971213, 0.00392131, 0.003851247, 0.003781231, 0.003796627, 
    0.003984944, 0.003879256, 0.003812062, 0.00398943, 0.003971563,
  0.003993856, 0.003823977, 0.003802353, 0.00376048, 0.003841701, 
    0.003881025, 0.003885631, 0.003816816, 0.003736178, 0.003722272, 
    0.00381624, 0.003801961, 0.003750767, 0.003947758, 0.003889849,
  0.004212066, 0.004061363, 0.003914405, 0.003700516, 0.003768937, 
    0.003864372, 0.003849174, 0.003792631, 0.003780164, 0.003703214, 
    0.003734603, 0.003743112, 0.003685725, 0.003839007, 0.003768678,
  0.004326959, 0.004141533, 0.003963287, 0.003809733, 0.003706312, 
    0.003812286, 0.003937217, 0.003868839, 0.003819016, 0.003781791, 
    0.003743362, 0.003694304, 0.003619296, 0.003785633, 0.003691998,
  0.004392824, 0.004064004, 0.003924957, 0.003751608, 0.003757241, 
    0.003770059, 0.003817619, 0.004028707, 0.003929878, 0.003827085, 
    0.003763839, 0.003662435, 0.003699958, 0.003702495, 0.003602243,
  0.004352686, 0.004066572, 0.003831753, 0.003717409, 0.003728528, 
    0.003788194, 0.003786933, 0.003752233, 0.003763689, 0.003766812, 
    0.003773813, 0.003708658, 0.003677643, 0.00363601, 0.003559669,
  0.004329206, 0.004095177, 0.003755212, 0.003684125, 0.003708854, 
    0.003716838, 0.003730165, 0.003739126, 0.003747339, 0.003740234, 
    0.003740231, 0.003692644, 0.003617893, 0.003521527, 0.003445684,
  0.004184198, 0.003929361, 0.003646911, 0.003607558, 0.003641099, 
    0.003671836, 0.003682391, 0.003697367, 0.003701276, 0.003697479, 
    0.003663113, 0.003588716, 0.003488896, 0.003402669, 0.003368798,
  0.003977186, 0.003781708, 0.003556854, 0.003551945, 0.003563548, 
    0.003573032, 0.003590703, 0.003594719, 0.003601589, 0.003599282, 
    0.003556496, 0.003510351, 0.003456013, 0.003453292, 0.003478991,
  0.003879569, 0.003758856, 0.003594476, 0.003580739, 0.003563931, 
    0.003552637, 0.003536957, 0.003540478, 0.003596399, 0.003607374, 
    0.003579453, 0.00350443, 0.003445049, 0.003457369, 0.003581242,
  0.004317152, 0.00398067, 0.004445626, 0.004023666, 0.004055714, 
    0.004405046, 0.004211536, 0.004006306, 0.004153015, 0.003730841, 
    0.003895445, 0.00405925, 0.004006664, 0.004093372, 0.004022195,
  0.004007159, 0.003866175, 0.003846607, 0.003756748, 0.003872087, 
    0.003996195, 0.004032813, 0.003890364, 0.003864457, 0.003546306, 
    0.00371449, 0.003914732, 0.003976148, 0.004066919, 0.003947868,
  0.004164326, 0.004097636, 0.003984497, 0.003692859, 0.003775004, 
    0.003932491, 0.003930435, 0.003840405, 0.003816568, 0.003489369, 
    0.003653127, 0.003830735, 0.00389926, 0.003943107, 0.003846948,
  0.004074844, 0.003984732, 0.003927835, 0.003814843, 0.003716295, 
    0.003805553, 0.003930227, 0.003760698, 0.003703421, 0.003505626, 
    0.003701715, 0.003799413, 0.003795248, 0.00388409, 0.003794706,
  0.003924906, 0.003867961, 0.003841036, 0.00375792, 0.003728265, 0.00375333, 
    0.003817082, 0.00392073, 0.003860109, 0.003609046, 0.003714954, 
    0.00378048, 0.003782782, 0.003846907, 0.0038668,
  0.003817841, 0.003830642, 0.00377073, 0.003657811, 0.003714004, 
    0.003754117, 0.003804781, 0.003731028, 0.003728393, 0.003673384, 
    0.003722268, 0.003765983, 0.00376635, 0.00381959, 0.00381292,
  0.00373009, 0.003791478, 0.003718395, 0.003654317, 0.003701611, 0.00376203, 
    0.003810661, 0.003758056, 0.003699627, 0.003629721, 0.003673865, 
    0.003675584, 0.003739316, 0.003811101, 0.003750171,
  0.003634324, 0.003702805, 0.003624951, 0.003669, 0.003718747, 0.003775891, 
    0.003772006, 0.003743508, 0.003701734, 0.003613905, 0.003630196, 
    0.00362447, 0.003703556, 0.003716701, 0.003650578,
  0.003484901, 0.003510553, 0.003503283, 0.003641015, 0.003735327, 
    0.00376666, 0.003738907, 0.003654582, 0.003605261, 0.003626899, 
    0.003715702, 0.003624249, 0.0036712, 0.003675255, 0.003641885,
  0.003312474, 0.003284479, 0.003364612, 0.003518698, 0.003661979, 
    0.003703272, 0.003657736, 0.003620238, 0.00362495, 0.003659979, 
    0.003608948, 0.003635683, 0.003615428, 0.003606881, 0.003617145,
  0.004017376, 0.003728673, 0.003898028, 0.003658428, 0.003743894, 
    0.003885835, 0.00379466, 0.003760903, 0.003857755, 0.003805212, 
    0.004086569, 0.004072133, 0.00395415, 0.004068504, 0.004020636,
  0.003882137, 0.003715515, 0.003673499, 0.003583245, 0.003694941, 
    0.003718453, 0.003726827, 0.003726784, 0.003749799, 0.003732353, 
    0.00394848, 0.003922866, 0.003946194, 0.004010011, 0.003986678,
  0.003844634, 0.003755188, 0.003727192, 0.003581643, 0.003656742, 
    0.00369926, 0.003746296, 0.003775641, 0.003784765, 0.003685263, 
    0.00367342, 0.003739315, 0.003903314, 0.003958145, 0.003979824,
  0.003951812, 0.003915233, 0.003860228, 0.003751668, 0.003666076, 
    0.003697522, 0.003715442, 0.003703279, 0.003786366, 0.003605111, 
    0.003695829, 0.003789471, 0.00387956, 0.003905153, 0.003841358,
  0.004034906, 0.003964266, 0.003917701, 0.003771702, 0.003736542, 
    0.003691747, 0.003682792, 0.003750677, 0.003990491, 0.003635402, 
    0.003645429, 0.003787551, 0.003856586, 0.003891964, 0.003931068,
  0.004067614, 0.004009947, 0.003890082, 0.003706903, 0.003728251, 
    0.003719199, 0.003715601, 0.003683015, 0.003717191, 0.003606913, 
    0.003747207, 0.003793027, 0.003843577, 0.003856929, 0.003842615,
  0.004057255, 0.00408119, 0.003835494, 0.003596677, 0.00365957, 0.003698497, 
    0.00372132, 0.003735279, 0.003646491, 0.003598605, 0.003714545, 
    0.003787953, 0.003807101, 0.003777683, 0.003711094,
  0.004089961, 0.004014657, 0.003664046, 0.003576278, 0.003645486, 
    0.003688793, 0.003701624, 0.003710938, 0.003671749, 0.003646782, 
    0.003725498, 0.003742008, 0.003746546, 0.003680649, 0.003628526,
  0.003974634, 0.003926645, 0.003656902, 0.003669611, 0.003681615, 
    0.003705068, 0.003696301, 0.003679474, 0.003672734, 0.003659782, 
    0.00373025, 0.003707092, 0.003705522, 0.003674492, 0.003666236,
  0.003857675, 0.003912207, 0.003765777, 0.00374277, 0.003724763, 
    0.003711639, 0.003654299, 0.003634853, 0.003654998, 0.003698232, 
    0.00367519, 0.0036874, 0.003684616, 0.003659198, 0.003662176,
  0.005225115, 0.004439325, 0.004885283, 0.004091873, 0.003995848, 
    0.004167886, 0.003864588, 0.003744609, 0.003663691, 0.003592907, 
    0.003712787, 0.003738593, 0.003720863, 0.003750117, 0.003697298,
  0.004310056, 0.00401032, 0.004044116, 0.003767733, 0.003899463, 
    0.003990655, 0.003824504, 0.003745253, 0.0036711, 0.003620469, 
    0.003721163, 0.003725723, 0.003720827, 0.003797182, 0.003865519,
  0.004322732, 0.004117075, 0.00389953, 0.003589005, 0.003649232, 
    0.003706954, 0.003647225, 0.003677393, 0.003671647, 0.003624532, 
    0.00363026, 0.003696595, 0.003708771, 0.003750275, 0.00381832,
  0.004085425, 0.004004641, 0.003911672, 0.00380678, 0.003666534, 
    0.003699852, 0.003694057, 0.003688128, 0.003624372, 0.003640221, 
    0.003661508, 0.003695382, 0.003717584, 0.003720125, 0.003755274,
  0.004101302, 0.00411399, 0.004045532, 0.003832079, 0.003788905, 0.00374761, 
    0.003733135, 0.003479643, 0.003431128, 0.003625123, 0.003629656, 
    0.003714254, 0.003748298, 0.003737635, 0.003803155,
  0.004358937, 0.004248704, 0.004049819, 0.003741979, 0.003740364, 
    0.003752433, 0.003744869, 0.003614471, 0.003588168, 0.003613062, 
    0.003689026, 0.00366293, 0.00365263, 0.003713379, 0.003793334,
  0.004433581, 0.004272909, 0.003836646, 0.003520786, 0.003572743, 
    0.003665821, 0.003717029, 0.003708779, 0.003623699, 0.003539205, 
    0.003585749, 0.003632672, 0.003683517, 0.003681564, 0.003711364,
  0.004330311, 0.003859418, 0.003624454, 0.003485213, 0.003594313, 
    0.003664124, 0.003685941, 0.00365505, 0.003617452, 0.003634899, 
    0.003638204, 0.003687085, 0.003687503, 0.00365676, 0.003632079,
  0.004015577, 0.003869516, 0.003613665, 0.003646438, 0.003664023, 
    0.00368339, 0.003663947, 0.003613045, 0.003656716, 0.003698698, 
    0.003729407, 0.003701608, 0.003669989, 0.003633809, 0.003591408,
  0.003965264, 0.003860351, 0.003724774, 0.003701794, 0.003688221, 
    0.003667859, 0.003618967, 0.003557749, 0.00369661, 0.003752948, 
    0.003749351, 0.003691938, 0.003641135, 0.003590642, 0.003521488,
  0.006779321, 0.005142569, 0.005927658, 0.004443092, 0.004358677, 
    0.004907922, 0.004252255, 0.003984889, 0.004144134, 0.004758029, 
    0.004586207, 0.004264683, 0.00366784, 0.003741747, 0.003687793,
  0.00505955, 0.004660718, 0.004621404, 0.004121403, 0.004622187, 
    0.004865791, 0.003914837, 0.00379615, 0.003889195, 0.004219634, 
    0.003987107, 0.003703974, 0.003608104, 0.003530452, 0.003588706,
  0.004621478, 0.004485135, 0.004185619, 0.003892804, 0.004090715, 
    0.004096819, 0.003763991, 0.003667128, 0.003634596, 0.003615023, 
    0.003432221, 0.003448001, 0.003482326, 0.003531145, 0.003644202,
  0.004277708, 0.004200398, 0.00403059, 0.003929795, 0.003764968, 
    0.003821156, 0.00377376, 0.003565766, 0.003459903, 0.003385419, 
    0.003366387, 0.003413593, 0.003470119, 0.003516747, 0.003652421,
  0.00419755, 0.0041037, 0.003995244, 0.003766144, 0.003718772, 0.003680384, 
    0.003687945, 0.003724983, 0.003592358, 0.00335384, 0.003368203, 
    0.003373991, 0.003505519, 0.003531158, 0.00357225,
  0.004327164, 0.004225425, 0.003934636, 0.003649937, 0.003673212, 0.0037056, 
    0.003681754, 0.00366186, 0.003587724, 0.003476776, 0.003425515, 
    0.003408471, 0.003239624, 0.003506703, 0.003562019,
  0.004375311, 0.004314355, 0.003904435, 0.003601145, 0.003553986, 
    0.003641594, 0.00368813, 0.003705048, 0.003660801, 0.003498167, 
    0.003583145, 0.003512563, 0.003266441, 0.003499931, 0.003436625,
  0.004440296, 0.004228078, 0.003819734, 0.003633258, 0.003614704, 
    0.003631022, 0.003643676, 0.003648952, 0.003681099, 0.003626132, 
    0.00360752, 0.003479991, 0.003314551, 0.003461615, 0.003318906,
  0.004323624, 0.004101267, 0.003757518, 0.003722172, 0.003693939, 
    0.003675542, 0.003653776, 0.003657503, 0.003693342, 0.00369124, 
    0.003592697, 0.003429657, 0.003472095, 0.003499897, 0.003254799,
  0.004189234, 0.004038902, 0.003826181, 0.003761722, 0.003717867, 
    0.003683522, 0.003627555, 0.003623528, 0.003688587, 0.003675482, 
    0.003549737, 0.003443113, 0.003575601, 0.003464645, 0.003165409,
  0.004797311, 0.004591998, 0.005549639, 0.004272943, 0.004522379, 
    0.004897947, 0.004234114, 0.00421886, 0.004682174, 0.005663034, 
    0.00502969, 0.004205684, 0.003757468, 0.003630539, 0.003804195,
  0.004274101, 0.004387013, 0.004512896, 0.004321691, 0.004947383, 
    0.004744755, 0.004038999, 0.004082529, 0.004211407, 0.004466791, 
    0.004183263, 0.003528035, 0.003292959, 0.003379778, 0.003685762,
  0.00439127, 0.004511352, 0.004324462, 0.0041536, 0.00424961, 0.004020671, 
    0.003947197, 0.003841301, 0.003833243, 0.003637712, 0.00346665, 
    0.003280777, 0.003219166, 0.003508525, 0.003677287,
  0.00433214, 0.004390488, 0.004296163, 0.004176734, 0.003933277, 
    0.004006227, 0.003897837, 0.003766798, 0.00361874, 0.003417987, 
    0.003318158, 0.00324237, 0.00321471, 0.003437595, 0.003579085,
  0.00424604, 0.004182588, 0.004158094, 0.003961439, 0.003895193, 0.00387839, 
    0.003866448, 0.003939265, 0.003659312, 0.003402361, 0.003303362, 
    0.003226198, 0.003167051, 0.003360372, 0.003484132,
  0.004144898, 0.004079465, 0.003885134, 0.00373461, 0.003772134, 
    0.003841082, 0.003810189, 0.003724258, 0.003626433, 0.00344796, 
    0.00327332, 0.003166443, 0.003127942, 0.003252079, 0.003397017,
  0.004040016, 0.00402952, 0.0037159, 0.003582298, 0.003606562, 0.003790606, 
    0.003823849, 0.003715027, 0.003524993, 0.003377635, 0.003309368, 
    0.003115452, 0.002980613, 0.002928345, 0.002992298,
  0.004179524, 0.003850871, 0.003700726, 0.003595924, 0.003647693, 
    0.003746418, 0.003749481, 0.003619488, 0.003490871, 0.00346413, 
    0.003369247, 0.003185489, 0.002938938, 0.002860625, 0.002783315,
  0.004263597, 0.003807824, 0.00363674, 0.003722352, 0.003729795, 
    0.003743174, 0.00371995, 0.003631265, 0.003584778, 0.003553041, 
    0.003409743, 0.003056723, 0.002904914, 0.00279737, 0.0027214,
  0.004198238, 0.003920384, 0.003714445, 0.003736897, 0.003749542, 
    0.003736197, 0.003691946, 0.003633653, 0.003637934, 0.003601142, 
    0.003389983, 0.003019732, 0.002935508, 0.002752542, 0.002603386,
  0.003663004, 0.003788437, 0.004396066, 0.003841618, 0.004213545, 
    0.004442162, 0.003995018, 0.00414126, 0.004320701, 0.005022061, 
    0.005107011, 0.004613657, 0.004163635, 0.004022573, 0.004134074,
  0.003772837, 0.003917601, 0.004055291, 0.003939236, 0.004510188, 
    0.004385501, 0.00389936, 0.003937828, 0.004003893, 0.004165758, 
    0.004452001, 0.003818069, 0.003700931, 0.0036541, 0.003786535,
  0.003972259, 0.004062309, 0.004106872, 0.003896768, 0.004024317, 
    0.003876689, 0.003813941, 0.003747132, 0.003715794, 0.003643613, 
    0.003579869, 0.003530995, 0.003566619, 0.003711377, 0.003755905,
  0.004148727, 0.004076741, 0.004093442, 0.003967358, 0.003664797, 
    0.003732446, 0.003626279, 0.00353498, 0.003389232, 0.003401155, 
    0.003436575, 0.00346521, 0.003472072, 0.003543558, 0.003470018,
  0.004226859, 0.004014644, 0.004025347, 0.003859944, 0.003700488, 
    0.003624757, 0.003565877, 0.003382508, 0.002923619, 0.003276244, 
    0.003292202, 0.003249548, 0.003159194, 0.003180006, 0.003092516,
  0.004282606, 0.00402614, 0.003882759, 0.003757674, 0.003685588, 
    0.003644893, 0.003518837, 0.003402057, 0.003276994, 0.003153969, 
    0.003142625, 0.00303277, 0.002909831, 0.002786257, 0.002795663,
  0.004297456, 0.004108677, 0.0037422, 0.003624691, 0.003585065, 0.003616424, 
    0.003528292, 0.003398557, 0.003210346, 0.003103254, 0.003046454, 
    0.002855653, 0.002659914, 0.002625499, 0.002561667,
  0.004178014, 0.004124686, 0.00356871, 0.003540706, 0.003579398, 
    0.003630735, 0.003459726, 0.003315536, 0.003112443, 0.003007608, 
    0.002884988, 0.002616307, 0.002492561, 0.002406268, 0.002379506,
  0.004420948, 0.004057494, 0.003586331, 0.00365448, 0.003661117, 0.00365293, 
    0.003435899, 0.003270665, 0.003087058, 0.00297547, 0.002713851, 
    0.002544272, 0.002448017, 0.002404144, 0.002433505,
  0.00445765, 0.004051869, 0.003719359, 0.003750788, 0.003743307, 
    0.003679271, 0.003394109, 0.003261576, 0.003039806, 0.002848955, 
    0.002628804, 0.002528028, 0.002432629, 0.002371121, 0.002453376,
  0.005853028, 0.004310134, 0.00463291, 0.003892678, 0.004087208, 
    0.004399817, 0.003968023, 0.004130744, 0.004366331, 0.005293381, 
    0.00517423, 0.004765355, 0.004605495, 0.00450968, 0.00442926,
  0.004419203, 0.004142478, 0.004186285, 0.003948925, 0.00456107, 
    0.004320932, 0.003877302, 0.003926256, 0.003921362, 0.004259254, 
    0.004450481, 0.00404704, 0.003904115, 0.003738046, 0.003909385,
  0.004521651, 0.004274802, 0.004154145, 0.003926228, 0.004331545, 
    0.003837966, 0.003807031, 0.00372776, 0.003733019, 0.003691751, 
    0.003803033, 0.003575078, 0.003503979, 0.003482125, 0.003393803,
  0.004599418, 0.004364075, 0.004157765, 0.004023421, 0.003792324, 
    0.003776699, 0.003710056, 0.003631323, 0.003626846, 0.003642953, 
    0.003609651, 0.00345356, 0.003275035, 0.003167728, 0.003103575,
  0.004532485, 0.004253005, 0.004131925, 0.003891869, 0.003675224, 
    0.003629655, 0.003627535, 0.003331305, 0.003181813, 0.003576174, 
    0.003421772, 0.003062405, 0.002861684, 0.002841055, 0.002934158,
  0.004454643, 0.004202331, 0.003996707, 0.003701456, 0.003612146, 
    0.003626566, 0.003537756, 0.003416239, 0.003400752, 0.003355443, 
    0.003077338, 0.002749939, 0.00265007, 0.002619589, 0.002756467,
  0.004380819, 0.004188192, 0.003796852, 0.003582665, 0.003543033, 
    0.003548545, 0.003534937, 0.003361244, 0.003292121, 0.003029105, 
    0.002803107, 0.002612757, 0.002535854, 0.002472328, 0.002661997,
  0.004300545, 0.004078026, 0.003598072, 0.003514207, 0.003498524, 
    0.003515675, 0.00338238, 0.003317478, 0.003147189, 0.002858264, 
    0.002560144, 0.002431949, 0.002289902, 0.002486414, 0.002792762,
  0.004252626, 0.003876944, 0.003520142, 0.003562152, 0.003571418, 
    0.003536889, 0.003346133, 0.003234541, 0.002974481, 0.002694041, 
    0.002463048, 0.002332424, 0.002379881, 0.002808249, 0.003136676,
  0.004294202, 0.003904822, 0.003644444, 0.003679612, 0.003670902, 
    0.003548342, 0.003254489, 0.003093967, 0.002866569, 0.002557038, 
    0.002398103, 0.002352141, 0.002541754, 0.003015813, 0.003267439,
  0.004651412, 0.003974164, 0.004232773, 0.003774706, 0.004150323, 
    0.00447804, 0.004041263, 0.003963464, 0.004178569, 0.005855378, 
    0.005635452, 0.004752561, 0.004464049, 0.004185088, 0.004144765,
  0.003977223, 0.003846189, 0.003806909, 0.003709936, 0.004137252, 
    0.004236963, 0.003866463, 0.003913113, 0.003948994, 0.00458177, 
    0.00520255, 0.004409042, 0.003889269, 0.003508599, 0.00356225,
  0.003968964, 0.003864472, 0.003740528, 0.003599783, 0.003764995, 
    0.00363753, 0.003799123, 0.003827536, 0.003881744, 0.003979273, 
    0.00436048, 0.003949197, 0.003620218, 0.003278836, 0.003233419,
  0.003859699, 0.003843043, 0.003678062, 0.003696886, 0.003582262, 
    0.003691157, 0.003620993, 0.003675976, 0.003735898, 0.003832164, 
    0.003893199, 0.003716753, 0.00337172, 0.003124437, 0.003078873,
  0.003645729, 0.003626011, 0.003641182, 0.003582121, 0.003512276, 
    0.003511278, 0.00368554, 0.003534575, 0.003544625, 0.003784693, 
    0.003739335, 0.00354599, 0.003236367, 0.003032596, 0.003014948,
  0.003620132, 0.003647493, 0.003655936, 0.003511527, 0.003477886, 
    0.003543543, 0.003620464, 0.003615555, 0.003606891, 0.00364851, 
    0.003591746, 0.003366055, 0.00309458, 0.002907549, 0.00303193,
  0.004014716, 0.003992471, 0.003722949, 0.003511009, 0.003484266, 
    0.003495716, 0.003614116, 0.003632787, 0.003587936, 0.003539426, 
    0.003408467, 0.003164991, 0.002897528, 0.002769571, 0.002753141,
  0.004144042, 0.004026317, 0.003656528, 0.003496232, 0.003462713, 
    0.003500608, 0.003591717, 0.003580174, 0.003570342, 0.003518101, 
    0.003280558, 0.002956922, 0.002748806, 0.002703466, 0.002781146,
  0.004071941, 0.003825642, 0.003581631, 0.003523861, 0.003492948, 
    0.003534228, 0.003590858, 0.003596156, 0.003573106, 0.003404017, 
    0.003038697, 0.00281498, 0.002735224, 0.002934718, 0.003010811,
  0.004061535, 0.003902613, 0.003620504, 0.003603724, 0.003644962, 
    0.003631821, 0.003588185, 0.003526682, 0.003395526, 0.003070162, 
    0.002772018, 0.002702198, 0.003054029, 0.003352098, 0.003469491,
  0.006528313, 0.00526787, 0.006091077, 0.004491266, 0.004406638, 
    0.004444389, 0.0041456, 0.004095568, 0.004384747, 0.005541279, 
    0.006305137, 0.006005729, 0.005834167, 0.004920316, 0.004343819,
  0.004256694, 0.004182772, 0.004113325, 0.0039147, 0.004095772, 0.003830702, 
    0.003698929, 0.003760457, 0.003801082, 0.004105416, 0.005065346, 
    0.004737635, 0.004801223, 0.004499238, 0.004239298,
  0.004117718, 0.004017309, 0.003861938, 0.003707784, 0.00377665, 
    0.003358073, 0.003343109, 0.003290634, 0.003516922, 0.003595208, 
    0.003899058, 0.003977385, 0.004010956, 0.00409036, 0.004020117,
  0.003953766, 0.003774997, 0.003580177, 0.003441629, 0.003331664, 
    0.003329653, 0.003104954, 0.003158053, 0.003263071, 0.00332229, 
    0.003553327, 0.003711967, 0.003820917, 0.003841335, 0.003755915,
  0.00360228, 0.003469837, 0.003421544, 0.003397403, 0.003321832, 
    0.003263413, 0.003147263, 0.002912031, 0.002866863, 0.003249204, 
    0.003231746, 0.00350401, 0.003728668, 0.003701167, 0.003596552,
  0.003557546, 0.003606831, 0.003603383, 0.00346614, 0.003384326, 
    0.003429625, 0.003472789, 0.003422934, 0.003317625, 0.003202993, 
    0.003201464, 0.003384435, 0.003637643, 0.003622391, 0.003492506,
  0.003675473, 0.003729044, 0.003628377, 0.003471536, 0.003450444, 
    0.003423989, 0.003521452, 0.003576518, 0.003559545, 0.003438844, 
    0.003394204, 0.003450501, 0.003610282, 0.003539144, 0.003421667,
  0.003857005, 0.003608497, 0.003611489, 0.003519512, 0.003468557, 
    0.003441432, 0.003536551, 0.003602629, 0.003607588, 0.003604402, 
    0.003542873, 0.003542195, 0.003590715, 0.003439088, 0.003222986,
  0.003509229, 0.003816601, 0.003643135, 0.003581417, 0.003455492, 
    0.003493522, 0.003567609, 0.003635272, 0.003661984, 0.003629792, 
    0.003592377, 0.003594813, 0.003541498, 0.003285243, 0.003102438,
  0.003687562, 0.003879077, 0.003761601, 0.003550166, 0.003564735, 
    0.003625246, 0.003551885, 0.003635004, 0.003672707, 0.003630876, 
    0.003599564, 0.003551626, 0.003403991, 0.003174417, 0.003077863,
  0.003797268, 0.003768719, 0.00428535, 0.003933571, 0.00406978, 0.004521029, 
    0.004296311, 0.004246464, 0.004345674, 0.005834336, 0.006568232, 
    0.006531525, 0.007065004, 0.00680187, 0.005909367,
  0.003824772, 0.003811854, 0.003893779, 0.003786735, 0.004276691, 
    0.004328167, 0.004041849, 0.004056883, 0.004062954, 0.004449677, 
    0.005355439, 0.004845622, 0.005095398, 0.005693929, 0.005630817,
  0.003897174, 0.00386021, 0.003795813, 0.003746842, 0.004101778, 
    0.003853149, 0.003928494, 0.0038764, 0.003877855, 0.003907633, 
    0.004176721, 0.004090431, 0.004099742, 0.00442567, 0.004814136,
  0.003772102, 0.00368972, 0.003584573, 0.003621996, 0.00361039, 0.003862736, 
    0.003590423, 0.003659681, 0.003611026, 0.003643752, 0.003675866, 
    0.003666993, 0.003801126, 0.003903294, 0.004064377,
  0.003680364, 0.003575217, 0.00343858, 0.003416253, 0.003340037, 
    0.003419536, 0.003531603, 0.003321982, 0.003120666, 0.003428919, 
    0.003412595, 0.00336554, 0.003526542, 0.003766593, 0.003882392,
  0.003791316, 0.003474897, 0.003450199, 0.003373202, 0.003324304, 
    0.003355903, 0.00341718, 0.003426072, 0.003378577, 0.003249917, 
    0.00317999, 0.003141838, 0.003322686, 0.003702252, 0.003752034,
  0.003739352, 0.003434288, 0.003509094, 0.003394401, 0.003386662, 
    0.00338942, 0.003413571, 0.003398827, 0.003391803, 0.00324474, 
    0.003209475, 0.003181953, 0.003266077, 0.003621038, 0.0037362,
  0.003744011, 0.003528888, 0.003541989, 0.003421327, 0.003382198, 
    0.003432039, 0.003411111, 0.003358061, 0.003464996, 0.003360403, 
    0.003368237, 0.003412163, 0.003556643, 0.003667732, 0.003684111,
  0.0034511, 0.003659027, 0.003527536, 0.003474434, 0.003446637, 0.003456572, 
    0.003534402, 0.003601565, 0.00362511, 0.00361475, 0.003598635, 
    0.003573923, 0.003599278, 0.003579868, 0.00343827,
  0.003389167, 0.003651994, 0.003570351, 0.003512242, 0.003577911, 
    0.003554711, 0.003464933, 0.003449074, 0.003576697, 0.003618674, 
    0.003574216, 0.003563882, 0.003536892, 0.00337072, 0.00320932,
  0.003733405, 0.003605075, 0.003602934, 0.003319036, 0.003425287, 
    0.003528783, 0.003366405, 0.003352433, 0.003426629, 0.003798881, 
    0.00402482, 0.004093037, 0.004298054, 0.004656576, 0.005217423,
  0.003709339, 0.003552347, 0.003385196, 0.003301159, 0.003395648, 
    0.003384573, 0.003259423, 0.003345854, 0.003405832, 0.003596157, 
    0.003907762, 0.003927755, 0.003968508, 0.004121465, 0.004470911,
  0.00380134, 0.003462567, 0.003313386, 0.003208558, 0.003166625, 
    0.003090569, 0.003243809, 0.00334046, 0.003392398, 0.003397319, 
    0.003576059, 0.003807105, 0.003821456, 0.003893076, 0.004151531,
  0.004075019, 0.003645386, 0.003484328, 0.003131071, 0.003196563, 
    0.003079101, 0.003115917, 0.003272906, 0.00322922, 0.003326416, 
    0.003636717, 0.003796761, 0.003809989, 0.00381616, 0.003913225,
  0.004197241, 0.003972064, 0.003378728, 0.003102351, 0.003141875, 
    0.003299714, 0.003218172, 0.003004161, 0.00296821, 0.003372368, 
    0.003732172, 0.003825726, 0.003814204, 0.003798617, 0.003849152,
  0.004286928, 0.004108909, 0.003590101, 0.003407062, 0.003362402, 
    0.003378297, 0.003405674, 0.003167744, 0.003124773, 0.003477318, 
    0.003777725, 0.003811812, 0.003801339, 0.003847765, 0.003898275,
  0.004177825, 0.003889229, 0.003612535, 0.003434359, 0.003422202, 
    0.003394906, 0.003396441, 0.003309485, 0.003359962, 0.003558249, 
    0.003706011, 0.00375459, 0.003725548, 0.00374225, 0.003731537,
  0.004015086, 0.003364007, 0.003428434, 0.003446886, 0.003453798, 
    0.003431936, 0.003472481, 0.003406643, 0.003522576, 0.003629529, 
    0.003736774, 0.003720136, 0.003650817, 0.003626627, 0.003606127,
  0.003653858, 0.003522151, 0.003512588, 0.00349022, 0.003490684, 
    0.003456989, 0.003522073, 0.003523329, 0.003580209, 0.003666971, 
    0.003726478, 0.003698716, 0.003600632, 0.003525403, 0.003469937,
  0.003666021, 0.003514032, 0.003568191, 0.003534216, 0.003493497, 
    0.003500598, 0.003446056, 0.00350593, 0.003419542, 0.003626061, 
    0.003679344, 0.003651808, 0.003550004, 0.003446834, 0.003431701,
  0.004837724, 0.004692601, 0.006111139, 0.004626386, 0.004693931, 
    0.005593006, 0.004472414, 0.004112347, 0.004094479, 0.004654168, 
    0.004473598, 0.004045814, 0.003989719, 0.004057277, 0.004223429,
  0.003977145, 0.00408721, 0.004301192, 0.004217466, 0.004936396, 
    0.004617619, 0.003890807, 0.003802735, 0.003756912, 0.003913513, 
    0.0040734, 0.003813071, 0.003706226, 0.003818189, 0.004064944,
  0.003873046, 0.003990192, 0.003989534, 0.003930838, 0.004129092, 
    0.003669231, 0.003659521, 0.003582219, 0.003522594, 0.003505645, 
    0.003628293, 0.003686792, 0.003549779, 0.003634477, 0.003948524,
  0.00364435, 0.003692391, 0.003667753, 0.00366451, 0.003610672, 0.003603637, 
    0.003353795, 0.003410565, 0.003358395, 0.003395263, 0.003627887, 
    0.003609745, 0.003396054, 0.003587947, 0.003897787,
  0.003509503, 0.003437229, 0.003356514, 0.00338165, 0.003391364, 
    0.003480557, 0.003341467, 0.003061729, 0.002913338, 0.003392623, 
    0.00362847, 0.003524791, 0.00336545, 0.003566266, 0.003618636,
  0.003475478, 0.00334505, 0.003331879, 0.003344346, 0.00331229, 0.003342269, 
    0.003395281, 0.00319466, 0.003225733, 0.003539335, 0.003522871, 
    0.003533294, 0.003394705, 0.003548868, 0.003537155,
  0.003461898, 0.003307765, 0.003309801, 0.003315689, 0.003317915, 
    0.003332324, 0.003323993, 0.003373385, 0.003449676, 0.003511597, 
    0.003534186, 0.003520784, 0.003418922, 0.00345906, 0.003473134,
  0.003505071, 0.003221611, 0.003321157, 0.003296124, 0.003289122, 
    0.003247411, 0.003184507, 0.003160188, 0.003472193, 0.003545571, 
    0.003588906, 0.003480007, 0.003398788, 0.00350488, 0.003448412,
  0.003621781, 0.00349292, 0.003460904, 0.003439093, 0.003349918, 
    0.003276612, 0.003171873, 0.00316572, 0.003465204, 0.00359694, 
    0.003494621, 0.003407879, 0.003478816, 0.003509799, 0.00345942,
  0.003582309, 0.003544456, 0.003534077, 0.003508355, 0.003388566, 
    0.003364061, 0.003084685, 0.003167444, 0.003429565, 0.003295234, 
    0.003450447, 0.003420065, 0.003265726, 0.003458113, 0.00333579,
  0.003855289, 0.003945656, 0.004564035, 0.004004606, 0.004329359, 
    0.005993624, 0.005129867, 0.005063323, 0.00551952, 0.00931668, 
    0.00861134, 0.006841415, 0.00583503, 0.00507152, 0.004798797,
  0.003755238, 0.003883244, 0.003986083, 0.00391839, 0.005060511, 
    0.006224781, 0.00443305, 0.00445823, 0.004643641, 0.006141597, 
    0.007954011, 0.00550977, 0.004678096, 0.004703329, 0.00458598,
  0.003638122, 0.003818526, 0.004013005, 0.003912694, 0.004809811, 
    0.004648738, 0.004461102, 0.004075918, 0.004161717, 0.004563871, 
    0.005082532, 0.004516353, 0.004135147, 0.003996288, 0.004130342,
  0.003489723, 0.003679475, 0.003811918, 0.00397632, 0.003993939, 
    0.004951133, 0.004218844, 0.004053088, 0.003985474, 0.004059883, 
    0.004108961, 0.003975621, 0.003794435, 0.003693335, 0.003944161,
  0.003377462, 0.003465407, 0.003653508, 0.00372458, 0.003692659, 
    0.003956163, 0.004197345, 0.004318238, 0.004376594, 0.004428461, 
    0.003906073, 0.00383046, 0.003631303, 0.003605479, 0.003702424,
  0.00326587, 0.003382175, 0.003430818, 0.003571256, 0.003574607, 
    0.003709141, 0.003909198, 0.004055106, 0.004439919, 0.004023845, 
    0.003816549, 0.00365453, 0.003546176, 0.003534647, 0.003422322,
  0.003290004, 0.003323911, 0.003268599, 0.003424658, 0.003529276, 
    0.003572982, 0.003663416, 0.003866889, 0.003852171, 0.003701698, 
    0.003671698, 0.003600375, 0.003497001, 0.00342697, 0.003311712,
  0.003458063, 0.003299872, 0.003184594, 0.003329211, 0.003418531, 
    0.003504819, 0.003554154, 0.003670917, 0.003663389, 0.003631869, 
    0.003583187, 0.00348914, 0.003453467, 0.003371556, 0.003329176,
  0.00361955, 0.003302894, 0.003165669, 0.003232981, 0.003302942, 
    0.003373879, 0.003541681, 0.003640155, 0.003612692, 0.003564109, 
    0.00347511, 0.003393287, 0.003328393, 0.003333658, 0.003443307,
  0.003663944, 0.003517177, 0.003129216, 0.003178922, 0.003222178, 
    0.003288272, 0.003396096, 0.003498699, 0.003503521, 0.003428845, 
    0.003314585, 0.003232606, 0.00316272, 0.003266587, 0.003405401,
  0.003685011, 0.003879458, 0.004269832, 0.003945498, 0.004605622, 
    0.005713613, 0.004925458, 0.004945342, 0.005555459, 0.01079451, 
    0.01104336, 0.009472773, 0.009699243, 0.008324606, 0.007469548,
  0.003593748, 0.003619878, 0.00370472, 0.003870196, 0.004932858, 
    0.005224013, 0.004013399, 0.004271525, 0.004294327, 0.006143617, 
    0.01034843, 0.007922011, 0.006907204, 0.008235756, 0.007086581,
  0.003408382, 0.003469625, 0.003605745, 0.003610117, 0.003935212, 
    0.00393946, 0.004282555, 0.003988026, 0.004043411, 0.004287405, 
    0.005557167, 0.005189542, 0.004904166, 0.00557052, 0.005966696,
  0.00333759, 0.003310634, 0.00336197, 0.003520059, 0.003471625, 0.003904599, 
    0.003913743, 0.0042893, 0.00399452, 0.004017107, 0.00425638, 0.004499582, 
    0.004201565, 0.004719961, 0.005239985,
  0.00336465, 0.003188058, 0.003210372, 0.003414421, 0.003364896, 
    0.003419853, 0.003707448, 0.003980679, 0.004379422, 0.004789571, 
    0.003982256, 0.004113233, 0.004090056, 0.004178906, 0.004316712,
  0.003406653, 0.003240013, 0.003143536, 0.003378296, 0.003313791, 
    0.00334976, 0.00343273, 0.003577499, 0.004063977, 0.00404483, 
    0.004431411, 0.004001676, 0.003951963, 0.003940624, 0.004011942,
  0.003598749, 0.003390792, 0.003115222, 0.003355924, 0.003321134, 
    0.003337053, 0.003374861, 0.003497845, 0.003586513, 0.003697615, 
    0.003840206, 0.003934927, 0.003876776, 0.003843362, 0.003861466,
  0.003656671, 0.003521736, 0.003104179, 0.003329327, 0.003294171, 
    0.003331043, 0.003377794, 0.003489336, 0.00359736, 0.003712142, 
    0.003780954, 0.003831114, 0.003837934, 0.003794062, 0.003784593,
  0.003816271, 0.003412215, 0.003076857, 0.003337678, 0.003331289, 
    0.003266655, 0.00340015, 0.003568341, 0.003680429, 0.003761227, 
    0.003792219, 0.003798687, 0.003788329, 0.003747658, 0.003748578,
  0.003905533, 0.003383199, 0.003130707, 0.003325296, 0.003336754, 
    0.003308287, 0.003363923, 0.003532497, 0.003673096, 0.003765515, 
    0.003802769, 0.003767986, 0.003732257, 0.003704884, 0.003748195,
  0.003850346, 0.00404425, 0.004991103, 0.004737658, 0.005380753, 
    0.006601301, 0.0051316, 0.005030091, 0.006580524, 0.01119078, 0.01150998, 
    0.01029137, 0.01129228, 0.01041108, 0.01013341,
  0.003724327, 0.003785484, 0.004031555, 0.004642287, 0.006404015, 
    0.006151134, 0.004434456, 0.004538123, 0.005075237, 0.006889544, 
    0.01095957, 0.007584006, 0.006963092, 0.0108165, 0.01017104,
  0.003672775, 0.003730277, 0.003788477, 0.003958452, 0.004822031, 
    0.00426187, 0.00440153, 0.004223675, 0.004430359, 0.004668441, 
    0.005612204, 0.005422794, 0.004791189, 0.005706744, 0.008170893,
  0.003591676, 0.00359688, 0.003567605, 0.003661535, 0.00384321, 0.004609004, 
    0.004086253, 0.004298786, 0.004022995, 0.00406803, 0.004144238, 
    0.004114322, 0.004123753, 0.004546187, 0.006688714,
  0.003594699, 0.003467497, 0.003422292, 0.003405982, 0.003402457, 
    0.003693526, 0.004222478, 0.004179848, 0.004007407, 0.004106039, 
    0.003904185, 0.003903655, 0.003927322, 0.003938755, 0.004456148,
  0.003626887, 0.003518897, 0.003260115, 0.003253625, 0.003257057, 
    0.003346866, 0.00349209, 0.003652036, 0.003707305, 0.003712484, 
    0.003912199, 0.003731989, 0.003805955, 0.003813225, 0.003878187,
  0.003713483, 0.00383728, 0.003324896, 0.003183759, 0.0031215, 0.003179289, 
    0.003248258, 0.00335573, 0.003370908, 0.003422009, 0.003502179, 
    0.003663321, 0.003696759, 0.003728866, 0.003760961,
  0.004015473, 0.004182907, 0.003642043, 0.003144759, 0.003014605, 
    0.003065328, 0.003077911, 0.003186986, 0.003243014, 0.003391919, 
    0.003470297, 0.003590264, 0.003618427, 0.003627426, 0.003705938,
  0.00405049, 0.003755702, 0.003515343, 0.003346521, 0.002894508, 
    0.002828786, 0.002941168, 0.003039374, 0.003142113, 0.003232021, 
    0.003354044, 0.00347393, 0.003510299, 0.003562666, 0.003640904,
  0.004198946, 0.004055617, 0.003681662, 0.003423079, 0.003183301, 
    0.002851529, 0.002824774, 0.002898844, 0.002985392, 0.003094113, 
    0.003191799, 0.003284679, 0.003347973, 0.003431258, 0.003565686,
  0.004023871, 0.004105258, 0.004351567, 0.004038975, 0.004611154, 
    0.005942853, 0.005094214, 0.005190107, 0.006138201, 0.01105648, 
    0.01121232, 0.01028356, 0.01120334, 0.01036802, 0.01037729,
  0.003910614, 0.00403764, 0.0040758, 0.004021073, 0.005849987, 0.00656944, 
    0.00450231, 0.004893174, 0.00546834, 0.006829595, 0.01086233, 
    0.007792918, 0.00812799, 0.01080112, 0.01069372,
  0.00395435, 0.004088139, 0.00413138, 0.004159377, 0.005885946, 0.004599595, 
    0.004713749, 0.00448954, 0.004879147, 0.005244444, 0.00642986, 
    0.00669763, 0.005803511, 0.006139253, 0.009217522,
  0.00392467, 0.003927086, 0.004067918, 0.004331164, 0.004671389, 
    0.005613855, 0.004473573, 0.00502964, 0.004633381, 0.004676378, 
    0.004865831, 0.005042133, 0.004738844, 0.005077135, 0.007078908,
  0.003795662, 0.00372616, 0.003796139, 0.003916365, 0.003987591, 
    0.004591019, 0.004985896, 0.004778714, 0.005001607, 0.005257593, 
    0.00456077, 0.004595912, 0.004515543, 0.004467403, 0.004932785,
  0.003938273, 0.003597276, 0.00354519, 0.003569922, 0.003685047, 
    0.003989304, 0.004477633, 0.00472686, 0.005789388, 0.005105447, 
    0.004993484, 0.00437089, 0.004280351, 0.004184009, 0.004182503,
  0.003929187, 0.00354265, 0.003365789, 0.003367235, 0.003555988, 
    0.003697169, 0.003935373, 0.004272341, 0.004529286, 0.004218505, 
    0.004224596, 0.004133691, 0.00409587, 0.004058583, 0.00401845,
  0.00386844, 0.00356233, 0.00329054, 0.003249667, 0.003355109, 0.003573809, 
    0.003612873, 0.003890421, 0.00406429, 0.00403075, 0.004034976, 
    0.003951485, 0.003920003, 0.003869516, 0.003955847,
  0.003811145, 0.003679619, 0.003362873, 0.003177135, 0.0031367, 0.003303402, 
    0.003515891, 0.003697933, 0.003792387, 0.003822026, 0.003842022, 
    0.00379274, 0.003733392, 0.003678499, 0.003758931,
  0.00402038, 0.003992262, 0.003465307, 0.003323159, 0.003123809, 
    0.003073641, 0.003269169, 0.003459828, 0.00357319, 0.003633407, 
    0.003647032, 0.003586128, 0.00352853, 0.003474938, 0.003514434,
  0.003866677, 0.00391637, 0.004193766, 0.003958089, 0.004047876, 
    0.004213444, 0.003865599, 0.004004826, 0.004466728, 0.01091296, 
    0.01079896, 0.009519359, 0.01001713, 0.009369325, 0.009040846,
  0.003861233, 0.003895503, 0.004031448, 0.003939218, 0.004246192, 
    0.004353972, 0.0039759, 0.004067258, 0.004268444, 0.006494997, 
    0.01044801, 0.008033818, 0.007955531, 0.009642051, 0.009411842,
  0.003862004, 0.003986234, 0.004136659, 0.003949569, 0.004265129, 
    0.003950498, 0.004240151, 0.0041195, 0.004114913, 0.005277447, 
    0.006928584, 0.006891948, 0.005837682, 0.005365967, 0.008551666,
  0.003781697, 0.003848037, 0.004058294, 0.004099178, 0.004035166, 
    0.00457739, 0.004228771, 0.004576492, 0.004151735, 0.00460432, 
    0.004982912, 0.004954162, 0.004810101, 0.005079193, 0.007121265,
  0.003710749, 0.003687725, 0.00377256, 0.003994837, 0.003893207, 
    0.003965132, 0.004650872, 0.004510793, 0.00467959, 0.005180036, 
    0.00455155, 0.004537554, 0.004587272, 0.004525877, 0.004733809,
  0.00398071, 0.00357186, 0.003593774, 0.003603137, 0.003757707, 0.003799586, 
    0.003935449, 0.004277907, 0.005588823, 0.005216605, 0.005238127, 
    0.004420199, 0.004364324, 0.004396567, 0.004218682,
  0.003664025, 0.00347523, 0.003482223, 0.003479981, 0.00361751, 0.00375302, 
    0.00385537, 0.004004628, 0.00429818, 0.004175764, 0.00434884, 
    0.004338165, 0.00424852, 0.004287458, 0.004174955,
  0.003511115, 0.003403017, 0.003359486, 0.003412195, 0.003488892, 
    0.003621625, 0.003696038, 0.003881705, 0.004055026, 0.004130019, 
    0.004161078, 0.004233522, 0.004173432, 0.004230306, 0.00419153,
  0.003577895, 0.003389717, 0.00330505, 0.003299642, 0.003354367, 
    0.003473219, 0.003659618, 0.003852679, 0.004001212, 0.004088083, 
    0.004113615, 0.004112953, 0.004141281, 0.004141227, 0.004180904,
  0.003801725, 0.003451837, 0.003317756, 0.003286403, 0.003297613, 
    0.003354308, 0.003638913, 0.003793674, 0.003924753, 0.004021948, 
    0.004113134, 0.004074271, 0.004051307, 0.003994623, 0.004133043,
  0.003909171, 0.003728815, 0.003930378, 0.003840366, 0.003752419, 
    0.003893807, 0.003725272, 0.003675812, 0.003747024, 0.006361892, 
    0.008897002, 0.008174461, 0.007903298, 0.007708987, 0.007782138,
  0.003905132, 0.003797938, 0.00376686, 0.003762352, 0.003880844, 
    0.003908335, 0.003722216, 0.003702999, 0.003682997, 0.004656288, 
    0.0083287, 0.007118522, 0.0068936, 0.007750343, 0.008034582,
  0.003994422, 0.003933364, 0.00391358, 0.003814889, 0.003954625, 
    0.003748467, 0.003931739, 0.003789994, 0.003778189, 0.00412533, 
    0.0060497, 0.006499897, 0.005392725, 0.005108977, 0.00753658,
  0.004122571, 0.003875389, 0.003809693, 0.003859311, 0.003846598, 
    0.004070425, 0.003856268, 0.004115009, 0.003970113, 0.004146488, 
    0.004513535, 0.00446529, 0.004198572, 0.005049737, 0.007027236,
  0.004120284, 0.003712169, 0.00371992, 0.003926433, 0.003759906, 
    0.003854691, 0.004321751, 0.004103151, 0.004297956, 0.004772096, 
    0.004122849, 0.004106523, 0.003979817, 0.004336783, 0.004707993,
  0.004218637, 0.003573445, 0.00359999, 0.003685929, 0.003733861, 
    0.003735736, 0.003725303, 0.00400801, 0.005006844, 0.0050496, 
    0.004773432, 0.00407314, 0.003987845, 0.004074575, 0.004129449,
  0.004041937, 0.003445518, 0.003485426, 0.003509095, 0.00370388, 
    0.003750538, 0.003670094, 0.003694767, 0.003955889, 0.004177605, 
    0.004076072, 0.003972908, 0.004051998, 0.004062969, 0.004086233,
  0.003882741, 0.003373286, 0.00341171, 0.003478165, 0.003548617, 0.00370028, 
    0.003549418, 0.003603323, 0.003839894, 0.004020141, 0.004002954, 
    0.004062068, 0.004086454, 0.003997829, 0.003922372,
  0.003933262, 0.003317531, 0.003333692, 0.003419057, 0.003441741, 
    0.003501674, 0.00348403, 0.003644736, 0.003832595, 0.003957141, 
    0.003953471, 0.004055496, 0.004047768, 0.00406031, 0.004135339,
  0.004019734, 0.003424104, 0.003283049, 0.003303637, 0.003422029, 
    0.003444012, 0.003555438, 0.003656062, 0.003797261, 0.003868585, 
    0.003997931, 0.004008973, 0.003983081, 0.003980203, 0.004209472,
  0.004064866, 0.003875114, 0.004095922, 0.003716289, 0.003636429, 
    0.003557174, 0.003346733, 0.003353163, 0.003468577, 0.004216614, 
    0.005545596, 0.007156952, 0.007971506, 0.007918334, 0.007907867,
  0.003979325, 0.003852707, 0.003837878, 0.003702823, 0.003651657, 
    0.003544864, 0.003320152, 0.003381945, 0.003436325, 0.003922211, 
    0.005138685, 0.006587908, 0.00716678, 0.007776647, 0.007951519,
  0.004075447, 0.004073229, 0.004020643, 0.003720186, 0.003667325, 
    0.003440979, 0.003302024, 0.003367505, 0.003506302, 0.003702638, 
    0.004761968, 0.006250926, 0.005770283, 0.005487892, 0.007124272,
  0.004306993, 0.004236782, 0.004041594, 0.003810883, 0.003533963, 
    0.003393579, 0.003289989, 0.003551132, 0.00351246, 0.003849357, 
    0.003875281, 0.004169865, 0.004402518, 0.00518429, 0.00646593,
  0.004459398, 0.004266905, 0.003871469, 0.003502465, 0.003308592, 
    0.003302228, 0.00340531, 0.003160332, 0.003365658, 0.004119575, 
    0.003914501, 0.003758822, 0.004161495, 0.004660011, 0.005063234,
  0.004567116, 0.004130423, 0.003596196, 0.003357707, 0.003299495, 
    0.003299413, 0.003363166, 0.003381141, 0.003570936, 0.003905605, 
    0.004117053, 0.003670906, 0.003961579, 0.004301138, 0.004579076,
  0.004390055, 0.003948854, 0.003656586, 0.003489124, 0.003510689, 
    0.003499595, 0.003437543, 0.003373174, 0.003353406, 0.003458925, 
    0.003618838, 0.003683021, 0.003951904, 0.004166996, 0.004289485,
  0.004226296, 0.004075443, 0.003756311, 0.003585269, 0.003540652, 
    0.003546117, 0.003462834, 0.003419703, 0.003368813, 0.003464537, 
    0.003580344, 0.003713115, 0.003941125, 0.004065525, 0.004116254,
  0.004338141, 0.004168054, 0.003723569, 0.00352681, 0.003461333, 
    0.003423512, 0.003353768, 0.003491334, 0.003487228, 0.003573862, 
    0.003614001, 0.003724499, 0.003857281, 0.004002362, 0.004241135,
  0.004436906, 0.004290433, 0.003685254, 0.003436793, 0.003469037, 
    0.003359029, 0.003391381, 0.003474202, 0.003474073, 0.003697004, 
    0.003712084, 0.003750931, 0.003839497, 0.003950357, 0.004315779,
  0.003914619, 0.003871237, 0.003867427, 0.003653501, 0.003575881, 
    0.003343848, 0.003227726, 0.003412024, 0.003680477, 0.004690233, 
    0.006939432, 0.007945639, 0.00873948, 0.009152628, 0.009537729,
  0.004039139, 0.003869885, 0.003802045, 0.003612559, 0.00369036, 
    0.003416413, 0.003252866, 0.003267246, 0.003551546, 0.00404494, 
    0.006220207, 0.007215368, 0.007461271, 0.008960775, 0.009362794,
  0.004157203, 0.004035825, 0.003987421, 0.003730637, 0.003601213, 
    0.00326656, 0.003254301, 0.003243784, 0.00341423, 0.003700785, 
    0.004852145, 0.006441742, 0.006070239, 0.00535595, 0.007699552,
  0.004434297, 0.004212331, 0.003997938, 0.003950467, 0.003688953, 
    0.003321735, 0.003038352, 0.003180022, 0.003224182, 0.003433061, 
    0.003610718, 0.004015783, 0.004141239, 0.00485939, 0.006756961,
  0.004585173, 0.004341973, 0.004037062, 0.003828758, 0.003518979, 
    0.003366826, 0.003158514, 0.002978744, 0.002953495, 0.003230783, 
    0.003463991, 0.003615703, 0.00396694, 0.004412157, 0.005089546,
  0.004504573, 0.004377133, 0.004123049, 0.003832836, 0.003620841, 
    0.003477279, 0.003334162, 0.003164869, 0.003141739, 0.003138134, 
    0.003265288, 0.003450186, 0.00375384, 0.004052563, 0.004675598,
  0.004287852, 0.004310204, 0.003964846, 0.003752275, 0.003724232, 
    0.003698251, 0.003560559, 0.003346474, 0.003286002, 0.003110623, 
    0.00306238, 0.003301208, 0.003628566, 0.003885286, 0.004177291,
  0.003900056, 0.004050318, 0.003802713, 0.003645574, 0.003625094, 
    0.003683025, 0.00361888, 0.003533996, 0.003448843, 0.003306027, 
    0.003142396, 0.003195352, 0.003532556, 0.003760111, 0.003965139,
  0.003708094, 0.003716772, 0.003618621, 0.003543385, 0.003482637, 
    0.003504047, 0.003484118, 0.003543298, 0.003575483, 0.003412887, 
    0.003241214, 0.003194373, 0.003409244, 0.003693517, 0.004018453,
  0.003672285, 0.003650319, 0.003556414, 0.003528291, 0.003512886, 
    0.003417205, 0.003394474, 0.003506209, 0.003546659, 0.003530687, 
    0.003397214, 0.003247583, 0.003393465, 0.003651729, 0.004123297 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;
}
