netcdf tracer_level.0002-0002.radon {
dimensions:
	bnds = 2 ;
	lat = 18 ;
	lon = 29 ;
	pfull = 65 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	float radon(time, pfull, lat, lon) ;
		radon:_FillValue = -1.e+10f ;
		radon:missing_value = -1.e+10f ;
		radon:units = "vmr*1e21" ;
		radon:long_name = "radon-222" ;
		radon:interp_method = "conserve_order1" ;
		radon:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 17:15:31 2024" ;
		:hostname = "pp329" ;
		:history = "Tue Aug 12 16:31:13 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0002-0002.radon.nc reduced/tracer_level.0002-0002.radon.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00020101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 radon =
  5.84339e-21, 5.84339e-21, 5.84339e-21, 5.84339e-21, 5.84339e-21, 
    5.84339e-21, 5.84339e-21, 5.85205e-21, 5.85205e-21, 5.85205e-21, 
    5.85205e-21, 5.85205e-21, 5.85205e-21, 5.85205e-21, 5.599931e-21, 
    5.599931e-21, 5.599931e-21, 5.599931e-21, 5.599931e-21, 5.599931e-21, 
    5.599931e-21, 5.548771e-21, 5.548771e-21, 5.548771e-21, 5.548771e-21, 
    5.548771e-21, 5.548771e-21, 5.548771e-21, 5.84339e-21,
  1.198741e-20, 1.299412e-20, 1.395899e-20, 1.41411e-20, 1.44535e-20, 
    1.441263e-20, 1.422459e-20, 1.413948e-20, 1.395243e-20, 1.382196e-20, 
    1.385767e-20, 1.356916e-20, 1.342116e-20, 1.309725e-20, 1.223367e-20, 
    1.132538e-20, 1.055133e-20, 9.848495e-21, 8.995003e-21, 8.414929e-21, 
    8.158891e-21, 8.272644e-21, 8.636143e-21, 8.988981e-21, 9.159225e-21, 
    9.668289e-21, 1.03914e-20, 1.115577e-20, 1.17925e-20,
  3.988212e-20, 4.192882e-20, 4.235576e-20, 4.312869e-20, 4.347288e-20, 
    4.301136e-20, 4.148279e-20, 3.984913e-20, 3.773708e-20, 3.562445e-20, 
    3.3724e-20, 3.150882e-20, 3.049929e-20, 2.94706e-20, 2.798438e-20, 
    2.682879e-20, 2.511883e-20, 2.309388e-20, 2.138211e-20, 2.008185e-20, 
    2.097233e-20, 2.439631e-20, 2.506329e-20, 2.674843e-20, 3.110935e-20, 
    3.530936e-20, 3.747691e-20, 3.845483e-20, 3.929381e-20,
  9.23977e-20, 8.989233e-20, 8.9078e-20, 8.494835e-20, 7.88697e-20, 
    7.185045e-20, 6.958999e-20, 6.886071e-20, 6.775045e-20, 6.822258e-20, 
    6.768512e-20, 6.54755e-20, 6.390265e-20, 6.282017e-20, 6.01831e-20, 
    5.848478e-20, 5.845113e-20, 5.612616e-20, 6.12331e-20, 6.632685e-20, 
    6.852493e-20, 7.516223e-20, 7.436023e-20, 7.682494e-20, 8.144852e-20, 
    8.587138e-20, 8.673109e-20, 8.954943e-20, 9.353769e-20,
  1.676626e-19, 1.600606e-19, 1.576191e-19, 1.575593e-19, 1.611268e-19, 
    1.581065e-19, 1.487266e-19, 1.5056e-19, 1.457768e-19, 1.433591e-19, 
    1.476282e-19, 1.489915e-19, 1.504677e-19, 1.581947e-19, 1.610768e-19, 
    1.662772e-19, 1.694416e-19, 1.643467e-19, 1.632436e-19, 1.68068e-19, 
    1.656754e-19, 1.645962e-19, 1.739198e-19, 1.728013e-19, 1.665438e-19, 
    1.666085e-19, 1.60743e-19, 1.61974e-19, 1.644189e-19,
  5.017099e-19, 4.677956e-19, 4.884215e-19, 4.654161e-19, 4.419133e-19, 
    4.394227e-19, 4.101568e-19, 4.166481e-19, 4.188666e-19, 4.211412e-19, 
    4.174287e-19, 4.103794e-19, 4.105997e-19, 4.174788e-19, 4.282823e-19, 
    4.233993e-19, 4.435461e-19, 4.492687e-19, 4.732326e-19, 4.733919e-19, 
    4.663231e-19, 4.668501e-19, 4.771285e-19, 4.6415e-19, 4.637538e-19, 
    4.70485e-19, 4.914007e-19, 4.968845e-19, 4.93063e-19,
  7.159445e-19, 7.0666e-19, 7.315589e-19, 7.256269e-19, 7.31208e-19, 
    7.773026e-19, 7.291497e-19, 7.126458e-19, 6.763248e-19, 6.460242e-19, 
    6.370277e-19, 6.332769e-19, 6.325801e-19, 6.452814e-19, 6.616452e-19, 
    6.68401e-19, 6.812757e-19, 6.784512e-19, 6.693791e-19, 6.612863e-19, 
    6.51095e-19, 6.447277e-19, 6.36117e-19, 6.390991e-19, 6.653711e-19, 
    7.085907e-19, 7.518243e-19, 7.394156e-19, 7.164423e-19,
  1.256679e-18, 1.284313e-18, 1.296225e-18, 1.263281e-18, 1.333639e-18, 
    1.367417e-18, 1.401715e-18, 1.378492e-18, 1.323475e-18, 1.22865e-18, 
    1.174052e-18, 1.059855e-18, 1.011895e-18, 1.014956e-18, 1.004562e-18, 
    1.002404e-18, 1.012907e-18, 1.018147e-18, 9.778554e-19, 1.023645e-18, 
    1.046083e-18, 1.09245e-18, 1.140773e-18, 1.186175e-18, 1.173745e-18, 
    1.220771e-18, 1.247251e-18, 1.292161e-18, 1.246758e-18,
  1.933289e-18, 2.010366e-18, 1.962795e-18, 1.876074e-18, 1.923072e-18, 
    1.913945e-18, 1.84059e-18, 1.829779e-18, 1.772057e-18, 1.663342e-18, 
    1.588365e-18, 1.488312e-18, 1.339947e-18, 1.297808e-18, 1.265664e-18, 
    1.329685e-18, 1.372561e-18, 1.394841e-18, 1.409629e-18, 1.535438e-18, 
    1.579933e-18, 1.571549e-18, 1.700445e-18, 1.741679e-18, 1.809356e-18, 
    1.867685e-18, 1.942781e-18, 1.958211e-18, 1.936998e-18,
  2.254025e-18, 2.340263e-18, 2.300781e-18, 2.472096e-18, 2.233653e-18, 
    1.993895e-18, 2.124191e-18, 1.997922e-18, 2.016187e-18, 1.884663e-18, 
    1.718078e-18, 1.598761e-18, 1.485849e-18, 1.450272e-18, 1.38919e-18, 
    1.354577e-18, 1.410564e-18, 1.436808e-18, 1.482563e-18, 1.607155e-18, 
    1.667475e-18, 1.866273e-18, 1.991495e-18, 2.100921e-18, 2.027615e-18, 
    2.000152e-18, 2.083874e-18, 2.157436e-18, 2.199004e-18,
  1.910091e-18, 1.892556e-18, 1.843853e-18, 1.932534e-18, 2.045345e-18, 
    1.830165e-18, 1.876093e-18, 1.864876e-18, 1.891418e-18, 1.751256e-18, 
    1.623613e-18, 1.471139e-18, 1.405307e-18, 1.305212e-18, 1.30293e-18, 
    1.273433e-18, 1.314838e-18, 1.250777e-18, 1.34168e-18, 1.398566e-18, 
    1.431248e-18, 1.564259e-18, 1.691422e-18, 1.688176e-18, 1.589839e-18, 
    1.636006e-18, 1.650379e-18, 1.731339e-18, 1.819367e-18,
  1.124006e-18, 1.214729e-18, 1.190516e-18, 1.216969e-18, 1.241422e-18, 
    1.229622e-18, 1.176128e-18, 1.201278e-18, 1.240727e-18, 1.234497e-18, 
    1.188991e-18, 1.157493e-18, 1.099372e-18, 1.082613e-18, 1.016631e-18, 
    9.708385e-19, 9.517844e-19, 9.624285e-19, 9.513399e-19, 9.943577e-19, 
    9.969322e-19, 1.011609e-18, 9.903212e-19, 1.052326e-18, 1.011325e-18, 
    9.774881e-19, 9.90129e-19, 1.00032e-18, 1.084322e-18,
  5.714814e-19, 5.740148e-19, 5.678875e-19, 5.687421e-19, 5.889092e-19, 
    6.171778e-19, 6.18418e-19, 6.292414e-19, 6.113904e-19, 6.195642e-19, 
    6.188271e-19, 6.099353e-19, 6.418947e-19, 6.675075e-19, 6.69934e-19, 
    6.485724e-19, 6.586832e-19, 6.393117e-19, 6.272148e-19, 6.200668e-19, 
    6.017179e-19, 5.800767e-19, 5.824525e-19, 5.902714e-19, 5.918825e-19, 
    5.957305e-19, 5.857419e-19, 5.792533e-19, 5.69676e-19,
  3.33498e-19, 3.282898e-19, 3.323145e-19, 3.375877e-19, 3.53432e-19, 
    3.256791e-19, 3.304914e-19, 3.275893e-19, 3.097313e-19, 3.045691e-19, 
    3.124289e-19, 3.194567e-19, 3.380362e-19, 3.501267e-19, 3.548766e-19, 
    3.599535e-19, 3.581268e-19, 3.570578e-19, 3.650124e-19, 3.758646e-19, 
    3.672109e-19, 3.64748e-19, 3.589337e-19, 3.668835e-19, 3.81445e-19, 
    3.925614e-19, 3.750466e-19, 3.69311e-19, 3.628528e-19,
  2.373749e-19, 2.325169e-19, 2.34159e-19, 2.368427e-19, 2.375816e-19, 
    2.305828e-19, 2.276798e-19, 2.230612e-19, 2.127191e-19, 2.003248e-19, 
    2.021949e-19, 1.928761e-19, 1.886081e-19, 1.879712e-19, 1.856532e-19, 
    1.883481e-19, 1.881563e-19, 1.842456e-19, 1.806791e-19, 1.811443e-19, 
    1.792848e-19, 1.799122e-19, 1.833879e-19, 1.879286e-19, 2.01725e-19, 
    2.115259e-19, 2.279945e-19, 2.344891e-19, 2.367071e-19,
  1.529449e-19, 1.65292e-19, 1.689644e-19, 1.78333e-19, 1.838897e-19, 
    1.767373e-19, 1.752229e-19, 1.726593e-19, 1.717012e-19, 1.691492e-19, 
    1.676185e-19, 1.643526e-19, 1.546848e-19, 1.423153e-19, 1.432375e-19, 
    1.311745e-19, 1.225036e-19, 1.159216e-19, 1.141783e-19, 1.079945e-19, 
    1.026344e-19, 1.001708e-19, 9.785487e-20, 1.033884e-19, 1.078638e-19, 
    1.160255e-19, 1.210624e-19, 1.304348e-19, 1.386956e-19,
  9.454434e-20, 1.011526e-19, 1.087208e-19, 1.181045e-19, 1.237857e-19, 
    1.331372e-19, 1.312209e-19, 1.315192e-19, 1.342567e-19, 1.319524e-19, 
    1.25826e-19, 1.208904e-19, 1.177443e-19, 1.152348e-19, 1.077108e-19, 
    1.024004e-19, 9.895595e-20, 9.693264e-20, 9.163443e-20, 8.636474e-20, 
    8.627093e-20, 8.400422e-20, 8.466875e-20, 8.279168e-20, 8.304315e-20, 
    8.361411e-20, 8.158932e-20, 8.349756e-20, 8.830607e-20,
  7.049846e-20, 7.507717e-20, 7.990289e-20, 8.293483e-20, 8.503609e-20, 
    8.550144e-20, 8.58254e-20, 8.724467e-20, 8.958452e-20, 8.875779e-20, 
    8.735089e-20, 8.667962e-20, 8.652562e-20, 8.495816e-20, 8.239288e-20, 
    7.949362e-20, 7.647031e-20, 7.308275e-20, 7.057199e-20, 6.871842e-20, 
    6.725071e-20, 6.602716e-20, 6.711956e-20, 6.738065e-20, 6.856526e-20, 
    6.992131e-20, 6.818808e-20, 6.797335e-20, 6.881146e-20,
  1.185919e-20, 1.185919e-20, 1.185919e-20, 1.185919e-20, 1.185919e-20, 
    1.185919e-20, 1.185919e-20, 1.208638e-20, 1.208638e-20, 1.208638e-20, 
    1.208638e-20, 1.208638e-20, 1.208638e-20, 1.208638e-20, 1.152267e-20, 
    1.152267e-20, 1.152267e-20, 1.152267e-20, 1.152267e-20, 1.152267e-20, 
    1.152267e-20, 1.135162e-20, 1.135162e-20, 1.135162e-20, 1.135162e-20, 
    1.135162e-20, 1.135162e-20, 1.135162e-20, 1.185919e-20,
  2.707962e-20, 2.905326e-20, 2.980403e-20, 2.988591e-20, 3.159022e-20, 
    3.214779e-20, 3.280329e-20, 3.290715e-20, 3.338785e-20, 3.369146e-20, 
    3.434866e-20, 3.322639e-20, 3.195334e-20, 3.130187e-20, 3.001608e-20, 
    2.786248e-20, 2.549224e-20, 2.259379e-20, 1.954434e-20, 1.735624e-20, 
    1.583031e-20, 1.578698e-20, 1.610511e-20, 1.658809e-20, 1.698009e-20, 
    1.857542e-20, 2.036513e-20, 2.287169e-20, 2.604007e-20,
  1.23809e-19, 1.293425e-19, 1.32349e-19, 1.36319e-19, 1.371649e-19, 
    1.355689e-19, 1.319779e-19, 1.26972e-19, 1.222209e-19, 1.173505e-19, 
    1.092137e-19, 1.02436e-19, 1.020149e-19, 1.002714e-19, 9.679182e-20, 
    9.29953e-20, 8.591047e-20, 7.664754e-20, 6.918082e-20, 6.226031e-20, 
    5.651796e-20, 5.326771e-20, 5.453421e-20, 6.155005e-20, 7.787226e-20, 
    9.392817e-20, 1.015409e-19, 1.088599e-19, 1.173068e-19,
  4.609579e-19, 4.644202e-19, 4.613056e-19, 4.415146e-19, 3.995059e-19, 
    3.631393e-19, 3.329895e-19, 3.19562e-19, 3.008677e-19, 2.978356e-19, 
    3.017658e-19, 2.935436e-19, 2.851914e-19, 2.713931e-19, 2.58183e-19, 
    2.445813e-19, 2.310291e-19, 2.13177e-19, 2.093895e-19, 2.188581e-19, 
    2.344673e-19, 2.626575e-19, 2.841175e-19, 3.097684e-19, 3.36386e-19, 
    3.756469e-19, 4.011706e-19, 4.360166e-19, 4.573192e-19,
  8.620944e-19, 8.234886e-19, 8.071626e-19, 7.895268e-19, 8.046996e-19, 
    8.30295e-19, 8.27618e-19, 8.32158e-19, 8.435626e-19, 8.338157e-19, 
    8.713345e-19, 8.74859e-19, 8.753936e-19, 8.793461e-19, 9.143705e-19, 
    9.005902e-19, 8.41627e-19, 8.193221e-19, 8.349696e-19, 8.248268e-19, 
    8.47791e-19, 8.371562e-19, 8.353733e-19, 8.192377e-19, 8.5443e-19, 
    8.75559e-19, 8.57255e-19, 8.264584e-19, 8.515639e-19,
  2.220719e-18, 2.253939e-18, 2.255894e-18, 2.166642e-18, 2.147533e-18, 
    2.087051e-18, 2.045625e-18, 2.07671e-18, 2.028562e-18, 2.105859e-18, 
    2.058137e-18, 2.070441e-18, 2.048906e-18, 2.065468e-18, 2.073347e-18, 
    2.069909e-18, 2.038022e-18, 2.03833e-18, 2.072334e-18, 2.08255e-18, 
    2.016392e-18, 2.031872e-18, 2.072792e-18, 2.086386e-18, 2.07855e-18, 
    2.10674e-18, 2.212336e-18, 2.264133e-18, 2.296892e-18,
  3.504275e-18, 3.513177e-18, 3.438844e-18, 3.394736e-18, 3.351176e-18, 
    3.308358e-18, 3.389212e-18, 3.233967e-18, 3.15889e-18, 3.051358e-18, 
    3.018303e-18, 2.91569e-18, 2.989164e-18, 2.983739e-18, 3.006068e-18, 
    2.983992e-18, 3.022316e-18, 3.08781e-18, 2.973029e-18, 3.002232e-18, 
    3.021137e-18, 3.01642e-18, 3.013112e-18, 3.022437e-18, 3.098948e-18, 
    3.289958e-18, 3.335777e-18, 3.319996e-18, 3.42475e-18,
  5.590849e-18, 5.55269e-18, 5.668937e-18, 6.042864e-18, 6.055307e-18, 
    6.106279e-18, 6.128899e-18, 6.092841e-18, 5.860204e-18, 5.665532e-18, 
    5.668252e-18, 4.966193e-18, 4.82342e-18, 4.788701e-18, 4.624032e-18, 
    4.319714e-18, 4.375419e-18, 4.200488e-18, 4.238741e-18, 4.363111e-18, 
    4.645226e-18, 4.714267e-18, 4.937322e-18, 5.179848e-18, 5.213051e-18, 
    5.587021e-18, 5.482319e-18, 5.418035e-18, 5.515932e-18,
  8.371234e-18, 8.793145e-18, 8.761938e-18, 8.608266e-18, 8.422631e-18, 
    8.155201e-18, 8.145283e-18, 8.345602e-18, 8.073777e-18, 7.772584e-18, 
    7.533275e-18, 7.30093e-18, 6.684877e-18, 6.355826e-18, 6.049754e-18, 
    5.872622e-18, 5.770742e-18, 5.846888e-18, 6.287328e-18, 6.823553e-18, 
    6.958977e-18, 7.44261e-18, 7.892287e-18, 8.256529e-18, 8.522762e-18, 
    8.32479e-18, 8.740065e-18, 7.986353e-18, 8.419408e-18,
  8.751752e-18, 8.873683e-18, 9.164531e-18, 9.489986e-18, 9.380382e-18, 
    8.881326e-18, 8.75369e-18, 9.132705e-18, 8.771671e-18, 8.515462e-18, 
    7.891765e-18, 7.294376e-18, 6.857647e-18, 6.370113e-18, 6.316319e-18, 
    6.398892e-18, 6.246027e-18, 6.275202e-18, 6.479502e-18, 7.105089e-18, 
    7.412745e-18, 7.85932e-18, 8.561985e-18, 8.700535e-18, 8.352943e-18, 
    8.270181e-18, 8.687162e-18, 8.384117e-18, 8.683482e-18,
  7.191244e-18, 6.986222e-18, 7.616118e-18, 7.86035e-18, 7.882755e-18, 
    7.414226e-18, 7.990207e-18, 7.990461e-18, 7.859966e-18, 7.792495e-18, 
    7.218109e-18, 6.811194e-18, 6.23609e-18, 5.992788e-18, 5.66366e-18, 
    5.566447e-18, 5.512399e-18, 5.635751e-18, 5.804163e-18, 6.01425e-18, 
    6.308238e-18, 6.79403e-18, 6.848035e-18, 7.131796e-18, 7.328849e-18, 
    7.207631e-18, 7.137037e-18, 7.164227e-18, 7.047129e-18,
  4.782836e-18, 4.813305e-18, 4.735694e-18, 4.769134e-18, 4.900859e-18, 
    4.900398e-18, 4.64675e-18, 4.620817e-18, 4.737683e-18, 4.833437e-18, 
    4.995046e-18, 4.883178e-18, 4.776741e-18, 4.520365e-18, 4.426598e-18, 
    4.374325e-18, 4.202566e-18, 4.065589e-18, 4.087422e-18, 4.202438e-18, 
    4.182047e-18, 4.24604e-18, 4.246617e-18, 4.200805e-18, 4.348669e-18, 
    4.420393e-18, 4.355143e-18, 4.490684e-18, 4.567121e-18,
  2.555731e-18, 2.656728e-18, 2.636204e-18, 2.742888e-18, 2.73926e-18, 
    2.733799e-18, 2.62188e-18, 2.654622e-18, 2.542771e-18, 2.40005e-18, 
    2.437376e-18, 2.583454e-18, 2.825939e-18, 2.952761e-18, 2.860488e-18, 
    2.745602e-18, 2.715331e-18, 2.672581e-18, 2.654126e-18, 2.693531e-18, 
    2.655976e-18, 2.690813e-18, 2.730797e-18, 2.701066e-18, 2.64072e-18, 
    2.748501e-18, 2.662758e-18, 2.538994e-18, 2.550945e-18,
  1.624111e-18, 1.645151e-18, 1.736122e-18, 1.775624e-18, 1.775097e-18, 
    1.735036e-18, 1.732962e-18, 1.683789e-18, 1.623182e-18, 1.545376e-18, 
    1.60216e-18, 1.52529e-18, 1.542921e-18, 1.504336e-18, 1.465288e-18, 
    1.468299e-18, 1.480683e-18, 1.428695e-18, 1.452159e-18, 1.490037e-18, 
    1.525317e-18, 1.575456e-18, 1.590679e-18, 1.692172e-18, 1.75986e-18, 
    1.809442e-18, 1.735127e-18, 1.695839e-18, 1.673556e-18,
  1.040316e-18, 1.07455e-18, 1.108352e-18, 1.206379e-18, 1.276653e-18, 
    1.215275e-18, 1.216359e-18, 1.224965e-18, 1.206288e-18, 1.09284e-18, 
    1.116806e-18, 1.148394e-18, 9.751913e-19, 8.873719e-19, 8.621195e-19, 
    8.183905e-19, 8.018185e-19, 7.922155e-19, 7.473181e-19, 7.157828e-19, 
    7.042099e-19, 7.296942e-19, 7.438525e-19, 7.768757e-19, 8.506742e-19, 
    8.795363e-19, 9.589968e-19, 1.021083e-18, 1.056169e-18,
  5.343008e-19, 5.902574e-19, 6.340668e-19, 6.661261e-19, 7.399694e-19, 
    7.268791e-19, 7.416042e-19, 7.577694e-19, 7.891242e-19, 8.198663e-19, 
    8.219861e-19, 8.011135e-19, 7.937513e-19, 6.848651e-19, 6.530885e-19, 
    6.062458e-19, 5.479265e-19, 4.925101e-19, 4.840998e-19, 4.574231e-19, 
    4.4381e-19, 4.259706e-19, 4.281715e-19, 4.358963e-19, 4.298682e-19, 
    4.51201e-19, 4.466847e-19, 4.642206e-19, 5.096833e-19,
  2.844974e-19, 2.975986e-19, 3.240214e-19, 3.81569e-19, 4.112748e-19, 
    4.475874e-19, 4.562926e-19, 4.704515e-19, 4.786623e-19, 5.094932e-19, 
    5.181861e-19, 5.165314e-19, 5.116919e-19, 4.83201e-19, 4.527447e-19, 
    4.284883e-19, 4.036346e-19, 3.952462e-19, 3.704336e-19, 3.341393e-19, 
    3.076546e-19, 2.965337e-19, 2.972282e-19, 2.912745e-19, 2.842698e-19, 
    2.835105e-19, 2.841933e-19, 2.8985e-19, 2.866417e-19,
  2.139712e-19, 2.177625e-19, 2.27246e-19, 2.322934e-19, 2.335477e-19, 
    2.437643e-19, 2.585626e-19, 2.632354e-19, 2.683956e-19, 2.713639e-19, 
    2.729648e-19, 2.733534e-19, 2.791158e-19, 2.819586e-19, 2.783923e-19, 
    2.70201e-19, 2.608449e-19, 2.503838e-19, 2.458972e-19, 2.336908e-19, 
    2.240074e-19, 2.199597e-19, 2.136146e-19, 2.094429e-19, 2.116189e-19, 
    2.119441e-19, 2.091216e-19, 2.081945e-19, 2.120859e-19,
  3.511195e-20, 3.511195e-20, 3.511195e-20, 3.511195e-20, 3.511195e-20, 
    3.511195e-20, 3.511195e-20, 3.683615e-20, 3.683615e-20, 3.683615e-20, 
    3.683615e-20, 3.683615e-20, 3.683615e-20, 3.683615e-20, 3.553514e-20, 
    3.553514e-20, 3.553514e-20, 3.553514e-20, 3.553514e-20, 3.553514e-20, 
    3.553514e-20, 3.405742e-20, 3.405742e-20, 3.405742e-20, 3.405742e-20, 
    3.405742e-20, 3.405742e-20, 3.405742e-20, 3.511195e-20,
  6.797557e-20, 7.752918e-20, 8.378107e-20, 8.648182e-20, 9.250627e-20, 
    9.281318e-20, 9.435022e-20, 9.497133e-20, 9.680672e-20, 1.004698e-19, 
    1.030624e-19, 9.921878e-20, 9.85607e-20, 9.913604e-20, 9.586824e-20, 
    9.193446e-20, 8.376938e-20, 7.32414e-20, 5.973088e-20, 5.029052e-20, 
    4.29404e-20, 3.910392e-20, 3.924608e-20, 4.001912e-20, 4.221015e-20, 
    4.633971e-20, 4.886731e-20, 5.354411e-20, 6.378665e-20,
  3.143575e-19, 3.416411e-19, 3.676746e-19, 3.902803e-19, 3.935601e-19, 
    4.007468e-19, 4.095146e-19, 4.070865e-19, 4.116053e-19, 4.159644e-19, 
    4.099406e-19, 4.019576e-19, 3.977015e-19, 3.872939e-19, 3.781921e-19, 
    3.607969e-19, 3.359845e-19, 3.023034e-19, 2.712356e-19, 2.360612e-19, 
    2.075646e-19, 1.784793e-19, 1.666308e-19, 1.570074e-19, 1.728923e-19, 
    2.121524e-19, 2.560324e-19, 2.942486e-19, 3.02108e-19,
  1.931975e-18, 2.000229e-18, 2.041798e-18, 2.054761e-18, 2.003897e-18, 
    1.984425e-18, 1.926371e-18, 1.863756e-18, 1.803289e-18, 1.786591e-18, 
    1.772779e-18, 1.748262e-18, 1.724747e-18, 1.661309e-18, 1.573988e-18, 
    1.437506e-18, 1.292576e-18, 1.16149e-18, 1.040891e-18, 9.369812e-19, 
    8.759952e-19, 9.330191e-19, 1.098688e-18, 1.282426e-18, 1.395052e-18, 
    1.53774e-18, 1.663187e-18, 1.762999e-18, 1.871792e-18,
  5.409764e-18, 5.251639e-18, 5.015069e-18, 4.732593e-18, 4.62965e-18, 
    4.744715e-18, 4.713624e-18, 4.827051e-18, 4.94733e-18, 5.154155e-18, 
    5.127374e-18, 5.175868e-18, 5.299192e-18, 5.043778e-18, 4.929783e-18, 
    4.934343e-18, 4.782016e-18, 4.607948e-18, 4.58407e-18, 4.583882e-18, 
    4.612211e-18, 4.582867e-18, 4.721586e-18, 4.776076e-18, 4.977466e-18, 
    5.113132e-18, 5.384005e-18, 5.491616e-18, 5.322937e-18,
  1.24427e-17, 1.24934e-17, 1.248227e-17, 1.193303e-17, 1.180164e-17, 
    1.187915e-17, 1.157738e-17, 1.140837e-17, 1.142231e-17, 1.198432e-17, 
    1.186393e-17, 1.184219e-17, 1.200309e-17, 1.185566e-17, 1.1503e-17, 
    1.151193e-17, 1.178456e-17, 1.191645e-17, 1.176074e-17, 1.164456e-17, 
    1.150339e-17, 1.164974e-17, 1.131296e-17, 1.121586e-17, 1.162394e-17, 
    1.22188e-17, 1.264471e-17, 1.26317e-17, 1.264873e-17,
  2.17654e-17, 2.181623e-17, 2.045369e-17, 2.040588e-17, 2.006994e-17, 
    1.9887e-17, 2.004497e-17, 1.931473e-17, 1.936159e-17, 1.813606e-17, 
    1.810552e-17, 1.77748e-17, 1.752155e-17, 1.717151e-17, 1.708641e-17, 
    1.795748e-17, 1.845197e-17, 1.872323e-17, 1.898065e-17, 1.87574e-17, 
    1.907719e-17, 1.922524e-17, 1.996936e-17, 2.025369e-17, 2.078483e-17, 
    2.195817e-17, 2.147813e-17, 2.184054e-17, 2.155031e-17,
  2.992028e-17, 3.087789e-17, 3.242845e-17, 3.245987e-17, 3.365187e-17, 
    3.378062e-17, 3.339795e-17, 3.33327e-17, 3.118843e-17, 2.953351e-17, 
    2.868219e-17, 2.862649e-17, 2.794173e-17, 2.700943e-17, 2.618747e-17, 
    2.484223e-17, 2.39596e-17, 2.369959e-17, 2.426419e-17, 2.438779e-17, 
    2.5471e-17, 2.635045e-17, 2.721679e-17, 2.794006e-17, 2.999269e-17, 
    2.924454e-17, 2.969888e-17, 2.915113e-17, 2.969686e-17,
  4.579302e-17, 4.907349e-17, 4.769741e-17, 5.007499e-17, 4.84023e-17, 
    4.465835e-17, 4.531215e-17, 4.659883e-17, 4.650991e-17, 4.385449e-17, 
    4.13788e-17, 3.92741e-17, 3.671814e-17, 3.445082e-17, 3.47252e-17, 
    3.255161e-17, 3.111898e-17, 3.154369e-17, 3.353046e-17, 3.419613e-17, 
    3.629479e-17, 3.939554e-17, 4.22603e-17, 4.515493e-17, 4.897993e-17, 
    4.973815e-17, 4.967481e-17, 4.762845e-17, 4.521251e-17,
  4.901516e-17, 5.07387e-17, 5.161308e-17, 5.078571e-17, 4.93307e-17, 
    4.659961e-17, 4.736826e-17, 4.745489e-17, 4.675777e-17, 4.407051e-17, 
    4.156648e-17, 3.812498e-17, 3.487822e-17, 3.281984e-17, 3.168664e-17, 
    3.219192e-17, 3.210463e-17, 3.241331e-17, 3.129476e-17, 3.301757e-17, 
    3.545295e-17, 3.826343e-17, 4.070946e-17, 4.423764e-17, 4.49985e-17, 
    4.607659e-17, 4.76962e-17, 5.013882e-17, 4.908901e-17,
  3.841225e-17, 3.901256e-17, 4.011534e-17, 3.92935e-17, 3.976606e-17, 
    4.145306e-17, 4.05373e-17, 4.032028e-17, 3.784544e-17, 3.750618e-17, 
    3.741166e-17, 3.580617e-17, 3.427108e-17, 3.243082e-17, 2.977588e-17, 
    2.92728e-17, 2.868005e-17, 3.03553e-17, 3.186147e-17, 3.153355e-17, 
    3.200667e-17, 3.360213e-17, 3.530622e-17, 3.800624e-17, 4.00453e-17, 
    3.976487e-17, 3.817089e-17, 3.837397e-17, 3.825952e-17,
  2.596551e-17, 2.5629e-17, 2.734861e-17, 2.632042e-17, 2.536915e-17, 
    2.539952e-17, 2.501211e-17, 2.44642e-17, 2.420559e-17, 2.45737e-17, 
    2.6136e-17, 2.636699e-17, 2.669792e-17, 2.626331e-17, 2.506233e-17, 
    2.388114e-17, 2.303261e-17, 2.295144e-17, 2.276558e-17, 2.259383e-17, 
    2.272624e-17, 2.295296e-17, 2.391477e-17, 2.486356e-17, 2.697058e-17, 
    2.756905e-17, 2.69919e-17, 2.752812e-17, 2.619525e-17,
  1.763806e-17, 1.836953e-17, 1.788345e-17, 1.751669e-17, 1.583388e-17, 
    1.546035e-17, 1.504235e-17, 1.49463e-17, 1.485683e-17, 1.462354e-17, 
    1.457358e-17, 1.469364e-17, 1.526888e-17, 1.54737e-17, 1.543711e-17, 
    1.549628e-17, 1.575084e-17, 1.558216e-17, 1.552429e-17, 1.581544e-17, 
    1.607875e-17, 1.591936e-17, 1.629411e-17, 1.636267e-17, 1.677824e-17, 
    1.686026e-17, 1.665941e-17, 1.66669e-17, 1.709478e-17,
  1.075961e-17, 1.126461e-17, 1.149439e-17, 1.294e-17, 1.357698e-17, 
    1.359848e-17, 1.283007e-17, 1.198098e-17, 1.105696e-17, 1.076089e-17, 
    1.087548e-17, 1.096748e-17, 9.728329e-18, 9.195036e-18, 8.668625e-18, 
    8.195157e-18, 7.590612e-18, 7.214573e-18, 7.359808e-18, 7.575321e-18, 
    8.159854e-18, 8.650262e-18, 9.118574e-18, 9.731259e-18, 9.819119e-18, 
    1.010037e-17, 1.020618e-17, 1.035297e-17, 1.023836e-17,
  5.570154e-18, 6.115842e-18, 6.338269e-18, 6.906305e-18, 7.340127e-18, 
    7.566139e-18, 7.987394e-18, 7.911199e-18, 7.661679e-18, 7.561585e-18, 
    7.482547e-18, 7.478302e-18, 6.576801e-18, 5.655201e-18, 4.956855e-18, 
    4.392662e-18, 4.136179e-18, 4.1461e-18, 3.917383e-18, 3.728755e-18, 
    3.670991e-18, 3.603911e-18, 3.54548e-18, 3.651218e-18, 3.874512e-18, 
    4.294314e-18, 4.562688e-18, 5.080024e-18, 5.023535e-18,
  2.228575e-18, 2.465187e-18, 2.681833e-18, 2.864751e-18, 3.024048e-18, 
    3.379841e-18, 3.636619e-18, 3.787482e-18, 4.043055e-18, 4.334695e-18, 
    4.481796e-18, 4.861036e-18, 4.491108e-18, 3.748696e-18, 3.509963e-18, 
    3.253538e-18, 2.953484e-18, 2.628202e-18, 2.304785e-18, 2.171787e-18, 
    2.11838e-18, 2.093148e-18, 2.121602e-18, 2.082383e-18, 2.216352e-18, 
    2.181398e-18, 2.209532e-18, 2.128496e-18, 2.181839e-18,
  1.153643e-18, 1.096513e-18, 1.139061e-18, 1.246044e-18, 1.398708e-18, 
    1.495194e-18, 1.721032e-18, 1.876284e-18, 2.010334e-18, 2.247719e-18, 
    2.564489e-18, 2.686642e-18, 2.427991e-18, 2.219133e-18, 2.140839e-18, 
    1.997507e-18, 1.809255e-18, 1.734248e-18, 1.562466e-18, 1.399607e-18, 
    1.350433e-18, 1.331118e-18, 1.382904e-18, 1.460029e-18, 1.436156e-18, 
    1.329343e-18, 1.287482e-18, 1.228867e-18, 1.223722e-18,
  8.173409e-19, 7.569217e-19, 7.393803e-19, 7.786027e-19, 8.207501e-19, 
    8.535274e-19, 8.759789e-19, 9.590726e-19, 1.130395e-18, 1.203365e-18, 
    1.271137e-18, 1.309013e-18, 1.261052e-18, 1.202222e-18, 1.217919e-18, 
    1.223441e-18, 1.163123e-18, 1.137518e-18, 1.119388e-18, 1.083398e-18, 
    1.098676e-18, 1.118872e-18, 1.099868e-18, 1.083335e-18, 1.045709e-18, 
    1.008321e-18, 9.4416e-19, 9.070591e-19, 8.487973e-19,
  1.002282e-19, 1.002282e-19, 1.002282e-19, 1.002282e-19, 1.002282e-19, 
    1.002282e-19, 1.002282e-19, 1.038349e-19, 1.038349e-19, 1.038349e-19, 
    1.038349e-19, 1.038349e-19, 1.038349e-19, 1.038349e-19, 9.979833e-20, 
    9.979833e-20, 9.979833e-20, 9.979833e-20, 9.979833e-20, 9.979833e-20, 
    9.979833e-20, 9.68647e-20, 9.68647e-20, 9.68647e-20, 9.68647e-20, 
    9.68647e-20, 9.68647e-20, 9.68647e-20, 1.002282e-19,
  1.787181e-19, 1.90655e-19, 2.029319e-19, 2.116916e-19, 2.278889e-19, 
    2.399766e-19, 2.483835e-19, 2.534163e-19, 2.552579e-19, 2.601388e-19, 
    2.701329e-19, 2.665497e-19, 2.620147e-19, 2.556897e-19, 2.414795e-19, 
    2.148033e-19, 1.942782e-19, 1.792368e-19, 1.428272e-19, 1.177183e-19, 
    1.02743e-19, 9.457519e-20, 9.3296e-20, 9.443759e-20, 9.79789e-20, 
    1.057609e-19, 1.20107e-19, 1.41197e-19, 1.681359e-19,
  7.474381e-19, 8.543573e-19, 8.867539e-19, 9.42779e-19, 9.711431e-19, 
    1.010841e-18, 1.007622e-18, 1.036529e-18, 1.004369e-18, 1.007008e-18, 
    1.001767e-18, 9.670778e-19, 9.872503e-19, 9.782181e-19, 8.880396e-19, 
    7.882312e-19, 6.951572e-19, 5.862244e-19, 4.986947e-19, 4.049522e-19, 
    3.380558e-19, 2.758617e-19, 2.53276e-19, 2.537437e-19, 2.810835e-19, 
    3.115427e-19, 4.047148e-19, 5.190901e-19, 6.674272e-19,
  7.05767e-18, 6.865743e-18, 6.895692e-18, 7.073624e-18, 7.120801e-18, 
    7.528479e-18, 7.884757e-18, 7.975197e-18, 7.774248e-18, 7.828816e-18, 
    7.944573e-18, 7.641832e-18, 7.483757e-18, 7.458564e-18, 7.315677e-18, 
    6.918591e-18, 6.508949e-18, 5.838539e-18, 5.309487e-18, 4.913313e-18, 
    4.580729e-18, 4.402924e-18, 4.256371e-18, 4.518336e-18, 4.906796e-18, 
    5.972919e-18, 6.040646e-18, 6.340463e-18, 7.002252e-18,
  2.522745e-17, 2.564824e-17, 2.565691e-17, 2.497246e-17, 2.387112e-17, 
    2.348214e-17, 2.262568e-17, 2.2567e-17, 2.301787e-17, 2.377452e-17, 
    2.340792e-17, 2.311599e-17, 2.352979e-17, 2.293182e-17, 2.147379e-17, 
    2.075714e-17, 2.021139e-17, 2.054234e-17, 1.989015e-17, 1.952166e-17, 
    1.931147e-17, 1.918556e-17, 2.025008e-17, 2.181582e-17, 2.389161e-17, 
    2.470884e-17, 2.522149e-17, 2.562466e-17, 2.48825e-17,
  5.818827e-17, 6.040543e-17, 5.953148e-17, 5.746726e-17, 5.604416e-17, 
    5.460786e-17, 5.652573e-17, 5.515101e-17, 5.538904e-17, 5.584049e-17, 
    5.555654e-17, 5.517126e-17, 5.779969e-17, 5.611847e-17, 5.274214e-17, 
    5.311796e-17, 5.333353e-17, 5.336407e-17, 5.366745e-17, 5.302874e-17, 
    5.185632e-17, 5.497657e-17, 5.373011e-17, 5.346694e-17, 5.451881e-17, 
    5.724848e-17, 5.948534e-17, 5.855041e-17, 5.918952e-17,
  1.050475e-16, 1.079909e-16, 1.072426e-16, 1.040219e-16, 1.050629e-16, 
    1.070188e-16, 1.03721e-16, 9.964944e-17, 9.849265e-17, 9.619308e-17, 
    9.201715e-17, 9.433633e-17, 9.1727e-17, 9.263653e-17, 9.252601e-17, 
    9.56301e-17, 9.382949e-17, 9.407627e-17, 9.339736e-17, 9.66998e-17, 
    9.776565e-17, 1.012007e-16, 1.047618e-16, 1.062747e-16, 1.070339e-16, 
    1.089481e-16, 1.07695e-16, 1.107202e-16, 1.08251e-16,
  1.577338e-16, 1.57275e-16, 1.642038e-16, 1.763859e-16, 1.674907e-16, 
    1.701167e-16, 1.739851e-16, 1.625828e-16, 1.599175e-16, 1.533318e-16, 
    1.457194e-16, 1.403314e-16, 1.384926e-16, 1.331095e-16, 1.255588e-16, 
    1.244191e-16, 1.248526e-16, 1.238922e-16, 1.26184e-16, 1.266479e-16, 
    1.282564e-16, 1.315413e-16, 1.406314e-16, 1.425265e-16, 1.53392e-16, 
    1.519852e-16, 1.468261e-16, 1.449558e-16, 1.528949e-16,
  2.337489e-16, 2.305018e-16, 2.271799e-16, 2.294833e-16, 2.33884e-16, 
    2.233753e-16, 2.144345e-16, 2.197559e-16, 2.267011e-16, 2.219472e-16, 
    2.037647e-16, 1.933847e-16, 1.748809e-16, 1.636865e-16, 1.583669e-16, 
    1.509087e-16, 1.437523e-16, 1.484833e-16, 1.509136e-16, 1.539241e-16, 
    1.619214e-16, 1.689838e-16, 1.842126e-16, 1.96836e-16, 2.123825e-16, 
    2.291791e-16, 2.348728e-16, 2.323398e-16, 2.340552e-16,
  2.303209e-16, 2.369914e-16, 2.343313e-16, 2.329797e-16, 2.272818e-16, 
    2.236026e-16, 2.221412e-16, 2.179102e-16, 2.137185e-16, 2.020381e-16, 
    1.881746e-16, 1.763663e-16, 1.650083e-16, 1.615434e-16, 1.484234e-16, 
    1.461074e-16, 1.474421e-16, 1.466636e-16, 1.348461e-16, 1.412657e-16, 
    1.534155e-16, 1.575657e-16, 1.606562e-16, 1.715291e-16, 1.863898e-16, 
    2.110728e-16, 2.072303e-16, 2.341074e-16, 2.282403e-16,
  1.91857e-16, 1.930086e-16, 1.870693e-16, 1.862712e-16, 1.894879e-16, 
    1.90106e-16, 1.930511e-16, 1.94543e-16, 1.923124e-16, 1.862866e-16, 
    1.779715e-16, 1.70257e-16, 1.622095e-16, 1.572762e-16, 1.503426e-16, 
    1.459911e-16, 1.465384e-16, 1.428106e-16, 1.52401e-16, 1.510638e-16, 
    1.586387e-16, 1.669836e-16, 1.742466e-16, 1.808987e-16, 1.755994e-16, 
    1.797896e-16, 1.807486e-16, 1.834644e-16, 1.861859e-16,
  1.405625e-16, 1.330732e-16, 1.306445e-16, 1.253936e-16, 1.225868e-16, 
    1.179119e-16, 1.180224e-16, 1.183565e-16, 1.224303e-16, 1.257098e-16, 
    1.349186e-16, 1.386409e-16, 1.341256e-16, 1.270205e-16, 1.205991e-16, 
    1.162336e-16, 1.146258e-16, 1.165294e-16, 1.17761e-16, 1.240371e-16, 
    1.304204e-16, 1.404323e-16, 1.397675e-16, 1.455084e-16, 1.511909e-16, 
    1.538049e-16, 1.451007e-16, 1.406604e-16, 1.409135e-16,
  1.092202e-16, 1.237953e-16, 1.200738e-16, 1.103093e-16, 9.954805e-17, 
    9.911594e-17, 9.886324e-17, 1.004614e-16, 9.783024e-17, 9.814669e-17, 
    8.836667e-17, 8.518567e-17, 8.479668e-17, 8.340464e-17, 8.129416e-17, 
    8.038786e-17, 7.830973e-17, 7.575929e-17, 7.33262e-17, 7.503024e-17, 
    7.751864e-17, 7.814905e-17, 8.306782e-17, 9.032575e-17, 9.651931e-17, 
    1.018615e-16, 1.065219e-16, 1.018546e-16, 1.010677e-16,
  7.346155e-17, 8.943609e-17, 9.59219e-17, 9.699192e-17, 9.10943e-17, 
    8.765419e-17, 8.394204e-17, 8.454956e-17, 8.752106e-17, 8.766863e-17, 
    7.266755e-17, 5.978231e-17, 5.190123e-17, 4.878885e-17, 4.284779e-17, 
    3.798538e-17, 3.536903e-17, 3.469026e-17, 3.49248e-17, 3.468209e-17, 
    3.502163e-17, 3.757924e-17, 3.909906e-17, 3.906359e-17, 4.190244e-17, 
    4.92522e-17, 5.213632e-17, 6.138642e-17, 6.522294e-17,
  2.598463e-17, 3.054876e-17, 3.579904e-17, 3.95221e-17, 4.152886e-17, 
    4.097858e-17, 4.083359e-17, 3.9407e-17, 4.492036e-17, 5.057355e-17, 
    4.89191e-17, 3.828033e-17, 3.32015e-17, 3.123013e-17, 2.797835e-17, 
    2.564203e-17, 2.299268e-17, 2.093672e-17, 1.74752e-17, 1.654746e-17, 
    1.671093e-17, 1.581243e-17, 1.663645e-17, 1.654016e-17, 1.743174e-17, 
    1.888076e-17, 2.151642e-17, 2.23832e-17, 2.382386e-17,
  9.20797e-18, 9.500177e-18, 1.007291e-17, 1.070267e-17, 1.129384e-17, 
    1.274601e-17, 1.40876e-17, 1.559745e-17, 1.647875e-17, 1.971639e-17, 
    2.108486e-17, 2.277851e-17, 2.204054e-17, 2.035868e-17, 1.859288e-17, 
    1.717924e-17, 1.586284e-17, 1.408911e-17, 1.162817e-17, 1.022644e-17, 
    9.769758e-18, 9.845888e-18, 1.049531e-17, 1.063253e-17, 1.059545e-17, 
    1.015837e-17, 9.408572e-18, 9.268395e-18, 9.801152e-18,
  4.678007e-18, 4.411665e-18, 4.288983e-18, 4.296142e-18, 3.986972e-18, 
    4.410271e-18, 4.975029e-18, 6.16426e-18, 7.327934e-18, 8.279766e-18, 
    9.156822e-18, 1.031781e-17, 1.139011e-17, 1.078733e-17, 1.040332e-17, 
    1.010505e-17, 9.092928e-18, 8.158592e-18, 7.491661e-18, 6.803963e-18, 
    6.196644e-18, 6.561507e-18, 6.904189e-18, 6.817556e-18, 6.674606e-18, 
    6.388305e-18, 5.83353e-18, 5.454154e-18, 5.003668e-18,
  3.669048e-18, 3.039071e-18, 2.701336e-18, 2.653049e-18, 2.624069e-18, 
    2.765919e-18, 3.030582e-18, 3.307294e-18, 3.924984e-18, 4.416166e-18, 
    4.934792e-18, 5.184756e-18, 5.308342e-18, 5.306932e-18, 5.38463e-18, 
    5.39296e-18, 5.146515e-18, 4.914754e-18, 4.823813e-18, 4.957202e-18, 
    5.204772e-18, 5.314114e-18, 5.426404e-18, 5.295985e-18, 4.853615e-18, 
    4.562157e-18, 4.274747e-18, 4.126534e-18, 3.88501e-18,
  2.568689e-19, 2.568689e-19, 2.568689e-19, 2.568689e-19, 2.568689e-19, 
    2.568689e-19, 2.568689e-19, 2.706009e-19, 2.706009e-19, 2.706009e-19, 
    2.706009e-19, 2.706009e-19, 2.706009e-19, 2.706009e-19, 2.573365e-19, 
    2.573365e-19, 2.573365e-19, 2.573365e-19, 2.573365e-19, 2.573365e-19, 
    2.573365e-19, 2.472184e-19, 2.472184e-19, 2.472184e-19, 2.472184e-19, 
    2.472184e-19, 2.472184e-19, 2.472184e-19, 2.568689e-19,
  3.396632e-19, 4.168067e-19, 4.813706e-19, 5.300602e-19, 5.810034e-19, 
    6.192389e-19, 6.366067e-19, 6.45719e-19, 6.45808e-19, 6.449241e-19, 
    6.675817e-19, 6.677785e-19, 6.639509e-19, 6.46074e-19, 6.031987e-19, 
    5.208753e-19, 4.498272e-19, 4.02687e-19, 3.555542e-19, 2.954102e-19, 
    2.571948e-19, 2.392855e-19, 2.253367e-19, 2.238034e-19, 2.23625e-19, 
    2.226435e-19, 2.402776e-19, 2.657763e-19, 3.135684e-19,
  1.569529e-18, 2.048053e-18, 2.333046e-18, 2.467659e-18, 2.675355e-18, 
    2.591961e-18, 2.521683e-18, 2.510357e-18, 2.482626e-18, 2.481188e-18, 
    2.480499e-18, 2.489184e-18, 2.521743e-18, 2.596769e-18, 2.425935e-18, 
    2.044399e-18, 1.704078e-18, 1.315041e-18, 9.524456e-19, 7.526295e-19, 
    6.147437e-19, 5.033992e-19, 4.463944e-19, 4.029998e-19, 4.517591e-19, 
    5.689755e-19, 7.07211e-19, 9.89891e-19, 1.328208e-18,
  2.254491e-17, 2.232016e-17, 2.175056e-17, 2.11099e-17, 2.082852e-17, 
    2.155038e-17, 2.14974e-17, 2.088472e-17, 2.07409e-17, 2.079409e-17, 
    2.091903e-17, 1.974747e-17, 1.924652e-17, 1.954108e-17, 1.826708e-17, 
    1.691743e-17, 1.666696e-17, 1.42166e-17, 1.216525e-17, 1.213007e-17, 
    1.219534e-17, 1.241935e-17, 1.192378e-17, 1.187557e-17, 1.110399e-17, 
    1.326024e-17, 1.652935e-17, 1.80139e-17, 2.136541e-17,
  8.542387e-17, 8.604148e-17, 8.33578e-17, 8.442921e-17, 8.501324e-17, 
    8.314638e-17, 8.104006e-17, 8.022874e-17, 8.358994e-17, 8.746554e-17, 
    9.086138e-17, 8.932489e-17, 8.977545e-17, 9.026336e-17, 8.996947e-17, 
    8.521053e-17, 8.128067e-17, 7.860881e-17, 7.689616e-17, 7.260596e-17, 
    6.97823e-17, 6.778313e-17, 6.834772e-17, 7.523115e-17, 8.374654e-17, 
    9.382237e-17, 9.532063e-17, 8.755786e-17, 8.403261e-17,
  2.179767e-16, 2.243404e-16, 2.207546e-16, 2.177802e-16, 2.196125e-16, 
    2.139154e-16, 2.157506e-16, 2.092851e-16, 2.217664e-16, 2.211231e-16, 
    2.170214e-16, 2.147264e-16, 2.268503e-16, 2.146308e-16, 2.081762e-16, 
    2.019845e-16, 1.993963e-16, 1.934356e-16, 1.929886e-16, 1.882033e-16, 
    1.796353e-16, 1.930939e-16, 2.010442e-16, 2.05456e-16, 2.117031e-16, 
    2.106177e-16, 2.259031e-16, 2.246265e-16, 2.254891e-16,
  4.058763e-16, 4.107989e-16, 4.270884e-16, 4.28042e-16, 4.363085e-16, 
    4.181141e-16, 4.219474e-16, 4.106671e-16, 3.994076e-16, 3.843722e-16, 
    3.903498e-16, 3.811612e-16, 3.765484e-16, 3.7827e-16, 3.814432e-16, 
    3.849506e-16, 3.835419e-16, 3.73712e-16, 3.88316e-16, 3.902239e-16, 
    3.964357e-16, 4.07294e-16, 4.175738e-16, 4.151292e-16, 4.151427e-16, 
    4.132361e-16, 4.090545e-16, 4.03171e-16, 3.986166e-16,
  7.35418e-16, 7.517271e-16, 7.752885e-16, 7.882499e-16, 8.519834e-16, 
    8.252911e-16, 8.148732e-16, 8.275994e-16, 7.781467e-16, 7.12317e-16, 
    7.19612e-16, 6.947381e-16, 6.412e-16, 6.27293e-16, 6.091021e-16, 
    5.859224e-16, 5.819367e-16, 5.868236e-16, 6.007963e-16, 6.177071e-16, 
    6.469546e-16, 6.648969e-16, 6.700564e-16, 6.983982e-16, 6.955205e-16, 
    6.71398e-16, 6.970119e-16, 6.854741e-16, 6.836909e-16,
  9.926429e-16, 1.028034e-15, 1.047185e-15, 9.831838e-16, 9.822744e-16, 
    9.309856e-16, 9.36201e-16, 9.162767e-16, 9.282747e-16, 9.445043e-16, 
    9.150121e-16, 8.632932e-16, 8.084234e-16, 7.69148e-16, 7.43653e-16, 
    7.300038e-16, 6.986544e-16, 7.018535e-16, 7.319474e-16, 7.280164e-16, 
    7.366264e-16, 7.675425e-16, 8.116617e-16, 8.951731e-16, 9.320893e-16, 
    9.564403e-16, 1.011531e-15, 1.01585e-15, 9.461288e-16,
  9.558013e-16, 9.262232e-16, 9.312004e-16, 9.255713e-16, 9.258863e-16, 
    8.988595e-16, 8.934365e-16, 9.081425e-16, 8.854678e-16, 8.651415e-16, 
    8.610282e-16, 8.617386e-16, 7.927493e-16, 7.479931e-16, 7.117779e-16, 
    7.057023e-16, 6.758104e-16, 6.60907e-16, 6.726848e-16, 6.823153e-16, 
    7.11121e-16, 7.283638e-16, 7.686011e-16, 7.92459e-16, 8.207189e-16, 
    8.861665e-16, 9.698721e-16, 9.826522e-16, 9.333073e-16,
  7.7603e-16, 7.64764e-16, 7.535909e-16, 7.498476e-16, 7.308029e-16, 
    7.373244e-16, 7.637259e-16, 7.827402e-16, 7.727771e-16, 7.790644e-16, 
    7.674476e-16, 7.520417e-16, 7.342196e-16, 7.040154e-16, 6.596534e-16, 
    6.532171e-16, 6.573827e-16, 6.596782e-16, 6.534383e-16, 6.70414e-16, 
    6.771506e-16, 6.994375e-16, 7.279712e-16, 7.972412e-16, 7.857101e-16, 
    7.445907e-16, 7.658447e-16, 7.697622e-16, 7.7435e-16,
  6.383935e-16, 6.11545e-16, 5.762922e-16, 5.635944e-16, 5.757426e-16, 
    5.701348e-16, 5.723998e-16, 5.50402e-16, 5.694728e-16, 5.915165e-16, 
    6.436803e-16, 6.309337e-16, 6.027023e-16, 6.114901e-16, 5.884816e-16, 
    5.965092e-16, 5.823246e-16, 6.018413e-16, 6.144138e-16, 6.227419e-16, 
    6.362222e-16, 6.389936e-16, 6.437971e-16, 6.367291e-16, 6.283401e-16, 
    6.142603e-16, 6.124335e-16, 6.174608e-16, 6.203653e-16,
  5.15208e-16, 6.034217e-16, 5.860226e-16, 5.773838e-16, 5.602019e-16, 
    5.938926e-16, 6.07052e-16, 5.718842e-16, 5.467959e-16, 4.810751e-16, 
    4.177073e-16, 3.566353e-16, 3.707392e-16, 3.689178e-16, 3.539476e-16, 
    3.476981e-16, 3.532567e-16, 3.477831e-16, 3.529057e-16, 4.022285e-16, 
    4.385258e-16, 4.421762e-16, 4.453257e-16, 4.590729e-16, 5.167171e-16, 
    5.105835e-16, 4.746845e-16, 4.815666e-16, 4.79177e-16,
  3.725992e-16, 4.781445e-16, 5.452797e-16, 5.05534e-16, 4.605043e-16, 
    4.677614e-16, 4.793408e-16, 4.866989e-16, 4.817969e-16, 5.131096e-16, 
    3.658234e-16, 2.604026e-16, 2.185173e-16, 1.983585e-16, 1.66874e-16, 
    1.489356e-16, 1.326532e-16, 1.319542e-16, 1.33609e-16, 1.328895e-16, 
    1.307181e-16, 1.369648e-16, 1.47987e-16, 1.773955e-16, 2.128472e-16, 
    2.525568e-16, 2.942936e-16, 3.066887e-16, 3.278923e-16,
  1.435163e-16, 1.660059e-16, 1.839141e-16, 1.951721e-16, 1.839967e-16, 
    1.677755e-16, 1.668243e-16, 1.962075e-16, 2.275148e-16, 2.477294e-16, 
    2.480111e-16, 1.826536e-16, 1.327268e-16, 1.342631e-16, 1.156773e-16, 
    1.008343e-16, 9.333901e-17, 8.80225e-17, 6.931079e-17, 6.261461e-17, 
    6.203898e-17, 6.167835e-17, 6.566883e-17, 6.676229e-17, 6.708363e-17, 
    6.514493e-17, 7.241676e-17, 9.404807e-17, 1.125487e-16,
  3.589236e-17, 3.451385e-17, 3.40748e-17, 3.696046e-17, 3.895963e-17, 
    4.531935e-17, 5.230503e-17, 5.943746e-17, 6.723307e-17, 7.197361e-17, 
    8.771253e-17, 1.030388e-16, 9.937951e-17, 9.685431e-17, 8.556556e-17, 
    8.225137e-17, 7.573607e-17, 6.458201e-17, 5.043492e-17, 4.285414e-17, 
    3.885291e-17, 3.714619e-17, 3.522079e-17, 3.799102e-17, 3.829503e-17, 
    3.655541e-17, 3.661111e-17, 3.789342e-17, 3.756039e-17,
  1.754412e-17, 1.644396e-17, 1.497546e-17, 1.375527e-17, 1.310682e-17, 
    1.29021e-17, 1.493243e-17, 1.903929e-17, 2.564943e-17, 3.04293e-17, 
    3.591587e-17, 4.002013e-17, 5.228462e-17, 5.765312e-17, 5.565111e-17, 
    5.10927e-17, 4.394079e-17, 4.050533e-17, 3.535226e-17, 3.367096e-17, 
    3.004184e-17, 2.979406e-17, 2.833364e-17, 2.666252e-17, 2.367015e-17, 
    2.02044e-17, 1.963905e-17, 2.116785e-17, 1.885104e-17,
  1.585811e-17, 1.509252e-17, 1.349914e-17, 1.175899e-17, 1.070948e-17, 
    1.035633e-17, 9.707199e-18, 9.513434e-18, 1.144084e-17, 1.366111e-17, 
    1.53299e-17, 1.787498e-17, 1.977859e-17, 2.137142e-17, 2.325366e-17, 
    2.294147e-17, 2.275539e-17, 2.233693e-17, 2.240516e-17, 2.180453e-17, 
    2.185863e-17, 2.157142e-17, 2.119238e-17, 2.068237e-17, 2.070009e-17, 
    2.028987e-17, 1.877005e-17, 1.749869e-17, 1.630261e-17,
  6.702528e-19, 6.702528e-19, 6.702528e-19, 6.702528e-19, 6.702528e-19, 
    6.702528e-19, 6.702528e-19, 7.092562e-19, 7.092562e-19, 7.092562e-19, 
    7.092562e-19, 7.092562e-19, 7.092562e-19, 7.092562e-19, 6.940363e-19, 
    6.940363e-19, 6.940363e-19, 6.940363e-19, 6.940363e-19, 6.940363e-19, 
    6.940363e-19, 6.619364e-19, 6.619364e-19, 6.619364e-19, 6.619364e-19, 
    6.619364e-19, 6.619364e-19, 6.619364e-19, 6.702528e-19,
  5.990152e-19, 7.488989e-19, 9.190379e-19, 1.075272e-18, 1.344044e-18, 
    1.510993e-18, 1.706112e-18, 1.791994e-18, 1.706995e-18, 1.686028e-18, 
    1.768838e-18, 1.824302e-18, 1.877213e-18, 1.796105e-18, 1.654267e-18, 
    1.483811e-18, 1.29184e-18, 1.133623e-18, 1.019168e-18, 8.669296e-19, 
    8.111053e-19, 7.791482e-19, 7.031308e-19, 5.816162e-19, 4.836453e-19, 
    4.53621e-19, 4.399653e-19, 4.940621e-19, 5.64729e-19,
  3.444882e-18, 4.711691e-18, 5.68484e-18, 6.371747e-18, 7.053466e-18, 
    7.471624e-18, 7.676013e-18, 6.93578e-18, 6.388622e-18, 6.189855e-18, 
    6.474581e-18, 6.861136e-18, 7.206886e-18, 7.475451e-18, 7.329787e-18, 
    6.022353e-18, 4.64645e-18, 3.453612e-18, 2.421192e-18, 2.069368e-18, 
    1.67268e-18, 1.335845e-18, 1.068971e-18, 8.947437e-19, 8.617712e-19, 
    1.016267e-18, 1.379353e-18, 2.086105e-18, 2.968645e-18,
  5.770714e-17, 5.663296e-17, 5.629766e-17, 5.510467e-17, 5.218701e-17, 
    5.263283e-17, 5.236518e-17, 5.243692e-17, 5.135069e-17, 5.058783e-17, 
    4.965692e-17, 4.942516e-17, 4.826598e-17, 4.806464e-17, 4.288867e-17, 
    3.520184e-17, 3.240461e-17, 2.190853e-17, 1.350323e-17, 1.136646e-17, 
    1.012847e-17, 1.071776e-17, 1.202394e-17, 1.297655e-17, 1.418909e-17, 
    1.643683e-17, 2.706305e-17, 3.879878e-17, 5.216641e-17,
  2.327029e-16, 2.373756e-16, 2.153146e-16, 1.998691e-16, 1.953872e-16, 
    1.988017e-16, 1.984225e-16, 1.891063e-16, 2.017845e-16, 2.095462e-16, 
    2.301559e-16, 2.329993e-16, 2.410639e-16, 2.529587e-16, 2.651569e-16, 
    2.592631e-16, 2.530149e-16, 2.380082e-16, 2.218749e-16, 2.135225e-16, 
    1.953622e-16, 1.871077e-16, 1.789579e-16, 1.989242e-16, 2.063266e-16, 
    2.345729e-16, 2.698529e-16, 2.436593e-16, 2.27775e-16,
  7.68746e-16, 7.684518e-16, 7.54676e-16, 7.534237e-16, 7.734948e-16, 
    7.727958e-16, 7.483991e-16, 7.174753e-16, 7.338672e-16, 6.850489e-16, 
    6.907202e-16, 6.703394e-16, 6.719686e-16, 6.559773e-16, 6.654121e-16, 
    6.3501e-16, 6.100771e-16, 5.8271e-16, 6.013833e-16, 5.937614e-16, 
    5.802224e-16, 5.957243e-16, 6.354104e-16, 6.580188e-16, 7.051304e-16, 
    7.036826e-16, 7.437787e-16, 7.642137e-16, 7.578286e-16,
  1.664905e-15, 1.640784e-15, 1.675716e-15, 1.67248e-15, 1.651287e-15, 
    1.665925e-15, 1.638118e-15, 1.66737e-15, 1.562028e-15, 1.495094e-15, 
    1.483034e-15, 1.427057e-15, 1.39562e-15, 1.42438e-15, 1.45901e-15, 
    1.484415e-15, 1.542521e-15, 1.540091e-15, 1.557885e-15, 1.508072e-15, 
    1.532287e-15, 1.62806e-15, 1.651717e-15, 1.619215e-15, 1.650239e-15, 
    1.680764e-15, 1.646664e-15, 1.626966e-15, 1.639817e-15,
  3.361137e-15, 3.520987e-15, 3.632256e-15, 3.568125e-15, 3.718786e-15, 
    3.655485e-15, 3.488792e-15, 3.504452e-15, 3.481472e-15, 3.357096e-15, 
    3.222782e-15, 3.264201e-15, 3.156913e-15, 3.053262e-15, 3.040533e-15, 
    3.024992e-15, 2.944227e-15, 2.880107e-15, 2.996505e-15, 3.156272e-15, 
    3.216788e-15, 3.446836e-15, 3.421824e-15, 3.511436e-15, 3.479504e-15, 
    3.365954e-15, 3.302174e-15, 3.343838e-15, 3.313333e-15,
  3.935523e-15, 4.056479e-15, 4.249684e-15, 4.313589e-15, 3.989695e-15, 
    4.067771e-15, 3.87782e-15, 3.957812e-15, 3.974848e-15, 4.112383e-15, 
    4.101042e-15, 3.804065e-15, 3.446567e-15, 3.394654e-15, 3.356635e-15, 
    3.253882e-15, 3.051804e-15, 3.065345e-15, 3.161051e-15, 3.327609e-15, 
    3.348342e-15, 3.463568e-15, 3.836418e-15, 3.957134e-15, 3.91075e-15, 
    4.019922e-15, 4.283411e-15, 4.351774e-15, 3.936445e-15,
  3.590385e-15, 3.570606e-15, 3.480707e-15, 3.55463e-15, 3.484526e-15, 
    3.17429e-15, 3.222975e-15, 3.270279e-15, 3.474297e-15, 3.648413e-15, 
    3.593038e-15, 3.234054e-15, 3.094458e-15, 2.872428e-15, 2.789139e-15, 
    2.65765e-15, 2.67526e-15, 2.584522e-15, 2.513315e-15, 2.571384e-15, 
    2.557051e-15, 2.688682e-15, 2.854901e-15, 2.950171e-15, 3.034391e-15, 
    3.281823e-15, 3.562749e-15, 3.619681e-15, 3.575306e-15,
  2.815747e-15, 2.825178e-15, 2.722596e-15, 2.738567e-15, 2.85274e-15, 
    2.8845e-15, 2.96233e-15, 2.921021e-15, 3.032872e-15, 3.069521e-15, 
    3.099092e-15, 2.932191e-15, 2.834294e-15, 2.725047e-15, 2.691401e-15, 
    2.743743e-15, 2.657121e-15, 2.632476e-15, 2.52262e-15, 2.513893e-15, 
    2.536216e-15, 2.658697e-15, 2.583857e-15, 2.76216e-15, 2.84667e-15, 
    2.897715e-15, 2.943833e-15, 2.789999e-15, 2.959669e-15,
  2.581705e-15, 2.502794e-15, 2.688868e-15, 2.785987e-15, 2.754664e-15, 
    2.552297e-15, 2.519783e-15, 2.660483e-15, 2.774949e-15, 2.671898e-15, 
    2.655541e-15, 2.792905e-15, 2.819343e-15, 2.792474e-15, 2.742598e-15, 
    2.792158e-15, 2.85515e-15, 2.929825e-15, 2.918686e-15, 2.838364e-15, 
    2.859136e-15, 2.714401e-15, 2.625899e-15, 2.49984e-15, 2.432891e-15, 
    2.465704e-15, 2.497828e-15, 2.548466e-15, 2.567381e-15,
  1.945481e-15, 2.005683e-15, 2.022625e-15, 2.115585e-15, 2.204957e-15, 
    2.249699e-15, 2.162837e-15, 2.037711e-15, 2.042971e-15, 1.851879e-15, 
    1.603752e-15, 1.421928e-15, 1.496398e-15, 1.538215e-15, 1.687167e-15, 
    1.840256e-15, 1.778504e-15, 1.765043e-15, 1.882301e-15, 2.099293e-15, 
    2.348733e-15, 2.25703e-15, 2.02913e-15, 1.993008e-15, 1.951148e-15, 
    1.932727e-15, 1.950522e-15, 1.898322e-15, 1.887284e-15,
  1.301016e-15, 1.4299e-15, 1.484474e-15, 1.598921e-15, 1.579048e-15, 
    1.479033e-15, 1.487374e-15, 1.451013e-15, 1.518023e-15, 1.632021e-15, 
    1.331905e-15, 1.01012e-15, 7.918966e-16, 7.019453e-16, 5.966777e-16, 
    5.510456e-16, 5.174781e-16, 4.419146e-16, 4.811201e-16, 5.079576e-16, 
    4.869188e-16, 5.177565e-16, 6.774357e-16, 8.216779e-16, 9.939454e-16, 
    1.158302e-15, 1.130333e-15, 9.637675e-16, 1.131116e-15,
  6.122233e-16, 6.914517e-16, 7.559182e-16, 6.055299e-16, 4.912664e-16, 
    5.265776e-16, 6.283761e-16, 7.087501e-16, 7.667162e-16, 8.966479e-16, 
    9.399676e-16, 7.637179e-16, 5.604284e-16, 4.567469e-16, 3.63269e-16, 
    2.946113e-16, 2.709313e-16, 2.613767e-16, 2.318047e-16, 2.08474e-16, 
    1.999697e-16, 1.967671e-16, 2.024082e-16, 2.205835e-16, 2.267112e-16, 
    2.386173e-16, 2.971584e-16, 4.327507e-16, 5.337622e-16,
  1.227217e-16, 1.153255e-16, 1.276639e-16, 1.291311e-16, 1.261255e-16, 
    1.414832e-16, 1.646065e-16, 1.890866e-16, 1.95499e-16, 2.133356e-16, 
    2.887494e-16, 3.464631e-16, 3.583424e-16, 3.567489e-16, 3.234064e-16, 
    2.896388e-16, 2.636939e-16, 2.100531e-16, 1.747322e-16, 1.336988e-16, 
    1.205297e-16, 1.084412e-16, 1.011227e-16, 1.001991e-16, 1.054946e-16, 
    1.036998e-16, 1.02836e-16, 1.155357e-16, 1.20977e-16,
  5.171643e-17, 5.58904e-17, 5.770989e-17, 4.902152e-17, 4.339376e-17, 
    4.156834e-17, 4.226082e-17, 6.030188e-17, 8.39426e-17, 1.069171e-16, 
    1.224777e-16, 1.534823e-16, 1.911201e-16, 2.048873e-16, 1.968826e-16, 
    1.749658e-16, 1.500674e-16, 1.345178e-16, 1.181342e-16, 1.148847e-16, 
    1.047852e-16, 9.644999e-17, 9.184493e-17, 8.603843e-17, 7.557828e-17, 
    6.083289e-17, 5.839335e-17, 5.751933e-17, 4.610114e-17,
  5.290143e-17, 5.132156e-17, 4.682543e-17, 3.938491e-17, 3.537971e-17, 
    3.381828e-17, 3.252095e-17, 3.19683e-17, 3.462821e-17, 3.908628e-17, 
    4.587925e-17, 5.56584e-17, 6.342989e-17, 7.299849e-17, 8.490582e-17, 
    8.901162e-17, 8.614326e-17, 8.267989e-17, 7.895133e-17, 7.430841e-17, 
    7.475366e-17, 7.647009e-17, 7.743305e-17, 7.470773e-17, 6.861118e-17, 
    6.108131e-17, 5.322117e-17, 5.041397e-17, 5.294534e-17,
  2.00547e-18, 2.00547e-18, 2.00547e-18, 2.00547e-18, 2.00547e-18, 
    2.00547e-18, 2.00547e-18, 1.974109e-18, 1.974109e-18, 1.974109e-18, 
    1.974109e-18, 1.974109e-18, 1.974109e-18, 1.974109e-18, 1.987059e-18, 
    1.987059e-18, 1.987059e-18, 1.987059e-18, 1.987059e-18, 1.987059e-18, 
    1.987059e-18, 2.023051e-18, 2.023051e-18, 2.023051e-18, 2.023051e-18, 
    2.023051e-18, 2.023051e-18, 2.023051e-18, 2.00547e-18,
  1.299381e-18, 1.545818e-18, 1.954178e-18, 2.643496e-18, 3.097243e-18, 
    3.189643e-18, 3.547272e-18, 4.03801e-18, 4.579586e-18, 4.825279e-18, 
    5.264691e-18, 5.391157e-18, 5.406425e-18, 5.377715e-18, 4.839027e-18, 
    4.275578e-18, 3.714027e-18, 3.401148e-18, 2.900264e-18, 2.574916e-18, 
    2.548072e-18, 2.432083e-18, 1.963399e-18, 1.539572e-18, 1.198263e-18, 
    1.079008e-18, 1.029032e-18, 1.046434e-18, 1.178617e-18,
  8.063314e-18, 1.086962e-17, 1.279476e-17, 1.493027e-17, 1.665609e-17, 
    1.917945e-17, 2.028704e-17, 1.945343e-17, 1.82639e-17, 1.653227e-17, 
    1.59869e-17, 1.716311e-17, 1.827211e-17, 2.057968e-17, 2.136815e-17, 
    1.964014e-17, 1.566811e-17, 1.082529e-17, 7.113285e-18, 5.939352e-18, 
    4.870333e-18, 3.705732e-18, 2.8231e-18, 2.083049e-18, 2.076069e-18, 
    2.233577e-18, 2.997763e-18, 4.182243e-18, 6.637539e-18,
  1.514905e-16, 1.504096e-16, 1.676375e-16, 1.716208e-16, 1.548526e-16, 
    1.475496e-16, 1.496119e-16, 1.513691e-16, 1.466178e-16, 1.457995e-16, 
    1.570319e-16, 1.532722e-16, 1.518109e-16, 1.449998e-16, 1.338887e-16, 
    1.156564e-16, 1.066007e-16, 7.279287e-17, 3.260053e-17, 2.127045e-17, 
    1.43693e-17, 1.335756e-17, 1.208827e-17, 1.433462e-17, 2.163945e-17, 
    2.99257e-17, 4.831155e-17, 8.185366e-17, 1.360058e-16,
  7.545791e-16, 7.576954e-16, 6.199251e-16, 5.173377e-16, 4.133913e-16, 
    3.857306e-16, 3.727051e-16, 3.744268e-16, 3.550367e-16, 3.709389e-16, 
    3.630198e-16, 3.738911e-16, 4.125025e-16, 4.234354e-16, 4.434574e-16, 
    4.163527e-16, 3.807631e-16, 3.447316e-16, 3.510099e-16, 3.203059e-16, 
    3.040992e-16, 3.111781e-16, 3.233069e-16, 3.604195e-16, 4.955315e-16, 
    6.129271e-16, 7.366432e-16, 7.648927e-16, 7.712498e-16,
  2.335395e-15, 2.418831e-15, 2.318728e-15, 2.363417e-15, 2.242005e-15, 
    2.212949e-15, 2.156285e-15, 2.264077e-15, 2.260602e-15, 2.102842e-15, 
    1.990431e-15, 1.927633e-15, 1.971371e-15, 2.057903e-15, 2.079181e-15, 
    2.060228e-15, 1.8625e-15, 1.676101e-15, 1.718672e-15, 1.759246e-15, 
    1.740557e-15, 1.768161e-15, 1.892193e-15, 1.978971e-15, 2.157801e-15, 
    2.239034e-15, 2.268055e-15, 2.397756e-15, 2.423644e-15,
  6.08073e-15, 6.166678e-15, 6.297265e-15, 6.208868e-15, 6.136232e-15, 
    5.753289e-15, 6.049316e-15, 5.82477e-15, 5.812346e-15, 5.483172e-15, 
    5.306923e-15, 5.196445e-15, 5.317747e-15, 5.279331e-15, 5.368423e-15, 
    5.208511e-15, 5.267122e-15, 5.443113e-15, 5.237932e-15, 5.231773e-15, 
    5.569792e-15, 5.631222e-15, 5.766315e-15, 5.931625e-15, 5.988722e-15, 
    6.089481e-15, 6.287233e-15, 6.315565e-15, 6.127657e-15,
  1.510084e-14, 1.513104e-14, 1.538868e-14, 1.568541e-14, 1.468116e-14, 
    1.452429e-14, 1.450081e-14, 1.405265e-14, 1.379707e-14, 1.363147e-14, 
    1.348123e-14, 1.358025e-14, 1.289564e-14, 1.289394e-14, 1.306933e-14, 
    1.327015e-14, 1.359349e-14, 1.392374e-14, 1.38169e-14, 1.445965e-14, 
    1.512024e-14, 1.517631e-14, 1.556179e-14, 1.579461e-14, 1.604301e-14, 
    1.576933e-14, 1.542242e-14, 1.541581e-14, 1.543393e-14,
  1.6902e-14, 1.682848e-14, 1.736317e-14, 1.695523e-14, 1.698343e-14, 
    1.676246e-14, 1.737439e-14, 1.775699e-14, 1.783047e-14, 1.746672e-14, 
    1.689764e-14, 1.576605e-14, 1.459488e-14, 1.421837e-14, 1.375867e-14, 
    1.357613e-14, 1.34488e-14, 1.345042e-14, 1.38704e-14, 1.453346e-14, 
    1.499179e-14, 1.553447e-14, 1.587901e-14, 1.68451e-14, 1.651725e-14, 
    1.63788e-14, 1.595343e-14, 1.623997e-14, 1.645032e-14,
  1.146037e-14, 1.161644e-14, 1.175977e-14, 1.202523e-14, 1.244994e-14, 
    1.232664e-14, 1.28472e-14, 1.332316e-14, 1.355775e-14, 1.41893e-14, 
    1.408871e-14, 1.269782e-14, 1.1782e-14, 1.174148e-14, 1.154323e-14, 
    1.157241e-14, 1.174714e-14, 1.183648e-14, 1.198899e-14, 1.208619e-14, 
    1.172222e-14, 1.175649e-14, 1.170305e-14, 1.11446e-14, 1.089959e-14, 
    1.155581e-14, 1.156982e-14, 1.128385e-14, 1.153773e-14,
  1.24709e-14, 1.239096e-14, 1.156066e-14, 1.185256e-14, 1.188909e-14, 
    1.319967e-14, 1.338535e-14, 1.365034e-14, 1.421641e-14, 1.39375e-14, 
    1.361701e-14, 1.274653e-14, 1.171986e-14, 1.155419e-14, 1.206336e-14, 
    1.246507e-14, 1.276789e-14, 1.296243e-14, 1.30349e-14, 1.328197e-14, 
    1.331479e-14, 1.265954e-14, 1.266986e-14, 1.23932e-14, 1.220203e-14, 
    1.209003e-14, 1.208664e-14, 1.2297e-14, 1.277199e-14,
  9.78719e-15, 1.037563e-14, 1.049485e-14, 9.669182e-15, 9.276161e-15, 
    9.511424e-15, 1.014303e-14, 1.083022e-14, 9.936654e-15, 9.648743e-15, 
    1.053731e-14, 1.01402e-14, 1.075195e-14, 1.072611e-14, 1.087e-14, 
    1.130958e-14, 1.149455e-14, 1.15516e-14, 1.217681e-14, 1.256934e-14, 
    1.276728e-14, 1.196738e-14, 1.069216e-14, 1.033268e-14, 1.063113e-14, 
    1.043134e-14, 9.865511e-15, 9.787396e-15, 9.957186e-15,
  5.655591e-15, 5.71951e-15, 5.518425e-15, 6.209311e-15, 6.291918e-15, 
    5.901829e-15, 5.600377e-15, 5.913057e-15, 6.036509e-15, 5.237428e-15, 
    4.986222e-15, 5.05071e-15, 5.207248e-15, 5.38459e-15, 6.30142e-15, 
    6.944629e-15, 6.17832e-15, 6.143438e-15, 6.144729e-15, 6.492106e-15, 
    6.889321e-15, 7.173957e-15, 6.827125e-15, 6.701604e-15, 6.793513e-15, 
    7.065737e-15, 6.719269e-15, 6.051928e-15, 5.333585e-15,
  3.254671e-15, 3.023208e-15, 3.324312e-15, 4.145675e-15, 4.106885e-15, 
    3.465745e-15, 3.377287e-15, 3.026835e-15, 3.692589e-15, 3.440967e-15, 
    2.882097e-15, 2.566744e-15, 2.158554e-15, 1.997349e-15, 2.028983e-15, 
    1.824808e-15, 1.517057e-15, 1.182188e-15, 1.405538e-15, 1.43961e-15, 
    1.435357e-15, 1.794379e-15, 2.168656e-15, 2.232937e-15, 2.790978e-15, 
    3.26878e-15, 2.922079e-15, 2.546223e-15, 3.133404e-15,
  1.674837e-15, 1.922067e-15, 1.917449e-15, 1.699706e-15, 1.28469e-15, 
    1.336018e-15, 1.648964e-15, 1.783442e-15, 1.935862e-15, 2.447295e-15, 
    2.291427e-15, 1.909499e-15, 1.634901e-15, 1.063348e-15, 8.512284e-16, 
    6.739019e-16, 5.662395e-16, 5.717481e-16, 5.173171e-16, 5.154854e-16, 
    4.763997e-16, 4.598154e-16, 4.5938e-16, 5.349865e-16, 6.256856e-16, 
    8.405357e-16, 1.051125e-15, 1.457218e-15, 1.593676e-15,
  3.087112e-16, 3.272674e-16, 3.357232e-16, 3.225701e-16, 3.107017e-16, 
    3.258273e-16, 3.770522e-16, 4.475212e-16, 4.806402e-16, 6.230136e-16, 
    8.595915e-16, 1.007808e-15, 9.798188e-16, 9.465272e-16, 8.877013e-16, 
    7.781101e-16, 7.071448e-16, 5.785618e-16, 5.042854e-16, 4.301021e-16, 
    3.788071e-16, 3.444512e-16, 3.082379e-16, 2.731652e-16, 2.671557e-16, 
    2.593377e-16, 2.74711e-16, 2.889286e-16, 3.135799e-16,
  1.15617e-16, 1.337694e-16, 1.755378e-16, 1.813632e-16, 1.241359e-16, 
    9.939769e-17, 1.08535e-16, 1.449407e-16, 2.036488e-16, 3.022856e-16, 
    3.279898e-16, 4.265055e-16, 5.091358e-16, 5.997723e-16, 6.296143e-16, 
    5.759665e-16, 5.088408e-16, 4.464932e-16, 3.773903e-16, 3.587095e-16, 
    3.302923e-16, 3.139052e-16, 2.701922e-16, 2.344476e-16, 1.968595e-16, 
    1.643535e-16, 1.581666e-16, 1.312641e-16, 1.171476e-16,
  1.077997e-16, 1.039697e-16, 1.000944e-16, 9.108993e-17, 8.430679e-17, 
    7.956922e-17, 6.724426e-17, 6.675249e-17, 7.788127e-17, 9.275895e-17, 
    1.126194e-16, 1.348995e-16, 1.526969e-16, 1.853677e-16, 2.208768e-16, 
    2.398723e-16, 2.458363e-16, 2.379422e-16, 2.255306e-16, 2.098124e-16, 
    2.1004e-16, 2.142815e-16, 2.16858e-16, 2.107614e-16, 1.801288e-16, 
    1.424815e-16, 1.217122e-16, 1.137777e-16, 1.091331e-16,
  5.258524e-18, 5.258524e-18, 5.258524e-18, 5.258524e-18, 5.258524e-18, 
    5.258524e-18, 5.258524e-18, 6.030217e-18, 6.030217e-18, 6.030217e-18, 
    6.030217e-18, 6.030217e-18, 6.030217e-18, 6.030217e-18, 5.824785e-18, 
    5.824785e-18, 5.824785e-18, 5.824785e-18, 5.824785e-18, 5.824785e-18, 
    5.824785e-18, 5.131814e-18, 5.131814e-18, 5.131814e-18, 5.131814e-18, 
    5.131814e-18, 5.131814e-18, 5.131814e-18, 5.258524e-18,
  3.388956e-18, 3.675393e-18, 5.293733e-18, 6.711811e-18, 7.821629e-18, 
    9.404795e-18, 1.08197e-17, 1.141201e-17, 1.129875e-17, 1.26982e-17, 
    1.485493e-17, 1.574497e-17, 1.586207e-17, 1.553788e-17, 1.490883e-17, 
    1.266856e-17, 1.026652e-17, 8.831376e-18, 8.274757e-18, 7.444654e-18, 
    6.6939e-18, 5.739259e-18, 4.374356e-18, 3.84295e-18, 2.90378e-18, 
    2.759157e-18, 2.818152e-18, 2.982901e-18, 3.25817e-18,
  2.081845e-17, 2.519371e-17, 3.326851e-17, 3.883094e-17, 4.354286e-17, 
    5.106039e-17, 6.183274e-17, 6.607206e-17, 5.422169e-17, 4.396043e-17, 
    3.926443e-17, 4.162877e-17, 4.908408e-17, 6.086051e-17, 6.346279e-17, 
    5.808849e-17, 5.494973e-17, 3.63431e-17, 2.449601e-17, 1.80149e-17, 
    1.338642e-17, 1.006895e-17, 7.262354e-18, 5.451809e-18, 5.069212e-18, 
    6.272248e-18, 6.778703e-18, 9.316594e-18, 1.621506e-17,
  6.3979e-16, 6.320339e-16, 7.246233e-16, 7.649481e-16, 6.90816e-16, 
    5.959413e-16, 5.880549e-16, 5.675695e-16, 5.318845e-16, 5.077228e-16, 
    5.904527e-16, 5.86682e-16, 5.725994e-16, 5.5134e-16, 4.874119e-16, 
    4.30525e-16, 4.265404e-16, 2.799122e-16, 1.060635e-16, 6.60661e-17, 
    4.17205e-17, 3.677268e-17, 3.322439e-17, 3.188974e-17, 5.029493e-17, 
    8.393227e-17, 1.446101e-16, 3.686463e-16, 5.73452e-16,
  3.187514e-15, 2.95539e-15, 2.887392e-15, 2.031307e-15, 1.739831e-15, 
    1.230212e-15, 1.034265e-15, 1.175809e-15, 1.11766e-15, 1.126266e-15, 
    1.066407e-15, 1.062673e-15, 1.079585e-15, 1.101622e-15, 1.009404e-15, 
    8.933559e-16, 8.813766e-16, 6.6462e-16, 6.223826e-16, 5.120361e-16, 
    3.520945e-16, 3.426784e-16, 4.318561e-16, 6.565547e-16, 1.35295e-15, 
    2.333197e-15, 3.312881e-15, 3.447377e-15, 3.151673e-15,
  6.115039e-15, 6.195752e-15, 6.000391e-15, 5.98859e-15, 4.736287e-15, 
    4.644394e-15, 4.100522e-15, 4.463471e-15, 4.661997e-15, 4.636031e-15, 
    4.547813e-15, 4.630423e-15, 4.926717e-15, 5.347035e-15, 5.495375e-15, 
    5.488314e-15, 5.105541e-15, 4.743368e-15, 4.418779e-15, 4.325695e-15, 
    4.35274e-15, 4.785866e-15, 4.845808e-15, 5.106733e-15, 5.787364e-15, 
    5.646906e-15, 5.977267e-15, 6.16114e-15, 6.538929e-15,
  1.92156e-14, 1.89515e-14, 1.93064e-14, 1.928367e-14, 1.838135e-14, 
    1.753504e-14, 1.781297e-14, 1.824198e-14, 1.804659e-14, 1.695488e-14, 
    1.624963e-14, 1.603416e-14, 1.615792e-14, 1.613308e-14, 1.575839e-14, 
    1.567163e-14, 1.582179e-14, 1.588352e-14, 1.610551e-14, 1.736634e-14, 
    1.81256e-14, 1.711228e-14, 1.735411e-14, 1.875048e-14, 1.871e-14, 
    1.873298e-14, 1.959443e-14, 1.902566e-14, 1.88866e-14,
  5.607849e-14, 5.763772e-14, 5.696446e-14, 5.670508e-14, 5.515809e-14, 
    5.4813e-14, 5.404851e-14, 5.342679e-14, 5.211662e-14, 5.051618e-14, 
    4.996043e-14, 4.846404e-14, 4.693437e-14, 4.684268e-14, 4.752052e-14, 
    4.824378e-14, 4.902467e-14, 5.046466e-14, 5.313925e-14, 5.581524e-14, 
    5.774357e-14, 5.916579e-14, 5.969028e-14, 6.081103e-14, 6.082938e-14, 
    5.931655e-14, 5.746314e-14, 5.478706e-14, 5.497482e-14,
  7.382589e-14, 7.351256e-14, 7.557874e-14, 7.515342e-14, 7.35584e-14, 
    7.384169e-14, 7.354486e-14, 7.446636e-14, 7.287857e-14, 7.229793e-14, 
    7.039257e-14, 6.764056e-14, 6.501223e-14, 6.402966e-14, 6.410894e-14, 
    6.447536e-14, 6.442735e-14, 6.668458e-14, 6.875679e-14, 6.96536e-14, 
    7.059509e-14, 7.232869e-14, 7.265119e-14, 7.170301e-14, 7.403794e-14, 
    7.43e-14, 7.570539e-14, 7.446023e-14, 7.487287e-14,
  6.819587e-14, 6.571603e-14, 6.366024e-14, 6.342688e-14, 6.365103e-14, 
    6.386808e-14, 6.468259e-14, 6.516397e-14, 6.671183e-14, 6.831033e-14, 
    6.764352e-14, 6.689523e-14, 6.495398e-14, 6.260543e-14, 6.207959e-14, 
    6.236796e-14, 6.227045e-14, 6.415563e-14, 6.829944e-14, 7.037308e-14, 
    7.173077e-14, 7.256024e-14, 7.29181e-14, 7.369908e-14, 7.336329e-14, 
    7.270793e-14, 7.21328e-14, 7.129452e-14, 6.989273e-14,
  5.664844e-14, 5.31658e-14, 5.119287e-14, 4.881764e-14, 4.795565e-14, 
    4.85745e-14, 5.119274e-14, 5.248168e-14, 5.352202e-14, 5.559231e-14, 
    5.665667e-14, 5.691877e-14, 5.434593e-14, 5.27774e-14, 5.213056e-14, 
    5.151997e-14, 5.431688e-14, 5.637006e-14, 5.635976e-14, 5.815358e-14, 
    5.762583e-14, 5.796673e-14, 5.929557e-14, 6.06116e-14, 6.23922e-14, 
    5.990499e-14, 5.919424e-14, 5.870787e-14, 5.764054e-14,
  3.345914e-14, 3.382583e-14, 3.289319e-14, 3.169527e-14, 3.092578e-14, 
    3.259802e-14, 3.199437e-14, 3.253619e-14, 3.034588e-14, 2.976104e-14, 
    3.291294e-14, 3.313195e-14, 3.379848e-14, 3.415078e-14, 3.41734e-14, 
    3.469453e-14, 3.443976e-14, 3.530833e-14, 3.788249e-14, 3.938349e-14, 
    4.202907e-14, 4.05866e-14, 3.838861e-14, 3.922278e-14, 4.064597e-14, 
    4.016125e-14, 3.738819e-14, 3.506821e-14, 3.451462e-14,
  1.558331e-14, 1.551431e-14, 1.522159e-14, 1.566727e-14, 1.555395e-14, 
    1.401495e-14, 1.304183e-14, 1.41605e-14, 1.404199e-14, 1.228103e-14, 
    1.211799e-14, 1.313046e-14, 1.322959e-14, 1.358557e-14, 1.517949e-14, 
    1.597308e-14, 1.572538e-14, 1.528061e-14, 1.519106e-14, 1.565747e-14, 
    1.603727e-14, 1.643055e-14, 1.803253e-14, 1.761247e-14, 1.949067e-14, 
    1.906777e-14, 1.788007e-14, 1.620777e-14, 1.42738e-14,
  6.350498e-15, 5.621662e-15, 6.974404e-15, 7.922032e-15, 8.233892e-15, 
    7.53177e-15, 6.75655e-15, 5.68794e-15, 6.371719e-15, 5.665873e-15, 
    5.618473e-15, 4.819853e-15, 4.559657e-15, 3.934388e-15, 4.753888e-15, 
    4.048934e-15, 3.016135e-15, 2.431382e-15, 2.659989e-15, 2.752301e-15, 
    2.833787e-15, 3.908697e-15, 5.017235e-15, 5.068978e-15, 6.385259e-15, 
    6.642233e-15, 5.789543e-15, 5.543665e-15, 6.308436e-15,
  2.984665e-15, 4.005378e-15, 3.513342e-15, 3.10121e-15, 2.428071e-15, 
    2.647909e-15, 3.060444e-15, 3.208125e-15, 3.558193e-15, 4.059521e-15, 
    3.481624e-15, 3.237911e-15, 2.994293e-15, 2.297906e-15, 1.794707e-15, 
    1.37503e-15, 1.147581e-15, 1.190779e-15, 1.052298e-15, 1.070061e-15, 
    1.055921e-15, 1.003774e-15, 9.604133e-16, 1.026157e-15, 1.429118e-15, 
    1.894053e-15, 2.20906e-15, 2.742968e-15, 2.69271e-15,
  6.160063e-16, 6.253963e-16, 5.900574e-16, 5.568397e-16, 7.171387e-16, 
    7.026991e-16, 7.421615e-16, 9.386932e-16, 1.041932e-15, 1.450483e-15, 
    1.781127e-15, 2.024433e-15, 1.862258e-15, 1.765407e-15, 1.803831e-15, 
    1.70487e-15, 1.584403e-15, 1.301764e-15, 1.14986e-15, 1.094709e-15, 
    9.543696e-16, 8.564149e-16, 7.622594e-16, 6.500435e-16, 6.236351e-16, 
    5.62307e-16, 5.556366e-16, 5.968346e-16, 6.38359e-16,
  2.339175e-16, 2.591358e-16, 2.913211e-16, 2.820683e-16, 2.225139e-16, 
    1.662145e-16, 1.992123e-16, 2.423202e-16, 3.401015e-16, 5.294177e-16, 
    6.666658e-16, 8.486158e-16, 1.051081e-15, 1.322088e-15, 1.326874e-15, 
    1.184712e-15, 1.127144e-15, 1.070928e-15, 9.81576e-16, 9.105705e-16, 
    8.792028e-16, 7.703932e-16, 6.403416e-16, 4.78718e-16, 4.108216e-16, 
    3.297277e-16, 2.920261e-16, 2.568094e-16, 2.441667e-16,
  1.384552e-16, 1.629372e-16, 1.800199e-16, 1.722956e-16, 1.457765e-16, 
    1.347895e-16, 1.324006e-16, 1.301501e-16, 1.414433e-16, 1.633836e-16, 
    2.122493e-16, 2.633349e-16, 3.068152e-16, 3.642912e-16, 4.104934e-16, 
    4.407938e-16, 4.588221e-16, 4.85769e-16, 4.750445e-16, 4.444364e-16, 
    4.202378e-16, 4.026789e-16, 3.843802e-16, 3.589944e-16, 2.933248e-16, 
    2.311311e-16, 1.791505e-16, 1.451287e-16, 1.349195e-16,
  1.187743e-17, 1.187743e-17, 1.187743e-17, 1.187743e-17, 1.187743e-17, 
    1.187743e-17, 1.187743e-17, 1.212573e-17, 1.212573e-17, 1.212573e-17, 
    1.212573e-17, 1.212573e-17, 1.212573e-17, 1.212573e-17, 1.194063e-17, 
    1.194063e-17, 1.194063e-17, 1.194063e-17, 1.194063e-17, 1.194063e-17, 
    1.194063e-17, 1.170687e-17, 1.170687e-17, 1.170687e-17, 1.170687e-17, 
    1.170687e-17, 1.170687e-17, 1.170687e-17, 1.187743e-17,
  1.118741e-17, 1.088408e-17, 1.097672e-17, 1.391476e-17, 2.010704e-17, 
    2.20309e-17, 2.544273e-17, 2.808632e-17, 2.948477e-17, 3.256534e-17, 
    3.721348e-17, 3.853303e-17, 3.829368e-17, 3.655238e-17, 3.317333e-17, 
    2.928362e-17, 2.485438e-17, 2.058292e-17, 1.992531e-17, 1.7583e-17, 
    1.400118e-17, 1.216279e-17, 1.112296e-17, 1.053393e-17, 8.347401e-18, 
    9.679634e-18, 1.114028e-17, 1.14787e-17, 1.15808e-17,
  3.475303e-17, 8.000879e-17, 7.776191e-17, 9.80247e-17, 1.120636e-16, 
    1.326416e-16, 1.588015e-16, 1.853357e-16, 1.624114e-16, 1.198461e-16, 
    1.068965e-16, 1.207783e-16, 1.395961e-16, 1.728814e-16, 1.732356e-16, 
    1.402899e-16, 1.283399e-16, 1.05509e-16, 8.162664e-17, 5.450363e-17, 
    3.133447e-17, 2.235699e-17, 1.77428e-17, 1.509734e-17, 1.591088e-17, 
    1.681585e-17, 1.625143e-17, 1.818388e-17, 2.505318e-17,
  3.159006e-15, 2.856386e-15, 2.709902e-15, 2.489831e-15, 2.317235e-15, 
    2.008042e-15, 1.822599e-15, 1.718833e-15, 1.537805e-15, 1.463172e-15, 
    1.708837e-15, 1.766341e-15, 1.919657e-15, 2.063227e-15, 1.871853e-15, 
    1.664418e-15, 1.717839e-15, 1.048269e-15, 3.190505e-16, 2.037954e-16, 
    1.410512e-16, 1.073542e-16, 8.299457e-17, 8.262924e-17, 1.059678e-16, 
    2.117865e-16, 6.352165e-16, 1.789989e-15, 2.908946e-15,
  9.376185e-15, 7.940392e-15, 8.114875e-15, 6.463615e-15, 6.044143e-15, 
    3.914046e-15, 3.09039e-15, 3.347021e-15, 3.318083e-15, 3.464736e-15, 
    3.624825e-15, 3.557155e-15, 3.326324e-15, 3.310573e-15, 2.870542e-15, 
    2.303654e-15, 2.249966e-15, 2.033191e-15, 1.896648e-15, 1.681734e-15, 
    9.27042e-16, 8.05897e-16, 1.044433e-15, 1.983706e-15, 4.2867e-15, 
    7.669146e-15, 9.85356e-15, 8.658209e-15, 8.12168e-15,
  1.604187e-14, 1.545202e-14, 1.481154e-14, 1.466561e-14, 1.162372e-14, 
    1.028795e-14, 9.454069e-15, 9.34362e-15, 9.605447e-15, 9.979806e-15, 
    9.175492e-15, 9.370326e-15, 1.061259e-14, 1.133291e-14, 1.175468e-14, 
    1.136923e-14, 1.117338e-14, 1.138442e-14, 1.04424e-14, 1.042601e-14, 
    1.159319e-14, 1.145969e-14, 1.250926e-14, 1.54886e-14, 1.661277e-14, 
    1.343579e-14, 1.384713e-14, 1.71184e-14, 1.68779e-14,
  5.203256e-14, 5.353449e-14, 5.348684e-14, 5.135398e-14, 4.902718e-14, 
    4.687906e-14, 4.832715e-14, 4.958399e-14, 4.893192e-14, 4.809236e-14, 
    4.387282e-14, 4.379255e-14, 4.247841e-14, 4.03433e-14, 3.922409e-14, 
    3.955739e-14, 3.929979e-14, 4.199528e-14, 4.472112e-14, 4.697653e-14, 
    4.96179e-14, 5.064583e-14, 5.326265e-14, 5.497049e-14, 5.147798e-14, 
    5.406559e-14, 5.516069e-14, 5.241838e-14, 5.158302e-14,
  1.864404e-13, 1.897342e-13, 1.937351e-13, 1.910313e-13, 1.904173e-13, 
    1.886508e-13, 1.885709e-13, 1.865116e-13, 1.731901e-13, 1.689667e-13, 
    1.657896e-13, 1.624995e-13, 1.604254e-13, 1.617839e-13, 1.632903e-13, 
    1.651138e-13, 1.680231e-13, 1.692311e-13, 1.783179e-13, 1.853382e-13, 
    1.947115e-13, 1.99757e-13, 2.029169e-13, 2.067994e-13, 2.011332e-13, 
    1.962713e-13, 1.914235e-13, 1.900257e-13, 1.872105e-13,
  3.118109e-13, 3.091458e-13, 3.01615e-13, 2.902532e-13, 2.895847e-13, 
    2.915009e-13, 2.893786e-13, 2.838547e-13, 2.779036e-13, 2.699809e-13, 
    2.64432e-13, 2.670971e-13, 2.671572e-13, 2.666486e-13, 2.664328e-13, 
    2.661603e-13, 2.706923e-13, 2.748055e-13, 2.817914e-13, 2.93739e-13, 
    2.981094e-13, 3.011599e-13, 3.040097e-13, 3.129949e-13, 3.128987e-13, 
    3.159835e-13, 3.125137e-13, 3.179468e-13, 3.145177e-13,
  3.21479e-13, 3.201848e-13, 3.162148e-13, 3.021719e-13, 3.018713e-13, 
    2.920553e-13, 2.92451e-13, 2.923845e-13, 2.839331e-13, 2.812639e-13, 
    2.855074e-13, 2.875318e-13, 2.860669e-13, 2.918918e-13, 2.865182e-13, 
    2.782735e-13, 2.723593e-13, 2.700483e-13, 2.681367e-13, 2.70462e-13, 
    2.792624e-13, 2.779819e-13, 2.756484e-13, 2.886218e-13, 2.99361e-13, 
    3.073826e-13, 3.114248e-13, 3.187855e-13, 3.238979e-13,
  2.021362e-13, 1.984659e-13, 1.868636e-13, 1.705919e-13, 1.606882e-13, 
    1.614514e-13, 1.592167e-13, 1.616253e-13, 1.589699e-13, 1.665519e-13, 
    1.80681e-13, 1.854423e-13, 1.920871e-13, 1.920888e-13, 1.910946e-13, 
    1.840302e-13, 1.756294e-13, 1.760616e-13, 1.802316e-13, 1.763408e-13, 
    1.729434e-13, 1.826782e-13, 1.907118e-13, 1.960213e-13, 1.970087e-13, 
    2.073368e-13, 2.061572e-13, 2.181012e-13, 2.090725e-13,
  1.190081e-13, 1.110677e-13, 1.01077e-13, 1.012098e-13, 1.013083e-13, 
    9.874583e-14, 9.71161e-14, 9.890535e-14, 9.58793e-14, 9.534845e-14, 
    9.70904e-14, 1.039894e-13, 1.074329e-13, 1.143098e-13, 1.160229e-13, 
    1.131728e-13, 1.096594e-13, 1.169135e-13, 1.200737e-13, 1.206474e-13, 
    1.233086e-13, 1.257616e-13, 1.271799e-13, 1.222923e-13, 1.237089e-13, 
    1.281635e-13, 1.275038e-13, 1.275078e-13, 1.238662e-13,
  4.370994e-14, 4.026492e-14, 3.95705e-14, 4.015485e-14, 3.911699e-14, 
    3.672807e-14, 3.435458e-14, 3.452682e-14, 3.203716e-14, 3.092972e-14, 
    2.997158e-14, 2.920787e-14, 3.114572e-14, 3.109582e-14, 3.442759e-14, 
    3.893294e-14, 4.08092e-14, 4.292132e-14, 4.150425e-14, 4.357864e-14, 
    4.518879e-14, 4.586589e-14, 5.111585e-14, 5.394399e-14, 5.086458e-14, 
    4.757718e-14, 4.655906e-14, 4.597133e-14, 4.22276e-14,
  1.399905e-14, 1.40892e-14, 1.4175e-14, 1.514006e-14, 1.568516e-14, 
    1.462908e-14, 1.356708e-14, 1.183444e-14, 1.144115e-14, 1.033861e-14, 
    1.102335e-14, 9.824406e-15, 9.729073e-15, 7.597415e-15, 7.989997e-15, 
    6.804395e-15, 5.746584e-15, 5.206876e-15, 5.082193e-15, 5.20924e-15, 
    5.838732e-15, 6.431288e-15, 8.887502e-15, 1.094709e-14, 1.223934e-14, 
    1.240879e-14, 1.185848e-14, 1.099817e-14, 1.407421e-14,
  4.126054e-15, 6.086547e-15, 5.859995e-15, 5.525944e-15, 4.650814e-15, 
    4.387776e-15, 4.968117e-15, 5.531931e-15, 6.07194e-15, 6.003769e-15, 
    5.911048e-15, 6.255663e-15, 6.520279e-15, 6.224791e-15, 4.262462e-15, 
    3.3027e-15, 2.40163e-15, 2.518358e-15, 2.426529e-15, 2.552943e-15, 
    2.128378e-15, 1.992193e-15, 1.976982e-15, 2.053063e-15, 2.346022e-15, 
    2.739403e-15, 3.022995e-15, 3.598362e-15, 3.75763e-15,
  1.011492e-15, 1.148434e-15, 9.280526e-16, 8.549911e-16, 1.397028e-15, 
    1.504379e-15, 1.531136e-15, 1.843433e-15, 2.122708e-15, 2.56873e-15, 
    3.397743e-15, 3.604341e-15, 3.516754e-15, 3.377006e-15, 3.58209e-15, 
    3.222203e-15, 3.096001e-15, 2.75179e-15, 2.478336e-15, 2.518968e-15, 
    2.23841e-15, 1.987962e-15, 1.963602e-15, 1.46559e-15, 1.329451e-15, 
    1.111907e-15, 1.071157e-15, 1.01293e-15, 9.860344e-16,
  4.654583e-16, 4.916965e-16, 4.899546e-16, 4.65585e-16, 3.520012e-16, 
    2.970022e-16, 3.001927e-16, 4.026977e-16, 5.633809e-16, 7.882756e-16, 
    1.095006e-15, 1.399739e-15, 1.915291e-15, 2.357271e-15, 2.113562e-15, 
    2.26813e-15, 2.33107e-15, 2.28596e-15, 2.150312e-15, 2.093662e-15, 
    2.12504e-15, 1.830302e-15, 1.385611e-15, 9.563437e-16, 7.656981e-16, 
    5.76818e-16, 5.160754e-16, 4.422525e-16, 4.572966e-16,
  2.052945e-16, 2.251042e-16, 2.571141e-16, 2.689677e-16, 2.538795e-16, 
    2.407404e-16, 2.143344e-16, 2.146608e-16, 2.245647e-16, 2.628572e-16, 
    3.57649e-16, 4.336375e-16, 4.729413e-16, 5.334287e-16, 6.14393e-16, 
    7.404995e-16, 8.858952e-16, 1.009789e-15, 9.844811e-16, 9.006386e-16, 
    7.641471e-16, 6.414803e-16, 5.499046e-16, 5.10493e-16, 4.246131e-16, 
    3.068523e-16, 2.31709e-16, 2.118375e-16, 2.026396e-16,
  2.72789e-17, 2.72789e-17, 2.72789e-17, 2.72789e-17, 2.72789e-17, 
    2.72789e-17, 2.72789e-17, 2.73463e-17, 2.73463e-17, 2.73463e-17, 
    2.73463e-17, 2.73463e-17, 2.73463e-17, 2.73463e-17, 2.697088e-17, 
    2.697088e-17, 2.697088e-17, 2.697088e-17, 2.697088e-17, 2.697088e-17, 
    2.697088e-17, 2.685846e-17, 2.685846e-17, 2.685846e-17, 2.685846e-17, 
    2.685846e-17, 2.685846e-17, 2.685846e-17, 2.72789e-17,
  3.127639e-17, 3.732474e-17, 4.578252e-17, 3.113836e-17, 3.49383e-17, 
    4.441927e-17, 4.743222e-17, 5.362744e-17, 5.886523e-17, 6.800903e-17, 
    7.781299e-17, 8.065724e-17, 8.006582e-17, 7.55457e-17, 6.707258e-17, 
    6.069497e-17, 5.743696e-17, 5.200766e-17, 4.255998e-17, 3.643948e-17, 
    2.946116e-17, 2.571063e-17, 2.581582e-17, 2.65525e-17, 2.286146e-17, 
    3.225108e-17, 3.41893e-17, 3.098461e-17, 2.980638e-17,
  6.002412e-17, 1.069252e-16, 1.953958e-16, 1.802195e-16, 2.189972e-16, 
    2.398546e-16, 2.957098e-16, 3.709363e-16, 3.726161e-16, 2.915953e-16, 
    2.58423e-16, 3.356131e-16, 3.493279e-16, 3.847881e-16, 3.742753e-16, 
    3.257852e-16, 3.225038e-16, 2.837012e-16, 2.448621e-16, 2.008649e-16, 
    1.060532e-16, 6.279559e-17, 4.882172e-17, 4.246183e-17, 4.879624e-17, 
    4.704337e-17, 4.466384e-17, 4.714155e-17, 5.474362e-17,
  6.890621e-15, 6.567263e-15, 6.291316e-15, 5.214076e-15, 5.10474e-15, 
    4.641368e-15, 3.828221e-15, 3.741635e-15, 3.450564e-15, 3.39442e-15, 
    3.807572e-15, 4.075632e-15, 4.740471e-15, 5.390374e-15, 5.02538e-15, 
    4.656002e-15, 4.680997e-15, 2.727342e-15, 9.576381e-16, 6.728581e-16, 
    4.571471e-16, 3.964812e-16, 2.611832e-16, 2.300691e-16, 2.531337e-16, 
    5.412507e-16, 1.588407e-15, 3.616165e-15, 6.178844e-15,
  1.803936e-14, 1.646834e-14, 1.705245e-14, 1.52339e-14, 1.454808e-14, 
    8.954309e-15, 6.535243e-15, 7.541226e-15, 7.890496e-15, 8.809554e-15, 
    9.839917e-15, 9.750187e-15, 7.9753e-15, 6.629391e-15, 5.982884e-15, 
    5.739886e-15, 5.493709e-15, 5.218508e-15, 4.821128e-15, 4.417394e-15, 
    2.550229e-15, 2.094034e-15, 2.381238e-15, 4.23051e-15, 8.554594e-15, 
    1.565399e-14, 1.896061e-14, 1.603662e-14, 1.61512e-14,
  4.530788e-14, 3.784294e-14, 3.635946e-14, 3.824539e-14, 3.046452e-14, 
    2.704191e-14, 2.808789e-14, 2.514089e-14, 2.497797e-14, 2.630253e-14, 
    2.052887e-14, 1.8861e-14, 2.16268e-14, 2.405474e-14, 2.451253e-14, 
    2.366626e-14, 2.200538e-14, 2.108111e-14, 2.027959e-14, 2.238223e-14, 
    2.489406e-14, 2.3752e-14, 2.822027e-14, 3.687394e-14, 4.128727e-14, 
    3.767541e-14, 3.908473e-14, 4.88612e-14, 4.884322e-14,
  1.460789e-13, 1.52852e-13, 1.368131e-13, 1.284911e-13, 1.29067e-13, 
    1.26633e-13, 1.25339e-13, 1.393121e-13, 1.380315e-13, 1.285344e-13, 
    1.234615e-13, 1.227469e-13, 1.156895e-13, 1.097259e-13, 1.047476e-13, 
    1.024409e-13, 9.904436e-14, 1.13126e-13, 1.198526e-13, 1.287766e-13, 
    1.390043e-13, 1.468632e-13, 1.578105e-13, 1.612478e-13, 1.543766e-13, 
    1.566852e-13, 1.496635e-13, 1.387595e-13, 1.404299e-13,
  6.221716e-13, 6.454263e-13, 6.511946e-13, 6.550007e-13, 6.382931e-13, 
    6.296749e-13, 6.074068e-13, 5.912514e-13, 5.959886e-13, 5.812358e-13, 
    5.696135e-13, 5.481019e-13, 5.413581e-13, 5.295529e-13, 5.454472e-13, 
    5.474972e-13, 5.393484e-13, 5.723497e-13, 5.982161e-13, 6.102715e-13, 
    6.420884e-13, 6.670906e-13, 6.515851e-13, 6.635461e-13, 6.526768e-13, 
    6.362153e-13, 6.246788e-13, 6.082896e-13, 6.345407e-13,
  1.101923e-12, 1.075471e-12, 1.060389e-12, 1.037511e-12, 1.034703e-12, 
    9.836812e-13, 1.009912e-12, 1.018801e-12, 1.003772e-12, 9.614856e-13, 
    9.076661e-13, 8.662743e-13, 8.680529e-13, 8.724406e-13, 8.681275e-13, 
    8.6392e-13, 8.668795e-13, 8.875951e-13, 9.277627e-13, 9.608438e-13, 
    9.977258e-13, 1.032779e-12, 1.047832e-12, 1.046225e-12, 1.076452e-12, 
    1.076297e-12, 1.098589e-12, 1.092718e-12, 1.103666e-12,
  9.394598e-13, 9.549914e-13, 9.632125e-13, 9.527076e-13, 9.697359e-13, 
    9.485418e-13, 9.969707e-13, 1.005425e-12, 1.008568e-12, 1.02931e-12, 
    1.030611e-12, 9.818832e-13, 9.799781e-13, 9.505079e-13, 9.6825e-13, 
    9.505399e-13, 9.160135e-13, 9.125236e-13, 9.113687e-13, 9.093326e-13, 
    9.282301e-13, 9.329833e-13, 9.379988e-13, 9.514158e-13, 9.320321e-13, 
    9.074256e-13, 9.343261e-13, 9.213848e-13, 9.392472e-13,
  6.492252e-13, 6.650062e-13, 6.214202e-13, 6.002975e-13, 5.784105e-13, 
    5.531367e-13, 5.49706e-13, 5.447562e-13, 5.478137e-13, 5.642205e-13, 
    5.831599e-13, 6.055997e-13, 6.092952e-13, 6.246962e-13, 6.319933e-13, 
    6.297755e-13, 6.332768e-13, 6.232947e-13, 6.145244e-13, 6.179567e-13, 
    6.124878e-13, 6.059892e-13, 6.165622e-13, 6.240931e-13, 6.189469e-13, 
    6.332307e-13, 6.43909e-13, 6.505274e-13, 6.696573e-13,
  4.156564e-13, 3.998407e-13, 3.705612e-13, 3.658956e-13, 3.632261e-13, 
    3.506697e-13, 3.348226e-13, 3.351169e-13, 3.339799e-13, 3.388316e-13, 
    3.465532e-13, 3.811088e-13, 4.078049e-13, 4.311725e-13, 4.234887e-13, 
    4.301369e-13, 4.679846e-13, 4.795862e-13, 4.744169e-13, 4.514638e-13, 
    4.456992e-13, 4.466296e-13, 4.414494e-13, 4.252751e-13, 4.206594e-13, 
    4.167457e-13, 4.155599e-13, 4.268194e-13, 4.241346e-13,
  1.330857e-13, 1.268708e-13, 1.155124e-13, 1.160872e-13, 1.112792e-13, 
    1.083507e-13, 1.037285e-13, 9.821177e-14, 9.401781e-14, 9.34366e-14, 
    8.989691e-14, 8.29345e-14, 8.332853e-14, 8.313863e-14, 1.053211e-13, 
    1.18405e-13, 1.252365e-13, 1.289837e-13, 1.271464e-13, 1.308388e-13, 
    1.439707e-13, 1.66223e-13, 1.9475e-13, 1.962285e-13, 1.858003e-13, 
    1.69468e-13, 1.568341e-13, 1.418862e-13, 1.356528e-13,
  3.635838e-14, 3.884551e-14, 3.821515e-14, 3.547121e-14, 3.281788e-14, 
    3.030646e-14, 2.865964e-14, 2.543655e-14, 2.507789e-14, 2.419851e-14, 
    2.548139e-14, 2.496208e-14, 2.370764e-14, 2.456611e-14, 2.07177e-14, 
    1.819943e-14, 1.623777e-14, 1.623764e-14, 1.653118e-14, 1.790264e-14, 
    1.590701e-14, 1.55316e-14, 1.760396e-14, 2.250102e-14, 2.519326e-14, 
    2.913112e-14, 2.96881e-14, 2.85494e-14, 3.248937e-14,
  6.297185e-15, 8.514146e-15, 1.110126e-14, 1.241838e-14, 1.170249e-14, 
    9.437967e-15, 1.043864e-14, 1.113516e-14, 1.141232e-14, 1.224995e-14, 
    1.271926e-14, 1.339605e-14, 1.458751e-14, 1.704865e-14, 1.354729e-14, 
    9.20487e-15, 6.382354e-15, 6.728856e-15, 6.755358e-15, 5.951559e-15, 
    5.570807e-15, 5.187332e-15, 5.39525e-15, 5.993073e-15, 4.968016e-15, 
    5.347203e-15, 5.019433e-15, 5.966071e-15, 6.227222e-15,
  2.134547e-15, 2.175083e-15, 2.196225e-15, 1.717957e-15, 2.225472e-15, 
    3.176418e-15, 3.258397e-15, 3.629224e-15, 4.561825e-15, 5.373392e-15, 
    7.573638e-15, 7.990419e-15, 9.65287e-15, 1.085854e-14, 9.987408e-15, 
    8.284017e-15, 7.016029e-15, 6.240123e-15, 6.269289e-15, 6.546309e-15, 
    6.188737e-15, 5.962591e-15, 5.679865e-15, 4.836216e-15, 3.012335e-15, 
    2.939526e-15, 2.560114e-15, 2.648094e-15, 2.130564e-15,
  1.229603e-15, 1.184779e-15, 1.405828e-15, 1.152704e-15, 8.778922e-16, 
    6.876812e-16, 5.857814e-16, 6.911777e-16, 9.164841e-16, 1.193032e-15, 
    2.033039e-15, 2.446811e-15, 4.025912e-15, 4.899933e-15, 4.59012e-15, 
    4.952877e-15, 4.908362e-15, 5.029425e-15, 4.619124e-15, 4.535442e-15, 
    4.769446e-15, 4.387439e-15, 3.857432e-15, 2.586008e-15, 1.762836e-15, 
    1.445256e-15, 1.348358e-15, 1.302574e-15, 1.311496e-15,
  5.398552e-16, 5.114861e-16, 5.026341e-16, 5.073215e-16, 4.781745e-16, 
    4.349011e-16, 4.134499e-16, 3.7855e-16, 3.793962e-16, 4.201145e-16, 
    5.616675e-16, 7.488668e-16, 8.729991e-16, 9.656143e-16, 1.202778e-15, 
    1.558115e-15, 1.919704e-15, 2.238902e-15, 2.323894e-15, 2.230037e-15, 
    1.887618e-15, 1.439801e-15, 1.085105e-15, 9.35005e-16, 7.643834e-16, 
    5.77053e-16, 5.050853e-16, 5.137864e-16, 5.379323e-16,
  6.386993e-17, 6.386993e-17, 6.386993e-17, 6.386993e-17, 6.386993e-17, 
    6.386993e-17, 6.386993e-17, 6.514379e-17, 6.514379e-17, 6.514379e-17, 
    6.514379e-17, 6.514379e-17, 6.514379e-17, 6.514379e-17, 6.427956e-17, 
    6.427956e-17, 6.427956e-17, 6.427956e-17, 6.427956e-17, 6.427956e-17, 
    6.427956e-17, 6.237695e-17, 6.237695e-17, 6.237695e-17, 6.237695e-17, 
    6.237695e-17, 6.237695e-17, 6.237695e-17, 6.386993e-17,
  5.399635e-17, 6.145649e-17, 7.353218e-17, 8.395274e-17, 1.036111e-16, 
    1.008034e-16, 9.645129e-17, 1.125443e-16, 1.29014e-16, 1.418518e-16, 
    1.655332e-16, 1.727689e-16, 1.736604e-16, 1.706169e-16, 1.670374e-16, 
    1.569432e-16, 1.438467e-16, 1.333594e-16, 1.171946e-16, 1.064563e-16, 
    9.027498e-17, 7.703739e-17, 6.910095e-17, 7.704885e-17, 7.868372e-17, 
    7.071191e-17, 5.723579e-17, 5.239099e-17, 5.273041e-17,
  1.516194e-16, 1.832833e-16, 2.750754e-16, 3.648217e-16, 4.409474e-16, 
    4.725071e-16, 5.224111e-16, 5.892204e-16, 6.656405e-16, 6.095999e-16, 
    5.712047e-16, 8.286943e-16, 1.00965e-15, 9.078355e-16, 9.211191e-16, 
    9.682805e-16, 9.764066e-16, 8.300282e-16, 6.868124e-16, 7.050931e-16, 
    5.028642e-16, 2.147248e-16, 1.699911e-16, 1.567723e-16, 1.507708e-16, 
    1.329843e-16, 1.222834e-16, 1.294429e-16, 1.415002e-16,
  7.869748e-15, 8.971832e-15, 1.083026e-14, 9.594517e-15, 8.617051e-15, 
    7.992703e-15, 6.651888e-15, 6.089726e-15, 6.316442e-15, 6.909869e-15, 
    6.978576e-15, 7.746704e-15, 8.511328e-15, 1.023103e-14, 9.78166e-15, 
    9.488197e-15, 9.064277e-15, 5.142145e-15, 3.038064e-15, 2.526215e-15, 
    1.85567e-15, 1.45976e-15, 1.091538e-15, 8.339739e-16, 8.246413e-16, 
    1.852905e-15, 2.865991e-15, 4.427954e-15, 6.65841e-15,
  3.508022e-14, 3.414881e-14, 3.473024e-14, 3.503225e-14, 3.137526e-14, 
    2.100016e-14, 1.502563e-14, 1.620755e-14, 1.733132e-14, 2.067128e-14, 
    2.263503e-14, 2.349181e-14, 2.022174e-14, 1.62588e-14, 1.456838e-14, 
    1.541397e-14, 1.379929e-14, 1.371499e-14, 1.31021e-14, 1.074588e-14, 
    8.589742e-15, 7.717085e-15, 7.530784e-15, 8.14769e-15, 1.167752e-14, 
    2.131015e-14, 3.201363e-14, 2.92569e-14, 3.113157e-14,
  1.144964e-13, 1.012461e-13, 9.794453e-14, 1.083775e-13, 1.048756e-13, 
    8.127405e-14, 9.600827e-14, 9.025259e-14, 8.355098e-14, 8.029097e-14, 
    6.372217e-14, 5.435475e-14, 5.378919e-14, 5.652046e-14, 5.269944e-14, 
    5.041253e-14, 4.647689e-14, 4.172282e-14, 3.911072e-14, 4.121285e-14, 
    4.607553e-14, 4.725174e-14, 5.088459e-14, 6.470147e-14, 7.934794e-14, 
    8.629127e-14, 1.023843e-13, 1.219335e-13, 1.208142e-13,
  4.862479e-13, 4.40786e-13, 4.118751e-13, 3.912854e-13, 3.886343e-13, 
    3.942887e-13, 4.146222e-13, 4.201379e-13, 4.420568e-13, 3.998767e-13, 
    3.952637e-13, 3.633295e-13, 3.328136e-13, 3.085478e-13, 3.072994e-13, 
    3.204128e-13, 3.231514e-13, 3.519912e-13, 3.810652e-13, 3.942286e-13, 
    4.262216e-13, 4.30794e-13, 4.561759e-13, 4.913581e-13, 4.793081e-13, 
    4.735543e-13, 4.164967e-13, 4.011408e-13, 4.291493e-13,
  2.147522e-12, 2.141813e-12, 2.219612e-12, 2.200408e-12, 2.164494e-12, 
    2.143047e-12, 2.038178e-12, 2.035211e-12, 1.997967e-12, 2.0115e-12, 
    1.998719e-12, 1.91372e-12, 1.89059e-12, 1.82126e-12, 1.816064e-12, 
    1.793469e-12, 1.847175e-12, 1.891682e-12, 1.951497e-12, 2.013075e-12, 
    2.103108e-12, 2.152989e-12, 2.212375e-12, 2.26084e-12, 2.216467e-12, 
    2.154592e-12, 2.115519e-12, 2.124904e-12, 2.10538e-12,
  3.562183e-12, 3.547177e-12, 3.451847e-12, 3.549445e-12, 3.555072e-12, 
    3.335538e-12, 3.22576e-12, 3.379527e-12, 3.392697e-12, 3.362525e-12, 
    3.225389e-12, 3.149774e-12, 3.038132e-12, 2.954731e-12, 2.867383e-12, 
    2.831309e-12, 2.777938e-12, 2.759446e-12, 2.878915e-12, 3.015025e-12, 
    3.026433e-12, 3.13069e-12, 3.305719e-12, 3.35373e-12, 3.40483e-12, 
    3.43946e-12, 3.637431e-12, 3.610249e-12, 3.596606e-12,
  3.052508e-12, 3.000262e-12, 2.978378e-12, 2.956002e-12, 2.944261e-12, 
    2.896662e-12, 2.876508e-12, 2.96681e-12, 3.106566e-12, 3.210769e-12, 
    3.277605e-12, 3.353876e-12, 3.248727e-12, 3.142228e-12, 3.107545e-12, 
    3.110952e-12, 3.070827e-12, 3.006831e-12, 2.9875e-12, 2.925394e-12, 
    2.929784e-12, 3.074329e-12, 3.156972e-12, 3.155387e-12, 3.120056e-12, 
    3.06765e-12, 3.038247e-12, 2.977341e-12, 2.997682e-12,
  2.393714e-12, 2.325095e-12, 2.228308e-12, 2.231911e-12, 2.103455e-12, 
    1.979699e-12, 1.926771e-12, 1.972847e-12, 1.99748e-12, 2.041894e-12, 
    2.117619e-12, 2.132901e-12, 2.141538e-12, 2.11413e-12, 2.121116e-12, 
    2.153188e-12, 2.21326e-12, 2.227219e-12, 2.226844e-12, 2.267818e-12, 
    2.225055e-12, 2.18949e-12, 2.226074e-12, 2.272387e-12, 2.358758e-12, 
    2.385155e-12, 2.308755e-12, 2.400232e-12, 2.356556e-12,
  1.436728e-12, 1.431776e-12, 1.377474e-12, 1.306858e-12, 1.346896e-12, 
    1.262903e-12, 1.306289e-12, 1.246149e-12, 1.306486e-12, 1.344588e-12, 
    1.402935e-12, 1.423111e-12, 1.450167e-12, 1.442223e-12, 1.475578e-12, 
    1.705968e-12, 1.669511e-12, 1.685217e-12, 1.64961e-12, 1.632045e-12, 
    1.6374e-12, 1.537254e-12, 1.540638e-12, 1.508897e-12, 1.532061e-12, 
    1.516282e-12, 1.445506e-12, 1.425261e-12, 1.465367e-12,
  4.428687e-13, 4.211454e-13, 3.711049e-13, 3.679461e-13, 3.620087e-13, 
    3.441876e-13, 3.534227e-13, 3.520219e-13, 3.363298e-13, 3.231874e-13, 
    2.936366e-13, 2.693298e-13, 2.792767e-13, 2.917002e-13, 3.168752e-13, 
    3.865182e-13, 4.881497e-13, 4.764144e-13, 4.313908e-13, 4.516831e-13, 
    5.028904e-13, 6.206077e-13, 6.66808e-13, 5.889128e-13, 5.417557e-13, 
    5.170276e-13, 5.035365e-13, 4.558885e-13, 4.480928e-13,
  8.123182e-14, 9.918866e-14, 1.05201e-13, 1.007005e-13, 8.681368e-14, 
    8.041921e-14, 7.447513e-14, 6.808538e-14, 6.506247e-14, 6.65142e-14, 
    6.347851e-14, 6.795491e-14, 6.747619e-14, 6.987752e-14, 6.372921e-14, 
    6.05421e-14, 5.40479e-14, 5.375389e-14, 5.737404e-14, 5.264154e-14, 
    4.328416e-14, 4.35639e-14, 4.509956e-14, 6.410891e-14, 7.480338e-14, 
    6.907438e-14, 6.481028e-14, 6.470159e-14, 7.497218e-14,
  1.258297e-14, 1.565293e-14, 2.142793e-14, 2.670854e-14, 2.687729e-14, 
    2.537859e-14, 2.649391e-14, 2.854003e-14, 2.82417e-14, 3.325748e-14, 
    3.474158e-14, 3.649701e-14, 3.620207e-14, 4.226771e-14, 4.257175e-14, 
    3.197332e-14, 2.604475e-14, 2.621341e-14, 2.410168e-14, 1.869562e-14, 
    1.821958e-14, 1.620256e-14, 1.660497e-14, 1.96866e-14, 1.791255e-14, 
    1.553283e-14, 1.446817e-14, 1.256188e-14, 1.236644e-14,
  7.955987e-15, 7.342694e-15, 6.003495e-15, 5.269045e-15, 5.599523e-15, 
    6.342386e-15, 7.125846e-15, 8.085431e-15, 9.908486e-15, 1.352765e-14, 
    1.858051e-14, 2.430658e-14, 3.200754e-14, 3.514289e-14, 3.288456e-14, 
    2.930447e-14, 2.53243e-14, 2.090035e-14, 1.862078e-14, 1.866188e-14, 
    1.767898e-14, 1.79343e-14, 1.710611e-14, 1.81913e-14, 1.277138e-14, 
    8.842761e-15, 7.461735e-15, 7.494435e-15, 7.649166e-15,
  4.665884e-15, 3.745017e-15, 3.526841e-15, 3.743029e-15, 2.921862e-15, 
    2.092336e-15, 1.652836e-15, 1.686741e-15, 2.063986e-15, 2.694337e-15, 
    4.656513e-15, 5.575497e-15, 1.036082e-14, 1.247297e-14, 1.399718e-14, 
    1.209043e-14, 1.157945e-14, 1.339128e-14, 1.377516e-14, 1.418844e-14, 
    1.405495e-14, 1.176194e-14, 1.181086e-14, 1.123015e-14, 5.045018e-15, 
    5.336717e-15, 5.381553e-15, 5.621198e-15, 4.99839e-15,
  1.722561e-15, 1.492303e-15, 1.436305e-15, 1.379386e-15, 1.185236e-15, 
    1.021073e-15, 9.18239e-16, 9.118473e-16, 9.255567e-16, 1.096718e-15, 
    1.290938e-15, 1.677867e-15, 2.038603e-15, 2.401224e-15, 3.184888e-15, 
    3.985142e-15, 4.949164e-15, 6.517563e-15, 7.314204e-15, 7.347807e-15, 
    6.484888e-15, 5.030421e-15, 3.083581e-15, 2.024625e-15, 1.653991e-15, 
    1.410625e-15, 1.332811e-15, 1.588886e-15, 1.744037e-15,
  2.272603e-16, 2.272603e-16, 2.272603e-16, 2.272603e-16, 2.272603e-16, 
    2.272603e-16, 2.272603e-16, 2.360814e-16, 2.360814e-16, 2.360814e-16, 
    2.360814e-16, 2.360814e-16, 2.360814e-16, 2.360814e-16, 2.433287e-16, 
    2.433287e-16, 2.433287e-16, 2.433287e-16, 2.433287e-16, 2.433287e-16, 
    2.433287e-16, 2.313079e-16, 2.313079e-16, 2.313079e-16, 2.313079e-16, 
    2.313079e-16, 2.313079e-16, 2.313079e-16, 2.272603e-16,
  1.596789e-16, 1.650774e-16, 1.75024e-16, 1.786915e-16, 2.017231e-16, 
    2.602506e-16, 3.018847e-16, 3.141911e-16, 3.057642e-16, 3.492627e-16, 
    4.400454e-16, 4.760932e-16, 4.993781e-16, 5.095064e-16, 5.226542e-16, 
    5.408812e-16, 5.112206e-16, 4.627e-16, 4.09975e-16, 3.619354e-16, 
    3.343716e-16, 3.301687e-16, 3.600314e-16, 4.088089e-16, 3.224885e-16, 
    2.222971e-16, 1.856226e-16, 1.679641e-16, 1.628073e-16,
  4.402493e-16, 5.342362e-16, 6.813365e-16, 9.141483e-16, 9.622582e-16, 
    1.206474e-15, 1.257465e-15, 1.314844e-15, 1.605386e-15, 1.653199e-15, 
    1.659173e-15, 2.162308e-15, 2.686367e-15, 2.853744e-15, 2.919489e-15, 
    3.117667e-15, 3.25647e-15, 2.60336e-15, 1.904118e-15, 2.398567e-15, 
    1.567431e-15, 6.816292e-16, 6.905584e-16, 7.45469e-16, 6.059467e-16, 
    4.434514e-16, 3.979294e-16, 3.902783e-16, 4.010345e-16,
  1.245854e-14, 1.464261e-14, 1.903622e-14, 1.707179e-14, 1.487052e-14, 
    1.433154e-14, 1.194537e-14, 1.125492e-14, 1.261997e-14, 1.484617e-14, 
    1.629108e-14, 1.707914e-14, 1.814655e-14, 2.336604e-14, 2.489379e-14, 
    2.333716e-14, 2.198571e-14, 1.491437e-14, 1.181466e-14, 1.015295e-14, 
    8.069622e-15, 5.958036e-15, 4.565163e-15, 3.837158e-15, 3.416957e-15, 
    5.963618e-15, 8.35135e-15, 9.990352e-15, 1.140371e-14,
  7.954602e-14, 8.243735e-14, 8.153076e-14, 8.371435e-14, 7.19472e-14, 
    5.376299e-14, 3.867855e-14, 4.072327e-14, 4.530797e-14, 5.211262e-14, 
    6.183024e-14, 6.485123e-14, 6.335193e-14, 5.909556e-14, 5.173531e-14, 
    5.272315e-14, 4.602698e-14, 4.265749e-14, 4.200349e-14, 3.5405e-14, 
    3.49972e-14, 3.195441e-14, 2.823791e-14, 2.508086e-14, 2.808922e-14, 
    3.709058e-14, 7.254742e-14, 7.003798e-14, 6.78475e-14,
  3.250209e-13, 3.112283e-13, 3.427742e-13, 3.762543e-13, 3.505678e-13, 
    2.489729e-13, 3.132136e-13, 3.520723e-13, 2.582025e-13, 2.178166e-13, 
    1.703178e-13, 1.636801e-13, 1.397055e-13, 1.427847e-13, 1.480849e-13, 
    1.411325e-13, 1.299214e-13, 1.167574e-13, 9.319359e-14, 8.92121e-14, 
    9.500868e-14, 1.113086e-13, 1.243752e-13, 1.671163e-13, 2.487116e-13, 
    2.416116e-13, 2.679082e-13, 3.54223e-13, 3.933628e-13,
  1.445421e-12, 1.427387e-12, 1.369875e-12, 1.34959e-12, 1.354148e-12, 
    1.416237e-12, 1.447991e-12, 1.423401e-12, 1.445901e-12, 1.357564e-12, 
    1.302811e-12, 1.170992e-12, 1.105304e-12, 1.052652e-12, 1.091066e-12, 
    1.092919e-12, 1.137396e-12, 1.324051e-12, 1.433887e-12, 1.435759e-12, 
    1.446935e-12, 1.478458e-12, 1.59407e-12, 1.671945e-12, 1.541976e-12, 
    1.403784e-12, 1.322194e-12, 1.356228e-12, 1.531976e-12,
  7.758927e-12, 7.836811e-12, 7.880254e-12, 7.75378e-12, 7.400142e-12, 
    7.442457e-12, 7.538727e-12, 7.277959e-12, 7.401288e-12, 7.410485e-12, 
    7.009791e-12, 6.827649e-12, 6.617453e-12, 6.751817e-12, 6.738755e-12, 
    6.692762e-12, 6.707581e-12, 6.962797e-12, 7.038395e-12, 7.275442e-12, 
    7.463811e-12, 7.360879e-12, 7.645328e-12, 8.096056e-12, 8.03933e-12, 
    7.773772e-12, 7.70686e-12, 7.819233e-12, 8.000449e-12,
  1.222842e-11, 1.231883e-11, 1.172585e-11, 1.158795e-11, 1.20385e-11, 
    1.135761e-11, 1.131699e-11, 1.107366e-11, 1.14808e-11, 1.187299e-11, 
    1.134168e-11, 1.066125e-11, 1.057138e-11, 9.948554e-12, 9.746122e-12, 
    9.547841e-12, 9.55862e-12, 9.67075e-12, 9.772363e-12, 1.021198e-11, 
    1.040908e-11, 1.052517e-11, 1.064553e-11, 1.110836e-11, 1.121339e-11, 
    1.176369e-11, 1.161315e-11, 1.174819e-11, 1.194871e-11,
  1.063161e-11, 1.04734e-11, 1.050603e-11, 1.035606e-11, 1.018186e-11, 
    1.024041e-11, 1.041604e-11, 1.03815e-11, 1.063514e-11, 1.102471e-11, 
    1.121521e-11, 1.121357e-11, 1.12786e-11, 1.096862e-11, 1.064599e-11, 
    1.055795e-11, 1.080786e-11, 1.101892e-11, 1.107773e-11, 1.10439e-11, 
    1.095329e-11, 1.090508e-11, 1.09764e-11, 1.09575e-11, 1.124171e-11, 
    1.10787e-11, 1.111606e-11, 1.122013e-11, 1.097345e-11,
  8.864776e-12, 8.615569e-12, 8.257269e-12, 8.005947e-12, 7.849514e-12, 
    7.235231e-12, 7.190319e-12, 7.173486e-12, 7.286985e-12, 7.291025e-12, 
    7.752434e-12, 7.55204e-12, 7.561531e-12, 7.613642e-12, 7.742177e-12, 
    7.830202e-12, 7.770377e-12, 8.051899e-12, 8.271995e-12, 8.166097e-12, 
    7.936031e-12, 7.98816e-12, 7.940502e-12, 8.048385e-12, 8.351333e-12, 
    8.495645e-12, 8.674202e-12, 8.866459e-12, 8.861163e-12,
  5.414932e-12, 5.276757e-12, 5.119361e-12, 4.99241e-12, 4.907848e-12, 
    4.7294e-12, 4.462785e-12, 4.626323e-12, 4.96896e-12, 4.868973e-12, 
    4.967152e-12, 4.816774e-12, 4.957468e-12, 4.93306e-12, 5.441612e-12, 
    5.578816e-12, 5.144491e-12, 5.481626e-12, 5.627604e-12, 5.650849e-12, 
    5.760353e-12, 5.470146e-12, 5.150995e-12, 5.228483e-12, 5.310692e-12, 
    5.213485e-12, 5.176811e-12, 5.579193e-12, 5.471052e-12,
  1.415852e-12, 1.383432e-12, 1.327637e-12, 1.196267e-12, 1.127171e-12, 
    1.193257e-12, 1.234738e-12, 1.31255e-12, 1.249955e-12, 1.088151e-12, 
    9.583383e-13, 8.752753e-13, 8.905719e-13, 9.522272e-13, 9.724009e-13, 
    1.392385e-12, 1.800416e-12, 1.791665e-12, 1.447493e-12, 1.399672e-12, 
    1.550729e-12, 1.816316e-12, 1.766002e-12, 1.64425e-12, 1.494726e-12, 
    1.42477e-12, 1.496464e-12, 1.499062e-12, 1.425409e-12,
  2.140587e-13, 2.601168e-13, 3.048178e-13, 3.354346e-13, 2.968324e-13, 
    2.847108e-13, 2.643035e-13, 2.702564e-13, 2.293888e-13, 2.149069e-13, 
    2.087284e-13, 2.073329e-13, 2.458996e-13, 1.881488e-13, 1.661393e-13, 
    1.700263e-13, 1.590344e-13, 1.712918e-13, 1.691375e-13, 1.528408e-13, 
    1.232733e-13, 1.264843e-13, 1.607459e-13, 2.023026e-13, 2.455487e-13, 
    1.978255e-13, 1.65997e-13, 1.83202e-13, 1.961518e-13,
  3.498125e-14, 4.524178e-14, 5.823079e-14, 7.790268e-14, 7.71287e-14, 
    7.53113e-14, 7.967895e-14, 1.005406e-13, 9.379401e-14, 1.005479e-13, 
    1.194633e-13, 1.452796e-13, 1.545982e-13, 1.632016e-13, 1.454002e-13, 
    1.150103e-13, 1.103698e-13, 1.136195e-13, 1.042381e-13, 9.951009e-14, 
    8.498914e-14, 6.495693e-14, 5.505457e-14, 6.124325e-14, 6.78777e-14, 
    5.251038e-14, 5.305024e-14, 4.569728e-14, 3.49966e-14,
  3.243259e-14, 3.094497e-14, 2.715561e-14, 2.257946e-14, 1.996004e-14, 
    1.909648e-14, 1.931508e-14, 2.103951e-14, 2.291387e-14, 3.629e-14, 
    5.298385e-14, 7.247162e-14, 9.89888e-14, 1.085702e-13, 1.336327e-13, 
    1.331206e-13, 1.19359e-13, 9.519864e-14, 7.629503e-14, 6.438066e-14, 
    5.685818e-14, 5.382867e-14, 5.43489e-14, 5.234085e-14, 6.21492e-14, 
    2.964567e-14, 2.704981e-14, 2.595819e-14, 3.040129e-14,
  1.963073e-14, 1.874204e-14, 1.256666e-14, 1.110264e-14, 1.195279e-14, 
    9.449899e-15, 6.869776e-15, 6.639317e-15, 6.532116e-15, 9.092836e-15, 
    1.447362e-14, 1.786488e-14, 3.20424e-14, 4.515588e-14, 5.526345e-14, 
    4.158438e-14, 4.11293e-14, 4.327026e-14, 4.391646e-14, 4.58675e-14, 
    4.454651e-14, 4.044579e-14, 3.435744e-14, 5.196037e-14, 2.203464e-14, 
    2.239443e-14, 1.904585e-14, 1.882215e-14, 2.041123e-14,
  6.942966e-15, 6.416535e-15, 4.968774e-15, 4.192798e-15, 3.517244e-15, 
    3.401611e-15, 3.183977e-15, 3.13675e-15, 3.362958e-15, 3.797909e-15, 
    4.835146e-15, 5.915694e-15, 7.255285e-15, 8.397446e-15, 1.15527e-14, 
    1.508701e-14, 2.034528e-14, 3.16171e-14, 3.568749e-14, 3.616492e-14, 
    3.297134e-14, 2.70962e-14, 1.547425e-14, 7.197991e-15, 5.545025e-15, 
    4.791632e-15, 5.053895e-15, 6.755658e-15, 7.054927e-15,
  9.672524e-16, 9.672524e-16, 9.672524e-16, 9.672524e-16, 9.672524e-16, 
    9.672524e-16, 9.672524e-16, 9.826549e-16, 9.826549e-16, 9.826549e-16, 
    9.826549e-16, 9.826549e-16, 9.826549e-16, 9.826549e-16, 9.961765e-16, 
    9.961765e-16, 9.961765e-16, 9.961765e-16, 9.961765e-16, 9.961765e-16, 
    9.961765e-16, 9.788376e-16, 9.788376e-16, 9.788376e-16, 9.788376e-16, 
    9.788376e-16, 9.788376e-16, 9.788376e-16, 9.672524e-16,
  8.529583e-16, 7.466007e-16, 6.89719e-16, 6.57357e-16, 6.963503e-16, 
    8.023495e-16, 8.701831e-16, 9.774809e-16, 1.186565e-15, 1.503872e-15, 
    1.673107e-15, 1.789602e-15, 1.945605e-15, 1.977607e-15, 1.958546e-15, 
    2.065851e-15, 2.039074e-15, 1.805625e-15, 1.451887e-15, 9.928461e-16, 
    7.986241e-16, 7.930932e-16, 1.017635e-15, 1.338051e-15, 1.283621e-15, 
    1.250016e-15, 1.241025e-15, 1.115475e-15, 9.055223e-16,
  1.412823e-15, 1.655293e-15, 2.110893e-15, 2.814528e-15, 3.398099e-15, 
    3.911433e-15, 4.64412e-15, 4.68377e-15, 5.168878e-15, 5.881491e-15, 
    5.910565e-15, 7.304217e-15, 7.682158e-15, 8.814875e-15, 9.721849e-15, 
    1.122766e-14, 1.173735e-14, 9.264672e-15, 6.40825e-15, 6.821323e-15, 
    5.534501e-15, 2.092283e-15, 2.081732e-15, 2.561841e-15, 2.6735e-15, 
    2.504277e-15, 1.729027e-15, 1.54572e-15, 1.393369e-15,
  3.594381e-14, 3.812792e-14, 4.655852e-14, 5.041783e-14, 4.256336e-14, 
    3.757659e-14, 3.069791e-14, 3.23439e-14, 3.671314e-14, 4.16787e-14, 
    4.71998e-14, 5.063431e-14, 5.670619e-14, 7.256776e-14, 8.595842e-14, 
    8.434756e-14, 8.194108e-14, 6.116708e-14, 5.262964e-14, 4.445651e-14, 
    3.198136e-14, 2.358504e-14, 2.038975e-14, 1.649543e-14, 1.555918e-14, 
    2.242161e-14, 3.190848e-14, 3.182216e-14, 3.311393e-14,
  2.604996e-13, 2.761888e-13, 2.451655e-13, 2.365274e-13, 1.813912e-13, 
    1.495542e-13, 1.208235e-13, 1.247346e-13, 1.348713e-13, 1.895058e-13, 
    2.157319e-13, 2.336659e-13, 2.438678e-13, 2.551496e-13, 2.287016e-13, 
    2.210036e-13, 1.853708e-13, 1.543812e-13, 1.518745e-13, 1.223339e-13, 
    1.288145e-13, 1.290026e-13, 1.138523e-13, 1.030275e-13, 1.0557e-13, 
    1.132743e-13, 2.333657e-13, 2.329716e-13, 2.237337e-13,
  1.303545e-12, 1.185572e-12, 1.262727e-12, 1.248015e-12, 9.994103e-13, 
    7.866873e-13, 9.846279e-13, 1.070592e-12, 6.351082e-13, 5.212389e-13, 
    5.199848e-13, 4.826626e-13, 4.476082e-13, 4.460716e-13, 4.669816e-13, 
    4.42519e-13, 4.133131e-13, 3.820561e-13, 3.406134e-13, 2.899923e-13, 
    2.874157e-13, 3.235868e-13, 3.887051e-13, 5.639422e-13, 1.021518e-12, 
    9.062089e-13, 1.010637e-12, 1.166063e-12, 1.395628e-12,
  4.972377e-12, 5.05687e-12, 4.974054e-12, 4.795732e-12, 5.123728e-12, 
    5.496152e-12, 5.362127e-12, 4.924548e-12, 4.854782e-12, 4.704638e-12, 
    4.405195e-12, 3.924976e-12, 3.804749e-12, 3.892352e-12, 4.039923e-12, 
    4.012051e-12, 4.419768e-12, 4.859276e-12, 5.0864e-12, 5.257049e-12, 
    5.571526e-12, 5.720904e-12, 5.782457e-12, 6.029485e-12, 5.787955e-12, 
    4.946185e-12, 4.732214e-12, 5.122546e-12, 5.041438e-12,
  2.790856e-11, 2.869652e-11, 2.861493e-11, 2.86756e-11, 2.854368e-11, 
    2.798458e-11, 2.750718e-11, 2.750357e-11, 2.750915e-11, 2.704129e-11, 
    2.623663e-11, 2.596739e-11, 2.56955e-11, 2.418923e-11, 2.330699e-11, 
    2.385648e-11, 2.486562e-11, 2.424361e-11, 2.524955e-11, 2.689476e-11, 
    2.777422e-11, 2.866733e-11, 2.977183e-11, 2.912586e-11, 2.894669e-11, 
    2.831685e-11, 2.772591e-11, 2.852025e-11, 2.788465e-11,
  4.011083e-11, 4.095413e-11, 4.183416e-11, 4.268345e-11, 4.16588e-11, 
    3.941499e-11, 4.006561e-11, 4.034044e-11, 3.955436e-11, 4.07844e-11, 
    4.049713e-11, 3.931275e-11, 3.770153e-11, 3.762655e-11, 3.506359e-11, 
    3.365826e-11, 3.350191e-11, 3.365961e-11, 3.411529e-11, 3.566769e-11, 
    3.623864e-11, 3.731427e-11, 3.954853e-11, 3.928014e-11, 3.906568e-11, 
    3.971676e-11, 4.258592e-11, 4.226678e-11, 4.104258e-11,
  3.914598e-11, 3.759789e-11, 3.738977e-11, 3.808253e-11, 3.873917e-11, 
    3.871976e-11, 3.771693e-11, 3.85803e-11, 3.979518e-11, 4.059943e-11, 
    4.190659e-11, 4.341081e-11, 4.189979e-11, 4.260656e-11, 4.233726e-11, 
    4.202899e-11, 4.197135e-11, 4.18622e-11, 4.194258e-11, 4.302622e-11, 
    4.445361e-11, 4.563587e-11, 4.384699e-11, 4.30715e-11, 4.177457e-11, 
    4.153934e-11, 4.099314e-11, 4.147341e-11, 4.083954e-11,
  3.184391e-11, 3.044483e-11, 2.932622e-11, 2.982373e-11, 2.816621e-11, 
    2.656688e-11, 2.579299e-11, 2.533327e-11, 2.489357e-11, 2.579303e-11, 
    2.718561e-11, 2.714347e-11, 2.785474e-11, 2.872584e-11, 2.969311e-11, 
    2.949559e-11, 2.896761e-11, 2.956163e-11, 2.981594e-11, 2.906154e-11, 
    2.798977e-11, 2.755676e-11, 2.677914e-11, 2.651064e-11, 2.790849e-11, 
    2.894351e-11, 2.961444e-11, 3.110199e-11, 3.220463e-11,
  2.011034e-11, 2.023793e-11, 1.954281e-11, 1.801452e-11, 1.723918e-11, 
    1.787185e-11, 1.766571e-11, 1.712252e-11, 1.710521e-11, 1.649028e-11, 
    1.675723e-11, 1.635985e-11, 1.692462e-11, 1.7361e-11, 1.932394e-11, 
    1.987433e-11, 1.897299e-11, 1.911496e-11, 2.004921e-11, 1.886104e-11, 
    1.913306e-11, 1.979599e-11, 2.012404e-11, 1.972056e-11, 1.966908e-11, 
    1.934192e-11, 1.983152e-11, 1.957903e-11, 2.070213e-11,
  4.679006e-12, 4.926639e-12, 4.700496e-12, 4.026892e-12, 3.837481e-12, 
    4.1972e-12, 4.320559e-12, 4.394564e-12, 4.357446e-12, 4.073841e-12, 
    3.607524e-12, 3.222743e-12, 3.058458e-12, 3.231475e-12, 3.304679e-12, 
    3.99289e-12, 4.822225e-12, 4.516232e-12, 3.887755e-12, 3.724158e-12, 
    4.023412e-12, 4.59683e-12, 4.454687e-12, 4.595556e-12, 4.536084e-12, 
    4.513376e-12, 5.003659e-12, 4.913912e-12, 4.602302e-12,
  9.139784e-13, 1.008292e-12, 1.147588e-12, 1.102937e-12, 1.035608e-12, 
    1.047202e-12, 1.000776e-12, 1.035708e-12, 8.989259e-13, 8.20765e-13, 
    7.088815e-13, 7.434821e-13, 9.553093e-13, 6.57502e-13, 4.866065e-13, 
    4.877748e-13, 4.268076e-13, 5.885925e-13, 5.316379e-13, 5.280078e-13, 
    4.315352e-13, 4.543542e-13, 6.623509e-13, 6.910404e-13, 7.803398e-13, 
    6.618828e-13, 5.879557e-13, 6.853459e-13, 9.054931e-13,
  1.284972e-13, 1.382963e-13, 1.88335e-13, 2.591096e-13, 2.899049e-13, 
    2.598724e-13, 2.488795e-13, 3.257291e-13, 3.562518e-13, 4.036173e-13, 
    5.415163e-13, 6.533877e-13, 6.872588e-13, 8.026844e-13, 6.076546e-13, 
    4.343116e-13, 4.209906e-13, 4.561592e-13, 4.175367e-13, 3.734682e-13, 
    3.320382e-13, 2.848461e-13, 2.258363e-13, 2.240654e-13, 2.224927e-13, 
    1.839519e-13, 2.059993e-13, 1.827597e-13, 1.365826e-13,
  1.089015e-13, 9.395148e-14, 1.017983e-13, 8.428553e-14, 6.732408e-14, 
    6.565559e-14, 6.118361e-14, 5.714174e-14, 5.676743e-14, 1.035898e-13, 
    1.765096e-13, 2.289925e-13, 3.422015e-13, 4.074508e-13, 5.580726e-13, 
    6.375392e-13, 6.18387e-13, 4.865634e-13, 3.473298e-13, 2.668414e-13, 
    1.973481e-13, 1.94024e-13, 1.658851e-13, 1.723395e-13, 2.131391e-13, 
    1.263192e-13, 1.119199e-13, 1.102774e-13, 1.025416e-13,
  5.827195e-14, 4.988503e-14, 5.169023e-14, 3.322076e-14, 4.139402e-14, 
    4.012277e-14, 2.609924e-14, 2.780217e-14, 2.219318e-14, 3.256176e-14, 
    4.966749e-14, 6.383643e-14, 1.018253e-13, 1.631437e-13, 1.927998e-13, 
    1.560262e-13, 1.517886e-13, 1.596201e-13, 1.596324e-13, 1.557657e-13, 
    1.451711e-13, 1.321144e-13, 1.116829e-13, 1.619288e-13, 1.249443e-13, 
    6.432746e-14, 5.788433e-14, 5.769215e-14, 5.557315e-14,
  3.36802e-14, 2.718187e-14, 2.025419e-14, 1.403883e-14, 9.333312e-15, 
    1.049276e-14, 1.16429e-14, 1.333313e-14, 1.22653e-14, 1.397917e-14, 
    1.710145e-14, 2.221119e-14, 2.744353e-14, 3.230395e-14, 4.363867e-14, 
    5.751265e-14, 8.394496e-14, 1.206228e-13, 1.264103e-13, 1.253918e-13, 
    1.230884e-13, 1.14933e-13, 7.507132e-14, 3.101939e-14, 2.01306e-14, 
    1.75126e-14, 2.515424e-14, 3.277888e-14, 3.466267e-14,
  4.591861e-15, 4.591861e-15, 4.591861e-15, 4.591861e-15, 4.591861e-15, 
    4.591861e-15, 4.591861e-15, 4.452135e-15, 4.452135e-15, 4.452135e-15, 
    4.452135e-15, 4.452135e-15, 4.452135e-15, 4.452135e-15, 4.323085e-15, 
    4.323085e-15, 4.323085e-15, 4.323085e-15, 4.323085e-15, 4.323085e-15, 
    4.323085e-15, 4.469816e-15, 4.469816e-15, 4.469816e-15, 4.469816e-15, 
    4.469816e-15, 4.469816e-15, 4.469816e-15, 4.591861e-15,
  6.189363e-15, 4.978484e-15, 4.237863e-15, 3.887072e-15, 3.858633e-15, 
    4.120116e-15, 4.247341e-15, 4.476316e-15, 4.735701e-15, 5.314549e-15, 
    6.509293e-15, 7.297559e-15, 7.892685e-15, 7.940831e-15, 7.806719e-15, 
    7.301704e-15, 6.786081e-15, 5.764213e-15, 3.819412e-15, 2.764054e-15, 
    1.997342e-15, 1.57161e-15, 1.348498e-15, 1.897773e-15, 3.731834e-15, 
    5.72309e-15, 6.613323e-15, 6.852431e-15, 6.709079e-15,
  5.662443e-15, 6.258735e-15, 8.08454e-15, 1.183202e-14, 1.388325e-14, 
    1.357435e-14, 1.494281e-14, 1.788788e-14, 1.91916e-14, 2.243471e-14, 
    2.478983e-14, 2.734484e-14, 2.736894e-14, 2.865779e-14, 3.158509e-14, 
    3.743282e-14, 3.885561e-14, 3.014044e-14, 1.95241e-14, 1.902167e-14, 
    1.657765e-14, 1.007609e-14, 6.114539e-15, 7.385046e-15, 1.191516e-14, 
    1.171404e-14, 1.120081e-14, 8.233138e-15, 6.290205e-15,
  1.250514e-13, 1.341477e-13, 1.472249e-13, 1.800236e-13, 1.759974e-13, 
    1.56672e-13, 1.215103e-13, 1.249244e-13, 1.309067e-13, 1.407357e-13, 
    1.521806e-13, 1.675784e-13, 1.996988e-13, 2.676901e-13, 3.247753e-13, 
    3.308336e-13, 3.311086e-13, 2.365147e-13, 2.072164e-13, 1.919396e-13, 
    1.32129e-13, 9.538442e-14, 9.481234e-14, 8.565623e-14, 7.370846e-14, 
    1.002457e-13, 1.282785e-13, 1.18433e-13, 1.186853e-13,
  9.349249e-13, 1.166924e-12, 9.359792e-13, 7.877029e-13, 5.803958e-13, 
    5.192658e-13, 4.509453e-13, 4.425489e-13, 4.483343e-13, 7.214183e-13, 
    8.607467e-13, 9.90384e-13, 1.17141e-12, 1.101899e-12, 9.782715e-13, 
    9.611775e-13, 7.695793e-13, 6.675331e-13, 5.814322e-13, 5.209704e-13, 
    4.967095e-13, 5.37299e-13, 5.005195e-13, 4.350745e-13, 4.32207e-13, 
    4.722678e-13, 9.403849e-13, 8.961186e-13, 8.786352e-13,
  3.79758e-12, 3.81049e-12, 3.81052e-12, 3.557401e-12, 2.966798e-12, 
    2.963508e-12, 3.299735e-12, 3.567785e-12, 2.357518e-12, 1.939142e-12, 
    2.104326e-12, 1.8444e-12, 1.653427e-12, 1.602819e-12, 1.520087e-12, 
    1.379286e-12, 1.362231e-12, 1.381156e-12, 1.359285e-12, 1.147754e-12, 
    1.211638e-12, 1.436291e-12, 1.583581e-12, 2.172381e-12, 3.272521e-12, 
    3.396502e-12, 3.496496e-12, 3.689929e-12, 4.079632e-12,
  1.786335e-11, 1.737577e-11, 1.731458e-11, 1.844524e-11, 2.002369e-11, 
    2.08123e-11, 1.88497e-11, 1.776632e-11, 1.709241e-11, 1.576388e-11, 
    1.540843e-11, 1.498073e-11, 1.37713e-11, 1.4149e-11, 1.391191e-11, 
    1.416886e-11, 1.588578e-11, 1.652972e-11, 1.699973e-11, 1.809321e-11, 
    1.935255e-11, 1.968808e-11, 2.089252e-11, 2.168023e-11, 2.001703e-11, 
    1.772247e-11, 1.763203e-11, 1.874755e-11, 1.764613e-11,
  1.076524e-10, 1.081026e-10, 1.080819e-10, 1.066765e-10, 1.070963e-10, 
    1.08343e-10, 1.045819e-10, 1.015176e-10, 1.058759e-10, 1.064918e-10, 
    1.018643e-10, 9.498751e-11, 9.391551e-11, 9.308363e-11, 9.152086e-11, 
    9.201565e-11, 9.313453e-11, 9.175373e-11, 9.769782e-11, 1.004675e-10, 
    1.016566e-10, 1.076454e-10, 1.125271e-10, 1.132832e-10, 1.154098e-10, 
    1.139364e-10, 1.100556e-10, 1.074558e-10, 1.074633e-10,
  1.496796e-10, 1.453922e-10, 1.465075e-10, 1.492716e-10, 1.534643e-10, 
    1.56132e-10, 1.484306e-10, 1.467828e-10, 1.5139e-10, 1.596216e-10, 
    1.537279e-10, 1.476564e-10, 1.445166e-10, 1.394046e-10, 1.388792e-10, 
    1.278372e-10, 1.267553e-10, 1.251662e-10, 1.258034e-10, 1.32229e-10, 
    1.367545e-10, 1.383337e-10, 1.430056e-10, 1.493932e-10, 1.52398e-10, 
    1.511355e-10, 1.5139e-10, 1.48873e-10, 1.505544e-10,
  1.35154e-10, 1.354649e-10, 1.302304e-10, 1.25761e-10, 1.299694e-10, 
    1.320154e-10, 1.386652e-10, 1.414089e-10, 1.435958e-10, 1.500176e-10, 
    1.559529e-10, 1.599758e-10, 1.623732e-10, 1.616213e-10, 1.599071e-10, 
    1.644041e-10, 1.60289e-10, 1.54851e-10, 1.511717e-10, 1.524167e-10, 
    1.530441e-10, 1.553886e-10, 1.528713e-10, 1.56737e-10, 1.499792e-10, 
    1.50426e-10, 1.43675e-10, 1.385583e-10, 1.365935e-10,
  1.096894e-10, 1.059385e-10, 1.016234e-10, 1.020813e-10, 1.007096e-10, 
    9.734108e-11, 9.69262e-11, 9.401341e-11, 9.445936e-11, 9.492241e-11, 
    1.015728e-10, 1.061552e-10, 1.055985e-10, 1.068923e-10, 1.08628e-10, 
    1.126209e-10, 1.142057e-10, 1.140986e-10, 1.13686e-10, 1.14382e-10, 
    1.114159e-10, 1.098659e-10, 1.058316e-10, 1.018041e-10, 1.052611e-10, 
    1.047802e-10, 1.045603e-10, 1.049778e-10, 1.101091e-10,
  7.535018e-11, 7.342273e-11, 7.098699e-11, 7.052039e-11, 6.691216e-11, 
    6.773033e-11, 6.861078e-11, 6.954136e-11, 6.79858e-11, 6.426285e-11, 
    6.264838e-11, 6.335995e-11, 6.35975e-11, 6.600481e-11, 6.870221e-11, 
    7.537609e-11, 7.439347e-11, 7.582299e-11, 7.910752e-11, 7.900858e-11, 
    8.066262e-11, 7.804427e-11, 7.86107e-11, 7.865677e-11, 7.786801e-11, 
    7.483889e-11, 7.517914e-11, 7.651503e-11, 7.820529e-11,
  1.656661e-11, 1.801706e-11, 1.683869e-11, 1.450278e-11, 1.437485e-11, 
    1.471591e-11, 1.474993e-11, 1.425705e-11, 1.382207e-11, 1.450147e-11, 
    1.370532e-11, 1.165964e-11, 1.171097e-11, 1.227363e-11, 1.262711e-11, 
    1.283194e-11, 1.406802e-11, 1.335974e-11, 1.23496e-11, 1.248999e-11, 
    1.279723e-11, 1.464118e-11, 1.4909e-11, 1.627907e-11, 1.581854e-11, 
    1.651078e-11, 1.689947e-11, 1.742131e-11, 1.722308e-11,
  3.486028e-12, 4.098138e-12, 4.452919e-12, 4.134018e-12, 3.366297e-12, 
    3.162936e-12, 3.24448e-12, 3.245417e-12, 3.026861e-12, 3.089093e-12, 
    2.756592e-12, 2.863845e-12, 3.143101e-12, 2.259035e-12, 1.482027e-12, 
    1.522497e-12, 1.38485e-12, 1.841288e-12, 1.867728e-12, 1.897446e-12, 
    1.603382e-12, 1.788462e-12, 2.568913e-12, 2.600562e-12, 2.432012e-12, 
    2.496107e-12, 2.184291e-12, 2.290466e-12, 3.120551e-12,
  4.295291e-13, 4.84225e-13, 5.422167e-13, 6.75739e-13, 8.815433e-13, 
    8.852805e-13, 9.122149e-13, 1.177506e-12, 1.556867e-12, 1.786671e-12, 
    2.148615e-12, 2.474293e-12, 2.54625e-12, 2.863922e-12, 2.390219e-12, 
    1.693789e-12, 1.282974e-12, 1.471406e-12, 1.411326e-12, 1.425727e-12, 
    1.142494e-12, 1.065193e-12, 8.619177e-13, 8.247362e-13, 7.899413e-13, 
    7.414328e-13, 6.094847e-13, 4.855009e-13, 4.201857e-13,
  3.09483e-13, 2.5881e-13, 2.646812e-13, 2.985208e-13, 2.494155e-13, 
    1.872394e-13, 1.741668e-13, 1.548256e-13, 1.508997e-13, 2.759509e-13, 
    5.938199e-13, 8.310006e-13, 1.079043e-12, 1.531494e-12, 2.230408e-12, 
    2.667996e-12, 2.730806e-12, 2.643145e-12, 2.222732e-12, 1.413135e-12, 
    7.656163e-13, 6.558363e-13, 5.156669e-13, 5.493979e-13, 6.357031e-13, 
    4.504387e-13, 3.696807e-13, 3.720763e-13, 3.268559e-13,
  1.327815e-13, 1.408727e-13, 1.275052e-13, 1.218491e-13, 1.002846e-13, 
    1.312024e-13, 8.677001e-14, 9.014564e-14, 6.917859e-14, 9.732878e-14, 
    1.535126e-13, 2.088152e-13, 2.949696e-13, 5.318282e-13, 6.287912e-13, 
    5.733286e-13, 5.346881e-13, 5.304988e-13, 5.431109e-13, 5.004234e-13, 
    4.921055e-13, 4.159376e-13, 3.571466e-13, 4.394599e-13, 4.577063e-13, 
    1.711252e-13, 1.706785e-13, 1.506394e-13, 1.385359e-13,
  8.76493e-14, 8.266446e-14, 5.677702e-14, 3.721672e-14, 2.638148e-14, 
    3.651758e-14, 4.394155e-14, 4.622841e-14, 4.3031e-14, 4.368126e-14, 
    4.717731e-14, 6.580476e-14, 8.34048e-14, 1.138778e-13, 1.607276e-13, 
    2.215144e-13, 3.079685e-13, 3.747538e-13, 3.797296e-13, 3.765874e-13, 
    3.742226e-13, 3.602022e-13, 2.59381e-13, 1.127103e-13, 6.21869e-14, 
    5.349038e-14, 7.332228e-14, 8.666118e-14, 8.882135e-14,
  1.61205e-14, 1.61205e-14, 1.61205e-14, 1.61205e-14, 1.61205e-14, 
    1.61205e-14, 1.61205e-14, 1.580792e-14, 1.580792e-14, 1.580792e-14, 
    1.580792e-14, 1.580792e-14, 1.580792e-14, 1.580792e-14, 1.502787e-14, 
    1.502787e-14, 1.502787e-14, 1.502787e-14, 1.502787e-14, 1.502787e-14, 
    1.502787e-14, 1.528823e-14, 1.528823e-14, 1.528823e-14, 1.528823e-14, 
    1.528823e-14, 1.528823e-14, 1.528823e-14, 1.61205e-14,
  2.657154e-14, 2.419917e-14, 2.205841e-14, 1.993587e-14, 1.845152e-14, 
    1.760713e-14, 1.705839e-14, 1.688105e-14, 1.654078e-14, 1.746899e-14, 
    2.099094e-14, 2.370948e-14, 2.574501e-14, 2.786766e-14, 2.910234e-14, 
    3.000526e-14, 2.561399e-14, 1.976898e-14, 1.085497e-14, 7.167818e-15, 
    6.276732e-15, 5.692949e-15, 4.78534e-15, 4.663067e-15, 7.253432e-15, 
    1.17116e-14, 1.67529e-14, 2.454448e-14, 2.748111e-14,
  3.009428e-14, 2.648682e-14, 3.130825e-14, 4.263302e-14, 6.104282e-14, 
    6.27818e-14, 6.483664e-14, 6.838268e-14, 7.642927e-14, 8.619251e-14, 
    9.219502e-14, 8.881546e-14, 8.831916e-14, 9.452304e-14, 1.114337e-13, 
    1.334766e-13, 1.346228e-13, 1.025804e-13, 7.661217e-14, 7.326484e-14, 
    6.209978e-14, 4.475385e-14, 2.332558e-14, 2.162683e-14, 3.508384e-14, 
    3.889525e-14, 5.42473e-14, 5.374348e-14, 3.644957e-14,
  4.718251e-13, 4.484285e-13, 5.025333e-13, 6.516566e-13, 6.981237e-13, 
    7.278149e-13, 5.394734e-13, 4.808429e-13, 4.758353e-13, 4.662888e-13, 
    4.825807e-13, 5.651839e-13, 6.857658e-13, 9.3931e-13, 1.176906e-12, 
    1.282646e-12, 1.340153e-12, 1.018239e-12, 9.837415e-13, 8.854422e-13, 
    6.240676e-13, 4.408962e-13, 3.67982e-13, 3.945715e-13, 3.213426e-13, 
    4.324211e-13, 4.908042e-13, 4.440061e-13, 4.392262e-13,
  3.632861e-12, 4.067979e-12, 4.567803e-12, 2.710682e-12, 2.163926e-12, 
    1.98085e-12, 1.757768e-12, 1.825231e-12, 1.831245e-12, 2.611323e-12, 
    3.181406e-12, 3.623027e-12, 4.375109e-12, 3.966253e-12, 3.867349e-12, 
    3.644946e-12, 2.960432e-12, 3.37309e-12, 2.186218e-12, 1.84518e-12, 
    1.842227e-12, 2.140167e-12, 2.121944e-12, 1.812752e-12, 1.814504e-12, 
    2.275456e-12, 3.809769e-12, 3.734177e-12, 3.623287e-12,
  9.649911e-12, 1.089522e-11, 1.196872e-11, 1.134726e-11, 1.052263e-11, 
    9.402322e-12, 1.209469e-11, 1.476762e-11, 9.786488e-12, 7.950925e-12, 
    8.371825e-12, 7.197692e-12, 6.22696e-12, 5.869599e-12, 5.104768e-12, 
    4.733891e-12, 4.778659e-12, 5.43327e-12, 5.860334e-12, 4.779074e-12, 
    5.289718e-12, 6.724378e-12, 6.745413e-12, 8.880684e-12, 1.324652e-11, 
    1.443647e-11, 1.176661e-11, 1.066548e-11, 1.06515e-11,
  6.030681e-11, 5.980401e-11, 5.975833e-11, 6.276137e-11, 6.84573e-11, 
    7.32097e-11, 6.325872e-11, 5.781696e-11, 5.62952e-11, 5.604913e-11, 
    5.499066e-11, 5.478502e-11, 5.377512e-11, 4.940538e-11, 4.683638e-11, 
    4.947142e-11, 5.38633e-11, 6.117776e-11, 6.238e-11, 6.305593e-11, 
    6.487653e-11, 7.146345e-11, 7.728714e-11, 8.103551e-11, 7.385637e-11, 
    6.629264e-11, 6.451797e-11, 6.328233e-11, 5.958228e-11,
  4.131215e-10, 4.060512e-10, 4.117025e-10, 3.96971e-10, 4.005874e-10, 
    3.890722e-10, 3.961445e-10, 3.977421e-10, 3.945353e-10, 3.974981e-10, 
    3.791815e-10, 3.645113e-10, 3.518351e-10, 3.357032e-10, 3.370585e-10, 
    3.400525e-10, 3.559301e-10, 3.649026e-10, 3.80306e-10, 3.882196e-10, 
    4.000512e-10, 4.195982e-10, 4.369525e-10, 4.383672e-10, 4.466163e-10, 
    4.36254e-10, 4.444455e-10, 4.293746e-10, 4.132402e-10,
  5.344192e-10, 5.549607e-10, 5.664621e-10, 5.661034e-10, 5.581238e-10, 
    5.266031e-10, 5.488495e-10, 5.748188e-10, 5.782093e-10, 5.868385e-10, 
    5.646244e-10, 5.400418e-10, 5.197288e-10, 5.088292e-10, 4.950564e-10, 
    4.831206e-10, 4.67184e-10, 4.684154e-10, 4.939977e-10, 5.049097e-10, 
    5.178671e-10, 5.485239e-10, 5.528578e-10, 5.723099e-10, 5.834982e-10, 
    5.937768e-10, 5.875139e-10, 5.560042e-10, 5.401876e-10,
  4.664627e-10, 4.631689e-10, 4.691389e-10, 4.62288e-10, 4.515061e-10, 
    4.737749e-10, 4.872706e-10, 5.232228e-10, 5.416723e-10, 5.609749e-10, 
    5.909763e-10, 6.057186e-10, 6.110604e-10, 5.978982e-10, 5.87122e-10, 
    5.79934e-10, 5.575185e-10, 5.446277e-10, 5.302223e-10, 5.268014e-10, 
    5.221363e-10, 5.1658e-10, 5.138198e-10, 5.175664e-10, 5.157304e-10, 
    5.171089e-10, 5.018851e-10, 4.876153e-10, 4.690685e-10,
  3.767371e-10, 3.511886e-10, 3.670913e-10, 3.628862e-10, 3.492857e-10, 
    3.592639e-10, 3.695637e-10, 3.894849e-10, 3.854397e-10, 3.896862e-10, 
    4.131555e-10, 4.58049e-10, 4.623571e-10, 4.707699e-10, 4.659869e-10, 
    4.720747e-10, 4.719747e-10, 4.720378e-10, 4.557288e-10, 4.342453e-10, 
    4.145097e-10, 4.111495e-10, 3.983096e-10, 3.80595e-10, 3.768566e-10, 
    3.813945e-10, 3.737177e-10, 3.759101e-10, 3.851635e-10,
  2.951846e-10, 2.85025e-10, 2.698327e-10, 2.565109e-10, 2.466494e-10, 
    2.60735e-10, 2.660847e-10, 2.485504e-10, 2.434197e-10, 2.363041e-10, 
    2.405529e-10, 2.498493e-10, 2.672226e-10, 2.872743e-10, 3.009914e-10, 
    3.245378e-10, 3.221814e-10, 3.274219e-10, 3.257319e-10, 3.230539e-10, 
    3.315668e-10, 3.267959e-10, 3.113438e-10, 2.925586e-10, 2.908256e-10, 
    3.020708e-10, 3.088767e-10, 3.114152e-10, 3.124221e-10,
  6.251569e-11, 6.37276e-11, 5.905221e-11, 4.8701e-11, 4.676897e-11, 
    4.945314e-11, 4.833497e-11, 4.752294e-11, 4.704336e-11, 4.951303e-11, 
    4.653402e-11, 4.16519e-11, 4.25673e-11, 4.563229e-11, 5.032279e-11, 
    4.496055e-11, 4.751313e-11, 4.488554e-11, 4.354321e-11, 4.401458e-11, 
    4.450454e-11, 4.910887e-11, 5.918736e-11, 6.022269e-11, 6.013779e-11, 
    5.934221e-11, 5.785902e-11, 5.682155e-11, 6.636568e-11,
  1.039176e-11, 1.48866e-11, 1.60707e-11, 1.537854e-11, 1.133545e-11, 
    9.383868e-12, 1.033799e-11, 9.708316e-12, 9.083498e-12, 8.900297e-12, 
    9.028775e-12, 9.589525e-12, 9.988645e-12, 6.869697e-12, 5.380255e-12, 
    5.166633e-12, 5.377802e-12, 6.958904e-12, 7.444778e-12, 7.385379e-12, 
    6.698236e-12, 7.706583e-12, 8.483933e-12, 8.873737e-12, 8.127243e-12, 
    9.770229e-12, 9.219166e-12, 7.473476e-12, 9.416212e-12,
  1.134877e-12, 1.307524e-12, 1.26672e-12, 1.511466e-12, 2.320533e-12, 
    3.129113e-12, 3.223164e-12, 3.456191e-12, 5.094618e-12, 6.052401e-12, 
    6.594251e-12, 7.517867e-12, 8.007208e-12, 7.800455e-12, 6.548506e-12, 
    4.966352e-12, 4.874165e-12, 4.849165e-12, 5.265758e-12, 5.749989e-12, 
    5.699312e-12, 5.082742e-12, 3.398726e-12, 2.625475e-12, 2.663778e-12, 
    2.576877e-12, 2.064716e-12, 1.31215e-12, 1.160801e-12,
  1.079125e-12, 8.849154e-13, 7.819379e-13, 7.345886e-13, 7.275772e-13, 
    5.513308e-13, 4.230115e-13, 3.976572e-13, 3.96023e-13, 7.041526e-13, 
    1.61169e-12, 2.697664e-12, 3.608731e-12, 5.522196e-12, 7.84581e-12, 
    9.097852e-12, 9.311828e-12, 9.128893e-12, 1.012088e-11, 8.889087e-12, 
    5.805742e-12, 2.519595e-12, 1.589076e-12, 1.619232e-12, 1.762379e-12, 
    1.497077e-12, 1.208255e-12, 1.076687e-12, 1.138321e-12,
  3.145656e-13, 3.351542e-13, 3.349163e-13, 3.352101e-13, 2.653428e-13, 
    2.769261e-13, 2.623012e-13, 2.064955e-13, 2.043227e-13, 2.664318e-13, 
    4.371214e-13, 5.505476e-13, 8.118871e-13, 1.603749e-12, 2.135996e-12, 
    2.264432e-12, 1.970714e-12, 1.769018e-12, 1.690168e-12, 1.572948e-12, 
    1.463915e-12, 1.213512e-12, 1.067504e-12, 1.176432e-12, 1.209649e-12, 
    4.373959e-13, 3.795561e-13, 3.328187e-13, 3.174549e-13,
  1.431686e-13, 1.468087e-13, 1.444062e-13, 9.846683e-14, 6.5041e-14, 
    7.758748e-14, 1.272122e-13, 1.118075e-13, 1.23739e-13, 1.314955e-13, 
    1.515971e-13, 2.023153e-13, 2.667365e-13, 3.355157e-13, 4.824127e-13, 
    6.78069e-13, 9.051057e-13, 1.049459e-12, 1.024833e-12, 9.821793e-13, 
    9.548879e-13, 8.815757e-13, 6.655262e-13, 3.128043e-13, 1.503009e-13, 
    1.19616e-13, 1.338296e-13, 1.435173e-13, 1.439575e-13,
  5.170192e-14, 5.170192e-14, 5.170192e-14, 5.170192e-14, 5.170192e-14, 
    5.170192e-14, 5.170192e-14, 4.955567e-14, 4.955567e-14, 4.955567e-14, 
    4.955567e-14, 4.955567e-14, 4.955567e-14, 4.955567e-14, 4.024347e-14, 
    4.024347e-14, 4.024347e-14, 4.024347e-14, 4.024347e-14, 4.024347e-14, 
    4.024347e-14, 4.198124e-14, 4.198124e-14, 4.198124e-14, 4.198124e-14, 
    4.198124e-14, 4.198124e-14, 4.198124e-14, 5.170192e-14,
  9.461897e-14, 9.876561e-14, 9.521563e-14, 7.969796e-14, 6.608922e-14, 
    5.974697e-14, 5.870455e-14, 5.667309e-14, 5.464785e-14, 5.508055e-14, 
    6.358717e-14, 6.979337e-14, 8.101746e-14, 9.48348e-14, 9.935114e-14, 
    9.872981e-14, 7.637093e-14, 5.259125e-14, 3.082233e-14, 2.205678e-14, 
    2.016078e-14, 1.956829e-14, 1.799311e-14, 1.608476e-14, 1.700093e-14, 
    2.572901e-14, 3.696756e-14, 5.538596e-14, 9.384006e-14,
  1.493936e-13, 1.283086e-13, 1.324086e-13, 1.660151e-13, 2.460922e-13, 
    2.342664e-13, 2.335145e-13, 2.435186e-13, 2.726632e-13, 3.316861e-13, 
    3.896072e-13, 3.537299e-13, 3.453376e-13, 3.68762e-13, 4.435606e-13, 
    5.32992e-13, 4.977548e-13, 3.669259e-13, 2.909519e-13, 2.625869e-13, 
    2.345144e-13, 1.756766e-13, 1.023007e-13, 9.282631e-14, 1.157126e-13, 
    1.447779e-13, 1.884967e-13, 2.273612e-13, 1.760646e-13,
  1.653863e-12, 1.564433e-12, 1.55204e-12, 1.87204e-12, 2.399247e-12, 
    2.670763e-12, 2.103479e-12, 1.780253e-12, 1.7774e-12, 1.644354e-12, 
    1.567452e-12, 1.769319e-12, 2.150964e-12, 2.977915e-12, 4.06957e-12, 
    5.049045e-12, 5.489531e-12, 4.757955e-12, 4.246164e-12, 3.578561e-12, 
    2.596355e-12, 1.828313e-12, 1.513324e-12, 1.554625e-12, 1.674659e-12, 
    1.718719e-12, 1.908383e-12, 1.706555e-12, 1.628393e-12,
  1.299253e-11, 1.456333e-11, 1.743112e-11, 1.273557e-11, 7.888078e-12, 
    6.670035e-12, 6.309234e-12, 7.06401e-12, 7.71608e-12, 8.780876e-12, 
    1.017568e-11, 1.193987e-11, 1.516239e-11, 1.403474e-11, 1.42787e-11, 
    1.286021e-11, 1.085182e-11, 1.419544e-11, 8.286693e-12, 6.33299e-12, 
    6.439876e-12, 7.020048e-12, 7.463025e-12, 7.321686e-12, 6.844804e-12, 
    1.14483e-11, 1.403392e-11, 1.516351e-11, 1.254278e-11,
  2.922435e-11, 3.161366e-11, 3.759442e-11, 3.704365e-11, 3.846869e-11, 
    3.266288e-11, 5.17809e-11, 5.287426e-11, 3.785745e-11, 3.200383e-11, 
    3.683699e-11, 2.870937e-11, 2.208001e-11, 2.035109e-11, 1.819752e-11, 
    1.666773e-11, 1.725235e-11, 2.030132e-11, 2.285699e-11, 1.930858e-11, 
    2.206152e-11, 2.760904e-11, 2.970874e-11, 4.013468e-11, 5.330901e-11, 
    5.788343e-11, 4.661808e-11, 3.50769e-11, 3.250312e-11,
  2.150125e-10, 2.223294e-10, 2.203449e-10, 2.246443e-10, 2.405988e-10, 
    2.326936e-10, 2.114683e-10, 2.139162e-10, 1.964358e-10, 2.093482e-10, 
    2.043312e-10, 1.946544e-10, 1.947584e-10, 1.766255e-10, 1.686744e-10, 
    1.721881e-10, 1.945419e-10, 2.20323e-10, 2.264064e-10, 2.264265e-10, 
    2.415931e-10, 2.693117e-10, 3.025179e-10, 3.027338e-10, 2.725669e-10, 
    2.451932e-10, 2.311442e-10, 2.255043e-10, 2.132839e-10,
  1.566765e-09, 1.531677e-09, 1.521214e-09, 1.511025e-09, 1.508665e-09, 
    1.541305e-09, 1.520491e-09, 1.459958e-09, 1.495664e-09, 1.486305e-09, 
    1.46367e-09, 1.390022e-09, 1.362125e-09, 1.328637e-09, 1.301612e-09, 
    1.281583e-09, 1.324368e-09, 1.39755e-09, 1.433728e-09, 1.475583e-09, 
    1.537165e-09, 1.605967e-09, 1.684927e-09, 1.76429e-09, 1.70828e-09, 
    1.672368e-09, 1.646069e-09, 1.597286e-09, 1.555054e-09,
  2.152029e-09, 2.07497e-09, 2.063674e-09, 2.159478e-09, 2.121131e-09, 
    2.196138e-09, 2.145992e-09, 2.242901e-09, 2.325278e-09, 2.308101e-09, 
    2.207241e-09, 2.035808e-09, 1.953347e-09, 1.915711e-09, 1.939551e-09, 
    1.84858e-09, 1.819986e-09, 1.816099e-09, 1.884869e-09, 1.944356e-09, 
    2.064392e-09, 2.110409e-09, 2.213748e-09, 2.228775e-09, 2.305232e-09, 
    2.308663e-09, 2.173553e-09, 2.151263e-09, 2.190932e-09,
  1.734851e-09, 1.731355e-09, 1.738024e-09, 1.779076e-09, 1.801725e-09, 
    1.752702e-09, 1.952512e-09, 2.041621e-09, 2.090823e-09, 2.191176e-09, 
    2.277301e-09, 2.287156e-09, 2.216923e-09, 2.185928e-09, 2.076279e-09, 
    1.956355e-09, 1.890002e-09, 1.874439e-09, 1.808322e-09, 1.746452e-09, 
    1.723834e-09, 1.728504e-09, 1.710545e-09, 1.737618e-09, 1.807789e-09, 
    1.774071e-09, 1.722866e-09, 1.690969e-09, 1.68952e-09,
  1.351602e-09, 1.284058e-09, 1.310431e-09, 1.385926e-09, 1.391507e-09, 
    1.452107e-09, 1.548243e-09, 1.553234e-09, 1.628974e-09, 1.72504e-09, 
    1.889128e-09, 1.936769e-09, 1.910227e-09, 1.841089e-09, 1.832529e-09, 
    1.795886e-09, 1.757704e-09, 1.687166e-09, 1.634845e-09, 1.530944e-09, 
    1.482947e-09, 1.490682e-09, 1.399544e-09, 1.37706e-09, 1.415707e-09, 
    1.461692e-09, 1.450782e-09, 1.353422e-09, 1.373531e-09,
  1.054497e-09, 1.010615e-09, 1.071827e-09, 1.029478e-09, 1.014184e-09, 
    1.036323e-09, 1.048294e-09, 1.02578e-09, 9.711761e-10, 9.52522e-10, 
    9.889362e-10, 1.096117e-09, 1.218346e-09, 1.294676e-09, 1.31007e-09, 
    1.301187e-09, 1.291423e-09, 1.27657e-09, 1.246129e-09, 1.182441e-09, 
    1.114951e-09, 1.1112e-09, 1.169161e-09, 1.13983e-09, 1.155886e-09, 
    1.158613e-09, 1.209718e-09, 1.173784e-09, 1.127711e-09,
  2.361376e-10, 2.276592e-10, 1.941134e-10, 1.678846e-10, 1.738168e-10, 
    1.730864e-10, 1.724423e-10, 1.661097e-10, 1.632002e-10, 1.792237e-10, 
    1.751055e-10, 1.636671e-10, 1.717913e-10, 1.821149e-10, 1.948829e-10, 
    1.887496e-10, 1.857773e-10, 1.713631e-10, 1.612582e-10, 1.585559e-10, 
    1.616653e-10, 1.761905e-10, 2.059961e-10, 2.021289e-10, 1.974503e-10, 
    2.026959e-10, 1.908356e-10, 2.045706e-10, 2.247319e-10,
  2.619446e-11, 3.191063e-11, 4.31967e-11, 4.365294e-11, 3.519324e-11, 
    2.695185e-11, 3.511019e-11, 2.836262e-11, 2.756226e-11, 2.418719e-11, 
    2.855688e-11, 2.927378e-11, 2.874805e-11, 1.974132e-11, 1.902543e-11, 
    1.708547e-11, 1.821341e-11, 2.457783e-11, 2.768518e-11, 2.728788e-11, 
    2.715305e-11, 3.318624e-11, 3.175976e-11, 3.16004e-11, 3.100674e-11, 
    3.494068e-11, 3.408551e-11, 2.978724e-11, 3.094671e-11,
  3.937313e-12, 3.95945e-12, 3.575834e-12, 3.549161e-12, 4.487028e-12, 
    8.295389e-12, 9.058815e-12, 9.34414e-12, 1.241625e-11, 1.839839e-11, 
    2.008205e-11, 1.87703e-11, 2.115944e-11, 2.043488e-11, 1.543644e-11, 
    1.256254e-11, 1.463308e-11, 1.353704e-11, 1.542837e-11, 1.701063e-11, 
    1.929686e-11, 2.047829e-11, 1.79434e-11, 8.855672e-12, 9.850616e-12, 
    9.50533e-12, 7.184644e-12, 4.580696e-12, 3.547726e-12,
  3.435168e-12, 2.908854e-12, 2.600998e-12, 2.228984e-12, 2.023213e-12, 
    1.899305e-12, 1.295991e-12, 1.308353e-12, 1.250356e-12, 2.032141e-12, 
    3.400934e-12, 8.512889e-12, 1.330196e-11, 1.83462e-11, 2.106861e-11, 
    1.974073e-11, 1.851924e-11, 1.797741e-11, 2.111208e-11, 2.528865e-11, 
    2.355211e-11, 1.543099e-11, 4.990685e-12, 4.727771e-12, 5.574975e-12, 
    5.384153e-12, 4.265163e-12, 3.740168e-12, 3.669271e-12,
  9.338505e-13, 9.304495e-13, 1.095059e-12, 1.038431e-12, 9.583629e-13, 
    8.272336e-13, 7.447491e-13, 6.22357e-13, 6.083707e-13, 7.98917e-13, 
    1.320972e-12, 1.571458e-12, 2.094697e-12, 4.038843e-12, 6.720608e-12, 
    8.823085e-12, 9.454808e-12, 1.007474e-11, 7.884577e-12, 5.953107e-12, 
    4.030916e-12, 3.424057e-12, 2.898005e-12, 2.848e-12, 2.95121e-12, 
    9.986815e-13, 8.428736e-13, 7.824134e-13, 9.067832e-13,
  5.315609e-13, 4.974049e-13, 4.487528e-13, 4.29659e-13, 3.091593e-13, 
    2.4805e-13, 3.369833e-13, 3.329304e-13, 2.663858e-13, 3.273092e-13, 
    4.562328e-13, 6.357006e-13, 8.110971e-13, 8.945938e-13, 1.068541e-12, 
    1.513391e-12, 2.073737e-12, 2.524683e-12, 2.550546e-12, 2.379935e-12, 
    2.186272e-12, 1.935179e-12, 1.430656e-12, 6.632614e-13, 3.537327e-13, 
    3.419222e-13, 3.780123e-13, 4.593411e-13, 5.264658e-13,
  8.748715e-14, 8.748715e-14, 8.748715e-14, 8.748715e-14, 8.748715e-14, 
    8.748715e-14, 8.748715e-14, 8.477162e-14, 8.477162e-14, 8.477162e-14, 
    8.477162e-14, 8.477162e-14, 8.477162e-14, 8.477162e-14, 5.636055e-14, 
    5.636055e-14, 5.636055e-14, 5.636055e-14, 5.636055e-14, 5.636055e-14, 
    5.636055e-14, 6.140132e-14, 6.140132e-14, 6.140132e-14, 6.140132e-14, 
    6.140132e-14, 6.140132e-14, 6.140132e-14, 8.748715e-14,
  2.660231e-13, 2.979323e-13, 2.812544e-13, 2.718527e-13, 2.427256e-13, 
    2.171409e-13, 2.318981e-13, 2.253177e-13, 2.227237e-13, 2.208875e-13, 
    2.186269e-13, 2.147674e-13, 2.520101e-13, 2.914314e-13, 2.941088e-13, 
    2.492577e-13, 1.946948e-13, 1.381985e-13, 9.547086e-14, 8.320782e-14, 
    7.696971e-14, 7.312329e-14, 6.967684e-14, 6.22645e-14, 5.087604e-14, 
    6.201951e-14, 8.445564e-14, 1.184102e-13, 2.208045e-13,
  6.866829e-13, 5.585876e-13, 5.607224e-13, 6.073149e-13, 8.703988e-13, 
    9.703192e-13, 9.135027e-13, 9.467927e-13, 1.061695e-12, 1.120429e-12, 
    1.37758e-12, 1.458104e-12, 1.414979e-12, 1.505955e-12, 1.769156e-12, 
    2.05214e-12, 1.687638e-12, 1.28174e-12, 1.056526e-12, 9.396104e-13, 
    8.732586e-13, 6.728676e-13, 4.389271e-13, 4.107082e-13, 4.105488e-13, 
    5.261409e-13, 5.784404e-13, 7.127582e-13, 7.364177e-13,
  5.974546e-12, 4.924014e-12, 4.777671e-12, 5.675285e-12, 7.75819e-12, 
    9.070069e-12, 8.089017e-12, 7.134654e-12, 6.285265e-12, 5.770073e-12, 
    5.269888e-12, 5.087411e-12, 7.067106e-12, 1.006882e-11, 1.296752e-11, 
    1.6773e-11, 1.958382e-11, 1.811698e-11, 1.659293e-11, 1.394683e-11, 
    1.021839e-11, 7.082881e-12, 7.389616e-12, 7.418162e-12, 7.861865e-12, 
    7.703093e-12, 8.953762e-12, 7.059529e-12, 5.540342e-12,
  4.74635e-11, 5.231895e-11, 5.130472e-11, 5.306302e-11, 3.2612e-11, 
    2.480524e-11, 2.356332e-11, 2.410861e-11, 2.746399e-11, 2.426675e-11, 
    3.017846e-11, 4.055534e-11, 5.953561e-11, 4.903113e-11, 4.939272e-11, 
    4.726905e-11, 4.479516e-11, 5.244051e-11, 3.221449e-11, 2.246311e-11, 
    2.354727e-11, 2.425548e-11, 2.455323e-11, 2.602197e-11, 2.44991e-11, 
    4.672057e-11, 4.998071e-11, 5.277782e-11, 4.633887e-11,
  1.246842e-10, 1.032343e-10, 1.219849e-10, 1.213636e-10, 1.140509e-10, 
    1.072118e-10, 1.858389e-10, 1.943331e-10, 1.477002e-10, 1.155542e-10, 
    1.426278e-10, 1.094159e-10, 7.762316e-11, 6.842242e-11, 6.375922e-11, 
    5.981429e-11, 6.142659e-11, 7.388751e-11, 8.073529e-11, 7.802035e-11, 
    8.481819e-11, 1.102081e-10, 1.120667e-10, 1.591361e-10, 2.300601e-10, 
    2.478776e-10, 1.889557e-10, 1.411593e-10, 1.302804e-10,
  7.71851e-10, 7.834688e-10, 7.794155e-10, 8.027498e-10, 8.872129e-10, 
    8.566239e-10, 8.072583e-10, 7.787732e-10, 8.098571e-10, 8.130712e-10, 
    7.92038e-10, 7.469473e-10, 7.057954e-10, 6.575664e-10, 6.360614e-10, 
    6.458563e-10, 7.354887e-10, 7.950315e-10, 8.475273e-10, 8.387236e-10, 
    8.783572e-10, 9.488167e-10, 1.027902e-09, 1.017096e-09, 9.169453e-10, 
    8.499272e-10, 8.361323e-10, 8.197522e-10, 7.754838e-10,
  5.920456e-09, 5.862892e-09, 5.820764e-09, 5.595527e-09, 5.601554e-09, 
    5.912645e-09, 5.674995e-09, 5.661144e-09, 5.903873e-09, 5.719776e-09, 
    5.616885e-09, 5.6765e-09, 5.38504e-09, 5.062884e-09, 5.082358e-09, 
    5.324541e-09, 5.376356e-09, 5.329884e-09, 5.512164e-09, 5.76474e-09, 
    6.032212e-09, 6.217483e-09, 6.27334e-09, 6.198369e-09, 6.377123e-09, 
    6.425636e-09, 6.308184e-09, 6.021137e-09, 5.93282e-09,
  8.466161e-09, 8.328495e-09, 8.163414e-09, 8.368682e-09, 8.367461e-09, 
    8.338364e-09, 8.463173e-09, 8.769846e-09, 8.762754e-09, 8.675249e-09, 
    8.391652e-09, 8.120621e-09, 7.542945e-09, 7.334522e-09, 7.380114e-09, 
    7.237364e-09, 6.80896e-09, 7.081415e-09, 7.433154e-09, 7.906857e-09, 
    8.176921e-09, 8.613495e-09, 8.833065e-09, 9.217914e-09, 9.016198e-09, 
    8.787604e-09, 8.696734e-09, 8.624633e-09, 8.427171e-09,
  6.735504e-09, 6.823785e-09, 6.494777e-09, 6.606277e-09, 6.729895e-09, 
    7.47966e-09, 7.976769e-09, 8.392293e-09, 8.352939e-09, 8.466251e-09, 
    8.318641e-09, 8.337985e-09, 7.586564e-09, 7.3827e-09, 7.069864e-09, 
    6.803976e-09, 6.654986e-09, 6.582584e-09, 6.46958e-09, 6.227813e-09, 
    6.556009e-09, 6.603211e-09, 6.75942e-09, 6.786317e-09, 6.935644e-09, 
    6.64535e-09, 6.495788e-09, 6.560705e-09, 6.553358e-09,
  5.396705e-09, 5.508924e-09, 5.747906e-09, 6.070966e-09, 6.169463e-09, 
    6.511268e-09, 6.600168e-09, 7.00626e-09, 7.090863e-09, 7.086855e-09, 
    7.240505e-09, 7.085987e-09, 6.688996e-09, 6.640062e-09, 6.578504e-09, 
    6.462564e-09, 6.275723e-09, 6.288758e-09, 5.839467e-09, 5.490283e-09, 
    5.529876e-09, 5.802827e-09, 5.58039e-09, 5.6088e-09, 5.700418e-09, 
    5.405238e-09, 5.453912e-09, 5.120532e-09, 5.248432e-09,
  3.85642e-09, 3.798541e-09, 3.991044e-09, 3.780708e-09, 3.739882e-09, 
    3.920631e-09, 3.899248e-09, 3.714581e-09, 3.765599e-09, 4.042571e-09, 
    4.226356e-09, 4.73429e-09, 4.929949e-09, 4.759085e-09, 4.684277e-09, 
    4.700436e-09, 4.603881e-09, 4.292795e-09, 4.27335e-09, 4.189069e-09, 
    4.13304e-09, 4.070416e-09, 4.063162e-09, 4.014326e-09, 4.152156e-09, 
    4.212838e-09, 4.316291e-09, 4.355695e-09, 4.105763e-09,
  8.184105e-10, 7.570531e-10, 6.560965e-10, 6.01863e-10, 6.506394e-10, 
    6.696942e-10, 6.256572e-10, 5.916878e-10, 5.937055e-10, 6.624981e-10, 
    7.104368e-10, 6.883453e-10, 7.830885e-10, 7.397956e-10, 7.312081e-10, 
    7.50318e-10, 7.337349e-10, 6.514762e-10, 6.066966e-10, 6.113398e-10, 
    6.258333e-10, 6.94708e-10, 7.160929e-10, 6.566386e-10, 6.676397e-10, 
    6.63865e-10, 6.338266e-10, 6.681453e-10, 7.457562e-10,
  9.480637e-11, 8.448344e-11, 1.01932e-10, 1.380534e-10, 1.093339e-10, 
    9.089468e-11, 1.040384e-10, 8.844676e-11, 9.194767e-11, 7.81756e-11, 
    9.091676e-11, 9.975246e-11, 9.948045e-11, 7.753579e-11, 6.71134e-11, 
    6.67069e-11, 7.340305e-11, 9.513278e-11, 9.83654e-11, 9.475061e-11, 
    9.830946e-11, 1.209015e-10, 1.12057e-10, 1.119188e-10, 1.110018e-10, 
    1.164737e-10, 1.103145e-10, 1.22818e-10, 1.082097e-10,
  1.872591e-11, 1.717458e-11, 1.65124e-11, 1.689144e-11, 1.682225e-11, 
    2.088528e-11, 2.713523e-11, 2.810676e-11, 3.013797e-11, 5.199269e-11, 
    5.219501e-11, 4.782369e-11, 5.497689e-11, 4.629741e-11, 3.328987e-11, 
    2.986414e-11, 3.377731e-11, 3.284978e-11, 3.50411e-11, 3.522305e-11, 
    3.960988e-11, 4.629391e-11, 4.939168e-11, 4.266444e-11, 4.031178e-11, 
    3.99685e-11, 3.343492e-11, 2.28462e-11, 1.679507e-11,
  1.156807e-11, 1.029383e-11, 8.712427e-12, 7.990477e-12, 6.464359e-12, 
    6.617349e-12, 6.193389e-12, 5.337356e-12, 4.410449e-12, 6.439915e-12, 
    7.701124e-12, 2.53635e-11, 3.619148e-11, 5.048528e-11, 4.739195e-11, 
    4.026559e-11, 3.65245e-11, 3.69087e-11, 3.780916e-11, 4.079641e-11, 
    4.778645e-11, 4.968572e-11, 2.314903e-11, 1.348957e-11, 1.769725e-11, 
    1.765997e-11, 1.285146e-11, 1.134713e-11, 1.150016e-11,
  3.332315e-12, 3.336073e-12, 3.431944e-12, 4.38499e-12, 3.665162e-12, 
    3.479349e-12, 2.408685e-12, 2.391812e-12, 2.01367e-12, 2.505525e-12, 
    3.840318e-12, 4.825209e-12, 5.905396e-12, 9.873793e-12, 2.006701e-11, 
    3.038293e-11, 3.591373e-11, 4.079465e-11, 3.719332e-11, 2.938158e-11, 
    1.477425e-11, 9.406895e-12, 7.519047e-12, 7.989197e-12, 7.835157e-12, 
    3.052551e-12, 2.706218e-12, 3.179902e-12, 3.250282e-12,
  2.298647e-12, 2.656327e-12, 2.605661e-12, 2.022297e-12, 1.683625e-12, 
    1.373259e-12, 1.151298e-12, 1.177818e-12, 9.955825e-13, 9.931414e-13, 
    1.493957e-12, 2.225022e-12, 2.455361e-12, 2.520826e-12, 2.722807e-12, 
    3.489602e-12, 4.614206e-12, 5.966703e-12, 6.394195e-12, 6.096693e-12, 
    5.243632e-12, 4.262378e-12, 2.839895e-12, 1.562959e-12, 1.317273e-12, 
    1.755702e-12, 1.941677e-12, 2.010231e-12, 2.160897e-12,
  1.323306e-13, 1.323306e-13, 1.323306e-13, 1.323306e-13, 1.323306e-13, 
    1.323306e-13, 1.323306e-13, 1.151073e-13, 1.151073e-13, 1.151073e-13, 
    1.151073e-13, 1.151073e-13, 1.151073e-13, 1.151073e-13, 9.917767e-14, 
    9.917767e-14, 9.917767e-14, 9.917767e-14, 9.917767e-14, 9.917767e-14, 
    9.917767e-14, 1.027419e-13, 1.027419e-13, 1.027419e-13, 1.027419e-13, 
    1.027419e-13, 1.027419e-13, 1.027419e-13, 1.323306e-13,
  5.338106e-13, 6.930059e-13, 7.947201e-13, 8.112363e-13, 7.714558e-13, 
    7.538741e-13, 9.176515e-13, 9.675872e-13, 9.127618e-13, 8.871027e-13, 
    8.464764e-13, 8.041901e-13, 7.977091e-13, 7.187035e-13, 6.028625e-13, 
    6.228384e-13, 5.850202e-13, 4.92202e-13, 4.138496e-13, 3.651588e-13, 
    3.415124e-13, 3.187196e-13, 2.812538e-13, 2.491465e-13, 1.951275e-13, 
    1.65117e-13, 2.320187e-13, 2.897292e-13, 4.539046e-13,
  2.24272e-12, 2.014639e-12, 1.929894e-12, 2.22259e-12, 3.279989e-12, 
    3.469839e-12, 3.193116e-12, 3.033783e-12, 3.482519e-12, 3.70804e-12, 
    4.504579e-12, 5.132004e-12, 5.449641e-12, 5.722023e-12, 6.510732e-12, 
    7.110363e-12, 5.725692e-12, 4.722661e-12, 4.08019e-12, 3.561715e-12, 
    3.449883e-12, 2.511935e-12, 1.921722e-12, 1.815289e-12, 1.865125e-12, 
    2.042745e-12, 2.285849e-12, 2.114389e-12, 2.293566e-12,
  1.931394e-11, 1.710293e-11, 1.57289e-11, 1.677307e-11, 2.200683e-11, 
    2.66101e-11, 2.684326e-11, 2.488083e-11, 2.355186e-11, 2.119094e-11, 
    1.783821e-11, 1.68121e-11, 2.179707e-11, 3.116817e-11, 3.912625e-11, 
    5.218069e-11, 5.964398e-11, 5.444315e-11, 5.461581e-11, 5.272413e-11, 
    4.313878e-11, 3.153765e-11, 2.794696e-11, 2.663729e-11, 2.801666e-11, 
    2.850976e-11, 3.129167e-11, 2.803132e-11, 2.204884e-11,
  1.61995e-10, 1.712932e-10, 1.57599e-10, 1.756373e-10, 1.36465e-10, 
    1.078679e-10, 1.046966e-10, 8.973392e-11, 8.798175e-11, 7.402592e-11, 
    8.576984e-11, 1.20885e-10, 2.298886e-10, 1.78633e-10, 1.831825e-10, 
    1.81294e-10, 1.737798e-10, 1.913086e-10, 1.31969e-10, 7.624443e-11, 
    7.795735e-11, 8.370834e-11, 8.950354e-11, 9.438583e-11, 9.295147e-11, 
    1.594255e-10, 1.617053e-10, 1.7046e-10, 1.636066e-10,
  4.473721e-10, 3.855473e-10, 4.184055e-10, 4.030705e-10, 3.515713e-10, 
    3.132602e-10, 4.984512e-10, 6.685804e-10, 4.474533e-10, 4.031423e-10, 
    5.303536e-10, 3.63122e-10, 2.861255e-10, 2.35856e-10, 2.305559e-10, 
    2.163254e-10, 2.133451e-10, 2.881869e-10, 3.261366e-10, 3.181942e-10, 
    3.212029e-10, 4.036191e-10, 3.922425e-10, 4.592894e-10, 7.935753e-10, 
    8.841834e-10, 6.949282e-10, 5.714448e-10, 4.976488e-10,
  2.866571e-09, 2.962939e-09, 2.967017e-09, 2.943645e-09, 3.061721e-09, 
    3.08641e-09, 2.956688e-09, 2.920278e-09, 3.403978e-09, 3.133367e-09, 
    2.963767e-09, 2.627629e-09, 2.562632e-09, 2.493866e-09, 2.449248e-09, 
    2.563733e-09, 2.846692e-09, 2.967581e-09, 3.226036e-09, 3.179668e-09, 
    3.294749e-09, 3.464851e-09, 3.637997e-09, 3.893556e-09, 3.704013e-09, 
    3.287305e-09, 3.084127e-09, 2.910208e-09, 2.825719e-09,
  2.267728e-08, 2.212673e-08, 2.155148e-08, 2.156692e-08, 2.162608e-08, 
    2.145152e-08, 2.11934e-08, 2.137423e-08, 2.196199e-08, 2.289675e-08, 
    2.184601e-08, 2.117164e-08, 2.037155e-08, 2.035377e-08, 1.989627e-08, 
    1.995995e-08, 2.080118e-08, 2.071204e-08, 2.105212e-08, 2.188488e-08, 
    2.284007e-08, 2.368401e-08, 2.447922e-08, 2.445029e-08, 2.378704e-08, 
    2.297674e-08, 2.249488e-08, 2.271731e-08, 2.299319e-08,
  3.413898e-08, 3.395757e-08, 3.418822e-08, 3.475855e-08, 3.602055e-08, 
    3.488416e-08, 3.457577e-08, 3.541246e-08, 3.46884e-08, 3.381445e-08, 
    3.157046e-08, 2.90564e-08, 2.963679e-08, 2.973269e-08, 2.958274e-08, 
    2.790715e-08, 2.670829e-08, 2.84005e-08, 3.007837e-08, 3.208455e-08, 
    3.32627e-08, 3.616458e-08, 3.69465e-08, 3.560159e-08, 3.528117e-08, 
    3.469268e-08, 3.485962e-08, 3.588059e-08, 3.657469e-08,
  2.759779e-08, 2.774676e-08, 2.822932e-08, 2.870964e-08, 2.971091e-08, 
    3.217847e-08, 3.368626e-08, 3.303343e-08, 3.449282e-08, 3.452191e-08, 
    3.25285e-08, 3.145289e-08, 3.011796e-08, 3.02207e-08, 2.843474e-08, 
    2.724099e-08, 2.704046e-08, 2.693981e-08, 2.660239e-08, 2.692149e-08, 
    2.718556e-08, 2.786592e-08, 2.668842e-08, 2.658717e-08, 2.713458e-08, 
    2.65128e-08, 2.653165e-08, 2.614891e-08, 2.701496e-08,
  2.247809e-08, 2.25843e-08, 2.390262e-08, 2.563385e-08, 2.590577e-08, 
    2.640826e-08, 2.762749e-08, 2.670679e-08, 2.775418e-08, 2.732104e-08, 
    2.676381e-08, 2.549355e-08, 2.512871e-08, 2.54769e-08, 2.51641e-08, 
    2.429864e-08, 2.465056e-08, 2.355396e-08, 2.316814e-08, 2.209291e-08, 
    2.205689e-08, 2.072136e-08, 2.040219e-08, 2.170819e-08, 2.123051e-08, 
    2.052434e-08, 2.091486e-08, 2.011541e-08, 2.152015e-08,
  1.433671e-08, 1.430631e-08, 1.571273e-08, 1.536926e-08, 1.47558e-08, 
    1.504183e-08, 1.487824e-08, 1.470378e-08, 1.598765e-08, 1.630665e-08, 
    1.677349e-08, 1.729663e-08, 1.715615e-08, 1.641889e-08, 1.637624e-08, 
    1.699024e-08, 1.650139e-08, 1.60272e-08, 1.560011e-08, 1.4708e-08, 
    1.41379e-08, 1.397938e-08, 1.41244e-08, 1.43218e-08, 1.476651e-08, 
    1.464129e-08, 1.451274e-08, 1.557827e-08, 1.478891e-08,
  2.445678e-09, 2.630879e-09, 2.306389e-09, 2.104694e-09, 2.243241e-09, 
    2.38629e-09, 2.216758e-09, 2.109497e-09, 2.286908e-09, 2.705846e-09, 
    2.868461e-09, 3.060377e-09, 3.463643e-09, 2.931126e-09, 2.845445e-09, 
    2.783964e-09, 2.733431e-09, 2.456127e-09, 2.342331e-09, 2.292658e-09, 
    2.324003e-09, 2.57737e-09, 2.58387e-09, 2.352877e-09, 2.341214e-09, 
    2.269487e-09, 2.21551e-09, 2.157561e-09, 2.349287e-09,
  3.212788e-10, 2.709138e-10, 2.717775e-10, 3.824473e-10, 3.965498e-10, 
    3.948283e-10, 3.752549e-10, 2.881734e-10, 3.053198e-10, 2.598269e-10, 
    2.934363e-10, 3.891459e-10, 4.775261e-10, 3.233082e-10, 2.883489e-10, 
    2.923047e-10, 3.352336e-10, 4.107665e-10, 3.657578e-10, 3.41783e-10, 
    3.387894e-10, 3.969901e-10, 3.884675e-10, 3.610172e-10, 3.693567e-10, 
    3.588828e-10, 3.623345e-10, 4.094571e-10, 3.598616e-10,
  9.242819e-11, 7.961033e-11, 8.144228e-11, 8.159639e-11, 7.668081e-11, 
    7.707698e-11, 7.915553e-11, 7.454422e-11, 8.275571e-11, 1.530313e-10, 
    1.410512e-10, 1.427351e-10, 1.742628e-10, 1.625374e-10, 1.060546e-10, 
    7.332889e-11, 8.50028e-11, 8.400704e-11, 9.205284e-11, 9.686466e-11, 
    9.640415e-11, 1.136936e-10, 1.192211e-10, 1.479075e-10, 1.545827e-10, 
    1.495849e-10, 1.367739e-10, 1.11464e-10, 9.554e-11,
  3.884517e-11, 3.911401e-11, 3.636973e-11, 2.817853e-11, 3.03093e-11, 
    3.356761e-11, 2.919107e-11, 2.334031e-11, 1.87414e-11, 2.11784e-11, 
    2.615514e-11, 5.805258e-11, 1.100012e-10, 1.120521e-10, 1.129674e-10, 
    9.578132e-11, 8.462522e-11, 9.646001e-11, 9.543134e-11, 9.483914e-11, 
    1.080896e-10, 1.150145e-10, 1.012726e-10, 4.599102e-11, 5.57183e-11, 
    5.785082e-11, 4.507976e-11, 3.825228e-11, 3.784145e-11,
  2.098412e-11, 2.146811e-11, 1.887712e-11, 1.834221e-11, 1.778149e-11, 
    1.626573e-11, 1.202832e-11, 9.811213e-12, 9.228959e-12, 9.463558e-12, 
    1.311843e-11, 1.723492e-11, 2.095846e-11, 3.395788e-11, 7.298426e-11, 
    9.223568e-11, 1.069081e-10, 1.203241e-10, 1.227739e-10, 1.147083e-10, 
    6.879869e-11, 3.046375e-11, 2.28456e-11, 2.356513e-11, 2.296974e-11, 
    1.133121e-11, 1.291102e-11, 1.474783e-11, 1.883468e-11,
  7.758605e-12, 9.132762e-12, 1.111376e-11, 1.070761e-11, 7.771031e-12, 
    6.40462e-12, 5.727385e-12, 4.594802e-12, 4.14023e-12, 3.869347e-12, 
    4.982112e-12, 7.483692e-12, 8.12047e-12, 8.813886e-12, 9.816651e-12, 
    1.136481e-11, 1.370478e-11, 1.717568e-11, 1.778293e-11, 1.585514e-11, 
    1.281859e-11, 9.845806e-12, 6.182142e-12, 5.061925e-12, 6.484706e-12, 
    7.524308e-12, 6.958443e-12, 6.857417e-12, 7.283451e-12,
  3.53954e-13, 3.53954e-13, 3.53954e-13, 3.53954e-13, 3.53954e-13, 
    3.53954e-13, 3.53954e-13, 3.623851e-13, 3.623851e-13, 3.623851e-13, 
    3.623851e-13, 3.623851e-13, 3.623851e-13, 3.623851e-13, 3.613755e-13, 
    3.613755e-13, 3.613755e-13, 3.613755e-13, 3.613755e-13, 3.613755e-13, 
    3.613755e-13, 3.483862e-13, 3.483862e-13, 3.483862e-13, 3.483862e-13, 
    3.483862e-13, 3.483862e-13, 3.483862e-13, 3.53954e-13,
  1.325008e-12, 1.546789e-12, 1.622344e-12, 1.632529e-12, 1.852763e-12, 
    2.038594e-12, 2.442345e-12, 2.785355e-12, 2.717181e-12, 2.528347e-12, 
    2.193338e-12, 1.996891e-12, 1.869832e-12, 1.721194e-12, 1.743423e-12, 
    1.909684e-12, 1.967833e-12, 1.888718e-12, 1.740801e-12, 1.653956e-12, 
    1.699286e-12, 1.550215e-12, 1.42621e-12, 1.212931e-12, 9.637874e-13, 
    7.21661e-13, 6.521536e-13, 9.555918e-13, 1.252091e-12,
  7.817822e-12, 7.667407e-12, 6.990848e-12, 7.565905e-12, 1.000295e-11, 
    1.293899e-11, 1.237494e-11, 1.14392e-11, 1.273156e-11, 1.341339e-11, 
    1.457985e-11, 1.757792e-11, 1.884336e-11, 2.003889e-11, 2.097265e-11, 
    2.253955e-11, 1.981312e-11, 1.788401e-11, 1.56883e-11, 1.313303e-11, 
    1.198313e-11, 9.355173e-12, 7.902349e-12, 7.561896e-12, 7.835657e-12, 
    7.934956e-12, 8.3327e-12, 7.979803e-12, 7.576165e-12,
  6.785527e-11, 5.539744e-11, 4.424687e-11, 4.43528e-11, 5.58442e-11, 
    7.043683e-11, 7.871636e-11, 8.178971e-11, 7.843661e-11, 7.402853e-11, 
    6.668076e-11, 6.5064e-11, 7.871882e-11, 1.01317e-10, 1.294377e-10, 
    1.627357e-10, 1.701114e-10, 1.586362e-10, 1.524575e-10, 1.577696e-10, 
    1.516964e-10, 1.208193e-10, 8.968657e-11, 7.910718e-11, 8.276849e-11, 
    8.460024e-11, 8.352179e-11, 8.123456e-11, 7.270112e-11,
  5.375929e-10, 5.369315e-10, 5.175887e-10, 5.726021e-10, 5.033389e-10, 
    4.480823e-10, 4.172724e-10, 3.634955e-10, 3.224514e-10, 2.710434e-10, 
    3.233331e-10, 4.656638e-10, 7.386712e-10, 7.583459e-10, 7.604232e-10, 
    7.651834e-10, 6.595924e-10, 6.411284e-10, 4.671681e-10, 2.482331e-10, 
    2.464031e-10, 2.882035e-10, 3.537638e-10, 4.220543e-10, 3.78334e-10, 
    5.07231e-10, 4.974428e-10, 4.912394e-10, 5.146489e-10,
  1.53893e-09, 1.416792e-09, 1.458439e-09, 1.525595e-09, 1.422747e-09, 
    1.28133e-09, 1.400791e-09, 1.893161e-09, 1.293665e-09, 1.534525e-09, 
    2.02432e-09, 1.510217e-09, 9.99502e-10, 9.233141e-10, 8.473386e-10, 
    7.959712e-10, 8.059736e-10, 1.047742e-09, 1.253506e-09, 1.256226e-09, 
    1.317566e-09, 1.41005e-09, 1.246316e-09, 1.34247e-09, 2.355279e-09, 
    2.761019e-09, 2.349697e-09, 2.068657e-09, 1.720883e-09,
  1.180641e-08, 1.186672e-08, 1.153628e-08, 1.18969e-08, 1.132929e-08, 
    1.139571e-08, 1.121364e-08, 1.072115e-08, 1.255167e-08, 1.19188e-08, 
    1.054311e-08, 1.002165e-08, 9.653694e-09, 9.188795e-09, 9.402775e-09, 
    1.004636e-08, 1.034682e-08, 1.07906e-08, 1.169514e-08, 1.196536e-08, 
    1.214216e-08, 1.264379e-08, 1.415153e-08, 1.558234e-08, 1.492984e-08, 
    1.338321e-08, 1.237173e-08, 1.206524e-08, 1.150362e-08,
  8.734356e-08, 8.539636e-08, 8.332882e-08, 8.226612e-08, 8.294916e-08, 
    8.136755e-08, 8.188853e-08, 8.512821e-08, 8.684184e-08, 8.537252e-08, 
    8.361354e-08, 8.009561e-08, 7.644515e-08, 7.696975e-08, 7.970142e-08, 
    7.769896e-08, 7.870056e-08, 8.260637e-08, 8.564849e-08, 8.80183e-08, 
    9.049879e-08, 9.22149e-08, 9.289786e-08, 9.333872e-08, 9.476593e-08, 
    9.323716e-08, 9.050545e-08, 8.75737e-08, 8.660722e-08,
  1.49198e-07, 1.409663e-07, 1.348758e-07, 1.414175e-07, 1.398645e-07, 
    1.460238e-07, 1.456824e-07, 1.381418e-07, 1.370733e-07, 1.317348e-07, 
    1.271098e-07, 1.216635e-07, 1.23891e-07, 1.239872e-07, 1.205069e-07, 
    1.1322e-07, 1.122989e-07, 1.193574e-07, 1.266283e-07, 1.35872e-07, 
    1.428492e-07, 1.448186e-07, 1.432313e-07, 1.502711e-07, 1.493376e-07, 
    1.476133e-07, 1.459333e-07, 1.457956e-07, 1.474159e-07,
  1.148761e-07, 1.13358e-07, 1.170416e-07, 1.214169e-07, 1.279828e-07, 
    1.298176e-07, 1.319994e-07, 1.345335e-07, 1.366408e-07, 1.412442e-07, 
    1.479283e-07, 1.437086e-07, 1.443802e-07, 1.413901e-07, 1.334587e-07, 
    1.291001e-07, 1.230411e-07, 1.202873e-07, 1.184267e-07, 1.165378e-07, 
    1.159539e-07, 1.154468e-07, 1.12427e-07, 1.104785e-07, 1.110284e-07, 
    1.120504e-07, 1.145443e-07, 1.187455e-07, 1.167097e-07,
  9.002557e-08, 9.291156e-08, 9.445181e-08, 9.767797e-08, 1.042351e-07, 
    1.041264e-07, 1.059734e-07, 1.10143e-07, 1.106101e-07, 1.090467e-07, 
    1.096151e-07, 1.027107e-07, 1.046733e-07, 1.062184e-07, 1.005383e-07, 
    9.619547e-08, 8.875493e-08, 8.67958e-08, 7.918068e-08, 8.161747e-08, 
    8.463911e-08, 8.716287e-08, 8.477808e-08, 8.541014e-08, 8.374597e-08, 
    8.238348e-08, 8.399219e-08, 7.918226e-08, 8.537617e-08,
  5.268643e-08, 5.332549e-08, 5.301494e-08, 5.345656e-08, 5.321332e-08, 
    5.529724e-08, 5.558365e-08, 5.716739e-08, 6.513332e-08, 6.721115e-08, 
    6.865317e-08, 6.761515e-08, 6.500849e-08, 5.999397e-08, 5.89395e-08, 
    5.938971e-08, 5.74234e-08, 5.601813e-08, 5.507842e-08, 5.425903e-08, 
    5.446489e-08, 5.2645e-08, 5.053703e-08, 5.003771e-08, 5.094567e-08, 
    5.103031e-08, 5.314554e-08, 5.3991e-08, 5.326854e-08,
  8.115665e-09, 8.495586e-09, 8.820596e-09, 8.067234e-09, 8.84397e-09, 
    8.53076e-09, 8.118392e-09, 8.060806e-09, 9.334833e-09, 1.126548e-08, 
    1.312455e-08, 1.361756e-08, 1.442363e-08, 1.235708e-08, 1.18123e-08, 
    1.158466e-08, 1.130823e-08, 1.027633e-08, 9.614576e-09, 9.168131e-09, 
    8.836755e-09, 9.47911e-09, 9.098391e-09, 8.70429e-09, 8.791576e-09, 
    8.361549e-09, 7.968401e-09, 7.647962e-09, 7.678038e-09,
  1.293215e-09, 1.100999e-09, 9.593719e-10, 1.094816e-09, 1.248342e-09, 
    1.392728e-09, 1.315517e-09, 1.053837e-09, 1.042328e-09, 8.969427e-10, 
    1.34333e-09, 1.585563e-09, 2.417399e-09, 1.653409e-09, 1.613856e-09, 
    1.272059e-09, 1.42057e-09, 1.683091e-09, 1.44279e-09, 1.374973e-09, 
    1.368715e-09, 1.473218e-09, 1.441802e-09, 1.409297e-09, 1.405153e-09, 
    1.322873e-09, 1.33233e-09, 1.380819e-09, 1.35907e-09,
  4.513595e-10, 3.784911e-10, 3.758575e-10, 3.546584e-10, 3.227359e-10, 
    3.711789e-10, 3.424527e-10, 2.467295e-10, 2.508486e-10, 4.240681e-10, 
    4.568054e-10, 4.582771e-10, 6.609315e-10, 7.176809e-10, 4.852561e-10, 
    2.810629e-10, 3.042631e-10, 3.001277e-10, 3.638003e-10, 3.722434e-10, 
    3.496844e-10, 4.145231e-10, 4.518349e-10, 5.155293e-10, 5.999147e-10, 
    7.237492e-10, 6.94063e-10, 5.409055e-10, 4.787171e-10,
  1.545019e-10, 1.795482e-10, 1.89775e-10, 1.403874e-10, 1.832157e-10, 
    1.422525e-10, 1.108418e-10, 1.296954e-10, 9.521594e-11, 7.917086e-11, 
    1.032608e-10, 1.799727e-10, 3.820566e-10, 3.449331e-10, 3.227397e-10, 
    2.943095e-10, 2.679804e-10, 2.973134e-10, 3.323294e-10, 3.487892e-10, 
    3.865395e-10, 4.272703e-10, 3.324106e-10, 2.128271e-10, 2.161562e-10, 
    2.282576e-10, 1.978048e-10, 1.548825e-10, 1.428374e-10,
  1.019494e-10, 9.162526e-11, 9.446207e-11, 8.483288e-11, 1.004004e-10, 
    8.418901e-11, 8.037897e-11, 6.048975e-11, 5.006606e-11, 4.042819e-11, 
    5.457139e-11, 6.951643e-11, 8.013294e-11, 1.440087e-10, 2.333514e-10, 
    2.748071e-10, 3.305016e-10, 3.740177e-10, 3.84836e-10, 3.734921e-10, 
    3.012306e-10, 1.35213e-10, 8.708968e-11, 8.276278e-11, 8.977074e-11, 
    5.683822e-11, 5.72529e-11, 1.019231e-10, 1.147242e-10,
  3.436915e-11, 4.048637e-11, 5.286548e-11, 5.920878e-11, 5.387439e-11, 
    3.183264e-11, 2.573189e-11, 2.163908e-11, 1.791997e-11, 1.578016e-11, 
    1.765796e-11, 3.077784e-11, 3.709277e-11, 3.794623e-11, 4.342923e-11, 
    5.549838e-11, 6.534449e-11, 7.128193e-11, 6.62361e-11, 4.849123e-11, 
    3.460588e-11, 2.645926e-11, 1.959025e-11, 2.253313e-11, 3.148614e-11, 
    3.130877e-11, 2.821073e-11, 2.800585e-11, 3.233328e-11,
  1.563455e-12, 1.563455e-12, 1.563455e-12, 1.563455e-12, 1.563455e-12, 
    1.563455e-12, 1.563455e-12, 1.66084e-12, 1.66084e-12, 1.66084e-12, 
    1.66084e-12, 1.66084e-12, 1.66084e-12, 1.66084e-12, 1.66483e-12, 
    1.66483e-12, 1.66483e-12, 1.66483e-12, 1.66483e-12, 1.66483e-12, 
    1.66483e-12, 1.57459e-12, 1.57459e-12, 1.57459e-12, 1.57459e-12, 
    1.57459e-12, 1.57459e-12, 1.57459e-12, 1.563455e-12,
  5.538631e-12, 5.603272e-12, 5.031783e-12, 4.878094e-12, 5.121185e-12, 
    5.412774e-12, 5.675141e-12, 6.435939e-12, 7.03605e-12, 6.40707e-12, 
    6.033363e-12, 6.022729e-12, 5.851243e-12, 5.861027e-12, 6.949911e-12, 
    8.112123e-12, 8.51532e-12, 8.697491e-12, 8.6019e-12, 7.603004e-12, 
    7.070935e-12, 7.234641e-12, 6.557448e-12, 6.041948e-12, 4.872599e-12, 
    3.680229e-12, 2.962811e-12, 3.290034e-12, 5.02178e-12,
  2.94849e-11, 2.885403e-11, 2.74583e-11, 2.899343e-11, 3.298332e-11, 
    4.102725e-11, 4.133491e-11, 3.637209e-11, 3.94216e-11, 4.358445e-11, 
    4.749976e-11, 6.09632e-11, 6.74354e-11, 7.29078e-11, 7.768499e-11, 
    7.907498e-11, 7.30788e-11, 7.017945e-11, 6.227906e-11, 5.121917e-11, 
    4.507849e-11, 3.356158e-11, 3.308572e-11, 3.212839e-11, 3.352479e-11, 
    3.426756e-11, 3.577544e-11, 3.668673e-11, 3.197477e-11,
  1.834633e-10, 1.74864e-10, 1.42529e-10, 1.519577e-10, 1.788342e-10, 
    2.16966e-10, 2.410691e-10, 2.594951e-10, 2.538705e-10, 2.293926e-10, 
    2.380122e-10, 2.641696e-10, 3.045767e-10, 3.930217e-10, 4.935363e-10, 
    5.662646e-10, 5.530847e-10, 5.232805e-10, 4.808448e-10, 4.545849e-10, 
    4.563188e-10, 4.012926e-10, 3.460598e-10, 2.932066e-10, 2.848252e-10, 
    2.589043e-10, 2.286312e-10, 2.224851e-10, 1.94621e-10,
  1.480341e-09, 1.571593e-09, 1.685835e-09, 1.916314e-09, 1.855601e-09, 
    1.867722e-09, 1.576496e-09, 1.402684e-09, 1.256154e-09, 1.284589e-09, 
    1.518998e-09, 1.557014e-09, 2.089299e-09, 2.609569e-09, 2.638565e-09, 
    2.485078e-09, 2.198453e-09, 2.015756e-09, 1.515511e-09, 9.108211e-10, 
    8.233312e-10, 1.133158e-09, 1.376104e-09, 1.679195e-09, 1.667172e-09, 
    1.758077e-09, 1.608521e-09, 1.415617e-09, 1.48229e-09,
  5.416106e-09, 5.424508e-09, 5.685867e-09, 6.257402e-09, 6.666592e-09, 
    6.454803e-09, 5.358625e-09, 5.74358e-09, 4.64067e-09, 4.898772e-09, 
    6.3085e-09, 6.161602e-09, 4.297012e-09, 3.643687e-09, 3.15829e-09, 
    2.877348e-09, 3.272064e-09, 3.589738e-09, 4.428961e-09, 5.091547e-09, 
    4.911795e-09, 5.137164e-09, 4.481068e-09, 4.716572e-09, 7.018381e-09, 
    9.096763e-09, 9.161417e-09, 7.944566e-09, 6.138225e-09,
  5.232252e-08, 5.015372e-08, 4.762578e-08, 4.596759e-08, 4.368191e-08, 
    4.358282e-08, 4.301681e-08, 4.347131e-08, 4.516345e-08, 4.487922e-08, 
    4.174936e-08, 3.907823e-08, 3.963276e-08, 3.923831e-08, 3.863325e-08, 
    3.985914e-08, 4.073129e-08, 4.287219e-08, 4.59508e-08, 4.76202e-08, 
    4.804671e-08, 4.887469e-08, 5.254284e-08, 5.776868e-08, 5.320778e-08, 
    4.889995e-08, 4.811055e-08, 4.949045e-08, 5.20627e-08,
  3.460206e-07, 3.336791e-07, 3.273543e-07, 3.316467e-07, 3.24985e-07, 
    3.215299e-07, 3.180564e-07, 3.175974e-07, 3.273857e-07, 3.311155e-07, 
    3.215519e-07, 3.050139e-07, 2.99946e-07, 3.007808e-07, 3.035636e-07, 
    3.027324e-07, 3.110922e-07, 3.156818e-07, 3.381594e-07, 3.496113e-07, 
    3.634979e-07, 3.722878e-07, 3.818948e-07, 3.8678e-07, 3.687521e-07, 
    3.610353e-07, 3.581872e-07, 3.695826e-07, 3.551185e-07,
  5.878754e-07, 5.694627e-07, 5.969791e-07, 6.148874e-07, 6.406078e-07, 
    6.223239e-07, 6.01408e-07, 5.641153e-07, 5.591247e-07, 5.404074e-07, 
    5.100835e-07, 4.721639e-07, 4.622493e-07, 4.333009e-07, 4.138313e-07, 
    4.232175e-07, 4.442009e-07, 4.785301e-07, 5.081304e-07, 5.540754e-07, 
    5.909712e-07, 6.074695e-07, 5.966841e-07, 6.010508e-07, 5.840137e-07, 
    5.942426e-07, 6.252106e-07, 6.357305e-07, 6.314755e-07,
  4.751791e-07, 4.587709e-07, 4.656575e-07, 4.702004e-07, 4.584979e-07, 
    4.93584e-07, 5.086085e-07, 5.06497e-07, 5.431917e-07, 5.883415e-07, 
    5.917977e-07, 6.079281e-07, 6.289455e-07, 6.676866e-07, 6.564599e-07, 
    6.392356e-07, 6.217732e-07, 5.593075e-07, 5.394102e-07, 4.719401e-07, 
    4.675548e-07, 4.835373e-07, 5.031808e-07, 4.732346e-07, 4.390544e-07, 
    4.371101e-07, 4.459702e-07, 4.854628e-07, 4.889584e-07,
  3.597288e-07, 3.592437e-07, 3.642167e-07, 3.732986e-07, 3.984692e-07, 
    3.959195e-07, 4.117908e-07, 4.27351e-07, 4.649878e-07, 4.676168e-07, 
    4.799255e-07, 4.526992e-07, 4.366105e-07, 4.460641e-07, 4.110859e-07, 
    3.801644e-07, 3.743828e-07, 3.525144e-07, 3.200462e-07, 3.243699e-07, 
    3.188537e-07, 3.21107e-07, 3.379581e-07, 3.450326e-07, 3.411369e-07, 
    3.413774e-07, 3.484916e-07, 3.454169e-07, 3.561436e-07,
  2.025331e-07, 2.05278e-07, 2.096866e-07, 2.093921e-07, 2.085832e-07, 
    2.07623e-07, 2.108904e-07, 2.267586e-07, 2.555073e-07, 2.54226e-07, 
    2.909765e-07, 2.871635e-07, 2.556941e-07, 2.47702e-07, 2.282086e-07, 
    2.336417e-07, 2.265465e-07, 2.250383e-07, 2.104992e-07, 2.02354e-07, 
    1.982696e-07, 1.965689e-07, 1.970257e-07, 1.974395e-07, 1.973862e-07, 
    1.932769e-07, 2.003153e-07, 2.065512e-07, 2.08469e-07,
  3.353867e-08, 3.672274e-08, 3.655388e-08, 3.640849e-08, 3.82066e-08, 
    3.378698e-08, 3.231452e-08, 3.277122e-08, 3.931801e-08, 4.483625e-08, 
    5.33665e-08, 6.153817e-08, 6.254218e-08, 5.503536e-08, 5.36285e-08, 
    5.019144e-08, 5.089286e-08, 4.477712e-08, 4.056786e-08, 3.804839e-08, 
    3.796816e-08, 3.75425e-08, 3.562236e-08, 3.718245e-08, 3.534618e-08, 
    3.432915e-08, 3.393997e-08, 3.235856e-08, 3.152592e-08,
  5.482669e-09, 5.135804e-09, 4.25716e-09, 4.103334e-09, 5.731208e-09, 
    5.568863e-09, 5.506914e-09, 4.248946e-09, 4.051519e-09, 3.591088e-09, 
    5.615093e-09, 7.521931e-09, 1.488139e-08, 1.013126e-08, 8.541583e-09, 
    6.474774e-09, 6.573012e-09, 7.120931e-09, 6.506248e-09, 5.770009e-09, 
    5.822431e-09, 5.72449e-09, 6.074748e-09, 6.231699e-09, 5.902764e-09, 
    5.563878e-09, 5.512136e-09, 5.911479e-09, 5.827614e-09,
  2.078047e-09, 1.660967e-09, 1.75414e-09, 1.41966e-09, 1.32997e-09, 
    1.7311e-09, 1.505335e-09, 1.091706e-09, 8.780632e-10, 1.348508e-09, 
    1.534592e-09, 1.568664e-09, 2.384923e-09, 3.308216e-09, 2.613856e-09, 
    1.468288e-09, 1.243211e-09, 1.338297e-09, 1.374603e-09, 1.544994e-09, 
    1.529609e-09, 1.755051e-09, 2.198856e-09, 1.966425e-09, 2.477424e-09, 
    3.116303e-09, 3.087598e-09, 2.897917e-09, 2.417827e-09,
  6.96053e-10, 8.216317e-10, 8.708869e-10, 8.597743e-10, 7.792142e-10, 
    6.045893e-10, 4.884247e-10, 5.302706e-10, 4.393449e-10, 3.4582e-10, 
    3.760892e-10, 7.906051e-10, 9.449377e-10, 1.162987e-09, 1.112827e-09, 
    1.264134e-09, 1.091643e-09, 1.235562e-09, 1.391585e-09, 1.654353e-09, 
    1.654072e-09, 1.929104e-09, 1.26773e-09, 1.07678e-09, 9.306226e-10, 
    9.379778e-10, 8.981472e-10, 6.900943e-10, 6.750346e-10,
  3.83684e-10, 3.603128e-10, 3.338293e-10, 3.740691e-10, 3.797993e-10, 
    4.293863e-10, 4.03456e-10, 3.427894e-10, 2.252024e-10, 1.702547e-10, 
    2.090869e-10, 2.706904e-10, 3.478475e-10, 5.69999e-10, 6.949899e-10, 
    1.059772e-09, 1.356586e-09, 1.376808e-09, 1.306161e-09, 1.281194e-09, 
    1.130925e-09, 6.140201e-10, 3.692205e-10, 3.004108e-10, 4.125829e-10, 
    2.697929e-10, 3.692814e-10, 5.289694e-10, 4.177766e-10,
  2.378921e-10, 3.243485e-10, 3.635907e-10, 3.558741e-10, 3.245706e-10, 
    2.597724e-10, 1.586289e-10, 1.063717e-10, 7.981141e-11, 7.568412e-11, 
    8.808936e-11, 1.357539e-10, 1.626378e-10, 1.848783e-10, 2.68137e-10, 
    3.220111e-10, 3.491736e-10, 3.622091e-10, 3.297539e-10, 2.199353e-10, 
    1.233327e-10, 9.732627e-11, 8.601446e-11, 1.108801e-10, 1.358468e-10, 
    1.307582e-10, 1.1894e-10, 1.38414e-10, 1.977597e-10,
  8.223117e-12, 8.223117e-12, 8.223117e-12, 8.223117e-12, 8.223117e-12, 
    8.223117e-12, 8.223117e-12, 8.599698e-12, 8.599698e-12, 8.599698e-12, 
    8.599698e-12, 8.599698e-12, 8.599698e-12, 8.599698e-12, 8.82966e-12, 
    8.82966e-12, 8.82966e-12, 8.82966e-12, 8.82966e-12, 8.82966e-12, 
    8.82966e-12, 8.528646e-12, 8.528646e-12, 8.528646e-12, 8.528646e-12, 
    8.528646e-12, 8.528646e-12, 8.528646e-12, 8.223117e-12,
  1.895778e-11, 2.092674e-11, 1.9508e-11, 1.904566e-11, 1.952548e-11, 
    2.033039e-11, 2.030101e-11, 2.076401e-11, 2.2779e-11, 2.180364e-11, 
    2.47601e-11, 2.586512e-11, 2.769675e-11, 2.765316e-11, 2.878587e-11, 
    3.501456e-11, 3.785275e-11, 3.811518e-11, 3.651258e-11, 3.701783e-11, 
    3.680952e-11, 3.559888e-11, 3.43222e-11, 3.163615e-11, 2.63864e-11, 
    2.030743e-11, 1.610411e-11, 1.450552e-11, 1.719083e-11,
  1.170561e-10, 1.057109e-10, 1.027678e-10, 1.106634e-10, 1.269147e-10, 
    1.433236e-10, 1.449695e-10, 1.324247e-10, 1.305515e-10, 1.391684e-10, 
    1.516603e-10, 1.823008e-10, 2.33745e-10, 2.784821e-10, 2.997492e-10, 
    3.133319e-10, 2.979016e-10, 2.879781e-10, 2.558278e-10, 2.14749e-10, 
    1.895472e-10, 1.616781e-10, 1.552669e-10, 1.546285e-10, 1.56006e-10, 
    1.58006e-10, 1.559885e-10, 1.520645e-10, 1.281625e-10,
  5.92708e-10, 5.577823e-10, 4.832998e-10, 5.504414e-10, 6.179406e-10, 
    6.901804e-10, 7.256862e-10, 8.002297e-10, 7.988462e-10, 8.182486e-10, 
    9.229014e-10, 1.169862e-09, 1.482569e-09, 1.777402e-09, 2.221625e-09, 
    2.413542e-09, 2.234136e-09, 1.987696e-09, 1.800631e-09, 1.593345e-09, 
    1.406595e-09, 1.253751e-09, 1.211878e-09, 1.161775e-09, 1.135707e-09, 
    1.049017e-09, 8.860417e-10, 7.764486e-10, 6.695396e-10,
  4.523127e-09, 4.767062e-09, 6.253611e-09, 6.627652e-09, 7.237356e-09, 
    8.045914e-09, 6.579822e-09, 5.332099e-09, 4.260313e-09, 5.185954e-09, 
    5.831585e-09, 5.598242e-09, 7.143343e-09, 8.095506e-09, 8.448927e-09, 
    8.257008e-09, 6.959529e-09, 6.186477e-09, 4.80353e-09, 3.341858e-09, 
    2.892582e-09, 4.187906e-09, 4.895216e-09, 5.994689e-09, 6.283603e-09, 
    6.272738e-09, 5.822698e-09, 4.406476e-09, 4.653734e-09,
  2.431481e-08, 2.108021e-08, 2.514644e-08, 2.559812e-08, 2.716471e-08, 
    2.543684e-08, 2.475008e-08, 2.250543e-08, 2.271083e-08, 2.095054e-08, 
    2.409206e-08, 2.29876e-08, 1.843146e-08, 1.632593e-08, 1.417886e-08, 
    1.218869e-08, 1.221885e-08, 1.360478e-08, 1.693574e-08, 1.929027e-08, 
    1.817044e-08, 2.010334e-08, 1.79038e-08, 1.771025e-08, 2.342155e-08, 
    3.229397e-08, 3.6384e-08, 3.290273e-08, 2.754112e-08,
  2.333601e-07, 2.201078e-07, 2.040803e-07, 2.004899e-07, 1.880392e-07, 
    1.815387e-07, 1.78474e-07, 1.701583e-07, 1.77777e-07, 1.73937e-07, 
    1.559457e-07, 1.518386e-07, 1.511278e-07, 1.50075e-07, 1.540367e-07, 
    1.652543e-07, 1.69951e-07, 1.818149e-07, 1.966044e-07, 2.007168e-07, 
    2.092034e-07, 2.131213e-07, 2.176452e-07, 2.291382e-07, 2.163395e-07, 
    2.088399e-07, 2.116425e-07, 2.249921e-07, 2.242202e-07,
  1.48367e-06, 1.401045e-06, 1.343319e-06, 1.275706e-06, 1.271086e-06, 
    1.271288e-06, 1.238208e-06, 1.279586e-06, 1.20883e-06, 1.207988e-06, 
    1.192934e-06, 1.163848e-06, 1.158762e-06, 1.1822e-06, 1.190256e-06, 
    1.195673e-06, 1.230372e-06, 1.29274e-06, 1.346631e-06, 1.412971e-06, 
    1.447516e-06, 1.525102e-06, 1.516628e-06, 1.535195e-06, 1.558945e-06, 
    1.546834e-06, 1.515636e-06, 1.462468e-06, 1.475922e-06,
  2.69833e-06, 2.497178e-06, 2.542426e-06, 2.648814e-06, 2.761229e-06, 
    2.934444e-06, 2.705329e-06, 2.507968e-06, 2.302506e-06, 2.304999e-06, 
    2.15105e-06, 1.9852e-06, 1.806326e-06, 1.691656e-06, 1.617868e-06, 
    1.596818e-06, 1.705879e-06, 1.890326e-06, 2.043718e-06, 2.185515e-06, 
    2.329414e-06, 2.466315e-06, 2.576465e-06, 2.548376e-06, 2.473009e-06, 
    2.471306e-06, 2.566739e-06, 2.673039e-06, 2.683461e-06,
  1.913795e-06, 1.900041e-06, 1.853585e-06, 1.889455e-06, 1.918085e-06, 
    1.884912e-06, 1.921826e-06, 2.020875e-06, 2.055966e-06, 2.136633e-06, 
    2.396969e-06, 2.583465e-06, 2.794008e-06, 2.830212e-06, 2.775758e-06, 
    2.940484e-06, 2.820122e-06, 2.609311e-06, 2.440188e-06, 2.172085e-06, 
    2.220083e-06, 2.191807e-06, 2.151811e-06, 2.003729e-06, 1.889894e-06, 
    1.892457e-06, 1.790008e-06, 1.838527e-06, 1.953138e-06,
  1.556175e-06, 1.553498e-06, 1.489852e-06, 1.494879e-06, 1.56968e-06, 
    1.649045e-06, 1.609999e-06, 1.718304e-06, 1.824587e-06, 1.982787e-06, 
    2.065287e-06, 2.074531e-06, 1.998229e-06, 1.887849e-06, 1.655109e-06, 
    1.55214e-06, 1.489234e-06, 1.40766e-06, 1.330301e-06, 1.331429e-06, 
    1.40627e-06, 1.429438e-06, 1.406634e-06, 1.416105e-06, 1.391836e-06, 
    1.438686e-06, 1.431745e-06, 1.435867e-06, 1.486746e-06,
  8.727992e-07, 8.47229e-07, 8.054665e-07, 8.260816e-07, 8.301193e-07, 
    8.425232e-07, 8.879742e-07, 9.930777e-07, 1.031946e-06, 1.1871e-06, 
    1.292564e-06, 1.167017e-06, 1.063106e-06, 9.652699e-07, 9.02814e-07, 
    8.586288e-07, 8.403833e-07, 8.592946e-07, 8.695337e-07, 8.672521e-07, 
    8.602383e-07, 8.322939e-07, 8.019817e-07, 7.993902e-07, 8.203556e-07, 
    8.224588e-07, 8.605519e-07, 8.465807e-07, 8.698394e-07,
  1.626463e-07, 1.808328e-07, 1.759553e-07, 1.834895e-07, 1.735281e-07, 
    1.541576e-07, 1.40775e-07, 1.406736e-07, 1.728634e-07, 1.88625e-07, 
    2.168323e-07, 2.618719e-07, 3.105295e-07, 2.6364e-07, 2.491752e-07, 
    2.314517e-07, 2.203898e-07, 2.006663e-07, 1.741256e-07, 1.632446e-07, 
    1.579139e-07, 1.633836e-07, 1.648168e-07, 1.687249e-07, 1.722839e-07, 
    1.626611e-07, 1.546747e-07, 1.54649e-07, 1.540928e-07,
  2.87449e-08, 2.588516e-08, 2.165998e-08, 2.334363e-08, 2.622411e-08, 
    2.053142e-08, 2.251631e-08, 1.907258e-08, 1.758756e-08, 1.702262e-08, 
    2.400155e-08, 3.458359e-08, 7.664228e-08, 6.320077e-08, 5.331684e-08, 
    3.860271e-08, 2.940785e-08, 2.939597e-08, 2.875714e-08, 2.549471e-08, 
    2.666273e-08, 2.731467e-08, 2.832678e-08, 2.94584e-08, 2.864256e-08, 
    2.748899e-08, 2.652111e-08, 2.932244e-08, 3.22299e-08,
  9.509065e-09, 8.379441e-09, 7.52275e-09, 6.093382e-09, 5.899473e-09, 
    8.510816e-09, 7.682184e-09, 5.667962e-09, 3.54709e-09, 4.738599e-09, 
    6.974717e-09, 6.625948e-09, 8.172272e-09, 1.525593e-08, 1.347508e-08, 
    9.385033e-09, 6.071499e-09, 5.565849e-09, 6.180431e-09, 6.368699e-09, 
    7.360828e-09, 8.93621e-09, 1.031193e-08, 8.762373e-09, 1.071431e-08, 
    1.124749e-08, 1.030507e-08, 1.106687e-08, 9.977013e-09,
  3.364856e-09, 3.701566e-09, 3.938756e-09, 4.549663e-09, 3.621563e-09, 
    2.982321e-09, 2.102318e-09, 1.902629e-09, 1.569155e-09, 1.75811e-09, 
    1.374918e-09, 2.462275e-09, 2.726493e-09, 3.883608e-09, 4.608207e-09, 
    5.505132e-09, 6.687851e-09, 6.418429e-09, 5.897722e-09, 6.81306e-09, 
    8.368601e-09, 7.88082e-09, 5.396184e-09, 5.265567e-09, 4.104116e-09, 
    3.779415e-09, 4.250255e-09, 3.545176e-09, 3.268689e-09,
  2.091469e-09, 1.538576e-09, 1.356176e-09, 1.399998e-09, 1.821068e-09, 
    2.048168e-09, 1.687673e-09, 1.353729e-09, 1.044549e-09, 7.595547e-10, 
    8.248714e-10, 1.189351e-09, 1.464697e-09, 2.149205e-09, 3.543053e-09, 
    4.47687e-09, 5.911736e-09, 6.507923e-09, 4.940848e-09, 5.227931e-09, 
    4.550709e-09, 2.943828e-09, 1.486456e-09, 1.135156e-09, 1.618623e-09, 
    1.317011e-09, 1.900785e-09, 2.303849e-09, 2.333227e-09,
  1.216238e-09, 1.334828e-09, 1.379464e-09, 1.466927e-09, 1.610349e-09, 
    1.305056e-09, 9.131501e-10, 6.475035e-10, 4.026801e-10, 3.367152e-10, 
    3.770511e-10, 5.438309e-10, 6.516928e-10, 9.778667e-10, 1.324255e-09, 
    1.541386e-09, 1.657899e-09, 1.673117e-09, 1.490996e-09, 1.011893e-09, 
    5.128185e-10, 3.73327e-10, 3.680481e-10, 5.252777e-10, 5.680247e-10, 
    4.590925e-10, 4.798492e-10, 5.983125e-10, 1.051936e-09,
  5.810028e-11, 5.810028e-11, 5.810028e-11, 5.810028e-11, 5.810028e-11, 
    5.810028e-11, 5.810028e-11, 5.998692e-11, 5.998692e-11, 5.998692e-11, 
    5.998692e-11, 5.998692e-11, 5.998692e-11, 5.998692e-11, 5.744665e-11, 
    5.744665e-11, 5.744665e-11, 5.744665e-11, 5.744665e-11, 5.744665e-11, 
    5.744665e-11, 5.58125e-11, 5.58125e-11, 5.58125e-11, 5.58125e-11, 
    5.58125e-11, 5.58125e-11, 5.58125e-11, 5.810028e-11,
  7.823552e-11, 9.149771e-11, 8.949004e-11, 8.83988e-11, 9.329554e-11, 
    9.505625e-11, 9.570111e-11, 9.975876e-11, 1.079457e-10, 1.081321e-10, 
    1.442614e-10, 1.560022e-10, 1.503889e-10, 1.47638e-10, 1.412979e-10, 
    1.418716e-10, 1.582414e-10, 1.777213e-10, 1.881681e-10, 1.914295e-10, 
    1.992487e-10, 1.986157e-10, 1.764312e-10, 1.549048e-10, 1.242592e-10, 
    1.089553e-10, 8.780212e-11, 7.349578e-11, 7.197074e-11,
  4.832629e-10, 4.304589e-10, 4.127027e-10, 4.310184e-10, 4.851611e-10, 
    5.187501e-10, 5.093568e-10, 4.690273e-10, 4.493635e-10, 4.644418e-10, 
    5.320794e-10, 6.326e-10, 8.033436e-10, 1.104175e-09, 1.348512e-09, 
    1.363839e-09, 1.372401e-09, 1.243918e-09, 1.165539e-09, 1.07398e-09, 
    9.598052e-10, 8.337397e-10, 7.873914e-10, 7.65813e-10, 7.767594e-10, 
    7.227041e-10, 6.933423e-10, 6.501515e-10, 5.430337e-10,
  2.411029e-09, 2.205357e-09, 2.156202e-09, 2.241603e-09, 2.496418e-09, 
    2.64376e-09, 2.745688e-09, 2.781573e-09, 2.939229e-09, 2.980151e-09, 
    3.315788e-09, 5.169135e-09, 7.041005e-09, 8.815596e-09, 9.773561e-09, 
    9.780991e-09, 8.656533e-09, 7.661085e-09, 6.953595e-09, 6.182812e-09, 
    5.269448e-09, 4.310558e-09, 4.438298e-09, 4.694755e-09, 4.745184e-09, 
    4.591298e-09, 3.952164e-09, 3.211914e-09, 2.758641e-09,
  1.531255e-08, 1.714136e-08, 2.189658e-08, 2.358657e-08, 2.784144e-08, 
    3.394284e-08, 2.869868e-08, 1.939013e-08, 1.621518e-08, 1.760983e-08, 
    2.277827e-08, 2.726433e-08, 3.188529e-08, 3.125122e-08, 3.301077e-08, 
    3.219147e-08, 2.59914e-08, 2.076651e-08, 1.62454e-08, 1.313628e-08, 
    1.195675e-08, 1.614645e-08, 1.88881e-08, 2.439189e-08, 2.419597e-08, 
    2.317577e-08, 2.167332e-08, 1.646904e-08, 1.545397e-08,
  1.111926e-07, 1.013387e-07, 1.054089e-07, 1.145725e-07, 1.112794e-07, 
    1.11339e-07, 1.075059e-07, 1.142008e-07, 1.082802e-07, 1.157194e-07, 
    1.158441e-07, 1.108259e-07, 9.521094e-08, 8.440916e-08, 7.191781e-08, 
    5.859752e-08, 4.813966e-08, 5.351563e-08, 7.402096e-08, 7.517377e-08, 
    8.269451e-08, 9.254442e-08, 7.79327e-08, 7.483658e-08, 9.576111e-08, 
    1.098413e-07, 1.434457e-07, 1.466983e-07, 1.186168e-07,
  1.045195e-06, 1.020212e-06, 9.420758e-07, 8.955344e-07, 8.477242e-07, 
    8.239416e-07, 7.990819e-07, 7.943455e-07, 7.605333e-07, 7.189111e-07, 
    6.650853e-07, 6.118008e-07, 6.11911e-07, 6.13505e-07, 6.179367e-07, 
    6.466533e-07, 6.802838e-07, 7.619432e-07, 8.192798e-07, 8.796427e-07, 
    9.087864e-07, 9.240515e-07, 9.609697e-07, 1.005381e-06, 9.452179e-07, 
    9.197857e-07, 9.590891e-07, 1.02779e-06, 1.061418e-06,
  6.14431e-06, 5.844502e-06, 5.793006e-06, 5.739106e-06, 5.327875e-06, 
    5.318311e-06, 4.916329e-06, 4.762975e-06, 4.781446e-06, 4.519713e-06, 
    4.423262e-06, 4.284873e-06, 4.428279e-06, 4.498702e-06, 4.538321e-06, 
    4.80888e-06, 5.086486e-06, 5.40868e-06, 5.805322e-06, 6.103283e-06, 
    6.553629e-06, 6.675169e-06, 6.714442e-06, 6.355761e-06, 6.314007e-06, 
    6.24201e-06, 6.462526e-06, 6.619451e-06, 6.441966e-06,
  1.06515e-05, 1.030565e-05, 1.04122e-05, 1.125006e-05, 1.19127e-05, 
    1.19557e-05, 1.205456e-05, 1.161634e-05, 1.135643e-05, 1.005527e-05, 
    9.340372e-06, 8.29539e-06, 7.500297e-06, 6.55622e-06, 6.178297e-06, 
    6.235854e-06, 6.454262e-06, 7.09597e-06, 7.92908e-06, 8.777221e-06, 
    9.980134e-06, 1.031829e-05, 1.028579e-05, 1.02033e-05, 1.006685e-05, 
    1.034126e-05, 1.079161e-05, 1.148149e-05, 1.162063e-05,
  7.461611e-06, 7.445995e-06, 7.539083e-06, 7.772003e-06, 7.827238e-06, 
    7.618985e-06, 7.919864e-06, 8.056675e-06, 8.432617e-06, 9.387727e-06, 
    1.000565e-05, 1.070813e-05, 1.083694e-05, 1.164249e-05, 1.275602e-05, 
    1.207322e-05, 1.152019e-05, 1.097816e-05, 1.082361e-05, 1.105697e-05, 
    1.046815e-05, 9.69802e-06, 8.999683e-06, 8.63925e-06, 7.745987e-06, 
    7.555089e-06, 7.39796e-06, 7.503056e-06, 7.339205e-06,
  6.70073e-06, 6.671669e-06, 6.754452e-06, 6.494977e-06, 6.87663e-06, 
    6.829722e-06, 6.934072e-06, 7.151632e-06, 7.525512e-06, 8.012775e-06, 
    8.987804e-06, 9.210495e-06, 8.919317e-06, 8.062198e-06, 7.163284e-06, 
    6.534609e-06, 5.994537e-06, 5.679438e-06, 5.285624e-06, 5.316531e-06, 
    5.387057e-06, 5.760204e-06, 5.930009e-06, 5.947392e-06, 5.884985e-06, 
    6.199218e-06, 6.369042e-06, 6.432301e-06, 6.890206e-06,
  4.031212e-06, 3.841898e-06, 3.669024e-06, 3.762312e-06, 3.518611e-06, 
    3.580028e-06, 4.054243e-06, 3.982317e-06, 4.283046e-06, 5.289298e-06, 
    6.082552e-06, 6.067934e-06, 4.976055e-06, 4.145724e-06, 3.907363e-06, 
    3.620868e-06, 3.702306e-06, 3.664313e-06, 3.522603e-06, 3.487674e-06, 
    3.565414e-06, 3.621978e-06, 3.660256e-06, 3.639706e-06, 3.63211e-06, 
    3.748294e-06, 3.889284e-06, 4.060311e-06, 4.060631e-06,
  8.541641e-07, 8.77076e-07, 8.653416e-07, 9.715751e-07, 7.757178e-07, 
    6.706263e-07, 6.39234e-07, 6.180284e-07, 6.539317e-07, 6.935003e-07, 
    9.156172e-07, 1.228134e-06, 1.467903e-06, 1.372818e-06, 1.145845e-06, 
    1.099599e-06, 9.408835e-07, 8.731437e-07, 7.893339e-07, 7.608357e-07, 
    7.459763e-07, 7.572979e-07, 7.546055e-07, 8.409235e-07, 8.630684e-07, 
    8.541059e-07, 8.165208e-07, 8.139051e-07, 8.09012e-07,
  1.611267e-07, 1.512989e-07, 1.35263e-07, 1.319803e-07, 1.335924e-07, 
    9.462519e-08, 8.373532e-08, 8.191648e-08, 7.544897e-08, 7.597905e-08, 
    1.003456e-07, 1.512803e-07, 3.354101e-07, 3.33433e-07, 2.988596e-07, 
    2.445857e-07, 1.803174e-07, 1.337748e-07, 1.300963e-07, 1.142811e-07, 
    1.171704e-07, 1.216703e-07, 1.286283e-07, 1.409222e-07, 1.376861e-07, 
    1.396599e-07, 1.405412e-07, 1.533732e-07, 1.783344e-07,
  4.40129e-08, 4.290805e-08, 3.736977e-08, 2.73538e-08, 2.767922e-08, 
    3.608939e-08, 3.481628e-08, 2.684423e-08, 1.712974e-08, 1.922423e-08, 
    3.060348e-08, 2.834182e-08, 3.498375e-08, 6.555123e-08, 5.935229e-08, 
    4.450794e-08, 3.03661e-08, 2.662168e-08, 2.699667e-08, 3.118285e-08, 
    3.222638e-08, 4.099575e-08, 4.616674e-08, 3.772403e-08, 4.365905e-08, 
    4.636648e-08, 4.626047e-08, 4.950574e-08, 4.475103e-08,
  1.671631e-08, 1.854426e-08, 1.941739e-08, 2.090884e-08, 1.469856e-08, 
    1.13005e-08, 8.191597e-09, 7.545564e-09, 6.444866e-09, 5.807499e-09, 
    5.209057e-09, 1.020599e-08, 1.282121e-08, 2.210686e-08, 2.0503e-08, 
    2.464815e-08, 3.482129e-08, 3.028423e-08, 2.581524e-08, 2.672097e-08, 
    3.264795e-08, 3.311032e-08, 2.225183e-08, 2.31658e-08, 1.924095e-08, 
    1.556278e-08, 2.057628e-08, 2.12547e-08, 1.754095e-08,
  1.078114e-08, 8.613658e-09, 5.408824e-09, 5.521498e-09, 7.499574e-09, 
    7.746837e-09, 7.608217e-09, 5.723884e-09, 4.838265e-09, 3.453247e-09, 
    3.361381e-09, 4.992631e-09, 5.998891e-09, 1.212939e-08, 1.501664e-08, 
    1.580763e-08, 2.066471e-08, 2.859043e-08, 2.674972e-08, 2.29116e-08, 
    2.114007e-08, 1.315528e-08, 5.850914e-09, 3.811884e-09, 5.807184e-09, 
    6.538186e-09, 9.269908e-09, 1.286297e-08, 1.16413e-08,
  4.786045e-09, 4.736517e-09, 4.798391e-09, 5.153353e-09, 6.246551e-09, 
    5.968055e-09, 4.390238e-09, 3.494858e-09, 2.347199e-09, 1.62815e-09, 
    1.487542e-09, 1.638111e-09, 2.405488e-09, 3.89035e-09, 5.294324e-09, 
    6.281109e-09, 6.591e-09, 6.415067e-09, 5.669142e-09, 3.749395e-09, 
    2.190763e-09, 1.306509e-09, 1.375074e-09, 2.143099e-09, 2.587299e-09, 
    2.150539e-09, 2.082698e-09, 2.972176e-09, 4.502559e-09,
  3.209372e-10, 3.209372e-10, 3.209372e-10, 3.209372e-10, 3.209372e-10, 
    3.209372e-10, 3.209372e-10, 3.261481e-10, 3.261481e-10, 3.261481e-10, 
    3.261481e-10, 3.261481e-10, 3.261481e-10, 3.261481e-10, 3.284654e-10, 
    3.284654e-10, 3.284654e-10, 3.284654e-10, 3.284654e-10, 3.284654e-10, 
    3.284654e-10, 3.29559e-10, 3.29559e-10, 3.29559e-10, 3.29559e-10, 
    3.29559e-10, 3.29559e-10, 3.29559e-10, 3.209372e-10,
  4.049505e-10, 4.375319e-10, 4.786965e-10, 4.851897e-10, 5.055883e-10, 
    5.182114e-10, 5.047731e-10, 4.98992e-10, 4.946856e-10, 4.900276e-10, 
    6.695688e-10, 7.210867e-10, 7.134735e-10, 7.374039e-10, 7.639646e-10, 
    7.846966e-10, 7.787816e-10, 8.247154e-10, 8.343214e-10, 8.553997e-10, 
    9.008768e-10, 8.938811e-10, 8.135354e-10, 7.592964e-10, 6.929487e-10, 
    6.309229e-10, 5.686361e-10, 4.789466e-10, 4.133363e-10,
  1.955055e-09, 1.727914e-09, 1.633175e-09, 1.752491e-09, 1.924999e-09, 
    1.943208e-09, 1.78643e-09, 1.66849e-09, 1.612692e-09, 1.674385e-09, 
    1.711047e-09, 2.237549e-09, 2.957836e-09, 4.579811e-09, 5.843841e-09, 
    6.285123e-09, 6.335291e-09, 5.935565e-09, 5.500344e-09, 5.044405e-09, 
    4.236749e-09, 3.676612e-09, 3.631366e-09, 3.576842e-09, 3.719609e-09, 
    3.44715e-09, 3.287086e-09, 2.956225e-09, 2.229868e-09,
  1.015515e-08, 8.422775e-09, 8.832495e-09, 9.830702e-09, 1.088922e-08, 
    1.182724e-08, 1.127244e-08, 1.06702e-08, 1.181839e-08, 1.321817e-08, 
    1.255315e-08, 2.115541e-08, 3.180921e-08, 4.30124e-08, 4.834619e-08, 
    4.305746e-08, 3.553878e-08, 3.106338e-08, 2.826638e-08, 2.405713e-08, 
    2.101577e-08, 1.88149e-08, 1.915037e-08, 1.941265e-08, 2.185011e-08, 
    2.120815e-08, 1.778449e-08, 1.534051e-08, 1.251082e-08,
  5.920394e-08, 6.801505e-08, 8.457007e-08, 9.169326e-08, 1.100182e-07, 
    1.355125e-07, 1.288909e-07, 8.559226e-08, 6.650228e-08, 6.44151e-08, 
    9.724295e-08, 1.244908e-07, 1.553955e-07, 1.444978e-07, 1.492144e-07, 
    1.508857e-07, 1.169105e-07, 8.370024e-08, 6.624904e-08, 5.342791e-08, 
    4.956317e-08, 6.211094e-08, 7.088319e-08, 9.782153e-08, 1.064238e-07, 
    9.746881e-08, 8.545561e-08, 7.000673e-08, 5.729065e-08,
  5.974302e-07, 5.510254e-07, 4.987314e-07, 5.233397e-07, 5.486809e-07, 
    5.211804e-07, 4.442753e-07, 4.536016e-07, 6.286127e-07, 6.391419e-07, 
    6.812277e-07, 5.994946e-07, 5.769929e-07, 4.703777e-07, 3.898523e-07, 
    3.146934e-07, 2.270343e-07, 2.312471e-07, 3.056482e-07, 3.241413e-07, 
    3.501175e-07, 4.70218e-07, 4.14853e-07, 3.775234e-07, 4.267105e-07, 
    3.801155e-07, 4.373826e-07, 6.135667e-07, 6.350223e-07,
  4.911429e-06, 4.791599e-06, 4.642823e-06, 4.749412e-06, 4.512139e-06, 
    4.24218e-06, 4.128517e-06, 3.88686e-06, 3.839757e-06, 3.410728e-06, 
    3.004713e-06, 2.555899e-06, 2.360759e-06, 2.276121e-06, 2.382883e-06, 
    2.688885e-06, 3.001481e-06, 3.35018e-06, 3.803506e-06, 3.986931e-06, 
    4.112427e-06, 4.08228e-06, 4.229155e-06, 4.676304e-06, 4.66345e-06, 
    4.666849e-06, 4.353222e-06, 4.462806e-06, 4.795945e-06,
  2.989994e-05, 2.878631e-05, 2.63433e-05, 2.524346e-05, 2.53065e-05, 
    2.403797e-05, 2.265658e-05, 2.088005e-05, 1.93314e-05, 1.825923e-05, 
    1.763596e-05, 1.804123e-05, 1.73753e-05, 1.747367e-05, 1.754319e-05, 
    1.808124e-05, 1.957507e-05, 2.091185e-05, 2.321812e-05, 2.505058e-05, 
    2.66192e-05, 2.733413e-05, 2.747223e-05, 2.768234e-05, 2.851204e-05, 
    2.885173e-05, 2.907607e-05, 2.919669e-05, 3.015943e-05,
  5.099401e-05, 4.731012e-05, 4.494853e-05, 4.814104e-05, 5.172318e-05, 
    5.739157e-05, 5.408258e-05, 5.350114e-05, 5.072773e-05, 4.724196e-05, 
    4.016409e-05, 3.710046e-05, 3.18029e-05, 2.753072e-05, 2.535962e-05, 
    2.424088e-05, 2.456552e-05, 2.684691e-05, 3.080988e-05, 3.395385e-05, 
    3.867225e-05, 4.354687e-05, 4.613653e-05, 4.379265e-05, 4.038955e-05, 
    4.074047e-05, 4.528544e-05, 4.870749e-05, 5.174649e-05,
  2.899924e-05, 3.011688e-05, 3.158509e-05, 3.059216e-05, 3.188918e-05, 
    3.301176e-05, 3.276904e-05, 3.407485e-05, 3.723054e-05, 3.994324e-05, 
    4.526719e-05, 5.117871e-05, 5.726362e-05, 5.97627e-05, 6.251017e-05, 
    5.831606e-05, 5.774197e-05, 5.37231e-05, 4.944509e-05, 4.47823e-05, 
    3.974887e-05, 3.71124e-05, 3.300006e-05, 3.097395e-05, 3.059249e-05, 
    2.974556e-05, 2.91934e-05, 2.847415e-05, 2.851483e-05,
  3.092983e-05, 3.018324e-05, 3.0659e-05, 3.142262e-05, 2.990459e-05, 
    2.911128e-05, 3.153261e-05, 3.294004e-05, 3.243589e-05, 3.546273e-05, 
    4.063708e-05, 4.159606e-05, 3.875614e-05, 3.49955e-05, 2.979408e-05, 
    2.64668e-05, 2.508775e-05, 2.482358e-05, 2.36095e-05, 2.30788e-05, 
    2.373338e-05, 2.46818e-05, 2.493404e-05, 2.359203e-05, 2.445004e-05, 
    2.548069e-05, 2.758136e-05, 2.85003e-05, 3.071863e-05,
  1.889859e-05, 1.759226e-05, 1.71135e-05, 1.668236e-05, 1.586421e-05, 
    1.551601e-05, 1.850656e-05, 1.797077e-05, 1.830214e-05, 2.132117e-05, 
    2.757634e-05, 2.60968e-05, 2.218881e-05, 1.906662e-05, 1.729015e-05, 
    1.590112e-05, 1.626244e-05, 1.634319e-05, 1.673999e-05, 1.657168e-05, 
    1.6663e-05, 1.647706e-05, 1.573376e-05, 1.580072e-05, 1.635366e-05, 
    1.685933e-05, 1.758921e-05, 1.838666e-05, 1.876491e-05,
  4.695508e-06, 4.89482e-06, 5.208678e-06, 4.632228e-06, 4.249617e-06, 
    4.203805e-06, 3.503697e-06, 2.995436e-06, 2.799429e-06, 3.11086e-06, 
    3.829375e-06, 5.305595e-06, 8.024802e-06, 6.754119e-06, 5.229274e-06, 
    4.87741e-06, 4.257428e-06, 4.014629e-06, 3.63702e-06, 3.369151e-06, 
    3.306928e-06, 3.542454e-06, 3.687023e-06, 3.850695e-06, 4.140961e-06, 
    4.182899e-06, 4.232007e-06, 4.454411e-06, 4.603095e-06,
  1.0105e-06, 8.541638e-07, 8.481605e-07, 7.752534e-07, 7.162012e-07, 
    6.004105e-07, 4.623107e-07, 4.375614e-07, 3.760665e-07, 3.604088e-07, 
    4.103162e-07, 6.768623e-07, 1.295694e-06, 1.731597e-06, 1.630613e-06, 
    1.197468e-06, 1.024811e-06, 7.353818e-07, 6.632559e-07, 5.490962e-07, 
    4.77507e-07, 4.645999e-07, 5.127433e-07, 6.090331e-07, 6.604623e-07, 
    6.988303e-07, 7.523257e-07, 8.290899e-07, 1.063627e-06,
  2.147723e-07, 1.931725e-07, 1.709656e-07, 1.442277e-07, 1.264604e-07, 
    1.451927e-07, 1.361423e-07, 1.239342e-07, 8.403303e-08, 8.810836e-08, 
    1.284106e-07, 1.337931e-07, 1.773561e-07, 2.802991e-07, 2.766452e-07, 
    2.810931e-07, 2.291373e-07, 1.618477e-07, 1.198599e-07, 1.427091e-07, 
    1.394924e-07, 1.498731e-07, 1.778063e-07, 1.569989e-07, 1.631621e-07, 
    1.902923e-07, 2.058988e-07, 2.298124e-07, 2.124643e-07,
  8.40899e-08, 8.811242e-08, 9.295505e-08, 9.449151e-08, 6.402753e-08, 
    4.302232e-08, 3.111485e-08, 2.722387e-08, 2.532599e-08, 2.265549e-08, 
    2.050898e-08, 4.818798e-08, 5.944764e-08, 1.066305e-07, 9.661105e-08, 
    1.099303e-07, 1.468596e-07, 1.337931e-07, 1.084933e-07, 1.065731e-07, 
    1.068106e-07, 1.120409e-07, 8.773235e-08, 8.687407e-08, 8.199378e-08, 
    7.335635e-08, 9.860812e-08, 1.126421e-07, 8.401072e-08,
  3.687936e-08, 3.439335e-08, 2.880236e-08, 2.097145e-08, 2.83402e-08, 
    3.021398e-08, 2.86692e-08, 2.184847e-08, 1.751366e-08, 1.429572e-08, 
    1.290819e-08, 1.873512e-08, 2.569118e-08, 6.660826e-08, 4.785407e-08, 
    5.465798e-08, 6.497918e-08, 1.054918e-07, 1.282709e-07, 8.206685e-08, 
    7.394623e-08, 4.627768e-08, 2.543069e-08, 1.370433e-08, 2.275258e-08, 
    3.11582e-08, 4.91703e-08, 5.087145e-08, 4.049512e-08,
  1.947252e-08, 1.951162e-08, 1.953264e-08, 1.890451e-08, 2.122684e-08, 
    2.166263e-08, 2.16283e-08, 2.180125e-08, 1.582563e-08, 9.863963e-09, 
    6.55107e-09, 6.902968e-09, 9.544635e-09, 1.480353e-08, 2.174522e-08, 
    2.7698e-08, 2.689406e-08, 2.372181e-08, 2.000457e-08, 1.284163e-08, 
    7.778065e-09, 5.069658e-09, 5.120531e-09, 7.822724e-09, 9.889765e-09, 
    9.059365e-09, 8.663013e-09, 1.626331e-08, 1.927224e-08,
  1.591832e-09, 1.591832e-09, 1.591832e-09, 1.591832e-09, 1.591832e-09, 
    1.591832e-09, 1.591832e-09, 1.590417e-09, 1.590417e-09, 1.590417e-09, 
    1.590417e-09, 1.590417e-09, 1.590417e-09, 1.590417e-09, 1.820406e-09, 
    1.820406e-09, 1.820406e-09, 1.820406e-09, 1.820406e-09, 1.820406e-09, 
    1.820406e-09, 1.810847e-09, 1.810847e-09, 1.810847e-09, 1.810847e-09, 
    1.810847e-09, 1.810847e-09, 1.810847e-09, 1.591832e-09,
  2.469798e-09, 2.333356e-09, 2.504216e-09, 2.745518e-09, 2.854252e-09, 
    2.884201e-09, 2.857905e-09, 2.713711e-09, 2.451695e-09, 2.305596e-09, 
    2.411704e-09, 2.382549e-09, 2.726496e-09, 3.3224e-09, 3.814172e-09, 
    4.431198e-09, 4.30926e-09, 4.17706e-09, 3.377117e-09, 3.394156e-09, 
    3.553983e-09, 3.705733e-09, 3.804654e-09, 3.872309e-09, 3.641971e-09, 
    3.502376e-09, 3.090344e-09, 2.741141e-09, 2.565581e-09,
  7.623957e-09, 6.86328e-09, 6.582759e-09, 7.098813e-09, 8.285334e-09, 
    8.424339e-09, 7.24779e-09, 6.254777e-09, 5.929377e-09, 6.338414e-09, 
    6.051086e-09, 6.909109e-09, 1.051895e-08, 1.425924e-08, 2.360103e-08, 
    2.710273e-08, 2.775761e-08, 2.671559e-08, 2.368456e-08, 2.056339e-08, 
    1.727114e-08, 1.590526e-08, 1.556756e-08, 1.565965e-08, 1.661349e-08, 
    1.642777e-08, 1.493944e-08, 1.335464e-08, 8.664582e-09,
  4.396214e-08, 3.931298e-08, 3.738572e-08, 4.275836e-08, 4.685668e-08, 
    5.327938e-08, 5.168902e-08, 4.786973e-08, 5.217489e-08, 6.168298e-08, 
    5.536086e-08, 7.148822e-08, 1.35364e-07, 2.007889e-07, 2.357494e-07, 
    1.964002e-07, 1.618509e-07, 1.347977e-07, 1.160239e-07, 9.419392e-08, 
    8.425452e-08, 7.958889e-08, 8.317898e-08, 9.35977e-08, 1.091394e-07, 
    1.057931e-07, 8.882864e-08, 7.362106e-08, 5.622457e-08,
  2.500911e-07, 2.698498e-07, 3.408317e-07, 3.692444e-07, 4.748312e-07, 
    5.818593e-07, 5.902101e-07, 4.175349e-07, 3.019314e-07, 2.666905e-07, 
    3.971539e-07, 5.391967e-07, 6.86333e-07, 7.929603e-07, 6.979948e-07, 
    8.081992e-07, 5.854918e-07, 4.142772e-07, 2.803406e-07, 2.407126e-07, 
    2.290307e-07, 2.68058e-07, 2.897911e-07, 4.00705e-07, 4.694496e-07, 
    4.605317e-07, 3.996956e-07, 3.057083e-07, 2.459256e-07,
  3.148722e-06, 3.13503e-06, 2.999835e-06, 2.216849e-06, 2.360201e-06, 
    2.812377e-06, 2.323417e-06, 1.881974e-06, 2.667728e-06, 3.479667e-06, 
    3.570067e-06, 3.273125e-06, 3.329512e-06, 2.69237e-06, 2.568097e-06, 
    1.820434e-06, 1.28191e-06, 1.077066e-06, 1.252256e-06, 1.389177e-06, 
    1.318767e-06, 2.137515e-06, 2.222404e-06, 1.919555e-06, 2.001897e-06, 
    1.689082e-06, 1.573977e-06, 2.293052e-06, 2.758565e-06,
  2.460174e-05, 2.477595e-05, 2.411167e-05, 2.370335e-05, 2.382526e-05, 
    2.428704e-05, 2.472428e-05, 2.370588e-05, 2.102531e-05, 1.999348e-05, 
    1.724736e-05, 1.370243e-05, 1.067715e-05, 9.36924e-06, 8.489313e-06, 
    9.290254e-06, 1.172171e-05, 1.458424e-05, 1.640181e-05, 1.779102e-05, 
    1.844178e-05, 1.811588e-05, 1.862295e-05, 2.031e-05, 2.008365e-05, 
    2.053182e-05, 2.209353e-05, 2.25043e-05, 2.39131e-05,
  0.000136254, 0.0001398843, 0.000138687, 0.0001274261, 0.0001217752, 
    0.0001182988, 0.0001080613, 9.743594e-05, 8.897957e-05, 7.852629e-05, 
    6.607208e-05, 6.198644e-05, 6.302857e-05, 6.728829e-05, 7.038261e-05, 
    7.591562e-05, 7.860028e-05, 8.425368e-05, 9.151817e-05, 0.0001011913, 
    0.0001098135, 0.0001124116, 0.0001136011, 0.0001133161, 0.0001166245, 
    0.0001190862, 0.0001282328, 0.0001387681, 0.0001370877,
  0.0002057848, 0.0002059843, 0.0002080945, 0.0002118992, 0.0002306777, 
    0.0002435854, 0.0002603804, 0.0002474296, 0.0002581868, 0.0002335387, 
    0.0001802699, 0.0001492478, 0.0001305989, 0.0001121602, 0.0001007589, 
    9.893277e-05, 0.0001022899, 0.0001092407, 0.0001240063, 0.0001410949, 
    0.0001644498, 0.0001835247, 0.0001837143, 0.0001926131, 0.0001808594, 
    0.0001784017, 0.0001826465, 0.0001967008, 0.0002089139,
  0.0001191184, 0.0001389477, 0.0001520565, 0.0001483903, 0.0001462295, 
    0.0001409036, 0.0001490231, 0.0001606653, 0.0001787936, 0.000219674, 
    0.0002418808, 0.0002655193, 0.0002802582, 0.0002807731, 0.0002681838, 
    0.000262131, 0.0002215537, 0.0001943264, 0.0001641799, 0.0001475189, 
    0.0001261882, 0.0001131351, 0.000105293, 0.000112018, 0.0001236712, 
    0.000127708, 0.0001217182, 0.0001161934, 0.000115223,
  0.0001434052, 0.0001505985, 0.0001364014, 0.0001408724, 0.000148253, 
    0.0001414379, 0.0001436613, 0.0001525861, 0.0001549294, 0.000174464, 
    0.0001933646, 0.0001759472, 0.0001540961, 0.0001535316, 0.0001256537, 
    0.0001125303, 0.000101605, 9.872446e-05, 9.86037e-05, 9.698929e-05, 
    9.803126e-05, 0.0001020709, 0.0001023885, 0.0001065753, 0.0001087021, 
    0.0001142019, 0.0001216293, 0.0001328656, 0.0001400669,
  9.420435e-05, 9.125416e-05, 8.810619e-05, 8.527934e-05, 8.018594e-05, 
    7.869612e-05, 7.890844e-05, 9.317745e-05, 8.182873e-05, 0.0001036393, 
    0.0001215326, 0.0001158832, 0.000110741, 9.103363e-05, 8.012921e-05, 
    6.999969e-05, 6.706401e-05, 6.940648e-05, 7.00212e-05, 7.246408e-05, 
    7.779187e-05, 8.224558e-05, 8.343358e-05, 8.325782e-05, 8.479952e-05, 
    8.294461e-05, 8.652134e-05, 9.107365e-05, 9.454824e-05,
  2.72576e-05, 2.985417e-05, 3.192442e-05, 2.945079e-05, 2.530819e-05, 
    2.547828e-05, 2.136183e-05, 1.695792e-05, 1.469161e-05, 1.423639e-05, 
    1.68636e-05, 2.132316e-05, 3.849898e-05, 3.151772e-05, 2.696296e-05, 
    2.319139e-05, 1.995149e-05, 1.920738e-05, 1.752859e-05, 1.768787e-05, 
    1.675081e-05, 1.677076e-05, 1.802882e-05, 1.936664e-05, 2.042169e-05, 
    2.200773e-05, 2.268472e-05, 2.406466e-05, 2.561456e-05,
  6.18539e-06, 5.658614e-06, 5.24734e-06, 4.732855e-06, 4.495386e-06, 
    4.401393e-06, 3.280321e-06, 2.725634e-06, 2.291378e-06, 2.016665e-06, 
    2.063438e-06, 2.813936e-06, 5.212808e-06, 7.820426e-06, 8.608227e-06, 
    6.34187e-06, 5.582473e-06, 4.70027e-06, 3.727363e-06, 3.313296e-06, 
    2.356021e-06, 2.063229e-06, 2.07063e-06, 2.725134e-06, 3.140526e-06, 
    3.428101e-06, 3.71792e-06, 4.303351e-06, 5.5969e-06,
  1.138156e-06, 1.02528e-06, 8.755727e-07, 7.753117e-07, 6.774395e-07, 
    6.214205e-07, 6.264905e-07, 6.093347e-07, 4.64619e-07, 4.189289e-07, 
    5.754606e-07, 6.811329e-07, 8.583601e-07, 1.551445e-06, 1.425467e-06, 
    1.397659e-06, 1.290188e-06, 1.120241e-06, 7.877436e-07, 7.84618e-07, 
    7.04606e-07, 5.8249e-07, 6.093504e-07, 6.109928e-07, 6.352763e-07, 
    7.797868e-07, 8.256354e-07, 9.090377e-07, 9.662286e-07,
  4.085688e-07, 3.913011e-07, 4.166026e-07, 4.168905e-07, 3.29271e-07, 
    2.168689e-07, 1.48077e-07, 1.081566e-07, 1.028948e-07, 9.47031e-08, 
    8.908793e-08, 2.179523e-07, 2.659181e-07, 4.214036e-07, 4.519589e-07, 
    3.970697e-07, 5.38686e-07, 5.456628e-07, 5.129271e-07, 4.039567e-07, 
    3.876813e-07, 3.811832e-07, 2.965087e-07, 2.884667e-07, 3.090572e-07, 
    3.478422e-07, 3.966987e-07, 4.791472e-07, 4.180409e-07,
  1.957074e-07, 1.175589e-07, 1.024511e-07, 8.473086e-08, 9.545359e-08, 
    1.124075e-07, 1.291587e-07, 9.077928e-08, 6.449892e-08, 5.338212e-08, 
    4.590505e-08, 6.938848e-08, 1.113529e-07, 2.320822e-07, 1.820578e-07, 
    1.742675e-07, 1.90223e-07, 2.93598e-07, 4.254548e-07, 2.659576e-07, 
    2.097189e-07, 1.414613e-07, 9.164113e-08, 8.919126e-08, 1.299695e-07, 
    1.579685e-07, 2.318169e-07, 2.469329e-07, 2.351856e-07,
  7.815628e-08, 8.432929e-08, 8.507227e-08, 8.280055e-08, 8.713593e-08, 
    8.452496e-08, 8.453903e-08, 9.669758e-08, 8.618158e-08, 5.366616e-08, 
    2.962403e-08, 3.220097e-08, 4.600439e-08, 6.540478e-08, 1.054941e-07, 
    1.394873e-07, 1.323664e-07, 9.658617e-08, 7.155298e-08, 4.526055e-08, 
    2.736258e-08, 1.980423e-08, 2.173979e-08, 3.133263e-08, 3.065979e-08, 
    2.892981e-08, 3.845492e-08, 6.860014e-08, 7.61077e-08,
  8.500012e-09, 8.500012e-09, 8.500012e-09, 8.500012e-09, 8.500012e-09, 
    8.500012e-09, 8.500012e-09, 8.440455e-09, 8.440455e-09, 8.440455e-09, 
    8.440455e-09, 8.440455e-09, 8.440455e-09, 8.440455e-09, 9.083859e-09, 
    9.083859e-09, 9.083859e-09, 9.083859e-09, 9.083859e-09, 9.083859e-09, 
    9.083859e-09, 8.977735e-09, 8.977735e-09, 8.977735e-09, 8.977735e-09, 
    8.977735e-09, 8.977735e-09, 8.977735e-09, 8.500012e-09,
  1.236298e-08, 1.171917e-08, 1.241853e-08, 1.433933e-08, 1.603305e-08, 
    1.643527e-08, 1.543526e-08, 1.403959e-08, 1.288394e-08, 1.202964e-08, 
    1.135679e-08, 1.084944e-08, 1.101333e-08, 1.263885e-08, 1.443665e-08, 
    1.734687e-08, 1.902432e-08, 1.961155e-08, 1.866117e-08, 1.661804e-08, 
    1.662973e-08, 1.729017e-08, 1.850185e-08, 2.048175e-08, 1.917484e-08, 
    1.859565e-08, 1.672803e-08, 1.481642e-08, 1.295353e-08,
  3.155963e-08, 2.883595e-08, 2.884239e-08, 3.289884e-08, 3.992524e-08, 
    4.020269e-08, 3.329819e-08, 2.760956e-08, 2.584248e-08, 2.734689e-08, 
    2.760016e-08, 2.881462e-08, 3.761274e-08, 5.745026e-08, 8.010211e-08, 
    1.07923e-07, 1.159412e-07, 1.17409e-07, 1.147814e-07, 1.010734e-07, 
    8.760983e-08, 8.242331e-08, 7.939079e-08, 8.242187e-08, 9.293734e-08, 
    9.668801e-08, 8.04101e-08, 6.303283e-08, 3.966491e-08,
  2.201837e-07, 1.759451e-07, 1.812035e-07, 1.987459e-07, 2.137185e-07, 
    2.22337e-07, 2.242188e-07, 2.104739e-07, 2.424155e-07, 2.502892e-07, 
    2.419084e-07, 2.970938e-07, 4.809309e-07, 6.980455e-07, 9.25227e-07, 
    9.258999e-07, 7.663081e-07, 6.147403e-07, 5.519369e-07, 4.40124e-07, 
    3.77054e-07, 3.615652e-07, 4.030404e-07, 4.786916e-07, 5.429538e-07, 
    5.142225e-07, 4.277132e-07, 3.563468e-07, 2.814569e-07,
  1.274136e-06, 1.221075e-06, 1.494805e-06, 1.700241e-06, 2.178478e-06, 
    2.653446e-06, 2.641636e-06, 1.953312e-06, 1.369136e-06, 1.260095e-06, 
    1.325263e-06, 2.60366e-06, 3.005097e-06, 3.929393e-06, 3.986249e-06, 
    4.013602e-06, 2.974564e-06, 2.134617e-06, 1.397156e-06, 1.14327e-06, 
    1.085618e-06, 1.196936e-06, 1.35407e-06, 1.584245e-06, 2.048916e-06, 
    2.060256e-06, 1.865294e-06, 1.466518e-06, 1.212221e-06,
  1.128346e-05, 1.165001e-05, 1.520882e-05, 1.276038e-05, 9.939038e-06, 
    1.380944e-05, 1.108015e-05, 8.670796e-06, 9.495764e-06, 1.757962e-05, 
    1.974063e-05, 1.730651e-05, 1.991729e-05, 1.742438e-05, 1.486819e-05, 
    1.161721e-05, 7.672493e-06, 5.810083e-06, 5.430558e-06, 6.266617e-06, 
    5.123447e-06, 7.550868e-06, 9.572782e-06, 8.661682e-06, 1.066238e-05, 
    9.701468e-06, 8.116285e-06, 7.84964e-06, 1.02219e-05,
  0.0001140648, 0.0001156262, 0.0001145604, 0.0001234098, 0.0001227272, 
    0.0001217968, 0.000127298, 0.0001302915, 0.0001415124, 0.0001337772, 
    0.000109263, 8.191257e-05, 6.034641e-05, 4.698296e-05, 3.698276e-05, 
    3.368637e-05, 3.710045e-05, 5.270571e-05, 6.457489e-05, 7.125914e-05, 
    7.360706e-05, 7.596773e-05, 7.905557e-05, 8.737046e-05, 8.426647e-05, 
    8.376534e-05, 8.822882e-05, 9.932734e-05, 0.000109029,
  0.0006288398, 0.0006192607, 0.0006302245, 0.0006569066, 0.0006765724, 
    0.0006846797, 0.0006395376, 0.0006395178, 0.0005620344, 0.0004489166, 
    0.0003528303, 0.0002699832, 0.0002345819, 0.0002223523, 0.0002382709, 
    0.0002638332, 0.0003004182, 0.000327182, 0.0003634343, 0.0004095751, 
    0.0004417082, 0.0004744144, 0.0004873026, 0.000509778, 0.0005113721, 
    0.0005078585, 0.0005203135, 0.000556869, 0.0006094888,
  0.0009455283, 0.0009264402, 0.0009682499, 0.001054079, 0.001164255, 
    0.001272677, 0.001236246, 0.001295258, 0.001313969, 0.001147571, 
    0.0008925815, 0.0007321337, 0.000586113, 0.0004938514, 0.0004448412, 
    0.0004020105, 0.0004041463, 0.0004251283, 0.0004772846, 0.0005709875, 
    0.0007167701, 0.0008399065, 0.000872378, 0.0008069474, 0.00078023, 
    0.0008058342, 0.0008385524, 0.0008699569, 0.0009631916,
  0.0005890243, 0.0006835902, 0.0007138448, 0.0006613149, 0.0006254977, 
    0.0006712044, 0.0006914591, 0.0007960685, 0.001022759, 0.001129723, 
    0.001377337, 0.001550136, 0.001536826, 0.00139029, 0.001125413, 
    0.0008953993, 0.0006763001, 0.0005508327, 0.0004700208, 0.00042326, 
    0.0003745251, 0.0003889606, 0.0004751419, 0.0005478397, 0.0005667001, 
    0.0005360064, 0.0005089222, 0.0004916, 0.0005148027,
  0.0006670664, 0.0007251771, 0.000721001, 0.0007149652, 0.0007099576, 
    0.0006967997, 0.0007856204, 0.0007566086, 0.0008351767, 0.0009827767, 
    0.0009858049, 0.0008367938, 0.0007300259, 0.0005834269, 0.0005118484, 
    0.0004889813, 0.0004640079, 0.0004408936, 0.0004047358, 0.0003926789, 
    0.0004130707, 0.0004245184, 0.0004282526, 0.0004133105, 0.0004459244, 
    0.0004876902, 0.0005338354, 0.0006003806, 0.0006641141,
  0.0005189366, 0.000534185, 0.0005234469, 0.0004820327, 0.0004488447, 
    0.0004307752, 0.0004716152, 0.000434451, 0.0003591972, 0.0004596383, 
    0.0005502357, 0.0006104594, 0.0005546423, 0.0004156776, 0.0003655677, 
    0.0003251823, 0.0002940703, 0.0003042148, 0.0003078704, 0.0003137352, 
    0.0003228395, 0.0003452731, 0.0003601127, 0.000388033, 0.0004139367, 
    0.0004275769, 0.0004400168, 0.0004719325, 0.0005154251,
  0.0001678822, 0.0001807438, 0.0001895189, 0.0001789954, 0.0001710267, 
    0.0001561434, 0.0001458338, 0.0001146502, 9.482702e-05, 8.523979e-05, 
    7.651682e-05, 9.697704e-05, 0.0001544395, 0.0001344494, 0.0001103875, 
    0.0001040979, 8.492553e-05, 7.982561e-05, 7.986029e-05, 7.535171e-05, 
    7.675556e-05, 8.046812e-05, 8.300058e-05, 8.94033e-05, 9.863149e-05, 
    0.0001064047, 0.0001195065, 0.0001323484, 0.000152529,
  3.413183e-05, 3.196423e-05, 3.245256e-05, 2.847878e-05, 2.572104e-05, 
    2.370775e-05, 2.621598e-05, 2.131101e-05, 1.353258e-05, 1.202004e-05, 
    1.222709e-05, 1.434728e-05, 1.967911e-05, 3.059734e-05, 3.283004e-05, 
    2.716915e-05, 2.524441e-05, 2.319625e-05, 2.00772e-05, 1.648665e-05, 
    1.323836e-05, 9.768886e-06, 8.932315e-06, 1.239017e-05, 1.315947e-05, 
    1.50741e-05, 1.738656e-05, 2.138934e-05, 2.911017e-05,
  5.131739e-06, 5.712016e-06, 4.980288e-06, 3.777858e-06, 3.693296e-06, 
    3.101304e-06, 3.11751e-06, 2.6353e-06, 2.309818e-06, 2.351944e-06, 
    2.992674e-06, 3.713645e-06, 4.050794e-06, 6.228804e-06, 6.784693e-06, 
    6.507369e-06, 5.763118e-06, 5.256361e-06, 5.428223e-06, 5.054721e-06, 
    4.30129e-06, 2.77787e-06, 2.224795e-06, 2.100511e-06, 2.317941e-06, 
    2.959127e-06, 3.310366e-06, 3.782679e-06, 4.45506e-06,
  1.739589e-06, 1.64327e-06, 1.592727e-06, 1.636327e-06, 1.477671e-06, 
    1.159131e-06, 8.635899e-07, 5.291603e-07, 5.333981e-07, 5.327021e-07, 
    4.319053e-07, 9.320585e-07, 1.204665e-06, 1.617487e-06, 1.631191e-06, 
    1.513056e-06, 1.662447e-06, 1.841789e-06, 1.963003e-06, 1.731158e-06, 
    1.761426e-06, 1.534047e-06, 1.127852e-06, 1.162914e-06, 1.221125e-06, 
    1.262594e-06, 1.352851e-06, 1.573784e-06, 2.024753e-06,
  1.066923e-06, 6.725595e-07, 4.273089e-07, 3.846937e-07, 3.998158e-07, 
    4.389257e-07, 5.116722e-07, 3.477953e-07, 2.538849e-07, 2.375429e-07, 
    1.786432e-07, 2.813837e-07, 4.183061e-07, 7.637622e-07, 6.840417e-07, 
    5.13571e-07, 4.918311e-07, 7.134407e-07, 9.089155e-07, 7.783798e-07, 
    5.672262e-07, 4.411436e-07, 3.023537e-07, 6.376177e-07, 7.249242e-07, 
    8.301332e-07, 1.04875e-06, 1.197412e-06, 1.216981e-06,
  3.870574e-07, 3.617488e-07, 3.560413e-07, 3.633225e-07, 3.832072e-07, 
    3.888843e-07, 3.412711e-07, 3.131097e-07, 2.974407e-07, 2.254813e-07, 
    1.596676e-07, 1.619802e-07, 2.219746e-07, 2.901252e-07, 3.784577e-07, 
    4.444063e-07, 4.41336e-07, 3.339986e-07, 2.374499e-07, 1.542176e-07, 
    1.030354e-07, 8.670732e-08, 1.059536e-07, 1.308743e-07, 1.362385e-07, 
    1.443864e-07, 2.30928e-07, 3.923549e-07, 4.15143e-07,
  5.857941e-08, 5.857941e-08, 5.857941e-08, 5.857941e-08, 5.857941e-08, 
    5.857941e-08, 5.857941e-08, 5.872547e-08, 5.872547e-08, 5.872547e-08, 
    5.872547e-08, 5.872547e-08, 5.872547e-08, 5.872547e-08, 6.120026e-08, 
    6.120026e-08, 6.120026e-08, 6.120026e-08, 6.120026e-08, 6.120026e-08, 
    6.120026e-08, 6.143682e-08, 6.143682e-08, 6.143682e-08, 6.143682e-08, 
    6.143682e-08, 6.143682e-08, 6.143682e-08, 5.857941e-08,
  6.779644e-08, 6.766712e-08, 7.067862e-08, 7.711986e-08, 8.353386e-08, 
    8.417005e-08, 7.686649e-08, 6.820419e-08, 6.060448e-08, 5.096163e-08, 
    4.863338e-08, 4.986508e-08, 5.148968e-08, 5.410787e-08, 5.979548e-08, 
    6.923264e-08, 7.9656e-08, 8.256725e-08, 8.68848e-08, 8.749307e-08, 
    8.67896e-08, 8.965506e-08, 9.363931e-08, 1.002393e-07, 9.586101e-08, 
    9.312033e-08, 8.589602e-08, 7.732692e-08, 6.88033e-08,
  1.866951e-07, 1.46221e-07, 1.376738e-07, 1.562483e-07, 1.903312e-07, 
    1.993048e-07, 1.55542e-07, 1.225023e-07, 1.157987e-07, 1.243348e-07, 
    1.174284e-07, 1.301727e-07, 1.581351e-07, 2.436155e-07, 3.801492e-07, 
    4.18528e-07, 4.763164e-07, 4.922978e-07, 4.907824e-07, 5.007056e-07, 
    4.852423e-07, 4.509154e-07, 4.627276e-07, 4.538898e-07, 4.582693e-07, 
    4.799586e-07, 4.039756e-07, 3.034341e-07, 2.175543e-07,
  1.117271e-06, 9.40833e-07, 8.736912e-07, 9.392499e-07, 9.906147e-07, 
    1.085283e-06, 1.026935e-06, 9.303521e-07, 1.044782e-06, 1.078783e-06, 
    1.051647e-06, 1.336364e-06, 1.757746e-06, 2.565642e-06, 3.563283e-06, 
    3.814168e-06, 3.32399e-06, 2.818184e-06, 2.441574e-06, 2.018571e-06, 
    1.651137e-06, 1.666123e-06, 1.852941e-06, 2.239265e-06, 2.486143e-06, 
    2.072865e-06, 1.772052e-06, 1.606321e-06, 1.42742e-06,
  5.801122e-06, 5.280924e-06, 6.572511e-06, 8.148586e-06, 9.412462e-06, 
    1.098747e-05, 1.117005e-05, 8.305259e-06, 5.962425e-06, 5.279118e-06, 
    5.772062e-06, 1.043831e-05, 1.212018e-05, 1.63181e-05, 1.98573e-05, 
    2.328135e-05, 1.825238e-05, 1.204553e-05, 8.219113e-06, 5.844187e-06, 
    5.361395e-06, 5.525671e-06, 6.213229e-06, 7.375524e-06, 8.97201e-06, 
    9.342603e-06, 8.44964e-06, 7.272554e-06, 5.957445e-06,
  4.392455e-05, 4.395329e-05, 5.4185e-05, 7.232597e-05, 5.187738e-05, 
    5.614496e-05, 6.251838e-05, 4.292359e-05, 4.144715e-05, 7.38871e-05, 
    9.851985e-05, 9.69603e-05, 9.790649e-05, 9.730054e-05, 9.079609e-05, 
    6.857231e-05, 4.585308e-05, 3.378205e-05, 2.759181e-05, 2.904709e-05, 
    2.805964e-05, 3.36027e-05, 4.252272e-05, 4.412905e-05, 5.686101e-05, 
    5.52032e-05, 4.512387e-05, 3.462937e-05, 3.974442e-05,
  0.000439007, 0.0004444767, 0.0004127123, 0.0004703079, 0.0005814514, 
    0.0006147179, 0.000719085, 0.0007713039, 0.0008235874, 0.0009359402, 
    0.0008148037, 0.000659853, 0.0004404031, 0.0003072294, 0.0002392245, 
    0.0001609058, 0.0001497949, 0.0001705063, 0.0002183189, 0.0002568085, 
    0.0003025305, 0.0003267181, 0.0003323283, 0.0003748785, 0.000400538, 
    0.0003724276, 0.0003561949, 0.0003660242, 0.0004174991,
  0.002452331, 0.002499606, 0.00273045, 0.002731599, 0.002781128, 
    0.003046817, 0.003335435, 0.003340026, 0.003336324, 0.002930594, 
    0.002182928, 0.001553683, 0.001133821, 0.0009100092, 0.0008014613, 
    0.0008168529, 0.0009270109, 0.00107418, 0.001237636, 0.001442886, 
    0.001681119, 0.001795069, 0.001804525, 0.001846652, 0.00190185, 
    0.001947677, 0.002116716, 0.002221513, 0.002288076,
  0.00466784, 0.004570714, 0.004746271, 0.005017328, 0.005320365, 
    0.005776304, 0.006330625, 0.006312879, 0.006639414, 0.006681722, 
    0.00487133, 0.003358783, 0.00242402, 0.00214458, 0.001821822, 
    0.001541981, 0.00138437, 0.001404126, 0.001707423, 0.002249992, 
    0.003093368, 0.003658907, 0.003666024, 0.00369485, 0.003467216, 
    0.003380664, 0.003565121, 0.004032261, 0.004295592,
  0.003394886, 0.003391148, 0.003353902, 0.003134303, 0.002893142, 
    0.003126987, 0.003378051, 0.004528722, 0.005556052, 0.006912713, 
    0.008433945, 0.007533637, 0.006223011, 0.004566752, 0.003200778, 
    0.002486055, 0.002156715, 0.001910307, 0.001730197, 0.001669716, 
    0.001873171, 0.002201809, 0.002614499, 0.00308457, 0.002652672, 
    0.002481793, 0.002502718, 0.002370899, 0.002996823,
  0.00310149, 0.003194296, 0.003515978, 0.003756515, 0.003915469, 0.00396176, 
    0.004368243, 0.004168548, 0.004886118, 0.00552304, 0.004669731, 
    0.003366917, 0.002911425, 0.0021411, 0.001883805, 0.001925191, 
    0.00176348, 0.001740745, 0.00176481, 0.001797367, 0.00195493, 
    0.002040947, 0.002278784, 0.001997025, 0.001966407, 0.002113574, 
    0.002221136, 0.002844458, 0.00290269,
  0.002432782, 0.002718534, 0.003092507, 0.003361948, 0.003341212, 
    0.003093101, 0.003013208, 0.002628157, 0.002253873, 0.002248284, 
    0.002920536, 0.002818269, 0.00236185, 0.001756496, 0.001488567, 
    0.001327828, 0.001156608, 0.0011584, 0.001156165, 0.001249501, 
    0.00132764, 0.001449604, 0.001551756, 0.001583465, 0.00163951, 
    0.001681962, 0.001828582, 0.002007289, 0.002192507,
  0.0008363786, 0.000980138, 0.001037078, 0.001105294, 0.001117129, 
    0.001140614, 0.001033475, 0.0008148407, 0.0006949771, 0.000567825, 
    0.0004579335, 0.0004550882, 0.0006671855, 0.0005721031, 0.0004172615, 
    0.0003782873, 0.00033838, 0.0002891902, 0.0002791312, 0.000262894, 
    0.0002514981, 0.0002841002, 0.0003579944, 0.0003849645, 0.0004105349, 
    0.0004591878, 0.0004835864, 0.0005604137, 0.0007114828,
  0.0001847424, 0.0001910129, 0.0002083477, 0.0001946129, 0.0001694548, 
    0.0001477352, 0.0001929267, 0.0001849485, 0.0001022909, 6.632737e-05, 
    7.060682e-05, 8.665652e-05, 8.854567e-05, 0.0001128651, 0.0001197306, 
    9.083275e-05, 8.447813e-05, 9.499094e-05, 8.603474e-05, 7.382369e-05, 
    6.85272e-05, 4.800523e-05, 4.110828e-05, 5.122586e-05, 4.848807e-05, 
    5.429229e-05, 6.288201e-05, 8.422103e-05, 0.0001371253,
  2.148748e-05, 3.358223e-05, 2.889081e-05, 2.058798e-05, 2.099449e-05, 
    1.76453e-05, 1.806538e-05, 1.506687e-05, 1.400604e-05, 1.253287e-05, 
    1.652088e-05, 1.945869e-05, 2.23358e-05, 2.511752e-05, 3.056286e-05, 
    2.701024e-05, 2.365295e-05, 2.549567e-05, 2.516161e-05, 2.816323e-05, 
    2.085528e-05, 1.225688e-05, 8.998196e-06, 7.678796e-06, 9.118648e-06, 
    1.181778e-05, 1.30208e-05, 1.367386e-05, 1.692566e-05,
  5.803916e-06, 6.52678e-06, 7.410573e-06, 6.221434e-06, 7.455463e-06, 
    6.098544e-06, 5.330687e-06, 3.170255e-06, 2.88795e-06, 2.759368e-06, 
    2.62546e-06, 3.707936e-06, 5.580541e-06, 6.664179e-06, 6.953098e-06, 
    5.454423e-06, 5.42732e-06, 6.196356e-06, 7.409286e-06, 7.72461e-06, 
    6.557743e-06, 5.557994e-06, 4.444191e-06, 4.426036e-06, 4.322521e-06, 
    4.239459e-06, 5.520395e-06, 6.120707e-06, 6.925858e-06,
  3.666933e-06, 2.791546e-06, 2.188596e-06, 1.901741e-06, 1.880366e-06, 
    2.174407e-06, 2.273616e-06, 1.590586e-06, 1.168126e-06, 1.111785e-06, 
    1.365777e-06, 1.021762e-06, 1.325433e-06, 2.21915e-06, 2.19581e-06, 
    1.598491e-06, 1.494796e-06, 1.762098e-06, 1.810398e-06, 2.007209e-06, 
    1.514838e-06, 1.350637e-06, 1.179189e-06, 2.416883e-06, 2.656243e-06, 
    2.890501e-06, 3.59528e-06, 3.898077e-06, 3.994714e-06,
  1.784873e-06, 1.418318e-06, 1.319073e-06, 1.345317e-06, 1.382932e-06, 
    1.398397e-06, 1.337449e-06, 1.141195e-06, 9.794659e-07, 8.071424e-07, 
    6.916862e-07, 8.535012e-07, 9.375082e-07, 8.647522e-07, 8.86193e-07, 
    9.964851e-07, 1.023824e-06, 8.761277e-07, 6.926421e-07, 5.080891e-07, 
    3.43804e-07, 3.41751e-07, 4.111566e-07, 5.052038e-07, 6.398852e-07, 
    8.572708e-07, 1.336056e-06, 1.850524e-06, 1.934567e-06,
  3.12504e-07, 3.12504e-07, 3.12504e-07, 3.12504e-07, 3.12504e-07, 
    3.12504e-07, 3.12504e-07, 3.117875e-07, 3.117875e-07, 3.117875e-07, 
    3.117875e-07, 3.117875e-07, 3.117875e-07, 3.117875e-07, 3.148462e-07, 
    3.148462e-07, 3.148462e-07, 3.148462e-07, 3.148462e-07, 3.148462e-07, 
    3.148462e-07, 3.286316e-07, 3.286316e-07, 3.286316e-07, 3.286316e-07, 
    3.286316e-07, 3.286316e-07, 3.286316e-07, 3.12504e-07,
  3.301741e-07, 3.471152e-07, 3.710489e-07, 4.3967e-07, 5.370691e-07, 
    5.272037e-07, 4.72165e-07, 4.236023e-07, 3.697624e-07, 2.667354e-07, 
    2.442824e-07, 2.321262e-07, 2.312947e-07, 2.604161e-07, 2.858878e-07, 
    3.181821e-07, 3.696588e-07, 4.097227e-07, 4.343699e-07, 4.45384e-07, 
    4.665e-07, 4.752284e-07, 4.842073e-07, 5.059712e-07, 4.67282e-07, 
    4.412847e-07, 4.106881e-07, 3.731714e-07, 3.334029e-07,
  1.303898e-06, 1.065519e-06, 8.24507e-07, 9.026937e-07, 1.040319e-06, 
    1.089242e-06, 8.44001e-07, 6.696577e-07, 6.182797e-07, 5.814449e-07, 
    5.612119e-07, 6.767475e-07, 7.585218e-07, 9.258544e-07, 1.728375e-06, 
    1.834944e-06, 1.805234e-06, 2.050725e-06, 2.17011e-06, 2.217094e-06, 
    2.193426e-06, 2.13515e-06, 2.082573e-06, 2.024202e-06, 2.071621e-06, 
    2.168406e-06, 1.923315e-06, 1.528992e-06, 1.303438e-06,
  5.543566e-06, 4.575447e-06, 4.236394e-06, 4.764416e-06, 4.549068e-06, 
    4.873936e-06, 5.059014e-06, 4.524162e-06, 4.399311e-06, 3.995645e-06, 
    4.075895e-06, 5.095711e-06, 6.518176e-06, 1.033531e-05, 1.620688e-05, 
    1.911728e-05, 1.423331e-05, 1.027003e-05, 9.174642e-06, 8.02102e-06, 
    7.081152e-06, 6.74813e-06, 7.866717e-06, 9.336618e-06, 1.102577e-05, 
    9.643661e-06, 8.002893e-06, 6.526805e-06, 6.942843e-06,
  2.537253e-05, 2.400094e-05, 2.794489e-05, 3.807666e-05, 4.404825e-05, 
    4.68078e-05, 4.120832e-05, 3.808734e-05, 2.768073e-05, 2.209124e-05, 
    2.461502e-05, 4.261809e-05, 5.473217e-05, 7.172041e-05, 0.0001062776, 
    0.0001353221, 9.570314e-05, 6.687546e-05, 4.302206e-05, 3.013137e-05, 
    2.678886e-05, 2.652051e-05, 3.036993e-05, 3.418794e-05, 3.876079e-05, 
    4.049233e-05, 3.436485e-05, 3.211341e-05, 2.802394e-05,
  0.0001659673, 0.0001795738, 0.0002141969, 0.0002813233, 0.0002606554, 
    0.0002348092, 0.0003518256, 0.0002431742, 0.0001838235, 0.000239902, 
    0.0004383088, 0.0004257543, 0.0004305731, 0.0003955752, 0.000443729, 
    0.0004076424, 0.0003528681, 0.0002098203, 0.000138168, 0.0001294602, 
    0.0001440379, 0.0001733915, 0.0001936655, 0.0002299615, 0.0002818954, 
    0.0002693761, 0.0002321504, 0.0001724067, 0.0001669487,
  0.001987076, 0.001884868, 0.001569255, 0.001437799, 0.001917313, 
    0.002332663, 0.003358415, 0.004205957, 0.004716828, 0.005044765, 
    0.004442196, 0.004583756, 0.002875473, 0.001800844, 0.001562065, 
    0.001064083, 0.0007096175, 0.0006951219, 0.0008158199, 0.0009751123, 
    0.001196965, 0.00153609, 0.001700739, 0.002083227, 0.002186564, 
    0.001586781, 0.001607804, 0.001549825, 0.001576706,
  0.009513591, 0.009404593, 0.009623173, 0.01082181, 0.01059308, 0.01106281, 
    0.01342559, 0.01715366, 0.01782249, 0.01907616, 0.01529714, 0.01272571, 
    0.008133963, 0.005503328, 0.003829656, 0.002726599, 0.002666443, 
    0.002883146, 0.003479064, 0.004560563, 0.005990956, 0.007653317, 
    0.008168336, 0.008008608, 0.007442123, 0.006475079, 0.007005989, 
    0.008251509, 0.009343663,
  0.01794833, 0.01860093, 0.01822674, 0.01976869, 0.02177808, 0.02526226, 
    0.02869011, 0.03560802, 0.03679873, 0.03892151, 0.02985905, 0.0204911, 
    0.01542508, 0.01269582, 0.01171329, 0.007654424, 0.005167237, 
    0.004340081, 0.005029705, 0.007665359, 0.01343584, 0.01876449, 0.020145, 
    0.01811868, 0.01494002, 0.01335677, 0.01386496, 0.01548766, 0.01905096,
  0.02034116, 0.01778628, 0.01694014, 0.01564602, 0.01548589, 0.01645909, 
    0.02050203, 0.02514697, 0.03079902, 0.03725656, 0.03972039, 0.03148018, 
    0.02503829, 0.02053183, 0.01546019, 0.01236813, 0.009986592, 0.008277071, 
    0.007280075, 0.008857005, 0.01262072, 0.01472665, 0.01720642, 0.01604231, 
    0.01435864, 0.01411557, 0.01465358, 0.01392985, 0.01909509,
  0.01657215, 0.01549724, 0.01761363, 0.0175547, 0.02136891, 0.02171575, 
    0.02336084, 0.02783269, 0.0278329, 0.03019086, 0.02329851, 0.01584607, 
    0.01445248, 0.01314752, 0.01239544, 0.009639712, 0.008270093, 
    0.007493459, 0.006451219, 0.007127885, 0.009170191, 0.009848359, 
    0.01125803, 0.009602661, 0.01002949, 0.01082598, 0.01139546, 0.01412541, 
    0.0157625,
  0.009577685, 0.01262951, 0.01525983, 0.01614964, 0.01798273, 0.01898467, 
    0.01796107, 0.01727191, 0.01413191, 0.01316143, 0.01469814, 0.01420465, 
    0.01217308, 0.009649262, 0.007495977, 0.006066739, 0.004743438, 
    0.004290455, 0.003589112, 0.003416857, 0.003942873, 0.005028651, 
    0.00605003, 0.006300424, 0.006607735, 0.006265962, 0.006289771, 
    0.007275558, 0.008481087,
  0.003286852, 0.004547493, 0.005427477, 0.005578173, 0.00618141, 
    0.006856555, 0.007164434, 0.005606224, 0.005170626, 0.004961129, 
    0.00297763, 0.002297248, 0.002841253, 0.002649435, 0.001783159, 
    0.001334623, 0.001212519, 0.001123413, 0.0009831856, 0.0009897425, 
    0.000990134, 0.0009553506, 0.001115887, 0.001399249, 0.001537521, 
    0.001613095, 0.001718354, 0.001917785, 0.002573793,
  0.0009037484, 0.001016216, 0.001194034, 0.001267043, 0.001145038, 
    0.0008609003, 0.0010218, 0.00112788, 0.0006945697, 0.0003717715, 
    0.0003731806, 0.0004735186, 0.000463519, 0.0004861248, 0.0004802987, 
    0.0003128643, 0.0002659672, 0.0003085755, 0.0003155344, 0.0003064451, 
    0.0003269405, 0.0003051358, 0.0002033779, 0.0001656256, 0.0002459577, 
    0.0001562714, 0.0001711513, 0.0002453393, 0.0005153844,
  7.697652e-05, 0.0001822903, 0.0001712169, 0.0001204573, 0.0001193867, 
    8.713959e-05, 9.464985e-05, 0.0001068179, 8.206739e-05, 8.702652e-05, 
    0.0001031147, 0.0001210336, 0.00012909, 0.0001225352, 0.0001206358, 
    0.0001025435, 8.532017e-05, 9.221695e-05, 0.0001032107, 0.0001247152, 
    8.521394e-05, 5.520225e-05, 4.000334e-05, 3.284476e-05, 4.201171e-05, 
    4.660962e-05, 5.411548e-05, 5.622687e-05, 5.225012e-05,
  2.319655e-05, 2.629488e-05, 4.156347e-05, 3.247894e-05, 3.47473e-05, 
    3.165717e-05, 3.301501e-05, 2.497452e-05, 1.891257e-05, 1.565645e-05, 
    1.685326e-05, 1.874923e-05, 2.379239e-05, 2.641515e-05, 2.642844e-05, 
    2.134378e-05, 2.142868e-05, 2.054326e-05, 2.404175e-05, 2.70927e-05, 
    2.17645e-05, 1.750842e-05, 1.470276e-05, 1.298049e-05, 1.612585e-05, 
    1.742013e-05, 2.383168e-05, 2.974115e-05, 2.705658e-05,
  9.872597e-06, 8.821434e-06, 8.123715e-06, 1.19571e-05, 8.075297e-06, 
    8.90106e-06, 8.733345e-06, 8.312296e-06, 5.5774e-06, 5.109349e-06, 
    8.398847e-06, 4.955572e-06, 4.716204e-06, 6.6679e-06, 7.139614e-06, 
    5.8874e-06, 4.831075e-06, 5.347648e-06, 5.591447e-06, 6.194433e-06, 
    5.340728e-06, 4.444499e-06, 4.591127e-06, 6.520439e-06, 6.455281e-06, 
    8.844192e-06, 1.133738e-05, 1.157838e-05, 1.025785e-05,
  4.978866e-06, 4.754008e-06, 4.829935e-06, 4.847029e-06, 4.811418e-06, 
    4.536181e-06, 4.251076e-06, 3.928328e-06, 3.53869e-06, 3.546053e-06, 
    3.568276e-06, 3.666933e-06, 2.996293e-06, 2.169314e-06, 1.91354e-06, 
    2.048416e-06, 2.22511e-06, 2.100823e-06, 1.8529e-06, 1.616779e-06, 
    1.386592e-06, 1.281005e-06, 1.664948e-06, 2.326921e-06, 2.900738e-06, 
    3.583356e-06, 4.282806e-06, 4.92152e-06, 5.069943e-06,
  1.958516e-06, 1.958516e-06, 1.958516e-06, 1.958516e-06, 1.958516e-06, 
    1.958516e-06, 1.958516e-06, 1.791175e-06, 1.791175e-06, 1.791175e-06, 
    1.791175e-06, 1.791175e-06, 1.791175e-06, 1.791175e-06, 1.754707e-06, 
    1.754707e-06, 1.754707e-06, 1.754707e-06, 1.754707e-06, 1.754707e-06, 
    1.754707e-06, 1.869377e-06, 1.869377e-06, 1.869377e-06, 1.869377e-06, 
    1.869377e-06, 1.869377e-06, 1.869377e-06, 1.958516e-06,
  1.62583e-06, 1.74109e-06, 2.107263e-06, 2.776072e-06, 2.947424e-06, 
    2.672812e-06, 2.397529e-06, 2.234417e-06, 1.917814e-06, 1.359319e-06, 
    1.30568e-06, 1.315057e-06, 1.213928e-06, 1.356994e-06, 1.486241e-06, 
    1.609094e-06, 1.818237e-06, 1.988961e-06, 2.125308e-06, 2.199153e-06, 
    2.324894e-06, 2.371539e-06, 2.563574e-06, 2.497478e-06, 2.279886e-06, 
    2.254319e-06, 2.036999e-06, 1.852446e-06, 1.639284e-06,
  3.82715e-06, 3.878873e-06, 4.778783e-06, 4.599789e-06, 5.367535e-06, 
    5.410542e-06, 4.115498e-06, 3.289593e-06, 3.192868e-06, 2.912474e-06, 
    2.804429e-06, 3.170321e-06, 3.589636e-06, 4.080003e-06, 5.400698e-06, 
    8.108256e-06, 8.625481e-06, 8.710179e-06, 9.490793e-06, 8.407871e-06, 
    7.975328e-06, 8.247748e-06, 8.665341e-06, 8.642426e-06, 9.237239e-06, 
    9.251858e-06, 8.506517e-06, 7.15897e-06, 4.549748e-06,
  2.843354e-05, 2.282802e-05, 1.830093e-05, 1.982687e-05, 2.066549e-05, 
    2.178131e-05, 2.26284e-05, 2.008408e-05, 1.71892e-05, 1.564782e-05, 
    1.579546e-05, 1.984002e-05, 3.250565e-05, 4.687976e-05, 7.33815e-05, 
    7.417409e-05, 5.938791e-05, 4.111645e-05, 3.58293e-05, 3.137211e-05, 
    2.820048e-05, 2.990778e-05, 3.024231e-05, 3.640025e-05, 4.39223e-05, 
    4.101495e-05, 3.265215e-05, 2.675315e-05, 2.429201e-05,
  0.0001124084, 0.000103619, 0.000114601, 0.0001371517, 0.0001844882, 
    0.0001872342, 0.0001665341, 0.0001447395, 0.0001287631, 0.0001017276, 
    0.0001153662, 0.0001975956, 0.000323709, 0.0004026688, 0.0005509502, 
    0.0006454759, 0.0004648864, 0.0002901809, 0.0001692575, 0.0001155894, 
    0.0001062251, 0.0001203283, 0.0001314091, 0.0001452921, 0.0001653995, 
    0.0001638713, 0.0001432021, 0.0001323836, 0.0001314278,
  0.0006477858, 0.000724093, 0.0009831218, 0.001003014, 0.0009608711, 
    0.0009175014, 0.001220961, 0.001139161, 0.0008776459, 0.001194843, 
    0.002312799, 0.002449131, 0.002268364, 0.002015834, 0.002537636, 
    0.00245718, 0.002040204, 0.001191424, 0.0007680603, 0.0006049401, 
    0.0006854247, 0.0007690946, 0.0007092824, 0.0009128216, 0.001264328, 
    0.001081427, 0.0009324828, 0.0007675994, 0.0006729173,
  0.007584499, 0.008655318, 0.007786477, 0.006423475, 0.005520491, 
    0.009068802, 0.01705047, 0.02188403, 0.02901024, 0.03780846, 0.03732141, 
    0.03083732, 0.02188337, 0.01196604, 0.009761773, 0.007503362, 
    0.004436135, 0.002953695, 0.003318209, 0.003968379, 0.004892206, 
    0.005426038, 0.007472956, 0.009536668, 0.01045442, 0.007613653, 
    0.00629758, 0.005834961, 0.005709078,
  0.0367212, 0.03967365, 0.03591872, 0.0340642, 0.04111185, 0.05132816, 
    0.07303645, 0.1189869, 0.1408233, 0.1825889, 0.1814617, 0.1484395, 
    0.0904057, 0.05222952, 0.03402713, 0.02008131, 0.01126044, 0.008050933, 
    0.008631295, 0.01201586, 0.02111759, 0.02838861, 0.03764914, 0.04095976, 
    0.03688606, 0.02695139, 0.02236625, 0.02527422, 0.03272266,
  0.08848865, 0.07508942, 0.0657433, 0.06564432, 0.07909802, 0.1078921, 
    0.1396559, 0.1829016, 0.2113809, 0.2403494, 0.2562993, 0.2366008, 
    0.1594232, 0.1236608, 0.09190873, 0.06079875, 0.03933368, 0.02418393, 
    0.02245723, 0.02661989, 0.04071167, 0.06775946, 0.09924942, 0.1209719, 
    0.09670568, 0.05837413, 0.0451137, 0.05533312, 0.07631736,
  0.1055854, 0.09452714, 0.08473237, 0.07375075, 0.07935736, 0.08832012, 
    0.1076173, 0.1275276, 0.1544657, 0.1783177, 0.202122, 0.1940544, 
    0.1459739, 0.1234493, 0.1036072, 0.08387729, 0.06489346, 0.04801891, 
    0.04059161, 0.03884819, 0.05491634, 0.06833779, 0.08352109, 0.08762152, 
    0.07368241, 0.06916498, 0.06243597, 0.06284413, 0.07984255,
  0.07985778, 0.09279373, 0.1032552, 0.130616, 0.1341424, 0.133048, 
    0.1435034, 0.1521543, 0.1667381, 0.1787452, 0.1496339, 0.1209844, 
    0.1075537, 0.09319262, 0.07683852, 0.05744418, 0.04377423, 0.04155604, 
    0.0341391, 0.02728678, 0.03419838, 0.04316702, 0.0443358, 0.03865431, 
    0.03662515, 0.04017362, 0.04408037, 0.05090991, 0.06780466,
  0.04647778, 0.06806315, 0.09685263, 0.1252178, 0.1365876, 0.1388215, 
    0.1414614, 0.1596237, 0.1286879, 0.1016445, 0.08938098, 0.08543765, 
    0.06750993, 0.04778647, 0.03527029, 0.02730338, 0.02039137, 0.01757323, 
    0.01586931, 0.01348496, 0.01259408, 0.01505014, 0.01744062, 0.01854104, 
    0.01977458, 0.02116507, 0.02234646, 0.02559988, 0.03365621,
  0.01602475, 0.02457202, 0.03135889, 0.03871426, 0.04306677, 0.04251378, 
    0.05108759, 0.0543225, 0.05280622, 0.03924027, 0.02141719, 0.01385783, 
    0.01196454, 0.01213908, 0.007675717, 0.004901269, 0.004168263, 
    0.004462791, 0.003966677, 0.004404755, 0.004833205, 0.004322106, 
    0.003927785, 0.004358059, 0.004852857, 0.004811373, 0.004788956, 
    0.006925664, 0.01057826,
  0.003452856, 0.004387477, 0.005063917, 0.006080682, 0.005831243, 
    0.004147286, 0.00529718, 0.006133537, 0.004254591, 0.002652838, 
    0.002336521, 0.002509495, 0.002537669, 0.002106441, 0.001927359, 
    0.001169497, 0.0009252715, 0.000974403, 0.001083729, 0.001256226, 
    0.001516383, 0.001340594, 0.0009592054, 0.0006497533, 0.001137492, 
    0.0005774921, 0.0005058986, 0.0006016758, 0.001559107,
  0.0002393177, 0.0005281342, 0.0007603577, 0.0007130235, 0.0004559016, 
    0.0003748478, 0.0003933798, 0.000471423, 0.00047035, 0.0004572041, 
    0.0006049742, 0.000651225, 0.0006274943, 0.0006138408, 0.0004830318, 
    0.0004385473, 0.0002903893, 0.0002874661, 0.0003558621, 0.0003643431, 
    0.0003348206, 0.0002453472, 0.0001799766, 0.0001457779, 0.0001454237, 
    0.0001831493, 0.0002014856, 0.000202004, 0.0001691899,
  7.3406e-05, 8.547234e-05, 0.0001852205, 0.0001857559, 0.0001675913, 
    0.000143951, 0.0001470463, 0.0001844616, 0.0001063618, 9.882201e-05, 
    9.39652e-05, 0.0001038683, 0.0001031221, 0.0001077158, 0.0001036949, 
    7.912937e-05, 6.986621e-05, 6.759453e-05, 7.888361e-05, 8.478512e-05, 
    7.388525e-05, 5.452372e-05, 4.310601e-05, 4.203002e-05, 6.589148e-05, 
    6.551413e-05, 7.946837e-05, 0.000101982, 9.039854e-05,
  2.797629e-05, 2.52085e-05, 2.675618e-05, 4.867624e-05, 5.270451e-05, 
    4.81108e-05, 3.085753e-05, 3.436915e-05, 3.257811e-05, 3.075518e-05, 
    3.205539e-05, 2.466284e-05, 1.919722e-05, 2.269234e-05, 2.353203e-05, 
    2.059286e-05, 1.878513e-05, 1.981179e-05, 2.267682e-05, 2.319911e-05, 
    1.998042e-05, 1.573426e-05, 1.540083e-05, 1.725032e-05, 1.899041e-05, 
    2.844725e-05, 3.40937e-05, 3.520018e-05, 3.340296e-05,
  1.554238e-05, 1.75415e-05, 2.052131e-05, 1.98281e-05, 2.075282e-05, 
    1.936382e-05, 1.623973e-05, 1.592615e-05, 1.565292e-05, 1.669335e-05, 
    1.735998e-05, 1.594579e-05, 1.11703e-05, 7.731369e-06, 6.559928e-06, 
    5.675095e-06, 5.070492e-06, 4.862366e-06, 5.130104e-06, 5.310943e-06, 
    5.372897e-06, 6.120258e-06, 7.926279e-06, 9.26028e-06, 1.042526e-05, 
    1.143812e-05, 1.370033e-05, 1.440072e-05, 1.510068e-05,
  8.129346e-06, 8.129346e-06, 8.129346e-06, 8.129346e-06, 8.129346e-06, 
    8.129346e-06, 8.129346e-06, 7.850588e-06, 7.850588e-06, 7.850588e-06, 
    7.850588e-06, 7.850588e-06, 7.850588e-06, 7.850588e-06, 8.65819e-06, 
    8.65819e-06, 8.65819e-06, 8.65819e-06, 8.65819e-06, 8.65819e-06, 
    8.65819e-06, 8.524074e-06, 8.524074e-06, 8.524074e-06, 8.524074e-06, 
    8.524074e-06, 8.524074e-06, 8.524074e-06, 8.129346e-06,
  7.850933e-06, 8.773354e-06, 1.076125e-05, 1.266633e-05, 1.337158e-05, 
    1.263073e-05, 1.03937e-05, 9.0487e-06, 8.558112e-06, 5.999753e-06, 
    5.009843e-06, 5.437528e-06, 5.906003e-06, 6.114904e-06, 7.118002e-06, 
    8.284441e-06, 8.393941e-06, 8.912157e-06, 9.567887e-06, 9.997781e-06, 
    1.062e-05, 1.059105e-05, 1.08089e-05, 1.039344e-05, 1.031039e-05, 
    1.020682e-05, 9.730852e-06, 8.756603e-06, 8.306309e-06,
  1.343629e-05, 1.093519e-05, 1.341319e-05, 1.611435e-05, 2.18447e-05, 
    2.68613e-05, 1.813705e-05, 1.499632e-05, 1.39193e-05, 1.349755e-05, 
    1.301738e-05, 1.29419e-05, 1.479683e-05, 1.717636e-05, 1.932172e-05, 
    2.390429e-05, 2.569344e-05, 2.840785e-05, 2.899749e-05, 2.828519e-05, 
    2.938063e-05, 2.999658e-05, 3.280631e-05, 3.404761e-05, 3.419923e-05, 
    3.300572e-05, 3.111488e-05, 2.590394e-05, 1.967624e-05,
  9.491881e-05, 9.301825e-05, 8.343404e-05, 8.497998e-05, 9.462951e-05, 
    9.585283e-05, 9.192296e-05, 8.43441e-05, 6.525939e-05, 5.796975e-05, 
    5.716276e-05, 7.626936e-05, 9.893369e-05, 0.000166019, 0.0002270486, 
    0.0002485486, 0.0001977837, 0.0001510141, 0.0001207431, 9.452536e-05, 
    8.644429e-05, 0.0001024645, 0.0001071233, 0.0001247806, 0.0001448378, 
    0.0001414304, 0.0001206338, 0.0001059736, 9.34836e-05,
  0.0004307971, 0.0003510042, 0.0003452188, 0.000411556, 0.0005790244, 
    0.0006742704, 0.0005925534, 0.0005331404, 0.0004899453, 0.0004708522, 
    0.0004479914, 0.0006375181, 0.001164099, 0.001900302, 0.002318537, 
    0.002523928, 0.002008745, 0.001140284, 0.0006330175, 0.0004692086, 
    0.0004546789, 0.0005253222, 0.0005845767, 0.0006525081, 0.0006053625, 
    0.000574838, 0.0005350175, 0.0004958917, 0.0004748,
  0.002294396, 0.002541481, 0.003187524, 0.003696497, 0.003118337, 
    0.003081861, 0.003486013, 0.003524601, 0.003088613, 0.004609293, 
    0.008566282, 0.01151455, 0.01444292, 0.009790765, 0.01447449, 0.01414621, 
    0.009313934, 0.006013905, 0.003946988, 0.002569159, 0.002564097, 
    0.003057034, 0.002340098, 0.002835533, 0.004338397, 0.003699351, 
    0.002845126, 0.002731493, 0.002280312,
  0.02399371, 0.0345671, 0.03892901, 0.03388855, 0.02094049, 0.0288769, 
    0.06816449, 0.1113333, 0.1396803, 0.2258212, 0.2322663, 0.1868875, 
    0.1251694, 0.08251632, 0.06026765, 0.03601779, 0.02447734, 0.01346765, 
    0.009548972, 0.01306605, 0.01688105, 0.01881786, 0.02187976, 0.03015072, 
    0.04056858, 0.03601918, 0.02370502, 0.01930788, 0.0202958,
  0.1492908, 0.2099547, 0.224276, 0.1762363, 0.1413892, 0.1816424, 0.2972517, 
    0.4576443, 0.6611061, 1.039862, 1.092166, 0.7640465, 0.4609886, 
    0.2955933, 0.1943562, 0.1226534, 0.0655122, 0.03445587, 0.02913085, 
    0.03052876, 0.05172355, 0.09133168, 0.144794, 0.2257421, 0.2449572, 
    0.1933188, 0.09817124, 0.08802502, 0.1221512,
  0.3681111, 0.3480568, 0.286389, 0.2413776, 0.2685845, 0.3596581, 0.5326987, 
    0.6493213, 0.8500754, 1.115179, 1.256101, 1.107509, 0.6824631, 0.5077117, 
    0.3612491, 0.260091, 0.1790856, 0.1237763, 0.09820586, 0.09124728, 
    0.09488494, 0.1389597, 0.2863734, 0.4864733, 0.5639279, 0.383544, 
    0.1512055, 0.1753152, 0.2888417,
  0.3635964, 0.4200625, 0.3719551, 0.2940368, 0.2853142, 0.3225457, 
    0.4427718, 0.5384439, 0.7087657, 0.8867304, 0.845242, 0.6926674, 
    0.4542029, 0.3798825, 0.3267584, 0.2697356, 0.2341989, 0.1894178, 
    0.1534476, 0.1260337, 0.1359456, 0.1839075, 0.2345806, 0.3174624, 
    0.268124, 0.2461666, 0.2044819, 0.1862619, 0.2497026,
  0.2557167, 0.3701183, 0.4168488, 0.5417352, 0.574053, 0.6355011, 0.8001335, 
    0.7508568, 0.9890171, 0.8255445, 0.6622556, 0.513077, 0.425172, 0.341121, 
    0.2652973, 0.2145445, 0.1639254, 0.1578737, 0.1623653, 0.1255601, 
    0.1223464, 0.1296392, 0.1426628, 0.1347585, 0.09958019, 0.1020701, 
    0.1458725, 0.1564799, 0.2113754,
  0.164882, 0.2582845, 0.4386607, 0.6585239, 0.7863477, 0.863685, 1.055773, 
    1.08052, 1.030878, 0.607838, 0.4444049, 0.362592, 0.2687304, 0.1867487, 
    0.1185353, 0.08680242, 0.07058089, 0.06700169, 0.07444715, 0.08516593, 
    0.07667527, 0.05524118, 0.05927657, 0.05457333, 0.04745113, 0.0484079, 
    0.05831851, 0.08148959, 0.1115403,
  0.06307267, 0.1124748, 0.1539009, 0.2294403, 0.2574833, 0.2877817, 
    0.3698564, 0.4173728, 0.3097955, 0.1846617, 0.112421, 0.07230031, 
    0.06023282, 0.05214253, 0.03077295, 0.01722783, 0.01381518, 0.01632989, 
    0.01778552, 0.02227876, 0.02976158, 0.02096637, 0.01577839, 0.01392255, 
    0.01277171, 0.01164279, 0.01040683, 0.01428252, 0.03550841,
  0.008244531, 0.01523123, 0.01727285, 0.02167013, 0.02406089, 0.01894471, 
    0.02483917, 0.02890931, 0.02353797, 0.01528256, 0.01265673, 0.01253217, 
    0.01598659, 0.01005831, 0.008089394, 0.005780953, 0.003511617, 
    0.003142346, 0.003678383, 0.005015804, 0.007515417, 0.005420886, 
    0.003736468, 0.002349746, 0.002386144, 0.002047906, 0.001477129, 
    0.00148523, 0.003182047,
  0.0005090595, 0.0008591739, 0.001641915, 0.002472805, 0.001899615, 
    0.001409458, 0.001459929, 0.001474801, 0.001858875, 0.002241099, 
    0.002859347, 0.0028823, 0.00254007, 0.002893603, 0.002067815, 
    0.001587196, 0.001226546, 0.001048998, 0.001053132, 0.001047889, 
    0.001080499, 0.0008674318, 0.0006153531, 0.0005146725, 0.0004901303, 
    0.0006624737, 0.0006551889, 0.0006020289, 0.0005999665,
  0.0001829722, 0.0002666889, 0.0004149197, 0.0005362694, 0.0005754373, 
    0.0006677055, 0.0006402332, 0.0005967416, 0.0005164318, 0.0003790846, 
    0.0003991842, 0.0004197805, 0.0004462549, 0.0003807702, 0.0003939225, 
    0.000296371, 0.000290028, 0.0002562483, 0.0002804101, 0.000259566, 
    0.0002115484, 0.0001723124, 0.0001375688, 0.0001443855, 0.0001928548, 
    0.0002178703, 0.000256472, 0.0002786433, 0.0002412536,
  8.073515e-05, 7.227701e-05, 9.253401e-05, 0.0001186983, 0.0001991801, 
    0.0001949464, 0.0001672961, 0.0001464655, 0.0001442945, 0.0001267643, 
    0.0001167605, 9.173074e-05, 7.166096e-05, 8.016695e-05, 8.748103e-05, 
    8.073197e-05, 8.308091e-05, 8.443382e-05, 9.171006e-05, 8.903474e-05, 
    7.374978e-05, 5.47698e-05, 5.704823e-05, 5.795625e-05, 6.604088e-05, 
    8.184673e-05, 0.0001080961, 0.0001084158, 9.23378e-05,
  4.586608e-05, 4.926444e-05, 5.202076e-05, 5.392388e-05, 5.421723e-05, 
    6.840485e-05, 7.232126e-05, 7.019097e-05, 6.664434e-05, 6.373004e-05, 
    6.399232e-05, 6.043127e-05, 4.114956e-05, 3.152174e-05, 2.818541e-05, 
    2.236157e-05, 1.807633e-05, 1.460521e-05, 1.814738e-05, 2.01985e-05, 
    2.534226e-05, 2.943936e-05, 3.00091e-05, 3.294954e-05, 3.524811e-05, 
    3.910082e-05, 4.524039e-05, 4.506049e-05, 4.486337e-05,
  3.785294e-05, 3.785294e-05, 3.785294e-05, 3.785294e-05, 3.785294e-05, 
    3.785294e-05, 3.785294e-05, 3.66391e-05, 3.66391e-05, 3.66391e-05, 
    3.66391e-05, 3.66391e-05, 3.66391e-05, 3.66391e-05, 3.835928e-05, 
    3.835928e-05, 3.835928e-05, 3.835928e-05, 3.835928e-05, 3.835928e-05, 
    3.835928e-05, 4.12934e-05, 4.12934e-05, 4.12934e-05, 4.12934e-05, 
    4.12934e-05, 4.12934e-05, 4.12934e-05, 3.785294e-05,
  3.667513e-05, 3.924871e-05, 4.567593e-05, 5.317755e-05, 5.75594e-05, 
    5.330252e-05, 4.254732e-05, 3.328822e-05, 3.107276e-05, 2.315224e-05, 
    1.684366e-05, 1.651256e-05, 2.073367e-05, 2.451096e-05, 2.933395e-05, 
    3.230652e-05, 3.35503e-05, 3.641284e-05, 3.817375e-05, 3.997239e-05, 
    4.55176e-05, 4.541859e-05, 4.911261e-05, 4.948404e-05, 4.530124e-05, 
    4.218243e-05, 4.079325e-05, 4.188512e-05, 3.709177e-05,
  5.051922e-05, 3.203779e-05, 3.659061e-05, 5.208247e-05, 0.0001045948, 
    0.0001197235, 7.286618e-05, 5.374059e-05, 4.618564e-05, 4.105059e-05, 
    4.142559e-05, 4.243359e-05, 5.168128e-05, 5.359502e-05, 5.55768e-05, 
    6.146507e-05, 7.014183e-05, 7.340338e-05, 7.162825e-05, 8.144852e-05, 
    8.959598e-05, 0.000110456, 0.0001306104, 0.0001298055, 0.0001240522, 
    0.0001204341, 0.0001045073, 8.770431e-05, 6.992434e-05,
  0.0002827593, 0.0003046642, 0.0002768324, 0.0002837613, 0.0003220941, 
    0.0003160039, 0.0002831677, 0.0002570481, 0.0002185276, 0.0001954088, 
    0.0001924982, 0.0002106477, 0.0003031467, 0.0004173562, 0.000715015, 
    0.0007887221, 0.0006217568, 0.0004681219, 0.0003756648, 0.0002977891, 
    0.0002859502, 0.0003442071, 0.0003553526, 0.0003990655, 0.0004443778, 
    0.0004518711, 0.0004587965, 0.0003847319, 0.0003343126,
  0.001305501, 0.001116814, 0.001078864, 0.001171451, 0.001742032, 
    0.002255795, 0.001927203, 0.001702605, 0.00152196, 0.001366198, 
    0.001368123, 0.001717854, 0.004494698, 0.006419723, 0.008642692, 
    0.009241073, 0.006499079, 0.003505848, 0.002101872, 0.001624402, 
    0.001775643, 0.001844291, 0.001969253, 0.002175514, 0.001887821, 
    0.001667465, 0.001534722, 0.001379927, 0.001311135,
  0.007087128, 0.007556155, 0.009972622, 0.0137031, 0.01268573, 0.01084895, 
    0.01115599, 0.01005535, 0.0098408, 0.01481014, 0.03148848, 0.05017845, 
    0.04991813, 0.03440156, 0.05181674, 0.05479342, 0.03655199, 0.02341601, 
    0.01519207, 0.009815079, 0.007279731, 0.008175321, 0.006538269, 
    0.007830145, 0.01018425, 0.009261695, 0.007222014, 0.007371406, 
    0.007391428,
  0.07214225, 0.141107, 0.1943605, 0.189835, 0.1138897, 0.07660191, 
    0.1732595, 0.2866161, 0.4066054, 0.619807, 0.7292686, 0.6054723, 
    0.4137043, 0.2922981, 0.2055455, 0.1216671, 0.08781539, 0.05279282, 
    0.02853594, 0.02601643, 0.04087114, 0.05494991, 0.06061758, 0.08730124, 
    0.1275665, 0.1503888, 0.09798217, 0.06889816, 0.06003853,
  0.6017647, 0.9716393, 1.10124, 0.8489406, 0.5593815, 0.4897842, 0.6854569, 
    1.058074, 1.655901, 2.425157, 2.653533, 2.028147, 1.130268, 0.7474961, 
    0.5233094, 0.3609463, 0.2361705, 0.1228493, 0.09012967, 0.07706526, 
    0.09059057, 0.1943646, 0.4325985, 0.9279484, 1.377347, 1.136283, 
    0.4378668, 0.2622712, 0.4138399,
  1.12407, 1.722147, 1.13671, 0.849202, 0.7568559, 0.8599304, 1.171951, 
    1.537799, 2.019667, 2.505956, 2.643166, 2.326054, 1.368444, 0.9860991, 
    0.7359958, 0.5581379, 0.4310992, 0.3091205, 0.2530378, 0.2282726, 
    0.2026577, 0.2268843, 0.5453699, 1.214262, 2.104385, 1.784924, 0.6307526, 
    0.4452299, 0.7798264,
  0.9686348, 1.476695, 1.188795, 0.83332, 0.7543529, 0.8937687, 1.194791, 
    1.64011, 2.110323, 2.242568, 1.893954, 1.353684, 0.7613827, 0.6679184, 
    0.5636933, 0.4854996, 0.4382088, 0.4119546, 0.3516378, 0.2941775, 
    0.2766919, 0.3147368, 0.4984457, 0.6941499, 0.8264392, 0.7501405, 
    0.5913385, 0.5105256, 0.7160136,
  0.6808956, 0.9598599, 1.127018, 1.224681, 1.351396, 1.852152, 2.370403, 
    2.795481, 2.989189, 2.13495, 1.458858, 0.9755213, 0.8121945, 0.639225, 
    0.5447406, 0.4525246, 0.3784603, 0.3763043, 0.3914226, 0.3695178, 
    0.408076, 0.3902099, 0.4680354, 0.3944268, 0.2913473, 0.3250046, 
    0.4617269, 0.5540213, 0.5879531,
  0.4039363, 0.6272584, 1.066224, 1.587264, 2.092087, 2.502613, 3.460428, 
    3.469731, 3.092592, 1.985431, 1.358279, 0.9052042, 0.7017914, 0.5248543, 
    0.3448135, 0.2237386, 0.1858399, 0.1827118, 0.2442192, 0.3628989, 
    0.3920824, 0.2170917, 0.2062122, 0.1567008, 0.1211793, 0.117176, 
    0.1565986, 0.2338522, 0.3172978,
  0.147236, 0.2972832, 0.483439, 0.6892799, 0.8441941, 0.9318373, 1.359638, 
    1.614628, 1.111733, 0.6072319, 0.3697904, 0.2730609, 0.2312921, 
    0.1765491, 0.1010432, 0.05146149, 0.03594503, 0.04327397, 0.06084819, 
    0.08775602, 0.129685, 0.07089231, 0.06726343, 0.04547818, 0.03817711, 
    0.02969518, 0.02096065, 0.02446599, 0.06951594,
  0.01678267, 0.03551867, 0.04234381, 0.05943808, 0.08386677, 0.07347926, 
    0.07911529, 0.1021785, 0.09071065, 0.05821932, 0.04549532, 0.05047328, 
    0.06473634, 0.0423975, 0.03106879, 0.02261751, 0.01165673, 0.009249956, 
    0.01075794, 0.01541727, 0.02456146, 0.02001463, 0.01227929, 0.008350641, 
    0.006815255, 0.007478561, 0.005190868, 0.005615376, 0.00600728,
  0.001586531, 0.001867272, 0.003556208, 0.006728166, 0.006255106, 
    0.003881961, 0.003453224, 0.003743457, 0.005034473, 0.008632094, 
    0.01134204, 0.01159288, 0.009331797, 0.009927595, 0.007384156, 
    0.004512278, 0.004323582, 0.003906883, 0.00294769, 0.002948673, 
    0.003152844, 0.002663025, 0.001965007, 0.001538637, 0.001619819, 
    0.002029697, 0.002199526, 0.0017853, 0.001564873,
  0.0004388596, 0.0004835861, 0.0007599944, 0.001298803, 0.001580057, 
    0.001936566, 0.002070138, 0.00151419, 0.001372467, 0.001283893, 
    0.001181831, 0.001464579, 0.001461309, 0.00116564, 0.001111428, 
    0.001112721, 0.000959307, 0.00090774, 0.0009191032, 0.0007855843, 
    0.0006897806, 0.0006300037, 0.0004461199, 0.0004198057, 0.0004783058, 
    0.0006257372, 0.0007661842, 0.0007095023, 0.0005646834,
  0.0002072845, 0.0001718423, 0.0002208017, 0.0002268191, 0.0003385801, 
    0.0004514151, 0.0004926474, 0.0004391729, 0.0004024089, 0.0004179216, 
    0.0003850091, 0.0002851144, 0.0002402371, 0.0002375531, 0.0002471076, 
    0.0003207558, 0.0003531923, 0.0003803376, 0.000371913, 0.0003598423, 
    0.0002988822, 0.0002045801, 0.0002105773, 0.000200571, 0.0002208159, 
    0.0002548529, 0.0003248239, 0.0003312042, 0.000250244,
  0.0001204569, 0.0001121865, 0.0001188674, 0.0001250304, 0.0001228164, 
    0.0001510236, 0.0001796161, 0.0002020143, 0.0002017849, 0.0002023481, 
    0.0002031861, 0.0002004049, 0.0001439859, 0.0001083747, 9.012462e-05, 
    6.97779e-05, 7.02305e-05, 6.683197e-05, 7.827315e-05, 9.211057e-05, 
    0.0001071211, 0.0001075886, 0.0001060936, 0.0001235762, 0.0001318298, 
    0.0001423144, 0.0001505998, 0.0001335977, 0.0001249376,
  0.00016837, 0.00016837, 0.00016837, 0.00016837, 0.00016837, 0.00016837, 
    0.00016837, 0.0001441926, 0.0001441926, 0.0001441926, 0.0001441926, 
    0.0001441926, 0.0001441926, 0.0001441926, 0.0001580813, 0.0001580813, 
    0.0001580813, 0.0001580813, 0.0001580813, 0.0001580813, 0.0001580813, 
    0.0001663036, 0.0001663036, 0.0001663036, 0.0001663036, 0.0001663036, 
    0.0001663036, 0.0001663036, 0.00016837,
  0.000165512, 0.0001391753, 0.0001713224, 0.0002337921, 0.0002738443, 
    0.000248737, 0.0001684698, 0.0001270242, 0.0001033003, 7.844826e-05, 
    5.726703e-05, 5.019453e-05, 5.782908e-05, 7.289305e-05, 8.906325e-05, 
    0.0001062467, 0.0001431808, 0.0001564087, 0.0001417237, 0.0001386724, 
    0.0001618335, 0.0001669706, 0.0001924493, 0.0002098583, 0.0001928876, 
    0.000174196, 0.0001699105, 0.0001850393, 0.0001680838,
  0.0001663305, 0.0001063483, 0.0001282731, 0.0002044238, 0.0004705527, 
    0.0004700952, 0.0002576692, 0.0001463809, 0.0001180368, 0.0001045825, 
    0.0001123155, 0.0001182925, 0.0001458874, 0.0001637551, 0.0001553086, 
    0.0001718352, 0.0001974004, 0.000200762, 0.000183741, 0.0001979446, 
    0.0002646864, 0.0003575333, 0.0004178466, 0.00041653, 0.0004046582, 
    0.0003705871, 0.0003285731, 0.000283849, 0.0002246687,
  0.0006899168, 0.0006316947, 0.0006815236, 0.0007521592, 0.0008556612, 
    0.0008100963, 0.0007249428, 0.0006195468, 0.0005638495, 0.0004542593, 
    0.0004219888, 0.0004226506, 0.0005272759, 0.0008479965, 0.001413578, 
    0.001643333, 0.001480805, 0.001179705, 0.0009353276, 0.0008635022, 
    0.0007964412, 0.0008468759, 0.0009107724, 0.001121897, 0.001177768, 
    0.001214993, 0.001315179, 0.001058095, 0.0008873872,
  0.003489165, 0.003168552, 0.003192662, 0.003412756, 0.00537108, 
    0.007399887, 0.005690995, 0.005142569, 0.004590473, 0.004025622, 
    0.003650321, 0.004653043, 0.01201189, 0.02036655, 0.02215812, 0.02592278, 
    0.01854275, 0.009553579, 0.005747488, 0.004540564, 0.004914972, 
    0.00530802, 0.005559372, 0.00576199, 0.005341088, 0.004618384, 
    0.004034105, 0.00362065, 0.00327046,
  0.02335357, 0.01878341, 0.02761065, 0.03696054, 0.04421724, 0.04232745, 
    0.04117569, 0.02964457, 0.0266787, 0.03955682, 0.08252606, 0.1311782, 
    0.1216236, 0.09048829, 0.1153304, 0.126277, 0.09301687, 0.06610774, 
    0.04563421, 0.03211471, 0.01956331, 0.01923232, 0.01859046, 0.01985583, 
    0.02328928, 0.01966397, 0.01836839, 0.01920175, 0.021095,
  0.1992937, 0.451212, 0.7076672, 0.691013, 0.3431293, 0.2442824, 0.3480552, 
    0.4993435, 0.7592334, 1.15038, 1.391662, 1.227324, 0.8441944, 0.6226609, 
    0.4240949, 0.2733292, 0.2108809, 0.1490919, 0.07970595, 0.05462457, 
    0.06890182, 0.09329877, 0.1327094, 0.1895781, 0.3495108, 0.5051624, 
    0.3269144, 0.2510042, 0.1594933,
  1.582673, 2.674844, 2.776267, 2.170141, 1.32113, 1.028233, 1.196087, 
    1.68107, 2.489181, 3.553141, 3.97918, 3.357733, 1.919539, 1.169283, 
    0.8793969, 0.6594657, 0.4807527, 0.2961062, 0.199419, 0.1605825, 
    0.1643162, 0.3251894, 1.025942, 2.381774, 4.092618, 3.266107, 1.278084, 
    0.605508, 0.9256855,
  2.390531, 4.554895, 3.257707, 1.98106, 1.572688, 1.542977, 1.891281, 
    2.431709, 3.16389, 3.359123, 3.612141, 3.386017, 2.021439, 1.372873, 
    1.065812, 0.8206854, 0.6699973, 0.5165639, 0.440612, 0.4017841, 
    0.3540309, 0.3582804, 0.9124247, 2.549137, 4.889712, 4.194527, 1.676127, 
    0.9111168, 1.512637,
  2.194782, 3.965358, 2.954849, 1.805257, 1.589315, 1.882204, 2.311864, 
    3.007147, 3.998283, 4.133033, 2.675861, 2.017249, 1.023944, 0.8267136, 
    0.7354322, 0.6324973, 0.5778536, 0.5883304, 0.5646771, 0.5393164, 
    0.4897481, 0.5024323, 0.8614046, 1.562347, 2.197399, 1.984666, 1.415594, 
    1.193959, 1.547032,
  1.783831, 2.314875, 2.471797, 2.208293, 2.573545, 3.153931, 3.99552, 
    4.566509, 4.604065, 3.321661, 2.128936, 1.322278, 0.9756356, 0.8482354, 
    0.7644463, 0.6753438, 0.6034352, 0.6116719, 0.6653852, 0.7428091, 
    0.8848096, 1.048733, 1.373896, 1.148432, 0.955556, 1.064416, 1.291656, 
    1.524758, 1.750365,
  0.8976769, 1.192101, 1.762636, 2.57345, 3.293737, 4.209626, 5.726836, 
    5.769657, 4.996045, 3.482721, 2.512033, 1.587717, 1.24773, 1.011681, 
    0.7666786, 0.5264639, 0.401476, 0.3780108, 0.4960116, 0.8778399, 
    1.135021, 0.6942217, 0.5958711, 0.3689077, 0.3165808, 0.3102886, 
    0.456267, 0.8726956, 0.8554353,
  0.2633767, 0.5259087, 0.9021079, 1.215916, 1.474112, 1.696823, 2.891241, 
    3.38351, 2.434121, 1.444856, 0.9297882, 0.7364658, 0.5550811, 0.4327704, 
    0.2700239, 0.1595236, 0.103069, 0.09690175, 0.1386559, 0.2624375, 
    0.3212393, 0.2093689, 0.2577006, 0.1759795, 0.133053, 0.08692144, 
    0.05103138, 0.06211286, 0.1218875,
  0.02421259, 0.05421808, 0.07992616, 0.1263375, 0.2062116, 0.1882041, 
    0.1744543, 0.2419498, 0.2369336, 0.1492884, 0.1294694, 0.1554315, 
    0.1874354, 0.1304714, 0.09040271, 0.06614683, 0.04144812, 0.02632768, 
    0.0294701, 0.03918401, 0.06137489, 0.05638298, 0.03715173, 0.02466672, 
    0.02525262, 0.03348463, 0.02775976, 0.01767129, 0.01426943,
  0.00378228, 0.00341105, 0.006243026, 0.01112427, 0.01543662, 0.008552802, 
    0.006658855, 0.00684691, 0.01003942, 0.0213315, 0.02827938, 0.03638616, 
    0.02868041, 0.02933256, 0.02280753, 0.01231994, 0.01212379, 0.01223741, 
    0.00929046, 0.008386212, 0.008680094, 0.007651508, 0.005748461, 
    0.004193331, 0.004509538, 0.005875901, 0.007274854, 0.005366109, 
    0.003973627,
  0.001106739, 0.0009862018, 0.001206319, 0.002463821, 0.003330164, 
    0.004648288, 0.005125428, 0.003210237, 0.00255233, 0.003244757, 
    0.003034778, 0.004299165, 0.004393824, 0.003841809, 0.003406735, 
    0.003254194, 0.002847159, 0.002773449, 0.002486611, 0.002407466, 
    0.002114762, 0.001842553, 0.001269963, 0.001124897, 0.001301725, 
    0.00165462, 0.002005938, 0.001696896, 0.001222963,
  0.0004890177, 0.000394512, 0.0004215276, 0.000436689, 0.0005810553, 
    0.0008508648, 0.0009527034, 0.001075479, 0.0009686889, 0.0009631212, 
    0.000934021, 0.0008443895, 0.0006332655, 0.0006894709, 0.0006650381, 
    0.0009835977, 0.001151457, 0.001277244, 0.001226309, 0.001185743, 
    0.0008828157, 0.0007553506, 0.0005836467, 0.0005196601, 0.0006263838, 
    0.000662775, 0.0007304055, 0.0007448054, 0.0006014354,
  0.0003572052, 0.0003250858, 0.000312219, 0.0003246238, 0.0003415492, 
    0.00037004, 0.0004299015, 0.0004865935, 0.0005379991, 0.0005706383, 
    0.0005917365, 0.0005684409, 0.0004409023, 0.0003207796, 0.000293429, 
    0.0003397384, 0.0003429592, 0.0003378708, 0.0003741212, 0.0003603436, 
    0.0003486863, 0.0003553861, 0.0003756338, 0.0003825689, 0.0004141283, 
    0.0004295752, 0.0004052588, 0.0003953037, 0.0003774783,
  0.001031774, 0.001031774, 0.001031774, 0.001031774, 0.001031774, 
    0.001031774, 0.001031774, 0.0008537697, 0.0008537697, 0.0008537697, 
    0.0008537697, 0.0008537697, 0.0008537697, 0.0008537697, 0.0009564271, 
    0.0009564271, 0.0009564271, 0.0009564271, 0.0009564271, 0.0009564271, 
    0.0009564271, 0.00103126, 0.00103126, 0.00103126, 0.00103126, 0.00103126, 
    0.00103126, 0.00103126, 0.001031774,
  0.001068673, 0.001042599, 0.001115025, 0.001258979, 0.001435656, 
    0.001310868, 0.0008204622, 0.0004906079, 0.0003346064, 0.000282052, 
    0.0002218493, 0.0001726206, 0.0001715889, 0.0002487283, 0.0004063312, 
    0.0006528941, 0.0008836457, 0.0009179583, 0.0005726173, 0.000733137, 
    0.0007765456, 0.0007600301, 0.0008137383, 0.00106555, 0.001063555, 
    0.0008749487, 0.0007217196, 0.0007428895, 0.001077203,
  0.0005443341, 0.0004196659, 0.0004951573, 0.0007791163, 0.002676307, 
    0.003999679, 0.001074475, 0.0004355203, 0.0003229448, 0.0002978295, 
    0.0003056395, 0.0003150718, 0.0003984557, 0.000512152, 0.0005422132, 
    0.0005487893, 0.0005874104, 0.0005920984, 0.0005489244, 0.0006162591, 
    0.0008514477, 0.001153519, 0.001354225, 0.001335705, 0.001355564, 
    0.001218654, 0.001101564, 0.0008869211, 0.0006746058,
  0.00161799, 0.001298227, 0.001575636, 0.001794496, 0.002142755, 
    0.003787016, 0.002632086, 0.001606434, 0.001262928, 0.0009648316, 
    0.0008143238, 0.0009078305, 0.00116876, 0.001645431, 0.002712335, 
    0.003917215, 0.004144295, 0.003514034, 0.002406468, 0.002003389, 
    0.001828189, 0.002128209, 0.002429938, 0.002982398, 0.003439456, 
    0.003761365, 0.003434671, 0.002667231, 0.002091944,
  0.008732111, 0.008278049, 0.0087434, 0.009622669, 0.01945272, 0.02631613, 
    0.02042215, 0.01718776, 0.0160636, 0.01372572, 0.01166997, 0.01234036, 
    0.02535797, 0.04514374, 0.0488708, 0.05688674, 0.04501217, 0.02674186, 
    0.01598274, 0.01149844, 0.01291572, 0.01398238, 0.01498025, 0.01452369, 
    0.01273534, 0.009654922, 0.009394018, 0.008846916, 0.00837722,
  0.06633552, 0.04841735, 0.07815579, 0.09754978, 0.1181835, 0.1157162, 
    0.1144658, 0.0870047, 0.06386629, 0.08639248, 0.1700594, 0.2351577, 
    0.2244062, 0.1769247, 0.2004196, 0.2321832, 0.1959175, 0.1516418, 
    0.1125824, 0.08309094, 0.0497362, 0.04780027, 0.04727966, 0.03981712, 
    0.04592095, 0.03901694, 0.04052625, 0.06166229, 0.05719281,
  0.4473082, 1.07325, 1.672141, 1.458652, 0.7407532, 0.5268633, 0.6406925, 
    0.759617, 1.110987, 1.714036, 2.048965, 1.921446, 1.372537, 0.9715598, 
    0.6827516, 0.4605697, 0.3712128, 0.3160436, 0.1896605, 0.1182394, 
    0.1200548, 0.1329824, 0.2066986, 0.3197435, 0.7735556, 1.182884, 
    0.8810959, 0.6505113, 0.4285741,
  2.767131, 4.864307, 4.666913, 3.597505, 2.307043, 1.662907, 1.669037, 
    2.150351, 3.050264, 4.241547, 4.836067, 4.239116, 2.613072, 1.527113, 
    1.180313, 0.9308224, 0.7240663, 0.5326359, 0.3666448, 0.2916947, 
    0.2895599, 0.5118006, 1.873918, 3.951726, 6.57283, 5.559466, 2.560007, 
    1.257911, 1.569728,
  4.121706, 8.331096, 6.574606, 3.491006, 2.410454, 2.040482, 2.434866, 
    3.098775, 4.126081, 3.917189, 3.957772, 4.030132, 2.536386, 1.598768, 
    1.265674, 1.006845, 0.8361932, 0.6908461, 0.6011873, 0.5746177, 0.515102, 
    0.5298491, 1.53418, 4.71952, 7.749079, 6.509078, 3.279446, 1.587752, 
    2.394914,
  4.044291, 8.006962, 6.100003, 3.138576, 2.384378, 2.465086, 3.011395, 
    3.829971, 5.498542, 6.019589, 3.029078, 2.451708, 1.17728, 0.8931909, 
    0.8198912, 0.7244392, 0.6705971, 0.7241648, 0.7526165, 0.8107545, 
    0.7597101, 0.8133609, 1.367083, 3.237426, 4.486243, 3.880793, 2.627648, 
    2.212155, 2.831324,
  4.080462, 5.377981, 4.704665, 3.46916, 3.490816, 3.931968, 4.816358, 
    5.416343, 5.543294, 4.026439, 2.432766, 1.541981, 1.082477, 0.9697003, 
    0.8734012, 0.8349865, 0.761956, 0.7983288, 0.9192455, 1.172105, 1.443925, 
    1.93277, 2.702529, 2.689901, 2.193034, 2.256885, 2.670381, 3.173059, 
    4.041836,
  1.697021, 2.000406, 2.629664, 3.541032, 4.354189, 5.403506, 6.95544, 
    7.36502, 6.630531, 4.692927, 3.267786, 2.152437, 1.63847, 1.415365, 
    1.235394, 0.9260232, 0.7111262, 0.6052015, 0.7557281, 1.355215, 2.29117, 
    1.612086, 1.288863, 0.7498978, 0.7209492, 0.7073352, 1.056536, 2.026446, 
    2.056452,
  0.4178821, 0.7624434, 1.246032, 1.593479, 1.950575, 2.390578, 4.079564, 
    4.856044, 3.594231, 2.634474, 1.777405, 1.416935, 1.114559, 0.8633634, 
    0.6415762, 0.4539752, 0.2727937, 0.2233862, 0.3002435, 0.5771337, 
    0.7195931, 0.5391458, 0.712488, 0.6319786, 0.442117, 0.2752855, 
    0.1738484, 0.1582426, 0.2059441,
  0.05230269, 0.07855133, 0.1233716, 0.2091259, 0.3683317, 0.3134263, 
    0.2922941, 0.4651977, 0.4593671, 0.2932945, 0.3360644, 0.3638894, 
    0.4267738, 0.3294063, 0.269149, 0.2159482, 0.1485246, 0.08945864, 
    0.08169878, 0.08117891, 0.1401947, 0.1573697, 0.1055906, 0.06959172, 
    0.1263723, 0.1789002, 0.146044, 0.07272983, 0.04785635,
  0.01262518, 0.0101342, 0.01217596, 0.01794206, 0.02484602, 0.0172027, 
    0.01124336, 0.01166972, 0.01469715, 0.03011621, 0.04673406, 0.09036306, 
    0.08449307, 0.0823236, 0.06056914, 0.03301524, 0.03684104, 0.03367272, 
    0.02823312, 0.02287009, 0.02182474, 0.02052363, 0.01559799, 0.01057008, 
    0.01241167, 0.02073447, 0.02679668, 0.02029661, 0.01345572,
  0.002750172, 0.002629437, 0.002899383, 0.003979492, 0.0056079, 0.008277092, 
    0.008131527, 0.00573563, 0.004454411, 0.005089817, 0.005477913, 
    0.008458578, 0.009805031, 0.008749222, 0.008114359, 0.007316949, 
    0.006811637, 0.006883421, 0.006533867, 0.006470772, 0.005561499, 
    0.004448923, 0.002998476, 0.002783418, 0.003299379, 0.004427329, 
    0.005486389, 0.003930492, 0.003058516,
  0.001364979, 0.001067172, 0.0009577473, 0.0009698138, 0.001108042, 
    0.001355549, 0.001617325, 0.001890731, 0.00173405, 0.001873618, 
    0.00199648, 0.001748995, 0.001662564, 0.002010047, 0.001702705, 
    0.002133253, 0.002425789, 0.003081071, 0.002964318, 0.002595627, 
    0.001834469, 0.001656694, 0.001507099, 0.001303355, 0.001601277, 
    0.001714285, 0.00189082, 0.00197535, 0.001549491,
  0.0008464536, 0.0007884985, 0.0006997939, 0.0006971427, 0.0007702506, 
    0.0008084697, 0.0008589646, 0.0009288711, 0.001041685, 0.001260434, 
    0.0014083, 0.001201147, 0.001021622, 0.0009574166, 0.000843964, 
    0.0009198987, 0.0009839715, 0.001021675, 0.001165065, 0.001122882, 
    0.0009863101, 0.0009719669, 0.0008871536, 0.0009172696, 0.0009808346, 
    0.000942986, 0.0008811041, 0.0009200537, 0.0008875026,
  0.007043442, 0.007043442, 0.007043442, 0.007043442, 0.007043442, 
    0.007043442, 0.007043442, 0.006161894, 0.006161894, 0.006161894, 
    0.006161894, 0.006161894, 0.006161894, 0.006161894, 0.0069004, 0.0069004, 
    0.0069004, 0.0069004, 0.0069004, 0.0069004, 0.0069004, 0.007193029, 
    0.007193029, 0.007193029, 0.007193029, 0.007193029, 0.007193029, 
    0.007193029, 0.007043442,
  0.006093835, 0.00683558, 0.007961246, 0.009020133, 0.01067477, 0.008121607, 
    0.004668175, 0.003308439, 0.001705178, 0.001159137, 0.000919585, 
    0.0007961576, 0.0007362107, 0.001550943, 0.002746505, 0.002363513, 
    0.00373935, 0.00435937, 0.004305048, 0.006284474, 0.00512011, 0.00459056, 
    0.004618353, 0.006714622, 0.006403288, 0.004401155, 0.003813896, 
    0.003403453, 0.005286539,
  0.002336703, 0.001885888, 0.002314215, 0.006056737, 0.019954, 0.02713751, 
    0.006180323, 0.001501283, 0.0009097088, 0.0009136815, 0.0009115225, 
    0.0008467659, 0.001239549, 0.002451658, 0.003178311, 0.002309683, 
    0.001635817, 0.001720589, 0.001790197, 0.002867308, 0.004044039, 
    0.005144894, 0.006849281, 0.00709098, 0.006881002, 0.00521075, 
    0.00431068, 0.003743858, 0.002818847,
  0.004538618, 0.003861595, 0.004352657, 0.004897338, 0.01375428, 0.03255035, 
    0.01929844, 0.006250222, 0.003423261, 0.002576654, 0.002138807, 
    0.002339408, 0.003069327, 0.004438773, 0.008185873, 0.01203155, 
    0.0123291, 0.009593821, 0.006575432, 0.00496937, 0.004962435, 
    0.006359018, 0.00832442, 0.00874025, 0.0102051, 0.01097304, 0.009830103, 
    0.007794047, 0.005955348,
  0.02404609, 0.02132165, 0.02302885, 0.02773257, 0.06081837, 0.08930902, 
    0.08894128, 0.05951571, 0.05345252, 0.04378735, 0.03618684, 0.03369973, 
    0.06097103, 0.09858387, 0.1043804, 0.1308361, 0.09806651, 0.06546688, 
    0.04064098, 0.03176295, 0.03693971, 0.03682569, 0.04157572, 0.03609778, 
    0.03190842, 0.0243166, 0.0257348, 0.02529908, 0.02553952,
  0.1808721, 0.1415983, 0.2056941, 0.2351603, 0.2736468, 0.2655894, 
    0.2672913, 0.2605431, 0.1886898, 0.1778202, 0.2782082, 0.3682909, 
    0.379869, 0.3068608, 0.3351571, 0.4017023, 0.3645213, 0.3083599, 
    0.2495908, 0.2011115, 0.140536, 0.1183957, 0.1118925, 0.07581889, 
    0.08507358, 0.1024, 0.1304303, 0.20836, 0.1793497,
  0.8691427, 1.907778, 2.786379, 2.319654, 1.297457, 0.9952564, 1.010763, 
    1.037117, 1.370445, 2.155226, 2.574117, 2.48908, 1.850242, 1.283427, 
    0.9122134, 0.6781116, 0.5892478, 0.5352147, 0.404083, 0.2671047, 
    0.2196657, 0.2252232, 0.3216917, 0.4985853, 1.525463, 2.192402, 1.775534, 
    1.271708, 0.9243091,
  4.012699, 7.220873, 6.721888, 4.997764, 3.233349, 2.338382, 2.061949, 
    2.521517, 3.431282, 4.596916, 5.399055, 4.749897, 3.100329, 1.851424, 
    1.432529, 1.111887, 0.9404809, 0.7365489, 0.5516142, 0.4575856, 
    0.4598268, 0.7745771, 2.726531, 5.193817, 8.274952, 7.241297, 4.090118, 
    2.217302, 2.401935,
  6.182646, 11.94391, 10.19618, 5.223026, 3.028301, 2.220754, 2.597105, 
    3.401042, 4.743326, 4.34208, 4.090907, 4.373701, 2.804376, 1.65955, 
    1.338339, 1.102554, 0.929179, 0.8012334, 0.6945722, 0.7056805, 0.6702211, 
    0.7407602, 2.549276, 7.556787, 10.73254, 8.683981, 4.707904, 2.505005, 
    3.520967,
  6.169339, 12.63805, 9.975681, 4.675555, 2.857003, 2.698483, 3.148018, 
    3.9382, 6.375113, 7.509053, 3.213844, 2.622215, 1.194286, 0.8906807, 
    0.8310924, 0.7814986, 0.7292362, 0.8203993, 0.8548489, 0.9906834, 
    1.06831, 1.16468, 2.101697, 5.793824, 7.400343, 5.862851, 4.02346, 
    3.464642, 4.429479,
  7.299016, 9.654945, 7.726424, 4.746104, 4.042722, 4.189593, 5.086056, 
    5.813767, 6.076966, 4.411034, 2.563883, 1.556677, 1.123353, 1.038203, 
    0.9174342, 0.912791, 0.8585632, 0.9252438, 1.125098, 1.544374, 1.982923, 
    2.697839, 3.937804, 4.78568, 3.869346, 3.831774, 4.362123, 5.543949, 
    6.703146,
  2.830426, 3.229064, 4.02828, 4.73637, 5.253286, 6.213503, 7.587559, 
    8.264569, 7.915987, 5.520363, 3.790765, 2.580563, 1.945395, 1.695721, 
    1.548276, 1.27463, 1.01373, 0.88258, 1.005064, 1.67102, 2.963639, 
    2.686715, 1.951471, 1.479334, 1.30299, 1.332211, 1.830276, 3.371325, 
    3.506874,
  0.6592776, 0.9780514, 1.491669, 1.846585, 2.275014, 2.844694, 4.754204, 
    6.004613, 4.780118, 3.94947, 2.83088, 2.326936, 1.857217, 1.5147, 
    1.335522, 1.029689, 0.6861313, 0.5327492, 0.6048309, 0.9025639, 1.25804, 
    1.064635, 1.39165, 1.472625, 1.12727, 0.7530946, 0.4837886, 0.3956007, 
    0.3924016,
  0.167223, 0.1398107, 0.1855573, 0.2918764, 0.530374, 0.412082, 0.4127182, 
    0.6967021, 0.6730381, 0.4729518, 0.6483406, 0.784937, 0.9278967, 
    0.8710663, 0.752479, 0.6778064, 0.4984009, 0.3331563, 0.2382358, 
    0.1749917, 0.3001347, 0.3934587, 0.327188, 0.3425045, 0.5575974, 
    0.611501, 0.5363719, 0.3118922, 0.1993485,
  0.06008036, 0.03799067, 0.04274623, 0.04491844, 0.04959013, 0.03415508, 
    0.02065266, 0.01885826, 0.0202345, 0.04136678, 0.08222251, 0.2074491, 
    0.2623973, 0.283684, 0.2125908, 0.1146723, 0.1385535, 0.1393283, 
    0.09681011, 0.05911538, 0.05436139, 0.05342007, 0.0450988, 0.04703258, 
    0.05236928, 0.1050935, 0.1558272, 0.118804, 0.06815951,
  0.008577872, 0.008696394, 0.01035874, 0.01160403, 0.01302914, 0.01556956, 
    0.01383192, 0.01141121, 0.008467484, 0.008646048, 0.01211354, 0.0158709, 
    0.02045903, 0.02091472, 0.01591659, 0.01631459, 0.01466413, 0.01975897, 
    0.02292654, 0.02412776, 0.01991523, 0.01323126, 0.008287389, 0.007531261, 
    0.00852535, 0.01421411, 0.01896299, 0.01586199, 0.01063155,
  0.003713142, 0.002890462, 0.002414769, 0.002746192, 0.002982337, 
    0.002738707, 0.002848033, 0.003708545, 0.003830021, 0.003742752, 
    0.003779331, 0.003665925, 0.003764326, 0.004655036, 0.002744286, 
    0.00326083, 0.004310778, 0.004996845, 0.005327482, 0.005334962, 
    0.004180672, 0.003669252, 0.003483322, 0.00350651, 0.00485186, 
    0.004686928, 0.005237476, 0.006793494, 0.004544796,
  0.002077556, 0.001924373, 0.00177717, 0.001821288, 0.001937577, 
    0.002022099, 0.002168531, 0.002373744, 0.002567008, 0.003019305, 
    0.003290998, 0.002541269, 0.002286702, 0.002164358, 0.001963887, 
    0.002049658, 0.002201538, 0.002687289, 0.003008634, 0.002721355, 
    0.002676012, 0.002626681, 0.002132691, 0.002100071, 0.002183682, 
    0.002078009, 0.002055599, 0.002184378, 0.002153618,
  0.02378623, 0.02378623, 0.02378623, 0.02378623, 0.02378623, 0.02378623, 
    0.02378623, 0.02248622, 0.02248622, 0.02248622, 0.02248622, 0.02248622, 
    0.02248622, 0.02248622, 0.02360819, 0.02360819, 0.02360819, 0.02360819, 
    0.02360819, 0.02360819, 0.02360819, 0.02429589, 0.02429589, 0.02429589, 
    0.02429589, 0.02429589, 0.02429589, 0.02429589, 0.02378623,
  0.01572161, 0.01846066, 0.02568419, 0.03727169, 0.04937186, 0.03202864, 
    0.01620893, 0.01164625, 0.008175819, 0.004712277, 0.003630576, 
    0.003107148, 0.003355299, 0.006372291, 0.006860975, 0.006966758, 
    0.009017285, 0.01047027, 0.01352584, 0.01701093, 0.01769068, 0.01637443, 
    0.01924837, 0.02857408, 0.02551061, 0.01750355, 0.01654911, 0.01277575, 
    0.01419874,
  0.009631373, 0.008225481, 0.01553595, 0.03905389, 0.08276391, 0.08638199, 
    0.02927756, 0.005387811, 0.003267739, 0.003605132, 0.00307708, 
    0.003090629, 0.005806617, 0.01330087, 0.01447527, 0.0126165, 0.008494006, 
    0.00785448, 0.009492096, 0.01612714, 0.02094805, 0.0206523, 0.03070557, 
    0.02984841, 0.02955965, 0.02364587, 0.01969714, 0.01513404, 0.01137303,
  0.0177479, 0.01377726, 0.01237998, 0.01440838, 0.0673053, 0.1228273, 
    0.08028598, 0.03401462, 0.01564403, 0.009836601, 0.007300888, 0.00983302, 
    0.01349813, 0.02396059, 0.04006049, 0.05097793, 0.04511179, 0.02856759, 
    0.02087873, 0.01722604, 0.01587492, 0.02103954, 0.02649267, 0.02819118, 
    0.03132889, 0.03185023, 0.03421237, 0.02942886, 0.02121694,
  0.1012825, 0.07642463, 0.06800265, 0.09379743, 0.208581, 0.3293254, 
    0.3304209, 0.2043764, 0.128828, 0.1129003, 0.09977791, 0.09278591, 
    0.1530582, 0.2262722, 0.2694336, 0.3095474, 0.2440772, 0.1589741, 
    0.1031761, 0.1054529, 0.1140317, 0.1219296, 0.1227951, 0.0972018, 
    0.0911473, 0.08236478, 0.09748004, 0.1054811, 0.1130531,
  0.4989969, 0.3781531, 0.4603524, 0.5235537, 0.6725523, 0.6950203, 
    0.6983954, 0.6732009, 0.4713218, 0.3531044, 0.421747, 0.5301843, 
    0.610038, 0.562533, 0.615266, 0.7227987, 0.6542822, 0.5785465, 0.463625, 
    0.4052138, 0.30961, 0.2738881, 0.2423281, 0.1537774, 0.1733363, 0.269712, 
    0.4512933, 0.5982531, 0.5179274,
  1.533243, 2.672988, 3.723637, 3.433683, 2.113576, 1.695486, 1.503828, 
    1.36824, 1.618081, 2.438886, 2.955269, 2.885385, 2.254055, 1.620203, 
    1.172161, 0.9251617, 0.8462204, 0.7655067, 0.688979, 0.4914785, 
    0.3977605, 0.4296249, 0.5153003, 0.7576484, 2.360507, 3.230268, 2.919505, 
    2.203346, 1.60947,
  5.336156, 9.260505, 8.658177, 6.341576, 4.094179, 2.868634, 2.360611, 
    2.754468, 3.712803, 4.774116, 5.724006, 5.179744, 3.428282, 2.148115, 
    1.60992, 1.244878, 1.102714, 0.8579158, 0.6845912, 0.6082274, 0.6805248, 
    1.163726, 3.472714, 6.115976, 9.513625, 8.609018, 5.41484, 3.189362, 
    3.489399,
  8.081616, 14.81478, 13.21977, 7.085117, 3.484542, 2.252929, 2.488093, 
    3.352131, 4.934481, 4.643604, 4.10121, 4.543813, 2.821834, 1.654095, 
    1.321529, 1.136075, 0.9586905, 0.8447081, 0.7358208, 0.7447418, 
    0.7862805, 1.00052, 3.855877, 10.23271, 13.19069, 10.43264, 5.626361, 
    3.443907, 4.626178,
  8.322108, 16.18679, 13.44826, 6.022214, 3.184865, 2.765484, 2.965147, 
    3.661134, 6.79506, 8.47854, 3.274839, 2.56921, 1.143724, 0.8263943, 
    0.8005521, 0.7956554, 0.7551027, 0.8485391, 0.8999918, 1.039585, 
    1.302008, 1.511676, 3.125675, 9.10823, 10.23872, 7.734805, 5.065566, 
    4.703009, 5.885873,
  10.35148, 12.69366, 10.93727, 5.860357, 4.430011, 4.109775, 5.034729, 
    5.75309, 6.347586, 4.55286, 2.614647, 1.532358, 1.128343, 1.051481, 
    0.9379345, 0.9361244, 0.9151313, 0.9939706, 1.254368, 1.776354, 2.389029, 
    3.188274, 4.75144, 6.604491, 5.519797, 5.23523, 5.866068, 7.61434, 
    9.235745,
  4.190732, 4.61109, 5.648344, 5.996581, 6.106482, 6.83733, 7.965495, 
    8.696718, 8.806052, 6.010448, 4.173466, 2.863774, 2.213538, 1.902338, 
    1.772803, 1.570408, 1.291751, 1.121404, 1.169649, 1.852099, 3.240458, 
    3.564635, 2.593773, 2.348749, 2.210313, 2.183422, 2.687317, 4.638992, 
    4.864491,
  1.076452, 1.279927, 1.717839, 2.157422, 2.561802, 3.16686, 5.162899, 
    6.881102, 5.618738, 5.171692, 4.007854, 3.345813, 2.670584, 2.315035, 
    2.224895, 1.826039, 1.48285, 1.07865, 1.010849, 1.18912, 1.828495, 
    1.687792, 2.296002, 2.491548, 2.124467, 1.544257, 1.065517, 0.8525522, 
    0.8005153,
  0.5254202, 0.3354739, 0.321643, 0.39356, 0.7056636, 0.5129247, 0.5487262, 
    0.9480191, 0.8699781, 0.7622593, 1.097478, 1.432629, 1.742808, 1.898174, 
    1.708739, 1.625185, 1.30206, 0.9400148, 0.6653054, 0.4060715, 0.5975175, 
    0.804741, 0.9864834, 1.187514, 1.449082, 1.656548, 1.478255, 0.9765734, 
    0.6794374,
  0.2422705, 0.1577878, 0.2222248, 0.1899294, 0.1619779, 0.1271575, 
    0.05926237, 0.04504457, 0.04694263, 0.1552765, 0.3087496, 0.578538, 
    0.7957853, 0.8074632, 0.6371761, 0.4629416, 0.529022, 0.5706558, 
    0.3938525, 0.1720611, 0.1578276, 0.18393, 0.1924082, 0.2181724, 
    0.2659203, 0.4404849, 0.6585839, 0.4901327, 0.2944351,
  0.05056626, 0.04014127, 0.05506442, 0.05461153, 0.05194101, 0.04626035, 
    0.03936825, 0.03456579, 0.03408171, 0.05135043, 0.1080065, 0.07982063, 
    0.09646797, 0.09978523, 0.06317928, 0.06303681, 0.06787404, 0.08722553, 
    0.09404025, 0.1196749, 0.09453379, 0.0538305, 0.04192337, 0.04443577, 
    0.03650933, 0.0634438, 0.1025185, 0.104756, 0.06785139,
  0.01225487, 0.008871062, 0.007831855, 0.009117144, 0.009588471, 
    0.008243918, 0.008181841, 0.009352261, 0.008874631, 0.008051984, 
    0.009041279, 0.01341733, 0.01383593, 0.01478428, 0.006648138, 
    0.006491906, 0.00898843, 0.01260727, 0.01487275, 0.0151861, 0.01241368, 
    0.01033022, 0.008915085, 0.009164851, 0.01579077, 0.01417883, 0.01376764, 
    0.02871484, 0.01667742,
  0.006503441, 0.006477897, 0.006323551, 0.006299415, 0.006224668, 
    0.006246238, 0.006842399, 0.007341362, 0.008361778, 0.009243646, 
    0.009954083, 0.009239286, 0.007716683, 0.007631659, 0.007172126, 
    0.006429908, 0.006810184, 0.008943305, 0.009853711, 0.009550753, 
    0.008605369, 0.007437153, 0.006009243, 0.005609288, 0.005853993, 
    0.005146109, 0.005244994, 0.006372903, 0.006684361,
  0.04555744, 0.04555744, 0.04555744, 0.04555744, 0.04555744, 0.04555744, 
    0.04555744, 0.04446058, 0.04446058, 0.04446058, 0.04446058, 0.04446058, 
    0.04446058, 0.04446058, 0.04609259, 0.04609259, 0.04609259, 0.04609259, 
    0.04609259, 0.04609259, 0.04609259, 0.04794558, 0.04794558, 0.04794558, 
    0.04794558, 0.04794558, 0.04794558, 0.04794558, 0.04555744,
  0.03094472, 0.03610782, 0.05205704, 0.08488295, 0.1083729, 0.07037695, 
    0.03684892, 0.02587368, 0.02365202, 0.01399559, 0.01110564, 0.01210109, 
    0.01194309, 0.01969417, 0.0205844, 0.02177264, 0.02576301, 0.02850999, 
    0.03392671, 0.03852307, 0.04005696, 0.04380615, 0.05496405, 0.0762903, 
    0.06639129, 0.04698271, 0.04421759, 0.03499455, 0.03002584,
  0.02954113, 0.0274784, 0.05907543, 0.1199466, 0.1785477, 0.16692, 
    0.09003432, 0.01928782, 0.01352755, 0.01619912, 0.01312373, 0.01315898, 
    0.0283165, 0.04748524, 0.04516223, 0.05095354, 0.04532963, 0.04059535, 
    0.04511859, 0.05910585, 0.07066429, 0.06395677, 0.08474261, 0.08527091, 
    0.08238234, 0.07324777, 0.06412138, 0.0473019, 0.0342582,
  0.0627725, 0.04882297, 0.0427447, 0.05722166, 0.1872542, 0.249779, 
    0.2008573, 0.1120567, 0.06247119, 0.04041342, 0.02852508, 0.04771358, 
    0.06677846, 0.117412, 0.1692005, 0.186962, 0.1674388, 0.1138889, 
    0.08337818, 0.0703532, 0.06353638, 0.07220553, 0.0768719, 0.08518208, 
    0.09633505, 0.09636412, 0.1218949, 0.1137149, 0.07975262,
  0.3292331, 0.2722768, 0.2276016, 0.2662132, 0.5618688, 0.7907209, 
    0.7519016, 0.5240793, 0.3312298, 0.2694941, 0.220061, 0.2308466, 
    0.3748479, 0.4903995, 0.6217477, 0.6638003, 0.5970895, 0.4011525, 
    0.2853615, 0.2508593, 0.2682921, 0.287902, 0.2907618, 0.2284474, 
    0.2280186, 0.2504769, 0.311747, 0.3957385, 0.4026782,
  1.028166, 0.7778538, 0.891271, 1.052227, 1.457936, 1.457848, 1.457833, 
    1.304227, 0.9501029, 0.70468, 0.6940974, 0.7741423, 0.9242674, 0.9742154, 
    1.095848, 1.222494, 1.104045, 0.9206594, 0.7323738, 0.6681643, 0.5547907, 
    0.504724, 0.4314117, 0.2841511, 0.3655515, 0.6560165, 1.160894, 1.386638, 
    1.109877,
  2.373431, 3.278898, 4.455742, 4.678293, 3.277252, 2.55882, 2.130595, 
    1.802747, 1.909532, 2.630241, 3.153512, 3.162243, 2.630585, 2.051481, 
    1.498473, 1.204869, 1.120514, 0.9699442, 0.8953649, 0.698342, 0.5786156, 
    0.72927, 0.7794836, 1.057943, 3.042102, 4.087119, 4.163722, 3.434296, 
    2.62995,
  6.302745, 10.65595, 10.45152, 7.40037, 4.944425, 3.31505, 2.586331, 
    2.852819, 3.784307, 4.801041, 5.855256, 5.471003, 3.68496, 2.325956, 
    1.739717, 1.349427, 1.191074, 0.8988984, 0.7701885, 0.7026622, 0.8519488, 
    1.611362, 3.973346, 7.047125, 10.48737, 9.626252, 6.552931, 4.347806, 
    4.592908,
  9.345423, 16.92636, 15.38395, 8.731359, 3.877697, 2.291401, 2.280972, 
    3.137527, 4.881021, 4.812071, 4.159129, 4.559219, 2.733031, 1.581962, 
    1.264556, 1.118183, 0.9413909, 0.8542234, 0.7589741, 0.7566527, 
    0.8639923, 1.330747, 4.944619, 12.34511, 15.04769, 11.78051, 6.336263, 
    4.403825, 5.572846,
  9.999452, 18.30005, 15.94012, 7.020208, 3.581412, 2.797848, 2.766165, 
    3.333601, 6.983264, 9.062756, 3.302422, 2.385707, 1.083473, 0.7900578, 
    0.7373539, 0.7887824, 0.7413799, 0.8241659, 0.8827002, 1.075024, 
    1.454718, 1.828874, 4.441229, 12.34989, 12.45896, 9.076691, 5.790476, 
    5.759983, 7.227684,
  12.33871, 14.59318, 13.51447, 6.756875, 4.728765, 3.996447, 4.874787, 
    5.42694, 6.336727, 4.539265, 2.652452, 1.504037, 1.122916, 1.04417, 
    0.9521249, 0.9479728, 0.9429407, 1.010302, 1.28837, 1.848973, 2.573416, 
    3.459275, 5.424645, 8.074549, 6.982996, 6.259938, 6.859801, 8.630982, 
    11.18721,
  5.301262, 5.860077, 6.89149, 6.971783, 6.939583, 7.370231, 8.222403, 
    8.803583, 9.31878, 6.366497, 4.441611, 3.099662, 2.416208, 2.14098, 
    1.987504, 1.817068, 1.534534, 1.288529, 1.258211, 1.961854, 3.419701, 
    4.105474, 3.149621, 3.160707, 3.323738, 3.031832, 3.515826, 5.374875, 
    5.907415,
  1.610674, 1.797061, 2.085256, 2.604247, 2.922501, 3.47488, 5.509704, 
    7.496518, 6.423091, 6.223915, 5.184737, 4.392651, 3.584082, 3.088464, 
    3.016826, 2.59422, 2.231053, 1.677136, 1.433925, 1.487413, 2.516436, 
    2.307825, 3.177131, 3.411445, 3.015571, 2.382334, 1.780206, 1.426762, 
    1.401948,
  1.134474, 0.8347921, 0.6879012, 0.6515912, 1.132143, 0.7652896, 0.7318344, 
    1.398715, 1.334931, 1.441027, 2.049853, 2.413262, 2.846415, 3.121881, 
    2.939613, 2.675183, 2.304695, 1.78731, 1.41446, 0.8251536, 1.081359, 
    1.567769, 2.03031, 2.48137, 2.568921, 2.851479, 2.55216, 2.008177, 
    1.507634,
  0.729188, 0.6396763, 0.833451, 0.7732114, 0.6105391, 0.602592, 0.3354817, 
    0.1626817, 0.2419403, 0.7161781, 1.040745, 1.226475, 1.695535, 1.774312, 
    1.450945, 1.355631, 1.320355, 1.446624, 1.101978, 0.5632568, 0.4939238, 
    0.6239192, 0.6411173, 0.630644, 0.8808182, 1.210715, 1.57109, 1.222008, 
    0.8248468,
  0.2591394, 0.2152491, 0.2935246, 0.3216006, 0.3240156, 0.2592958, 
    0.2230523, 0.2388618, 0.2514711, 0.4249246, 0.6350212, 0.5007392, 
    0.4372053, 0.4546375, 0.3332351, 0.2594431, 0.2824567, 0.2858955, 
    0.3023347, 0.3887213, 0.3658154, 0.2752452, 0.2558405, 0.1970701, 
    0.1902553, 0.310343, 0.4708874, 0.4359156, 0.3126238,
  0.0629584, 0.04120319, 0.03117292, 0.03536539, 0.03725029, 0.03593183, 
    0.03816131, 0.04086873, 0.04136927, 0.04098788, 0.0576185, 0.08037248, 
    0.06209521, 0.06497031, 0.047348, 0.03193791, 0.04562432, 0.0692668, 
    0.07578787, 0.06714552, 0.05350802, 0.04946528, 0.04890873, 0.04313217, 
    0.09204087, 0.0514053, 0.04218412, 0.1346716, 0.08581898,
  0.03912995, 0.03491928, 0.03369682, 0.03202901, 0.03129553, 0.03184469, 
    0.0319407, 0.03282658, 0.03714433, 0.04015282, 0.04063616, 0.03882308, 
    0.03826471, 0.03553414, 0.03186368, 0.03139094, 0.0310558, 0.03447655, 
    0.03682555, 0.03668411, 0.03661322, 0.03443006, 0.02282895, 0.02064569, 
    0.02401036, 0.01837945, 0.02089464, 0.0348964, 0.04347958,
  0.07273281, 0.07273281, 0.07273281, 0.07273281, 0.07273281, 0.07273281, 
    0.07273281, 0.07000896, 0.07000896, 0.07000896, 0.07000896, 0.07000896, 
    0.07000896, 0.07000896, 0.07198328, 0.07198328, 0.07198328, 0.07198328, 
    0.07198328, 0.07198328, 0.07198328, 0.07622317, 0.07622317, 0.07622317, 
    0.07622317, 0.07622317, 0.07622317, 0.07622317, 0.07273281,
  0.05700063, 0.06288863, 0.08804005, 0.1413724, 0.1600323, 0.1190327, 
    0.07115284, 0.05194412, 0.04762325, 0.03471054, 0.02758169, 0.03183723, 
    0.03046376, 0.04978515, 0.05798578, 0.06492599, 0.07466191, 0.07388484, 
    0.07888316, 0.08008494, 0.08337637, 0.09080394, 0.1113405, 0.1515559, 
    0.1325153, 0.1004922, 0.09565628, 0.07585407, 0.05914243,
  0.07538559, 0.07454929, 0.1230493, 0.2401048, 0.2700653, 0.2597725, 
    0.1963215, 0.05742295, 0.0434725, 0.05719363, 0.04808625, 0.0458759, 
    0.09326902, 0.1295405, 0.1226821, 0.1466633, 0.1431325, 0.1246396, 
    0.1288776, 0.151706, 0.1666117, 0.1534686, 0.1722691, 0.1830313, 
    0.1673732, 0.1609091, 0.1442465, 0.1100725, 0.08919953,
  0.1709854, 0.1358235, 0.1246443, 0.2100069, 0.3896055, 0.4425068, 
    0.3887753, 0.2506731, 0.1720158, 0.1313853, 0.104661, 0.1608258, 
    0.2216279, 0.3906322, 0.4691254, 0.4875091, 0.4619356, 0.3576866, 
    0.2697789, 0.2433982, 0.2051593, 0.2048993, 0.1903354, 0.2110266, 
    0.2314478, 0.2487449, 0.2946291, 0.2620494, 0.21348,
  0.7158622, 0.6179997, 0.5421469, 0.6737664, 1.107035, 1.379813, 1.324187, 
    1.036276, 0.6854493, 0.5390736, 0.4432205, 0.5178401, 0.7049156, 
    0.9679254, 1.175779, 1.22722, 1.132937, 0.8079581, 0.6388425, 0.5036159, 
    0.4982804, 0.5145875, 0.4994542, 0.4058348, 0.4511175, 0.5480673, 
    0.747541, 0.8978593, 0.858826,
  1.71758, 1.378666, 1.427609, 1.879837, 2.454535, 2.380054, 2.307089, 
    1.976699, 1.558679, 1.213468, 1.150984, 1.19295, 1.446602, 1.590848, 
    1.707586, 1.781474, 1.556938, 1.288128, 1.029422, 0.9259883, 0.7921892, 
    0.7371221, 0.650518, 0.4982241, 0.7128704, 1.370919, 2.095286, 2.268448, 
    1.867718,
  3.207677, 3.749772, 5.021703, 5.833949, 4.521698, 3.372029, 2.744327, 
    2.287266, 2.162419, 2.740317, 3.206229, 3.395351, 2.928133, 2.514421, 
    1.901654, 1.515435, 1.378646, 1.153942, 1.015659, 0.8270762, 0.7008859, 
    0.94028, 0.9396781, 1.406859, 3.599358, 4.839165, 5.190342, 4.535502, 
    3.620785,
  6.744846, 11.17727, 11.71315, 8.21605, 5.680595, 3.761711, 2.730994, 
    2.806987, 3.635975, 4.702363, 5.851826, 5.627277, 3.832545, 2.447416, 
    1.85942, 1.442014, 1.219046, 0.9127898, 0.8212261, 0.7345885, 0.927729, 
    1.862804, 4.191681, 7.570435, 11.14635, 10.31414, 7.397843, 5.304058, 
    5.394865,
  10.05939, 17.68078, 16.77988, 9.879729, 4.357988, 2.38004, 2.10387, 
    2.923395, 4.660261, 4.853512, 4.165521, 4.441926, 2.667393, 1.514018, 
    1.199096, 1.054353, 0.9283792, 0.8388402, 0.7640265, 0.7877722, 
    0.9409674, 1.596852, 5.691404, 13.91818, 16.1801, 12.85322, 6.932506, 
    5.138738, 6.325437,
  10.99937, 19.79076, 18.00903, 7.792528, 3.996528, 2.857924, 2.622556, 
    3.118006, 7.041026, 9.454695, 3.326179, 2.196993, 1.038742, 0.7632268, 
    0.679822, 0.7552742, 0.7059065, 0.7830338, 0.8676759, 1.078904, 1.514537, 
    2.058817, 5.66298, 14.5874, 13.9341, 9.847619, 6.43903, 6.433288, 8.431609,
  13.33653, 15.68698, 14.91837, 7.533681, 4.94753, 3.991658, 4.761621, 
    5.151858, 6.210688, 4.409513, 2.681745, 1.481022, 1.097971, 1.036192, 
    0.9496254, 0.9660432, 0.9605727, 0.9973329, 1.276945, 1.82983, 2.602734, 
    3.551875, 5.954921, 9.460382, 8.068511, 6.870887, 7.31643, 8.910159, 
    12.21965,
  6.037723, 6.467799, 7.366572, 7.467526, 7.358656, 7.571571, 8.312318, 
    8.698137, 9.526542, 6.556549, 4.658712, 3.367129, 2.643459, 2.379589, 
    2.196507, 1.994729, 1.724975, 1.393142, 1.295639, 1.998359, 3.512881, 
    4.491318, 3.602554, 3.732087, 4.18461, 3.679575, 4.018643, 5.652649, 
    6.455042,
  2.091116, 2.476462, 2.596678, 2.939702, 3.239917, 3.785033, 5.813036, 
    8.000048, 7.240567, 7.254704, 6.26973, 5.303094, 4.375764, 3.715172, 
    3.561, 3.175904, 2.716731, 2.215393, 1.790462, 1.734051, 3.12379, 
    2.934535, 3.982716, 4.053238, 3.586284, 2.960888, 2.376182, 1.93788, 
    1.948186,
  1.831822, 1.564468, 1.518186, 1.201707, 2.164814, 1.457342, 1.109261, 
    2.292553, 2.454733, 2.755185, 3.493223, 3.774909, 4.085544, 4.257608, 
    3.996623, 3.590781, 3.077248, 2.565626, 2.204752, 1.40901, 1.660909, 
    2.494611, 3.138125, 3.673355, 3.62796, 3.7407, 3.425969, 2.958799, 
    2.350595,
  1.452407, 1.641653, 2.050856, 2.183435, 1.856224, 1.693319, 1.289458, 
    0.6819431, 1.085305, 2.088995, 2.655077, 2.343314, 2.813909, 2.969534, 
    2.586219, 2.582095, 2.299423, 2.361483, 1.939521, 1.242439, 1.290029, 
    1.47307, 1.467643, 1.338074, 1.733321, 2.168827, 2.479616, 2.176444, 
    1.588284,
  0.7403414, 0.7697095, 0.9675754, 1.144659, 1.23992, 1.086586, 1.073689, 
    0.9234868, 0.8927811, 1.347942, 1.670959, 1.321936, 1.145583, 1.302881, 
    1.089839, 0.7660602, 0.7168406, 0.7284735, 0.722438, 0.9539598, 
    0.8766758, 0.8229674, 0.7854131, 0.6231073, 0.6578316, 0.9607744, 
    1.137264, 0.9901984, 0.8076268,
  0.252549, 0.1803708, 0.134534, 0.1670209, 0.1866458, 0.213457, 0.2310311, 
    0.2606914, 0.2666008, 0.2807243, 0.3411976, 0.3851739, 0.3105897, 
    0.3113015, 0.2736954, 0.183591, 0.2296026, 0.2827711, 0.3210758, 
    0.2952046, 0.2385409, 0.2528138, 0.2831237, 0.2382616, 0.407133, 
    0.1878962, 0.1340153, 0.4494974, 0.3334415,
  0.1908056, 0.1665236, 0.1419291, 0.1397711, 0.1596185, 0.1710603, 
    0.1556668, 0.1703101, 0.1971865, 0.2313331, 0.2145243, 0.1973078, 
    0.2137522, 0.1933465, 0.184397, 0.1824191, 0.1686263, 0.1532177, 
    0.144105, 0.1605728, 0.1733414, 0.1714615, 0.1228257, 0.1114148, 
    0.1189717, 0.08060557, 0.09800513, 0.176028, 0.2039069,
  0.1068113, 0.1068113, 0.1068113, 0.1068113, 0.1068113, 0.1068113, 
    0.1068113, 0.1014925, 0.1014925, 0.1014925, 0.1014925, 0.1014925, 
    0.1014925, 0.1014925, 0.1031661, 0.1031661, 0.1031661, 0.1031661, 
    0.1031661, 0.1031661, 0.1031661, 0.1100907, 0.1100907, 0.1100907, 
    0.1100907, 0.1100907, 0.1100907, 0.1100907, 0.1068113,
  0.1022332, 0.1058445, 0.1387274, 0.2073901, 0.2138944, 0.1745247, 
    0.1210056, 0.09798064, 0.08198255, 0.07128331, 0.06024703, 0.06720344, 
    0.0651826, 0.1042177, 0.1277508, 0.1467344, 0.1612504, 0.1592553, 
    0.1538417, 0.1486744, 0.154485, 0.157188, 0.1868091, 0.2541313, 
    0.2318824, 0.1919426, 0.1853454, 0.1488381, 0.1106547,
  0.1738568, 0.1705094, 0.2334471, 0.3837151, 0.3651278, 0.3641971, 
    0.3345099, 0.1309415, 0.104449, 0.1369304, 0.1223318, 0.1287092, 
    0.2135667, 0.286727, 0.2735381, 0.302498, 0.304809, 0.2596368, 0.2639901, 
    0.2866053, 0.2986939, 0.2777593, 0.2890924, 0.3066329, 0.2830639, 
    0.2976521, 0.2684203, 0.2249648, 0.2083347,
  0.341518, 0.2731383, 0.2620528, 0.4617989, 0.6487655, 0.6807005, 0.629081, 
    0.4592383, 0.34204, 0.2896477, 0.2525876, 0.371455, 0.5205388, 0.8146623, 
    0.9442192, 0.9595149, 0.8769327, 0.7280852, 0.564875, 0.5209664, 
    0.4262654, 0.406976, 0.3573947, 0.3803408, 0.4136485, 0.4647752, 
    0.5042187, 0.4702983, 0.3925424,
  1.128464, 1.051597, 0.9096623, 1.227628, 1.698492, 1.984503, 1.829759, 
    1.518037, 1.08224, 0.8559458, 0.7665105, 0.9201182, 1.166421, 1.587084, 
    1.846503, 1.843836, 1.639852, 1.240335, 1.047604, 0.8678947, 0.8014295, 
    0.7668105, 0.7158177, 0.5897128, 0.6868619, 0.9405602, 1.175393, 
    1.379168, 1.372094,
  2.336983, 2.013739, 1.99539, 2.722582, 3.246842, 3.145472, 3.002597, 
    2.536534, 2.090201, 1.761006, 1.651561, 1.74069, 2.054202, 2.284681, 
    2.293776, 2.262559, 1.924887, 1.5975, 1.2865, 1.143669, 0.9662633, 
    0.8924066, 0.8299186, 0.7342409, 1.22949, 2.081258, 2.945801, 2.945081, 
    2.485259,
  3.839282, 4.041112, 5.525414, 6.630647, 5.347289, 4.014535, 3.289486, 
    2.805657, 2.398025, 2.760401, 3.277547, 3.693536, 3.277499, 2.899015, 
    2.257337, 1.78843, 1.550627, 1.276155, 1.082556, 0.8941371, 0.7614163, 
    1.021037, 0.9814064, 1.592214, 3.787827, 5.392747, 5.919939, 5.228283, 
    4.360467,
  6.918411, 11.01666, 12.19916, 8.620864, 6.252575, 4.194493, 2.844071, 
    2.701006, 3.416399, 4.539516, 5.814036, 5.714417, 3.922593, 2.543113, 
    1.988263, 1.502481, 1.209719, 0.913018, 0.8309574, 0.7335629, 0.9445924, 
    1.915414, 4.111956, 7.501689, 11.38712, 10.69244, 7.884523, 5.820926, 
    5.779555,
  10.08707, 17.54919, 17.41317, 10.42521, 4.933578, 2.527627, 2.023263, 
    2.735171, 4.40026, 4.747063, 4.130227, 4.279584, 2.623518, 1.459404, 
    1.148679, 0.991374, 0.9235993, 0.8053027, 0.757548, 0.7928965, 0.9826122, 
    1.793522, 6.121356, 14.74715, 16.86804, 13.44593, 7.406814, 5.641001, 
    6.786213,
  11.43638, 20.97889, 19.40871, 8.398413, 4.366763, 2.99489, 2.562547, 
    2.959858, 7.038629, 9.648513, 3.337336, 2.006117, 0.9970132, 0.7319649, 
    0.6402501, 0.694745, 0.6803166, 0.7474356, 0.8682464, 1.056639, 1.564145, 
    2.23005, 6.733963, 16.04635, 14.70421, 10.02992, 6.834335, 6.979609, 
    9.179541,
  13.65406, 16.05454, 15.66717, 8.279982, 5.12184, 3.985006, 4.704709, 
    4.954487, 5.991002, 4.24919, 2.675088, 1.452036, 1.061363, 1.03363, 
    0.939459, 0.9836705, 0.9814708, 0.9726458, 1.262007, 1.797316, 2.57017, 
    3.594332, 6.360296, 10.47333, 8.488967, 7.142161, 7.386165, 8.885127, 
    12.77757,
  6.336086, 6.490202, 7.218618, 7.497521, 7.452131, 7.558548, 8.258081, 
    8.531659, 9.648398, 6.611326, 4.771348, 3.624554, 2.87049, 2.570473, 
    2.383253, 2.095285, 1.831793, 1.444646, 1.33018, 2.013833, 3.520652, 
    4.747013, 3.922358, 4.098278, 4.506234, 3.946114, 4.135959, 5.654241, 
    6.535527,
  2.506706, 3.087049, 2.95845, 3.15206, 3.433624, 4.091163, 6.120589, 
    8.407858, 7.958648, 8.309496, 7.211516, 6.071563, 4.992352, 4.128158, 
    3.973517, 3.588529, 3.015609, 2.52688, 1.961189, 1.8958, 3.542405, 
    3.525978, 4.579181, 4.490899, 3.834306, 3.247887, 2.776593, 2.392066, 
    2.340556,
  2.505993, 2.478755, 2.769123, 2.179616, 3.648462, 2.790019, 1.879434, 
    3.604652, 4.196138, 4.496829, 5.166287, 5.088264, 5.256067, 5.206897, 
    4.86115, 4.286002, 3.573403, 3.171567, 2.802577, 1.986907, 2.266005, 
    3.397951, 4.244926, 4.692655, 4.460861, 4.33941, 4.054276, 3.625349, 
    3.007354,
  2.210361, 2.832316, 3.484311, 3.98734, 3.6013, 3.327677, 2.794425, 
    1.915396, 2.78435, 3.897274, 4.61008, 3.769258, 3.869699, 4.098748, 
    3.811486, 3.728238, 3.206965, 3.101177, 2.697323, 2.098818, 2.373556, 
    2.592428, 2.543175, 2.274588, 2.775092, 3.05056, 3.268964, 3.00599, 
    2.339759,
  1.4963, 1.62222, 1.968886, 2.392059, 2.596419, 2.533669, 2.551888, 
    2.135465, 2.007539, 2.761353, 3.154204, 2.453176, 2.280803, 2.50038, 
    2.216223, 1.590001, 1.444223, 1.455403, 1.347092, 1.720574, 1.717491, 
    1.555899, 1.621461, 1.346004, 1.529441, 1.894602, 1.93911, 1.621011, 
    1.498436,
  0.66492, 0.5267208, 0.4817217, 0.6541904, 0.6718564, 0.7493054, 0.8315716, 
    0.9306201, 0.876784, 0.9890704, 1.049797, 1.106794, 0.9771085, 1.003813, 
    0.8444962, 0.6904752, 0.7188398, 0.8045976, 0.8471062, 0.8398615, 
    0.7668059, 0.8174404, 0.8647083, 0.7626073, 1.038757, 0.5052856, 
    0.352527, 1.006448, 0.8237021,
  0.5250781, 0.4675131, 0.412277, 0.4514874, 0.5278492, 0.5701602, 0.582653, 
    0.6144216, 0.6663293, 0.7039201, 0.7016042, 0.7279723, 0.7753264, 
    0.7224199, 0.6721113, 0.6479008, 0.5717112, 0.4913971, 0.4678997, 
    0.492216, 0.5036464, 0.4934816, 0.3913764, 0.3828894, 0.3985298, 
    0.2727024, 0.3359005, 0.5261259, 0.5570222,
  0.154615, 0.154615, 0.154615, 0.154615, 0.154615, 0.154615, 0.154615, 
    0.1477723, 0.1477723, 0.1477723, 0.1477723, 0.1477723, 0.1477723, 
    0.1477723, 0.1481623, 0.1481623, 0.1481623, 0.1481623, 0.1481623, 
    0.1481623, 0.1481623, 0.1583794, 0.1583794, 0.1583794, 0.1583794, 
    0.1583794, 0.1583794, 0.1583794, 0.154615,
  0.1742871, 0.1678025, 0.2089578, 0.2734692, 0.2732025, 0.2338718, 
    0.1768876, 0.1512891, 0.1323769, 0.1204375, 0.1098086, 0.1213329, 
    0.1179484, 0.1792819, 0.2258375, 0.255994, 0.2699226, 0.2714984, 
    0.2627076, 0.2543684, 0.2506096, 0.243292, 0.2842405, 0.3666746, 
    0.3464019, 0.306456, 0.3030854, 0.2486174, 0.1852171,
  0.3243506, 0.3255761, 0.3975123, 0.5366889, 0.4693053, 0.4695436, 
    0.4750679, 0.2384559, 0.2011997, 0.2374311, 0.2455124, 0.2666091, 
    0.3761093, 0.4947651, 0.4857991, 0.4964443, 0.5160249, 0.4329206, 
    0.4233032, 0.4214761, 0.4265735, 0.4050249, 0.4169079, 0.4201828, 
    0.4240932, 0.4425826, 0.4384838, 0.3941096, 0.3736419,
  0.5478649, 0.4490802, 0.4461831, 0.6957963, 0.9132707, 0.9290904, 
    0.8685752, 0.6890249, 0.5411971, 0.4770938, 0.4503921, 0.6208469, 
    0.8711951, 1.188959, 1.396188, 1.373467, 1.232143, 1.07451, 0.8838341, 
    0.8033615, 0.6489362, 0.5979468, 0.5302098, 0.5407746, 0.5849349, 
    0.6502573, 0.7089138, 0.6538458, 0.6003483,
  1.434699, 1.398692, 1.235216, 1.5761, 2.086692, 2.349603, 2.193569, 
    1.875944, 1.401692, 1.105876, 1.051669, 1.250447, 1.65072, 2.093891, 
    2.49123, 2.334038, 2.052301, 1.604588, 1.362967, 1.180901, 1.067914, 
    0.974659, 0.9078275, 0.7639261, 0.882553, 1.271585, 1.472323, 1.71569, 
    1.718755,
  2.739578, 2.484158, 2.450328, 3.372961, 3.732768, 3.580231, 3.364446, 
    2.904315, 2.488872, 2.22919, 2.085852, 2.176589, 2.660148, 2.834796, 
    2.763829, 2.585746, 2.188931, 1.789976, 1.414932, 1.271402, 1.085281, 
    0.9837252, 0.9373607, 0.8915317, 1.784707, 2.622468, 3.317968, 3.275266, 
    2.828148,
  4.19157, 4.207529, 5.967222, 7.000205, 5.705392, 4.508296, 3.722047, 
    3.233927, 2.657192, 2.762844, 3.391101, 4.090607, 3.674133, 3.227955, 
    2.522638, 1.998476, 1.653733, 1.364539, 1.108964, 0.9038122, 0.7783287, 
    1.011327, 0.9754952, 1.513651, 3.82863, 5.664322, 6.165757, 5.446731, 
    4.685719,
  6.932293, 10.58447, 11.9852, 8.583066, 6.599717, 4.568063, 2.988062, 
    2.656246, 3.196698, 4.304435, 5.715083, 5.68258, 3.976259, 2.628641, 
    2.120415, 1.541117, 1.198611, 0.9096299, 0.8136705, 0.7098944, 0.9468198, 
    1.817955, 3.831883, 6.982414, 11.24631, 10.71464, 8.097399, 5.979345, 
    5.901431,
  9.875412, 16.71851, 17.57137, 10.45482, 5.265027, 2.712212, 2.007998, 
    2.58189, 4.110824, 4.541153, 4.024488, 4.093591, 2.574248, 1.417818, 
    1.102941, 0.9566794, 0.8983733, 0.7785121, 0.7411936, 0.7958436, 
    1.023894, 1.887064, 6.190258, 15.27975, 17.24312, 13.63008, 7.63643, 
    6.110436, 7.001098,
  11.26018, 21.73786, 19.87904, 8.544997, 4.685247, 3.146587, 2.539743, 
    2.791389, 6.943689, 9.686237, 3.243011, 1.826269, 0.9652281, 0.7034776, 
    0.6080732, 0.6345156, 0.6556212, 0.7152479, 0.8578039, 1.030317, 
    1.588223, 2.362823, 7.58441, 16.71283, 14.81741, 9.674829, 6.922724, 
    7.25852, 9.366803,
  13.74926, 15.89623, 15.80313, 9.002816, 5.278315, 3.975978, 4.680007, 
    4.789451, 5.729145, 4.05688, 2.626303, 1.425157, 1.041352, 1.031428, 
    0.9279984, 1.001255, 0.9939908, 0.9729244, 1.250245, 1.772406, 2.494147, 
    3.623764, 6.590894, 10.9417, 8.328977, 7.071609, 7.295954, 8.821176, 
    13.11392,
  6.286935, 6.272121, 6.732897, 7.053679, 7.314673, 7.555923, 8.161839, 
    8.38481, 9.680593, 6.577239, 4.83347, 3.808589, 3.02715, 2.69268, 
    2.489353, 2.155774, 1.866806, 1.473351, 1.352681, 2.007749, 3.447732, 
    4.884505, 4.016949, 4.274965, 4.414926, 3.811216, 4.008547, 5.408183, 
    6.273714,
  2.933845, 3.469703, 3.299579, 3.37215, 3.600792, 4.422485, 6.407755, 
    8.732576, 8.5679, 9.412405, 8.042457, 6.688204, 5.399309, 4.455381, 
    4.301945, 3.826991, 3.223818, 2.690687, 2.011859, 2.015742, 3.862778, 
    3.987476, 5.00702, 4.758083, 3.915428, 3.390134, 3.066097, 2.820334, 
    2.662182,
  3.165564, 3.390724, 4.053868, 3.599983, 5.332552, 4.527231, 3.192306, 
    5.210073, 6.247157, 6.417486, 6.900018, 6.388941, 6.319797, 6.045963, 
    5.568404, 4.825684, 3.936874, 3.548035, 3.192374, 2.441309, 2.761375, 
    4.150885, 5.188708, 5.447414, 5.092621, 4.752271, 4.475924, 4.041746, 
    3.488166,
  2.901605, 3.825615, 4.585734, 5.569538, 5.057281, 5.013116, 4.642222, 
    3.675114, 4.79943, 5.734765, 6.281106, 5.069069, 4.843159, 5.076283, 
    4.887522, 4.672262, 3.991356, 3.685236, 3.302767, 2.920146, 3.324559, 
    3.672634, 3.662381, 3.353564, 3.750139, 3.850677, 3.889644, 3.656024, 
    2.97329,
  2.28936, 2.409006, 2.959422, 3.54306, 3.932473, 3.971769, 4.027484, 
    3.515363, 3.307527, 4.158657, 4.640257, 3.680084, 3.618876, 3.751723, 
    3.459205, 2.639117, 2.3216, 2.27104, 2.030497, 2.519874, 2.652571, 
    2.471137, 2.632122, 2.2206, 2.55566, 2.723157, 2.683642, 2.292794, 
    2.238285,
  1.246035, 1.102222, 1.143862, 1.465208, 1.497017, 1.492151, 1.686502, 
    1.829253, 1.72822, 1.89534, 1.986314, 2.059071, 1.92586, 1.910149, 
    1.706768, 1.527928, 1.455989, 1.528955, 1.573084, 1.619979, 1.606581, 
    1.613251, 1.712147, 1.562044, 1.804085, 1.023445, 0.7467336, 1.710615, 
    1.479899,
  1.013867, 0.9348862, 0.9131973, 1.003257, 1.111285, 1.163298, 1.244941, 
    1.27699, 1.311814, 1.355227, 1.467574, 1.61017, 1.664966, 1.584695, 
    1.488556, 1.418224, 1.273188, 1.107164, 1.06492, 1.059861, 1.034989, 
    1.032414, 0.8764474, 0.8712973, 0.9088527, 0.670477, 0.789603, 1.083387, 
    1.085181,
  0.2110141, 0.2110141, 0.2110141, 0.2110141, 0.2110141, 0.2110141, 
    0.2110141, 0.2043426, 0.2043426, 0.2043426, 0.2043426, 0.2043426, 
    0.2043426, 0.2043426, 0.2055644, 0.2055644, 0.2055644, 0.2055644, 
    0.2055644, 0.2055644, 0.2055644, 0.2175779, 0.2175779, 0.2175779, 
    0.2175779, 0.2175779, 0.2175779, 0.2175779, 0.2110141,
  0.2683745, 0.242781, 0.2864949, 0.3350827, 0.3265613, 0.2891599, 0.2324896, 
    0.2047199, 0.1890366, 0.1742077, 0.1715359, 0.1885182, 0.1827526, 
    0.2616042, 0.3286465, 0.3599334, 0.3703977, 0.3838101, 0.3851869, 
    0.3726239, 0.3541279, 0.3379373, 0.3812001, 0.45352, 0.4416122, 
    0.4103646, 0.4080175, 0.3519283, 0.2833117,
  0.492127, 0.4987567, 0.5683957, 0.6839169, 0.5803102, 0.564316, 0.5933071, 
    0.3694834, 0.3167886, 0.3434686, 0.3884604, 0.41692, 0.5486077, 
    0.6879178, 0.6899458, 0.6883087, 0.7120931, 0.5986133, 0.5771461, 
    0.5494605, 0.5451776, 0.5229305, 0.5240721, 0.518496, 0.5653507, 
    0.5562897, 0.5811805, 0.5475161, 0.5258532,
  0.7269034, 0.6359779, 0.6403899, 0.8774329, 1.123888, 1.111961, 1.056681, 
    0.8749753, 0.7179685, 0.643792, 0.662675, 0.8461053, 1.119677, 1.48834, 
    1.710395, 1.670531, 1.495281, 1.350879, 1.125969, 1.010375, 0.8173853, 
    0.7432042, 0.6705969, 0.6711411, 0.7132369, 0.7913844, 0.8774765, 
    0.8180991, 0.8059417,
  1.634064, 1.59357, 1.447076, 1.773739, 2.324624, 2.526602, 2.348498, 
    2.056958, 1.571456, 1.25406, 1.229816, 1.452582, 1.951365, 2.497645, 
    2.930729, 2.641731, 2.365042, 1.860002, 1.576427, 1.402632, 1.255827, 
    1.124933, 1.041283, 0.8978513, 1.000905, 1.487313, 1.674416, 1.928423, 
    1.910532,
  2.983708, 2.769214, 2.727325, 3.693732, 3.891893, 3.72839, 3.495236, 
    3.08947, 2.693676, 2.505916, 2.331745, 2.435038, 3.106426, 3.220158, 
    3.126294, 2.815919, 2.37144, 1.909298, 1.492682, 1.346155, 1.158134, 
    1.028929, 0.9748776, 0.9921157, 2.221389, 2.927676, 3.36683, 3.330758, 
    2.973662,
  4.260259, 4.195508, 6.300781, 7.135911, 5.865664, 4.755796, 3.976907, 
    3.443685, 2.900587, 2.826491, 3.496582, 4.357912, 4.012916, 3.536194, 
    2.807427, 2.167154, 1.754711, 1.436542, 1.115371, 0.889335, 0.8026816, 
    0.9736226, 0.9647208, 1.290693, 3.915188, 5.680637, 6.174358, 5.378833, 
    4.683284,
  6.69824, 9.996332, 11.58561, 8.36039, 6.638813, 4.828235, 3.183274, 
    2.674097, 2.996734, 4.010588, 5.498071, 5.577727, 3.95584, 2.684724, 
    2.211527, 1.579184, 1.199174, 0.9071665, 0.7839312, 0.6862152, 0.9693566, 
    1.681453, 3.447269, 6.374674, 10.8462, 10.47645, 8.03381, 5.884724, 
    5.826023,
  9.488095, 15.48684, 17.35037, 9.980574, 5.342345, 2.967242, 2.045378, 
    2.465748, 3.792217, 4.265913, 3.795402, 3.88477, 2.547549, 1.397111, 
    1.072231, 0.9359739, 0.8632011, 0.748916, 0.713444, 0.7817748, 1.015472, 
    1.778125, 6.053404, 15.2585, 17.35014, 13.2802, 7.62434, 6.274471, 
    6.942811,
  10.83329, 21.59897, 19.16252, 8.365811, 4.849988, 3.260885, 2.52438, 
    2.621359, 6.725609, 9.471968, 3.133415, 1.654209, 0.9375327, 0.6743713, 
    0.5918034, 0.590877, 0.6318554, 0.6842827, 0.8210911, 1.024818, 1.610789, 
    2.520952, 7.703404, 16.63736, 14.31813, 9.075025, 6.785609, 7.055115, 
    9.087246,
  13.66756, 15.21141, 15.31952, 9.627211, 5.289084, 4.008492, 4.657145, 
    4.673989, 5.449531, 3.834886, 2.558969, 1.382428, 1.048629, 1.031158, 
    0.9269369, 1.006366, 0.9852024, 0.9807126, 1.23533, 1.734555, 2.427525, 
    3.556618, 6.597788, 10.72456, 7.771708, 6.83171, 7.091191, 8.631023, 
    13.18096,
  5.997379, 5.971634, 6.157435, 6.496817, 6.968182, 7.385827, 8.07165, 
    8.243061, 9.620605, 6.580389, 4.855916, 3.899654, 3.106637, 2.779272, 
    2.49825, 2.186474, 1.862606, 1.495775, 1.337072, 1.984172, 3.330257, 
    4.974045, 3.936425, 4.169765, 4.102201, 3.525468, 3.769714, 4.868487, 
    5.910227,
  3.337721, 3.825552, 3.72303, 3.600366, 3.761748, 4.705667, 6.686347, 
    8.982853, 9.169842, 10.35129, 8.82423, 7.048103, 5.64215, 4.707876, 
    4.548424, 3.941797, 3.358368, 2.774025, 2.025418, 2.11339, 4.069694, 
    4.261791, 5.210728, 4.830007, 3.918216, 3.426223, 3.294, 3.187208, 
    2.939013,
  3.680766, 4.143845, 5.099999, 5.334717, 7.064342, 6.177771, 4.800496, 
    7.099148, 8.363858, 8.374338, 8.563765, 7.657479, 7.231249, 6.75156, 
    6.114374, 5.254345, 4.244482, 3.747045, 3.425176, 2.785667, 3.162594, 
    4.758757, 5.858478, 5.966961, 5.514821, 5.045198, 4.736037, 4.272967, 
    3.843482,
  3.448456, 4.703344, 5.472704, 6.810833, 6.253474, 6.402055, 6.432818, 
    5.484677, 6.663951, 7.331388, 7.515093, 6.129117, 5.632715, 5.875918, 
    5.709735, 5.377823, 4.604761, 4.173897, 3.721534, 3.613708, 4.119291, 
    4.576447, 4.535781, 4.319407, 4.551771, 4.526204, 4.399363, 4.120812, 
    3.488352,
  3.044663, 3.116859, 3.710787, 4.494702, 5.043512, 5.147993, 5.164205, 
    4.655643, 4.528216, 5.214457, 5.749984, 4.808895, 4.737588, 4.765659, 
    4.453376, 3.515458, 3.072564, 2.945301, 2.655614, 3.213397, 3.390025, 
    3.326777, 3.500481, 3.133722, 3.472048, 3.469846, 3.303689, 2.921828, 
    2.878625,
  1.911136, 1.810496, 1.902106, 2.285259, 2.346882, 2.303731, 2.588824, 
    2.755759, 2.604765, 2.802373, 2.871317, 3.005195, 2.781696, 2.726484, 
    2.558604, 2.329249, 2.170128, 2.175525, 2.302869, 2.298321, 2.346624, 
    2.355969, 2.565961, 2.391079, 2.5578, 1.644473, 1.28951, 2.381339, 
    2.161356,
  1.623059, 1.564172, 1.581434, 1.649955, 1.800336, 1.922467, 1.998284, 
    2.026703, 2.043769, 2.130707, 2.345179, 2.455933, 2.525374, 2.42253, 
    2.242261, 2.132907, 1.990659, 1.768368, 1.694071, 1.661953, 1.637894, 
    1.637371, 1.447793, 1.428021, 1.473149, 1.203725, 1.388007, 1.727325, 
    1.71283,
  0.2746139, 0.2746139, 0.2746139, 0.2746139, 0.2746139, 0.2746139, 
    0.2746139, 0.2669078, 0.2669078, 0.2669078, 0.2669078, 0.2669078, 
    0.2669078, 0.2669078, 0.268806, 0.268806, 0.268806, 0.268806, 0.268806, 
    0.268806, 0.268806, 0.2820072, 0.2820072, 0.2820072, 0.2820072, 
    0.2820072, 0.2820072, 0.2820072, 0.2746139,
  0.3727483, 0.3279251, 0.3667935, 0.3930373, 0.3802522, 0.3414086, 
    0.2869694, 0.257936, 0.2454858, 0.2291353, 0.2333913, 0.2510113, 
    0.2466894, 0.3331363, 0.4088922, 0.4317844, 0.437504, 0.4701747, 
    0.4851283, 0.4689191, 0.4488498, 0.4314859, 0.4597307, 0.5072574, 
    0.5002428, 0.4815806, 0.4779985, 0.4366732, 0.3903904,
  0.6529615, 0.6500812, 0.7069261, 0.7970302, 0.6972423, 0.6455541, 
    0.6644306, 0.4965887, 0.4306032, 0.4394762, 0.5011855, 0.5532553, 
    0.6756762, 0.8093569, 0.8200565, 0.8297988, 0.841554, 0.7191065, 
    0.6993878, 0.6549487, 0.6578146, 0.6178854, 0.606054, 0.5956763, 
    0.6632734, 0.6440958, 0.6761244, 0.6791121, 0.6553273,
  0.864364, 0.8114491, 0.7869753, 1.002542, 1.257102, 1.225298, 1.182162, 
    0.9948078, 0.8335483, 0.7624599, 0.812209, 0.9935288, 1.273188, 1.673304, 
    1.893283, 1.839225, 1.676293, 1.515918, 1.263633, 1.151109, 0.9444056, 
    0.8348529, 0.761973, 0.7560676, 0.7878165, 0.9015617, 0.9913507, 
    0.9705431, 0.96962,
  1.782931, 1.694295, 1.549989, 1.853873, 2.3661, 2.536448, 2.337605, 
    2.075469, 1.624286, 1.322339, 1.312894, 1.592463, 2.158875, 2.751661, 
    3.137896, 2.784029, 2.521404, 2.013691, 1.718718, 1.518399, 1.369214, 
    1.216787, 1.1256, 0.9879959, 1.07358, 1.613604, 1.794502, 2.044766, 
    2.017936,
  3.08139, 2.897326, 2.874498, 3.771511, 3.8547, 3.671637, 3.454474, 
    3.096325, 2.73278, 2.575648, 2.420312, 2.576566, 3.353467, 3.478951, 
    3.363218, 2.926208, 2.486801, 2.000839, 1.589331, 1.391661, 1.204851, 
    1.055115, 0.9771026, 1.066164, 2.540178, 3.045556, 3.33585, 3.293874, 
    2.986559,
  4.192395, 4.042463, 6.481194, 7.152277, 5.884042, 4.774081, 4.093217, 
    3.527921, 3.08213, 2.903563, 3.611035, 4.509442, 4.288124, 3.715659, 
    3.017585, 2.276086, 1.854318, 1.495285, 1.115515, 0.9009638, 0.8197881, 
    0.9219947, 0.9534466, 1.106727, 4.018848, 5.633604, 6.006808, 5.123041, 
    4.494018,
  6.244009, 9.254482, 11.131, 7.910356, 6.410196, 4.832646, 3.304516, 
    2.719098, 2.845081, 3.769275, 5.193747, 5.389583, 3.843889, 2.741127, 
    2.265167, 1.623108, 1.212305, 0.9103191, 0.751439, 0.6775117, 0.9405102, 
    1.575109, 3.034609, 5.662814, 10.35857, 10.10115, 7.81204, 5.636977, 
    5.573764,
  8.679891, 13.87183, 16.75859, 9.248523, 5.177198, 3.211807, 2.098386, 
    2.381163, 3.432793, 3.917305, 3.493756, 3.656059, 2.509361, 1.417565, 
    1.069873, 0.9116797, 0.8317165, 0.7254353, 0.6862565, 0.7272811, 
    0.9460645, 1.631326, 5.544117, 14.69025, 17.13136, 12.68652, 7.391383, 
    6.08642, 6.673045,
  10.39121, 20.43636, 17.54593, 7.906588, 4.828282, 3.377623, 2.510323, 
    2.509314, 6.330221, 9.024141, 3.020681, 1.548315, 0.89254, 0.6383189, 
    0.587211, 0.5743074, 0.6094956, 0.6672013, 0.7667335, 1.020296, 1.594412, 
    2.43518, 6.883847, 15.8263, 13.04828, 8.35509, 6.556655, 6.644398, 
    8.548992,
  13.19108, 14.15629, 14.31734, 9.839259, 5.134442, 3.991423, 4.546385, 
    4.560201, 5.218657, 3.673978, 2.473958, 1.336138, 1.057054, 1.032005, 
    0.9424413, 1.004998, 0.9730946, 0.9801111, 1.211611, 1.686388, 2.344351, 
    3.427592, 6.495395, 9.964359, 6.78461, 6.366169, 6.655075, 8.324158, 
    13.02604,
  5.561621, 5.587502, 5.648064, 5.99306, 6.466777, 7.051443, 7.965269, 
    8.03332, 9.496622, 6.54891, 4.747293, 3.902757, 3.10435, 2.82454, 
    2.469143, 2.223869, 1.834654, 1.493073, 1.332837, 1.968755, 3.17979, 
    4.893115, 3.72377, 3.80079, 3.633866, 3.275546, 3.53312, 4.40308, 5.547342,
  3.75194, 4.207886, 4.123689, 3.829337, 3.980281, 4.919702, 6.785395, 
    9.181197, 9.836935, 10.96118, 9.324588, 7.308896, 5.767063, 4.955383, 
    4.732858, 4.007487, 3.416847, 2.79606, 2.0346, 2.161481, 4.167181, 
    4.377886, 5.289006, 4.827401, 3.878838, 3.418455, 3.434319, 3.433611, 
    3.124164,
  4.084047, 4.75402, 5.915174, 7.0999, 8.542314, 7.496537, 6.428251, 
    9.176188, 10.38709, 10.21955, 9.968326, 8.739987, 7.973156, 7.303757, 
    6.603507, 5.584297, 4.489537, 3.86311, 3.559246, 3.050935, 3.491424, 
    5.163095, 6.313702, 6.364197, 5.823569, 5.240937, 4.89834, 4.384838, 
    4.057524,
  3.903255, 5.327616, 6.111769, 7.610597, 7.105317, 7.343405, 7.678434, 
    7.009706, 8.152352, 8.593771, 8.339971, 7.026204, 6.398991, 6.500903, 
    6.348231, 5.927543, 5.060523, 4.516041, 4.021008, 4.133159, 4.726934, 
    5.271598, 5.176463, 5.065039, 5.151667, 5.101473, 4.752301, 4.50731, 
    3.886884,
  3.65714, 3.773757, 4.315784, 5.181315, 5.850537, 6.022058, 6.03004, 
    5.531911, 5.434173, 5.991747, 6.544762, 5.88263, 5.643823, 5.481918, 
    5.109142, 4.107209, 3.621578, 3.438653, 3.176524, 3.734779, 3.958969, 
    4.029148, 4.229733, 3.911562, 4.208015, 4.095506, 3.808868, 3.440623, 
    3.388155,
  2.523581, 2.468269, 2.629894, 3.025705, 3.121689, 3.115653, 3.461007, 
    3.602419, 3.434095, 3.599618, 3.633147, 3.765967, 3.49237, 3.438045, 
    3.210068, 2.936261, 2.726559, 2.709923, 2.913316, 2.801494, 2.842805, 
    2.931612, 3.218812, 3.15861, 3.276753, 2.256073, 1.884471, 2.972508, 
    2.773144,
  2.271557, 2.242809, 2.250515, 2.295397, 2.475657, 2.649923, 2.712171, 
    2.787659, 2.803746, 2.884641, 3.13602, 3.174772, 3.222007, 3.073692, 
    2.829038, 2.676485, 2.551195, 2.291808, 2.212017, 2.193499, 2.230403, 
    2.238768, 1.977594, 1.96102, 2.016762, 1.753417, 1.970261, 2.354553, 
    2.34466,
  0.3400338, 0.3400338, 0.3400338, 0.3400338, 0.3400338, 0.3400338, 
    0.3400338, 0.332891, 0.332891, 0.332891, 0.332891, 0.332891, 0.332891, 
    0.332891, 0.3328422, 0.3328422, 0.3328422, 0.3328422, 0.3328422, 
    0.3328422, 0.3328422, 0.3462513, 0.3462513, 0.3462513, 0.3462513, 
    0.3462513, 0.3462513, 0.3462513, 0.3400338,
  0.461947, 0.4135256, 0.4463409, 0.4524766, 0.43427, 0.3900225, 0.3376312, 
    0.311884, 0.2995372, 0.2833656, 0.2874164, 0.3016883, 0.2991545, 
    0.3796794, 0.4525154, 0.4756284, 0.4740666, 0.5171018, 0.5401474, 
    0.5300407, 0.5122544, 0.5033775, 0.5167809, 0.5323768, 0.5238485, 
    0.519143, 0.5171137, 0.498213, 0.4826456,
  0.782528, 0.7488516, 0.7821645, 0.8509312, 0.7878427, 0.7061973, 0.6831311, 
    0.5901217, 0.5144405, 0.5038047, 0.5700551, 0.6482576, 0.7310007, 
    0.8572671, 0.8708935, 0.8851436, 0.9020293, 0.7819328, 0.7702434, 
    0.7167761, 0.7264838, 0.666475, 0.650626, 0.6516398, 0.7124524, 
    0.7067428, 0.7328198, 0.7760863, 0.760368,
  0.9603355, 0.9469079, 0.910336, 1.076768, 1.319187, 1.255375, 1.2258, 
    1.05006, 0.8746718, 0.811664, 0.8613368, 1.050743, 1.336064, 1.782123, 
    1.979162, 1.914416, 1.764523, 1.614378, 1.357514, 1.226982, 1.013489, 
    0.8833833, 0.8009974, 0.8113582, 0.8316246, 0.9757532, 1.079377, 
    1.113292, 1.08423,
  1.868316, 1.731389, 1.573078, 1.88245, 2.289051, 2.419251, 2.244596, 
    2.009741, 1.605938, 1.328766, 1.317929, 1.650938, 2.268188, 2.8582, 
    3.19181, 2.799996, 2.552219, 2.091372, 1.791798, 1.570357, 1.427223, 
    1.262069, 1.163717, 1.045122, 1.139021, 1.680918, 1.863237, 2.073607, 
    2.059404,
  3.028414, 2.879964, 2.877973, 3.680354, 3.702185, 3.519213, 3.305761, 
    2.971454, 2.647566, 2.487768, 2.376138, 2.633884, 3.447652, 3.548643, 
    3.466093, 2.924054, 2.515041, 2.072115, 1.668626, 1.414678, 1.234547, 
    1.070825, 0.9806944, 1.136906, 2.704814, 3.062503, 3.242012, 3.185402, 
    2.901573,
  4.002122, 3.827251, 6.529246, 6.991426, 5.702297, 4.613176, 4.0151, 
    3.480552, 3.170731, 2.979302, 3.685622, 4.511773, 4.477025, 3.774545, 
    3.103997, 2.320198, 1.937785, 1.554799, 1.119678, 0.9274223, 0.8183216, 
    0.8646703, 0.91798, 0.9859015, 4.16011, 5.577082, 5.694052, 4.764986, 
    4.228337,
  5.636996, 8.467481, 10.54848, 7.288817, 5.978696, 4.587395, 3.388561, 
    2.785864, 2.768503, 3.555827, 4.922665, 5.165609, 3.686756, 2.785104, 
    2.288754, 1.667519, 1.226212, 0.9197465, 0.7262049, 0.6621994, 0.89269, 
    1.497217, 2.644593, 4.898136, 9.826302, 9.694384, 7.415865, 5.215246, 
    5.20643,
  7.649066, 12.20744, 15.87267, 8.289123, 4.830972, 3.293855, 2.113158, 
    2.277131, 3.028686, 3.591531, 3.235926, 3.431607, 2.452952, 1.4705, 
    1.07337, 0.9004093, 0.796994, 0.6982033, 0.6530756, 0.6511478, 0.8285424, 
    1.452801, 4.78916, 13.68872, 16.34949, 11.82795, 6.964976, 5.648858, 
    6.329668,
  9.802097, 18.76026, 15.35376, 7.34906, 4.721774, 3.471254, 2.523291, 
    2.465701, 5.700246, 8.383445, 2.904846, 1.491131, 0.8608062, 0.6160876, 
    0.5851133, 0.572737, 0.5972209, 0.6345483, 0.7007278, 0.9679255, 
    1.437844, 2.082745, 5.860304, 14.14685, 11.31962, 7.47193, 6.312641, 
    6.243688, 7.823165,
  12.40252, 13.06256, 13.43729, 9.591409, 4.916296, 3.902263, 4.446747, 
    4.463235, 4.962568, 3.568939, 2.373116, 1.32454, 1.081481, 1.060265, 
    0.9763439, 0.997943, 0.9626339, 0.9672514, 1.180171, 1.604212, 2.190611, 
    3.258795, 5.964619, 8.777264, 5.692736, 5.674991, 6.096435, 7.927472, 
    12.55848,
  5.144383, 5.132381, 5.154216, 5.439108, 5.831545, 6.595485, 7.739224, 
    7.839084, 9.229448, 6.381766, 4.630099, 3.836462, 3.061034, 2.832123, 
    2.43413, 2.250063, 1.802947, 1.486004, 1.348737, 1.95734, 3.037353, 
    4.638451, 3.50529, 3.420802, 3.12988, 2.954717, 3.29956, 4.034349, 5.14606,
  4.080594, 4.519977, 4.400373, 4.130804, 4.195192, 5.06147, 6.806229, 
    9.242518, 10.54526, 11.57006, 9.740415, 7.58363, 5.874583, 5.240223, 
    4.889306, 4.076392, 3.440705, 2.771564, 2.057069, 2.148024, 4.229412, 
    4.397471, 5.237851, 4.758554, 3.811382, 3.374568, 3.515692, 3.606483, 
    3.254585,
  4.417608, 5.183622, 6.523723, 8.456411, 9.5507, 8.494495, 8.040533, 
    11.28936, 12.05267, 11.68701, 10.99774, 9.497806, 8.568919, 7.713648, 
    6.996378, 5.820125, 4.6693, 3.950886, 3.60064, 3.25672, 3.787583, 
    5.411261, 6.574274, 6.637974, 6.039118, 5.353778, 5.003485, 4.421273, 
    4.179565,
  4.205989, 5.791854, 6.582055, 8.068937, 7.643147, 7.906718, 8.428435, 
    8.109058, 9.164827, 9.423868, 8.940636, 7.798676, 7.165462, 6.992316, 
    6.809652, 6.311984, 5.41172, 4.735216, 4.223241, 4.48268, 5.189944, 
    5.67053, 5.678479, 5.696064, 5.627611, 5.566831, 5.010749, 4.833437, 
    4.164663,
  4.119041, 4.340651, 4.797451, 5.643111, 6.373048, 6.567035, 6.653751, 
    6.142104, 6.111531, 6.5752, 7.162213, 6.793679, 6.385514, 6.009429, 
    5.538707, 4.519521, 4.033591, 3.813834, 3.605197, 4.12578, 4.415318, 
    4.471317, 4.916968, 4.584114, 4.835613, 4.668977, 4.22959, 3.86201, 
    3.800257,
  3.038974, 3.016536, 3.231172, 3.662642, 3.823312, 3.883177, 4.236118, 
    4.34058, 4.233106, 4.368762, 4.279008, 4.413491, 4.13687, 4.03594, 
    3.654457, 3.339379, 3.134542, 3.168387, 3.424748, 3.203589, 3.16861, 
    3.408651, 3.765612, 3.864192, 3.949398, 2.871576, 2.465052, 3.497424, 
    3.264322,
  2.830419, 2.804182, 2.785854, 2.866196, 3.12606, 3.310931, 3.40168, 
    3.485211, 3.444314, 3.524375, 3.773105, 3.709136, 3.723393, 3.513185, 
    3.208838, 3.053121, 2.978979, 2.724885, 2.67882, 2.701634, 2.816504, 
    2.834236, 2.524137, 2.506986, 2.544469, 2.256421, 2.487103, 2.928098, 
    2.902523,
  0.3937578, 0.3937578, 0.3937578, 0.3937578, 0.3937578, 0.3937578, 
    0.3937578, 0.3893113, 0.3893113, 0.3893113, 0.3893113, 0.3893113, 
    0.3893113, 0.3893113, 0.3864796, 0.3864796, 0.3864796, 0.3864796, 
    0.3864796, 0.3864796, 0.3864796, 0.3977277, 0.3977277, 0.3977277, 
    0.3977277, 0.3977277, 0.3977277, 0.3977277, 0.3937578,
  0.5203037, 0.4807975, 0.5140924, 0.5069697, 0.4796294, 0.4290342, 0.379979, 
    0.3601641, 0.3459292, 0.3294586, 0.3318241, 0.3398713, 0.3371812, 
    0.3998804, 0.4660767, 0.4945518, 0.4828868, 0.5295399, 0.5627665, 
    0.563212, 0.5529544, 0.5512285, 0.5575789, 0.5398476, 0.5252094, 
    0.5291954, 0.5335438, 0.5407133, 0.5451123,
  0.8631181, 0.8150939, 0.8197379, 0.867335, 0.8364619, 0.7409577, 0.6734882, 
    0.6387807, 0.5599678, 0.5338722, 0.6049219, 0.6930982, 0.7419091, 
    0.843004, 0.8637534, 0.8856853, 0.9041144, 0.801788, 0.7917714, 
    0.7363611, 0.7501655, 0.6775406, 0.6748823, 0.6882424, 0.733677, 
    0.7443761, 0.7726951, 0.8203545, 0.843023,
  1.037951, 1.033985, 0.9966789, 1.126294, 1.333334, 1.251396, 1.20891, 
    1.051262, 0.869121, 0.8107385, 0.8638486, 1.059492, 1.319171, 1.79335, 
    1.96637, 1.903457, 1.776887, 1.65598, 1.399722, 1.247457, 1.040015, 
    0.8949582, 0.8032045, 0.8372949, 0.8522878, 1.022499, 1.158418, 1.2144, 
    1.166356,
  1.909341, 1.709242, 1.559485, 1.842213, 2.14775, 2.255038, 2.097935, 
    1.892116, 1.5329, 1.281847, 1.265234, 1.636319, 2.299682, 2.847514, 
    3.163467, 2.729781, 2.492344, 2.111384, 1.815365, 1.592967, 1.442491, 
    1.273379, 1.171064, 1.083113, 1.188941, 1.71573, 1.927061, 2.029227, 
    2.060444,
  2.868641, 2.727828, 2.774162, 3.533611, 3.499821, 3.325083, 3.104258, 
    2.780075, 2.496888, 2.315445, 2.255345, 2.649422, 3.458749, 3.503747, 
    3.43469, 2.87674, 2.481935, 2.111387, 1.714248, 1.421225, 1.257032, 
    1.075109, 0.9730037, 1.144265, 2.745462, 3.010086, 3.143319, 3.025755, 
    2.774625,
  3.728014, 3.595913, 6.534954, 6.711183, 5.38967, 4.314017, 3.803649, 
    3.341867, 3.123055, 3.022126, 3.733983, 4.456272, 4.524298, 3.782051, 
    3.155024, 2.350579, 1.978984, 1.602984, 1.119228, 0.9376714, 0.8102317, 
    0.7967898, 0.8684233, 0.8745114, 4.328526, 5.436323, 5.249396, 4.356646, 
    3.901015,
  5.108815, 7.735427, 9.94899, 6.683212, 5.463837, 4.272382, 3.391276, 
    2.791222, 2.714808, 3.402889, 4.747637, 4.953676, 3.526489, 2.771909, 
    2.284595, 1.697838, 1.240863, 0.9226891, 0.7128472, 0.6616079, 0.8808852, 
    1.421973, 2.304515, 4.337835, 9.137362, 9.19207, 6.957777, 4.809241, 
    4.827336,
  6.546383, 10.79874, 14.62806, 7.286716, 4.400075, 3.173489, 2.099508, 
    2.20297, 2.656349, 3.337834, 3.060468, 3.286474, 2.385823, 1.484403, 
    1.056012, 0.9054735, 0.784151, 0.6788046, 0.618208, 0.6034804, 0.6846151, 
    1.352601, 4.058325, 12.13796, 15.04238, 10.75606, 6.389822, 5.162256, 
    5.715652,
  9.025406, 16.62432, 13.1185, 6.668154, 4.455058, 3.382239, 2.560083, 
    2.449451, 5.085874, 7.707156, 2.82867, 1.451568, 0.8314769, 0.6087615, 
    0.578274, 0.5623124, 0.5920873, 0.6008821, 0.6410131, 0.9054039, 
    1.193063, 1.684697, 4.741606, 12.32381, 9.337147, 6.596995, 5.935234, 
    5.825277, 7.05448,
  11.74451, 12.09549, 12.76612, 9.066947, 4.674119, 3.900149, 4.355653, 
    4.350357, 4.767793, 3.531685, 2.305302, 1.322021, 1.098312, 1.101872, 
    1.001488, 0.9872457, 0.9512258, 0.9482328, 1.145162, 1.509689, 2.023139, 
    3.093811, 5.279676, 7.555966, 4.711674, 4.827498, 5.402425, 7.394913, 
    11.88042,
  4.743558, 4.657585, 4.675557, 4.881647, 5.219533, 6.101622, 7.411067, 
    7.579707, 8.978621, 6.102695, 4.486382, 3.718322, 2.988409, 2.786789, 
    2.386257, 2.232935, 1.797256, 1.478615, 1.345408, 1.940541, 2.941641, 
    4.311755, 3.274554, 3.105735, 2.752428, 2.655333, 3.088485, 3.703566, 
    4.750679,
  4.272049, 4.748672, 4.630489, 4.449239, 4.427694, 5.198686, 6.882129, 
    9.31824, 11.19054, 12.46719, 10.18668, 7.795072, 5.993123, 5.499152, 
    5.063156, 4.157059, 3.428334, 2.748415, 2.082532, 2.168255, 4.216961, 
    4.409494, 5.058148, 4.631956, 3.682635, 3.285616, 3.581736, 3.691888, 
    3.35088,
  4.667713, 5.468772, 6.781874, 9.330561, 10.18737, 9.1983, 9.579682, 
    12.96513, 13.22436, 12.7689, 11.66879, 9.976063, 8.922718, 8.008839, 
    7.288532, 5.944773, 4.75174, 3.99499, 3.583911, 3.405127, 4.099966, 
    5.545724, 6.618448, 6.700903, 6.143085, 5.370852, 5.017449, 4.445456, 
    4.246196,
  4.428321, 6.071225, 6.9054, 8.255842, 7.963385, 8.185974, 8.834797, 
    8.86883, 9.840635, 9.874949, 9.368991, 8.414694, 7.772703, 7.373474, 
    7.115309, 6.5557, 5.63696, 4.862387, 4.366632, 4.693663, 5.450861, 
    5.875012, 6.115437, 6.337046, 6.047534, 5.910315, 5.214289, 5.031935, 
    4.369622,
  4.473182, 4.826387, 5.199755, 5.975164, 6.665314, 6.844779, 6.99542, 
    6.513265, 6.605614, 7.071177, 7.724676, 7.450423, 6.94845, 6.400595, 
    5.851624, 4.818705, 4.341331, 4.130782, 3.979763, 4.420893, 4.766941, 
    4.799395, 5.488884, 5.224802, 5.44028, 5.15935, 4.60205, 4.203956, 
    4.177738,
  3.477501, 3.449899, 3.706926, 4.164922, 4.439423, 4.555465, 4.927068, 
    5.033401, 4.949574, 5.043692, 4.867571, 4.940172, 4.714603, 4.551793, 
    4.002907, 3.632977, 3.467023, 3.577529, 3.804183, 3.542122, 3.446171, 
    3.827539, 4.272005, 4.437738, 4.545915, 3.495081, 2.995643, 3.947819, 
    3.671372,
  3.286565, 3.241853, 3.209231, 3.373708, 3.682331, 3.88864, 4.042772, 
    4.10978, 4.033033, 4.023966, 4.198084, 4.112487, 4.070609, 3.8555, 
    3.513114, 3.396853, 3.328157, 3.074981, 3.057006, 3.113786, 3.293121, 
    3.36481, 3.097118, 3.047353, 3.073616, 2.712594, 2.974453, 3.441652, 
    3.375371,
  0.4325204, 0.4325204, 0.4325204, 0.4325204, 0.4325204, 0.4325204, 
    0.4325204, 0.4310121, 0.4310121, 0.4310121, 0.4310121, 0.4310121, 
    0.4310121, 0.4310121, 0.4260753, 0.4260753, 0.4260753, 0.4260753, 
    0.4260753, 0.4260753, 0.4260753, 0.4354626, 0.4354626, 0.4354626, 
    0.4354626, 0.4354626, 0.4354626, 0.4354626, 0.4325204,
  0.5530845, 0.5221275, 0.556076, 0.5469766, 0.5114761, 0.4588769, 0.4137249, 
    0.4011768, 0.3815664, 0.3638915, 0.3649014, 0.3678188, 0.3624956, 
    0.3996578, 0.4545629, 0.4883169, 0.4729726, 0.5209468, 0.5630974, 
    0.577622, 0.5768669, 0.584053, 0.5800652, 0.5364559, 0.5146989, 
    0.5210072, 0.5336189, 0.5648348, 0.5830774,
  0.8784308, 0.8284522, 0.8243164, 0.8577892, 0.8524404, 0.7561739, 
    0.6540225, 0.6527709, 0.5742621, 0.5407292, 0.6209941, 0.7004344, 
    0.7210889, 0.7931874, 0.8220918, 0.8553354, 0.8596045, 0.7824497, 
    0.7579116, 0.7232425, 0.7413725, 0.6641707, 0.673441, 0.7027241, 
    0.7412553, 0.7488228, 0.7799458, 0.8258613, 0.8786144,
  1.099274, 1.089727, 1.034433, 1.138875, 1.315893, 1.231657, 1.163409, 
    1.012881, 0.8379458, 0.7843077, 0.8445558, 1.04039, 1.261508, 1.733783, 
    1.911886, 1.833832, 1.733258, 1.616644, 1.400908, 1.223145, 1.031245, 
    0.8758854, 0.787817, 0.840226, 0.8582979, 1.053355, 1.225309, 1.28859, 
    1.211248,
  1.901558, 1.666946, 1.539646, 1.791481, 2.012236, 2.079059, 1.933948, 
    1.743066, 1.427225, 1.209121, 1.185119, 1.592529, 2.275218, 2.776135, 
    3.045685, 2.618048, 2.381641, 2.082037, 1.80264, 1.586937, 1.429481, 
    1.262018, 1.152078, 1.096378, 1.227502, 1.729325, 1.97504, 1.977501, 
    2.0368,
  2.64362, 2.53726, 2.637818, 3.380511, 3.264285, 3.064141, 2.876552, 
    2.540281, 2.314992, 2.160046, 2.117398, 2.619422, 3.411747, 3.451015, 
    3.324591, 2.813598, 2.438023, 2.10086, 1.735358, 1.425513, 1.268569, 
    1.070061, 0.9666632, 1.115093, 2.719457, 2.90806, 3.055659, 2.877004, 
    2.596747,
  3.395198, 3.328271, 6.315257, 6.35939, 4.994778, 3.951138, 3.528095, 
    3.183634, 3.003001, 2.954626, 3.674074, 4.307233, 4.444459, 3.714036, 
    3.127932, 2.336431, 1.974022, 1.618728, 1.122732, 0.9253114, 0.7939896, 
    0.7198704, 0.811063, 0.8250797, 4.417448, 5.307276, 4.750098, 3.971572, 
    3.572085,
  4.71836, 7.105305, 9.434324, 6.179699, 4.945186, 3.930537, 3.257256, 
    2.700529, 2.633065, 3.337066, 4.697465, 4.88082, 3.386026, 2.713171, 
    2.24938, 1.709385, 1.253749, 0.9232731, 0.7317854, 0.6562095, 0.8740377, 
    1.306882, 2.001428, 3.94069, 8.50409, 8.590731, 6.403815, 4.337595, 
    4.433753,
  5.696567, 9.691069, 13.23312, 6.318211, 3.963343, 2.903451, 2.015294, 
    2.140941, 2.408309, 3.252484, 2.963545, 3.250189, 2.280615, 1.443133, 
    1.031895, 0.8982916, 0.7889514, 0.6575456, 0.5867811, 0.5810171, 
    0.5959433, 1.276441, 3.508183, 10.72565, 13.5293, 9.86881, 5.778311, 
    4.665468, 5.036414,
  8.242556, 14.64342, 11.43656, 5.91141, 4.0373, 3.186824, 2.612504, 2.42126, 
    4.628978, 7.162929, 2.811652, 1.462224, 0.8001531, 0.5860153, 0.5709838, 
    0.5800492, 0.5838824, 0.582876, 0.5866611, 0.8325326, 0.9850876, 
    1.366872, 3.772625, 10.59566, 7.802255, 5.761933, 5.372353, 5.292924, 
    6.39783,
  11.13785, 11.4197, 12.34663, 8.345603, 4.444668, 3.897576, 4.242194, 
    4.278856, 4.630316, 3.486744, 2.352701, 1.339932, 1.130513, 1.157509, 
    1.012455, 0.9876533, 0.9469056, 0.9236642, 1.096273, 1.418583, 1.86489, 
    2.944805, 4.693076, 6.537916, 3.808118, 4.082255, 4.723114, 6.838889, 
    11.20767,
  4.251633, 4.108899, 4.176141, 4.54794, 4.796462, 5.637872, 7.115407, 
    7.318758, 8.706761, 5.809544, 4.349022, 3.555854, 2.897539, 2.735958, 
    2.319088, 2.207668, 1.782851, 1.46367, 1.340096, 1.892683, 2.850398, 
    4.007439, 3.094939, 2.858375, 2.43304, 2.421839, 2.922376, 3.484999, 
    4.373023,
  4.411264, 4.943387, 4.877542, 4.728271, 4.649241, 5.397492, 7.300705, 
    9.452092, 11.78539, 13.78443, 10.77893, 7.983217, 6.170543, 5.696476, 
    5.150958, 4.163903, 3.352001, 2.721284, 2.0988, 2.25251, 4.176067, 
    4.34441, 4.909613, 4.468341, 3.526661, 3.179248, 3.62847, 3.687675, 
    3.402762,
  4.795475, 5.69818, 6.934415, 9.752322, 10.66306, 9.559731, 10.97169, 
    14.14744, 13.96693, 13.39215, 11.97785, 10.18861, 9.102845, 8.21279, 
    7.484132, 5.981049, 4.817616, 3.996555, 3.548661, 3.498795, 4.353454, 
    5.749053, 6.560233, 6.653193, 6.151642, 5.325995, 4.948149, 4.439757, 
    4.26171,
  4.599635, 6.235183, 7.087285, 8.298123, 8.075398, 8.270389, 8.955807, 
    9.38464, 10.29611, 10.20411, 9.638931, 8.977235, 8.258209, 7.652251, 
    7.320266, 6.663729, 5.727284, 4.968393, 4.470477, 4.832879, 5.664136, 
    6.11265, 6.495359, 6.827219, 6.473472, 6.147682, 5.414562, 5.162256, 
    4.510508,
  4.75684, 5.17554, 5.564558, 6.254543, 6.824498, 7.072005, 7.231897, 
    6.771847, 6.993881, 7.529334, 8.317775, 7.913552, 7.358452, 6.711216, 
    6.097567, 5.056541, 4.561369, 4.434012, 4.305553, 4.616304, 5.109983, 
    5.0802, 5.835326, 5.818944, 6.020712, 5.626283, 4.931209, 4.520707, 
    4.510167,
  3.837094, 3.815664, 4.105026, 4.609357, 5.024979, 5.258738, 5.645344, 
    5.755263, 5.582703, 5.618545, 5.438346, 5.395959, 5.20257, 5.019438, 
    4.287382, 3.897973, 3.802326, 3.973275, 4.097262, 3.845699, 3.69999, 
    4.207778, 4.774868, 4.943185, 4.997861, 4.095875, 3.470961, 4.29848, 
    3.985532,
  3.693497, 3.666705, 3.660012, 3.927458, 4.173444, 4.3672, 4.588754, 
    4.645626, 4.585178, 4.464188, 4.476119, 4.367301, 4.257061, 4.071689, 
    3.735711, 3.666884, 3.611382, 3.370675, 3.361062, 3.453127, 3.678566, 
    3.772087, 3.570629, 3.532796, 3.576403, 3.175147, 3.451523, 3.865098, 
    3.770058,
  0.4566895, 0.4566895, 0.4566895, 0.4566895, 0.4566895, 0.4566895, 
    0.4566895, 0.4574845, 0.4574845, 0.4574845, 0.4574845, 0.4574845, 
    0.4574845, 0.4574845, 0.4526393, 0.4526393, 0.4526393, 0.4526393, 
    0.4526393, 0.4526393, 0.4526393, 0.4604472, 0.4604472, 0.4604472, 
    0.4604472, 0.4604472, 0.4604472, 0.4604472, 0.4566895,
  0.5711287, 0.5427616, 0.5763441, 0.5694143, 0.5311898, 0.4793175, 0.439573, 
    0.4323424, 0.4059372, 0.3887679, 0.387179, 0.3846391, 0.3766477, 
    0.3863649, 0.4270599, 0.4674393, 0.4518604, 0.4941733, 0.54313, 
    0.5730301, 0.5855883, 0.5982819, 0.5811958, 0.5235308, 0.5016569, 
    0.5059797, 0.5332392, 0.5773697, 0.6030506,
  0.8542596, 0.8033665, 0.8049258, 0.8194463, 0.85559, 0.757603, 0.6212102, 
    0.6432828, 0.5672529, 0.5317793, 0.6186477, 0.6873453, 0.6811923, 
    0.7262602, 0.7603605, 0.8061819, 0.793813, 0.7434726, 0.7022779, 
    0.6941423, 0.7062951, 0.6424984, 0.6593451, 0.6915748, 0.7253641, 
    0.7183812, 0.7615727, 0.8177521, 0.8732135,
  1.137516, 1.123599, 1.045963, 1.122654, 1.279802, 1.200921, 1.105598, 
    0.9493628, 0.8003629, 0.7482378, 0.8156843, 0.9989235, 1.175014, 
    1.655611, 1.841192, 1.752632, 1.663448, 1.531057, 1.351953, 1.157254, 
    0.9855127, 0.8388664, 0.7662446, 0.8240913, 0.8591648, 1.066568, 
    1.249854, 1.298984, 1.22482,
  1.859027, 1.613671, 1.510182, 1.716821, 1.902417, 1.925008, 1.782382, 
    1.601498, 1.313118, 1.122846, 1.103915, 1.526797, 2.222612, 2.675726, 
    2.864108, 2.487446, 2.244328, 1.999093, 1.735635, 1.540222, 1.379027, 
    1.22854, 1.110551, 1.100843, 1.286248, 1.734438, 2.042218, 1.946027, 
    2.021415,
  2.394108, 2.351785, 2.485796, 3.229028, 3.031382, 2.781578, 2.626678, 
    2.288017, 2.099548, 2.004267, 2.013376, 2.551006, 3.326006, 3.394892, 
    3.18977, 2.730046, 2.369348, 2.041802, 1.732134, 1.429003, 1.254327, 
    1.062705, 0.9580288, 1.094798, 2.716784, 2.847116, 2.923985, 2.699009, 
    2.418091,
  3.061027, 3.062835, 5.960181, 6.015786, 4.590557, 3.57814, 3.184294, 
    2.97313, 2.848376, 2.863262, 3.720979, 4.269936, 4.283789, 3.623276, 
    3.023857, 2.258856, 1.919112, 1.607965, 1.119361, 0.9125839, 0.778891, 
    0.6616933, 0.7469282, 0.8072252, 4.540248, 5.240351, 4.314231, 3.538479, 
    3.203548,
  4.351953, 6.674463, 9.012124, 5.670794, 4.4591, 3.572324, 3.034633, 
    2.630286, 2.554917, 3.227822, 4.711426, 4.922196, 3.288652, 2.657356, 
    2.184316, 1.678421, 1.246114, 0.9137277, 0.736164, 0.6462807, 0.853148, 
    1.151818, 1.66632, 3.768085, 8.256317, 8.119293, 5.831427, 3.88992, 
    4.029309,
  5.046947, 8.939305, 11.79278, 5.715225, 3.51502, 2.599058, 1.904741, 
    2.039684, 2.281201, 3.233307, 2.887004, 3.155127, 2.179358, 1.33746, 
    1.001195, 0.8912127, 0.7811641, 0.6330927, 0.5428651, 0.5526796, 
    0.5624905, 1.190432, 3.185885, 9.923793, 12.20995, 9.039718, 5.121964, 
    4.163908, 4.495354,
  7.852869, 13.97919, 10.5828, 5.289619, 3.480814, 2.916604, 2.556282, 
    2.393167, 4.414092, 6.796532, 2.882729, 1.484176, 0.7597736, 0.5516783, 
    0.5529896, 0.6117288, 0.5709015, 0.5513504, 0.5452176, 0.7441347, 
    0.8798062, 1.142327, 3.145042, 9.585656, 7.07273, 5.069935, 4.784773, 
    4.752694, 5.826523,
  10.77478, 11.10744, 12.20858, 7.664881, 4.180099, 3.861644, 4.110362, 
    4.195029, 4.549469, 3.441076, 2.353522, 1.345798, 1.23208, 1.17987, 
    1.023713, 1.005519, 0.9381325, 0.903463, 1.082383, 1.359898, 1.763949, 
    2.774154, 4.323249, 5.810485, 3.111641, 3.373402, 4.176164, 6.378967, 
    10.9073,
  3.796856, 3.663868, 3.817134, 4.575102, 4.647007, 5.327573, 6.87278, 
    7.089942, 8.561265, 5.59989, 4.14162, 3.387687, 2.803016, 2.680532, 
    2.27474, 2.18555, 1.766302, 1.441547, 1.372632, 1.812768, 2.771352, 
    3.808831, 2.940766, 2.646292, 2.208874, 2.269232, 2.820445, 3.424783, 
    3.963856,
  4.55957, 5.193532, 5.173814, 4.973637, 4.814301, 5.691093, 7.912659, 
    9.642467, 12.29237, 15.37782, 11.37796, 8.255791, 6.458133, 5.896044, 
    5.187654, 4.113202, 3.269722, 2.670115, 2.114562, 2.310758, 4.116388, 
    4.263433, 4.815001, 4.310573, 3.343666, 3.05179, 3.618651, 3.65692, 
    3.483365,
  4.862641, 5.84576, 7.035777, 9.902555, 11.13786, 9.766607, 12.22998, 
    15.03611, 14.41878, 13.61545, 12.03297, 10.26447, 9.13161, 8.333636, 
    7.528257, 5.962193, 4.88043, 3.993531, 3.560468, 3.550073, 4.507407, 
    6.035593, 6.519628, 6.596922, 6.198939, 5.235445, 4.826378, 4.341347, 
    4.271193,
  4.712477, 6.375408, 7.134888, 8.194932, 8.065526, 8.313237, 8.881264, 
    9.689843, 10.5955, 10.48607, 9.903831, 9.470532, 8.634185, 7.811647, 
    7.478981, 6.687869, 5.775164, 5.059986, 4.546321, 4.937952, 5.846246, 
    6.36084, 6.854889, 7.220408, 6.98551, 6.321441, 5.570954, 5.320673, 
    4.601205,
  4.942847, 5.447204, 5.872201, 6.455339, 6.968751, 7.306682, 7.462204, 
    7.022607, 7.322061, 7.940141, 8.845492, 8.278555, 7.708845, 6.972486, 
    6.330331, 5.237732, 4.744461, 4.661531, 4.558434, 4.723095, 5.327284, 
    5.294932, 6.057848, 6.299499, 6.558009, 6.056461, 5.232868, 4.79917, 
    4.749617,
  4.125039, 4.16842, 4.438643, 4.970079, 5.57959, 5.897201, 6.288508, 
    6.488413, 6.197021, 6.112978, 5.930563, 5.825152, 5.564548, 5.397376, 
    4.547482, 4.172198, 4.057134, 4.275329, 4.317525, 4.121638, 3.970028, 
    4.529582, 5.160549, 5.362216, 5.351521, 4.61967, 3.8946, 4.575853, 
    4.215199,
  4.078656, 4.091588, 4.144245, 4.424631, 4.55011, 4.733267, 4.961396, 
    5.051036, 4.983548, 4.812764, 4.676078, 4.496138, 4.361832, 4.175205, 
    3.86121, 3.858229, 3.798719, 3.621141, 3.619735, 3.746908, 3.979288, 
    4.071201, 3.905928, 3.901141, 3.998456, 3.60855, 3.875726, 4.253025, 
    4.151702,
  0.4699539, 0.4699539, 0.4699539, 0.4699539, 0.4699539, 0.4699539, 
    0.4699539, 0.4701157, 0.4701157, 0.4701157, 0.4701157, 0.4701157, 
    0.4701157, 0.4701157, 0.4668365, 0.4668365, 0.4668365, 0.4668365, 
    0.4668365, 0.4668365, 0.4668365, 0.4714731, 0.4714731, 0.4714731, 
    0.4714731, 0.4714731, 0.4714731, 0.4714731, 0.4699539,
  0.5839799, 0.5554429, 0.5834219, 0.5722892, 0.5356314, 0.4897521, 
    0.4554337, 0.4489895, 0.4170688, 0.4028795, 0.398369, 0.3917546, 
    0.3809282, 0.3665041, 0.390607, 0.4311866, 0.4206865, 0.4567364, 
    0.5084146, 0.552249, 0.5742876, 0.5922484, 0.567172, 0.5027593, 
    0.4850186, 0.4914811, 0.5318471, 0.5811702, 0.6124994,
  0.812977, 0.7762913, 0.7635083, 0.7673215, 0.8478259, 0.7410184, 0.5743976, 
    0.6175874, 0.5484488, 0.5132927, 0.5992953, 0.6588254, 0.6249581, 
    0.6629385, 0.6953503, 0.7433149, 0.7225552, 0.6901164, 0.6418202, 
    0.6542487, 0.6541021, 0.6150223, 0.6345068, 0.6547831, 0.6933362, 
    0.6776059, 0.7342539, 0.80843, 0.8430674,
  1.14124, 1.133576, 1.04742, 1.093858, 1.230637, 1.159243, 1.042529, 
    0.8833058, 0.7550303, 0.7128133, 0.7731689, 0.9529107, 1.086817, 
    1.580155, 1.757321, 1.663604, 1.588856, 1.416665, 1.259167, 1.070065, 
    0.9087878, 0.7907515, 0.7354135, 0.7891794, 0.8547833, 1.051746, 
    1.244154, 1.253285, 1.213552,
  1.801213, 1.544331, 1.463848, 1.636062, 1.809656, 1.785978, 1.634355, 
    1.472532, 1.203657, 1.032711, 1.030801, 1.459018, 2.174246, 2.558165, 
    2.67189, 2.377548, 2.109674, 1.868633, 1.625935, 1.452621, 1.289726, 
    1.16769, 1.049773, 1.097845, 1.361739, 1.763582, 2.100877, 1.933591, 
    2.018628,
  2.184741, 2.175092, 2.319765, 3.109607, 2.814296, 2.51072, 2.361084, 
    2.06528, 1.885076, 1.873984, 1.923449, 2.486861, 3.295145, 3.34667, 
    3.028356, 2.584896, 2.289915, 1.979819, 1.696113, 1.412284, 1.24183, 
    1.052041, 0.9456539, 1.0786, 2.860064, 2.849957, 2.812329, 2.504746, 
    2.234355,
  2.769576, 2.80429, 5.62926, 5.795543, 4.235927, 3.203325, 2.862166, 2.7128, 
    2.672247, 2.776614, 3.804225, 4.34533, 4.168446, 3.546294, 2.875295, 
    2.161227, 1.802108, 1.547148, 1.094386, 0.8989028, 0.7452896, 0.622134, 
    0.6831788, 0.8377506, 4.921071, 5.228261, 3.972079, 3.137699, 2.876934,
  3.975917, 6.486623, 8.709361, 5.240482, 4.049073, 3.184502, 2.869919, 
    2.545635, 2.428331, 3.206706, 4.778995, 5.056442, 3.181198, 2.596652, 
    2.095997, 1.583984, 1.199734, 0.8962615, 0.7089842, 0.6668099, 0.812991, 
    0.9717089, 1.382428, 3.811913, 8.206704, 7.804356, 5.281414, 3.511148, 
    3.583665,
  4.550753, 8.531756, 10.67377, 5.351205, 3.109226, 2.296103, 1.782353, 
    1.925915, 2.12118, 3.178724, 2.852902, 3.080067, 2.112634, 1.243667, 
    0.9740933, 0.8772366, 0.7416499, 0.5933843, 0.503723, 0.5056056, 
    0.5859005, 1.206179, 3.047511, 9.786186, 11.20205, 8.255254, 4.400991, 
    3.642137, 4.03253,
  8.017497, 14.5126, 10.86951, 4.909446, 2.955675, 2.570158, 2.442113, 
    2.357221, 4.436761, 6.531197, 2.971211, 1.51374, 0.7358541, 0.5414076, 
    0.53172, 0.6108835, 0.5470682, 0.500547, 0.5380108, 0.6660923, 0.784121, 
    1.071194, 3.014425, 9.472933, 7.111104, 4.568059, 4.337126, 4.360242, 
    5.600994,
  10.7446, 11.15667, 12.09246, 7.328062, 4.042887, 3.779081, 4.035774, 
    4.186368, 4.514758, 3.406708, 2.309966, 1.326573, 1.299398, 1.166759, 
    1.003242, 0.9909721, 0.9090637, 0.8937061, 1.084681, 1.308066, 1.711851, 
    2.663901, 4.159007, 5.350575, 2.654284, 2.904933, 3.808538, 6.139402, 
    11.27189,
  3.704417, 3.500316, 3.695979, 5.062934, 4.75153, 5.298929, 6.689553, 
    6.873973, 8.600084, 5.449476, 3.921544, 3.202303, 2.690157, 2.58342, 
    2.226965, 2.149252, 1.709744, 1.417853, 1.426691, 1.737903, 2.76576, 
    3.720207, 2.80155, 2.423566, 2.083747, 2.237288, 2.764527, 3.414859, 
    3.802904,
  4.947374, 5.498234, 5.442049, 5.371847, 5.072678, 6.125146, 8.982223, 
    9.909881, 12.93021, 17.05208, 11.88967, 8.576835, 6.791417, 6.045424, 
    5.1813, 4.067083, 3.215824, 2.630363, 2.127177, 2.343163, 4.103227, 
    4.296757, 4.755686, 4.170743, 3.170841, 2.915768, 3.585602, 3.602459, 
    3.768256,
  5.010291, 6.042215, 7.132606, 9.905917, 11.6538, 9.930068, 13.33041, 
    15.81856, 14.74119, 13.58018, 11.94613, 10.28964, 9.13508, 8.334894, 
    7.454418, 5.944027, 4.897572, 4.013875, 3.585366, 3.592946, 4.734265, 
    6.609834, 6.606481, 6.612386, 6.312882, 5.186114, 4.695888, 4.214007, 
    4.288721,
  4.804242, 6.525459, 7.107881, 7.953917, 8.016752, 8.329775, 8.794777, 
    9.793442, 10.74761, 10.77964, 10.4468, 10.01029, 8.900847, 7.972919, 
    7.628987, 6.693358, 5.802443, 5.074379, 4.558937, 4.910013, 6.029697, 
    6.676072, 7.263497, 7.732676, 7.579132, 6.494808, 5.73106, 5.436979, 
    4.689396,
  5.056105, 5.657963, 6.096137, 6.582874, 7.104733, 7.497939, 7.711018, 
    7.343352, 7.680278, 8.373546, 9.306559, 8.667722, 8.04243, 7.2315, 
    6.555599, 5.386776, 4.897704, 4.810305, 4.707059, 4.856502, 5.432277, 
    5.489795, 6.28735, 6.621856, 6.988031, 6.419792, 5.547928, 5.030985, 
    4.92296,
  4.396319, 4.490349, 4.758777, 5.290122, 6.02793, 6.418196, 6.716961, 
    7.124038, 6.806823, 6.553972, 6.364434, 6.180657, 5.806173, 5.677464, 
    4.802919, 4.425048, 4.24649, 4.509094, 4.494838, 4.352341, 4.226938, 
    4.777161, 5.452688, 5.705951, 5.667251, 5.08615, 4.299075, 4.803057, 
    4.407687,
  4.391542, 4.395107, 4.539282, 4.753533, 4.819818, 4.984812, 5.236513, 
    5.371452, 5.193628, 5.026927, 4.858951, 4.639374, 4.480597, 4.247345, 
    3.974503, 4.042168, 3.927703, 3.792566, 3.803935, 3.958609, 4.199784, 
    4.296675, 4.162125, 4.207261, 4.357117, 3.991265, 4.257928, 4.637245, 
    4.480775,
  0.4766698, 0.4766698, 0.4766698, 0.4766698, 0.4766698, 0.4766698, 
    0.4766698, 0.471012, 0.471012, 0.471012, 0.471012, 0.471012, 0.471012, 
    0.471012, 0.4680237, 0.4680237, 0.4680237, 0.4680237, 0.4680237, 
    0.4680237, 0.4680237, 0.4715536, 0.4715536, 0.4715536, 0.4715536, 
    0.4715536, 0.4715536, 0.4715536, 0.4766698,
  0.5926505, 0.5604157, 0.5797786, 0.5603889, 0.524875, 0.4878571, 0.4587584, 
    0.4517039, 0.4198593, 0.4066033, 0.3973396, 0.3883115, 0.3766981, 
    0.3444407, 0.3539944, 0.3854815, 0.3842064, 0.4154218, 0.4689517, 
    0.523367, 0.5541945, 0.569901, 0.5455113, 0.4815719, 0.466411, 0.4742585, 
    0.5264774, 0.5742795, 0.6152055,
  0.7803352, 0.7389006, 0.7154014, 0.7126518, 0.8176958, 0.7051517, 
    0.5272009, 0.5833297, 0.5180351, 0.4907337, 0.5689426, 0.6211457, 
    0.5669785, 0.5978792, 0.6361549, 0.6734821, 0.651769, 0.6332565, 
    0.5849332, 0.6057189, 0.6018656, 0.5760337, 0.6049801, 0.6036525, 
    0.655931, 0.6403492, 0.7089605, 0.799409, 0.8017275,
  1.125272, 1.123545, 1.034037, 1.049652, 1.158788, 1.102177, 0.9757357, 
    0.8282362, 0.7051396, 0.6658728, 0.71873, 0.9021904, 0.9998171, 1.495196, 
    1.660933, 1.571764, 1.491622, 1.290849, 1.150059, 0.977647, 0.8308877, 
    0.7414401, 0.6949257, 0.746978, 0.8500191, 1.029805, 1.228206, 1.219225, 
    1.181272,
  1.751141, 1.477342, 1.398597, 1.555725, 1.717374, 1.651021, 1.4918, 
    1.338266, 1.10154, 0.9526736, 0.9668054, 1.382635, 2.097573, 2.423093, 
    2.515535, 2.250924, 1.986759, 1.727418, 1.509345, 1.339832, 1.185603, 
    1.077447, 0.9835991, 1.092899, 1.428825, 1.795496, 2.159406, 1.934187, 
    2.000286,
  2.034203, 1.989509, 2.167839, 3.017998, 2.630413, 2.282779, 2.091764, 
    1.876288, 1.694824, 1.735604, 1.855964, 2.454362, 3.347944, 3.303199, 
    2.89357, 2.409534, 2.195799, 1.921604, 1.654039, 1.389549, 1.212978, 
    1.026634, 0.9145305, 1.069963, 3.218853, 2.924179, 2.72041, 2.347016, 
    2.094606,
  2.516484, 2.59157, 5.475379, 5.718989, 3.95545, 2.889252, 2.596654, 
    2.425574, 2.466237, 2.696626, 3.986571, 4.404936, 4.126374, 3.51434, 
    2.678394, 2.059381, 1.666937, 1.468648, 1.071475, 0.8728585, 0.7139598, 
    0.6018159, 0.6428404, 0.9064614, 5.609509, 5.365659, 3.729697, 2.818956, 
    2.582103,
  3.540884, 6.551917, 8.559237, 4.88671, 3.762001, 2.798482, 2.702746, 
    2.387021, 2.284631, 3.292043, 5.051119, 5.202121, 3.085604, 2.520533, 
    2.012692, 1.442508, 1.108403, 0.8593519, 0.6843398, 0.6674194, 0.7729633, 
    0.8739584, 1.260212, 3.991319, 8.665265, 7.654593, 4.766534, 3.277206, 
    3.220579,
  4.146886, 8.656491, 10.19736, 5.098512, 2.773178, 2.042883, 1.613485, 
    1.815173, 1.97, 3.090216, 2.851975, 3.039169, 2.058175, 1.112854, 
    0.9159755, 0.8340179, 0.6750454, 0.5506753, 0.4845578, 0.4801794, 
    0.6190795, 1.269746, 3.30144, 10.29901, 10.62635, 7.932316, 3.855798, 
    3.186438, 3.566586,
  8.748143, 15.95902, 12.50192, 4.54919, 2.655874, 2.316686, 2.297144, 
    2.345254, 4.451712, 6.41601, 3.00214, 1.542748, 0.7272087, 0.5244916, 
    0.5039153, 0.5574408, 0.5063361, 0.4652764, 0.514979, 0.6481999, 
    0.7301158, 1.075874, 3.670371, 10.08045, 7.58885, 4.527048, 4.032783, 
    4.141278, 5.754125,
  11.17085, 11.43465, 12.22997, 7.622319, 4.20963, 3.741237, 4.137381, 
    4.256421, 4.476694, 3.365829, 2.291085, 1.268502, 1.284601, 1.125224, 
    0.95435, 0.9832091, 0.8835259, 0.9076332, 1.092106, 1.299558, 1.69234, 
    2.629452, 4.137124, 5.010365, 2.364892, 2.681204, 3.616113, 6.258617, 
    11.8486,
  4.336099, 3.751413, 3.909232, 6.570135, 5.232109, 5.618243, 6.615396, 
    6.824767, 8.601805, 5.341694, 3.732478, 3.035833, 2.567178, 2.482882, 
    2.173925, 2.073612, 1.654952, 1.448076, 1.474778, 1.737414, 2.877676, 
    3.78919, 2.690104, 2.204001, 1.98895, 2.219482, 2.839038, 3.69172, 
    4.300675,
  5.636118, 6.027264, 5.714109, 6.027271, 5.710399, 6.800815, 10.13827, 
    10.27866, 13.74857, 18.64916, 12.44326, 8.921369, 7.062357, 6.066636, 
    5.112845, 4.03733, 3.202675, 2.582065, 2.104651, 2.433676, 4.179052, 
    4.541543, 4.846489, 4.075306, 3.056915, 2.814897, 3.560799, 3.591737, 
    4.374545,
  5.290497, 6.383416, 7.258054, 9.978364, 12.5024, 10.13424, 14.3457, 
    16.65436, 15.07301, 13.49719, 11.91351, 10.29263, 9.147167, 8.207702, 
    7.339415, 5.95477, 4.816895, 4.010345, 3.568989, 3.604704, 5.271688, 
    7.526985, 6.876481, 6.786376, 6.586533, 5.192799, 4.58178, 4.109871, 
    4.36797,
  4.895421, 6.715327, 7.085254, 7.826522, 8.102341, 8.425992, 8.807813, 
    9.779819, 10.88582, 11.27015, 11.23276, 10.62467, 9.136477, 8.186093, 
    7.711472, 6.650942, 5.779974, 5.011487, 4.497973, 4.892419, 6.291799, 
    7.136055, 7.812615, 8.471246, 8.142515, 6.702418, 5.897441, 5.507174, 
    4.753832,
  5.184929, 5.857223, 6.31592, 6.731816, 7.28258, 7.711749, 7.947014, 
    7.741004, 8.222425, 8.823947, 9.837689, 9.137789, 8.331761, 7.481809, 
    6.750835, 5.49538, 5.015329, 4.929355, 4.90063, 5.082947, 5.542843, 
    5.784896, 6.543291, 6.905235, 7.442043, 6.764726, 5.832481, 5.206649, 
    5.069519,
  4.674776, 4.790226, 5.083358, 5.574837, 6.385663, 6.835801, 6.971652, 
    7.568056, 7.343653, 7.004836, 6.742162, 6.483757, 5.980071, 5.858423, 
    5.020136, 4.612715, 4.439556, 4.712922, 4.666876, 4.557816, 4.407651, 
    4.984712, 5.696652, 5.98582, 5.936888, 5.49395, 4.678697, 5.008869, 
    4.599174,
  4.604337, 4.547444, 4.795751, 4.940432, 5.028892, 5.170306, 5.496583, 
    5.588703, 5.321778, 5.133413, 4.969086, 4.74245, 4.58164, 4.278612, 
    4.046103, 4.113711, 4.018752, 3.901574, 3.907391, 4.082103, 4.374152, 
    4.477482, 4.383955, 4.501878, 4.671377, 4.326209, 4.587308, 4.947544, 
    4.706725,
  0.4749982, 0.4749982, 0.4749982, 0.4749982, 0.4749982, 0.4749982, 
    0.4749982, 0.4645359, 0.4645359, 0.4645359, 0.4645359, 0.4645359, 
    0.4645359, 0.4645359, 0.4605221, 0.4605221, 0.4605221, 0.4605221, 
    0.4605221, 0.4605221, 0.4605221, 0.4649793, 0.4649793, 0.4649793, 
    0.4649793, 0.4649793, 0.4649793, 0.4649793, 0.4749982,
  0.5966731, 0.5570363, 0.5678756, 0.5415238, 0.5064216, 0.4745297, 0.449858, 
    0.4438086, 0.4164468, 0.3995266, 0.3853038, 0.3749329, 0.3678446, 
    0.3202361, 0.3220128, 0.3438917, 0.3482691, 0.3775717, 0.4300057, 
    0.4920928, 0.5271313, 0.5477555, 0.5232764, 0.4668871, 0.4505792, 
    0.458984, 0.5173393, 0.5574056, 0.6131986,
  0.7458328, 0.6876853, 0.6653336, 0.6571238, 0.7745381, 0.6584947, 0.480255, 
    0.5437572, 0.4851277, 0.4618633, 0.5317921, 0.5859125, 0.5164876, 
    0.5364054, 0.5818872, 0.6091763, 0.5851395, 0.5734202, 0.5300022, 
    0.5485466, 0.5493328, 0.5273955, 0.577208, 0.5603887, 0.6228695, 
    0.6072914, 0.6824022, 0.7852635, 0.7617489,
  1.093178, 1.094083, 1.002709, 0.9912186, 1.088476, 1.041929, 0.9076102, 
    0.7665887, 0.6483049, 0.6133454, 0.6654645, 0.8468695, 0.9283509, 
    1.399797, 1.567056, 1.499075, 1.388331, 1.181021, 1.039604, 0.8866774, 
    0.765395, 0.6986542, 0.6495163, 0.7036347, 0.8425292, 1.029184, 1.22178, 
    1.213746, 1.147952,
  1.697073, 1.419907, 1.339326, 1.474449, 1.623466, 1.530664, 1.363139, 
    1.217404, 1.006962, 0.8752428, 0.9061118, 1.313548, 2.00376, 2.272384, 
    2.405501, 2.107524, 1.850238, 1.585846, 1.393887, 1.219764, 1.082344, 
    0.9777809, 0.899717, 1.072831, 1.470643, 1.868271, 2.215857, 1.942746, 
    1.951772,
  1.898664, 1.841836, 2.020777, 2.954955, 2.495671, 2.067268, 1.850701, 
    1.677841, 1.524286, 1.582089, 1.81918, 2.469388, 3.474826, 3.230136, 
    2.77249, 2.234808, 2.086641, 1.827149, 1.593847, 1.355737, 1.171647, 
    0.9769747, 0.8849006, 1.062694, 3.772709, 3.060987, 2.661633, 2.251563, 
    1.978282,
  2.292392, 2.491791, 5.668032, 5.881447, 3.783429, 2.687109, 2.315882, 
    2.185626, 2.24172, 2.680243, 4.273811, 4.647846, 4.202462, 3.488654, 
    2.471768, 1.955085, 1.57258, 1.38111, 1.058366, 0.8350188, 0.6911973, 
    0.5835425, 0.6153647, 0.9760028, 6.609177, 5.571939, 3.501674, 2.606929, 
    2.291466,
  3.229089, 6.935664, 8.692479, 4.677368, 3.598944, 2.510919, 2.451262, 
    2.200563, 2.161129, 3.572072, 5.584081, 5.514449, 3.062308, 2.374481, 
    1.90406, 1.298325, 1.026381, 0.8172199, 0.6330573, 0.6665795, 0.7419336, 
    0.7689735, 1.207175, 4.287922, 9.533909, 7.635406, 4.386235, 3.095783, 
    3.015401,
  3.845778, 9.325099, 10.20839, 5.122003, 2.472875, 1.820285, 1.493068, 
    1.683563, 1.826575, 2.979807, 2.87138, 3.043921, 2.060629, 1.015877, 
    0.8434327, 0.7725915, 0.6033076, 0.5055855, 0.4598607, 0.4900373, 
    0.7028252, 1.400812, 4.043551, 11.23519, 10.71771, 7.896157, 3.448293, 
    2.852141, 3.176109,
  9.970213, 17.99129, 16.11723, 4.412662, 2.503506, 2.162273, 2.208709, 
    2.358088, 4.362659, 6.440028, 3.023451, 1.577255, 0.7176328, 0.4961319, 
    0.4606664, 0.4878267, 0.4662515, 0.4531605, 0.4804461, 0.623791, 
    0.7757388, 1.341503, 5.339626, 11.61744, 8.860375, 4.547874, 3.83004, 
    4.128545, 6.221515,
  11.95541, 12.20622, 12.70474, 8.865808, 4.891988, 4.003232, 4.478158, 
    4.4366, 4.446417, 3.318624, 2.263559, 1.234122, 1.210522, 1.07163, 
    0.8924587, 0.9743537, 0.8727807, 0.9468053, 1.104576, 1.350846, 1.74009, 
    2.667631, 4.242493, 4.904932, 2.198063, 2.66173, 3.672089, 6.616161, 
    12.71546,
  7.150325, 4.782622, 4.641602, 9.062119, 6.255053, 6.350884, 6.862213, 
    7.088072, 8.778878, 5.346342, 3.663944, 2.945102, 2.483201, 2.394094, 
    2.091278, 2.008811, 1.624926, 1.455486, 1.542389, 1.816573, 3.198295, 
    4.07528, 2.612383, 2.065371, 1.944015, 2.207373, 3.059684, 4.620621, 
    6.291802,
  6.860375, 6.904902, 6.09432, 6.7796, 6.924997, 7.887481, 11.50296, 
    10.74448, 14.78378, 20.3221, 12.91362, 9.160332, 7.204391, 6.098732, 
    4.984911, 3.997507, 3.223883, 2.557182, 2.085058, 2.599135, 4.516323, 
    5.195385, 5.132148, 4.033928, 2.950478, 2.76137, 3.540268, 3.761225, 
    5.535153,
  5.697429, 6.926678, 7.524383, 10.19744, 13.72085, 10.46639, 15.43927, 
    17.57598, 15.61957, 13.56826, 12.03227, 10.34172, 9.176367, 8.056739, 
    7.27543, 5.933781, 4.747779, 3.979612, 3.510153, 3.620076, 6.26847, 
    8.807782, 7.442849, 7.210013, 7.043756, 5.256713, 4.53813, 4.028833, 
    4.463912,
  4.997267, 6.892731, 7.247006, 7.876278, 8.33227, 8.773682, 8.986202, 
    9.786572, 11.11594, 12.01056, 12.10947, 11.25714, 9.439803, 8.43446, 
    7.778152, 6.622134, 5.703778, 4.907228, 4.409136, 4.913193, 6.738947, 
    7.855064, 8.454815, 9.308414, 8.70905, 7.003919, 6.014705, 5.508895, 
    4.85407,
  5.337352, 6.085739, 6.567849, 6.896806, 7.49325, 8.02409, 8.282839, 
    8.18914, 8.907677, 9.451908, 10.29643, 9.502032, 8.641982, 7.720194, 
    6.911887, 5.646837, 5.140912, 5.112026, 5.189793, 5.450563, 5.717045, 
    6.234643, 6.816654, 7.309367, 7.950948, 7.157768, 6.084639, 5.410041, 
    5.244427,
  4.912149, 5.034848, 5.385629, 5.849466, 6.762688, 7.229373, 7.189726, 
    7.944107, 7.881991, 7.47157, 7.084521, 6.758114, 6.204467, 5.967085, 
    5.190553, 4.712497, 4.645119, 4.879609, 4.819138, 4.77465, 4.565045, 
    5.159358, 5.949068, 6.240205, 6.202334, 5.892982, 4.990414, 5.237037, 
    4.801768,
  4.750857, 4.712909, 4.95795, 5.059063, 5.204669, 5.349894, 5.683633, 
    5.739722, 5.442209, 5.212239, 5.099885, 4.805651, 4.613845, 4.256139, 
    4.077658, 4.103478, 4.092396, 3.991691, 4.012371, 4.202813, 4.521494, 
    4.640576, 4.610257, 4.773211, 4.944688, 4.62871, 4.852817, 5.187362, 
    4.882563,
  0.4701429, 0.4701429, 0.4701429, 0.4701429, 0.4701429, 0.4701429, 
    0.4701429, 0.4546457, 0.4546457, 0.4546457, 0.4546457, 0.4546457, 
    0.4546457, 0.4546457, 0.4475154, 0.4475154, 0.4475154, 0.4475154, 
    0.4475154, 0.4475154, 0.4475154, 0.4571896, 0.4571896, 0.4571896, 
    0.4571896, 0.4571896, 0.4571896, 0.4571896, 0.4701429,
  0.5956888, 0.5484015, 0.5510916, 0.5184789, 0.482812, 0.4532831, 0.4321057, 
    0.4305238, 0.4094226, 0.3864131, 0.3659011, 0.354658, 0.3530925, 
    0.2952034, 0.2970747, 0.3114329, 0.3173669, 0.3467844, 0.3962358, 
    0.4560918, 0.4966329, 0.5265206, 0.5038396, 0.4631799, 0.4413825, 
    0.4477241, 0.5007871, 0.5378469, 0.606131,
  0.7053797, 0.6345483, 0.6074054, 0.6041222, 0.7270469, 0.6088977, 
    0.4325436, 0.5028834, 0.4553429, 0.4308408, 0.4920548, 0.5520179, 
    0.4686647, 0.4785828, 0.5342003, 0.5517886, 0.5344107, 0.5134151, 
    0.4810885, 0.4911279, 0.5040948, 0.4845733, 0.5421852, 0.5378792, 
    0.6030593, 0.5819904, 0.6692412, 0.7736282, 0.7344127,
  1.062878, 1.05513, 0.9632644, 0.934586, 1.027145, 0.9818081, 0.8378844, 
    0.6981575, 0.5910777, 0.5589699, 0.6189047, 0.7929843, 0.8726746, 
    1.308652, 1.464077, 1.431921, 1.286762, 1.086379, 0.9410939, 0.8029114, 
    0.7061764, 0.6542692, 0.606802, 0.6590945, 0.8330588, 1.051971, 1.225605, 
    1.224162, 1.122183,
  1.637505, 1.363349, 1.285387, 1.406264, 1.560445, 1.425665, 1.252806, 
    1.116643, 0.919468, 0.7975431, 0.8541508, 1.258135, 1.93358, 2.1368, 
    2.315934, 1.984888, 1.698483, 1.463889, 1.269944, 1.104836, 0.9761624, 
    0.8881719, 0.8108233, 1.042963, 1.527508, 2.004451, 2.294399, 1.96322, 
    1.885126,
  1.80404, 1.748224, 1.928704, 2.946946, 2.41241, 1.899107, 1.65095, 
    1.489116, 1.372749, 1.425519, 1.845589, 2.502633, 3.624699, 3.21857, 
    2.683504, 2.095961, 1.95958, 1.712039, 1.506143, 1.292723, 1.11626, 
    0.9265925, 0.8525249, 1.067246, 4.572562, 3.282207, 2.607483, 2.188175, 
    1.89501,
  2.107682, 2.438157, 6.287644, 6.384747, 3.763681, 2.531372, 2.073868, 
    1.960256, 2.052777, 2.792968, 4.779352, 5.204113, 4.513092, 3.48143, 
    2.296779, 1.806834, 1.500005, 1.287027, 1.031337, 0.8098853, 0.6723121, 
    0.565439, 0.6046534, 1.066652, 8.046205, 5.86531, 3.372184, 2.467094, 
    2.082139,
  3.113277, 8.048187, 9.351204, 4.760139, 3.601596, 2.338313, 2.232194, 
    2.015479, 2.126734, 4.140311, 6.689522, 5.927656, 3.084347, 2.216486, 
    1.763039, 1.159872, 0.9740565, 0.7762674, 0.6053052, 0.6528698, 
    0.6907071, 0.6749169, 1.154361, 4.560845, 10.59395, 7.967447, 4.130775, 
    2.908453, 2.807692,
  3.865927, 10.38312, 11.06362, 5.455521, 2.297873, 1.643942, 1.394748, 
    1.574406, 1.738981, 2.961382, 3.016405, 3.144215, 2.075788, 0.9392934, 
    0.7877029, 0.6917009, 0.5307564, 0.4481342, 0.432064, 0.5094917, 
    0.7984048, 1.552154, 5.012625, 12.38429, 11.54307, 8.60876, 3.074782, 
    2.528205, 2.931493,
  11.4194, 20.11927, 20.14484, 4.870982, 2.561645, 2.063161, 2.165444, 
    2.368822, 4.323874, 6.545996, 3.056571, 1.61215, 0.7076194, 0.4511891, 
    0.4101168, 0.4322921, 0.4278562, 0.4584455, 0.4753375, 0.62747, 
    0.9462462, 1.857909, 7.602282, 14.28256, 10.25136, 4.391102, 3.65242, 
    4.24358, 7.061691,
  13.87983, 13.84706, 14.09029, 10.90089, 5.966056, 4.670347, 5.238585, 
    4.847765, 4.453434, 3.327308, 2.225811, 1.245978, 1.133366, 0.9739631, 
    0.848732, 0.9580318, 0.8928882, 0.9929243, 1.149253, 1.445588, 1.890644, 
    2.866281, 4.459517, 5.01139, 2.111351, 2.729615, 3.972674, 7.266627, 
    13.94797,
  11.30495, 7.332525, 5.997029, 11.2576, 8.036894, 7.36275, 7.34804, 
    7.857997, 9.258168, 5.675993, 3.74416, 2.883882, 2.437271, 2.266169, 
    2.002279, 1.950954, 1.632285, 1.464601, 1.61363, 1.99172, 3.854737, 
    4.612178, 2.574483, 2.055544, 1.954076, 2.382996, 3.617095, 6.354759, 
    9.878737,
  8.400747, 8.103613, 6.796443, 7.845151, 8.938452, 9.73966, 13.63844, 
    11.40135, 16.24377, 21.84986, 13.04812, 9.285231, 7.240181, 6.132908, 
    4.879573, 3.936721, 3.256997, 2.566872, 2.070807, 2.757964, 5.286711, 
    6.300892, 5.703923, 4.079363, 2.888106, 2.786741, 3.512953, 3.87518, 
    6.740642,
  6.227923, 7.653373, 7.985773, 10.70183, 15.41007, 11.20175, 16.71359, 
    18.75501, 16.67616, 13.87528, 12.31707, 10.51097, 9.172623, 7.881523, 
    7.179332, 5.86315, 4.669548, 3.880549, 3.409147, 3.670375, 7.64219, 
    10.30679, 8.355181, 7.889146, 7.584904, 5.394438, 4.590694, 4.011182, 
    4.551131,
  5.129541, 7.142658, 7.647384, 8.214486, 8.908013, 9.40918, 9.415922, 
    9.867907, 11.55805, 12.95381, 13.10506, 11.89025, 9.902048, 8.70397, 
    7.947688, 6.631365, 5.606316, 4.773583, 4.349093, 5.012165, 7.464257, 
    8.791923, 9.196247, 10.19762, 9.448124, 7.374822, 6.207623, 5.526105, 
    4.970896,
  5.563809, 6.331647, 6.934031, 7.154369, 7.815291, 8.533533, 8.841211, 
    8.755137, 9.581142, 10.20836, 10.68316, 9.800327, 9.10085, 8.051299, 
    7.12208, 5.907565, 5.274432, 5.280396, 5.534848, 6.018879, 6.091264, 
    6.825853, 7.117693, 7.735107, 8.538446, 7.571468, 6.326071, 5.676672, 
    5.451394,
  5.126826, 5.296717, 5.697796, 6.181815, 7.189644, 7.602102, 7.464055, 
    8.379527, 8.443116, 7.956149, 7.470895, 7.154884, 6.495406, 6.076582, 
    5.398449, 4.849318, 4.878601, 5.038345, 5.049038, 5.027531, 4.818123, 
    5.321466, 6.18013, 6.545447, 6.48594, 6.22573, 5.253746, 5.465328, 
    4.987709,
  4.906882, 4.924721, 5.145611, 5.190497, 5.342454, 5.479787, 5.773409, 
    5.808411, 5.54584, 5.349728, 5.275153, 4.901166, 4.619685, 4.218513, 
    4.085203, 4.124502, 4.168424, 4.092285, 4.186259, 4.389549, 4.714589, 
    4.844609, 4.862435, 5.026146, 5.194379, 4.903528, 5.095495, 5.410861, 
    5.075343,
  0.4624002, 0.4624002, 0.4624002, 0.4624002, 0.4624002, 0.4624002, 
    0.4624002, 0.4452349, 0.4452349, 0.4452349, 0.4452349, 0.4452349, 
    0.4452349, 0.4452349, 0.437698, 0.437698, 0.437698, 0.437698, 0.437698, 
    0.437698, 0.437698, 0.4496841, 0.4496841, 0.4496841, 0.4496841, 
    0.4496841, 0.4496841, 0.4496841, 0.4624002,
  0.5916227, 0.5404015, 0.5327395, 0.4971243, 0.4589729, 0.4315211, 
    0.4127818, 0.4149648, 0.3994959, 0.3697396, 0.3438162, 0.3321577, 
    0.3353345, 0.2725757, 0.2756262, 0.2888737, 0.2934314, 0.3231712, 
    0.3687652, 0.4242347, 0.466236, 0.5053199, 0.4934034, 0.4567261, 
    0.4285967, 0.4398009, 0.4784552, 0.517907, 0.5977955,
  0.6517928, 0.5762699, 0.5440626, 0.5440261, 0.6768216, 0.5578752, 
    0.3842749, 0.4630009, 0.428542, 0.3996451, 0.4536674, 0.5161039, 
    0.4200688, 0.4265473, 0.4916784, 0.5061912, 0.4942218, 0.4590805, 
    0.4362568, 0.4429527, 0.466148, 0.452627, 0.5121806, 0.5308632, 
    0.6011995, 0.5742938, 0.6696076, 0.7611471, 0.7154054,
  1.040124, 1.007937, 0.9197407, 0.8744001, 0.9702973, 0.9200051, 0.7592578, 
    0.6273224, 0.5366974, 0.5065145, 0.5683582, 0.7335579, 0.8161682, 
    1.228109, 1.366664, 1.36009, 1.200966, 1.023223, 0.8626369, 0.7357532, 
    0.6566684, 0.613382, 0.5760543, 0.6154496, 0.834422, 1.102652, 1.256472, 
    1.240267, 1.105241,
  1.60506, 1.324624, 1.23403, 1.356315, 1.516955, 1.320186, 1.163215, 
    1.037273, 0.8406984, 0.7206826, 0.8015146, 1.218375, 1.891574, 2.028913, 
    2.232598, 1.906708, 1.584886, 1.345813, 1.148475, 0.9940926, 0.8793698, 
    0.8115214, 0.7349057, 1.013811, 1.631233, 2.188818, 2.35984, 1.998944, 
    1.852864,
  1.768097, 1.66629, 1.896604, 2.993496, 2.361101, 1.787873, 1.498737, 
    1.322213, 1.234589, 1.285885, 1.914577, 2.598986, 3.867998, 3.313483, 
    2.641445, 2.023404, 1.814982, 1.578927, 1.391049, 1.203642, 1.050676, 
    0.8673468, 0.8101098, 1.112937, 5.667129, 3.588114, 2.598687, 2.150591, 
    1.856568,
  1.930264, 2.405465, 7.28675, 7.120999, 3.821578, 2.4091, 1.915058, 1.72718, 
    1.84744, 3.068293, 5.544339, 6.030789, 5.103065, 3.529309, 2.201624, 
    1.632019, 1.403875, 1.180016, 1.007986, 0.8018784, 0.6643071, 0.565964, 
    0.5820554, 1.189831, 9.777843, 6.243383, 3.373648, 2.321715, 1.925279,
  3.226805, 9.787778, 10.63476, 5.068829, 3.765332, 2.213133, 2.077407, 
    1.89415, 2.281047, 5.172571, 7.927574, 6.548211, 3.229831, 2.090186, 
    1.629005, 1.048584, 0.9156335, 0.7531437, 0.6019952, 0.6029799, 
    0.6009053, 0.5986255, 1.072774, 4.888038, 11.80882, 8.590609, 3.973235, 
    2.729911, 2.63296,
  4.413432, 11.85816, 12.71018, 6.304842, 2.279923, 1.560839, 1.335147, 
    1.512423, 1.726994, 3.067213, 3.265049, 3.259016, 2.083215, 0.8865041, 
    0.726999, 0.5917908, 0.4655861, 0.4025045, 0.4196553, 0.5355863, 
    0.983484, 2.038871, 6.241687, 13.65402, 12.95865, 9.877392, 2.822198, 
    2.267966, 2.816936,
  12.80252, 21.83756, 23.20349, 5.980819, 3.1944, 2.124445, 2.162088, 
    2.379162, 4.447754, 6.778306, 3.119851, 1.655756, 0.70601, 0.4027702, 
    0.3646648, 0.3950492, 0.402182, 0.4512085, 0.5350618, 0.7624429, 
    1.236785, 2.992831, 10.4378, 16.52997, 11.3818, 4.141182, 3.548111, 
    4.577754, 8.101978,
  17.058, 17.31019, 16.6732, 13.11549, 7.142301, 5.55338, 6.394532, 5.48725, 
    4.659091, 3.388567, 2.228456, 1.259764, 1.078471, 0.892837, 0.8224974, 
    0.8825838, 0.915468, 1.012028, 1.208353, 1.559325, 2.101616, 3.249599, 
    4.855618, 5.346242, 2.182217, 3.020182, 4.581854, 8.486543, 15.71847,
  14.99583, 10.89593, 8.058225, 12.74059, 10.55619, 8.466098, 8.304778, 
    9.435631, 10.55512, 6.520323, 4.026339, 2.950972, 2.391332, 2.162009, 
    1.98381, 1.916086, 1.639865, 1.493891, 1.664654, 2.243984, 4.67563, 
    5.466245, 2.619794, 2.111238, 2.052459, 2.727318, 4.383609, 8.546917, 
    14.25891,
  10.15819, 9.641564, 7.752529, 9.834396, 11.57439, 12.08191, 16.66179, 
    12.33984, 18.19749, 23.11175, 12.98223, 9.238428, 7.183553, 6.08777, 
    4.815933, 3.968947, 3.240691, 2.550654, 2.10729, 2.955164, 6.559279, 
    7.822598, 6.387854, 4.24331, 2.933059, 2.913923, 3.552463, 4.009573, 
    7.756227,
  6.919485, 8.519901, 8.759501, 11.64122, 17.27908, 12.3975, 18.27708, 
    20.37328, 18.47881, 14.5674, 12.90591, 10.89921, 9.171683, 7.763893, 
    7.065827, 5.710721, 4.566527, 3.760067, 3.312473, 3.805754, 9.051415, 
    12.25517, 9.595218, 8.824876, 8.237609, 5.537519, 4.616716, 4.039116, 
    4.662199,
  5.326802, 7.537976, 8.229177, 8.814363, 9.895346, 10.37621, 10.06902, 
    10.14024, 12.26434, 14.16477, 14.2836, 12.67757, 10.58821, 9.032092, 
    8.199387, 6.696608, 5.558185, 4.675203, 4.312757, 5.171713, 8.61058, 
    10.01549, 10.29947, 11.0917, 10.32584, 7.863651, 6.486604, 5.645687, 
    5.092402,
  5.802347, 6.71782, 7.476941, 7.640175, 8.360193, 9.286669, 9.667616, 
    9.549946, 10.4253, 11.00003, 11.17678, 10.14308, 9.683762, 8.559908, 
    7.409244, 6.229319, 5.491794, 5.516637, 5.862614, 6.751841, 6.691554, 
    7.285195, 7.414052, 8.193321, 9.229856, 8.04395, 6.611866, 5.989978, 
    5.6565,
  5.346149, 5.58987, 6.077709, 6.581929, 7.707396, 8.003898, 7.88852, 
    8.958186, 9.106751, 8.422766, 7.931642, 7.727235, 6.794705, 6.252047, 
    5.655162, 5.1271, 5.122802, 5.342957, 5.481985, 5.413838, 5.212253, 
    5.484962, 6.430934, 6.864584, 6.73436, 6.524844, 5.466056, 5.703238, 
    5.166464,
  5.086865, 5.14332, 5.331967, 5.383984, 5.464365, 5.607613, 5.847682, 
    5.962524, 5.793573, 5.605757, 5.5207, 5.045899, 4.710403, 4.267448, 
    4.143627, 4.208972, 4.313951, 4.317655, 4.475384, 4.606941, 4.944644, 
    5.111042, 5.107057, 5.258941, 5.421364, 5.16503, 5.323988, 5.611199, 
    5.305443,
  0.451346, 0.451346, 0.451346, 0.451346, 0.451346, 0.451346, 0.451346, 
    0.4367347, 0.4367347, 0.4367347, 0.4367347, 0.4367347, 0.4367347, 
    0.4367347, 0.4305194, 0.4305194, 0.4305194, 0.4305194, 0.4305194, 
    0.4305194, 0.4305194, 0.4410538, 0.4410538, 0.4410538, 0.4410538, 
    0.4410538, 0.4410538, 0.4410538, 0.451346,
  0.5824398, 0.5350035, 0.5136908, 0.4747666, 0.4374119, 0.4130905, 
    0.3954117, 0.3983375, 0.3851147, 0.3515047, 0.3235184, 0.3098942, 
    0.3148716, 0.25159, 0.25514, 0.2693411, 0.271569, 0.3049405, 0.3476985, 
    0.4050386, 0.4506928, 0.49021, 0.4888118, 0.4473209, 0.4134157, 
    0.4315788, 0.4548221, 0.4984963, 0.5846022,
  0.5970496, 0.5182862, 0.4876779, 0.4791762, 0.6209737, 0.5047344, 
    0.3398415, 0.4255048, 0.4010514, 0.3692787, 0.4175673, 0.4765156, 
    0.37904, 0.3795522, 0.449629, 0.4683729, 0.4516884, 0.408477, 0.3954249, 
    0.4013171, 0.4236645, 0.426285, 0.4866972, 0.534918, 0.6238849, 
    0.5840278, 0.6681376, 0.7377946, 0.6936148,
  1.01055, 0.9574805, 0.8811499, 0.8196341, 0.9206149, 0.8594863, 0.6774209, 
    0.5552934, 0.4841056, 0.4558596, 0.5132374, 0.6751363, 0.7645391, 
    1.155206, 1.291285, 1.285722, 1.136246, 0.9637365, 0.7987367, 0.6701922, 
    0.6031795, 0.5749026, 0.5479708, 0.5816077, 0.8528078, 1.174143, 1.29469, 
    1.277269, 1.090259,
  1.556278, 1.265596, 1.200912, 1.322619, 1.470796, 1.226132, 1.089903, 
    0.9553205, 0.7667684, 0.6499918, 0.7402874, 1.188329, 1.892991, 1.996459, 
    2.175918, 1.839399, 1.502465, 1.254876, 1.045976, 0.8875115, 0.7972894, 
    0.7382154, 0.6718228, 0.99623, 1.871479, 2.443033, 2.441632, 2.032391, 
    1.812587,
  1.767963, 1.604054, 1.939807, 3.029856, 2.315005, 1.702929, 1.377068, 
    1.187709, 1.125487, 1.176179, 1.969136, 2.742353, 4.172366, 3.421483, 
    2.670542, 1.968685, 1.668891, 1.43987, 1.28022, 1.10409, 0.9706365, 
    0.7935506, 0.7568683, 1.231354, 6.893758, 3.940375, 2.700536, 2.147651, 
    1.841159,
  1.800554, 2.431879, 8.877794, 7.996663, 3.925864, 2.248578, 1.761651, 
    1.48859, 1.590895, 3.550444, 6.743558, 7.103293, 5.902477, 3.600853, 
    2.180692, 1.479418, 1.288738, 1.106463, 0.9754059, 0.801811, 0.648765, 
    0.577055, 0.5586284, 1.460462, 11.68125, 6.683449, 3.343956, 2.163851, 
    1.764298,
  3.331789, 11.61518, 12.63348, 5.665513, 4.029926, 2.042739, 1.945193, 
    1.870672, 2.656666, 6.533904, 9.302517, 7.713196, 3.676484, 2.045747, 
    1.502575, 0.9396812, 0.8292888, 0.7102705, 0.5998582, 0.5403364, 
    0.5445622, 0.5741043, 0.9632423, 5.20147, 13.39724, 9.332829, 4.005694, 
    2.429095, 2.553965,
  5.438422, 13.21532, 15.08559, 7.356643, 2.437172, 1.55933, 1.272708, 
    1.554152, 1.823468, 3.335385, 3.591802, 3.496246, 2.094604, 0.8274553, 
    0.6515307, 0.5083033, 0.4118938, 0.3798099, 0.4311622, 0.6238425, 
    1.24596, 2.919067, 7.524773, 15.08419, 14.76716, 11.54383, 2.738299, 
    2.197232, 2.968011,
  14.22311, 23.28401, 26.16696, 7.586555, 4.073416, 2.432401, 2.264666, 
    2.440093, 4.620504, 6.979315, 3.186055, 1.669285, 0.7127353, 0.3622388, 
    0.3259624, 0.3631818, 0.3953853, 0.4575067, 0.6469631, 1.0303, 1.801014, 
    4.741917, 13.50981, 18.01855, 12.15101, 4.036486, 3.474198, 5.117366, 
    9.217412,
  21.78315, 21.67299, 20.73214, 16.38229, 8.483586, 6.300307, 7.675487, 
    6.123244, 4.962618, 3.531293, 2.288504, 1.269641, 1.005097, 0.8543066, 
    0.764949, 0.8301962, 0.9026479, 1.013751, 1.319277, 1.715595, 2.408211, 
    3.688126, 5.41809, 5.973471, 2.493552, 3.589686, 5.68934, 10.43436, 
    18.9831,
  18.26987, 14.29922, 10.4152, 14.02755, 14.15294, 9.639691, 9.94147, 
    11.21423, 12.02019, 8.002055, 4.653684, 3.081103, 2.339934, 2.126374, 
    2.018506, 1.907096, 1.640052, 1.568655, 1.729234, 2.529426, 5.357135, 
    6.61233, 2.829232, 2.222178, 2.274675, 3.088141, 5.095322, 10.31442, 
    17.89417,
  12.33608, 11.47495, 8.737199, 12.80639, 14.55374, 14.91878, 20.09799, 
    13.79796, 20.76078, 23.86816, 12.66727, 9.017179, 6.960065, 5.78362, 
    4.765389, 4.047113, 3.263402, 2.545893, 2.145895, 3.129833, 8.182165, 
    9.498415, 7.170514, 4.506149, 3.042848, 3.076387, 3.701763, 4.227725, 
    8.92642,
  7.769128, 9.551853, 10.01596, 13.0513, 19.40941, 14.07703, 20.13997, 
    22.52666, 20.85583, 15.928, 14.00372, 11.50684, 9.32136, 7.746559, 
    6.870029, 5.57952, 4.481078, 3.68614, 3.225091, 4.042217, 10.62131, 
    14.70319, 11.07305, 10.02517, 9.218491, 5.758546, 4.653192, 4.180757, 
    4.876216,
  5.548027, 8.134175, 9.092886, 9.873658, 11.30602, 11.8193, 11.14425, 
    10.72718, 13.31118, 15.67616, 15.67427, 13.76868, 11.44415, 9.398313, 
    8.489855, 6.75361, 5.550845, 4.655154, 4.344064, 5.432002, 10.16756, 
    11.42927, 11.81848, 12.21381, 11.58465, 8.498548, 6.831647, 5.838451, 
    5.2379,
  6.157255, 7.32024, 8.1439, 8.426832, 9.255305, 10.28438, 10.77367, 
    10.63376, 11.62852, 12.04932, 12.03087, 10.66031, 10.26256, 9.157948, 
    7.834682, 6.631379, 5.691432, 5.801872, 6.237241, 7.628523, 7.503917, 
    7.811526, 7.826264, 8.736453, 9.964214, 8.598936, 6.926527, 6.31541, 
    5.918281,
  5.549238, 5.857417, 6.567544, 7.130415, 8.224169, 8.578524, 8.45637, 
    9.690554, 10.01187, 9.100336, 8.588367, 8.402626, 7.146683, 6.562562, 
    5.943521, 5.528489, 5.543434, 5.940884, 6.087148, 6.024064, 5.732368, 
    5.766533, 6.746162, 7.225163, 6.906954, 6.773511, 5.660417, 5.943815, 
    5.377168,
  5.358007, 5.337006, 5.550879, 5.628303, 5.665667, 5.853649, 6.003175, 
    6.288025, 6.227993, 5.986862, 5.823874, 5.322997, 4.921649, 4.50031, 
    4.345295, 4.450387, 4.578039, 4.564325, 4.785871, 4.851815, 5.167104, 
    5.423248, 5.385011, 5.509605, 5.679025, 5.419927, 5.516806, 5.808101, 
    5.58885,
  0.4358947, 0.4358947, 0.4358947, 0.4358947, 0.4358947, 0.4358947, 
    0.4358947, 0.425301, 0.425301, 0.425301, 0.425301, 0.425301, 0.425301, 
    0.425301, 0.4196342, 0.4196342, 0.4196342, 0.4196342, 0.4196342, 
    0.4196342, 0.4196342, 0.4272296, 0.4272296, 0.4272296, 0.4272296, 
    0.4272296, 0.4272296, 0.4272296, 0.4358947,
  0.5679162, 0.5242132, 0.4923705, 0.4501529, 0.4167866, 0.394699, 0.3778263, 
    0.380694, 0.3691618, 0.3348803, 0.3076506, 0.2906272, 0.2933211, 
    0.2332091, 0.2341187, 0.2481695, 0.249977, 0.2872441, 0.3319535, 
    0.3932292, 0.4469927, 0.4867839, 0.4856478, 0.4319811, 0.3945945, 
    0.4187384, 0.4267497, 0.4760024, 0.5671196,
  0.548016, 0.4615656, 0.4359372, 0.423144, 0.5594721, 0.4544999, 0.2992813, 
    0.3919177, 0.3701527, 0.3389463, 0.3819226, 0.4346829, 0.3471251, 
    0.3371594, 0.4065259, 0.4350031, 0.4109015, 0.3686892, 0.3613628, 
    0.3655099, 0.3833121, 0.4070507, 0.4709401, 0.5556257, 0.6572634, 
    0.6023238, 0.6564503, 0.7110897, 0.6656269,
  0.9797213, 0.9042049, 0.8378265, 0.7732363, 0.8673433, 0.7949903, 
    0.5991827, 0.4929464, 0.4329801, 0.4078189, 0.4613339, 0.6233557, 
    0.7310115, 1.111387, 1.250603, 1.234716, 1.085821, 0.9176126, 0.7480108, 
    0.6147617, 0.5568451, 0.5349697, 0.5138327, 0.5499228, 0.8931623, 
    1.271288, 1.320121, 1.313554, 1.079832,
  1.518647, 1.212017, 1.173633, 1.292396, 1.39898, 1.149732, 1.01528, 
    0.8633543, 0.6917054, 0.5774091, 0.6716855, 1.176074, 1.925766, 2.034662, 
    2.16373, 1.803826, 1.448174, 1.199272, 0.9693457, 0.815892, 0.7361432, 
    0.6664833, 0.6078326, 0.9981647, 2.314858, 2.75111, 2.592313, 2.092617, 
    1.76481,
  1.76787, 1.569864, 2.083663, 2.993639, 2.234186, 1.621174, 1.260165, 
    1.085423, 1.038494, 1.085996, 2.052678, 2.992865, 4.574361, 3.555346, 
    2.74921, 1.916507, 1.523077, 1.315073, 1.169164, 1.009769, 0.8816013, 
    0.7232485, 0.6906739, 1.44236, 8.110701, 4.377808, 2.82506, 2.161172, 
    1.836429,
  1.699131, 2.510351, 10.81791, 8.714327, 4.003167, 2.10424, 1.586639, 
    1.321963, 1.3631, 4.249129, 8.384107, 8.455672, 7.013856, 3.713501, 
    2.147385, 1.366302, 1.185927, 1.04955, 0.9222192, 0.7831492, 0.6145347, 
    0.5546859, 0.5455486, 1.906085, 13.69024, 7.194295, 3.292135, 1.981107, 
    1.647715,
  3.348774, 12.91891, 15.35188, 6.541142, 4.299269, 1.792647, 1.788004, 
    1.970956, 3.237712, 8.063038, 10.86353, 9.051821, 4.279092, 2.025417, 
    1.387317, 0.8417231, 0.7473997, 0.6570203, 0.5605636, 0.5034658, 
    0.5028096, 0.5292925, 0.909077, 5.367623, 15.51129, 10.38143, 3.993028, 
    2.166454, 2.45744,
  6.189981, 14.45802, 17.53058, 8.37707, 2.615448, 1.604138, 1.268304, 
    1.692116, 2.231356, 3.7494, 4.108293, 3.785942, 2.048471, 0.7426739, 
    0.5683149, 0.4504681, 0.3755476, 0.3882626, 0.4502722, 0.7962368, 
    1.640427, 3.570346, 8.642427, 16.66494, 16.39437, 12.88259, 2.62368, 
    2.233337, 3.279345,
  16.33678, 25.18219, 29.63402, 9.411866, 4.528722, 2.914058, 2.488789, 
    2.556926, 4.98568, 7.327482, 3.296968, 1.665466, 0.703796, 0.3291797, 
    0.305857, 0.3482704, 0.4000502, 0.524949, 0.825977, 1.41601, 2.635056, 
    6.707944, 15.80744, 19.3808, 13.60258, 4.357512, 3.665858, 5.918939, 
    10.88985,
  27.19468, 26.23141, 25.44278, 20.78083, 9.892333, 7.003456, 8.991758, 
    6.789603, 5.4419, 3.800001, 2.428736, 1.266246, 0.9119282, 0.7913114, 
    0.702085, 0.8131666, 0.8609134, 1.051966, 1.447266, 1.924724, 2.735627, 
    4.093091, 6.06867, 7.177538, 2.958255, 4.273289, 6.755916, 12.96545, 
    24.05312,
  20.90603, 16.97063, 12.47017, 15.45539, 18.01613, 10.85831, 12.15796, 
    12.99744, 13.48569, 10.03508, 5.613178, 3.279452, 2.350514, 2.152135, 
    2.123128, 1.963966, 1.710938, 1.643078, 1.795567, 2.734874, 6.079481, 
    7.988503, 3.198856, 2.528643, 2.540114, 3.47806, 5.489031, 11.31986, 
    20.84707,
  14.816, 13.27868, 9.652834, 16.09866, 17.64888, 17.72506, 23.53819, 
    15.59728, 23.74015, 24.30829, 12.38861, 8.73129, 6.74346, 5.461854, 
    4.725815, 4.059887, 3.294986, 2.588794, 2.177952, 3.163368, 9.739305, 
    11.29483, 7.970821, 4.871917, 3.215938, 3.232113, 3.854973, 4.399936, 
    10.45571,
  8.893478, 10.7426, 11.63691, 14.97979, 21.64458, 16.3511, 22.21222, 
    24.94281, 23.55835, 17.7899, 15.59729, 12.62709, 9.734243, 7.792697, 
    6.748586, 5.467974, 4.370008, 3.639451, 3.173863, 4.440567, 12.19221, 
    17.43212, 12.8341, 11.63825, 10.35141, 6.085016, 4.837386, 4.418691, 
    5.213048,
  5.899294, 9.012465, 10.4865, 11.3899, 12.98448, 13.63316, 12.72928, 
    11.58388, 14.68194, 17.65341, 17.63304, 15.36346, 12.39543, 10.01687, 
    8.790191, 6.83924, 5.607498, 4.722045, 4.551342, 5.915898, 12.3333, 
    13.37886, 13.95274, 14.06925, 13.11267, 9.342188, 7.220758, 6.072921, 
    5.434815,
  6.621116, 8.266451, 9.138803, 9.647646, 10.51258, 11.69249, 12.11886, 
    12.03294, 13.18249, 13.47752, 13.19125, 11.50657, 10.94194, 9.916891, 
    8.43583, 7.116991, 5.964849, 6.213969, 6.821498, 8.797099, 8.564277, 
    8.527749, 8.669906, 9.488973, 10.78548, 9.25677, 7.265464, 6.666012, 
    6.240058,
  5.76955, 6.391928, 7.213963, 7.9422, 8.951514, 9.273523, 9.246046, 10.7833, 
    11.21265, 10.15879, 9.583359, 9.160455, 7.571375, 6.984632, 6.341609, 
    6.040227, 6.18956, 6.780756, 6.886989, 6.956432, 6.357924, 6.18363, 
    7.156218, 7.589108, 7.027019, 6.979954, 5.809107, 6.192932, 5.670504,
  5.698559, 5.631623, 5.83375, 5.945838, 5.971449, 6.130066, 6.299925, 
    6.787864, 6.774674, 6.458154, 6.114198, 5.661951, 5.221375, 4.788865, 
    4.656479, 4.788943, 4.922543, 4.800202, 5.050928, 5.132619, 5.384148, 
    5.771595, 5.699323, 5.796262, 5.966484, 5.641517, 5.69698, 6.029144, 
    5.920204,
  0.4166179, 0.4166179, 0.4166179, 0.4166179, 0.4166179, 0.4166179, 
    0.4166179, 0.4097569, 0.4097569, 0.4097569, 0.4097569, 0.4097569, 
    0.4097569, 0.4097569, 0.4049671, 0.4049671, 0.4049671, 0.4049671, 
    0.4049671, 0.4049671, 0.4049671, 0.4101444, 0.4101444, 0.4101444, 
    0.4101444, 0.4101444, 0.4101444, 0.4101444, 0.4166179,
  0.5459655, 0.50828, 0.4693711, 0.4276339, 0.3977624, 0.3763118, 0.3609525, 
    0.3627824, 0.3525517, 0.3226024, 0.295343, 0.274554, 0.2738228, 
    0.2184681, 0.2118576, 0.2230559, 0.2279535, 0.2683477, 0.3179883, 
    0.384056, 0.44786, 0.4935638, 0.4789385, 0.4017712, 0.3697931, 0.3956556, 
    0.3949775, 0.4532108, 0.5433988,
  0.4967556, 0.4012423, 0.3867158, 0.3734257, 0.4993106, 0.4087584, 
    0.2617079, 0.3600565, 0.3377901, 0.309857, 0.349809, 0.3938909, 
    0.3194448, 0.2983631, 0.3650002, 0.3978465, 0.3733271, 0.3373878, 
    0.3281804, 0.33208, 0.3445616, 0.3843179, 0.4513492, 0.5894531, 
    0.6889845, 0.6240081, 0.646242, 0.6775681, 0.6236776,
  0.9516318, 0.8463782, 0.7922491, 0.7250971, 0.7994333, 0.7233214, 
    0.5402145, 0.444764, 0.3863063, 0.3622055, 0.412182, 0.5700831, 0.712517, 
    1.085739, 1.215362, 1.210212, 1.044985, 0.8746638, 0.6997955, 0.561906, 
    0.5090421, 0.49041, 0.4842297, 0.5312627, 0.9851831, 1.386871, 1.36255, 
    1.343529, 1.071388,
  1.472682, 1.172174, 1.138674, 1.258197, 1.321489, 1.086678, 0.9442028, 
    0.7724361, 0.6172161, 0.5129119, 0.6173164, 1.167954, 1.967833, 2.10555, 
    2.191129, 1.766315, 1.428306, 1.139724, 0.9061093, 0.7612193, 0.690225, 
    0.5985795, 0.5409251, 1.045053, 2.914635, 3.063237, 2.757539, 2.194715, 
    1.721117,
  1.747955, 1.525525, 2.230056, 2.970075, 2.150227, 1.521588, 1.144392, 
    0.9887909, 0.9413978, 1.025838, 2.122648, 3.282521, 5.0943, 3.758229, 
    2.905178, 1.896119, 1.383101, 1.200288, 1.062046, 0.9262103, 0.7865921, 
    0.6536888, 0.6246104, 1.764709, 9.308714, 4.946274, 2.925145, 2.152864, 
    1.807349,
  1.570593, 2.754818, 13.03673, 9.038671, 3.887248, 1.955361, 1.456943, 
    1.205147, 1.211645, 5.093325, 10.49268, 10.42791, 8.695949, 3.894077, 
    2.112214, 1.305875, 1.075771, 0.9693597, 0.852412, 0.7420676, 0.5717399, 
    0.5256632, 0.5688775, 2.466982, 16.18695, 7.932586, 3.269265, 1.869725, 
    1.545737,
  3.087049, 13.85117, 18.66929, 7.45621, 4.393618, 1.576073, 1.637332, 
    2.075229, 3.984499, 9.557726, 12.79992, 10.50575, 4.765865, 1.99597, 
    1.29196, 0.7563674, 0.6690779, 0.6088809, 0.5119306, 0.4913347, 
    0.4733295, 0.4844804, 0.7309616, 5.264712, 18.55502, 11.94369, 3.866538, 
    1.963731, 2.244555,
  6.486495, 15.88671, 20.02899, 9.864411, 2.732609, 1.556341, 1.313843, 
    2.013619, 2.911863, 4.390479, 4.846753, 4.061052, 2.021187, 0.6623769, 
    0.4929135, 0.4119643, 0.3709454, 0.4100387, 0.5145882, 1.010378, 
    1.961934, 3.868259, 8.954192, 18.8688, 18.2086, 14.13155, 2.582016, 
    2.239128, 3.448294,
  18.55313, 27.66367, 33.14874, 11.69285, 4.261321, 3.34238, 2.77381, 
    2.730955, 5.597005, 8.15209, 3.462143, 1.660895, 0.6755562, 0.3140482, 
    0.3072482, 0.3554951, 0.4391407, 0.6705457, 1.107833, 1.841365, 3.759047, 
    8.325026, 16.87226, 21.59865, 16.04328, 5.276202, 4.263714, 7.044237, 
    12.95565,
  32.94396, 31.55514, 29.54766, 24.70829, 11.26261, 7.393108, 10.55625, 
    7.521313, 6.198825, 4.229774, 2.679662, 1.27449, 0.8497245, 0.7223225, 
    0.6769799, 0.7716317, 0.8516838, 1.129224, 1.591709, 2.182555, 3.096873, 
    4.647758, 6.664256, 9.094699, 3.536052, 4.875781, 7.578901, 16.34034, 
    29.36752,
  22.59902, 19.50767, 14.48371, 17.43702, 22.09319, 12.25205, 14.89789, 
    15.21719, 15.46114, 12.19518, 6.615448, 3.569398, 2.452151, 2.257064, 
    2.186954, 1.980266, 1.786648, 1.665912, 1.837109, 2.909427, 6.793462, 
    9.51389, 3.780646, 3.033378, 2.746857, 3.847458, 5.719432, 11.9394, 
    22.4092,
  17.71485, 15.17947, 11.07892, 19.11688, 20.55006, 20.7277, 26.70213, 
    17.87568, 26.71705, 25.25847, 12.39815, 8.513455, 6.5817, 5.286972, 
    4.657183, 4.036975, 3.275047, 2.608584, 2.20039, 3.269826, 11.40179, 
    13.52736, 8.869132, 5.456437, 3.555881, 3.407375, 3.942204, 4.503122, 
    12.13377,
  10.36655, 12.02652, 13.83868, 17.38434, 24.36572, 19.17305, 24.49299, 
    27.62355, 26.60412, 19.87347, 17.82393, 14.44235, 10.37558, 7.882327, 
    6.737809, 5.380264, 4.284236, 3.616774, 3.168678, 5.150203, 13.76589, 
    20.46184, 15.12626, 13.8628, 11.57482, 6.649402, 5.177838, 4.721129, 
    5.749597,
  6.41687, 10.18778, 12.47568, 13.55468, 15.00503, 15.82481, 14.69722, 
    12.79211, 16.46929, 20.05522, 20.5317, 17.57003, 13.65501, 10.81192, 
    9.188501, 7.057305, 5.728103, 4.886877, 4.860539, 6.726265, 15.15304, 
    16.00106, 16.9236, 16.6717, 14.6948, 10.45194, 7.672951, 6.354183, 
    5.717163,
  7.247363, 9.584314, 10.3647, 11.16439, 12.18987, 13.48093, 13.89991, 
    14.07224, 15.12078, 15.47609, 14.73646, 12.67787, 11.83443, 10.902, 
    9.228724, 7.699266, 6.41814, 6.783576, 7.599793, 10.40617, 10.05883, 
    9.706105, 9.676588, 10.49775, 11.68628, 9.993281, 7.643715, 7.010314, 
    6.657457,
  6.139805, 6.996356, 8.072253, 8.941816, 9.676435, 10.0232, 10.07075, 
    11.76521, 12.54764, 11.52922, 10.74453, 10.0682, 8.123332, 7.663199, 
    6.996635, 6.561936, 6.971022, 7.917682, 7.99092, 8.238003, 7.130014, 
    6.750913, 7.539842, 8.017225, 7.209888, 7.142438, 5.915145, 6.407007, 
    6.061738,
  6.12454, 6.047068, 6.182497, 6.29401, 6.319715, 6.435412, 6.630904, 
    7.258207, 7.334367, 6.950861, 6.445329, 6.111039, 5.699679, 5.268013, 
    5.118411, 5.22852, 5.328337, 5.101885, 5.269715, 5.424399, 5.706299, 
    6.166396, 6.021245, 6.074375, 6.246861, 5.87112, 5.877216, 6.273757, 
    6.299896,
  0.3984487, 0.3984487, 0.3984487, 0.3984487, 0.3984487, 0.3984487, 
    0.3984487, 0.3953831, 0.3953831, 0.3953831, 0.3953831, 0.3953831, 
    0.3953831, 0.3953831, 0.3905486, 0.3905486, 0.3905486, 0.3905486, 
    0.3905486, 0.3905486, 0.3905486, 0.3953913, 0.3953913, 0.3953913, 
    0.3953913, 0.3953913, 0.3953913, 0.3953913, 0.3984487,
  0.5189677, 0.4884913, 0.4456709, 0.4046678, 0.3787532, 0.3576576, 
    0.3444825, 0.3438349, 0.3359609, 0.312745, 0.2861753, 0.2609253, 
    0.2581998, 0.2060002, 0.1915273, 0.1970449, 0.2068111, 0.249108, 
    0.305742, 0.3746728, 0.4506423, 0.4996994, 0.4640829, 0.3547262, 
    0.3395817, 0.3649687, 0.3654601, 0.4325094, 0.5163417,
  0.4490467, 0.3511694, 0.3401512, 0.3269494, 0.4464947, 0.3683173, 
    0.2291292, 0.3316873, 0.3057992, 0.2852812, 0.3222626, 0.3591835, 
    0.2959625, 0.2651512, 0.3220802, 0.354838, 0.3374757, 0.3104728, 
    0.3045842, 0.3061137, 0.3150878, 0.3623935, 0.4232379, 0.6104817, 
    0.7057668, 0.6476635, 0.6325027, 0.6428606, 0.5837346,
  0.9187388, 0.7986272, 0.7409952, 0.6786226, 0.7367496, 0.6501337, 
    0.4933361, 0.4007474, 0.3473609, 0.3236271, 0.3652508, 0.5195596, 
    0.6959615, 1.063701, 1.168242, 1.171892, 0.9934644, 0.8385313, 0.6529037, 
    0.5195855, 0.4696202, 0.4515614, 0.4559641, 0.5355984, 1.129741, 
    1.501727, 1.406533, 1.356585, 1.046903,
  1.404467, 1.147799, 1.103192, 1.225191, 1.238539, 1.022431, 0.8752776, 
    0.6850072, 0.5481699, 0.4591984, 0.5685517, 1.152298, 2.042789, 2.161381, 
    2.260214, 1.755583, 1.410032, 1.087996, 0.8596646, 0.7056993, 0.6436523, 
    0.5359183, 0.4845163, 1.176566, 3.657925, 3.336178, 2.893562, 2.2614, 
    1.671463,
  1.673478, 1.47626, 2.29551, 2.894436, 2.060799, 1.398891, 1.036147, 
    0.903049, 0.8380703, 0.9587979, 2.102872, 3.48474, 5.797407, 3.959264, 
    3.101938, 1.856303, 1.262323, 1.104375, 0.9617674, 0.8446741, 0.6973521, 
    0.5712525, 0.5601974, 2.226754, 10.78853, 5.545442, 3.086288, 2.122358, 
    1.781009,
  1.466566, 3.07208, 15.65668, 9.034243, 3.655318, 1.747138, 1.322138, 
    1.083938, 1.147431, 6.181088, 13.28317, 13.03187, 10.59657, 4.105237, 
    2.066879, 1.261003, 0.9711702, 0.8862756, 0.8043081, 0.6739514, 
    0.5259049, 0.4752215, 0.6071358, 3.22578, 19.17207, 8.722011, 3.147111, 
    1.818996, 1.486604,
  2.707603, 15.06629, 21.6807, 8.407033, 4.34542, 1.402639, 1.525194, 
    2.185358, 4.565084, 11.27824, 15.45964, 12.66806, 5.36505, 1.890867, 
    1.153028, 0.6905299, 0.5946342, 0.5577463, 0.4633762, 0.4729553, 
    0.444284, 0.4660149, 0.6062732, 5.24531, 22.18809, 13.91603, 3.556915, 
    1.854172, 1.977766,
  6.135055, 16.98421, 22.74812, 11.76113, 2.759933, 1.434081, 1.326125, 
    2.39081, 3.710555, 5.47069, 6.05842, 4.392343, 2.086513, 0.6073839, 
    0.4317492, 0.3897203, 0.3913247, 0.4432462, 0.6373263, 1.214005, 
    2.148175, 3.974837, 8.2977, 21.86011, 20.78524, 15.85231, 2.595571, 
    2.23235, 3.419478,
  20.29289, 30.91133, 36.45091, 14.76221, 3.82661, 3.344558, 3.017039, 
    2.884474, 6.405555, 9.466175, 3.668474, 1.656259, 0.6458443, 0.3182206, 
    0.333087, 0.3936835, 0.5384457, 0.878512, 1.442624, 2.393359, 4.783398, 
    9.460814, 16.98895, 24.55241, 18.85317, 6.561572, 5.106865, 8.246495, 
    14.81461,
  36.87286, 35.18812, 32.06027, 27.45358, 12.70126, 7.705986, 12.30379, 
    8.256194, 7.495923, 4.711476, 2.999479, 1.338277, 0.8145335, 0.675541, 
    0.6781734, 0.7571543, 0.8818407, 1.239831, 1.750959, 2.483635, 3.563869, 
    5.455102, 7.204723, 11.23081, 3.919749, 5.298284, 8.365515, 19.59606, 
    34.18354,
  24.26654, 22.15557, 16.57142, 20.13391, 25.77207, 14.04066, 17.85447, 
    17.94522, 18.19974, 13.68313, 7.397712, 3.807227, 2.627676, 2.421133, 
    2.166299, 2.004745, 1.848147, 1.667704, 1.888233, 2.896122, 7.171883, 
    11.17646, 4.394112, 3.755419, 3.007984, 4.077683, 5.856454, 12.16492, 
    23.32968,
  20.53953, 17.32812, 13.07375, 22.03391, 23.27485, 23.74318, 29.36949, 
    20.55548, 29.5816, 26.7072, 12.79363, 8.668318, 6.540674, 5.204111, 
    4.518366, 3.968597, 3.253341, 2.570776, 2.238105, 3.544799, 13.2541, 
    15.9989, 9.911629, 6.37314, 3.966567, 3.575547, 4.003356, 4.59738, 
    13.93842,
  12.13503, 13.60344, 16.814, 20.1941, 27.5256, 22.65849, 26.9775, 30.33513, 
    29.72493, 22.5359, 20.73744, 16.82527, 11.28919, 8.072392, 6.847134, 
    5.344268, 4.255867, 3.623014, 3.263218, 6.298736, 15.34353, 23.72318, 
    18.12937, 16.91557, 12.94476, 7.292594, 5.680798, 5.082811, 6.579854,
  7.157508, 11.96028, 15.3679, 16.1221, 17.55192, 18.30826, 17.16439, 
    14.26761, 18.67347, 22.95003, 24.0303, 20.37411, 15.29792, 11.71128, 
    9.805962, 7.406773, 5.984389, 5.163795, 5.285478, 7.936758, 18.44687, 
    19.48613, 20.54959, 19.66008, 16.48587, 11.75288, 8.229002, 6.682563, 
    6.07757,
  7.961988, 10.88698, 11.99682, 13.13851, 14.23609, 15.76374, 16.4157, 
    16.55846, 17.3875, 18.0301, 16.58999, 14.26009, 12.97351, 12.21547, 
    10.17174, 8.340565, 7.01545, 7.592986, 8.741837, 12.49946, 11.84995, 
    11.38443, 11.04987, 11.818, 12.69249, 10.69039, 8.0493, 7.369631, 7.159806,
  6.687086, 7.780337, 8.879145, 10.04912, 10.49986, 10.91548, 11.13767, 
    13.12206, 13.98386, 13.1603, 12.03609, 11.16882, 8.793093, 8.357296, 
    7.818082, 7.193128, 7.870294, 9.153779, 9.252534, 9.460589, 7.98998, 
    7.406197, 8.109261, 8.430635, 7.487708, 7.230182, 5.980449, 6.566087, 
    6.497423,
  6.578145, 6.545788, 6.644692, 6.749643, 6.858003, 6.917331, 7.106503, 
    7.784645, 8.017767, 7.621871, 6.975715, 6.73995, 6.307418, 5.837615, 
    5.692236, 5.675409, 5.623599, 5.408085, 5.491864, 5.811483, 6.099625, 
    6.653283, 6.305056, 6.361547, 6.49225, 6.092087, 6.044433, 6.514158, 
    6.633337,
  0.3832363, 0.3832363, 0.3832363, 0.3832363, 0.3832363, 0.3832363, 
    0.3832363, 0.3820756, 0.3820756, 0.3820756, 0.3820756, 0.3820756, 
    0.3820756, 0.3820756, 0.3793736, 0.3793736, 0.3793736, 0.3793736, 
    0.3793736, 0.3793736, 0.3793736, 0.3839518, 0.3839518, 0.3839518, 
    0.3839518, 0.3839518, 0.3839518, 0.3839518, 0.3832363,
  0.4899096, 0.4624029, 0.4202379, 0.3802632, 0.3579387, 0.337604, 0.3264754, 
    0.3225245, 0.3179919, 0.3031692, 0.2780287, 0.2504113, 0.2460543, 
    0.1963304, 0.1759618, 0.1757491, 0.1873678, 0.2296842, 0.2914754, 
    0.3663132, 0.4527061, 0.4992244, 0.438715, 0.3017027, 0.3065691, 0.33452, 
    0.3413621, 0.4103253, 0.4879413,
  0.4044054, 0.3033728, 0.2963744, 0.2830952, 0.3992035, 0.3325425, 0.203369, 
    0.305023, 0.277345, 0.2633605, 0.2990518, 0.3289972, 0.2735697, 
    0.2360589, 0.2842024, 0.3146939, 0.3007012, 0.2844258, 0.2841693, 
    0.2842548, 0.2907679, 0.3429525, 0.4088145, 0.6273406, 0.7244567, 
    0.6516713, 0.6153069, 0.6064183, 0.5414888,
  0.885241, 0.7523897, 0.693687, 0.6328033, 0.6761534, 0.5843587, 0.4440398, 
    0.3624651, 0.3140198, 0.2908084, 0.3231272, 0.4717853, 0.670896, 
    1.053337, 1.144096, 1.131832, 0.941299, 0.7944202, 0.6051133, 0.4740144, 
    0.4369059, 0.4178446, 0.4404194, 0.5741145, 1.298276, 1.59253, 1.45301, 
    1.357493, 1.0306,
  1.357117, 1.124512, 1.067259, 1.182987, 1.158342, 0.9569099, 0.7989311, 
    0.6030589, 0.4925699, 0.4147134, 0.5241905, 1.126398, 2.126367, 2.204551, 
    2.368854, 1.824086, 1.400103, 1.015933, 0.8134069, 0.6591733, 0.5855291, 
    0.4803548, 0.4406418, 1.489789, 4.461671, 3.606762, 2.974491, 2.251354, 
    1.62791,
  1.604343, 1.417054, 2.307228, 2.736397, 1.901823, 1.266767, 0.9370675, 
    0.8216289, 0.7237319, 0.870407, 2.015956, 3.601232, 6.618871, 4.074807, 
    3.452029, 1.813602, 1.144346, 1.009635, 0.8856802, 0.7695436, 0.6170646, 
    0.4970802, 0.4983637, 2.846368, 12.37223, 6.058254, 3.239754, 2.156894, 
    1.761698,
  1.344482, 3.396056, 18.60291, 8.655795, 3.338038, 1.50662, 1.121983, 
    0.9611779, 1.153103, 7.317776, 16.37161, 16.23593, 12.71395, 4.206285, 
    2.0286, 1.224177, 0.8927377, 0.807994, 0.7287461, 0.5980514, 0.479803, 
    0.4221528, 0.5772795, 4.30637, 22.26, 9.371544, 2.929219, 1.812318, 
    1.436096,
  2.478676, 16.70584, 25.16429, 9.323431, 4.207021, 1.183526, 1.373652, 
    2.213342, 4.925392, 13.6751, 19.40067, 16.523, 6.234447, 1.838058, 
    1.09287, 0.6485007, 0.5315251, 0.5101609, 0.4630382, 0.4203369, 
    0.4213906, 0.4483731, 0.6060815, 5.517804, 26.2364, 16.4755, 3.085003, 
    1.700222, 1.689037,
  5.362932, 18.26242, 25.79423, 13.60037, 2.60777, 1.338299, 1.346726, 
    2.679835, 4.663726, 6.932564, 7.92607, 4.85526, 2.204356, 0.5747242, 
    0.4031458, 0.3802089, 0.416705, 0.4753186, 0.7420189, 1.310914, 2.239328, 
    3.749348, 7.088876, 25.52165, 24.70309, 17.87877, 2.510877, 2.196773, 
    3.230926,
  21.2741, 34.8923, 39.77601, 17.44307, 3.738741, 3.255439, 3.175279, 
    3.03424, 7.408769, 11.20793, 3.86983, 1.648629, 0.6153924, 0.3284483, 
    0.369095, 0.4621482, 0.6824427, 1.105182, 1.840999, 3.039343, 5.512748, 
    9.758264, 16.60134, 27.55995, 21.2866, 7.635611, 5.831979, 9.242441, 
    15.7971,
  40.45536, 37.96, 33.43027, 29.34159, 13.97442, 8.37344, 14.19781, 9.030463, 
    9.013894, 5.25215, 3.386667, 1.390994, 0.8027158, 0.6659303, 0.6992704, 
    0.7766389, 0.9390062, 1.381549, 1.917418, 2.750042, 4.089434, 6.397778, 
    7.633229, 13.27069, 3.927611, 5.483296, 8.645574, 21.0999, 38.66949,
  27.08154, 25.28192, 18.87174, 23.07543, 28.7173, 16.11996, 21.00794, 
    20.76794, 22.11959, 14.4448, 7.657791, 3.844576, 2.655928, 2.46412, 
    2.180624, 2.009852, 1.899846, 1.761371, 2.019784, 2.934994, 7.231152, 
    12.93899, 5.079524, 4.492643, 3.115471, 4.255826, 5.97727, 12.14717, 
    24.72252,
  22.91254, 19.94258, 15.61046, 24.92221, 26.08474, 27.0714, 31.91392, 
    23.57844, 32.28889, 29.26031, 13.79697, 9.220464, 6.656037, 5.156769, 
    4.354654, 3.87157, 3.244992, 2.493988, 2.387487, 3.947398, 15.24037, 
    18.3751, 11.52911, 7.575526, 4.452265, 3.784936, 4.057501, 4.860924, 
    16.19494,
  14.14837, 15.53618, 20.37363, 23.14493, 30.77959, 26.35527, 29.80809, 
    33.43856, 33.11455, 26.02102, 24.53599, 19.79248, 12.51495, 8.461738, 
    6.946235, 5.391077, 4.308868, 3.689099, 3.419246, 8.215521, 17.05064, 
    27.25766, 21.80208, 20.66388, 14.45762, 8.041, 6.215219, 5.525047, 
    7.781336,
  8.120388, 14.22766, 19.07595, 19.43532, 20.71246, 20.9964, 20.1812, 
    16.18697, 21.34296, 26.52353, 28.47037, 23.90963, 17.40517, 12.76077, 
    10.44202, 7.78065, 6.400331, 5.501381, 5.786572, 9.477644, 21.93315, 
    23.92785, 24.74377, 23.23017, 18.94778, 13.36309, 8.938417, 7.05487, 
    6.607942,
  8.770526, 12.60324, 14.05229, 15.63515, 16.39507, 18.86638, 19.30643, 
    19.66471, 20.3422, 21.17217, 19.10759, 16.18901, 14.48853, 13.82787, 
    11.39625, 8.99253, 7.901891, 8.627339, 10.09458, 15.13679, 14.33234, 
    14.01215, 12.76638, 13.33084, 13.94618, 11.21888, 8.511889, 7.679687, 
    7.692115,
  7.209328, 8.588437, 9.675194, 11.45935, 11.57967, 12.15997, 12.38846, 
    14.9875, 15.57141, 14.97762, 13.71889, 12.56438, 9.684513, 9.151197, 
    8.675642, 7.975615, 8.932359, 10.54526, 10.63053, 10.72707, 9.10471, 
    8.230968, 8.809004, 8.821998, 7.828562, 7.282715, 6.043844, 6.679046, 
    6.913458,
  7.035, 7.254782, 7.302457, 7.489509, 7.610951, 7.615198, 7.662448, 
    8.359349, 8.73809, 8.474346, 7.898699, 7.522389, 7.051041, 6.49839, 
    6.236814, 6.15081, 6.112026, 5.922946, 5.959836, 6.255219, 6.558084, 
    7.235652, 6.675109, 6.660504, 6.695848, 6.306252, 6.235679, 6.731382, 
    6.990803,
  0.3667257, 0.3667257, 0.3667257, 0.3667257, 0.3667257, 0.3667257, 
    0.3667257, 0.3685054, 0.3685054, 0.3685054, 0.3685054, 0.3685054, 
    0.3685054, 0.3685054, 0.3699599, 0.3699599, 0.3699599, 0.3699599, 
    0.3699599, 0.3699599, 0.3699599, 0.3728617, 0.3728617, 0.3728617, 
    0.3728617, 0.3728617, 0.3728617, 0.3728617, 0.3667257,
  0.4574514, 0.4291912, 0.394164, 0.3568431, 0.3359155, 0.3160163, 0.3087613, 
    0.3023497, 0.3005219, 0.2920766, 0.2695379, 0.2446864, 0.2379205, 
    0.1913978, 0.1656415, 0.1587273, 0.1698378, 0.2141409, 0.2798944, 
    0.3622836, 0.4408643, 0.4857354, 0.4023469, 0.25365, 0.2737024, 
    0.3044178, 0.3216255, 0.3853572, 0.4556844,
  0.3542458, 0.2626303, 0.2553235, 0.2486712, 0.3562017, 0.3000707, 
    0.1841891, 0.2806011, 0.2531691, 0.2418619, 0.2776006, 0.3026238, 
    0.2520091, 0.2120994, 0.2541173, 0.2805907, 0.267989, 0.2614253, 
    0.2655049, 0.264277, 0.2736966, 0.3241136, 0.3999279, 0.6424609, 
    0.7255476, 0.6539515, 0.6006919, 0.5726715, 0.4912397,
  0.8582913, 0.7109588, 0.6447269, 0.5902295, 0.6178772, 0.5201873, 
    0.4007677, 0.3254013, 0.2835688, 0.2633156, 0.288418, 0.4241901, 
    0.6393705, 1.046992, 1.122564, 1.084315, 0.8893315, 0.7516857, 0.5595967, 
    0.440465, 0.413702, 0.3910812, 0.43733, 0.6615674, 1.53137, 1.69244, 
    1.502589, 1.357373, 1.016668,
  1.34357, 1.080929, 1.031083, 1.122588, 1.077267, 0.8642894, 0.7090699, 
    0.5331672, 0.4414493, 0.3768462, 0.479237, 1.105836, 2.165102, 2.211464, 
    2.498381, 1.910912, 1.348033, 0.9500659, 0.7687278, 0.6062427, 0.5379345, 
    0.4293957, 0.4112355, 2.031178, 5.290592, 3.978406, 3.071934, 2.250593, 
    1.58873,
  1.531617, 1.345262, 2.389089, 2.572446, 1.700919, 1.117976, 0.8354535, 
    0.7356476, 0.6260567, 0.7932659, 1.976169, 3.780631, 7.404168, 4.047686, 
    3.960117, 1.757777, 1.086758, 0.9251159, 0.825273, 0.7005875, 0.5448142, 
    0.4394912, 0.4447745, 3.860695, 14.05495, 6.584818, 3.366108, 2.165103, 
    1.755915,
  1.215661, 3.817953, 21.44972, 8.008595, 2.949216, 1.267839, 0.9064662, 
    0.8285385, 1.206176, 8.506853, 19.21519, 19.90723, 15.0744, 4.164995, 
    1.982156, 1.180028, 0.843457, 0.7334083, 0.6333186, 0.5364652, 0.4278041, 
    0.3775416, 0.5200117, 6.060381, 24.86408, 9.800185, 2.758905, 1.801934, 
    1.323465,
  2.455839, 18.57788, 29.0511, 10.0192, 3.876036, 1.030713, 1.192979, 
    2.131498, 5.288917, 16.77507, 25.44571, 21.48366, 7.025754, 1.92871, 
    1.066435, 0.6055843, 0.5046763, 0.484107, 0.4212742, 0.3646232, 
    0.3955965, 0.4337988, 0.6726713, 5.821026, 30.10073, 19.30542, 2.678189, 
    1.444262, 1.495382,
  4.620668, 19.28695, 29.08187, 14.82054, 2.370679, 1.304827, 1.36924, 
    2.85968, 5.322187, 8.085499, 9.970526, 5.297409, 2.381432, 0.5617358, 
    0.3860708, 0.3769598, 0.4387105, 0.502032, 0.7487975, 1.282566, 2.09739, 
    3.044463, 5.745752, 29.83631, 29.04722, 20.02066, 2.373699, 2.079779, 
    2.939798,
  21.07084, 39.00314, 42.91445, 19.27917, 3.934272, 3.340848, 3.329525, 
    3.194141, 8.62009, 13.38005, 4.07907, 1.658625, 0.5880765, 0.3373507, 
    0.3981131, 0.5243492, 0.7994668, 1.264269, 2.093786, 3.560509, 5.810071, 
    9.389239, 15.82424, 30.35279, 23.239, 8.484779, 6.322619, 9.914835, 
    16.25399,
  43.28202, 40.91094, 34.33698, 30.62278, 15.20993, 9.39865, 15.57221, 
    9.867632, 10.76473, 5.766772, 3.775033, 1.435884, 0.7913457, 0.675553, 
    0.7305834, 0.8115465, 1.020882, 1.532818, 2.071408, 2.961455, 4.548304, 
    7.374977, 7.91138, 14.89841, 3.880491, 5.607063, 9.239446, 21.46683, 
    42.54817,
  30.8562, 29.21225, 21.9433, 25.52228, 31.53077, 19.12131, 24.3898, 
    23.38928, 26.79556, 15.23486, 7.786148, 3.874858, 2.677786, 2.499191, 
    2.207991, 2.013404, 1.948131, 1.922307, 2.233807, 3.132107, 7.334923, 
    14.68695, 5.788487, 4.961314, 3.108633, 4.321728, 6.154844, 12.95741, 
    27.59772,
  25.37413, 22.86121, 18.38214, 28.27559, 28.82274, 30.61086, 34.38379, 
    26.22604, 34.89017, 33.34724, 15.46763, 10.11019, 6.951175, 5.198063, 
    4.268704, 3.798202, 3.272169, 2.540457, 2.72713, 4.728632, 17.44815, 
    20.79552, 13.99709, 9.017835, 4.931867, 4.04852, 4.173453, 5.421417, 
    18.80645,
  16.23282, 17.77622, 24.10018, 25.97779, 34.30159, 30.26506, 32.83125, 
    36.8998, 37.06647, 30.50228, 29.11271, 22.68177, 13.78284, 8.838976, 
    7.040266, 5.431226, 4.373853, 3.76941, 3.689238, 10.51638, 19.01406, 
    31.39, 26.47513, 25.40521, 16.17795, 8.6972, 6.739916, 5.914715, 9.332684,
  9.496808, 17.16258, 23.41527, 23.39575, 24.33611, 24.82932, 23.43552, 
    18.58679, 24.61406, 30.82045, 33.81417, 28.18447, 20.25916, 13.94689, 
    11.13019, 8.254499, 6.872941, 6.080224, 6.381222, 11.43473, 25.75702, 
    28.95134, 29.78518, 27.4511, 22.03591, 15.06525, 9.644139, 7.48894, 
    7.263213,
  9.587476, 14.73947, 16.83693, 18.87626, 19.48131, 23.16558, 23.35042, 
    23.44415, 24.43804, 25.08626, 22.73173, 18.69912, 16.16602, 15.58021, 
    13.01963, 9.827241, 9.081457, 9.951239, 11.68347, 18.26493, 18.05871, 
    16.94761, 15.08612, 15.28727, 15.48492, 11.49157, 8.939387, 8.014206, 
    8.13476,
  7.706934, 9.472034, 10.65186, 13.20557, 13.10193, 13.6838, 14.20504, 
    17.558, 17.45341, 17.04863, 15.84054, 14.31336, 10.70105, 10.27672, 
    9.802412, 8.954913, 10.24045, 12.19516, 12.11382, 12.41731, 10.50664, 
    9.35717, 9.676415, 9.246696, 8.157457, 7.286966, 6.10306, 6.703836, 
    7.388376,
  7.461308, 7.878256, 8.043123, 8.394089, 8.53938, 8.602348, 8.471208, 
    9.218724, 9.803187, 9.514413, 8.875523, 8.422179, 7.881443, 7.201825, 
    6.772885, 6.611806, 6.536366, 6.420842, 6.466784, 6.761983, 7.224706, 
    7.948883, 7.145464, 6.94827, 6.832455, 6.503559, 6.452115, 6.915193, 
    7.333494,
  0.3462757, 0.3462757, 0.3462757, 0.3462757, 0.3462757, 0.3462757, 
    0.3462757, 0.3495463, 0.3495463, 0.3495463, 0.3495463, 0.3495463, 
    0.3495463, 0.3495463, 0.355843, 0.355843, 0.355843, 0.355843, 0.355843, 
    0.355843, 0.355843, 0.3553828, 0.3553828, 0.3553828, 0.3553828, 
    0.3553828, 0.3553828, 0.3553828, 0.3462757,
  0.4236823, 0.3943839, 0.3672689, 0.3349462, 0.3134347, 0.296165, 0.293755, 
    0.2874056, 0.2853164, 0.2801884, 0.260725, 0.241383, 0.2321332, 
    0.1915144, 0.1598514, 0.1480212, 0.1576567, 0.2011716, 0.2701315, 0.3539, 
    0.4172223, 0.462125, 0.3611125, 0.2185568, 0.2447109, 0.2766556, 
    0.2992012, 0.3588043, 0.4235211,
  0.3111185, 0.2307027, 0.2217793, 0.2223802, 0.3186893, 0.2707035, 
    0.1730474, 0.2581228, 0.2337924, 0.2231082, 0.2567524, 0.2778741, 
    0.2333628, 0.1923703, 0.2323375, 0.256648, 0.2445917, 0.2400416, 
    0.2473281, 0.2439475, 0.260694, 0.3159688, 0.3973715, 0.6439781, 
    0.7048929, 0.6517961, 0.5804245, 0.5478678, 0.4391479,
  0.8290261, 0.6698864, 0.6008868, 0.5477772, 0.5580813, 0.4588512, 
    0.3566345, 0.2929993, 0.2572547, 0.2392156, 0.2601468, 0.3857266, 
    0.5973021, 1.016313, 1.077413, 1.045842, 0.8519537, 0.7241485, 0.5250114, 
    0.4136149, 0.3966953, 0.3660962, 0.4246188, 0.7468528, 1.775279, 
    1.809995, 1.550519, 1.350671, 1.011735,
  1.304128, 1.022298, 1.001862, 1.067882, 0.9804663, 0.7764918, 0.6235155, 
    0.4711208, 0.3977833, 0.3386725, 0.4303885, 1.065318, 2.188833, 2.184814, 
    2.633015, 1.97396, 1.287665, 0.8961787, 0.7187962, 0.5663822, 0.4996753, 
    0.3923282, 0.4029365, 2.88128, 6.204134, 4.346931, 3.183319, 2.235033, 
    1.560753,
  1.453739, 1.294906, 2.474543, 2.416565, 1.491149, 0.9983609, 0.7427954, 
    0.641924, 0.5444639, 0.7254828, 2.026619, 3.97099, 7.898492, 3.909817, 
    4.746253, 1.713672, 1.049441, 0.8554367, 0.7656273, 0.6416389, 0.4901829, 
    0.4004462, 0.3958946, 5.337112, 15.727, 6.937577, 3.374883, 2.135844, 
    1.698927,
  1.098862, 4.280504, 24.41059, 7.18603, 2.603429, 1.075636, 0.7601134, 
    0.7257814, 1.206381, 9.781746, 21.89525, 23.25068, 17.50946, 4.066898, 
    1.956592, 1.155042, 0.8083913, 0.6582178, 0.5504593, 0.474999, 0.3920539, 
    0.3422437, 0.4778291, 8.922709, 27.5569, 10.10947, 2.605178, 1.74538, 
    1.23749,
  2.645393, 20.71811, 32.32867, 10.30437, 3.421922, 0.9400714, 1.085965, 
    2.010328, 5.580694, 19.74032, 31.79512, 25.8655, 7.410388, 2.166964, 
    1.093121, 0.5905727, 0.4915293, 0.4539645, 0.3992115, 0.3346802, 
    0.3634879, 0.4484121, 0.8038743, 6.10745, 33.80865, 22.21694, 2.3053, 
    1.182494, 1.345206,
  4.40984, 19.69232, 32.30835, 15.64968, 2.104403, 1.283754, 1.393139, 
    2.959644, 5.759048, 8.938041, 11.79545, 5.681771, 2.538718, 0.5626586, 
    0.3760407, 0.3790862, 0.457431, 0.5254663, 0.7184663, 1.078315, 1.709772, 
    2.201853, 4.444524, 34.05693, 32.16734, 21.93473, 2.304546, 1.819506, 
    2.628636,
  20.07422, 43.04986, 46.1427, 20.5451, 4.070459, 3.489347, 3.582031, 
    3.377841, 9.93291, 15.77645, 4.262049, 1.710491, 0.5609954, 0.3446358, 
    0.4211998, 0.5709763, 0.8495892, 1.3214, 2.093626, 3.458328, 5.464911, 
    8.683701, 14.77247, 33.08001, 24.80404, 9.352555, 6.820048, 10.46006, 
    16.14051,
  44.66453, 43.83819, 36.36624, 31.50377, 17.06574, 10.15439, 16.41837, 
    10.65519, 12.85976, 6.13189, 4.17193, 1.472759, 0.7899065, 0.7021524, 
    0.7715862, 0.8615083, 1.102767, 1.680098, 2.224296, 3.155253, 5.016109, 
    8.406199, 8.124877, 16.16788, 3.878067, 5.574875, 9.965089, 21.64676, 
    45.09813,
  35.4838, 34.45292, 26.16484, 27.71416, 34.18635, 22.28388, 27.90285, 
    26.58454, 32.13401, 17.02295, 8.018797, 4.249341, 2.855486, 2.501021, 
    2.222167, 2.080895, 2.029919, 2.094383, 2.820071, 3.615696, 7.819006, 
    16.3723, 6.673151, 5.18052, 3.020288, 4.12641, 6.411469, 15.4842, 32.1269,
  28.46527, 25.91645, 21.53134, 31.55699, 31.5157, 34.40208, 37.32357, 
    28.66173, 37.52815, 38.85858, 17.91098, 11.01987, 7.287473, 5.359811, 
    4.178808, 3.773295, 3.3039, 2.644864, 3.16103, 6.008791, 20.10067, 
    23.9379, 17.39814, 10.46526, 5.509471, 4.354057, 4.263019, 6.334334, 
    22.04707,
  18.38602, 20.24333, 27.70908, 28.78536, 38.25917, 35.35644, 36.15292, 
    40.6102, 41.52788, 35.72441, 34.38867, 25.34962, 14.92418, 9.137508, 
    7.16148, 5.540689, 4.535516, 3.910046, 4.003147, 13.07222, 21.37402, 
    35.54132, 32.03426, 31.04863, 17.82271, 9.514213, 7.159223, 6.356985, 
    11.19221,
  11.36555, 21.09558, 28.52271, 28.66002, 28.54116, 29.94429, 27.63861, 
    21.48142, 28.59485, 35.93923, 40.80503, 33.78503, 23.35386, 15.35575, 
    11.8601, 8.864632, 7.419206, 6.742994, 7.258162, 13.94326, 29.68448, 
    34.97628, 36.34908, 32.76411, 25.87766, 16.69445, 10.21017, 7.897784, 
    8.098112,
  10.41047, 17.26632, 20.43291, 23.3175, 23.76575, 28.19465, 28.30293, 
    28.71336, 28.9307, 29.99661, 27.39299, 21.85447, 18.10973, 17.45434, 
    15.28438, 11.01285, 10.57159, 11.60562, 13.70783, 22.02791, 23.13647, 
    21.00633, 17.8952, 17.9303, 17.45518, 11.60838, 9.280901, 8.276714, 
    8.42634,
  8.211338, 10.50012, 11.74257, 15.29927, 15.136, 15.61109, 16.26198, 
    20.8723, 19.99639, 19.45288, 18.10363, 16.49919, 11.96111, 11.75704, 
    11.19747, 10.0947, 11.85749, 13.96628, 13.80989, 14.53255, 12.14585, 
    10.9032, 10.55405, 9.723451, 8.401114, 7.24875, 6.156647, 6.635741, 
    7.765688,
  7.932371, 8.404545, 8.717588, 9.166247, 9.391902, 9.510145, 9.452088, 
    10.28029, 10.89123, 10.65103, 9.941803, 9.267712, 8.673544, 7.960766, 
    7.348455, 7.073458, 7.035006, 6.973152, 7.0562, 7.41619, 7.924155, 
    8.579957, 7.613885, 7.209932, 6.896266, 6.621529, 6.631999, 7.036543, 
    7.634778,
  0.3244964, 0.3244964, 0.3244964, 0.3244964, 0.3244964, 0.3244964, 
    0.3244964, 0.3271607, 0.3271607, 0.3271607, 0.3271607, 0.3271607, 
    0.3271607, 0.3271607, 0.3375499, 0.3375499, 0.3375499, 0.3375499, 
    0.3375499, 0.3375499, 0.3375499, 0.3346604, 0.3346604, 0.3346604, 
    0.3346604, 0.3346604, 0.3346604, 0.3346604, 0.3244964,
  0.391773, 0.3641616, 0.3424391, 0.3168554, 0.292821, 0.2803345, 0.2827678, 
    0.2765504, 0.273129, 0.2675185, 0.2499967, 0.2364015, 0.2253762, 
    0.1940584, 0.1574671, 0.1415532, 0.1496173, 0.1909012, 0.2587089, 
    0.3339358, 0.3858699, 0.4331014, 0.3203408, 0.1941391, 0.2184076, 
    0.2523873, 0.2816573, 0.3332754, 0.3896173,
  0.2764772, 0.2070163, 0.1983167, 0.2044722, 0.2874594, 0.2451795, 
    0.1671257, 0.2374014, 0.2179208, 0.208743, 0.2378761, 0.2548732, 
    0.2161751, 0.177461, 0.2149107, 0.2421802, 0.2231118, 0.2216195, 
    0.2306386, 0.2264303, 0.2450825, 0.3146878, 0.3923477, 0.6335233, 
    0.6646957, 0.6405708, 0.5562404, 0.5259759, 0.3924679,
  0.7992578, 0.6308751, 0.5589734, 0.5097976, 0.5001655, 0.4028924, 
    0.3230627, 0.268932, 0.2373297, 0.2186882, 0.2365696, 0.3539045, 
    0.5554302, 0.9666269, 1.027765, 1.016654, 0.8315098, 0.7034906, 
    0.5018585, 0.3938207, 0.3772132, 0.3369278, 0.4140064, 0.7957342, 
    2.00516, 1.958931, 1.611436, 1.359007, 1.002461,
  1.253482, 0.9537882, 0.955713, 1.014349, 0.8771009, 0.6930505, 0.5518556, 
    0.4217963, 0.3651417, 0.3136337, 0.3927554, 1.047525, 2.190076, 2.103097, 
    2.719383, 1.960067, 1.240487, 0.855365, 0.6711187, 0.5310189, 0.4604116, 
    0.3614706, 0.4099751, 4.154278, 7.235686, 4.713137, 3.294953, 2.24549, 
    1.532162,
  1.37349, 1.249838, 2.522552, 2.237575, 1.315282, 0.8938813, 0.6610383, 
    0.5641226, 0.4820106, 0.6542497, 2.091426, 4.131217, 8.236808, 3.700481, 
    5.734743, 1.698852, 1.019892, 0.8041294, 0.7140177, 0.5893605, 0.4515062, 
    0.3708247, 0.3630847, 7.230724, 17.34609, 7.07256, 3.265384, 2.082263, 
    1.610244,
  1.020838, 4.795408, 27.47427, 6.362126, 2.264778, 0.9370927, 0.6807457, 
    0.6486016, 1.11328, 11.07504, 23.68792, 26.00743, 19.46078, 4.022589, 
    1.961774, 1.138123, 0.7762045, 0.6120303, 0.5066603, 0.4463006, 
    0.3762266, 0.3169618, 0.4654726, 12.66502, 30.22116, 10.22716, 2.453889, 
    1.632488, 1.155614,
  2.633666, 23.00751, 34.78015, 10.29066, 2.947056, 0.8889306, 1.0285, 
    1.904256, 5.384895, 21.41418, 35.83151, 28.77061, 7.309011, 2.231178, 
    1.129983, 0.5922453, 0.4830386, 0.4439882, 0.3884774, 0.3203078, 
    0.3317828, 0.4573924, 0.9319597, 6.572474, 37.57951, 25.39779, 1.944079, 
    0.9723887, 1.171552,
  4.378151, 19.97021, 34.75651, 16.14931, 1.873806, 1.271395, 1.429389, 
    3.061716, 6.157138, 9.748549, 13.40894, 6.05039, 2.663752, 0.5728459, 
    0.374493, 0.3854526, 0.473204, 0.5365762, 0.681553, 0.898434, 1.161418, 
    1.558144, 3.498665, 38.5986, 35.05719, 23.69142, 2.286236, 1.678656, 
    2.378527,
  19.10451, 45.73769, 48.58783, 21.60713, 4.226179, 3.711565, 3.884863, 
    3.568631, 11.24327, 18.27088, 4.459695, 1.790676, 0.5331821, 0.3490799, 
    0.4319998, 0.5981574, 0.8719444, 1.34088, 2.043723, 2.979912, 4.382503, 
    7.689887, 13.58928, 35.76878, 26.31118, 10.0697, 7.325376, 10.94744, 
    15.3069,
  45.51622, 45.93459, 40.4423, 32.19228, 18.62122, 10.63403, 17.04254, 
    11.6803, 15.66454, 6.509573, 4.610985, 1.496005, 0.7979457, 0.7370551, 
    0.8159936, 0.9090475, 1.167089, 1.78696, 2.359863, 3.35287, 5.54827, 
    9.521787, 8.356897, 17.18888, 3.918313, 5.500965, 10.5174, 22.10667, 
    46.48091,
  39.12715, 39.58943, 31.85941, 28.79021, 37.26564, 23.93793, 31.11972, 
    30.36345, 36.91997, 19.92497, 8.183193, 4.505254, 2.994521, 2.548875, 
    2.254117, 2.147141, 2.167638, 2.279025, 3.700128, 4.923031, 9.013468, 
    17.92537, 7.532234, 5.214803, 3.043668, 4.019678, 6.39076, 18.91237, 
    37.53944,
  31.907, 29.24637, 24.4835, 34.20125, 34.0885, 38.28404, 40.73328, 31.06764, 
    40.14557, 45.6109, 19.92288, 11.51329, 7.475352, 5.576447, 4.244038, 
    3.75108, 3.323383, 2.721256, 3.683075, 7.644316, 23.04862, 27.82862, 
    21.9214, 11.13097, 5.972847, 4.5946, 4.464247, 7.200501, 25.51722,
  20.66884, 22.71296, 30.76384, 31.55446, 42.61079, 41.66255, 39.33951, 
    44.95706, 46.10004, 40.99832, 39.3932, 27.37036, 15.55828, 9.497734, 
    7.380538, 5.705282, 4.710096, 4.091218, 4.293774, 15.86144, 24.15057, 
    39.68845, 38.43086, 35.96679, 18.84791, 10.14958, 7.531068, 6.830669, 
    12.96323,
  13.53843, 25.31721, 33.98457, 34.16428, 33.71641, 36.35735, 33.25582, 
    24.70456, 32.80097, 41.78598, 49.27696, 40.43228, 25.34147, 16.41875, 
    12.51231, 9.323329, 7.894077, 7.292753, 8.085351, 16.87054, 33.76046, 
    41.54997, 44.01992, 39.38029, 30.19443, 18.19746, 10.63082, 8.196397, 
    8.9414,
  11.15969, 20.25865, 24.51188, 28.64936, 29.37, 34.37211, 34.89632, 
    35.34592, 33.85913, 35.45825, 32.41059, 26.06371, 20.34761, 19.67717, 
    17.83248, 12.35802, 12.43354, 13.69675, 16.52717, 26.29335, 29.11024, 
    25.8321, 21.01519, 21.46037, 19.71992, 11.5497, 9.494921, 8.45011, 
    8.642234,
  8.611874, 11.69968, 13.14308, 17.59314, 17.37902, 17.92924, 18.91511, 
    24.7627, 23.0667, 21.97334, 21.01541, 19.12931, 13.60423, 13.44072, 
    12.76952, 11.34512, 13.78642, 16.17424, 16.03458, 17.34426, 14.12273, 
    12.76855, 11.45092, 10.32434, 8.680073, 7.232746, 6.203416, 6.496451, 
    8.049904,
  8.256494, 8.731441, 9.182814, 9.838589, 10.13735, 10.33243, 10.32986, 
    11.33131, 12.06312, 11.84785, 11.13786, 10.13213, 9.601747, 8.802797, 
    8.133006, 7.66065, 7.610837, 7.640581, 7.772218, 8.161711, 8.459115, 
    8.935887, 7.885978, 7.370434, 6.895183, 6.618686, 6.73756, 7.111141, 
    7.773888,
  0.3042182, 0.3042182, 0.3042182, 0.3042182, 0.3042182, 0.3042182, 
    0.3042182, 0.3045327, 0.3045327, 0.3045327, 0.3045327, 0.3045327, 
    0.3045327, 0.3045327, 0.3165859, 0.3165859, 0.3165859, 0.3165859, 
    0.3165859, 0.3165859, 0.3165859, 0.3126008, 0.3126008, 0.3126008, 
    0.3126008, 0.3126008, 0.3126008, 0.3126008, 0.3042182,
  0.3598081, 0.3389662, 0.3204632, 0.3011059, 0.2740952, 0.2664527, 
    0.2729438, 0.2664903, 0.2628672, 0.2563532, 0.2388533, 0.2294094, 
    0.2190409, 0.1968824, 0.1587093, 0.1374193, 0.1448015, 0.1830011, 
    0.2494668, 0.3076253, 0.3541478, 0.3950881, 0.2844414, 0.1829451, 
    0.2005426, 0.2329277, 0.2638656, 0.3112431, 0.3542174,
  0.2514772, 0.1937573, 0.1826557, 0.1939231, 0.2617526, 0.2242711, 
    0.1654208, 0.220079, 0.204718, 0.1985382, 0.2230889, 0.2342817, 
    0.2019821, 0.165979, 0.1994793, 0.2305296, 0.2075161, 0.2078409, 
    0.2164363, 0.2139327, 0.2303542, 0.3091355, 0.3781721, 0.6083161, 
    0.6059603, 0.6126113, 0.5351714, 0.506016, 0.3576965,
  0.7584079, 0.5903142, 0.5199007, 0.4826134, 0.45574, 0.3652961, 0.2987963, 
    0.2511743, 0.2249078, 0.2029665, 0.2198999, 0.3154815, 0.5173258, 
    0.9048182, 0.9751431, 0.9936121, 0.8174467, 0.678012, 0.4760698, 
    0.3721968, 0.3610301, 0.3192358, 0.4063998, 0.8694144, 2.300082, 
    2.067605, 1.650583, 1.346043, 0.9797221,
  1.204741, 0.9098136, 0.9120667, 0.9650774, 0.7967632, 0.6276692, 0.5046528, 
    0.3936452, 0.3402839, 0.2972783, 0.3731434, 1.029731, 2.1258, 2.012161, 
    2.769474, 1.930138, 1.197554, 0.818098, 0.6371862, 0.5073768, 0.431998, 
    0.341671, 0.4379859, 5.964336, 8.311462, 5.130583, 3.411195, 2.21828, 
    1.511379,
  1.302056, 1.20616, 2.52404, 2.064523, 1.183618, 0.8109131, 0.6022639, 
    0.5189288, 0.4478242, 0.58617, 2.178532, 4.258528, 8.414788, 3.465292, 
    6.900643, 1.702036, 0.9992411, 0.766403, 0.6751468, 0.5570089, 0.4384651, 
    0.3530422, 0.3438458, 9.757444, 19.06081, 7.1433, 3.10814, 1.999742, 
    1.519982,
  0.9753464, 5.156218, 30.26581, 5.639658, 1.977852, 0.837662, 0.6371118, 
    0.6183863, 0.9840247, 11.75764, 25.21932, 28.25764, 21.00768, 3.954033, 
    1.950506, 1.118505, 0.7584782, 0.5947343, 0.4897573, 0.4431737, 
    0.3684887, 0.3043181, 0.504033, 16.9378, 32.832, 9.960816, 2.30684, 
    1.53662, 1.104158,
  2.44992, 25.49116, 36.62617, 10.15763, 2.604913, 0.8506456, 0.9784275, 
    1.837216, 5.230605, 22.76706, 38.3168, 30.82746, 6.953207, 2.164598, 
    1.163765, 0.6026797, 0.4747803, 0.4347305, 0.3825863, 0.3145013, 
    0.325358, 0.4319537, 1.023163, 7.165503, 40.74234, 28.0911, 1.700952, 
    0.860339, 1.078165,
  4.739861, 20.76887, 36.42972, 16.58467, 1.731129, 1.260281, 1.470585, 
    3.166143, 6.476044, 10.5126, 14.38139, 6.371586, 2.815137, 0.5832995, 
    0.3737211, 0.3925418, 0.4884571, 0.534348, 0.6392863, 0.7909049, 
    0.8407732, 1.115339, 2.983891, 41.92464, 37.14077, 25.29472, 2.320505, 
    1.614104, 2.258805,
  17.98384, 46.7757, 49.45661, 22.95266, 4.395116, 3.935292, 4.294931, 
    3.831066, 12.27589, 20.39913, 4.704121, 1.952101, 0.5068527, 0.3493933, 
    0.4348164, 0.612842, 0.8815684, 1.342524, 1.993177, 2.715392, 3.494008, 
    5.916258, 12.16943, 37.89321, 27.72363, 10.63206, 7.718067, 11.10649, 
    13.94591,
  46.32918, 47.65565, 43.46571, 32.8498, 19.78027, 11.18892, 17.82436, 
    12.18606, 18.78336, 6.940464, 5.112776, 1.516226, 0.8118585, 0.7799311, 
    0.8596026, 0.9538842, 1.233467, 1.872536, 2.477616, 3.534, 6.061944, 
    10.74516, 8.515302, 18.06256, 3.967982, 5.537735, 10.52849, 22.86489, 
    47.33332,
  42.0294, 43.48303, 37.80313, 29.42884, 39.82442, 23.48878, 33.99272, 
    35.97006, 40.58111, 22.81445, 8.361444, 4.769053, 3.112118, 2.624705, 
    2.31326, 2.21079, 2.325146, 2.46443, 4.43157, 6.741044, 11.06624, 
    19.4646, 8.332366, 5.226314, 3.088146, 3.970469, 6.348716, 19.9438, 
    41.69567,
  35.47463, 32.46556, 26.71442, 36.81687, 36.47857, 42.27617, 44.49369, 
    33.64421, 42.85855, 52.01925, 21.15437, 11.74834, 7.587725, 5.72179, 
    4.301936, 3.76278, 3.352118, 2.813844, 4.145469, 9.852335, 26.37344, 
    31.38326, 27.05026, 11.40422, 6.267755, 4.723913, 4.608436, 7.623996, 
    28.67611,
  23.03545, 24.55968, 33.55698, 34.38274, 46.87876, 47.67617, 42.67406, 
    50.32087, 51.15213, 45.84823, 43.89033, 28.74938, 15.86518, 9.752125, 
    7.588384, 5.87275, 4.757351, 4.201238, 4.462192, 19.16214, 27.47751, 
    44.17853, 45.21088, 39.77172, 19.27468, 10.63955, 7.776706, 7.200526, 
    14.65254,
  15.75042, 29.31396, 39.55978, 40.48244, 40.94271, 43.29388, 39.7904, 
    28.27222, 37.36502, 48.70565, 58.80163, 48.79034, 26.63826, 17.0923, 
    12.97161, 9.64352, 8.177211, 7.638453, 8.684125, 20.21661, 38.4179, 
    48.59164, 51.90409, 46.39997, 35.33175, 19.17716, 10.87986, 8.342421, 
    9.689906,
  11.71109, 23.21225, 28.45724, 34.59143, 36.33212, 41.75967, 42.86722, 
    42.76359, 39.47213, 42.13169, 38.84315, 31.06284, 22.87666, 22.22546, 
    19.87702, 13.86382, 14.86897, 16.25365, 20.40725, 31.06891, 36.00279, 
    31.05059, 23.70353, 25.24035, 21.35777, 11.43564, 9.68549, 8.530881, 
    8.832488,
  8.82204, 12.74534, 14.76319, 19.63055, 19.51498, 20.61778, 22.41022, 
    29.0439, 26.46441, 24.29195, 24.44175, 22.02066, 15.39314, 15.25204, 
    14.77567, 12.92414, 15.82679, 18.67323, 18.58849, 20.38345, 16.47138, 
    14.7895, 12.62518, 11.07666, 9.003844, 7.258638, 6.24142, 6.280935, 
    8.111358,
  8.397864, 9.002821, 9.570478, 10.30867, 10.79427, 11.08134, 11.10872, 
    12.20619, 13.13973, 12.83199, 12.1702, 11.24895, 10.64168, 9.684171, 
    8.962807, 8.387337, 8.313643, 8.324678, 8.575678, 8.806074, 8.801497, 
    9.050574, 7.974895, 7.413306, 6.82783, 6.586723, 6.784679, 7.101698, 
    7.833189,
  0.2848201, 0.2848201, 0.2848201, 0.2848201, 0.2848201, 0.2848201, 
    0.2848201, 0.2853207, 0.2853207, 0.2853207, 0.2853207, 0.2853207, 
    0.2853207, 0.2853207, 0.2954123, 0.2954123, 0.2954123, 0.2954123, 
    0.2954123, 0.2954123, 0.2954123, 0.2915037, 0.2915037, 0.2915037, 
    0.2915037, 0.2915037, 0.2915037, 0.2915037, 0.2848201,
  0.328214, 0.3159839, 0.3009551, 0.2861495, 0.2580537, 0.2546437, 0.2626553, 
    0.2573209, 0.2535215, 0.2464537, 0.2290314, 0.2206717, 0.2130396, 
    0.2002725, 0.1607543, 0.1350675, 0.1422252, 0.1767493, 0.2430355, 
    0.2846609, 0.3255002, 0.3569874, 0.2556303, 0.1795599, 0.1884281, 
    0.2187402, 0.2483899, 0.2908886, 0.3215177,
  0.2319537, 0.1867531, 0.1741056, 0.1897164, 0.2413288, 0.2087543, 
    0.1671494, 0.2070488, 0.1953138, 0.191437, 0.2124885, 0.2168566, 
    0.1916699, 0.1584662, 0.1841617, 0.2179472, 0.1961908, 0.1964199, 
    0.2046892, 0.2039151, 0.2164849, 0.2993293, 0.3604947, 0.5712714, 
    0.5402873, 0.5830353, 0.5091495, 0.477457, 0.3294961,
  0.7255617, 0.5525207, 0.4875671, 0.4618173, 0.418374, 0.3430391, 0.2845437, 
    0.2405048, 0.2166741, 0.191884, 0.2077807, 0.2836664, 0.4857616, 
    0.8607853, 0.9196951, 0.9715925, 0.8008094, 0.6596695, 0.4608826, 
    0.3607454, 0.3511347, 0.3114126, 0.4014891, 0.9555766, 2.546522, 
    2.201622, 1.707622, 1.307364, 0.932372,
  1.177239, 0.8780333, 0.8739491, 0.9307455, 0.7305788, 0.5746399, 0.4781436, 
    0.3785091, 0.3257652, 0.287447, 0.3629949, 1.01227, 2.065769, 1.927347, 
    2.892163, 1.886042, 1.156631, 0.7841834, 0.6189372, 0.4963218, 0.412116, 
    0.3255108, 0.4616226, 8.126836, 9.232982, 5.423574, 3.48298, 2.207872, 
    1.503574,
  1.261651, 1.179619, 2.506665, 1.927972, 1.089291, 0.7613739, 0.5655699, 
    0.4969848, 0.4283532, 0.5324185, 2.21962, 4.35672, 8.478412, 3.232068, 
    8.297275, 1.704072, 0.9813619, 0.7420186, 0.6517177, 0.5420364, 
    0.4315515, 0.3460662, 0.3314552, 12.58041, 20.84625, 7.089902, 2.937351, 
    1.910686, 1.455757,
  0.9674364, 5.27687, 32.63173, 5.256682, 1.780033, 0.7827367, 0.610432, 
    0.6046397, 0.9298304, 12.12749, 26.79536, 30.30852, 22.62701, 3.818431, 
    1.930377, 1.09776, 0.7405856, 0.5853412, 0.4827967, 0.4370279, 0.3662704, 
    0.303593, 0.5017619, 21.79011, 35.35196, 9.738926, 2.237053, 1.471341, 
    1.092821,
  2.330058, 28.21202, 38.42311, 10.00895, 2.440206, 0.8291886, 0.9454231, 
    1.797202, 5.069509, 23.37657, 40.209, 32.51875, 6.747941, 2.143096, 
    1.20488, 0.6111263, 0.4742603, 0.4291987, 0.3795674, 0.3121178, 
    0.3203327, 0.4245932, 1.077489, 8.488098, 42.79178, 30.13301, 1.586102, 
    0.826175, 1.042714,
  4.818342, 21.83476, 37.42682, 17.26038, 1.682011, 1.254174, 1.477188, 
    3.177873, 6.678986, 11.10787, 14.9217, 6.753458, 3.016077, 0.595291, 
    0.3768674, 0.398588, 0.4989243, 0.5319319, 0.5984822, 0.7039786, 
    0.7286611, 0.88881, 2.781086, 43.33889, 38.04436, 26.80748, 2.405651, 
    1.570933, 2.20978,
  17.02281, 46.54697, 49.32448, 24.43706, 4.583351, 4.122298, 4.498985, 
    4.032191, 12.96312, 21.48101, 5.031422, 2.074767, 0.4858827, 0.3477224, 
    0.4334399, 0.6179803, 0.8818915, 1.319658, 1.919883, 2.533915, 3.087802, 
    4.34621, 10.10578, 38.97718, 28.94215, 10.66687, 7.945529, 10.94326, 
    12.84491,
  47.07737, 49.10597, 45.47515, 33.63222, 20.61031, 11.42634, 18.7565, 
    12.37162, 20.97658, 7.338499, 5.555515, 1.53908, 0.832505, 0.8133162, 
    0.8940274, 0.9844486, 1.274957, 1.93968, 2.593353, 3.699045, 6.521428, 
    11.81001, 8.818147, 18.88979, 3.988377, 5.498798, 10.41594, 23.23438, 
    48.13507,
  44.19991, 46.42988, 41.91668, 30.22941, 41.68923, 22.0345, 36.67386, 
    38.88928, 43.78784, 24.86266, 8.478871, 4.922456, 3.181205, 2.672165, 
    2.362152, 2.250964, 2.417647, 2.551205, 4.838921, 7.972688, 12.58275, 
    20.90033, 8.717979, 5.421079, 3.086641, 3.915947, 6.16843, 19.66055, 
    44.35947,
  38.94937, 34.93196, 28.29532, 39.17208, 38.82181, 46.33071, 48.49012, 
    36.28552, 45.80614, 57.71458, 21.84574, 11.83655, 7.649889, 5.806996, 
    4.361428, 3.779678, 3.379532, 2.855798, 4.419649, 12.29496, 29.81551, 
    34.07414, 30.63029, 11.45956, 6.410104, 4.77974, 4.66663, 7.745412, 
    31.52752,
  25.34064, 25.65455, 35.88467, 37.23389, 51.34424, 54.02834, 45.96957, 
    56.64428, 56.47652, 50.33121, 47.72612, 29.66925, 16.00705, 9.872635, 
    7.641372, 5.94629, 4.772717, 4.231951, 4.524663, 22.7568, 31.24129, 
    49.04654, 51.19083, 42.4637, 19.37064, 10.85328, 7.910151, 7.38133, 
    16.46055,
  17.82272, 33.25114, 45.06201, 47.57487, 49.83572, 52.07869, 46.90311, 
    31.98609, 42.33389, 56.11146, 67.47573, 57.5612, 27.42294, 17.49892, 
    13.17189, 9.749908, 8.277813, 7.876444, 9.234707, 23.91779, 43.50895, 
    55.61522, 58.66427, 53.19869, 40.34343, 19.64198, 10.92814, 8.350735, 
    10.21213,
  12.12502, 26.10118, 33.44315, 40.86784, 43.42749, 49.67326, 51.00963, 
    50.62502, 45.33061, 50.25719, 47.64653, 36.91753, 25.71255, 25.28255, 
    21.13272, 15.36988, 18.22034, 19.11168, 25.05661, 36.74577, 43.98434, 
    36.81606, 26.63387, 28.95285, 22.63338, 11.34918, 9.773049, 8.571839, 
    8.982517,
  8.966546, 13.31889, 16.44467, 21.04173, 21.80197, 23.40908, 25.99588, 
    34.32482, 30.15576, 26.34011, 28.60997, 25.49604, 17.54499, 17.50617, 
    17.46416, 14.87308, 18.22549, 21.43703, 21.38826, 23.75439, 19.00307, 
    16.91483, 14.12365, 11.98174, 9.273975, 7.24793, 6.255347, 6.071609, 
    8.12697,
  8.406294, 9.154147, 10.0247, 10.89933, 11.51485, 11.6928, 12.00886, 
    13.09348, 14.01229, 13.6839, 13.30748, 12.6229, 11.77669, 10.61445, 
    9.811783, 9.161313, 9.04131, 9.034889, 9.27831, 9.462022, 9.131634, 
    8.994911, 7.963368, 7.383852, 6.731857, 6.557935, 6.789924, 7.074039, 
    7.802053,
  0.2643491, 0.2643491, 0.2643491, 0.2643491, 0.2643491, 0.2643491, 
    0.2643491, 0.2675646, 0.2675646, 0.2675646, 0.2675646, 0.2675646, 
    0.2675646, 0.2675646, 0.2763406, 0.2763406, 0.2763406, 0.2763406, 
    0.2763406, 0.2763406, 0.2763406, 0.271569, 0.271569, 0.271569, 0.271569, 
    0.271569, 0.271569, 0.271569, 0.2643491,
  0.3016985, 0.293511, 0.282592, 0.2704626, 0.2440143, 0.2444737, 0.2529599, 
    0.2482225, 0.2448359, 0.2364043, 0.222544, 0.2162489, 0.2112859, 
    0.2037814, 0.1624362, 0.1348797, 0.1418017, 0.1724503, 0.2369255, 
    0.2680533, 0.3004127, 0.3151629, 0.2363587, 0.1799467, 0.1802451, 
    0.2098549, 0.2365231, 0.2720884, 0.2940034,
  0.2196669, 0.1845451, 0.1713288, 0.1887959, 0.2261702, 0.1983253, 
    0.1701694, 0.1978544, 0.189233, 0.1874725, 0.203249, 0.2018961, 
    0.1859385, 0.1550673, 0.1698541, 0.2017773, 0.1866301, 0.1854411, 
    0.1935236, 0.1973951, 0.2074009, 0.2830505, 0.3405721, 0.5320673, 
    0.4893391, 0.5542788, 0.4843939, 0.4531281, 0.3068564,
  0.694625, 0.522735, 0.465243, 0.4435947, 0.3929487, 0.3290735, 0.2765031, 
    0.2334038, 0.211251, 0.1862545, 0.2005943, 0.2622854, 0.4643226, 
    0.8374498, 0.8821031, 0.9453111, 0.7974671, 0.6535266, 0.4525589, 
    0.3520955, 0.3445022, 0.3086195, 0.3967634, 1.027511, 2.732824, 2.345578, 
    1.72839, 1.266995, 0.894883,
  1.157982, 0.8596433, 0.8540243, 0.9059428, 0.6828794, 0.5338032, 0.4569092, 
    0.3704274, 0.3180842, 0.282437, 0.3585025, 1.003089, 2.01184, 1.890693, 
    3.041364, 1.855657, 1.122574, 0.7617432, 0.6056296, 0.4836012, 0.4025551, 
    0.3179316, 0.4799087, 10.64109, 10.00797, 5.582157, 3.521964, 2.214328, 
    1.476038,
  1.240048, 1.167403, 2.493896, 1.840789, 1.026938, 0.7351165, 0.5500361, 
    0.4882198, 0.4187377, 0.5073674, 2.21312, 4.455188, 8.517133, 3.105235, 
    9.823333, 1.694084, 0.9711002, 0.7262396, 0.6403304, 0.5328646, 
    0.4274895, 0.3436127, 0.3274735, 15.7894, 22.85542, 7.042305, 2.815544, 
    1.855865, 1.423654,
  0.9750468, 5.043158, 35.09755, 5.057478, 1.674254, 0.7601942, 0.5983403, 
    0.6017339, 0.9069067, 12.41976, 28.95737, 32.60043, 24.82318, 3.722513, 
    1.91722, 1.09381, 0.7292337, 0.5790347, 0.4782935, 0.4355688, 0.3665451, 
    0.303228, 0.5032619, 26.38363, 38.40689, 9.520375, 2.201871, 1.43719, 
    1.083046,
  2.242319, 31.67682, 40.57703, 9.943361, 2.350475, 0.823185, 0.930521, 
    1.761703, 4.964942, 23.66951, 42.43407, 34.55591, 6.655594, 2.145237, 
    1.239172, 0.6155033, 0.4735352, 0.4281044, 0.3792526, 0.3124204, 
    0.3176592, 0.4228174, 1.075869, 9.830962, 44.9603, 32.32659, 1.530391, 
    0.8107896, 1.030217,
  4.799612, 22.98452, 38.57047, 18.60074, 1.683764, 1.251273, 1.475313, 
    3.171221, 6.735636, 11.36989, 15.19903, 6.96986, 3.249516, 0.6043499, 
    0.3786812, 0.3999646, 0.5012658, 0.5322401, 0.5918518, 0.6854553, 
    0.704837, 0.8657155, 2.731326, 44.18441, 38.85273, 28.78142, 2.517851, 
    1.555842, 2.177611,
  16.80425, 46.16981, 48.87495, 25.95897, 4.67197, 4.150812, 4.538848, 
    4.072289, 13.62669, 22.17964, 5.161646, 2.103071, 0.4824174, 0.3476226, 
    0.4324462, 0.619575, 0.8806391, 1.299013, 1.852477, 2.385837, 2.823227, 
    3.755303, 8.894305, 39.80634, 30.42128, 10.58171, 8.070773, 10.81067, 
    12.4591,
  48.05335, 50.90022, 47.57715, 34.80349, 21.44329, 11.48286, 19.5161, 
    12.39084, 22.22829, 7.605733, 5.880725, 1.5434, 0.8389134, 0.8273237, 
    0.9088133, 0.9977776, 1.296973, 1.972613, 2.66253, 3.743113, 6.659698, 
    12.28185, 9.525347, 19.84488, 3.99501, 5.476301, 10.39619, 23.11969, 
    49.25538,
  46.41351, 49.18454, 44.78851, 31.16456, 43.5715, 20.87883, 39.54539, 
    40.26649, 46.97399, 25.81751, 8.555178, 4.982316, 3.207499, 2.696949, 
    2.380386, 2.268211, 2.44004, 2.58385, 4.943064, 8.700827, 13.85678, 
    22.24865, 8.803237, 5.695571, 3.08745, 3.884266, 6.095516, 18.85947, 
    46.70704,
  42.36744, 37.30142, 29.82127, 41.63532, 41.14122, 50.35406, 52.93012, 
    39.29904, 49.2064, 62.80188, 22.1935, 11.87973, 7.695091, 5.860933, 
    4.383943, 3.788769, 3.396505, 2.872768, 4.526447, 14.43567, 33.28885, 
    36.71714, 33.42492, 11.46609, 6.488932, 4.810145, 4.686534, 7.855852, 
    34.38344,
  27.79109, 26.37812, 37.9346, 40.35255, 56.83127, 60.32638, 49.41063, 
    63.50257, 61.89266, 54.48797, 51.17472, 30.3849, 16.07142, 9.963263, 
    7.637814, 5.968881, 4.78069, 4.247889, 4.562441, 26.67672, 35.55798, 
    53.86489, 56.56631, 44.2982, 19.39226, 10.91021, 7.945294, 7.477545, 
    18.33268,
  19.99486, 37.41525, 50.65642, 54.93892, 58.73751, 61.90047, 54.61806, 
    35.91547, 47.68673, 63.45285, 74.89503, 66.20158, 27.83023, 17.78855, 
    13.13605, 9.746582, 8.311031, 8.036567, 9.628102, 27.97118, 48.90761, 
    62.28971, 64.12913, 59.64621, 44.56046, 19.85616, 10.89639, 8.325406, 
    10.55991,
  12.45895, 29.35383, 38.74793, 47.69278, 50.99899, 57.30144, 59.58133, 
    59.54703, 52.76276, 59.93537, 57.23224, 43.3834, 29.43277, 29.06728, 
    21.89334, 16.87856, 22.05182, 22.07954, 30.36628, 43.65044, 52.21376, 
    43.9899, 29.71479, 32.65876, 23.17162, 11.28761, 9.81911, 8.56704, 
    9.018302,
  9.076964, 13.58665, 18.43188, 22.17241, 24.14632, 26.47982, 29.54466, 
    39.96362, 33.90247, 28.75212, 32.87341, 29.63046, 20.10747, 20.94269, 
    20.47297, 16.89709, 20.58788, 24.35205, 24.08049, 27.4092, 21.5813, 
    18.95022, 15.83864, 13.24093, 9.644037, 7.238731, 6.239749, 5.908748, 
    8.111526,
  8.250496, 9.176017, 10.44145, 11.46322, 12.26367, 12.20157, 12.79921, 
    13.90728, 14.5853, 14.38464, 14.40241, 13.95728, 12.7167, 11.53021, 
    10.70857, 9.851741, 9.564271, 9.546189, 9.830907, 9.974317, 9.386044, 
    8.893042, 7.909238, 7.300377, 6.66262, 6.496212, 6.765296, 7.019972, 
    7.69917,
  0.2442631, 0.2442631, 0.2442631, 0.2442631, 0.2442631, 0.2442631, 
    0.2442631, 0.2490955, 0.2490955, 0.2490955, 0.2490955, 0.2490955, 
    0.2490955, 0.2490955, 0.2573162, 0.2573162, 0.2573162, 0.2573162, 
    0.2573162, 0.2573162, 0.2573162, 0.2520863, 0.2520863, 0.2520863, 
    0.2520863, 0.2520863, 0.2520863, 0.2520863, 0.2442631,
  0.2845521, 0.2755138, 0.2682624, 0.2565975, 0.2354496, 0.2365731, 
    0.2435335, 0.2381813, 0.235246, 0.2277571, 0.2184247, 0.2139565, 
    0.2123824, 0.2064091, 0.1641393, 0.1362659, 0.1435797, 0.1706015, 
    0.23475, 0.2522439, 0.2767163, 0.2799444, 0.2267375, 0.1822033, 
    0.1764432, 0.2008453, 0.2282802, 0.2573938, 0.2770554,
  0.2130943, 0.1845802, 0.1713609, 0.1892311, 0.2154074, 0.1920687, 
    0.1723012, 0.1916338, 0.1858525, 0.1853275, 0.1961021, 0.1909401, 
    0.1836102, 0.1543572, 0.1602582, 0.1914191, 0.1800863, 0.1783192, 
    0.1838466, 0.1901261, 0.1994722, 0.2713376, 0.3276335, 0.4963643, 
    0.4548014, 0.5308458, 0.4646198, 0.4336406, 0.2915112,
  0.6686062, 0.5045678, 0.4522541, 0.426893, 0.3776823, 0.3219377, 0.2719112, 
    0.2299677, 0.2079996, 0.1825128, 0.1964977, 0.2523297, 0.4501525, 
    0.8304835, 0.8701287, 0.9263296, 0.7980114, 0.6442166, 0.4441001, 
    0.3465557, 0.3407026, 0.3072058, 0.3935611, 1.078036, 2.926662, 2.469647, 
    1.737478, 1.250399, 0.8712059,
  1.143562, 0.848701, 0.8502575, 0.8850291, 0.6533093, 0.5124496, 0.4457095, 
    0.3669247, 0.3145007, 0.2800192, 0.3561922, 0.9962593, 1.974872, 
    1.884087, 3.226934, 1.820593, 1.102478, 0.7461961, 0.5994248, 0.4795814, 
    0.3993012, 0.315147, 0.4930993, 13.27955, 10.57006, 5.656201, 3.530576, 
    2.189503, 1.450294,
  1.227157, 1.161661, 2.47975, 1.800521, 0.9966208, 0.724218, 0.5428469, 
    0.4855393, 0.4144182, 0.4912384, 2.195136, 4.566549, 8.570848, 3.050004, 
    11.53439, 1.675934, 0.9665781, 0.7173855, 0.6331491, 0.5275934, 
    0.4253227, 0.3423531, 0.3261278, 19.305, 25.24659, 6.955924, 2.758103, 
    1.832086, 1.409048,
  0.9730382, 4.804256, 38.17801, 4.943917, 1.627471, 0.7516205, 0.59411, 
    0.5992448, 0.8993733, 12.51471, 31.64779, 35.43675, 27.67084, 3.679955, 
    1.912542, 1.092363, 0.723626, 0.5769466, 0.4757033, 0.4353296, 0.3667848, 
    0.3032187, 0.5032059, 29.81352, 41.777, 9.398008, 2.181621, 1.419168, 
    1.077883,
  2.213135, 35.71336, 43.41652, 9.950487, 2.322968, 0.8216015, 0.926236, 
    1.753382, 4.963067, 23.91445, 45.46107, 37.33237, 6.622656, 2.143993, 
    1.257941, 0.6162779, 0.4733815, 0.4278524, 0.3791607, 0.3123835, 
    0.3174078, 0.4225868, 1.075499, 10.49084, 47.02365, 34.94173, 1.508553, 
    0.8089787, 1.027344,
  4.801159, 24.28588, 40.15673, 20.64186, 1.682153, 1.250983, 1.47321, 
    3.170548, 6.742768, 11.40949, 15.32809, 7.022104, 3.520433, 0.6054746, 
    0.3789371, 0.4000733, 0.5014858, 0.5322382, 0.5905113, 0.6816898, 
    0.6993802, 0.8617557, 2.72129, 44.70964, 39.72011, 31.43259, 2.571301, 
    1.551215, 2.174532,
  16.76193, 45.93644, 48.70198, 27.2836, 4.69647, 4.155569, 4.546992, 
    4.078472, 14.37952, 22.58894, 5.189811, 2.109034, 0.4819297, 0.3474007, 
    0.4321623, 0.6190145, 0.8799077, 1.291093, 1.826091, 2.325722, 2.698739, 
    3.504353, 8.50903, 40.85594, 32.67306, 10.59282, 8.082343, 10.78928, 
    12.41054,
  49.66207, 53.17601, 50.01976, 36.83646, 22.49999, 11.49423, 20.21962, 
    12.4145, 22.82363, 7.650722, 6.023122, 1.545267, 0.8401829, 0.8297797, 
    0.9117902, 1.000047, 1.303107, 1.97901, 2.670545, 3.752184, 6.675849, 
    12.43203, 10.61414, 21.06849, 3.995095, 5.475249, 10.38924, 23.19658, 
    50.78331,
  48.88456, 52.60881, 47.72124, 32.3453, 46.22695, 20.58646, 42.70724, 
    40.88209, 50.82856, 26.18539, 8.578051, 5.003986, 3.213006, 2.70119, 
    2.384977, 2.273526, 2.444671, 2.595382, 4.972872, 9.100073, 14.91918, 
    23.55323, 8.826933, 5.886493, 3.08809, 3.880523, 6.086035, 18.4446, 
    49.6424,
  45.94132, 39.94695, 31.67689, 44.73713, 43.63325, 54.35427, 57.85082, 
    42.9348, 53.18973, 67.66798, 22.39507, 11.89561, 7.722994, 5.890955, 
    4.393888, 3.791167, 3.404515, 2.878716, 4.553942, 15.82182, 36.79464, 
    39.72989, 36.15262, 11.47208, 6.510838, 4.821714, 4.690066, 7.932489, 
    37.29792,
  30.49655, 27.06033, 40.06604, 43.66753, 63.81428, 65.49863, 53.12622, 
    70.64916, 67.20238, 58.51936, 54.52211, 30.98069, 16.11649, 10.04932, 
    7.62325, 5.961549, 4.777283, 4.249726, 4.573428, 30.96002, 40.47166, 
    58.87488, 61.41687, 45.59372, 19.3518, 10.92151, 7.962541, 7.512059, 
    20.45152,
  22.19171, 41.76133, 55.97446, 61.89213, 68.41628, 72.07244, 62.20905, 
    40.12724, 53.68941, 70.28386, 81.20641, 73.88564, 27.93602, 17.89378, 
    13.02266, 9.733407, 8.320027, 8.080949, 9.850144, 32.81764, 54.41109, 
    68.32799, 68.91396, 65.32973, 47.61218, 19.88543, 10.86797, 8.30469, 
    10.80731,
  12.74225, 33.22576, 42.84715, 55.28764, 58.32862, 64.5131, 67.89245, 
    69.64541, 62.3534, 70.05305, 65.70584, 50.68496, 34.34072, 33.76251, 
    22.34714, 18.16309, 26.51365, 25.08416, 36.77216, 51.41602, 59.84602, 
    51.79141, 32.19328, 36.81675, 23.43996, 11.27632, 9.829627, 8.56181, 
    9.009967,
  9.166538, 13.77402, 20.65789, 22.84224, 26.59957, 30.58219, 33.73346, 
    45.88122, 37.70385, 31.91364, 37.27285, 35.0674, 23.73523, 26.28537, 
    23.60791, 18.53409, 22.62813, 27.20932, 26.90788, 30.89677, 24.2497, 
    21.08018, 17.48003, 14.74078, 10.02557, 7.223883, 6.204144, 5.784432, 
    8.077038,
  8.157644, 9.176674, 10.57721, 11.75637, 12.74239, 12.72764, 13.21354, 
    14.25893, 14.859, 15.02844, 15.48285, 14.8717, 13.48862, 12.28891, 
    11.52114, 10.39103, 9.916151, 9.974962, 10.23322, 10.0488, 9.604025, 
    8.85449, 7.864571, 7.217093, 6.627211, 6.438487, 6.743498, 6.931252, 
    7.637196,
  0.2307505, 0.2307505, 0.2307505, 0.2307505, 0.2307505, 0.2307505, 
    0.2307505, 0.2341864, 0.2341864, 0.2341864, 0.2341864, 0.2341864, 
    0.2341864, 0.2341864, 0.2406562, 0.2406562, 0.2406562, 0.2406562, 
    0.2406562, 0.2406562, 0.2406562, 0.2372798, 0.2372798, 0.2372798, 
    0.2372798, 0.2372798, 0.2372798, 0.2372798, 0.2307505,
  0.2721483, 0.2620395, 0.2559921, 0.2473681, 0.231021, 0.2299041, 0.2348589, 
    0.2300058, 0.2287845, 0.2229038, 0.2151391, 0.2117721, 0.212258, 
    0.2079576, 0.167641, 0.1384561, 0.1457674, 0.1705901, 0.2355242, 
    0.2397843, 0.2578338, 0.2543192, 0.2211365, 0.1838866, 0.1745167, 
    0.1939287, 0.2253332, 0.2491345, 0.2668526,
  0.2097925, 0.1853456, 0.1725853, 0.1904367, 0.2074505, 0.1887092, 
    0.1736482, 0.1876695, 0.1850744, 0.1844356, 0.192215, 0.1840034, 
    0.1824706, 0.1551982, 0.1545711, 0.1843024, 0.1754508, 0.175335, 
    0.1777095, 0.1824564, 0.1937699, 0.2649812, 0.3211338, 0.4722159, 
    0.436038, 0.5186306, 0.4565465, 0.4185806, 0.2835163,
  0.6543143, 0.495061, 0.4466186, 0.4164368, 0.3698861, 0.3183144, 0.2691431, 
    0.2281696, 0.2058442, 0.1803759, 0.1939144, 0.2505511, 0.4421153, 
    0.8271077, 0.8658764, 0.9186561, 0.7969797, 0.633408, 0.4385783, 
    0.3444596, 0.3387897, 0.3063619, 0.3924302, 1.105178, 3.099497, 2.551893, 
    1.734439, 1.230443, 0.853146,
  1.134396, 0.8417563, 0.8546747, 0.8723739, 0.6397885, 0.5049752, 0.4404763, 
    0.3655593, 0.3124936, 0.2785411, 0.3570968, 0.9888831, 1.953141, 
    1.881112, 3.372238, 1.795137, 1.092622, 0.7402561, 0.5960183, 0.4779192, 
    0.3980738, 0.3141696, 0.4985252, 16.17471, 10.86156, 5.666274, 3.558796, 
    2.159978, 1.433342,
  1.220395, 1.159148, 2.464881, 1.780426, 0.9828619, 0.7197699, 0.539625, 
    0.4842893, 0.4128428, 0.4793087, 2.186166, 4.633715, 8.630954, 3.017523, 
    13.6222, 1.662869, 0.9640666, 0.7133189, 0.6298803, 0.5260814, 0.4241472, 
    0.341036, 0.3255411, 23.37931, 27.92474, 6.900717, 2.736148, 1.821785, 
    1.403085,
  0.9722143, 4.759559, 42.76807, 4.892202, 1.604885, 0.749153, 0.5927814, 
    0.5982779, 0.8970864, 12.5601, 35.26093, 39.41751, 31.7205, 3.663549, 
    1.909651, 1.090937, 0.7215973, 0.5762443, 0.4747329, 0.4352286, 
    0.3668703, 0.3032684, 0.5031263, 32.41614, 46.31416, 9.356019, 2.173025, 
    1.410716, 1.075609,
  2.205584, 40.26591, 47.56403, 9.961478, 2.32129, 0.8210768, 0.9246802, 
    1.750531, 4.963274, 24.08717, 50.35014, 41.5679, 6.629036, 2.144084, 
    1.261983, 0.6164567, 0.4732991, 0.4278094, 0.3791188, 0.3123793, 
    0.3173146, 0.4224218, 1.075626, 10.77156, 51.04208, 38.57246, 1.501281, 
    0.8084114, 1.026725,
  4.801605, 26.17433, 43.9122, 23.49714, 1.681716, 1.251046, 1.472633, 
    3.170271, 6.743998, 11.42398, 15.38778, 7.038903, 3.820407, 0.6059379, 
    0.3790525, 0.4000891, 0.5015461, 0.5322238, 0.5901285, 0.6806046, 
    0.6975007, 0.8604807, 2.719218, 46.37738, 41.93864, 35.7075, 2.604082, 
    1.549964, 2.173472,
  16.74723, 47.23307, 50.92859, 29.03879, 4.701005, 4.157592, 4.549456, 
    4.080575, 16.30539, 24.03987, 5.198709, 2.110796, 0.4817965, 0.3473371, 
    0.432115, 0.6189821, 0.8796303, 1.287713, 1.817929, 2.301643, 2.651823, 
    3.418882, 8.40175, 43.12578, 36.38548, 10.60065, 8.083958, 10.78467, 
    12.39523,
  53.20177, 56.89572, 53.65863, 40.36754, 23.95234, 11.49911, 21.14645, 
    12.42111, 23.1233, 7.661971, 6.105141, 1.545876, 0.8406585, 0.8305471, 
    0.9125595, 1.00078, 1.304432, 1.98078, 2.673002, 3.755151, 6.681878, 
    12.48492, 12.04548, 22.96771, 3.996096, 5.475271, 10.38766, 23.21371, 
    54.30812,
  53.53635, 57.648, 52.22072, 33.66648, 50.62346, 20.5729, 47.15237, 
    41.39288, 55.37629, 26.36031, 8.584337, 5.011084, 3.215574, 2.703368, 
    2.386523, 2.27529, 2.446135, 2.599869, 4.982844, 9.223972, 15.23134, 
    25.42161, 8.836962, 6.033796, 3.088254, 3.879228, 6.086451, 18.4388, 
    54.64853,
  50.86277, 43.99709, 34.56647, 49.65578, 47.0602, 59.15334, 64.61275, 
    47.61825, 57.89359, 73.91151, 22.52959, 11.90405, 7.738724, 5.90632, 
    4.40008, 3.79127, 3.40728, 2.881305, 4.562013, 16.82475, 41.22019, 
    43.62865, 39.76428, 11.47141, 6.518471, 4.825387, 4.691685, 7.967182, 
    41.36954,
  33.79115, 27.86503, 42.66955, 47.26025, 73.88573, 71.35648, 57.94695, 
    79.41269, 73.4164, 62.90287, 58.70834, 31.45111, 16.13362, 10.06651, 
    7.622897, 5.960462, 4.776524, 4.249005, 4.569726, 36.24068, 46.89374, 
    64.93649, 66.51282, 46.62876, 19.32009, 10.91981, 7.965252, 7.520266, 
    22.94987,
  24.14087, 46.44578, 61.85587, 69.57056, 80.4859, 84.66242, 71.14125, 
    45.28899, 61.30563, 76.95029, 87.64043, 81.44913, 27.82504, 17.8309, 
    12.93647, 9.707659, 8.341591, 8.098418, 9.954004, 38.58929, 60.62821, 
    74.31459, 73.98592, 71.16892, 50.03777, 19.82559, 10.856, 8.300155, 
    10.96323,
  12.92136, 37.71401, 46.01814, 63.47174, 65.86366, 71.868, 76.90226, 
    79.61608, 73.35751, 79.67065, 73.43864, 59.43943, 41.07576, 38.61901, 
    22.62798, 18.97889, 31.72805, 28.54455, 44.37355, 59.98322, 66.8103, 
    59.32022, 33.93404, 41.59402, 23.5567, 11.29764, 9.811057, 8.560516, 
    9.011073,
  9.200273, 13.87483, 23.35086, 23.23434, 28.65062, 34.59712, 38.96511, 
    51.89555, 42.23758, 36.24895, 41.42503, 41.46037, 28.65539, 32.92535, 
    26.32924, 19.74204, 24.84033, 29.6723, 29.79158, 34.10799, 27.74887, 
    24.01814, 19.10072, 16.6678, 10.27584, 7.182191, 6.147606, 5.694842, 
    8.007338,
  8.077063, 9.082121, 10.51815, 11.7718, 12.98189, 12.9727, 13.71138, 
    14.56839, 15.05814, 15.5995, 16.1771, 15.45149, 13.9949, 12.76036, 
    11.9274, 10.65622, 10.05336, 10.04949, 10.35922, 10.05087, 9.538676, 
    8.792247, 7.816166, 7.175088, 6.588481, 6.409289, 6.692918, 6.809655, 
    7.55153,
  0.2229644, 0.2229644, 0.2229644, 0.2229644, 0.2229644, 0.2229644, 
    0.2229644, 0.2251064, 0.2251064, 0.2251064, 0.2251064, 0.2251064, 
    0.2251064, 0.2251064, 0.2294156, 0.2294156, 0.2294156, 0.2294156, 
    0.2294156, 0.2294156, 0.2294156, 0.2280707, 0.2280707, 0.2280707, 
    0.2280707, 0.2280707, 0.2280707, 0.2280707, 0.2229644,
  0.2615055, 0.252426, 0.2467369, 0.2413559, 0.2273554, 0.2248869, 0.2277238, 
    0.2241565, 0.2243886, 0.2199245, 0.2128755, 0.2105571, 0.2108302, 
    0.2083814, 0.1720622, 0.141933, 0.145369, 0.1717467, 0.2359186, 
    0.2306772, 0.2475731, 0.2381476, 0.2180948, 0.1845524, 0.1726346, 
    0.1871214, 0.2234051, 0.2464673, 0.2597576,
  0.2086735, 0.1865734, 0.1734419, 0.1916071, 0.2016349, 0.1864974, 
    0.1743776, 0.1851769, 0.1851224, 0.1837085, 0.1900722, 0.1809182, 
    0.1824436, 0.1566402, 0.1515034, 0.1798075, 0.1728203, 0.1735661, 
    0.1741909, 0.1789999, 0.190325, 0.2612713, 0.3183487, 0.4590261, 
    0.426191, 0.5144891, 0.4518674, 0.4088362, 0.2793127,
  0.6475858, 0.4901983, 0.4435346, 0.4109817, 0.3661477, 0.3169281, 
    0.2678117, 0.2271793, 0.2045647, 0.1793592, 0.1926733, 0.2519775, 
    0.4383364, 0.8237859, 0.8636225, 0.9137418, 0.7947533, 0.6248544, 
    0.4361158, 0.3435781, 0.3377416, 0.3059005, 0.3921409, 1.114438, 
    3.219143, 2.584606, 1.730131, 1.219084, 0.8442113,
  1.129045, 0.8384777, 0.8581974, 0.8591693, 0.6306199, 0.5008267, 0.4371226, 
    0.3649329, 0.3114291, 0.2778297, 0.3607547, 0.9842203, 1.941584, 
    1.878363, 3.449766, 1.782407, 1.087529, 0.7378305, 0.5946182, 0.477188, 
    0.3976136, 0.3136978, 0.4992313, 19.63541, 10.9321, 5.668878, 3.565145, 
    2.143225, 1.422525,
  1.21778, 1.158346, 2.44876, 1.770444, 0.9760146, 0.7173391, 0.5381134, 
    0.4835699, 0.4122145, 0.4724841, 2.18384, 4.643908, 8.673843, 3.004534, 
    16.39644, 1.655711, 0.9626881, 0.7114542, 0.6283508, 0.5254139, 
    0.4235553, 0.3399576, 0.3252519, 28.86942, 30.56138, 6.866554, 2.727376, 
    1.816778, 1.400031,
  0.9718251, 4.762699, 49.88491, 4.870266, 1.593903, 0.7480918, 0.5922825, 
    0.5978861, 0.8960862, 12.70954, 40.37471, 45.52423, 37.71677, 3.657403, 
    1.907704, 1.089916, 0.7208298, 0.5760086, 0.4743631, 0.4351842, 
    0.3669068, 0.3032617, 0.5031493, 34.89211, 52.62496, 9.335473, 2.169162, 
    1.40739, 1.074719,
  2.20328, 45.67025, 53.66142, 9.960332, 2.32287, 0.8208426, 0.9240527, 
    1.749279, 4.961886, 24.15638, 58.43063, 48.34913, 6.633132, 2.144215, 
    1.26316, 0.6164898, 0.4732586, 0.4277892, 0.3790881, 0.3123704, 
    0.3172751, 0.4223392, 1.075714, 10.78748, 58.35473, 44.20338, 1.498371, 
    0.808174, 1.026463,
  4.802001, 29.16982, 52.16343, 27.77816, 1.681503, 1.25107, 1.472428, 
    3.169937, 6.74438, 11.43164, 15.41038, 7.046052, 4.17843, 0.6061543, 
    0.3791077, 0.4001048, 0.5015739, 0.5322082, 0.589943, 0.6801146, 
    0.6966301, 0.8599504, 2.71835, 52.54335, 47.94888, 42.78827, 2.618559, 
    1.549579, 2.173088,
  16.74133, 52.7064, 57.19209, 31.65089, 4.702784, 4.158401, 4.550425, 
    4.081343, 20.93052, 28.64805, 5.20283, 2.111451, 0.4817527, 0.3472987, 
    0.4320875, 0.618949, 0.8795124, 1.286865, 1.814913, 2.291324, 2.632097, 
    3.390613, 8.368831, 48.96877, 43.21756, 10.60248, 8.084414, 10.78283, 
    12.3889,
  60.26757, 63.19623, 59.21339, 47.01686, 26.37012, 11.50157, 22.45862, 
    12.42413, 23.25304, 7.666084, 6.149155, 1.546123, 0.8408571, 0.8308858, 
    0.9128814, 1.001089, 1.304951, 1.981442, 2.673856, 3.7562, 6.684104, 
    12.50449, 14.24331, 26.1598, 3.996418, 5.475087, 10.38718, 23.21988, 
    61.4445,
  61.58297, 64.85516, 59.31705, 34.79095, 58.25336, 20.57292, 53.41419, 
    41.76694, 63.03841, 26.45251, 8.586965, 5.014298, 3.216777, 2.704369, 
    2.387154, 2.275966, 2.446814, 2.600989, 4.987166, 9.259679, 15.30576, 
    28.44116, 8.841784, 6.138971, 3.088328, 3.878706, 6.087268, 18.47668, 
    62.61224,
  58.5687, 50.10917, 39.44748, 57.29027, 52.65376, 65.78986, 74.59106, 
    54.23064, 63.89388, 82.62093, 22.61045, 11.90945, 7.745965, 5.912606, 
    4.40274, 3.790809, 3.408272, 2.882359, 4.56352, 17.49868, 48.05033, 
    49.40268, 45.9678, 11.47183, 6.522, 4.826836, 4.692408, 7.975768, 47.6288,
  37.70655, 28.76339, 45.86963, 52.15116, 90.6663, 79.2471, 65.15463, 
    89.74791, 81.80257, 68.92895, 64.49128, 31.85031, 16.12601, 10.06885, 
    7.621076, 5.959278, 4.776607, 4.247926, 4.56794, 44.14618, 55.83076, 
    72.82364, 72.82079, 47.46301, 19.30413, 10.92029, 7.965036, 7.522423, 
    25.78808,
  25.93696, 52.0267, 69.15015, 77.70049, 95.09373, 98.94605, 81.23865, 
    52.93361, 71.05386, 84.78801, 95.5616, 89.68114, 27.56954, 17.69669, 
    12.90756, 9.696734, 8.365468, 8.105645, 9.995383, 45.79205, 68.23225, 
    81.2048, 80.22776, 77.86752, 52.22695, 19.74064, 10.84602, 8.299188, 
    11.0378,
  13.0149, 43.08073, 48.84341, 71.21839, 74.28593, 78.87361, 84.77783, 
    87.96375, 84.68799, 88.91813, 82.35267, 70.14789, 49.40724, 43.69222, 
    22.81296, 19.32307, 38.32976, 32.41765, 53.72483, 69.8923, 73.32157, 
    66.21916, 34.67565, 48.15132, 23.56161, 11.32077, 9.805299, 8.559052, 
    9.011127,
  9.207272, 13.91587, 26.1278, 23.43554, 30.24006, 37.38028, 44.31575, 
    58.01603, 47.53588, 41.70114, 45.09977, 48.70671, 35.09812, 37.61543, 
    28.60045, 20.48058, 27.29844, 31.78716, 31.90705, 36.20235, 32.0663, 
    27.35967, 20.81257, 19.5955, 10.39491, 7.112965, 6.089464, 5.63928, 
    7.927695,
  8.016405, 9.010994, 10.48796, 11.78505, 12.99837, 12.89574, 13.86396, 
    14.50686, 14.98453, 15.83752, 16.24439, 15.34557, 13.90995, 12.83872, 
    11.90238, 10.65807, 10.12914, 9.988202, 10.2948, 9.934958, 9.31484, 
    8.649586, 7.754925, 7.122393, 6.552009, 6.381419, 6.616971, 6.718473, 
    7.506337,
  0.2186493, 0.2186493, 0.2186493, 0.2186493, 0.2186493, 0.2186493, 
    0.2186493, 0.2215753, 0.2215753, 0.2215753, 0.2215753, 0.2215753, 
    0.2215753, 0.2215753, 0.2250614, 0.2250614, 0.2250614, 0.2250614, 
    0.2250614, 0.2250614, 0.2250614, 0.2228733, 0.2228733, 0.2228733, 
    0.2228733, 0.2228733, 0.2228733, 0.2228733, 0.2186493,
  0.2546053, 0.2472809, 0.2415814, 0.2364997, 0.223862, 0.221507, 0.2234758, 
    0.2207617, 0.2214115, 0.2179353, 0.2112535, 0.2096095, 0.2094006, 
    0.2084104, 0.1743602, 0.1445485, 0.1450306, 0.1739658, 0.2353456, 
    0.2264666, 0.2416028, 0.2298994, 0.2165019, 0.1844895, 0.1705948, 
    0.1820791, 0.2212182, 0.2460271, 0.2566295,
  0.2081207, 0.1875367, 0.1737199, 0.1923433, 0.1984612, 0.1850028, 
    0.1749556, 0.1842494, 0.1850787, 0.1834719, 0.1895187, 0.179679, 
    0.1824238, 0.1575903, 0.149915, 0.1772317, 0.1712542, 0.1723951, 
    0.1727342, 0.1777103, 0.188526, 0.2592587, 0.3153193, 0.452683, 
    0.4197682, 0.5105294, 0.4498671, 0.4034345, 0.2768214,
  0.6441337, 0.4878475, 0.4414714, 0.4085897, 0.3641728, 0.3161407, 
    0.2669555, 0.2266299, 0.2038585, 0.178906, 0.1922801, 0.2525066, 
    0.4353937, 0.8198634, 0.8626176, 0.9109139, 0.792703, 0.6189784, 
    0.4345716, 0.3430121, 0.3371531, 0.3056301, 0.3919799, 1.117313, 3.28774, 
    2.591136, 1.721901, 1.211815, 0.8386916,
  1.125621, 0.836571, 0.8608094, 0.8457114, 0.6254795, 0.4974293, 0.4346535, 
    0.3645542, 0.3107667, 0.2774278, 0.3616572, 0.9812635, 1.93366, 1.876022, 
    3.473949, 1.775367, 1.084609, 0.7365685, 0.5940413, 0.476878, 0.3973219, 
    0.3133864, 0.4991142, 24.40879, 10.92205, 5.647262, 3.552174, 2.131525, 
    1.415521,
  1.216423, 1.157983, 2.436449, 1.764993, 0.9725251, 0.7158557, 0.5372266, 
    0.4831421, 0.4118923, 0.4694361, 2.180882, 4.645805, 8.683422, 2.997772, 
    20.7263, 1.652058, 0.9619317, 0.7105079, 0.6275741, 0.5251295, 0.4233119, 
    0.3393495, 0.3250686, 38.18661, 32.40263, 6.847047, 2.722886, 1.813963, 
    1.39825,
  0.9715969, 4.756264, 63.13066, 4.861345, 1.588667, 0.7476015, 0.5920292, 
    0.597675, 0.8955824, 12.80578, 48.65623, 55.84777, 48.24639, 3.654569, 
    1.906898, 1.089591, 0.7205055, 0.5758791, 0.4741775, 0.4351481, 
    0.3669235, 0.3032485, 0.5031621, 37.62973, 62.64931, 9.322537, 2.167306, 
    1.406005, 1.074305,
  2.202202, 53.74871, 64.62136, 9.95806, 2.323667, 0.8207083, 0.9237196, 
    1.748593, 4.96072, 24.16308, 70.9837, 59.80415, 6.634441, 2.144237, 
    1.263525, 0.6165282, 0.4732279, 0.42777, 0.3790649, 0.3123615, 0.317252, 
    0.42229, 1.075768, 10.77785, 73.44, 54.7462, 1.496998, 0.8080448, 1.02632,
  4.802247, 35.28176, 69.92925, 34.89151, 1.681349, 1.251068, 1.472304, 
    3.169657, 6.744471, 11.43638, 15.42388, 7.049798, 4.600931, 0.6062595, 
    0.3791294, 0.4001093, 0.5015796, 0.5321892, 0.58983, 0.6798265, 0.696133, 
    0.859664, 2.717874, 69.88026, 63.25959, 55.58895, 2.626567, 1.54934, 
    2.172894,
  16.73882, 71.70437, 75.93913, 35.99635, 4.703521, 4.158733, 4.550887, 
    4.081649, 34.96244, 44.89287, 5.205221, 2.111777, 0.4817264, 0.3472801, 
    0.4320696, 0.6189196, 0.8794347, 1.286522, 1.813604, 2.286923, 2.62344, 
    3.381161, 8.356649, 64.10147, 57.16896, 10.6014, 8.084497, 10.78187, 
    12.38586,
  75.62, 76.25989, 69.80168, 60.96043, 30.63579, 11.50297, 24.98492, 
    12.42548, 23.32318, 7.667994, 6.17361, 1.546255, 0.84096, 0.8310593, 
    0.9130383, 1.001239, 1.305151, 1.981707, 2.674219, 3.756583, 6.685132, 
    12.51285, 19.2108, 30.86409, 3.996471, 5.47492, 10.38701, 23.22306, 
    78.34577,
  77.43043, 76.7947, 72.70758, 35.36396, 73.43124, 20.56703, 64.00452, 
    41.93524, 77.12669, 26.50347, 8.588246, 5.015929, 3.217396, 2.704874, 
    2.387488, 2.276283, 2.447113, 2.601453, 4.989159, 9.268361, 15.31986, 
    34.12655, 8.844466, 6.203157, 3.088346, 3.878384, 6.087458, 18.48292, 
    78.06009,
  73.73637, 61.82753, 49.48962, 70.69184, 63.99373, 77.60335, 89.72005, 
    64.77694, 73.47461, 97.00121, 22.63309, 11.91282, 7.749022, 5.91482, 
    4.403829, 3.790369, 3.408542, 2.88277, 4.563971, 17.70387, 61.70477, 
    57.83522, 57.5024, 11.47183, 6.523553, 4.827504, 4.692712, 7.977762, 
    59.61556,
  42.71867, 29.51159, 50.00597, 60.76216, 119.7086, 91.58904, 80.20596, 
    104.4863, 96.07129, 78.67876, 74.5344, 32.08748, 16.12014, 10.06931, 
    7.620382, 5.958332, 4.776248, 4.246809, 4.568531, 58.03792, 70.15143, 
    83.8474, 81.77579, 48.26873, 19.29548, 10.92116, 7.965022, 7.522986, 
    28.92578,
  27.61691, 59.65921, 78.84479, 87.83649, 110.6305, 114.8139, 94.3387, 
    69.47002, 84.43937, 95.78493, 106.8222, 100.297, 27.39799, 17.63576, 
    12.8819, 9.692119, 8.372313, 8.105747, 9.997209, 55.95961, 78.78628, 
    90.23605, 88.82954, 85.90729, 54.50065, 19.7014, 10.83688, 8.297532, 
    11.08294,
  13.06531, 49.4738, 51.86953, 77.34027, 82.42622, 85.18125, 91.62773, 
    94.8835, 94.51067, 97.94376, 91.73063, 82.58432, 59.0885, 48.46012, 
    22.8816, 19.40179, 45.36361, 37.25418, 64.59168, 81.25232, 79.47374, 
    73.28149, 34.75749, 57.75922, 23.54068, 11.33392, 9.806612, 8.556992, 
    9.010554,
  9.207324, 13.92863, 28.56002, 23.53951, 30.69762, 38.68145, 47.67991, 
    64.91161, 53.25886, 45.7672, 47.75529, 54.28667, 40.46976, 40.01307, 
    30.26431, 20.75385, 29.7399, 33.43459, 32.93195, 37.24878, 36.87843, 
    30.5428, 23.35666, 24.61692, 10.37281, 7.043863, 6.027721, 5.599058, 
    7.885869,
  7.999473, 8.995122, 10.47385, 11.76705, 12.93873, 12.78726, 13.84777, 
    14.34147, 14.83237, 15.8253, 16.05888, 15.08355, 13.66677, 12.68406, 
    11.80746, 10.67105, 10.06585, 9.814538, 10.14765, 9.757403, 9.119962, 
    8.54318, 7.681246, 7.05063, 6.503006, 6.343224, 6.523269, 6.631657, 
    7.480544,
  0.216563, 0.216563, 0.216563, 0.216563, 0.216563, 0.216563, 0.216563, 
    0.2205283, 0.2205283, 0.2205283, 0.2205283, 0.2205283, 0.2205283, 
    0.2205283, 0.2238842, 0.2238842, 0.2238842, 0.2238842, 0.2238842, 
    0.2238842, 0.2238842, 0.2205292, 0.2205292, 0.2205292, 0.2205292, 
    0.2205292, 0.2205292, 0.2205292, 0.216563,
  0.2524069, 0.2451792, 0.2395649, 0.2343972, 0.2217905, 0.2207001, 
    0.2217827, 0.2194007, 0.219594, 0.216723, 0.2108909, 0.209069, 0.2082332, 
    0.2081482, 0.1747936, 0.145895, 0.145279, 0.1750837, 0.2343171, 
    0.2248166, 0.2392324, 0.2273562, 0.2158087, 0.1842353, 0.1695205, 
    0.1796106, 0.2194759, 0.2455004, 0.2558319,
  0.2073721, 0.1877323, 0.1737692, 0.1925925, 0.1971661, 0.184581, 0.1752167, 
    0.1839336, 0.1850288, 0.1832698, 0.1892919, 0.1794109, 0.1822971, 
    0.1581374, 0.1490366, 0.1757766, 0.1704559, 0.171994, 0.1721481, 
    0.1772277, 0.1876494, 0.2582511, 0.31308, 0.4507427, 0.4152432, 
    0.5078963, 0.4484548, 0.4007315, 0.2753696,
  0.6420603, 0.4866797, 0.4401959, 0.4073668, 0.3631154, 0.3157421, 
    0.2663634, 0.2262794, 0.2034487, 0.178651, 0.1922281, 0.2520312, 
    0.4328296, 0.8157046, 0.8618873, 0.9084169, 0.7912288, 0.615002, 
    0.4332762, 0.3426002, 0.33686, 0.3054981, 0.3919589, 1.119571, 3.306999, 
    2.587558, 1.713907, 1.205954, 0.8354738,
  1.122881, 0.8353241, 0.8634856, 0.8319725, 0.6218821, 0.4954777, 0.4329431, 
    0.3642792, 0.3103457, 0.2771856, 0.3613695, 0.9789739, 1.927017, 
    1.875537, 3.481615, 1.770088, 1.082832, 0.7358288, 0.5937636, 0.4766413, 
    0.3971158, 0.3131881, 0.4988431, 32.58699, 10.90181, 5.615352, 3.530024, 
    2.124356, 1.411667,
  1.215588, 1.15793, 2.428363, 1.761688, 0.9704771, 0.7148801, 0.5367085, 
    0.4828595, 0.4117029, 0.4680635, 2.179122, 4.645604, 8.670521, 2.994136, 
    28.11686, 1.650199, 0.9615349, 0.709958, 0.6270943, 0.5250538, 0.4231917, 
    0.3389717, 0.3249684, 54.44349, 33.14612, 6.834514, 2.720111, 1.812225, 
    1.397064,
  0.9714519, 4.749606, 92.09241, 4.857379, 1.585843, 0.7473491, 0.5918913, 
    0.5975436, 0.8953038, 12.82399, 62.83666, 77.25015, 69.87774, 3.653045, 
    1.90652, 1.089474, 0.7203339, 0.5757815, 0.4740694, 0.4351164, 0.3669297, 
    0.3032362, 0.5031684, 40.079, 81.31528, 9.315841, 2.166384, 1.405461, 
    1.074092,
  2.201618, 66.07259, 87.21333, 9.95628, 2.323403, 0.8206257, 0.9235309, 
    1.748183, 4.959966, 24.16279, 92.10706, 83.12334, 6.634991, 2.144189, 
    1.263629, 0.6165466, 0.473207, 0.4277551, 0.3790487, 0.3123533, 
    0.3172369, 0.4222615, 1.075795, 10.77141, 106.4174, 76.8311, 1.496316, 
    0.8079748, 1.026235,
  4.802342, 48.00142, 111.3946, 47.25619, 1.681241, 1.251051, 1.472212, 
    3.169438, 6.744383, 11.44017, 15.43207, 7.051704, 5.197432, 0.6063113, 
    0.3791367, 0.4001072, 0.5015765, 0.5321701, 0.5897604, 0.6796677, 
    0.6958747, 0.8595164, 2.717599, 122.1879, 103.167, 80.7794, 2.630607, 
    1.549183, 2.172761,
  16.73752, 131.739, 131.7418, 42.38957, 4.703765, 4.158854, 4.551073, 
    4.081752, 72.45839, 88.9796, 5.207471, 2.11194, 0.4817106, 0.3472662, 
    0.4320526, 0.6188879, 0.8793712, 1.286332, 1.812994, 2.285268, 2.620396, 
    3.377972, 8.351719, 99.04272, 87.92728, 10.59983, 8.084364, 10.78122, 
    12.38415,
  108.3639, 101.9707, 86.90062, 89.57699, 37.06992, 11.50365, 30.56621, 
    12.42591, 23.36816, 7.668781, 6.190823, 1.546305, 0.8410018, 0.8311342, 
    0.9131035, 1.001298, 1.305214, 1.981795, 2.674348, 3.756685, 6.685478, 
    12.5166, 33.46801, 39.22448, 3.996414, 5.474722, 10.38679, 23.22471, 
    119.96,
  95.25408, 96.67449, 89.9272, 35.5331, 101.1411, 20.56364, 80.37724, 
    41.99739, 104.1873, 26.53121, 8.58885, 5.016776, 3.217714, 2.705128, 
    2.387654, 2.276415, 2.447215, 2.601624, 4.990057, 9.271708, 15.32487, 
    44.10493, 8.845881, 6.234868, 3.088319, 3.878146, 6.087386, 18.48195, 
    101.6866,
  100.7407, 80.40129, 67.85948, 90.24564, 86.10168, 97.56203, 113.1837, 
    77.49389, 90.22321, 123.3514, 22.63876, 11.91433, 7.750029, 5.915522, 
    4.404317, 3.789989, 3.408443, 2.882893, 4.564136, 17.72578, 87.83972, 
    73.58538, 81.72456, 11.47144, 6.524117, 4.827785, 4.692759, 7.978117, 
    78.01582,
  50.1019, 30.04091, 56.23397, 80.35539, 154.1334, 111.3256, 104.1474, 
    129.7464, 119.4887, 96.36922, 93.13641, 32.15056, 16.11646, 10.06957, 
    7.618654, 5.95694, 4.775693, 4.245711, 4.568624, 83.03971, 93.72541, 
    103.7107, 100.3286, 49.36451, 19.28938, 10.92068, 7.964008, 7.522645, 
    32.26499,
  29.54198, 74.47705, 97.2665, 108.5334, 132.5167, 138.6021, 116.5708, 
    96.44563, 103.4887, 116.44, 127.8368, 119.4117, 27.31807, 17.60597, 
    12.86393, 9.687935, 8.373286, 8.104364, 9.997294, 73.75516, 98.22646, 
    104.9219, 104.2522, 100.5589, 58.1271, 19.68304, 10.82975, 8.295594, 
    11.10436,
  13.08329, 59.25195, 56.73753, 85.71684, 93.88824, 94.18108, 101.4064, 
    104.2222, 108.317, 111.2683, 105.3609, 99.46453, 70.88293, 54.80457, 
    22.87546, 19.42122, 54.09762, 40.86845, 79.33712, 98.31652, 88.51984, 
    84.29832, 34.73164, 71.0625, 23.51215, 11.34146, 9.804412, 8.55585, 
    9.009805,
  9.206236, 13.93191, 30.32398, 23.57718, 30.74948, 39.09873, 49.6731, 
    74.34364, 59.22871, 47.79567, 49.38109, 57.57881, 44.25893, 40.63794, 
    31.08079, 20.77725, 31.40985, 34.50206, 33.24142, 37.61687, 43.74236, 
    31.92351, 25.32459, 32.59917, 10.34481, 6.999294, 5.997006, 5.58165, 
    7.869718,
  7.993111, 8.980096, 10.46856, 11.75339, 12.90022, 12.74117, 13.82655, 
    14.27335, 14.80169, 15.78934, 15.91248, 14.96273, 13.54382, 12.59387, 
    11.75914, 10.69717, 9.998465, 9.740543, 10.10436, 9.704138, 9.056081, 
    8.507159, 7.643522, 7.018068, 6.474077, 6.321802, 6.456017, 6.582062, 
    7.474211 ;

 time = 547.5 ;

 time_bnds =
  365, 730 ;
}
