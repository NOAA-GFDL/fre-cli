netcdf atmos.1980-1981.alb_sfc.10 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:22 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.10.nc reduced/atmos.1980-1981.alb_sfc.10.nc\n",
			"Mon Aug 25 14:40:09 2025: cdo -O -s -select,month=10 merged_output.nc monthly_nc_files/all_years.10.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.33449, 76.33449, 76.33449, 76.33449, 76.33449, 76.33449, 76.33449, 
    76.28231, 76.28231, 76.28231, 76.28231, 76.28231, 76.28231, 76.28231, 
    76.23557, 76.23557, 76.23557, 76.23557, 76.23557, 76.23557, 76.23557, 
    76.33238, 76.33238, 76.33238, 76.33238, 76.33238, 76.33238, 76.33238, 
    76.33449,
  64.89365, 64.60094, 64.62613, 64.91412, 64.72925, 64.83128, 64.80768, 
    64.69353, 64.78751, 64.80426, 64.42357, 64.74329, 64.83408, 64.97444, 
    65.00816, 65.40665, 64.99274, 64.86215, 65.00487, 64.80632, 64.74576, 
    64.71924, 65.08601, 65.72659, 65.76024, 65.28751, 65.41483, 65.09593, 
    64.82298,
  56.30526, 56.79601, 59.39198, 55.29308, 50.35805, 50.47821, 55.3756, 
    50.49345, 50.31135, 50.45788, 50.42206, 50.35148, 50.74648, 59.09888, 
    59.41391, 58.53436, 57.30656, 57.74013, 58.19674, 58.36672, 56.97602, 
    55.6699, 53.22737, 50.1631, 54.28902, 53.15627, 51.95485, 52.43283, 
    56.38609,
  43.65289, 45.8708, 41.94007, 17.36793, 10.41739, 17.95782, 43.85882, 
    21.45577, 23.72284, 4.709009, 4.923261, 4.973978, 4.763111, 4.693274, 
    4.901066, 4.707689, 4.484168, 4.314278, 4.535184, 4.634959, 4.858424, 
    4.893921, 4.869491, 4.753322, 4.574074, 29.41581, 39.7373, 41.81701, 
    42.60708,
  3.83607, 3.967484, 3.964263, 3.959356, 4.050488, 4.101132, 4.074278, 
    4.089469, 4.051799, 3.98153, 4.05492, 4.034421, 4.19336, 4.205874, 
    4.258635, 4.075782, 3.873711, 3.961206, 3.902529, 4.009511, 4.115092, 
    4.161087, 4.113496, 8.478819, 4.612352, 3.98701, 3.788815, 4.017158, 
    3.849496,
  3.668314, 3.804784, 3.915586, 3.969654, 3.887734, 3.809336, 3.7607, 
    3.691919, 3.730085, 3.709102, 3.890545, 3.983998, 4.151096, 3.838039, 
    13.27409, 3.749172, 3.576822, 3.746467, 3.613502, 3.868504, 3.684616, 
    3.854016, 3.862535, 11.35291, 4.312171, 3.903355, 3.862175, 3.920177, 
    3.914024,
  3.47544, 3.858366, 12.43369, 3.658632, 3.688557, 3.55559, 3.797017, 
    3.578522, 3.713913, 3.964096, 9.962275, 14.95204, 10.72287, 3.851408, 
    3.690404, 3.742199, 3.607705, 3.799831, 3.457982, 3.740146, 3.619228, 
    3.724531, 3.654555, 4.565013, 9.238891, 3.506716, 3.654079, 3.611954, 
    3.652737,
  3.407367, 10.03827, 10.24111, 3.902563, 3.711976, 3.715958, 3.904224, 
    3.572152, 3.605497, 3.676147, 12.16595, 11.58705, 3.756984, 3.738649, 
    3.658054, 3.647351, 3.436167, 3.570407, 3.465508, 3.813663, 3.646457, 
    3.586645, 3.291835, 3.703038, 9.198439, 9.049075, 3.508026, 3.497301, 
    3.588902,
  3.163558, 6.088051, 8.764066, 9.460228, 3.502448, 3.290087, 3.489283, 
    3.394534, 3.44349, 3.409374, 4.764651, 3.174836, 4.462643, 3.363357, 
    3.213201, 3.584055, 3.380014, 3.609385, 3.605475, 3.797937, 3.518559, 
    3.591338, 3.214479, 8.374235, 8.817045, 11.90966, 3.605053, 3.408043, 
    3.330478,
  3.279573, 8.054596, 8.133905, 9.983292, 3.449507, 3.433797, 3.485979, 
    3.304253, 8.452133, 8.421389, 3.22094, 3.205667, 3.314472, 3.353131, 
    3.488217, 3.650631, 3.599582, 3.747967, 3.634994, 3.769408, 3.477436, 
    3.118848, 3.222192, 8.435213, 8.465815, 3.482133, 3.566371, 3.425734, 
    3.350325,
  9.401318, 9.979445, 10.28362, 9.05938, 14.6164, 3.570421, 4.948544, 
    3.394856, 3.387215, 3.203587, 3.958858, 3.1696, 3.031856, 3.169187, 
    3.210605, 3.05199, 3.232244, 3.31694, 3.273671, 3.362318, 3.322351, 
    3.059923, 8.463055, 7.408549, 3.207694, 3.225554, 3.074302, 3.015416, 
    8.680962,
  16.94011, 19.35202, 21.31767, 3.383593, 21.5316, 3.628977, 10.32176, 
    3.418007, 8.999545, 3.50762, 3.315124, 3.360814, 3.348656, 3.482226, 
    3.651538, 3.521955, 3.716624, 3.542851, 3.628517, 3.366624, 3.583625, 
    5.941592, 3.451103, 4.208598, 3.398862, 3.628376, 3.414477, 3.269738, 
    21.95075,
  21.61691, 18.01588, 18.78199, 17.54185, 11.91949, 13.73728, 11.61217, 
    9.728458, 9.443087, 10.04087, 3.447944, 3.513157, 3.5361, 3.680428, 
    3.641797, 3.537591, 3.824213, 3.695109, 3.713941, 3.739687, 11.31065, 
    11.0418, 8.703667, 3.653294, 3.399177, 3.873982, 3.703648, 4.007224, 
    9.826793,
  6.966265, 3.860702, 5.848576, 9.510167, 1.799804, 13.46157, 8.500051, 
    13.76139, 11.61508, 10.81792, 6.839441, 3.925494, 3.55592, 3.411594, 
    3.512713, 3.573277, 3.658669, 3.289186, 3.5492, 11.02724, 10.23037, 
    12.132, 11.3145, 4.594079, 3.662359, 3.720324, 3.612163, 3.779814, 
    4.954942,
  5.200716, 9.760414, 10.87848, 11.3665, 10.63656, 9.959309, 7.159617, 
    14.19822, 8.601541, 6.851152, 8.030232, 7.631159, 3.702308, 3.892982, 
    3.884258, 3.692162, 3.696695, 3.434785, 3.56104, 7.801659, 8.737359, 
    8.261608, 7.175056, 7.500792, 4.626308, 3.448804, 3.490095, 3.67881, 
    3.832444,
  3.922763, 5.706948, 5.960257, 5.514321, 6.124828, 6.036503, 6.562703, 
    8.206805, 8.497008, 8.27655, 7.809693, 13.12139, 12.2827, 7.809515, 
    3.219304, 3.710072, 7.820669, 10.20123, 9.61092, 6.546225, 5.769936, 
    9.318075, 4.042863, 11.25973, 3.312636, 6.400282, 3.924871, 3.991752, 
    3.844339,
  3.326933, 3.783619, 7.061045, 3.36075, 3.179795, 4.014248, 11.77929, 
    12.55296, 17.70358, 24.46612, 13.99687, 7.75606, 9.729899, 25.94917, 
    30.15984, 3.31827, 20.07007, 17.77384, 9.796602, 5.840931, 21.24125, 
    22.78789, 22.67719, 23.88843, 3.306564, 28.53911, 28.49304, 18.01253, 
    2.922757,
  9.077251, 1.853443, 9.195395, 7.875948, 4.875147, 11.53121, 13.55694, 
    13.23315, 13.56532, 13.35256, 12.93416, 12.55337, 12.94472, 13.14573, 
    12.9847, 12.66494, 12.49049, 12.53083, 12.62221, 12.65725, 12.49406, 
    11.74651, 11.16045, 11.7965, 11.19992, 11.23822, 11.10759, 11.12378, 
    13.17749 ;

 average_DT = 730 ;

 average_T1 = 289.5 ;

 average_T2 = 1019.5 ;

 climatology_bounds =
  289.5, 1019.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
