netcdf tracer_level.0003-0003.radon {
dimensions:
	bnds = 2 ;
	lat = 2 ;
	lon = 2 ;
	pfull = 65 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	float radon(time, pfull, lat, lon) ;
		radon:_FillValue = -1.e+10f ;
		radon:missing_value = -1.e+10f ;
		radon:units = "vmr*1e21" ;
		radon:long_name = "radon-222" ;
		radon:interp_method = "conserve_order1" ;
		radon:cell_methods = "time: mean" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.02" ;
		:git_hash = "b86d27037f755a82c586e55073dd575245c144b1" ;
		:creationtime = "Fri Dec  6 16:33:51 2024" ;
		:hostname = "pp211" ;
		:history = "Tue Sep 23 14:27:37 2025: ncks -d lon,0,1 tracer_level.0003-0003.radon.nc_lat01 tracer_level.0003-0003.radon.nc_lat01_lon01\n",
			"Tue Sep 23 14:26:18 2025: ncks -d lat,0,1 tracer_level.0003-0003.radon.nc tracer_level.0003-0003.radon.nc_lat01\n",
			"Tue Aug 12 16:38:49 2025: ncks -d lat,,,10 -d lon,,,10 tracer_level.0003-0003.radon.nc reduced/tracer_level.0003-0003.radon.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 00030101.atmos_tracer --interp_method conserve_order1 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field bk,pk,radon,ssalt1_emis,ssalt2_emis,ssalt3_emis,ssalt4_emis,ssalt5_emis,ssalt1_setl,ssalt2_setl,ssalt3_setl,ssalt4_setl,ssalt5_setl,ssalt1_wet_dep,ssalt2_wet_dep,ssalt3_wet_dep,ssalt4_wet_dep,ssalt5_wet_dep,ssalt1_dvel,ssalt2_dvel,ssalt3_dvel,ssalt4_dvel,ssalt5_dvel,ssalt1_ddep,ssalt2_ddep,ssalt3_ddep,ssalt4_ddep,ssalt5_ddep,scale_salt_emis,time_bnds --output_file out.nc" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.3.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -89.5, -79.5 ;

 lat_bnds =
  -90, -89,
  -80, -79 ;

 lon = 0.625, 13.125 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 radon =
  1.529905e-20, 1.529905e-20,
  2.792644e-20, 2.94163e-20,
  3.242325e-20, 3.242325e-20,
  7.029581e-20, 8.047592e-20,
  6.112494e-20, 6.112494e-20,
  1.626581e-19, 1.928468e-19,
  1.096101e-19, 1.096101e-19,
  2.749104e-19, 3.449383e-19,
  2.335068e-19, 2.335068e-19,
  4.396797e-19, 5.745231e-19,
  7.670262e-19, 7.670262e-19,
  8.44475e-19, 9.234996e-19,
  3.003618e-18, 3.003618e-18,
  2.536947e-18, 2.52326e-18,
  8.734008e-18, 8.734008e-18,
  1.119383e-17, 1.005254e-17,
  2.687149e-17, 2.687149e-17,
  5.017255e-17, 3.859873e-17,
  7.383607e-17, 7.383607e-17,
  2.501018e-16, 2.084324e-16,
  2.126669e-16, 2.126669e-16,
  7.605858e-16, 7.466835e-16,
  7.15242e-16, 7.15242e-16,
  2.029833e-15, 2.382652e-15,
  2.061948e-15, 2.061948e-15,
  4.043051e-15, 5.290443e-15,
  6.156443e-15, 6.156443e-15,
  6.723339e-15, 1.066336e-14,
  1.635776e-14, 1.635776e-14,
  1.210668e-14, 1.835511e-14,
  5.917032e-14, 5.917032e-14,
  3.814151e-14, 4.551538e-14,
  1.942057e-13, 1.942057e-13,
  1.758452e-13, 1.729065e-13,
  8.420157e-13, 8.420157e-13,
  6.553611e-13, 6.849211e-13,
  3.676693e-12, 3.676693e-12,
  3.377821e-12, 3.22574e-12,
  1.324723e-11, 1.324723e-11,
  1.279997e-11, 1.367475e-11,
  5.244899e-11, 5.244899e-11,
  4.140589e-11, 4.331211e-11,
  1.622715e-10, 1.622715e-10,
  1.585583e-10, 1.691203e-10,
  6.46474e-10, 6.46474e-10,
  6.118613e-10, 5.785175e-10,
  3.054962e-09, 3.054962e-09,
  3.581226e-09, 2.907362e-09,
  1.791809e-08, 1.791809e-08,
  2.71468e-08, 2.06764e-08,
  9.061949e-08, 9.061949e-08,
  1.183366e-07, 1.092687e-07,
  3.910738e-07, 3.910738e-07,
  4.410547e-07, 4.059652e-07,
  1.3234e-06, 1.3234e-06,
  1.73945e-06, 1.61254e-06,
  4.982602e-06, 4.982602e-06,
  7.986441e-06, 6.262919e-06,
  2.935227e-05, 2.935227e-05,
  3.047991e-05, 2.411587e-05,
  0.0001150029, 0.0001150029,
  0.0001219315, 8.384464e-05,
  0.001580484, 0.001580484,
  0.0005094475, 0.0003166444,
  0.006951712, 0.006951712,
  0.001530386, 0.001031392,
  0.01511111, 0.01511111,
  0.005332128, 0.003749793,
  0.02353415, 0.02353415,
  0.01732665, 0.01451974,
  0.04405832, 0.04405832,
  0.04354375, 0.04125238,
  0.08071082, 0.08071082,
  0.09177209, 0.08587226,
  0.1330787, 0.1330787,
  0.1716765, 0.1484769,
  0.1946154, 0.1946154,
  0.272545, 0.2262737,
  0.2565826, 0.2565826,
  0.3724229, 0.3113475,
  0.3135954, 0.3135954,
  0.4482261, 0.3872498,
  0.3573337, 0.3573337,
  0.4966939, 0.4465986,
  0.3869947, 0.3869947,
  0.5298803, 0.4908582,
  0.4063181, 0.4063181,
  0.5524696, 0.516091,
  0.4189714, 0.4189714,
  0.5645616, 0.5260128,
  0.425905, 0.425905,
  0.564113, 0.530057,
  0.4269015, 0.4269015,
  0.5555304, 0.5293595,
  0.422201, 0.422201,
  0.5396417, 0.5166984,
  0.4085007, 0.4085007,
  0.5178865, 0.4952067,
  0.386014, 0.386014,
  0.4916043, 0.4708295,
  0.3577868, 0.3577868,
  0.4621152, 0.4425593,
  0.3326207, 0.3326207,
  0.432183, 0.4118441,
  0.3141891, 0.3141891,
  0.4043238, 0.3821345,
  0.2990493, 0.2990493,
  0.3825701, 0.354023,
  0.2843398, 0.2843398,
  0.363676, 0.3297343,
  0.2687275, 0.2687275,
  0.3479453, 0.3093624,
  0.2555091, 0.2555091,
  0.3332098, 0.2909473,
  0.2406541, 0.2406541,
  0.3152442, 0.2749273,
  0.2266015, 0.2266015,
  0.2942939, 0.2590224,
  0.2121684, 0.2121684,
  0.275326, 0.2455239,
  0.195764, 0.195764,
  0.2611513, 0.2370166,
  0.1867052, 0.1867052,
  0.2500449, 0.2307612,
  0.1845552, 0.1845552,
  0.2397681, 0.2250075,
  0.1836565, 0.1836565,
  0.2343223, 0.2209795,
  0.1830172, 0.1830172,
  0.2321628, 0.2189483 ;

 time = 912.5 ;

 time_bnds =
  730, 1095 ;
}
