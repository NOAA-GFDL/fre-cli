netcdf \00010101.ocean_cobalt_btm {
dimensions:
	xh = 1440 ;
	yh = 1161 ;
	time = UNLIMITED ; // (1 currently)
	nv = 2 ;
variables:
	double xh(xh) ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
		xh:units = "degrees_east" ;
	double yh(yh) ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
		yh:units = "degrees_north" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
		time_bnds:units = "days since 0001-01-01 00:00:00" ;
	float fcadet_arag_btm(time, yh, xh) ;
		fcadet_arag_btm:long_name = "Aragonite sinking flux at bottom" ;
		fcadet_arag_btm:units = "mol m-2 s-1" ;
		fcadet_arag_btm:missing_value = 1.e+20f ;
		fcadet_arag_btm:_FillValue = 1.e+20f ;
		fcadet_arag_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fcadet_arag_btm:cell_measures = "area: areacello" ;
	float fcadet_calc_btm(time, yh, xh) ;
		fcadet_calc_btm:long_name = "Calcite sinking flux at bottom" ;
		fcadet_calc_btm:units = "mol m-2 s-1" ;
		fcadet_calc_btm:missing_value = 1.e+20f ;
		fcadet_calc_btm:_FillValue = 1.e+20f ;
		fcadet_calc_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fcadet_calc_btm:cell_measures = "area: areacello" ;
	float fcased_burial(time, yh, xh) ;
		fcased_burial:long_name = "Calcite permanent burial flux" ;
		fcased_burial:units = "mol m-2 s-1" ;
		fcased_burial:missing_value = 1.e+20f ;
		fcased_burial:_FillValue = 1.e+20f ;
		fcased_burial:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fcased_burial:cell_measures = "area: areacello" ;
	float fcased_redis(time, yh, xh) ;
		fcased_redis:long_name = "Calcite redissolution from sediments" ;
		fcased_redis:units = "mol m-2 s-1" ;
		fcased_redis:missing_value = 1.e+20f ;
		fcased_redis:_FillValue = 1.e+20f ;
		fcased_redis:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fcased_redis:cell_measures = "area: areacello" ;
	float fcased_redis_surfresp(time, yh, xh) ;
		fcased_redis_surfresp:long_name = "Calcite redissolution rom sediments, surfresp" ;
		fcased_redis_surfresp:units = "mol m-2 s-1" ;
		fcased_redis_surfresp:missing_value = 1.e+20f ;
		fcased_redis_surfresp:_FillValue = 1.e+20f ;
		fcased_redis_surfresp:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fcased_redis_surfresp:cell_measures = "area: areacello" ;
	float cased_redis_coef(time, yh, xh) ;
		cased_redis_coef:long_name = "Calcite redissolution from sediments, deepresp coefficient," ;
		cased_redis_coef:units = "s-1" ;
		cased_redis_coef:missing_value = 1.e+20f ;
		cased_redis_coef:_FillValue = 1.e+20f ;
		cased_redis_coef:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		cased_redis_coef:cell_measures = "area: areacello" ;
	float cased_redis_delz(time, yh, xh) ;
		cased_redis_delz:long_name = "Calcite redissolution from sediments, effective depth" ;
		cased_redis_delz:units = "none (0-1)" ;
		cased_redis_delz:missing_value = 1.e+20f ;
		cased_redis_delz:_FillValue = 1.e+20f ;
		cased_redis_delz:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		cased_redis_delz:cell_measures = "area: areacello" ;
	float ffetot_btm(time, yh, xh) ;
		ffetot_btm:long_name = "Total Fe sinking flux to bottom" ;
		ffetot_btm:units = "mol m-2 s-1" ;
		ffetot_btm:missing_value = 1.e+20f ;
		ffetot_btm:_FillValue = 1.e+20f ;
		ffetot_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		ffetot_btm:cell_measures = "area: areacello" ;
	float ffe_sed(time, yh, xh) ;
		ffe_sed:long_name = "Sediment iron efflux" ;
		ffe_sed:units = "mol m-2 s-1" ;
		ffe_sed:missing_value = 1.e+20f ;
		ffe_sed:_FillValue = 1.e+20f ;
		ffe_sed:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		ffe_sed:cell_measures = "area: areacello" ;
	float ffe_geotherm(time, yh, xh) ;
		ffe_geotherm:long_name = "Geothermal iron efflux" ;
		ffe_geotherm:units = "mol m-2 s-1" ;
		ffe_geotherm:missing_value = 1.e+20f ;
		ffe_geotherm:_FillValue = 1.e+20f ;
		ffe_geotherm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		ffe_geotherm:cell_measures = "area: areacello" ;
	float flithdet_btm(time, yh, xh) ;
		flithdet_btm:long_name = "Lithogenic detrital sinking flux burial" ;
		flithdet_btm:units = "g m-2 s-1" ;
		flithdet_btm:missing_value = 1.e+20f ;
		flithdet_btm:_FillValue = 1.e+20f ;
		flithdet_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		flithdet_btm:cell_measures = "area: areacello" ;
	float fntot_btm(time, yh, xh) ;
		fntot_btm:long_name = "Total N sinking flux to bottom" ;
		fntot_btm:units = "mol m-2 s-1" ;
		fntot_btm:missing_value = 1.e+20f ;
		fntot_btm:_FillValue = 1.e+20f ;
		fntot_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fntot_btm:cell_measures = "area: areacello" ;
	float fno3denit_sed(time, yh, xh) ;
		fno3denit_sed:long_name = "Sediment denitrification flux" ;
		fno3denit_sed:units = "mol m-2 s-1" ;
		fno3denit_sed:missing_value = 1.e+20f ;
		fno3denit_sed:_FillValue = 1.e+20f ;
		fno3denit_sed:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fno3denit_sed:cell_measures = "area: areacello" ;
	float fnoxic_sed(time, yh, xh) ;
		fnoxic_sed:long_name = "Sediment oxic Ndet remineralization flux" ;
		fnoxic_sed:units = "mol m-2 s-1" ;
		fnoxic_sed:missing_value = 1.e+20f ;
		fnoxic_sed:_FillValue = 1.e+20f ;
		fnoxic_sed:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fnoxic_sed:cell_measures = "area: areacello" ;
	float fptot_btm(time, yh, xh) ;
		fptot_btm:long_name = "Total P sinking flux to bottom" ;
		fptot_btm:units = "mol m-2 s-1" ;
		fptot_btm:missing_value = 1.e+20f ;
		fptot_btm:_FillValue = 1.e+20f ;
		fptot_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fptot_btm:cell_measures = "area: areacello" ;
	float fsitot_btm(time, yh, xh) ;
		fsitot_btm:long_name = "Total Si sinking flux to bottom" ;
		fsitot_btm:units = "mol m-2 s-1" ;
		fsitot_btm:missing_value = 1.e+20f ;
		fsitot_btm:_FillValue = 1.e+20f ;
		fsitot_btm:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fsitot_btm:cell_measures = "area: areacello" ;
	float fn_burial(time, yh, xh) ;
		fn_burial:long_name = "ndet burial flux" ;
		fn_burial:units = "mol m-2 s-1" ;
		fn_burial:missing_value = 1.e+20f ;
		fn_burial:_FillValue = 1.e+20f ;
		fn_burial:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fn_burial:cell_measures = "area: areacello" ;
	float fp_burial(time, yh, xh) ;
		fp_burial:long_name = "pdet burial flux" ;
		fp_burial:units = "mol m-2 s-1" ;
		fp_burial:missing_value = 1.e+20f ;
		fp_burial:_FillValue = 1.e+20f ;
		fp_burial:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		fp_burial:cell_measures = "area: areacello" ;
	float btm_temp(time, yh, xh) ;
		btm_temp:long_name = "Bottom Temperature" ;
		btm_temp:units = "deg C" ;
		btm_temp:missing_value = 1.e+20f ;
		btm_temp:_FillValue = 1.e+20f ;
		btm_temp:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_temp:cell_measures = "area: areacello" ;
	float btm_o2(time, yh, xh) ;
		btm_o2:long_name = "Bottom Oxygen" ;
		btm_o2:units = "mol kg-1" ;
		btm_o2:missing_value = 1.e+20f ;
		btm_o2:_FillValue = 1.e+20f ;
		btm_o2:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_o2:cell_measures = "area: areacello" ;
	float btm_htotal(time, yh, xh) ;
		btm_htotal:long_name = "Bottom Htotal" ;
		btm_htotal:units = "mol kg-1" ;
		btm_htotal:missing_value = 1.e+20f ;
		btm_htotal:_FillValue = 1.e+20f ;
		btm_htotal:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_htotal:cell_measures = "area: areacello" ;
	float btm_co3_ion(time, yh, xh) ;
		btm_co3_ion:long_name = "Bottom Carbonate Ion" ;
		btm_co3_ion:units = "mol kg-1" ;
		btm_co3_ion:missing_value = 1.e+20f ;
		btm_co3_ion:_FillValue = 1.e+20f ;
		btm_co3_ion:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_co3_ion:cell_measures = "area: areacello" ;
	float btm_co3_sol_arag(time, yh, xh) ;
		btm_co3_sol_arag:long_name = "Bottom Aragonite Solubility" ;
		btm_co3_sol_arag:units = "mol kg-1" ;
		btm_co3_sol_arag:missing_value = 1.e+20f ;
		btm_co3_sol_arag:_FillValue = 1.e+20f ;
		btm_co3_sol_arag:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_co3_sol_arag:cell_measures = "area: areacello" ;
	float btm_co3_sol_calc(time, yh, xh) ;
		btm_co3_sol_calc:long_name = "Bottom Calcite Solubility" ;
		btm_co3_sol_calc:units = "mol kg-1" ;
		btm_co3_sol_calc:missing_value = 1.e+20f ;
		btm_co3_sol_calc:_FillValue = 1.e+20f ;
		btm_co3_sol_calc:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		btm_co3_sol_calc:cell_measures = "area: areacello" ;
	float cased(time, yh, xh) ;
		cased:long_name = "calcium carbonate in sediment" ;
		cased:units = "mol m-3" ;
		cased:missing_value = 1.e+20f ;
		cased:_FillValue = 1.e+20f ;
		cased:cell_methods = "xh:mean yh:mean area:mean time: mean" ;
		cased:cell_measures = "area: areacello" ;

// global attributes:
		:associated_files = "areacello: 00010101.ocean_static.nc" ;
data:

 xh = -299.875, -299.625, -299.375, -299.125, -298.875, -298.625, -298.375, 
    -298.125, -297.875, -297.625, -297.375, -297.125, -296.875, -296.625, 
    -296.375, -296.125, -295.875, -295.625, -295.375, -295.125, -294.875, 
    -294.625, -294.375, -294.125, -293.875, -293.625, -293.375, -293.125, 
    -292.875, -292.625, -292.375, -292.125, -291.875, -291.625, -291.375, 
    -291.125, -290.875, -290.625, -290.375, -290.125, -289.875, -289.625, 
    -289.375, -289.125, -288.875, -288.625, -288.375, -288.125, -287.875, 
    -287.625, -287.375, -287.125, -286.875, -286.625, -286.375, -286.125, 
    -285.875, -285.625, -285.375, -285.125, -284.875, -284.625, -284.375, 
    -284.125, -283.875, -283.625, -283.375, -283.125, -282.875, -282.625, 
    -282.375, -282.125, -281.875, -281.625, -281.375, -281.125, -280.875, 
    -280.625, -280.375, -280.125, -279.875, -279.625, -279.375, -279.125, 
    -278.875, -278.625, -278.375, -278.125, -277.875, -277.625, -277.375, 
    -277.125, -276.875, -276.625, -276.375, -276.125, -275.875, -275.625, 
    -275.375, -275.125, -274.875, -274.625, -274.375, -274.125, -273.875, 
    -273.625, -273.375, -273.125, -272.875, -272.625, -272.375, -272.125, 
    -271.875, -271.625, -271.375, -271.125, -270.875, -270.625, -270.375, 
    -270.125, -269.875, -269.625, -269.375, -269.125, -268.875, -268.625, 
    -268.375, -268.125, -267.875, -267.625, -267.375, -267.125, -266.875, 
    -266.625, -266.375, -266.125, -265.875, -265.625, -265.375, -265.125, 
    -264.875, -264.625, -264.375, -264.125, -263.875, -263.625, -263.375, 
    -263.125, -262.875, -262.625, -262.375, -262.125, -261.875, -261.625, 
    -261.375, -261.125, -260.875, -260.625, -260.375, -260.125, -259.875, 
    -259.625, -259.375, -259.125, -258.875, -258.625, -258.375, -258.125, 
    -257.875, -257.625, -257.375, -257.125, -256.875, -256.625, -256.375, 
    -256.125, -255.875, -255.625, -255.375, -255.125, -254.875, -254.625, 
    -254.375, -254.125, -253.875, -253.625, -253.375, -253.125, -252.875, 
    -252.625, -252.375, -252.125, -251.875, -251.625, -251.375, -251.125, 
    -250.875, -250.625, -250.375, -250.125, -249.875, -249.625, -249.375, 
    -249.125, -248.875, -248.625, -248.375, -248.125, -247.875, -247.625, 
    -247.375, -247.125, -246.875, -246.625, -246.375, -246.125, -245.875, 
    -245.625, -245.375, -245.125, -244.875, -244.625, -244.375, -244.125, 
    -243.875, -243.625, -243.375, -243.125, -242.875, -242.625, -242.375, 
    -242.125, -241.875, -241.625, -241.375, -241.125, -240.875, -240.625, 
    -240.375, -240.125, -239.875, -239.625, -239.375, -239.125, -238.875, 
    -238.625, -238.375, -238.125, -237.875, -237.625, -237.375, -237.125, 
    -236.875, -236.625, -236.375, -236.125, -235.875, -235.625, -235.375, 
    -235.125, -234.875, -234.625, -234.375, -234.125, -233.875, -233.625, 
    -233.375, -233.125, -232.875, -232.625, -232.375, -232.125, -231.875, 
    -231.625, -231.375, -231.125, -230.875, -230.625, -230.375, -230.125, 
    -229.875, -229.625, -229.375, -229.125, -228.875, -228.625, -228.375, 
    -228.125, -227.875, -227.625, -227.375, -227.125, -226.875, -226.625, 
    -226.375, -226.125, -225.875, -225.625, -225.375, -225.125, -224.875, 
    -224.625, -224.375, -224.125, -223.875, -223.625, -223.375, -223.125, 
    -222.875, -222.625, -222.375, -222.125, -221.875, -221.625, -221.375, 
    -221.125, -220.875, -220.625, -220.375, -220.125, -219.875, -219.625, 
    -219.375, -219.125, -218.875, -218.625, -218.375, -218.125, -217.875, 
    -217.625, -217.375, -217.125, -216.875, -216.625, -216.375, -216.125, 
    -215.875, -215.625, -215.375, -215.125, -214.875, -214.625, -214.375, 
    -214.125, -213.875, -213.625, -213.375, -213.125, -212.875, -212.625, 
    -212.375, -212.125, -211.875, -211.625, -211.375, -211.125, -210.875, 
    -210.625, -210.375, -210.125, -209.875, -209.625, -209.375, -209.125, 
    -208.875, -208.625, -208.375, -208.125, -207.875, -207.625, -207.375, 
    -207.125, -206.875, -206.625, -206.375, -206.125, -205.875, -205.625, 
    -205.375, -205.125, -204.875, -204.625, -204.375, -204.125, -203.875, 
    -203.625, -203.375, -203.125, -202.875, -202.625, -202.375, -202.125, 
    -201.875, -201.625, -201.375, -201.125, -200.875, -200.625, -200.375, 
    -200.125, -199.875, -199.625, -199.375, -199.125, -198.875, -198.625, 
    -198.375, -198.125, -197.875, -197.625, -197.375, -197.125, -196.875, 
    -196.625, -196.375, -196.125, -195.875, -195.625, -195.375, -195.125, 
    -194.875, -194.625, -194.375, -194.125, -193.875, -193.625, -193.375, 
    -193.125, -192.875, -192.625, -192.375, -192.125, -191.875, -191.625, 
    -191.375, -191.125, -190.875, -190.625, -190.375, -190.125, -189.875, 
    -189.625, -189.375, -189.125, -188.875, -188.625, -188.375, -188.125, 
    -187.875, -187.625, -187.375, -187.125, -186.875, -186.625, -186.375, 
    -186.125, -185.875, -185.625, -185.375, -185.125, -184.875, -184.625, 
    -184.375, -184.125, -183.875, -183.625, -183.375, -183.125, -182.875, 
    -182.625, -182.375, -182.125, -181.875, -181.625, -181.375, -181.125, 
    -180.875, -180.625, -180.375, -180.125, -179.875, -179.625, -179.375, 
    -179.125, -178.875, -178.625, -178.375, -178.125, -177.875, -177.625, 
    -177.375, -177.125, -176.875, -176.625, -176.375, -176.125, -175.875, 
    -175.625, -175.375, -175.125, -174.875, -174.625, -174.375, -174.125, 
    -173.875, -173.625, -173.375, -173.125, -172.875, -172.625, -172.375, 
    -172.125, -171.875, -171.625, -171.375, -171.125, -170.875, -170.625, 
    -170.375, -170.125, -169.875, -169.625, -169.375, -169.125, -168.875, 
    -168.625, -168.375, -168.125, -167.875, -167.625, -167.375, -167.125, 
    -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375, -163.125, -162.875, -162.625, -162.375, -162.125, -161.875, 
    -161.625, -161.375, -161.125, -160.875, -160.625, -160.375, -160.125, 
    -159.875, -159.625, -159.375, -159.125, -158.875, -158.625, -158.375, 
    -158.125, -157.875, -157.625, -157.375, -157.125, -156.875, -156.625, 
    -156.375, -156.125, -155.875, -155.625, -155.375, -155.125, -154.875, 
    -154.625, -154.375, -154.125, -153.875, -153.625, -153.375, -153.125, 
    -152.875, -152.625, -152.375, -152.125, -151.875, -151.625, -151.375, 
    -151.125, -150.875, -150.625, -150.375, -150.125, -149.875, -149.625, 
    -149.375, -149.125, -148.875, -148.625, -148.375, -148.125, -147.875, 
    -147.625, -147.375, -147.125, -146.875, -146.625, -146.375, -146.125, 
    -145.875, -145.625, -145.375, -145.125, -144.875, -144.625, -144.375, 
    -144.125, -143.875, -143.625, -143.375, -143.125, -142.875, -142.625, 
    -142.375, -142.125, -141.875, -141.625, -141.375, -141.125, -140.875, 
    -140.625, -140.375, -140.125, -139.875, -139.625, -139.375, -139.125, 
    -138.875, -138.625, -138.375, -138.125, -137.875, -137.625, -137.375, 
    -137.125, -136.875, -136.625, -136.375, -136.125, -135.875, -135.625, 
    -135.375, -135.125, -134.875, -134.625, -134.375, -134.125, -133.875, 
    -133.625, -133.375, -133.125, -132.875, -132.625, -132.375, -132.125, 
    -131.875, -131.625, -131.375, -131.125, -130.875, -130.625, -130.375, 
    -130.125, -129.875, -129.625, -129.375, -129.125, -128.875, -128.625, 
    -128.375, -128.125, -127.875, -127.625, -127.375, -127.125, -126.875, 
    -126.625, -126.375, -126.125, -125.875, -125.625, -125.375, -125.125, 
    -124.875, -124.625, -124.375, -124.125, -123.875, -123.625, -123.375, 
    -123.125, -122.875, -122.625, -122.375, -122.125, -121.875, -121.625, 
    -121.375, -121.125, -120.875, -120.625, -120.375, -120.125, -119.875, 
    -119.625, -119.375, -119.125, -118.875, -118.625, -118.375, -118.125, 
    -117.875, -117.625, -117.375, -117.125, -116.875, -116.625, -116.375, 
    -116.125, -115.875, -115.625, -115.375, -115.125, -114.875, -114.625, 
    -114.375, -114.125, -113.875, -113.625, -113.375, -113.125, -112.875, 
    -112.625, -112.375, -112.125, -111.875, -111.625, -111.375, -111.125, 
    -110.875, -110.625, -110.375, -110.125, -109.875, -109.625, -109.375, 
    -109.125, -108.875, -108.625, -108.375, -108.125, -107.875, -107.625, 
    -107.375, -107.125, -106.875, -106.625, -106.375, -106.125, -105.875, 
    -105.625, -105.375, -105.125, -104.875, -104.625, -104.375, -104.125, 
    -103.875, -103.625, -103.375, -103.125, -102.875, -102.625, -102.375, 
    -102.125, -101.875, -101.625, -101.375, -101.125, -100.875, -100.625, 
    -100.375, -100.125, -99.875, -99.625, -99.375, -99.125, -98.875, -98.625, 
    -98.375, -98.125, -97.875, -97.625, -97.375, -97.125, -96.875, -96.625, 
    -96.375, -96.125, -95.875, -95.625, -95.375, -95.125, -94.875, -94.625, 
    -94.375, -94.125, -93.875, -93.625, -93.375, -93.125, -92.875, -92.625, 
    -92.375, -92.125, -91.875, -91.625, -91.375, -91.125, -90.875, -90.625, 
    -90.375, -90.125, -89.875, -89.625, -89.375, -89.125, -88.875, -88.625, 
    -88.375, -88.125, -87.875, -87.625, -87.375, -87.125, -86.875, -86.625, 
    -86.375, -86.125, -85.875, -85.625, -85.375, -85.125, -84.875, -84.625, 
    -84.375, -84.125, -83.875, -83.625, -83.375, -83.125, -82.875, -82.625, 
    -82.375, -82.125, -81.875, -81.625, -81.375, -81.125, -80.875, -80.625, 
    -80.375, -80.125, -79.875, -79.625, -79.375, -79.125, -78.875, -78.625, 
    -78.375, -78.125, -77.875, -77.625, -77.375, -77.125, -76.875, -76.625, 
    -76.375, -76.125, -75.875, -75.625, -75.375, -75.125, -74.875, -74.625, 
    -74.375, -74.125, -73.875, -73.625, -73.375, -73.125, -72.875, -72.625, 
    -72.375, -72.125, -71.875, -71.625, -71.375, -71.125, -70.875, -70.625, 
    -70.375, -70.125, -69.875, -69.625, -69.375, -69.125, -68.875, -68.625, 
    -68.375, -68.125, -67.875, -67.625, -67.375, -67.125, -66.875, -66.625, 
    -66.375, -66.125, -65.875, -65.625, -65.375, -65.125, -64.875, -64.625, 
    -64.375, -64.125, -63.875, -63.625, -63.375, -63.125, -62.875, -62.625, 
    -62.375, -62.125, -61.875, -61.625, -61.375, -61.125, -60.875, -60.625, 
    -60.375, -60.125, -59.875, -59.625, -59.375, -59.125, -58.875, -58.625, 
    -58.375, -58.125, -57.875, -57.625, -57.375, -57.125, -56.875, -56.625, 
    -56.375, -56.125, -55.875, -55.625, -55.375, -55.125, -54.875, -54.625, 
    -54.375, -54.125, -53.875, -53.625, -53.375, -53.125, -52.875, -52.625, 
    -52.375, -52.125, -51.875, -51.625, -51.375, -51.125, -50.875, -50.625, 
    -50.375, -50.125, -49.875, -49.625, -49.375, -49.125, -48.875, -48.625, 
    -48.375, -48.125, -47.875, -47.625, -47.375, -47.125, -46.875, -46.625, 
    -46.375, -46.125, -45.875, -45.625, -45.375, -45.125, -44.875, -44.625, 
    -44.375, -44.125, -43.875, -43.625, -43.375, -43.125, -42.875, -42.625, 
    -42.375, -42.125, -41.875, -41.625, -41.375, -41.125, -40.875, -40.625, 
    -40.375, -40.125, -39.875, -39.625, -39.375, -39.125, -38.875, -38.625, 
    -38.375, -38.125, -37.875, -37.625, -37.375, -37.125, -36.875, -36.625, 
    -36.375, -36.125, -35.875, -35.625, -35.375, -35.125, -34.875, -34.625, 
    -34.375, -34.125, -33.875, -33.625, -33.375, -33.125, -32.875, -32.625, 
    -32.375, -32.125, -31.875, -31.625, -31.375, -31.125, -30.875, -30.625, 
    -30.375, -30.125, -29.875, -29.625, -29.375, -29.125, -28.875, -28.625, 
    -28.375, -28.125, -27.875, -27.625, -27.375, -27.125, -26.875, -26.625, 
    -26.375, -26.125, -25.875, -25.625, -25.375, -25.125, -24.875, -24.625, 
    -24.375, -24.125, -23.875, -23.625, -23.375, -23.125, -22.875, -22.625, 
    -22.375, -22.125, -21.875, -21.625, -21.375, -21.125, -20.875, -20.625, 
    -20.375, -20.125, -19.875, -19.625, -19.375, -19.125, -18.875, -18.625, 
    -18.375, -18.125, -17.875, -17.625, -17.375, -17.125, -16.875, -16.625, 
    -16.375, -16.125, -15.875, -15.625, -15.375, -15.125, -14.875, -14.625, 
    -14.375, -14.125, -13.875, -13.625, -13.375, -13.125, -12.875, -12.625, 
    -12.375, -12.125, -11.875, -11.625, -11.375, -11.125, -10.875, -10.625, 
    -10.375, -10.125, -9.875, -9.625, -9.375, -9.125, -8.875, -8.625, -8.375, 
    -8.125, -7.875, -7.625, -7.375, -7.125, -6.875, -6.625, -6.375, -6.125, 
    -5.875, -5.625, -5.375, -5.125, -4.875, -4.625, -4.375, -4.125, -3.875, 
    -3.625, -3.375, -3.125, -2.875, -2.625, -2.375, -2.125, -1.875, -1.625, 
    -1.375, -1.125, -0.875, -0.625, -0.375, -0.125, 0.125, 0.375, 0.625, 
    0.875, 1.125, 1.375, 1.625, 1.875, 2.125, 2.375, 2.625, 2.875, 3.125, 
    3.375, 3.625, 3.875, 4.125, 4.375, 4.625, 4.875, 5.125, 5.375, 5.625, 
    5.875, 6.125, 6.375, 6.625, 6.875, 7.125, 7.375, 7.625, 7.875, 8.125, 
    8.375, 8.625, 8.875, 9.125, 9.375, 9.625, 9.875, 10.125, 10.375, 10.625, 
    10.875, 11.125, 11.375, 11.625, 11.875, 12.125, 12.375, 12.625, 12.875, 
    13.125, 13.375, 13.625, 13.875, 14.125, 14.375, 14.625, 14.875, 15.125, 
    15.375, 15.625, 15.875, 16.125, 16.375, 16.625, 16.875, 17.125, 17.375, 
    17.625, 17.875, 18.125, 18.375, 18.625, 18.875, 19.125, 19.375, 19.625, 
    19.875, 20.125, 20.375, 20.625, 20.875, 21.125, 21.375, 21.625, 21.875, 
    22.125, 22.375, 22.625, 22.875, 23.125, 23.375, 23.625, 23.875, 24.125, 
    24.375, 24.625, 24.875, 25.125, 25.375, 25.625, 25.875, 26.125, 26.375, 
    26.625, 26.875, 27.125, 27.375, 27.625, 27.875, 28.125, 28.375, 28.625, 
    28.875, 29.125, 29.375, 29.625, 29.875, 30.125, 30.375, 30.625, 30.875, 
    31.125, 31.375, 31.625, 31.875, 32.125, 32.375, 32.625, 32.875, 33.125, 
    33.375, 33.625, 33.875, 34.125, 34.375, 34.625, 34.875, 35.125, 35.375, 
    35.625, 35.875, 36.125, 36.375, 36.625, 36.875, 37.125, 37.375, 37.625, 
    37.875, 38.125, 38.375, 38.625, 38.875, 39.125, 39.375, 39.625, 39.875, 
    40.125, 40.375, 40.625, 40.875, 41.125, 41.375, 41.625, 41.875, 42.125, 
    42.375, 42.625, 42.875, 43.125, 43.375, 43.625, 43.875, 44.125, 44.375, 
    44.625, 44.875, 45.125, 45.375, 45.625, 45.875, 46.125, 46.375, 46.625, 
    46.875, 47.125, 47.375, 47.625, 47.875, 48.125, 48.375, 48.625, 48.875, 
    49.125, 49.375, 49.625, 49.875, 50.125, 50.375, 50.625, 50.875, 51.125, 
    51.375, 51.625, 51.875, 52.125, 52.375, 52.625, 52.875, 53.125, 53.375, 
    53.625, 53.875, 54.125, 54.375, 54.625, 54.875, 55.125, 55.375, 55.625, 
    55.875, 56.125, 56.375, 56.625, 56.875, 57.125, 57.375, 57.625, 57.875, 
    58.125, 58.375, 58.625, 58.875, 59.125, 59.375, 59.625, 59.875 ;

 yh = -88.5208813286133, -88.4226439858398, -88.3244066430664, 
    -88.2261693002929, -88.1279319575195, -88.029694614746, 
    -87.9314572719726, -87.8332199291991, -87.7349825864257, 
    -87.6367452436523, -87.5385079008788, -87.4402705581054, 
    -87.3420332153319, -87.2437958725585, -87.145558529785, 
    -87.0473211870116, -86.9490838442381, -86.8508465014647, 
    -86.7526091586912, -86.6543718159178, -86.5561344731444, 
    -86.4578971303709, -86.3596597875975, -86.261422444824, 
    -86.1631851020506, -86.0649477592771, -85.9667104165037, 
    -85.8684730737302, -85.7702357309568, -85.6719983881833, 
    -85.5737610454099, -85.4755237026365, -85.377286359863, 
    -85.2790490170895, -85.1808116743161, -85.0825743315427, 
    -84.9843369887692, -84.8860996459958, -84.7878623032223, 
    -84.6896249604489, -84.5913876176754, -84.493150274902, 
    -84.3949129321285, -84.2966755893551, -84.1984382465816, 
    -84.1002009038082, -84.0019635610348, -83.9037262182613, 
    -83.8054888754879, -83.7072515327144, -83.609014189941, 
    -83.5107768471675, -83.4125395043941, -83.3143021616206, 
    -83.2160648188472, -83.1178274760737, -83.0195901333003, 
    -82.9213527905269, -82.8231154477534, -82.72487810498, -82.6266407622065, 
    -82.5284034194331, -82.4301660766596, -82.3319287338862, 
    -82.2336913911127, -82.1354540483393, -82.0372167055658, 
    -81.9389793627924, -81.840742020019, -81.7425046772455, -81.644267334472, 
    -81.5460299916986, -81.4477926489252, -81.3495553061517, 
    -81.2513179633783, -81.1530806206048, -81.0548432778314, 
    -80.9566059350579, -80.8583685922845, -80.760131249511, 
    -80.6618939067376, -80.5636565639641, -80.4654192211907, 
    -80.3671818784173, -80.2689445356438, -80.1707071928704, 
    -80.0724698500969, -79.9742325073235, -79.87599516455, -79.7777578217766, 
    -79.6795204790031, -79.5812831362297, -79.4830457934562, 
    -79.3848084506828, -79.2865711079094, -79.1883337651359, 
    -79.0900964223624, -78.991859079589, -78.8936217368156, 
    -78.7953843940421, -78.6971470512687, -78.5989097084952, 
    -78.5006723657218, -78.4024350229483, -78.3041976801749, 
    -78.2059603374015, -78.107722994628, -78.0094856518545, 
    -77.9112483090811, -77.8130109663077, -77.7147736235342, 
    -77.6165362807608, -77.5182989379873, -77.4200615952139, 
    -77.3218242524404, -77.223586909667, -77.1253495668935, 
    -77.0271122241201, -76.9288748813466, -76.8306375385732, 
    -76.7324001957998, -76.6341628530263, -76.5359255102529, 
    -76.4376881674794, -76.339450824706, -76.2412134819325, 
    -76.1429761391591, -76.0447387963856, -75.9465014536122, 
    -75.8482641108387, -75.7500267680653, -75.6517894252919, 
    -75.5535520825184, -75.4553147397449, -75.3570773969715, 
    -75.2588400541981, -75.1606027114246, -75.0623653686512, 
    -74.9641280258777, -74.8658906831043, -74.7676533403308, 
    -74.6694159975574, -74.5711786547839, -74.4729413120105, 
    -74.374703969237, -74.2764666264636, -74.1782292836902, 
    -74.0799919409167, -73.9817545981433, -73.8835172553698, 
    -73.7852799125964, -73.6870425698229, -73.5888052270495, 
    -73.490567884276, -73.3923305415026, -73.2940931987291, 
    -73.1958558559557, -73.0976185131823, -72.9993811704088, 
    -72.9011438276354, -72.8029064848619, -72.7046691420885, 
    -72.606431799315, -72.5081944565416, -72.4099571137681, 
    -72.3117197709947, -72.2134824282212, -72.1152450854478, 
    -72.0170077426744, -71.9187703999009, -71.8205330571274, 
    -71.722295714354, -71.6240583715806, -71.5258210288071, 
    -71.4275836860337, -71.3293463432602, -71.2311090004868, 
    -71.1328716577133, -71.0346343149399, -70.9363969721664, 
    -70.838159629393, -70.7399222866195, -70.6416849438461, 
    -70.5434476010727, -70.4452102582992, -70.3469729155258, 
    -70.2487355727523, -70.1504982299789, -70.0522608872054, 
    -69.954023544432, -69.8557862016585, -69.7575488588851, 
    -69.6593115161116, -69.5610741733382, -69.4628368305648, 
    -69.3645994877913, -69.2663621450179, -69.1681248022444, 
    -69.069887459471, -68.9716501166975, -68.8734127739241, 
    -68.7751754311506, -68.6769380883772, -68.5787007456037, 
    -68.4804634028303, -68.3822260600569, -68.2839887172834, 
    -68.1857513745099, -68.0875140317365, -67.9892766889631, 
    -67.8910393461896, -67.7928020034162, -67.6945646606427, 
    -67.5963273178693, -67.4980899750958, -67.3998526323224, 
    -67.3016152895489, -67.2033779467755, -67.105140604002, 
    -67.0069032612286, -66.9086659184552, -66.8103746406885, 
    -66.7117331375991, -66.6126955029787, -66.5132604431118, 
    -66.4134266638701, -66.3131928707682, -66.2125577690213, 
    -66.1115200636031, -66.0100784593041, -65.9082316607918, 
    -65.8059783726705, -65.7033172995429, -65.6002471460721, 
    -65.4967666170443, -65.3928744174327, -65.2885692524622, 
    -65.1838498276744, -65.0787148489947, -64.9731630227985, 
    -64.8671930559803, -64.760803656022, -64.6539935310628, 
    -64.5467613899703, -64.4391059424119, -64.3310258989275, 
    -64.2225199710027, -64.1135868711439, -64.0042253129527, 
    -63.894434011203, -63.784211681918, -63.6735570424482, -63.5624688115505, 
    -63.4509457094688, -63.3389864580144, -63.2265897806486, 
    -63.1137544025655, -63.0004790507758, -62.8867624541921, 
    -62.7726033437149, -62.6580004523194, -62.5429525151436, 
    -62.4274582695774, -62.3115164553525, -62.1951258146335, 
    -62.0782850921101, -61.9609930350901, -61.8432483935938, 
    -61.7250499204486, -61.6063963713863, -61.4872865051392, 
    -61.3677190835396, -61.2476928716185, -61.1272066377062, 
    -61.0062591535343, -60.884849194338, -60.7629755389598, 
    -60.6406369699546, -60.5178322736953, -60.3945602404801, 
    -60.2708196646404, -60.14660934465, -60.0219280832357, -59.8967746874882, 
    -59.7711479689751, -59.6450467438542, -59.5184698329885, 
    -59.3914160620619, -59.2638842616962, -59.1358732675693, 
    -59.0073819205344, -58.8784090667402, -58.7489535577527, 
    -58.6190142506776, -58.4885900082839, -58.3576796991292, 
    -58.2262821976854, -58.0943963844658, -57.9620211461538, 
    -57.8291553757318, -57.6957979726119, -57.5619478427679, 
    -57.4276038988677, -57.2927650604075, -57.1574302538468, 
    -57.0215984127446, -56.8852684778969, -56.7484393974749, 
    -56.6111101271648, -56.4732796303085, -56.3349468780456, 
    -56.1961108494559, -56.0567705317041, -55.9169249201846, 
    -55.7765730186677, -55.6357138394476, -55.4943464034902, 
    -55.3524697405834, -55.2100828894873, -55.0671848980862, 
    -54.9237748235415, -54.7798517324457, -54.6354147009772, 
    -54.4904628150566, -54.3449951705041, -54.199010873197, 
    -54.0525090392296, -53.9054887950733, -53.7579492777379, 
    -53.6098896349336, -53.4613090252352, -53.3122066182453, 
    -53.1625815947607, -53.0124331469381, -52.8617604784615, 
    -52.7105628047106, -52.5588393529298, -52.4065893623985, 
    -52.2538120846021, -52.1005067834039, -51.9466727352183, 
    -51.7923092291839, -51.637415567339, -51.4819910647963, 
    -51.3260350499197, -51.1695468645014, -51.0125258639398, 
    -50.8549714174182, -50.6968829080846, -50.5382597332318, 
    -50.3791013044785, -50.2194070479511, -50.0591764044664, 
    -49.8984088297146, -49.7371037944429, -49.5752607846407, 
    -49.412879301724, -49.2499588627218, -49.0864990004619, 
    -48.9224992637582, -48.7579592175979, -48.5928784433296, 
    -48.4272565388516, -48.2610931188013, -48.0943878147438, 
    -47.9271402753627, -47.7593501666492, -47.5910171720937, 
    -47.4221409928761, -47.2527213480571, -47.08275797477, -46.9122506284122, 
    -46.7411990828373, -46.5696031305474, -46.3974625828856, 
    -46.2247772702279, -46.0515470421768, -45.8777717677532, 
    -45.7034513355895, -45.5285856541224, -45.3531746517856, 
    -45.1772182772023, -45.0007164993782, -44.8236693078935, 
    -44.6460767130959, -44.4679387462917, -44.2892554599388, 
    -44.1100269278373, -43.9302532453218, -43.7499345294513, 
    -43.5690709192008, -43.3876625756504, -43.205709682176, 
    -43.0232124446377, -42.8401710915687, -42.6565858743633, 
    -42.4724570674644, -42.2877849685499, -42.1025698987191, 
    -41.9168122026777, -41.730512248922, -41.5436704299229, 
    -41.3562871623085, -41.1683628870455, -40.9798980696201, 
    -40.790893200218, -40.6013487939026, -40.4112653907925, 
    -40.2206435562383, -40.0294838809969, -39.8377869814059, 
    -39.6455534995561, -39.4527841034619, -39.2594794872318, 
    -39.0656403712361, -38.8712675022735, -38.6763616537367, 
    -38.4809236257751, -38.2849542454572, -38.0884543669302, 
    -37.8914248715784, -37.6938666681796, -37.4957806930597, 
    -37.2971679102448, -37.0980293116122, -36.8983659170386, 
    -36.6981787745468, -36.4974689604493, -36.2962375794908, 
    -36.0944857649878, -35.8922146789658, -35.6894255122942, 
    -35.4861194848192, -35.2822978454935, -35.0779618725039, 
    -34.8731128733961, -34.667752185197, -34.461881174534, -34.255501237752, 
    -34.0486138010269, -33.8412203204768, -33.6333222822699, 
    -33.4249212027298, -33.2160186284369, -33.0066161363278, 
    -32.7967153337909, -32.5863178587586, -32.3754253797966, 
    -32.1640395961899, -31.952162238025, -31.739795066269, -31.5269398728455, 
    -31.3135984807058, -31.0997727438981, -30.8854645476315, 
    -30.6706758083373, -30.4554084737265, -30.2396645228428, 
    -30.0234459661121, -29.8067548453888, -29.5895932339964, 
    -29.3719632367664, -29.1538669900706, -28.9353066618517, 
    -28.7162844516478, -28.496802590614, -28.2768633415386, 
    -28.0564689988566, -27.8356218886569, -27.6143243686867, 
    -27.3925788283504, -27.1703876887049, -26.9477534024496, 
    -26.7246784539123, -26.5011653590304, -26.2772166653272, 
    -26.0528349518839, -25.8280228293068, -25.6027829396893, 
    -25.3771179565698, -25.1510305848841, -24.9245235609136, 
    -24.6975996522279, -24.470261657623, -24.2425124070545, 
    -24.0143547615654, -23.7857916132091, -23.5568258849681, 
    -23.3274605306659, -23.0976985348757, -22.8675429128228, 
    -22.6369967102824, -22.4060630034717, -22.1747448989375, 
    -21.9430455334382, -21.7109680738206, -21.4785157168916, 
    -21.2456916892848, -21.0124992473213, -20.7789416768659, 
    -20.5450222931779, -20.3107444407557, -20.0761114931781, 
    -19.841126852938, -19.6057939512726, -19.3701162479875, 
    -19.1340972312755, -18.8977404175304, -18.6610493511555, 
    -18.4240276043667, -18.1866787769903, -17.9490064962555, 
    -17.7110144165822, -17.4727062193628, -17.2340856127391, 
    -16.9951563313743, -16.7559221362196, -16.5163868142751, 
    -16.2765541783467, -16.0364280667968, -15.7960123432904, 
    -15.5553108965366, -15.3143276400236, -15.0730665117507, 
    -14.8315314739535, -14.5897265128255, -14.3476556382336, 
    -14.1053228834302, -13.862732304759, -13.6198879813569, 
    -13.3767940148509, -13.1334545290505, -12.889873669635, 
    -12.6460556038367, -12.4020045201193, -12.1577246278516, 
    -11.9132201569774, -11.6684953576804, -11.4235545000447, 
    -11.1784018737118, -10.9330417875323, -10.6874785692145, 
    -10.4417165649682, -10.1957601391447, -9.9496136738729, 
    -9.70328156869134, -9.45676824017667, -9.21007812156814, 
    -8.96321566238849, -8.71618532806131, -8.46899159952477, 
    -8.22163897284192, -7.97413195880769, -7.72647508255252, 
    -7.4786728831428, -7.2307299131782, -6.98265073838595, -6.73443993721214, 
    -6.48610210041021, -6.23764183062656, -5.98906374198353, 
    -5.74037245965978, -5.49157261946812, -5.24266886743094, 
    -4.9936658593533, -4.74456826039377, -4.49538074463318, 
    -4.24610799464126, -3.9967547010414, -3.74732556207348, 
    -3.49782528315504, -3.2482585764407, -2.99863016038011, 
    -2.74894475927441, -2.49920710283131, -2.24942192571902, 
    -1.99959396711887, -1.74972797027709, -1.49982868205542, 
    -1.24990085248112, -0.999949234296017, -0.749978582505122, 
    -0.499993653924574, -0.249999206729245, 0, 0.249999206729245, 
    0.499993653924574, 0.749978582505122, 0.999949234296017, 
    1.24990085248112, 1.49982868205542, 1.74972797027709, 1.99959396711887, 
    2.24942192571902, 2.49920710283131, 2.74894475927441, 2.99863016038011, 
    3.2482585764407, 3.49782528315504, 3.74732556207348, 3.9967547010414, 
    4.24610799464126, 4.49538074463318, 4.74456826039377, 4.9936658593533, 
    5.24266886743094, 5.49157261946812, 5.74037245965978, 5.98906374198353, 
    6.23764183062656, 6.48610210041021, 6.73443993721214, 6.98265073838595, 
    7.2307299131782, 7.4786728831428, 7.72647508255252, 7.97413195880769, 
    8.22163897284192, 8.46899159952477, 8.71618532806131, 8.96321566238849, 
    9.21007812156814, 9.45676824017667, 9.70328156869134, 9.9496136738729, 
    10.1957601391447, 10.4417165649682, 10.6874785692145, 10.9330417875323, 
    11.1784018737118, 11.4235545000447, 11.6684953576804, 11.9132201569774, 
    12.1577246278516, 12.4020045201193, 12.6460556038367, 12.889873669635, 
    13.1334545290505, 13.3767940148509, 13.6198879813569, 13.862732304759, 
    14.1053228834302, 14.3476556382336, 14.5897265128255, 14.8315314739535, 
    15.0730665117507, 15.3143276400236, 15.5553108965366, 15.7960123432904, 
    16.0364280667968, 16.2765541783467, 16.5163868142751, 16.7559221362196, 
    16.9951563313743, 17.2340856127391, 17.4727062193628, 17.7110144165822, 
    17.9490064962555, 18.1866787769903, 18.4240276043667, 18.6610493511555, 
    18.8977404175304, 19.1340972312755, 19.3701162479875, 19.6057939512726, 
    19.841126852938, 20.0761114931781, 20.3107444407557, 20.5450222931779, 
    20.7789416768659, 21.0124992473213, 21.2456916892848, 21.4785157168916, 
    21.7109680738206, 21.9430455334382, 22.1747448989375, 22.4060630034717, 
    22.6369967102824, 22.8675429128228, 23.0976985348757, 23.3274605306659, 
    23.5568258849681, 23.7857916132091, 24.0143547615654, 24.2425124070545, 
    24.470261657623, 24.6975996522279, 24.9245235609136, 25.1510305848841, 
    25.3771179565698, 25.6027829396893, 25.8280228293068, 26.0528349518839, 
    26.2772166653272, 26.5011653590304, 26.7246784539123, 26.9477534024496, 
    27.1703876887049, 27.3925788283504, 27.6143243686867, 27.8356218886569, 
    28.0564689988566, 28.2768633415386, 28.496802590614, 28.7162844516478, 
    28.9353066618517, 29.1538669900706, 29.3719632367664, 29.5895932339964, 
    29.8067548453888, 30.0234459661121, 30.2396645228428, 30.4554084737265, 
    30.6706758083373, 30.8854645476315, 31.0997727438981, 31.3135984807058, 
    31.5269398728455, 31.739795066269, 31.952162238025, 32.1640395961899, 
    32.3754253797966, 32.5863178587586, 32.7967153337909, 33.0066161363278, 
    33.2160186284369, 33.4249212027298, 33.6333222822699, 33.8412203204768, 
    34.0486138010269, 34.255501237752, 34.461881174534, 34.667752185197, 
    34.8731128733961, 35.0779618725039, 35.2822978454935, 35.4861194848192, 
    35.6894255122942, 35.8922146789658, 36.0944857649878, 36.2962375794908, 
    36.4974689604493, 36.6981787745468, 36.8983659170386, 37.0980293116122, 
    37.2971679102448, 37.4957806930597, 37.6938666681796, 37.8914248715784, 
    38.0884543669302, 38.2849542454572, 38.4809236257751, 38.6763616537367, 
    38.8712675022735, 39.0656403712361, 39.2594794872318, 39.4527841034619, 
    39.6455534995561, 39.8377869814059, 40.0294838809969, 40.2206435562383, 
    40.4112653907925, 40.6013487939026, 40.790893200218, 40.9798980696201, 
    41.1683628870455, 41.3562871623085, 41.5436704299229, 41.730512248922, 
    41.9168122026777, 42.1025698987191, 42.2877849685499, 42.4724570674644, 
    42.6565858743633, 42.8401710915687, 43.0232124446377, 43.205709682176, 
    43.3876625756504, 43.5690709192008, 43.7499345294513, 43.9302532453218, 
    44.1100269278373, 44.2892554599388, 44.4679387462917, 44.6460767130959, 
    44.8236693078935, 45.0007164993782, 45.1772182772023, 45.3531746517856, 
    45.5285856541224, 45.7034513355895, 45.8777717677532, 46.0515470421768, 
    46.2247772702279, 46.3974625828856, 46.5696031305474, 46.7411990828373, 
    46.9122506284122, 47.08275797477, 47.2527213480571, 47.4221409928761, 
    47.5910171720937, 47.7593501666492, 47.9271402753627, 48.0943878147438, 
    48.2610931188013, 48.4272565388516, 48.5928784433296, 48.7579592175979, 
    48.9224992637582, 49.0864990004619, 49.2499588627218, 49.412879301724, 
    49.5752607846407, 49.7371037944429, 49.8984088297146, 50.0591764044664, 
    50.2194070479511, 50.3791013044785, 50.5382597332318, 50.6968829080846, 
    50.8549714174182, 51.0125258639398, 51.1695468645014, 51.3260350499197, 
    51.4819910647963, 51.637415567339, 51.7923092291839, 51.9466727352183, 
    52.1005067834039, 52.2538120846021, 52.4065893623985, 52.5588393529298, 
    52.7105628047106, 52.8617604784615, 53.0124331469381, 53.1625815947607, 
    53.3122066182453, 53.4613090252352, 53.6098896349336, 53.7579492777379, 
    53.9054887950733, 54.0525090392296, 54.199010873197, 54.3449951705041, 
    54.4904628150566, 54.6354147009772, 54.7798517324457, 54.9237748235415, 
    55.0671848980862, 55.2100828894873, 55.3524697405834, 55.4943464034902, 
    55.6357138394476, 55.7765730186677, 55.9169249201846, 56.0567705317041, 
    56.1961108494559, 56.3349468780456, 56.4732796303085, 56.6111101271648, 
    56.7484393974749, 56.8852684778969, 57.0215984127446, 57.1574302538468, 
    57.2927650604075, 57.4276038988677, 57.5619478427679, 57.6957979726119, 
    57.8291553757318, 57.9620211461538, 58.0943963844658, 58.2262821976854, 
    58.3576796991292, 58.4885900082839, 58.6190142506776, 58.7489535577527, 
    58.8784090667402, 59.0073819205344, 59.1358732675693, 59.2638842616962, 
    59.3914160620619, 59.5184698329885, 59.6450467438542, 59.7711479689751, 
    59.8967746874882, 60.0219280832357, 60.14660934465, 60.2708196646404, 
    60.3945602404801, 60.5178322736953, 60.6406369699546, 60.7629755389598, 
    60.884849194338, 61.0062591535343, 61.1272066377062, 61.2476928716185, 
    61.3677190835396, 61.4872865051392, 61.6063963713863, 61.7250499204486, 
    61.8432483935938, 61.9609930350901, 62.0782850921101, 62.1951258146335, 
    62.3115164553525, 62.4274582695774, 62.5429525151436, 62.6580004523194, 
    62.7726033437149, 62.8867624541921, 63.0004790507758, 63.1137544025655, 
    63.2265897806486, 63.3389864580144, 63.4509457094688, 63.5624688115505, 
    63.6735570424482, 63.784211681918, 63.894434011203, 64.0042253129527, 
    64.1130035635913, 64.2210912313842, 64.3291788991772, 64.4372665669701, 
    64.545354234763, 64.653441902556, 64.7615295703489, 64.8696172381418, 
    64.9777049059348, 65.0857925737277, 65.1938802415207, 65.3019679093136, 
    65.4100555771065, 65.5181432448995, 65.6262309126924, 65.7343185804854, 
    65.8424062482783, 65.9504939160712, 66.0585815838642, 66.1666692516571, 
    66.2747569194501, 66.382844587243, 66.4909322550359, 66.5990199228289, 
    66.7071075906218, 66.8151952584147, 66.9232829262077, 67.0313705940006, 
    67.1394582617935, 67.2475459295865, 67.3556335973794, 67.4637212651724, 
    67.5718089329653, 67.6798966007582, 67.7879842685512, 67.8960719363441, 
    68.0041596041371, 68.11224727193, 68.2203349397229, 68.3284226075159, 
    68.4365102753088, 68.5445979431017, 68.6526856108947, 68.7607732786876, 
    68.8688609464806, 68.9769486142735, 69.0850362820664, 69.1931239498594, 
    69.3012116176523, 69.4092992854453, 69.5173869532382, 69.6254746210311, 
    69.7335622888241, 69.841649956617, 69.9497376244099, 70.0578252922029, 
    70.1659129599958, 70.2740006277888, 70.3820882955817, 70.4901759633746, 
    70.5982636311676, 70.7063512989605, 70.8144389667535, 70.9225266345464, 
    71.0306143023393, 71.1387019701323, 71.2467896379252, 71.3548773057181, 
    71.4629649735111, 71.571052641304, 71.679140309097, 71.7872279768899, 
    71.8953156446828, 72.0034033124758, 72.1114909802687, 72.2195786480616, 
    72.3276663158546, 72.4357539836475, 72.5438416514405, 72.6519293192334, 
    72.7600169870263, 72.8681046548193, 72.9761923226122, 73.0842799904052, 
    73.1923676581981, 73.300455325991, 73.408542993784, 73.5166306615769, 
    73.6247183293698, 73.7328059971628, 73.8408936649557, 73.9489813327487, 
    74.0570690005416, 74.1651566683345, 74.2732443361275, 74.3813320039204, 
    74.4894196717133, 74.5975073395063, 74.7055950072992, 74.8136826750922, 
    74.9217703428851, 75.029858010678, 75.137945678471, 75.2460333462639, 
    75.3541210140569, 75.4622086818498, 75.5702963496427, 75.6783840174357, 
    75.7864716852286, 75.8945593530215, 76.0026470208145, 76.1107346886074, 
    76.2188223564004, 76.3269100241933, 76.4349976919862, 76.5430853597792, 
    76.6511730275721, 76.7592606953651, 76.867348363158, 76.9754360309509, 
    77.0835236987439, 77.1916113665368, 77.2996990343298, 77.4077867021227, 
    77.5158743699156, 77.6239620377086, 77.7320497055015, 77.8401373732944, 
    77.9482250410874, 78.0563127088803, 78.1644003766733, 78.2724880444662, 
    78.3805757122591, 78.4886633800521, 78.596751047845, 78.7048387156379, 
    78.8129263834309, 78.9210140512238, 79.0291017190168, 79.1371893868097, 
    79.2452770546026, 79.3533647223956, 79.4614523901885, 79.5695400579815, 
    79.6776277257744, 79.7857153935673, 79.8938030613603, 80.0018907291532, 
    80.1099783969461, 80.2180660647391, 80.326153732532, 80.434241400325, 
    80.5423290681179, 80.6504167359108, 80.7585044037038, 80.8665920714967, 
    80.9746797392897, 81.0827674070826, 81.1908550748755, 81.2989427426685, 
    81.4070304104614, 81.5151180782543, 81.6232057460473, 81.7312934138402, 
    81.8393810816331, 81.9474687494261, 82.055556417219, 82.163644085012, 
    82.2717317528049, 82.3798194205978, 82.4879070883908, 82.5959947561837, 
    82.7040824239767, 82.8121700917696, 82.9202577595625, 83.0283454273555, 
    83.1364330951484, 83.2445207629414, 83.3526084307343, 83.4606960985272, 
    83.5687837663202, 83.6768714341131, 83.7849591019061, 83.893046769699, 
    84.0011344374919, 84.1092221052849, 84.2173097730778, 84.3253974408707, 
    84.4334851086637, 84.5415727764566, 84.6496604442495, 84.7577481120425, 
    84.8658357798354, 84.9739234476284, 85.0820111154213, 85.1900987832142, 
    85.2981864510072, 85.4062741188001, 85.5143617865931, 85.622449454386, 
    85.7305371221789, 85.8386247899719, 85.9467124577648, 86.0548001255577, 
    86.1628877933507, 86.2709754611436, 86.3790631289366, 86.4871507967295, 
    86.5952384645225, 86.7033261323154, 86.8114138001083, 86.9195014679013, 
    87.0275891356942, 87.1356768034871, 87.2437644712801, 87.351852139073, 
    87.4599398068659, 87.5680274746589, 87.6761151424518, 87.7842028102448, 
    87.8922904780377, 88.0003781458306, 88.1084658136236, 88.2165534814165, 
    88.3246411492095, 88.4327288170024, 88.5408164847953, 88.6489041525883, 
    88.7569918203812, 88.8650794881741, 88.9731671559671, 89.08125482376, 
    89.189342491553, 89.2974301593459, 89.4055178271388, 89.5136054949318, 
    89.6216931627247, 89.7297808305177, 89.8378684983106, 89.9459561661037 ;

 time = 15.5 ;

 nv = 1, 2 ;
}
