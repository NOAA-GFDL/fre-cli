netcdf \00010101.atmos_daily.tile3.ps {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  101029.5, 100948.3, 101092.3, 101193.2, 101319.1, 101478.1, 101571.2, 
    101658.9, 101803.2, 101718.2, 101906.6, 102368.2, 102403.8, 102097.4, 
    102104.7,
  101050.6, 100974.8, 101005.8, 101039.6, 101224.7, 101266.9, 101544, 101637, 
    101711.9, 101941, 102128.6, 102298.6, 102470.6, 100668.1, 101518.5,
  101144.6, 101084.1, 101087.9, 101113.8, 101200.6, 97804.13, 101447, 
    101733.2, 101750.6, 101895.3, 102059.5, 102186, 102370, 102558, 102746.2,
  101119.9, 101170.1, 101196.4, 101235.1, 101367.2, 101346.1, 97669.09, 
    101535.7, 101818.3, 101942.3, 102061.7, 102136.3, 102298.3, 102513.6, 
    102752,
  101040.1, 101213.3, 101286.8, 101356, 101451.6, 101592.3, 101607, 95427.53, 
    94772.33, 101866.3, 102112.1, 102154.3, 102279, 102411.6, 102697.5,
  101068.9, 101231.6, 101349.8, 101432.3, 101497, 101609.6, 101769.8, 
    101826.5, 101807.8, 102130, 102174.2, 102194.7, 102303.8, 102432.7, 
    102643.9,
  101223.7, 101368, 101468, 101569.1, 101634, 101724, 101804.4, 101969.2, 
    102088.8, 102146, 102213.2, 102282.1, 102358.3, 102474.1, 102640.2,
  101497.7, 101573.7, 101626.4, 101702.4, 101753.8, 101851.1, 101945.8, 
    102033.4, 102116.4, 102222.7, 102307, 102381.8, 102442.9, 102540.2, 
    102662.9,
  101740, 101796.8, 101838, 101902.6, 101967.5, 102036.3, 102110, 102210.9, 
    102286.9, 102354.2, 102437.2, 102513.5, 102573.9, 102677.8, 102795.5,
  101975.2, 101993.4, 102023.2, 102064.9, 102105.7, 102191, 102283.9, 
    102374.7, 102478.8, 102547.5, 102613, 102688.4, 102752.8, 102828, 102883.5,
  100537.1, 100555.7, 100697.4, 100621.5, 100624.3, 100432.4, 100179.9, 
    99936.51, 99790.98, 99442.31, 99576.24, 100075.7, 100235.7, 100245, 100561,
  100556.9, 100481.4, 100575, 100650.8, 100717.6, 100402.3, 100424.5, 
    100181.8, 100008.1, 100028.6, 100096.5, 100349.3, 100620.7, 99122.48, 
    100219.4,
  100729.8, 100622.4, 100612.5, 100694.4, 100663.8, 97136.84, 100475.3, 
    100533.9, 100406.2, 100349.5, 100399.5, 100596.7, 100920, 101220.6, 
    101620.7,
  100933, 100864.2, 100828.8, 100820.8, 100882.9, 100657.2, 96918.36, 
    100489.6, 100613.5, 100660.1, 100711.7, 100864, 101167.1, 101551.7, 
    101913.1,
  101101.2, 101059.3, 101028.5, 101011.7, 101010.2, 101022.5, 100886.7, 
    94677.49, 94048.63, 100785.7, 101021.3, 101142, 101401.2, 101685, 102113.5,
  101268.6, 101230.3, 101188, 101166.6, 101144.2, 101126.6, 101165.3, 
    101126.3, 100961, 101222.7, 101295.4, 101394.4, 101627.9, 101917.3, 
    102265.1,
  101405.5, 101396.1, 101351.8, 101337.1, 101319.7, 101322.4, 101293.5, 
    101360.6, 101428, 101442.8, 101532.7, 101653, 101827.2, 102080.8, 102387,
  101556.9, 101546.7, 101510.2, 101481.9, 101435, 101430.6, 101441.1, 
    101442.1, 101480.2, 101614.6, 101760.2, 101887.9, 102053.3, 102277.8, 
    102548.1,
  101701, 101701.6, 101682.9, 101667, 101647.6, 101616.2, 101594.5, 101642, 
    101707.9, 101796.9, 101929, 102079.3, 102219.7, 102421.1, 102660.7,
  101854.8, 101852.3, 101835.5, 101827.6, 101801.2, 101816.8, 101834.2, 
    101847.5, 101895.2, 101966.2, 102094.7, 102246.5, 102373.6, 102559, 
    102759.1,
  100628.5, 100465, 100375.5, 100278.3, 100217.6, 100145.7, 99986.81, 
    99856.74, 99804.44, 99611.55, 99902.02, 100501.8, 100628, 100499.4, 100576,
  100602.7, 100477, 100332.9, 100206.7, 100089.1, 99797.42, 99879.91, 
    99692.3, 99602.45, 99854.79, 100132.6, 100506.1, 100765.2, 99172.52, 
    100109.8,
  100638.4, 100494.2, 100337.7, 100175.5, 99856.27, 96335.68, 99626.51, 
    99742.22, 99678.09, 99891.75, 100145.1, 100491.9, 100850.9, 101127.5, 
    101418.9,
  100655.5, 100517.4, 100378.3, 100181.2, 100001.6, 99580.81, 95923.34, 
    99457.01, 99644.83, 99909.08, 100206, 100513.3, 100885.5, 101284.1, 
    101606.8,
  100701.6, 100571.9, 100444.7, 100267.9, 100070.8, 99847.27, 99600.41, 
    93606.07, 93093.51, 99810.66, 100284, 100578.6, 100963, 101303, 101737.3,
  100760.6, 100650.2, 100517.5, 100370.6, 100166.3, 99931.4, 99810.04, 
    99767.23, 99613.07, 100089.5, 100346.4, 100684.2, 101063.7, 101464.8, 
    101845.8,
  100850.6, 100759.6, 100636.1, 100502.6, 100327.4, 100126.4, 99918.5, 
    99955.42, 100072.9, 100192.6, 100460, 100815.6, 101180.1, 101571.6, 
    101944.3,
  100968.6, 100889.3, 100774.1, 100651.3, 100471.4, 100305.8, 100171.6, 
    100087.8, 100127.5, 100339.5, 100649.4, 100972.9, 101346.9, 101725.2, 
    102156.4,
  101100.2, 101045.3, 100954.6, 100845.1, 100703.5, 100544.4, 100418.8, 
    100410, 100485.5, 100633.2, 100904.5, 101207, 101551.2, 101948.5, 102379.7,
  101264.4, 101203.2, 101131.4, 101042.2, 100914.1, 100794.7, 100707.1, 
    100664.7, 100724.4, 100887, 101179, 101486.3, 101821.5, 102229.4, 102579.2,
  101102.3, 100968.4, 100913, 100815, 100785.3, 100814.2, 100967.7, 101229.6, 
    101476.6, 101386.6, 101627.2, 102207.3, 102351.5, 102147.4, 102113.1,
  100910.8, 100802.4, 100756, 100703.5, 100704.4, 100579.9, 100866.7, 
    101068.5, 101291.5, 101625.7, 101893.1, 102274.1, 102538.9, 100813, 
    101658.5,
  100787, 100727.6, 100704.3, 100663.3, 100516.3, 97133.28, 100668.9, 
    101050.4, 101332, 101640, 101936.6, 102306.9, 102654.6, 102850.2, 102981.4,
  100669.7, 100652.6, 100626.8, 100580.1, 100550.3, 100390.8, 96920.89, 
    100806, 101277.3, 101659.6, 102034.8, 102355.8, 102694.4, 102960.3, 
    103119.3,
  100611.1, 100611.5, 100572.9, 100528.8, 100481.3, 100522.8, 100618.9, 
    94897.48, 94547.84, 101582.3, 102155, 102440.7, 102756.5, 102922.1, 
    103177.4,
  100574.1, 100568.5, 100503.4, 100446.4, 100408.8, 100417.5, 100779.9, 
    100991.9, 101146.6, 101849.8, 102203.5, 102523.9, 102807.2, 103018.6, 
    103236.3,
  100559.4, 100549.6, 100468.4, 100399.6, 100385.6, 100443.9, 100724.8, 
    101199.9, 101630.1, 101906.1, 102281.5, 102612, 102851.5, 103098.6, 
    103326.2,
  100573, 100538.9, 100438.2, 100348.1, 100344.9, 100471, 100829.9, 101155.5, 
    101523.5, 101965.5, 102376.8, 102682.8, 102968.5, 103244.1, 103512.3,
  100610.4, 100580, 100463, 100377.5, 100407.2, 100586.5, 100939, 101352.6, 
    101741, 102088.1, 102482.9, 102799.9, 103103, 103405.7, 103705.2,
  100674.2, 100626.7, 100494.2, 100429, 100493.2, 100744, 101088.1, 101407.8, 
    101771.6, 102188.7, 102612, 102947.4, 103286.2, 103622.9, 103899,
  102304.9, 102268.4, 102314, 102330.4, 102373.2, 102475.9, 102726.4, 
    103068.2, 103348.8, 103229.7, 103472.1, 103973.6, 103948.8, 103549.4, 
    103339.3,
  102071.6, 102032.6, 102041.2, 102077.5, 102267.2, 102358.4, 102831.1, 
    103084, 103286.2, 103577.3, 103800.7, 104047.4, 104143.2, 102191.2, 
    102902.4,
  101852.6, 101842.2, 101877.4, 101965.3, 102144.1, 98947.41, 102729.1, 
    103200.1, 103457.2, 103647.6, 103859.8, 104087.3, 104260.3, 104255.6, 
    104245.6,
  101656.5, 101671.6, 101738.4, 101854.5, 102196.9, 102246, 98853.62, 
    102898.7, 103361.6, 103647.4, 103947.5, 104125, 104297.1, 104371.8, 104388,
  101446.6, 101531.7, 101640, 101809.3, 102107, 102420.9, 102558.8, 96755.73, 
    96354.45, 103500.6, 104022.2, 104191.4, 104365.7, 104364.6, 104441.1,
  101278.2, 101410.6, 101554.7, 101739.3, 102016.6, 102282.7, 102718, 
    102918.7, 103036.4, 103748.3, 104028.8, 104251.8, 104404.5, 104464.8, 
    104495.8,
  101142.8, 101343.4, 101515.1, 101717.1, 101968.1, 102214.1, 102591.7, 
    103063.1, 103476, 103744.5, 104052.8, 104322.7, 104441.9, 104514.4, 
    104544.5,
  101048.9, 101292.6, 101482.4, 101685.1, 101890.3, 102139.5, 102586.6, 
    102921.6, 103309.6, 103719.4, 104118.3, 104363.6, 104500.6, 104582.9, 
    104645.3,
  101007.4, 101292.8, 101501.1, 101697.9, 101894.6, 102149.6, 102597.4, 
    103041.7, 103446.3, 103786.7, 104166.5, 104406.5, 104540.3, 104638, 104718,
  101006.8, 101298.2, 101498.9, 101691.1, 101902.4, 102218.5, 102679.4, 
    103024.9, 103414.4, 103817.7, 104213.5, 104444.3, 104598.3, 104727.2, 
    104799.7,
  103276.3, 103369, 103545, 103679.1, 103891.3, 104065.9, 104233.9, 104514, 
    104740.8, 104510.3, 104592.5, 104828.6, 104518.1, 103920.3, 103673.9,
  103084.7, 103187.5, 103361.6, 103523.7, 103777.9, 103837.1, 104251.1, 
    104476.5, 104638.3, 104845.5, 104913.3, 104904.4, 104722.9, 102611.2, 
    103268.3,
  102903.5, 103038.8, 103210.2, 103381.4, 103576, 100309.8, 104124.5, 
    104618.2, 104807.5, 104890, 104940.7, 104941.1, 104829, 104687.6, 104601.5,
  102748.3, 102875, 103054, 103209.6, 103547.1, 103620.9, 100162.9, 104226.6, 
    104636.8, 104853.9, 104982.8, 104956, 104871.7, 104763.5, 104736.5,
  102588, 102726.5, 102902.9, 103066.8, 103368.5, 103763.7, 103860.1, 
    97953.4, 97457.62, 104576.4, 105008.7, 104977.8, 104927.6, 104786.5, 
    104773.9,
  102411.9, 102553.8, 102730, 102900.6, 103183.8, 103542.9, 103941.9, 
    104139.7, 104156, 104807.3, 104950.3, 104996.6, 104942.6, 104884.5, 
    104835.4,
  102217.9, 102396.6, 102576.3, 102754.7, 103051.9, 103412, 103748.1, 
    104208.9, 104544.9, 104726.5, 104905.6, 105020.1, 104970.4, 104944.3, 
    104884.8,
  102010.2, 102216.4, 102400.3, 102611, 102914.3, 103261.6, 103636.4, 
    103940.5, 104270.2, 104634.7, 104900.7, 105006.6, 105007.5, 104996.6, 
    104955.5,
  101835.4, 102077.4, 102283.1, 102509.2, 102849.9, 103172.8, 103551.9, 
    103965.8, 104346.6, 104572, 104872.8, 105006.9, 105046.8, 105038.1, 
    104994.9,
  101681.7, 101926.9, 102170.8, 102422.2, 102771.7, 103099.2, 103489.6, 
    103815.1, 104164.2, 104483.3, 104843.2, 105000.2, 105068.7, 105069.6, 
    105015,
  103759.6, 103860.2, 104067.4, 104235.8, 104476.9, 104644.1, 104719.7, 
    104802.3, 104780.9, 104312.4, 104219.7, 104357, 104166, 103709, 103522.2,
  103626.9, 103729.1, 103935.5, 104150.2, 104422.8, 104437.4, 104734.8, 
    104795, 104748.2, 104717, 104576.7, 104473.6, 104377.3, 102413.7, 103143.1,
  103475.2, 103622.1, 103828.9, 104069.9, 104278.4, 100837.1, 104597, 
    104919.1, 104938.3, 104814.3, 104691, 104563.6, 104500.7, 104500.9, 
    104487.7,
  103316.2, 103484.1, 103699.5, 103941.2, 104302.1, 104248.4, 100639.9, 
    104555.7, 104812, 104856.4, 104798.6, 104646.9, 104577.7, 104580.8, 
    104627.2,
  103127.3, 103333, 103560.1, 103842.5, 104157.1, 104466.8, 104448.3, 
    98348.58, 97636.8, 104644.7, 104878, 104740, 104670.5, 104590.9, 104628.3,
  102924.6, 103142.6, 103382.4, 103693.2, 104018.8, 104280.7, 104583.6, 
    104603.8, 104506, 104879.4, 104896.6, 104833.9, 104746, 104697, 104661.1,
  102697.6, 102954.3, 103228.7, 103549.3, 103914.9, 104202.2, 104405.9, 
    104652.8, 104795.9, 104845.3, 104928.8, 104918.8, 104833.5, 104780.8, 
    104743.7,
  102462, 102735.1, 103037.6, 103389.8, 103741.7, 104064.9, 104303.5, 
    104447.5, 104612.9, 104831.8, 104971.2, 104974.2, 104922.4, 104852.9, 
    104817.4,
  102248.6, 102568.7, 102894.8, 103257.4, 103643.3, 103960.2, 104182.5, 
    104390.8, 104638.2, 104770.3, 104979.8, 105030.4, 105004.7, 104932, 
    104872.7,
  102060.8, 102375.1, 102726.6, 103108.9, 103483.5, 103827.2, 104065.3, 
    104207.8, 104451.2, 104672.2, 104951.6, 105041.3, 105063.1, 105006, 
    104938.3,
  103193.1, 103300.4, 103550.5, 103705.6, 103901.7, 103975.6, 103946.9, 
    103961, 103999.4, 103724.5, 103878.3, 104252.3, 104148.4, 103721.8, 
    103567.5,
  102986.9, 103108.9, 103390, 103605.1, 103862.6, 103802.8, 103997.9, 
    103973.4, 103960.8, 104064.6, 104151.6, 104289.9, 104329, 102403.7, 103171,
  102762.4, 102945.7, 103254.2, 103522.3, 103713.8, 100226.2, 103879.4, 
    104063.2, 104079.1, 104082.1, 104167.3, 104273.7, 104411, 104473.8, 
    104514.3,
  102569.1, 102779.1, 103114.1, 103396.1, 103748.6, 103644, 99957.77, 
    103786.7, 104005.3, 104102.4, 104179.2, 104267.7, 104397.2, 104532.8, 
    104627,
  102432.6, 102674.9, 103014, 103320.3, 103628.8, 103859.5, 103795, 97625.81, 
    96979.18, 103907.8, 104203.5, 104269.5, 104411.3, 104486, 104621.3,
  102351.6, 102595.2, 102916.1, 103236.6, 103529.9, 103696.1, 103946.2, 
    103926.8, 103814.8, 104112.1, 104203.5, 104270.9, 104392.8, 104482, 
    104574.9,
  102330.5, 102564.9, 102870.3, 103155.8, 103458.8, 103668.4, 103818.7, 
    103962.5, 104046.7, 104106.1, 104211, 104302, 104394.7, 104477, 104548.2,
  102292.8, 102505.9, 102769.5, 103060.3, 103336, 103563.9, 103783.5, 
    103872.4, 103965.9, 104119.4, 104249.2, 104325.7, 104413, 104513.6, 
    104603.1,
  102212.2, 102430.5, 102692.5, 102957.4, 103253.3, 103492.3, 103712.8, 
    103894.4, 104010, 104162.9, 104295.7, 104381.1, 104459.2, 104556.4, 
    104637.2,
  102069.9, 102268.6, 102526.6, 102821.1, 103118.2, 103379.9, 103635, 
    103816.2, 103954, 104139.8, 104314.3, 104429.4, 104511.1, 104609.2, 
    104670.3,
  102369.4, 102545.6, 102884.8, 103142.5, 103401.9, 103586.6, 103762.8, 
    103955.5, 104095.9, 103807.4, 103881.5, 104151.8, 103938.6, 103417.9, 
    103175.7,
  102214.1, 102386.4, 102736.4, 103040.6, 103353.3, 103395.6, 103762.7, 
    103932.7, 104045.2, 104196.7, 104238.6, 104278.1, 104202.2, 102184.5, 
    102809.8,
  102102.3, 102269.1, 102626.6, 102961.2, 103193.6, 99820.82, 103592.5, 
    103999.3, 104161.2, 104234.6, 104293.2, 104332.1, 104330.9, 104284.5, 
    104179,
  102023.8, 102165.7, 102539.1, 102853.9, 103260.8, 103182.2, 99665.33, 
    103614.1, 104032.3, 104203.5, 104329.6, 104349.8, 104384.5, 104375.5, 
    104326.7,
  101953, 102110.8, 102473.4, 102803.1, 103145.5, 103446.8, 103410.1, 
    97432.34, 96833.93, 103866.9, 104314, 104338, 104413.4, 104369.2, 104384,
  101917.8, 102090.1, 102434.4, 102770, 103051.2, 103246.8, 103549.2, 
    103601.5, 103552.9, 104033.5, 104202.4, 104311.6, 104392.8, 104410.3, 
    104413.9,
  101958.4, 102130.6, 102447.1, 102741.9, 103025.1, 103211.5, 103370.1, 
    103615.9, 103784, 103911.6, 104102.2, 104266.4, 104356.5, 104402.4, 104404,
  102010.8, 102193.3, 102463, 102740.4, 102954.5, 103129.2, 103300.3, 
    103394.5, 103542.2, 103785.7, 104040.7, 104198.9, 104326.5, 104399, 
    104446.3,
  102075.1, 102254.1, 102486.2, 102719.8, 102935.7, 103098.9, 103242, 
    103390.9, 103521.4, 103702.6, 103966.4, 104140.9, 104283.7, 104380.6, 
    104458.7,
  102083.9, 102236.4, 102454.2, 102685.2, 102875.5, 103017.9, 103179.8, 
    103279, 103395.3, 103607.3, 103895.3, 104081.8, 104239.6, 104372.3, 
    104477.4,
  102968.5, 103160.6, 103404.4, 103522.8, 103672.1, 103746.2, 103750.1, 
    103744.6, 103680.4, 103243.1, 103167.5, 103272.7, 102959, 102360.7, 
    102081.7,
  102918.8, 103093.1, 103336.6, 103534.5, 103732.3, 103634.2, 103845.9, 
    103819, 103735, 103703.2, 103567.8, 103445.4, 103228.2, 101138.1, 101674.3,
  102861.6, 103060.4, 103298.2, 103537.7, 103595.9, 100129.6, 103785.4, 
    104002.6, 103963.8, 103835.9, 103713.9, 103579.1, 103414, 103242.2, 
    103041.6,
  102810.4, 103009.6, 103263.6, 103455.2, 103745.3, 103569.3, 99880.36, 
    103685.7, 103866.9, 103929.6, 103851.3, 103704.6, 103564.6, 103410, 
    103247.5,
  102758.1, 102965.2, 103220, 103398.8, 103623.6, 103828.7, 103742.4, 
    97520.19, 96799.41, 103723.3, 103960.4, 103815.8, 103717.8, 103531, 
    103449.2,
  102727, 102915.4, 103145.9, 103343.8, 103530.6, 103656.3, 103843.4, 
    103833.9, 103711.7, 103940.8, 103993.7, 103926.6, 103851.4, 103723.7, 
    103621.2,
  102676.3, 102855.9, 103073.7, 103244.1, 103436, 103568.8, 103703.3, 
    103806.9, 103911.1, 103949.6, 104015.1, 104026.2, 103971.6, 103892.9, 
    103815,
  102625.5, 102775.8, 102971.7, 103142.8, 103314.9, 103432.8, 103564.1, 
    103658.4, 103734, 103891.3, 104039.5, 104084.7, 104096.3, 104061.6, 
    104024.5,
  102525.8, 102674.2, 102868.3, 103022.9, 103185.8, 103323.9, 103437.2, 
    103557.9, 103697.6, 103825, 104023.6, 104125, 104180.3, 104196.7, 104192.7,
  102407.9, 102520.1, 102700.9, 102879.7, 103063.4, 103176.8, 103316.1, 
    103416.5, 103516.2, 103699.6, 103955.9, 104122.5, 104228.5, 104300, 
    104328.6,
  103828.1, 103860.8, 103953.7, 103879.3, 103895.7, 103802, 103650.5, 
    103528.5, 103380.5, 102831.4, 102722, 102826.5, 102567.1, 102021, 101766.4,
  103768.9, 103787.6, 103859.4, 103875.6, 103923.1, 103620.6, 103765.5, 
    103550.1, 103387.1, 103261.8, 103079.7, 102966.2, 102806.1, 100781.3, 
    101350.2,
  103702.4, 103767.3, 103813.8, 103884.4, 103751.7, 100191.9, 103601.4, 
    103809, 103620.3, 103413.1, 103211.4, 103081.8, 102956.2, 102850, 102682.1,
  103637, 103701.2, 103772.9, 103814.8, 103882.4, 103590.8, 99810.02, 
    103428.6, 103562.9, 103540.9, 103376.5, 103218.3, 103103.6, 103001.5, 
    102880.3,
  103567.6, 103641.5, 103730.7, 103762.4, 103827.4, 103810.9, 103649.9, 
    97399.87, 96731.63, 103456, 103563, 103380.9, 103302.7, 103155.5, 103091.6,
  103443.2, 103531.8, 103611, 103683.5, 103728.3, 103744.7, 103745.4, 
    103726.3, 103572.8, 103762.9, 103695.1, 103569.1, 103490.5, 103387.5, 
    103292.3,
  103253.6, 103354.8, 103455.4, 103545.9, 103619.9, 103677, 103711.3, 
    103769.6, 103882.3, 103863.6, 103817.1, 103748.4, 103672.3, 103599.5, 
    103507.5,
  102999.5, 103087.1, 103195.1, 103315.9, 103426.2, 103527.1, 103603.8, 
    103644, 103738.1, 103884.7, 103933.9, 103893, 103854.8, 103795.6, 103726.2,
  102689, 102759.2, 102871.8, 103049.4, 103219.6, 103369, 103475.8, 103589.5, 
    103740.6, 103920, 104005, 104021.5, 104004.6, 103974.6, 103913.6,
  102347.1, 102375.8, 102452.7, 102662.4, 102945.5, 103171.8, 103350.6, 
    103459.7, 103604.3, 103825.5, 104001.3, 104099.8, 104126.3, 104127.8, 
    104073.6,
  104309.2, 104264.7, 104244.9, 104149.1, 104154.9, 104097.1, 103942.7, 
    103812.8, 103673.4, 103185.6, 103093.6, 103161.3, 102826.4, 102199.7, 
    101861.8,
  104193.5, 104169.9, 104088.2, 104039.3, 104083.5, 103869.4, 104019, 
    103859.4, 103708.6, 103605.2, 103438.7, 103288.1, 103045.2, 100925.3, 
    101379.8,
  104050.8, 104074.8, 104027.6, 104012.3, 103841.2, 100363.6, 103857.5, 
    104009, 103871.4, 103734.3, 103564.3, 103406.2, 103198.4, 102976.5, 
    102667.5,
  103889.9, 103933.5, 103951.1, 103918.7, 103877, 103678.8, 99996.54, 
    103733.4, 103876.9, 103830, 103705.6, 103529.4, 103339.7, 103112.9, 
    102820.3,
  103731.7, 103770.4, 103803.2, 103799.1, 103821.7, 103816, 103822, 97610.8, 
    96937.23, 103701.9, 103837.6, 103659.1, 103494.2, 103236.1, 103004.4,
  103508.1, 103558.1, 103617, 103665.7, 103690, 103731.1, 103854.9, 103940.9, 
    103800.3, 103976.9, 103918.4, 103796.1, 103631.7, 103409.3, 103167.3,
  103219.2, 103326.2, 103377.4, 103463.9, 103537.6, 103637.7, 103750.1, 
    103951.6, 104040, 104025.6, 103990.4, 103910.2, 103770.1, 103572.9, 
    103337.7,
  102802.4, 102947.8, 103103.5, 103260, 103347.9, 103479.3, 103617.5, 
    103777.2, 103895.7, 104003, 104040.1, 103991.4, 103897.6, 103736.1, 103534,
  102616.9, 102652.6, 102726, 102875.8, 103084.9, 103292.9, 103453.3, 
    103610.7, 103765.1, 103941.4, 104028.3, 104043.7, 103990.5, 103868.3, 
    103690,
  102722.2, 102683.4, 102643.2, 102670.7, 102796.5, 103027.3, 103257.9, 
    103413.8, 103554.4, 103741.6, 103941, 104026, 104036.5, 103973.9, 103836.7,
  104226.1, 104281.9, 104324.6, 104238.4, 104264.7, 104307.1, 104293, 
    104218.9, 104073.2, 103545, 103362.1, 103321.6, 102853.2, 102112.4, 
    101715.2,
  104166.2, 104200.7, 104151.2, 104073.2, 104149.8, 104075, 104262.1, 104194, 
    104056.7, 103928.7, 103690.1, 103437.2, 103065.2, 100861.9, 101239,
  104056.8, 104142.5, 104150.6, 104083.2, 103934.2, 100506.6, 104035, 
    104262.8, 104162.6, 104003.8, 103780.6, 103526.7, 103208.3, 102910.4, 
    102535,
  103922.4, 104036.3, 104082.2, 104061.7, 103972.1, 103834, 100106.4, 
    103868.3, 104037.9, 104030.8, 103869.7, 103615.8, 103338, 103031.4, 
    102698.3,
  103773, 103891.7, 103962, 103988.1, 103933.4, 103895.5, 103893.3, 97734.18, 
    97016.82, 103816.3, 103928.8, 103694.8, 103471.2, 103155.1, 102885.9,
  103602.4, 103729.6, 103803.3, 103856.3, 103839.6, 103795.9, 103881.1, 
    103929.6, 103823.5, 103994.2, 103923.5, 103755.8, 103563.4, 103303.4, 
    103031.4,
  103377.1, 103529.6, 103619.8, 103705.7, 103738.3, 103737.5, 103749, 
    103844.7, 103946.9, 103953.6, 103882.3, 103772.3, 103625, 103421.5, 
    103170.7,
  103127, 103315.5, 103421.9, 103526.9, 103560.7, 103589.8, 103604.9, 103659, 
    103697.8, 103766.5, 103771.1, 103718.2, 103629, 103493.5, 103307,
  102884.5, 103044.8, 103166.5, 103275.5, 103356.3, 103412, 103422.9, 
    103462.5, 103510.2, 103538.7, 103565.4, 103575.4, 103557.6, 103496.5, 
    103372.3,
  102777.8, 102872.5, 102942.7, 103024.4, 103080, 103130.7, 103174.1, 
    103200.1, 103225.2, 103245.3, 103318.7, 103368.4, 103397, 103410.4, 
    103362.6,
  102873.3, 103161.6, 103462.9, 103712.8, 103920.3, 104055.1, 104104, 
    104141.4, 104083.2, 103639.4, 103553.8, 103583.8, 103190.3, 102506.4, 
    102166.3,
  102965.5, 103195, 103452.3, 103677.1, 103860.5, 103836.2, 104051.3, 
    104047.5, 103988.1, 103951.9, 103824.3, 103656.9, 103379.4, 101230.4, 
    101667.1,
  103014.3, 103210.1, 103417.7, 103648.1, 103711.5, 100257.2, 103828.8, 
    104081.6, 104049.1, 103942.6, 103824.7, 103674.5, 103447, 103211, 102918.7,
  103058.7, 103236.1, 103422.4, 103580.6, 103752.5, 103601.2, 99929.71, 
    103663.4, 103805.8, 103851.2, 103799.5, 103662.3, 103461.7, 103244.8, 
    102986.9,
  103094.5, 103266, 103440.9, 103575.2, 103677.9, 103755.1, 103665.2, 
    97565.35, 96834.14, 103536.7, 103742.6, 103603.9, 103434.1, 103215, 103052,
  103093.8, 103269.4, 103417, 103546.5, 103615.6, 103652.7, 103682.9, 
    103635.6, 103490.9, 103651.3, 103634, 103520.8, 103371.8, 103186.2, 
    103049.7,
  103063.1, 103229.7, 103364.5, 103480.1, 103554.3, 103600.3, 103584.8, 
    103559.1, 103526.9, 103509.2, 103466.3, 103382.1, 103250.1, 103120.3, 
    103007.6,
  102993.4, 103151.7, 103261.4, 103362.1, 103400, 103430.3, 103430.2, 
    103401.4, 103347.2, 103311, 103262.5, 103190, 103104.6, 103027.4, 102958.9,
  102879.9, 103015.7, 103110.9, 103191, 103231.1, 103245.1, 103221.1, 
    103198.7, 103153.3, 103103.4, 103052.2, 102998.2, 102940.4, 102898.1, 
    102852.7,
  102709.5, 102825.6, 102896.1, 102946.2, 102956.6, 102960.6, 102950.4, 
    102917.3, 102868.4, 102808.6, 102803.1, 102776.1, 102746.9, 102730.6, 
    102713.4,
  102067.3, 102302.3, 102630.2, 102941.8, 103285.7, 103564.2, 103730.3, 
    103857, 103904.6, 103519.8, 103458, 103523.7, 103105.5, 102396, 102107.5,
  102063, 102278.6, 102602.6, 102958.5, 103269, 103385.8, 103723, 103828.8, 
    103784.7, 103778, 103642.6, 103498.3, 103206.1, 101079.7, 101632.3,
  102008, 102257.2, 102584.5, 102973.3, 103152.1, 99864.4, 103550.5, 
    103843.1, 103835.2, 103714.1, 103581, 103427.2, 103187.1, 103000.8, 
    102899.9,
  101969.5, 102226.3, 102568.8, 102904.1, 103258.2, 103189.8, 99653.16, 
    103441.5, 103635.3, 103600, 103535.9, 103368.9, 103165.6, 103004.6, 
    102983.3,
  101964.1, 102223.7, 102566.2, 102886.6, 103195, 103477.4, 103385.4, 
    97375.17, 96658.69, 103363.1, 103486.7, 103334.6, 103161.9, 102974.7, 
    103011.6,
  101982.8, 102247.6, 102556.5, 102861.5, 103103.7, 103312.5, 103543.8, 
    103508, 103437.3, 103524.9, 103430.1, 103299.3, 103144.4, 102991.1, 
    102956.1,
  102027.2, 102289.9, 102580.4, 102842.5, 103087.6, 103261.2, 103403.1, 
    103505.7, 103516.7, 103440.8, 103352.2, 103240.2, 103105.2, 102975.9, 
    102915,
  102088.2, 102335.1, 102583, 102812.2, 102996.2, 103168.4, 103292.5, 
    103350.4, 103339.3, 103317.4, 103246.1, 103156.4, 103047.8, 102937.5, 
    102859.8,
  102171.6, 102391.2, 102606.6, 102802.6, 102962.3, 103085.5, 103163, 
    103218.3, 103201.6, 103158.2, 103096, 103017.6, 102929.1, 102843.5, 
    102777.7,
  102242, 102416, 102580, 102729.8, 102846.6, 102940.7, 103000.1, 103005.5, 
    102978.4, 102919.8, 102890.2, 102829.7, 102758.7, 102700.1, 102646.5,
  102315.4, 102574.7, 102857, 103100.8, 103356.3, 103547.2, 103648.7, 
    103700.9, 103618, 103137.4, 103049.8, 103245.3, 103069.7, 102555.1, 
    102288.9,
  102295.6, 102546.5, 102837.4, 103121.7, 103348.4, 103381.8, 103665.6, 
    103708.1, 103605.4, 103506, 103333, 103250.5, 103182.2, 101182.6, 101741.8,
  102251.9, 102529.7, 102792.4, 103101, 103217.6, 99840.76, 103527.6, 
    103773.6, 103709.2, 103548.5, 103407.7, 103263.6, 103167.7, 103084.6, 
    102926.9,
  102217.8, 102479.6, 102729.9, 102990.6, 103275.2, 103185.2, 99605.99, 
    103400.6, 103610.5, 103555.1, 103475, 103323.8, 103169.9, 103060.4, 
    102948.5,
  102178.4, 102414.7, 102645.6, 102898.9, 103140.8, 103405.8, 103341.9, 
    97318.23, 96647.69, 103394.6, 103521.3, 103385.4, 103231.6, 103050.2, 
    102950.1,
  102126.9, 102337.2, 102535.9, 102777.9, 102984.8, 103194.2, 103427.9, 
    103444.6, 103395.5, 103614.2, 103539.1, 103426.8, 103278.3, 103089.5, 
    102943.6,
  102042.3, 102231.7, 102420.6, 102640.7, 102865.9, 103066.2, 103247.9, 
    103440.7, 103571.7, 103585.4, 103536.9, 103441, 103302.7, 103119, 102935.3,
  101951.8, 102113.1, 102290.5, 102497.9, 102698.3, 102908.5, 103098.9, 
    103236.6, 103369.9, 103475.1, 103487.7, 103414.6, 103287.9, 103127.8, 
    102948.2,
  101869.6, 102012.4, 102185.3, 102376.3, 102573.9, 102763.1, 102949.3, 
    103131.1, 103263.8, 103348.8, 103370, 103324.9, 103230.3, 103083.2, 
    102927.9,
  101829, 101957.3, 102115.3, 102280.3, 102453.1, 102627.4, 102795.2, 
    102936.1, 103047.9, 103127.9, 103205.1, 103194.9, 103122.5, 103014.6, 
    102890.9,
  102862, 103056.2, 103268.4, 103405.2, 103557.1, 103624.7, 103620.3, 
    103541.5, 103413.7, 102880.9, 102733.1, 102702.1, 102237.2, 101546.9, 
    101323.7,
  102841.3, 103021.8, 103227.9, 103414.2, 103544, 103467.8, 103643.5, 
    103541.8, 103411.5, 103266.3, 103057.1, 102824.1, 102476.6, 100351.5, 
    100932.7,
  102768.8, 102972.5, 103147.8, 103358.7, 103374.2, 99878.82, 103432.9, 
    103639.4, 103507.6, 103309.2, 103135.3, 102920.9, 102623.6, 102399, 
    102271.1,
  102681, 102881.5, 103053.5, 103213.4, 103387.6, 103243.2, 99524.21, 
    103163.1, 103350.8, 103315.1, 103191.9, 103003.6, 102747.9, 102549.1, 
    102447.4,
  102589.9, 102773.8, 102938.5, 103080.7, 103205.2, 103309.8, 103216.4, 
    97134.6, 96372.83, 103064.3, 103234.7, 103069.9, 102867.9, 102622.1, 
    102601.7,
  102474.2, 102652, 102802.7, 102939.7, 103028.4, 103096.9, 103169.6, 
    103143.2, 103035, 103232.8, 103211.4, 103114.8, 102964.3, 102754.2, 
    102707.8,
  102367, 102529.3, 102659.1, 102774.3, 102854.3, 102914.5, 102949.1, 103020, 
    103067.9, 103103.3, 103154, 103126.9, 103020.3, 102829.1, 102767.6,
  102255.2, 102388.2, 102496.4, 102599.6, 102659, 102714.7, 102758.9, 
    102778.5, 102820.9, 102934.8, 103039, 103079.6, 103053.8, 102917.5, 102834,
  102141.2, 102258.5, 102339.9, 102411.9, 102474.5, 102523, 102562.5, 
    102643.4, 102692.9, 102772.5, 102892.7, 102995.2, 103020.5, 102945.1, 
    102837.8,
  102037.4, 102101.3, 102160.3, 102213.7, 102250.3, 102298.9, 102350.4, 
    102387.4, 102458.8, 102530.2, 102712.8, 102857.6, 102938, 102943.6, 
    102860.9,
  103046.7, 103179.9, 103321.9, 103388.1, 103456.4, 103402.6, 103288.8, 
    103196.4, 103085.9, 102658, 102671.1, 102940.2, 102828.3, 102369.1, 
    102157.2,
  103108.6, 103232.1, 103361.5, 103451.5, 103456.3, 103203.4, 103314.3, 
    103125.1, 103010, 103020.8, 102995, 103044.2, 103056.8, 101102.2, 101801.8,
  103110.3, 103251.4, 103337.5, 103443.1, 103290.3, 99743.12, 103102.5, 
    103277.1, 103121.8, 103060.9, 103034.3, 103117.6, 103195.3, 103265.5, 
    103211.4,
  103094.5, 103226.1, 103290.8, 103327.4, 103315.6, 103069.5, 99267.49, 
    102788.4, 102911.4, 103053.5, 103069.1, 103137.8, 103246.8, 103379.6, 
    103383.6,
  103058.7, 103150.9, 103207.8, 103212.8, 103189.4, 103116.9, 102897.9, 
    96830.1, 96084.48, 102706.5, 103094.5, 103123.9, 103291.6, 103375.9, 
    103478.4,
  102942.5, 103042.1, 103072.3, 103083.6, 103022.5, 102968.5, 102890.8, 
    102779.6, 102596.4, 102808, 103043.5, 103095.8, 103270.5, 103401.4, 
    103493.4,
  102837.7, 102888.9, 102911.9, 102904.9, 102861.2, 102795.4, 102730.1, 
    102722.9, 102716.5, 102746.9, 102954.1, 103065.2, 103212.8, 103374.5, 
    103485.8,
  102708, 102735.5, 102725.9, 102718.5, 102661.5, 102621.2, 102593.4, 102572, 
    102590.4, 102669.7, 102861.5, 103004.9, 103137.7, 103320.6, 103460.4,
  102540.5, 102578.3, 102579.5, 102552.2, 102519.6, 102500.7, 102491, 
    102516.6, 102556, 102601.5, 102730.7, 102946.5, 103072.7, 103219.9, 
    103387.9,
  102347.6, 102379.6, 102386.2, 102382.6, 102372.8, 102366.3, 102367.5, 
    102338, 102354, 102417.7, 102585.9, 102801.4, 102974.1, 103126.8, 103230.6,
  103667.3, 103709.7, 103729.4, 103650.1, 103553.1, 103410.3, 103218.3, 
    103225.4, 103328.2, 103037.4, 103117.1, 103357.1, 103090.8, 102396.2, 
    101992.4,
  103682.3, 103712, 103710, 103642.3, 103506.5, 103139.9, 103181.1, 102991.7, 
    103079.5, 103255.6, 103321, 103340.8, 103219.6, 101068.7, 101524.1,
  103644.2, 103691.7, 103655.3, 103633.1, 103319.6, 99728.31, 102899.8, 
    103035, 103040.6, 103144.7, 103195.4, 103273.6, 103218.6, 103090.1, 
    102804.6,
  103573.9, 103640.2, 103619.2, 103547.4, 103370.8, 102987.4, 99118.8, 
    102555.6, 102809.9, 103029.5, 103122.8, 103173.8, 103185.8, 103106.2, 
    102877.3,
  103513.3, 103552.7, 103543.9, 103437.6, 103293.9, 103086.4, 102750.3, 
    96701.6, 95944.53, 102588.6, 103034.4, 103072.9, 103161.3, 103041.9, 
    102940.3,
  103387.8, 103430.3, 103411.6, 103314.6, 103159.2, 102981.5, 102832, 
    102667.7, 102486.6, 102718.6, 102936.7, 103003.1, 103087.7, 103043.7, 
    102954,
  103264.2, 103272.7, 103251.7, 103184, 103075.9, 102910, 102776, 102719.6, 
    102696.5, 102694.8, 102843.9, 102935.3, 103014.7, 103008.5, 102938.1,
  103159.8, 103164.5, 103129.8, 103075.7, 102949, 102824, 102734.8, 102642.3, 
    102599.9, 102634.2, 102747.8, 102828.7, 102919.9, 102970.9, 102948.1,
  102982.8, 103004.7, 102983.2, 102933.7, 102844.1, 102756.7, 102684.7, 
    102636.5, 102596, 102556.3, 102611.3, 102710.9, 102812, 102902.2, 102917.1,
  102779.7, 102806.9, 102811.4, 102774.9, 102710.6, 102667.4, 102616.8, 
    102538.2, 102465.5, 102393, 102421.4, 102518.9, 102655.2, 102803.4, 
    102888.8,
  103850.7, 103922.2, 103945, 103866.1, 103721.8, 103484.5, 103159, 102961, 
    102820, 102364.8, 102300.2, 102417, 102131.7, 101470.8, 101123.1,
  103761.4, 103818.7, 103821.1, 103762.3, 103602.6, 103182.4, 103154.2, 
    102846.6, 102669, 102581.1, 102460, 102354.2, 102202, 100118.3, 100586.6,
  103611, 103697.4, 103676.1, 103636.2, 103357, 99744.48, 102868.9, 102980.2, 
    102767.2, 102547.7, 102381.8, 102282.2, 102166.2, 102032.8, 101793.8,
  103471.1, 103551.7, 103540.2, 103494.5, 103359.4, 102966.5, 99122.48, 
    102479, 102518.3, 102465.8, 102325.5, 102212.4, 102126.5, 102024.5, 
    101824.5,
  103304.1, 103370.8, 103381.1, 103323.9, 103223.2, 103059.5, 102734.2, 
    96655.23, 95815.66, 102152.5, 102275.1, 102138, 102082.5, 101972.8, 101863,
  103186.8, 103196.8, 103186.5, 103145.9, 103029.4, 102910.6, 102781.3, 
    102548.8, 102258.8, 102306.6, 102201, 102092.4, 102028.9, 101979.7, 
    101877.3,
  103065.5, 103058.1, 103020.6, 102963.5, 102885.4, 102774.5, 102633, 
    102529.4, 102394.2, 102225.6, 102109.2, 102024, 101949.4, 101964.6, 
    101887.7,
  102899.4, 102887, 102843.8, 102789.6, 102692.6, 102591.6, 102471.1, 
    102322.6, 102190.7, 102117.8, 102034.2, 101947.4, 101896.1, 101960.3, 
    101919.1,
  102665, 102667.7, 102618.9, 102557.4, 102480.6, 102387.2, 102275, 102199.5, 
    102098, 102005.3, 101940.5, 101873.5, 101824.6, 101929.2, 101933.4,
  102439, 102414.5, 102363.7, 102319, 102221.5, 102131.5, 102047.4, 101937.6, 
    101851.2, 101802.7, 101825.8, 101796.8, 101748.6, 101871, 101948.7,
  103578, 103660.5, 103739.6, 103742.9, 103727.9, 103637.3, 103451.9, 
    103270.8, 103044.5, 102409.8, 102196.2, 102185.8, 101810.9, 101260, 
    101212.9,
  103410, 103469.4, 103497.3, 103520.2, 103476.2, 103196.3, 103248.1, 
    102957.9, 102701.2, 102527.6, 102277.2, 102070.6, 101847.4, 99876.09, 
    100667.2,
  103163.8, 103233.8, 103247, 103246.9, 103068.1, 99528.12, 102717.8, 
    102875.6, 102595.6, 102338.1, 102100.8, 101920.8, 101728.9, 101687.9, 
    101859.7,
  102995.6, 103009.6, 102994.9, 102967.5, 102880.3, 102580.7, 98790.79, 
    102115.5, 102199.1, 102121.6, 101916.1, 101736.7, 101597.4, 101629.8, 
    101865.2,
  102837.5, 102814.6, 102787.6, 102712, 102628.6, 102496.6, 102190.7, 
    96162.55, 95272.59, 101579.6, 101718.1, 101532.7, 101441.9, 101479.7, 
    101788.3,
  102700.6, 102631.6, 102534.3, 102447.4, 102292.1, 102167.8, 102015.9, 
    101786.2, 101504.5, 101572.2, 101431.8, 101315.4, 101263, 101370.3, 101702,
  102509.5, 102433.1, 102305.2, 102170.5, 102009.4, 101829.9, 101648, 
    101520.8, 101361.9, 101206.7, 101110.6, 101059.4, 101047.6, 101237.5, 
    101609.1,
  102236.6, 102120.9, 101948.7, 101806, 101605.6, 101441.3, 101257.8, 
    101090.3, 100956.8, 100895.3, 100810.7, 100780.4, 100829, 101118.3, 
    101554.8,
  101912.5, 101812.4, 101654.8, 101491.7, 101303.5, 101112.5, 100923.6, 
    100845.5, 100717.8, 100609.7, 100534, 100535.8, 100618.9, 100995.6, 
    101476.5,
  101637.6, 101507.8, 101337.9, 101179.7, 100958.2, 100781.1, 100683.8, 
    100545.3, 100411, 100319.2, 100292.6, 100331.5, 100462.9, 100908.6, 
    101415.1,
  102847.8, 102916.6, 103006.2, 103051.1, 103109, 103112.5, 103058, 103004.1, 
    102892.3, 102350, 102176.8, 102175.1, 101782.4, 101161.2, 101008.5,
  102585.7, 102635.2, 102695.9, 102764.6, 102801.4, 102633.8, 102764.6, 
    102583.7, 102388.9, 102237, 102024.1, 101783.1, 101554.3, 99559.16, 
    100260.8,
  102210.7, 102262, 102341.5, 102399, 102328.9, 98893.01, 102172.4, 102387.1, 
    102179.1, 101869.7, 101601.5, 101381.8, 101199.6, 101124.2, 101294.5,
  101823.5, 101876.3, 101955.7, 102013.6, 102064.1, 101860.8, 98167.88, 
    101526.4, 101557.7, 101445.4, 101200.8, 101001.3, 100939.9, 100893.4, 
    101240,
  101378.9, 101467, 101562.3, 101638.6, 101700.9, 101714.6, 101522.7, 
    95573.28, 94636.77, 100800.7, 100919.8, 100760.4, 100723.2, 100690.5, 
    101176.1,
  100899.3, 101005.1, 101120, 101229.7, 101281, 101314, 101290.1, 101093, 
    100812.2, 100830, 100703.8, 100611.6, 100542, 100568.9, 101138.2,
  100388.6, 100498.4, 100633.3, 100785.9, 100875.6, 100924.7, 100903.7, 
    100876.5, 100738.9, 100633.4, 100562, 100500.1, 100389.1, 100522.6, 
    101184.6,
  99937.68, 100002.3, 100107.4, 100288.8, 100416.1, 100530.6, 100562.6, 
    100536.2, 100510.7, 100524.3, 100451.6, 100395.6, 100302.9, 100555.5, 
    101280.5,
  99521, 99553.77, 99653.82, 99838.8, 100026, 100183.8, 100257.7, 100345, 
    100360.7, 100367.9, 100322.6, 100304.7, 100293.4, 100705, 101445.3,
  99159.09, 99145.91, 99225.46, 99405.06, 99610.88, 99815.99, 99961.91, 
    100072.9, 100139.4, 100192, 100211.7, 100238.7, 100385.2, 100887.5, 
    101531.2,
  101439, 101570.2, 101780.2, 101971.7, 102200.2, 102383.5, 102505.1, 
    102630.7, 102716.7, 102375.4, 102368.1, 102500.4, 102166.4, 101453.8, 
    101031.1,
  101009.8, 101121.1, 101338.1, 101556.3, 101790.4, 101819.7, 102145.5, 
    102239.5, 102279.7, 102376.3, 102340.3, 102268.2, 102086.3, 99959.77, 
    100411.9,
  100415.8, 100615, 100850.4, 101088.2, 101263.8, 98015.41, 101456.6, 101996, 
    102014.7, 102019.1, 102011.9, 101957.7, 101838.8, 101683.9, 101660.2,
  99899.41, 100091.8, 100348.1, 100562.3, 100857.6, 100838.2, 97445.66, 
    101082.9, 101554.3, 101674.7, 101719.2, 101654.8, 101637.5, 101596.4, 
    101768.8,
  99486.94, 99661.64, 99855.02, 100083.7, 100304, 100617.5, 100653.6, 
    95021.98, 94279.92, 100894.5, 101392.5, 101369.6, 101442.8, 101479.4, 
    101792.8,
  99209.64, 99340.76, 99456.8, 99612.22, 99773.03, 99978.74, 100307, 
    100392.1, 100480.7, 100973.4, 101087.4, 101164.3, 101290.8, 101478.1, 
    101820.4,
  99081.93, 99151.56, 99174.73, 99222.6, 99319.52, 99464.31, 99687.24, 
    100045.1, 100355.3, 100609.2, 100821.1, 100990.4, 101179.6, 101497.7, 
    101859.1,
  99044.73, 99041.7, 98965.03, 98921.07, 98897.24, 98987.54, 99165.36, 
    99420.09, 99776.75, 100228.3, 100567.5, 100812.9, 101110.1, 101524.9, 
    101933.4,
  99084.45, 99020.41, 98872.49, 98733.05, 98611.27, 98592.38, 98715.34, 
    99009.27, 99376.88, 99829.11, 100269, 100626.4, 101034.1, 101545.8, 
    102013.5,
  99155.59, 99023.45, 98821.36, 98615.36, 98383.07, 98233.92, 98291.94, 
    98545.89, 98946.53, 99429.63, 99992.58, 100451.9, 100974.4, 101566.5, 
    102042.4,
  100051.4, 100376.4, 100805, 101163.6, 101573, 101945.2, 102247.2, 102563.7, 
    102853.9, 102717.1, 102919.5, 103278.9, 103161.9, 102677.9, 102448.5,
  99718.92, 100030.5, 100450.2, 100887, 101298.4, 101520.8, 102021.4, 
    102304.3, 102547.7, 102824.5, 102995.9, 103141.2, 103197.1, 101246.6, 
    101879.8,
  99350.23, 99677.2, 100113.2, 100588.2, 100937.4, 97823.4, 101538.4, 
    102187.2, 102397.7, 102574.9, 102734.5, 102913.4, 103023, 103086, 103103.5,
  99003.02, 99361.84, 99783.64, 100203.3, 100759.2, 100806.7, 97564.94, 
    101471.6, 102040.7, 102296.2, 102512.6, 102642.6, 102847.8, 102956, 
    103104.6,
  98789.85, 99102.15, 99536.95, 99964.09, 100465.7, 100933.4, 100974, 
    95346.34, 94789.91, 101529.1, 102205.8, 102323.5, 102605.7, 102757.2, 
    103014.7,
  98935.91, 99001, 99365.5, 99755.54, 100178.6, 100542.8, 100934.9, 100989.6, 
    101080, 101624.1, 101836.5, 102025.1, 102331.9, 102591, 102887.4,
  99204.07, 99187.12, 99379.93, 99671.82, 100045.5, 100346.7, 100607, 
    100929.3, 101174.8, 101329.5, 101525.5, 101774.5, 102079.3, 102413.7, 
    102782.8,
  99509.89, 99439.94, 99465.11, 99625.92, 99851.39, 100082, 100305.4, 
    100501.3, 100712.3, 101030.2, 101312.6, 101571.1, 101901.1, 102273.6, 
    102715.6,
  99940.8, 99824.79, 99769.68, 99804.75, 99891.66, 99964.66, 100034.5, 
    100203.7, 100419.6, 100697.1, 101027.4, 101365.5, 101728, 102160.7, 
    102662.6,
  100269.6, 100209.4, 100156.8, 100110.3, 100051.9, 100015.1, 99939.05, 
    99921.28, 100035.3, 100290.9, 100721.6, 101144.9, 101577.2, 102072.1, 
    102617.6,
  100310, 100662.6, 101071.4, 101431.7, 101889.8, 102316.1, 102692.9, 103118, 
    103484, 103368.4, 103602.9, 103983.3, 103875.1, 103437.7, 103286.7,
  100216.8, 100543.1, 100960.1, 101376.5, 101801.1, 102091.8, 102644.6, 
    103045, 103354.2, 103676.9, 103868.8, 104023.3, 104071, 102105.2, 102885.7,
  100085.9, 100434.7, 100850.6, 101315.3, 101623.5, 98542.49, 102438, 
    103069.9, 103401.9, 103618.8, 103829.4, 103995.6, 104119.2, 104179, 
    104221.6,
  99955.05, 100305.7, 100724.8, 101157.8, 101673, 101697, 98547.7, 102614.4, 
    103231.8, 103551.2, 103789.9, 103923.3, 104099.4, 104200.8, 104338.6,
  99864.38, 100209.1, 100609.8, 101047.1, 101505.2, 101979.6, 102036.9, 
    96488.73, 96077.12, 103088.2, 103694.7, 103823.6, 104039.4, 104123.6, 
    104310.9,
  99818.57, 100149.1, 100507.1, 100926.9, 101348.3, 101723.1, 102188.7, 
    102315.8, 102483.6, 103191.6, 103484.7, 103695.4, 103910.6, 104069.9, 
    104230.9,
  99830.46, 100097.9, 100445.6, 100812, 101237.3, 101592.5, 101934.3, 
    102386.3, 102746.8, 102993.5, 103258.9, 103519.1, 103740.3, 103950.7, 
    104126.9,
  99929.55, 100148.7, 100411, 100738.5, 101094, 101438.7, 101773.8, 102030.6, 
    102317.2, 102716.9, 103048, 103305.9, 103562.9, 103810.6, 104041.6,
  100119.1, 100236.7, 100424.7, 100693.3, 101002.2, 101297.8, 101591.4, 
    101927.6, 102220.1, 102533.3, 102826.9, 103114.4, 103382.5, 103658.8, 
    103932.5,
  100479.5, 100498.7, 100561.3, 100717.5, 100937.2, 101169.8, 101421.1, 
    101667.2, 101928.8, 102240.8, 102621.5, 102933.8, 103210.4, 103520.3, 
    103828.2,
  101502.2, 101848.5, 102254.5, 102630, 103035.1, 103359.7, 103617, 103895.8, 
    104085.6, 103859.8, 104010.9, 104353.4, 104191.8, 103703.8, 103488.8,
  101566.2, 101913.7, 102323.6, 102744.7, 103108.2, 103290.6, 103770.8, 
    103991.5, 104114.3, 104319, 104402.6, 104518.9, 104464.7, 102487.6, 
    103145.1,
  101585, 101988.2, 102397.5, 102853, 103035.5, 99891.08, 103729.8, 104198.6, 
    104376, 104464.8, 104541.4, 104653.8, 104694.2, 104682.1, 104587.1,
  101578.2, 101991, 102413.4, 102826.7, 103266.7, 103224.9, 99947.38, 
    103938.1, 104348.8, 104548.2, 104686.1, 104748.1, 104826.2, 104854.1, 
    104803.3,
  101572, 101986.9, 102408.9, 102824.5, 103226.6, 103669, 103646.7, 97775.12, 
    97329.95, 104400.5, 104802.9, 104834.8, 104932, 104908.2, 104942.6,
  101542.3, 101956.3, 102354.2, 102784.4, 103158.5, 103534.2, 103930, 
    104020.7, 104080.9, 104655.6, 104798.4, 104898.4, 104986.6, 105006.5, 
    105012.2,
  101525.7, 101934.8, 102337.2, 102747.5, 103138.6, 103507, 103802.2, 
    104182.6, 104476.1, 104659.1, 104798.9, 104945.1, 105007.1, 105042.5, 
    105026.4,
  101487.9, 101882.1, 102273.1, 102676.6, 103053.7, 103427.8, 103755.4, 
    103998.7, 104258.7, 104585.4, 104788.9, 104929.9, 105018.7, 105074.9, 
    105076.2,
  101479.9, 101873, 102269.2, 102662.5, 103022.5, 103367.7, 103681.5, 
    104001.6, 104271.5, 104537.6, 104735, 104896.7, 104991.9, 105060.9, 
    105071.1,
  101458.7, 101828.3, 102209.9, 102596.4, 102966.2, 103308.4, 103600.5, 
    103847.5, 104094.2, 104375.4, 104627.1, 104812.4, 104932.2, 105024.4, 
    105064.6,
  102520, 102833.7, 103196.6, 103515.4, 103847.8, 104070.7, 104196.1, 
    104308.4, 104335.9, 103953.8, 103960, 104164.4, 103934.9, 103392.1, 
    103177.5,
  102579.6, 102911.9, 103293.3, 103683.1, 103958.1, 104018.9, 104382.2, 
    104432, 104417.4, 104467.6, 104407.2, 104390, 104232.7, 102197.6, 102829.1,
  102644.1, 103049.7, 103429.3, 103849.1, 103908.6, 100626.4, 104347.6, 
    104707.2, 104745.1, 104684.1, 104624.7, 104580, 104502.1, 104401.5, 104253,
  102726.3, 103143.5, 103540, 103885.2, 104227.3, 104057.8, 100618.7, 
    104482.9, 104760.2, 104854.3, 104840.9, 104739.7, 104680.3, 104580.6, 
    104473.7,
  102843.4, 103247.5, 103627.5, 103949.3, 104254.4, 104609.2, 104429.5, 
    98353.45, 97830.88, 104796.9, 105038.2, 104908.4, 104866.6, 104704.5, 
    104658,
  102971.6, 103347.6, 103692.2, 104018.1, 104268.7, 104523.5, 104832.8, 
    104808.3, 104783.9, 105152.8, 105155.3, 105088.6, 105008.7, 104888, 
    104777.6,
  103098.8, 103455.5, 103787.4, 104090.8, 104378.5, 104607.6, 104786.9, 
    105077.7, 105258.1, 105279.6, 105298.4, 105255.4, 105154.9, 105037.6, 
    104904.1,
  103208, 103547.4, 103876, 104159.4, 104413.6, 104660.9, 104887.4, 105060.2, 
    105220.4, 105392.9, 105436.5, 105390.3, 105302.6, 105178.4, 105039.2,
  103336.1, 103676.4, 103994.7, 104271.1, 104526.4, 104753.7, 104968.6, 
    105205.6, 105405.8, 105512, 105527, 105499, 105413.3, 105300, 105149.6,
  103428.5, 103754.7, 104066.8, 104344.8, 104599.7, 104829.8, 105040, 
    105219.1, 105397.1, 105496.1, 105567.5, 105552, 105487.3, 105399.2, 
    105272.7,
  103579.6, 103805.6, 103984.6, 104082.4, 104167.7, 104186.6, 104148.4, 
    104173, 104173.3, 103840.1, 103902.2, 104202.2, 104038, 103550.3, 103357.8,
  103589.4, 103834.7, 104034.6, 104228.9, 104294.6, 104122.5, 104324.5, 
    104250.2, 104179.7, 104219.6, 104215.9, 104249.4, 104193.2, 102169.8, 
    102828.2,
  103581.3, 103897.8, 104108.7, 104352.1, 104213.6, 100742.2, 104286.6, 
    104504.3, 104473.8, 104365, 104304.9, 104290.3, 104264.1, 104200.8, 
    104097.5,
  103567.4, 103898.6, 104152.3, 104349.2, 104521.3, 104236, 100583.1, 
    104293.4, 104407.7, 104473.2, 104415.1, 104330.7, 104287.9, 104219.8, 
    104164.4,
  103579.2, 103920.6, 104201.8, 104386.9, 104526.6, 104688.9, 104421.6, 
    98171.65, 97631.75, 104391, 104577.1, 104423.9, 104393.8, 104266.1, 104273,
  103578.1, 103942.9, 104224.9, 104466.9, 104600.1, 104713.8, 104865.5, 
    104792.4, 104592.3, 104769.8, 104701.1, 104582.4, 104506.2, 104417.3, 
    104376,
  103598.5, 103992.2, 104298, 104543.6, 104733.8, 104860.1, 104916.5, 105033, 
    105075.9, 104992.8, 104889.4, 104792.7, 104691.6, 104610.7, 104546,
  103619.7, 104012, 104342.9, 104621.4, 104821.8, 105010.9, 105141.1, 
    105187.7, 105198, 105191, 105105.6, 105001.8, 104904.2, 104820.5, 104761.8,
  103678.2, 104077.8, 104436.3, 104723.4, 104963.1, 105139.6, 105283.8, 
    105400.5, 105447.3, 105400.5, 105319.8, 105232.6, 105129, 105033.3, 
    104951.6,
  103719.6, 104117, 104479, 104790.8, 105054.5, 105278.2, 105453.6, 105541.5, 
    105552.9, 105496.2, 105484.5, 105445, 105354, 105266.1, 105177.4,
  103949.9, 103989.2, 104068, 104105.7, 104204.5, 104284.5, 104352, 104455.6, 
    104533.5, 104224.3, 104300.5, 104589.8, 104377.2, 103878.5, 103658.4,
  103965, 104031.6, 104107.9, 104210.8, 104279.3, 104162, 104412.7, 104456.3, 
    104469.5, 104594.8, 104642.2, 104713.6, 104647.5, 102654.5, 103339,
  103949, 104078.2, 104128.7, 104286.7, 104145.7, 100627.5, 104256.4, 
    104536.9, 104609.1, 104624, 104672.7, 104742.6, 104786.4, 104763.5, 
    104716.9,
  103943, 104051.6, 104116.1, 104212.2, 104319.2, 104084.4, 100378.4, 
    104205.9, 104458.3, 104589.2, 104700.1, 104743.1, 104820.8, 104861.1, 
    104897.9,
  103973.8, 104051.9, 104099.8, 104143, 104198.3, 104341.2, 104177.1, 
    98011.18, 97421, 104347.3, 104711.7, 104731.3, 104837.4, 104835.8, 104958,
  103995.7, 104088.3, 104123.5, 104184.2, 104215.6, 104271.4, 104390.3, 
    104386.8, 104217.2, 104589.1, 104680.1, 104746.9, 104851.3, 104922.5, 
    105009.4,
  104038.2, 104163.4, 104235.6, 104310.3, 104354.6, 104399.3, 104424.9, 
    104542.1, 104646, 104674.9, 104742.5, 104834.1, 104912, 105001.6, 105071.7,
  104092.9, 104262.7, 104374.6, 104475.4, 104525.1, 104581.7, 104633.2, 
    104663.9, 104715.8, 104801.1, 104871.9, 104945.1, 105030.1, 105111.1, 
    105176.6,
  104179, 104385.7, 104551.6, 104684.5, 104767.2, 104818.3, 104861.7, 
    104941.5, 105003.6, 105027, 105064.3, 105120.5, 105188, 105259.5, 105314.8,
  104256.7, 104508.1, 104719, 104882.8, 104988.9, 105073.3, 105123.5, 
    105144.6, 105173.8, 105188, 105279.2, 105341.9, 105391.5, 105453.1, 
    105494.2,
  104110.3, 104189.1, 104300.8, 104350.7, 104441.5, 104455.3, 104384.8, 
    104382.8, 104380.2, 104036.8, 104108.5, 104420.7, 104298.4, 103887.6, 
    103742,
  104097.1, 104197.3, 104316.3, 104440.4, 104514.7, 104327.9, 104516.9, 
    104452.4, 104405.4, 104484.7, 104496.2, 104587.3, 104547.5, 102665, 
    103408.4,
  104038.4, 104190.8, 104317, 104518, 104392.9, 100874.7, 104473.4, 104719.2, 
    104737.1, 104686.7, 104691.8, 104739.3, 104797.1, 104832.3, 104831.1,
  103977.8, 104135.8, 104292.4, 104440.2, 104639.6, 104338.4, 100717.7, 
    104497.2, 104734.6, 104840.5, 104900.2, 104893, 104966.5, 105036.7, 
    105094.2,
  103934.8, 104067.4, 104236.9, 104398.4, 104523.5, 104750.1, 104521.6, 
    98358.59, 97833.09, 104775.3, 105094.7, 105060.5, 105150.4, 105154.8, 
    105301.3,
  103884.3, 104023.7, 104146.5, 104328.1, 104441.2, 104602.5, 104844.9, 
    104782, 104654.7, 105103.7, 105180.2, 105223.4, 105299.1, 105358.6, 
    105455.6,
  103844.2, 103946.1, 104088.8, 104256.9, 104421.3, 104596.7, 104712.3, 
    104948.4, 105137.3, 105206.3, 105292.5, 105385.9, 105463.9, 105547.2, 
    105629.6,
  103802.3, 103929, 104062.8, 104223, 104360.1, 104561.8, 104754.4, 104878.2, 
    105061.9, 105271.6, 105411, 105514.6, 105621.7, 105733.9, 105843.9,
  103833.6, 103961.3, 104087.8, 104245.6, 104406.6, 104582.7, 104759, 
    105014.4, 105259.9, 105388.8, 105503.6, 105629.2, 105763.1, 105893.2, 
    106001.6,
  103926.5, 104062.5, 104190, 104318.6, 104451.2, 104636.7, 104839.8, 
    105028.7, 105238.4, 105381.5, 105573.9, 105738, 105890, 106034.8, 106152.1,
  104294.9, 104329.4, 104400.2, 104405, 104450.1, 104438.5, 104414.9, 
    104505.4, 104593.5, 104254.6, 104315.1, 104633.3, 104513.4, 104073.2, 
    103940.7,
  104232.1, 104270.6, 104318.2, 104375.2, 104373.5, 104212.9, 104428.9, 
    104479.4, 104512.1, 104622.4, 104690, 104801.8, 104817.8, 102923.1, 
    103732.6,
  104090.5, 104173, 104221.8, 104306.3, 104202.5, 100637.8, 104299.9, 
    104612.5, 104735.1, 104733.3, 104805.2, 104930.3, 105083, 105191.6, 
    105277.6,
  103969.5, 104031.9, 104099.8, 104133.9, 104293.5, 104066.3, 100469.8, 
    104305.8, 104643.2, 104799.1, 104969.8, 105073.9, 105293.2, 105496.8, 
    105607.8,
  103863.7, 103929.7, 103987.4, 104033.4, 104111.2, 104386.5, 104210.7, 
    98200.62, 97637.49, 104683.2, 105112.7, 105229.8, 105464.2, 105613, 
    105868.1,
  103793.5, 103885.4, 103918.1, 103967.9, 104042, 104212.3, 104492.2, 
    104453.7, 104387.4, 104950.2, 105162.8, 105365, 105594.8, 105788.4, 
    106003.1,
  103739.6, 103843.2, 103913.1, 103960.3, 104079.8, 104216.8, 104364.1, 
    104639.8, 104860.3, 104986.4, 105217.1, 105465.2, 105685.6, 105892.1, 
    106089.3,
  103691.9, 103822, 103928.8, 103989, 104080.4, 104235.7, 104405.3, 104497.3, 
    104717.8, 104997.5, 105276.5, 105517.6, 105763.8, 105981.1, 106187,
  103653.6, 103808.7, 103961.1, 104068.3, 104188, 104286.2, 104438, 104663.4, 
    104913.7, 105095.9, 105321.2, 105562.8, 105808.6, 106034.9, 106230.3,
  103595.8, 103761.8, 103948.5, 104085.9, 104209.4, 104345.8, 104500.2, 
    104654.2, 104874.6, 105059.3, 105334.1, 105581, 105827.7, 106061.4, 
    106247.9,
  104194.1, 104193, 104216.1, 104159.8, 104143.8, 104062.5, 103984.3, 
    104010.6, 104104, 103866.9, 104049.9, 104475.4, 104441.9, 104125.3, 
    104046.6,
  104126.5, 104135.1, 104141.6, 104145.3, 104136.7, 103902.1, 104078.3, 
    104011.8, 104048.1, 104220.5, 104360.2, 104559.2, 104672.5, 102833.2, 
    103675.4,
  103951.9, 104016.1, 104039.3, 104080.9, 103981.5, 100365.4, 103975.3, 
    104186.5, 104226.7, 104289.2, 104417.2, 104608, 104807.6, 104946.2, 
    105090.8,
  103772.9, 103840.2, 103884.4, 103904.3, 104001.3, 103840.4, 100079.2, 
    103940.4, 104194.1, 104348, 104534.4, 104696.8, 104928, 105171.7, 105349.2,
  103601.6, 103661.6, 103717.9, 103748.5, 103789.4, 103960.3, 103930.2, 
    97681.84, 97153.17, 104242.9, 104677.8, 104803.9, 105059.2, 105225.4, 
    105521.2,
  103434.7, 103483.6, 103535, 103592, 103639, 103764.7, 103994.6, 104066.6, 
    103964.5, 104498.3, 104721.9, 104913.6, 105160.1, 105370.5, 105600.3,
  103262.3, 103320.9, 103354.1, 103430.7, 103504.2, 103645.6, 103814, 
    104073.9, 104326.3, 104533.5, 104739.5, 104995.4, 105212.7, 105436.8, 
    105637.4,
  103092.7, 103157.1, 103195.9, 103272.7, 103349.1, 103502, 103724, 103928.4, 
    104181.5, 104480.6, 104753.7, 105017.8, 105253.7, 105487.5, 105693,
  102968.2, 103036.9, 103066.4, 103147.7, 103243.7, 103394.6, 103589.3, 
    103852.7, 104182.8, 104479.1, 104731.4, 105000.4, 105241.6, 105479.9, 
    105676.2,
  102858.8, 102942.8, 103014.6, 103087.8, 103171.1, 103314.9, 103504.9, 
    103731, 104061.2, 104344, 104650, 104925.1, 105175.3, 105423.9, 105623.6,
  103912.8, 103979, 104032.9, 104000.4, 104040.5, 104050.6, 104110.6, 
    104266.7, 104438.5, 104214.1, 104407.3, 104797, 104724.3, 104351.5, 
    104248.5,
  103768.6, 103862.5, 103937.1, 103956.1, 104035.6, 103887.5, 104148.2, 
    104219.9, 104364.4, 104535.9, 104686.6, 104835.7, 104914.7, 102987.6, 
    103780.7,
  103517.5, 103684, 103786.7, 103876.4, 103802.2, 100286.7, 103965.6, 
    104279.6, 104417, 104526.6, 104665.8, 104802.8, 104945.3, 105017, 105105.6,
  103221.5, 103449.2, 103573, 103680.9, 103749, 103670.4, 99929.32, 103912.7, 
    104279.3, 104448, 104626.1, 104749.1, 104919.8, 105078, 105221.3,
  102944.3, 103199.5, 103359.2, 103486.4, 103511.1, 103557.7, 103685.8, 
    97488.48, 96953.84, 104052.9, 104568.1, 104672.1, 104892.4, 104988.9, 
    105207.1,
  102663.5, 102939.1, 103118.9, 103285.9, 103356.1, 103362.5, 103535.2, 
    103762.6, 103649.2, 104132, 104384.8, 104570.7, 104797.6, 104965.2, 
    105149.7,
  102396.7, 102690.6, 102899.8, 103089.2, 103182.5, 103242.5, 103276.5, 
    103511.9, 103771.3, 103966.3, 104189.8, 104460.3, 104672.6, 104868.8, 
    105048.4,
  102140, 102443, 102668.2, 102875.3, 102997.8, 103090, 103148.1, 103289.5, 
    103516.8, 103810.1, 104064.6, 104313.7, 104539.6, 104758.3, 104965,
  101937.5, 102252.5, 102490.7, 102685, 102811.5, 102917.4, 102981.8, 
    103120.4, 103358.8, 103653.4, 103912.5, 104162.1, 104395.4, 104614.8, 
    104823.3,
  101768.5, 102070.3, 102301.5, 102490.6, 102626.1, 102749.1, 102843, 
    102967.1, 103186.5, 103440.3, 103728.9, 103988.5, 104221.3, 104465.2, 
    104679.1,
  102734.3, 103001.9, 103336.5, 103571.8, 103788.9, 104000.9, 104198.1, 
    104363.7, 104542.6, 104289.1, 104414.6, 104748.9, 104622.9, 104214.9, 
    104082.2,
  102500.4, 102738.5, 103102.5, 103392.6, 103657.3, 103746.3, 104137.9, 
    104281.4, 104412.5, 104587.8, 104692.4, 104773.8, 104812.3, 102819.6, 
    103603.9,
  102180.8, 102478.7, 102873.9, 103224.5, 103400.3, 100047.3, 103896.9, 
    104345.1, 104484.3, 104540, 104644.2, 104739.2, 104814.1, 104874.2, 
    104921.9,
  101794.9, 102159.3, 102565.4, 102951.1, 103362.8, 103347.1, 99836.62, 
    103863.4, 104289, 104462.4, 104605.9, 104678.3, 104789.6, 104895.2, 
    105016.5,
  101417.4, 101816.2, 102260.1, 102696.1, 103093.6, 103493.2, 103519.3, 
    97517.63, 96924.37, 103965.9, 104522.1, 104585.4, 104751.5, 104809.6, 
    104996.6,
  101096.1, 101481.8, 101922.2, 102411, 102815, 103161.6, 103514.7, 103609.3, 
    103587.8, 104047.6, 104295.8, 104453.8, 104647.2, 104773.6, 104913.3,
  100800.1, 101186.8, 101652.1, 102153.1, 102590.5, 102960.6, 103215.4, 
    103530.6, 103753.6, 103851.8, 104052.7, 104292.2, 104487.6, 104650.2, 
    104793.9,
  100559.8, 100916.1, 101363.3, 101886, 102326.2, 102724.9, 103015.7, 
    103214.3, 103413.3, 103667.2, 103901.1, 104123.5, 104322.1, 104501.9, 
    104662.8,
  100371, 100727.1, 101185.7, 101692.6, 102144.2, 102536.4, 102838.9, 103078, 
    103281.4, 103468.9, 103689, 103928.4, 104125.5, 104305.7, 104473.7,
  100232.7, 100547, 100980.8, 101491.9, 101941.3, 102338.1, 102656.9, 
    102888.1, 103065.1, 103234.8, 103462.5, 103691.6, 103900.9, 104101.8, 
    104274.6,
  101503.2, 101603.3, 101849.8, 102216.1, 102590.6, 102933.8, 103184.5, 
    103414.2, 103600, 103368.5, 103510.3, 103918, 103841.4, 103493.1, 103397.1,
  101253.6, 101377, 101634.6, 102044.5, 102420, 102641.5, 103096.7, 103311.8, 
    103446.7, 103676.7, 103784.4, 103944.4, 104023.6, 102092.4, 102897.7,
  100952.2, 101110.3, 101445.9, 101893.4, 102159.4, 98942.05, 102848.1, 
    103382.3, 103561.3, 103648, 103766.6, 103907.1, 104054, 104144.5, 104219.9,
  100683.5, 100811.7, 101205.6, 101645, 102135.4, 102150.4, 98834.71, 
    102884.3, 103372.3, 103589.7, 103758.5, 103858.8, 104025.8, 104173.9, 
    104322.5,
  100441.9, 100553.7, 100934.4, 101414.1, 101895, 102380.7, 102402, 96631.14, 
    96084.91, 103193.6, 103729.2, 103808, 104010.6, 104092.8, 104312.7,
  100256.3, 100338.7, 100662.1, 101157, 101607.8, 102062.7, 102523.1, 
    102620.3, 102694.1, 103329.9, 103579.9, 103746.9, 103944.3, 104089.5, 
    104266.8,
  100080.4, 100149.3, 100435.1, 100932.9, 101415.5, 101865, 102244.6, 
    102736.5, 103058.2, 103206.3, 103414.6, 103658, 103857.4, 104032.1, 
    104189.1,
  99960.6, 100014.7, 100239.1, 100725.3, 101176.4, 101653.4, 102051.6, 
    102394.2, 102706, 103040.9, 103323.9, 103558.3, 103766.2, 103958.1, 104128,
  99898.88, 99932.29, 100118.2, 100598.5, 101043.9, 101496.9, 101890.6, 
    102304.1, 102674.3, 102954.5, 103207.3, 103447.1, 103655, 103848.7, 
    104015.9,
  99910.28, 99907.87, 100049.7, 100465, 100906.4, 101347.9, 101734.3, 
    102096.4, 102481.1, 102783, 103072.4, 103309, 103520.9, 103721, 103891.2,
  100708.2, 100602.6, 100582.7, 100736.4, 101048.5, 101380.9, 101650.2, 
    101935.6, 102214.6, 102091.9, 102315.5, 102773.4, 102722.2, 102404.4, 
    102329.7,
  100498.5, 100377.8, 100387.3, 100614.6, 100994.8, 101166.4, 101643.9, 
    101885.2, 102118.4, 102380.3, 102563.1, 102764.3, 102882.5, 100993.4, 
    101816,
  100281.4, 100156.8, 100214.8, 100511.7, 100788.2, 97609.75, 101480, 
    101991.9, 102212.7, 102375, 102534.6, 102722.8, 102894.8, 103018.6, 
    103121.8,
  100054.8, 99954.93, 100016.3, 100344, 100781.4, 100817.4, 97509.61, 
    101590.4, 102075, 102323.6, 102523.6, 102678, 102883, 103074.6, 103236.2,
  99815.18, 99772.21, 99807.21, 100165.5, 100593.6, 101025, 101074.1, 
    95346.08, 94840.7, 101988.2, 102517.6, 102646.8, 102869.9, 102997.5, 
    103232,
  99610.56, 99603.66, 99616.02, 99961.7, 100391, 100799.5, 101230.6, 
    101386.2, 101484.9, 102145.9, 102414.4, 102618.2, 102842.6, 103015.9, 
    103204.4,
  99450.7, 99469.38, 99463.06, 99773.45, 100237.2, 100659.1, 101046.7, 
    101517.8, 101851.6, 102062.7, 102313.4, 102583.3, 102795.2, 102990.5, 
    103157.6,
  99395.54, 99411.27, 99371.24, 99637.97, 100099.2, 100525.9, 100922.3, 
    101294.8, 101606.8, 101974, 102279.2, 102547.4, 102771.7, 102974.5, 
    103144.8,
  99383.8, 99354.18, 99301.6, 99553.62, 100050.7, 100468.2, 100862.2, 101251, 
    101636.3, 101960.8, 102234.8, 102504, 102730, 102939.6, 103112.2,
  99393.2, 99303.12, 99248.07, 99551.05, 100044.3, 100416, 100789.4, 
    101172.6, 101562.2, 101872.7, 102190.2, 102462.1, 102685.1, 102904.5, 
    103085.8,
  99867.93, 99921.52, 100033, 100122.8, 100261.8, 100422.4, 100628.5, 
    100889.8, 101213, 101159.7, 101453.8, 101920.1, 101856.3, 101447.4, 
    101278.4,
  99530.75, 99604.08, 99758.73, 99896.12, 100078, 100189.9, 100629.3, 
    100838.5, 101104.2, 101444.4, 101679.4, 101910.7, 102023.9, 100094, 100830,
  99143.97, 99237.88, 99428.46, 99648.85, 99813.97, 96761.77, 100511.6, 
    101024.5, 101205.4, 101430.8, 101642.2, 101858.4, 102029.5, 102119.2, 
    102177.4,
  98808.94, 98907.12, 99084.11, 99342.16, 99732.41, 99824.95, 96621.56, 
    100617, 101123.7, 101386, 101612.1, 101802.9, 102020, 102199.5, 102310.8,
  98501.77, 98601.58, 98788.12, 99059.38, 99505.54, 99928.38, 99988.44, 
    94388.58, 93923.08, 101027.8, 101609.1, 101759.1, 102011.3, 102136.5, 
    102347.6,
  98271.64, 98344.7, 98528.79, 98821.31, 99270.46, 99745.88, 100104.7, 
    100245.7, 100371.3, 101140.2, 101480, 101719.4, 101989.8, 102168, 102359.3,
  98211.87, 98233.64, 98382.45, 98667.94, 99141.48, 99641.69, 99994.1, 
    100390.1, 100727.4, 101052.8, 101377.8, 101704.4, 101957.2, 102170.5, 
    102344.5,
  98238.72, 98270.78, 98379.96, 98662.52, 99121.3, 99581.28, 99965.95, 
    100281.1, 100627.2, 101061.7, 101396.5, 101709.5, 101962.7, 102191.5, 
    102368.1,
  98380.3, 98395.19, 98510.27, 98774.51, 99234.82, 99639.07, 100007.4, 
    100375.3, 100776.6, 101127.9, 101441.3, 101735.5, 101979.1, 102198.2, 
    102370.5,
  98529.79, 98565.74, 98696, 98975.49, 99396.82, 99741.23, 100118, 100482.3, 
    100884.9, 101173.6, 101496.9, 101772.8, 102002.9, 102216.9, 102388.3,
  99539.72, 99563.6, 99652.27, 99744.77, 99887.99, 100033.7, 100170.7, 
    100341.9, 100547.1, 100451.5, 100772.8, 101311.9, 101371.3, 101084, 
    100975.1,
  99192.59, 99231.55, 99344.41, 99476.48, 99615.67, 99649.31, 100004.4, 
    100147.8, 100354.2, 100672.8, 100947.8, 101255.6, 101475.2, 99612.24, 
    100346.3,
  98861.69, 98892.7, 99031.38, 99222.29, 99323.53, 96170.95, 99750.77, 
    100216.5, 100388.6, 100636.2, 100901.3, 101190.1, 101426.4, 101546, 
    101576.1,
  98632.57, 98647.28, 98751.74, 98979.59, 99284.66, 99303.27, 96047.91, 
    99871.64, 100347.7, 100632.4, 100882.5, 101143, 101403.6, 101574, 101585.7,
  98408.2, 98428.48, 98530.59, 98764, 99122.38, 99499.16, 99526.56, 93929.32, 
    93415.54, 100356.4, 100930.8, 101124.9, 101400.2, 101514.9, 101614.7,
  98243.81, 98240.07, 98337.62, 98622.98, 98997.47, 99369.77, 99711.02, 
    99796.13, 99860.33, 100527.7, 100845.3, 101117.7, 101397.8, 101542.3, 
    101625,
  98146.73, 98159.77, 98234.74, 98556.36, 98979.19, 99332.91, 99617.23, 
    99971.26, 100196.8, 100448, 100784.9, 101131.4, 101392.2, 101568.7, 101631,
  98135.73, 98160.47, 98258.97, 98648.59, 98993.9, 99351.94, 99622.72, 
    99847.86, 100099.2, 100489.8, 100830.3, 101171.8, 101423, 101617.9, 
    101685.6,
  98323.52, 98333.3, 98496.75, 98832.57, 99141.12, 99439.01, 99683.31, 
    99995.4, 100306.9, 100623.5, 100931.4, 101238.8, 101480.9, 101669.1, 
    101738.9,
  98837.12, 98790.72, 98896.74, 99129.02, 99335.96, 99590.23, 99867.42, 
    100188.4, 100480.3, 100741.7, 101036.6, 101334.9, 101550.5, 101735, 
    101802.9,
  100072.7, 100102.1, 100175.4, 100265, 100398.1, 100527.5, 100608.6, 
    100721.1, 100829.5, 100586.4, 100719.8, 101091.1, 101062, 100828.4, 
    100914.2,
  99716.95, 99748.09, 99827.89, 99948.54, 100047.7, 100038.4, 100345.2, 
    100441.4, 100525.6, 100686.2, 100782.5, 100959.3, 101114, 99403.55, 
    100300.6,
  99375.43, 99355.21, 99422.86, 99560.19, 99642.89, 96440.2, 99859.12, 
    100319.8, 100367.7, 100490.6, 100626.9, 100824.8, 101044.9, 101256.2, 
    101516.8,
  99163.98, 99083.56, 99081.81, 99159, 99401.87, 99413.68, 96072.98, 
    99757.03, 100218.6, 100366.2, 100536.3, 100726.1, 101024.2, 101313.6, 
    101601.3,
  99056.21, 98934.2, 98893.7, 98927.77, 99113.62, 99446.52, 99508.88, 
    93928.21, 93333.06, 100065.5, 100547.9, 100710.6, 101032.6, 101263.5, 
    101621.3,
  99074.99, 98894.2, 98787.45, 98804.73, 98950.43, 99298.72, 99643.61, 
    99713.31, 99764.02, 100299.2, 100497.7, 100750.5, 101077.7, 101332.1, 
    101646.5,
  99216.65, 99038.7, 98851.38, 98843.82, 99084.22, 99418.68, 99668.35, 
    99959.24, 100129.6, 100280.1, 100518, 100828.7, 101126, 101385.5, 101634.2,
  99431.89, 99355.08, 99294.89, 99303.16, 99439.83, 99608.22, 99789.32, 
    99928.11, 100141.5, 100396.1, 100634, 100932.5, 101203.3, 101459.1, 
    101659.9,
  99622.84, 99586.24, 99546.42, 99580.9, 99665.94, 99805.74, 99955.8, 
    100176.2, 100398, 100555.5, 100793.8, 101052.5, 101290.9, 101507.2, 
    101641.3,
  99842.53, 99783.9, 99789.88, 99823.65, 99888.9, 99995.59, 100152.4, 100348, 
    100529.3, 100681.1, 100918.6, 101162.5, 101371.3, 101542.8, 101617.4,
  100618, 100592.6, 100570.2, 100592.7, 100668.8, 100802, 100886.5, 101025.4, 
    101191.9, 101001.2, 101189.9, 101598.1, 101561.9, 101264.4, 101216.5,
  100424.9, 100341.9, 100267.1, 100274.3, 100319.1, 100325.6, 100638.8, 
    100767.3, 100889.2, 101100.8, 101244.5, 101413.2, 101521, 99742.28, 
    100507.3,
  100353.8, 100203.3, 100059.1, 99984.11, 99943.11, 96716.49, 100159.1, 
    100636.9, 100734.5, 100883.2, 101035.1, 101210.2, 101366.6, 101501, 
    101653.6,
  100344.2, 100150.6, 99951.65, 99779.59, 99776.74, 99749.21, 96335.45, 
    100038.8, 100509.7, 100692.5, 100870, 101018.8, 101226.4, 101434, 101641.3,
  100371.1, 100191.7, 99984.91, 99756.82, 99671.18, 99806.17, 99833.83, 
    94157.84, 93539.2, 100185.8, 100735.5, 100872.2, 101126.4, 101308.1, 
    101622.3,
  100415.8, 100271.8, 100055.6, 99877.48, 99692.65, 99742.94, 99968.38, 
    99954.07, 99906.52, 100287.4, 100529.7, 100769.2, 101057.5, 101312.8, 
    101630.9,
  100490.6, 100418.8, 100283.5, 100148.7, 100046.7, 99981.73, 100032.6, 
    100137.1, 100189.5, 100199.5, 100451.5, 100743.4, 101054.1, 101352.5, 
    101686.6,
  100532, 100514, 100436.1, 100356.5, 100262.9, 100230.7, 100229.5, 100212.5, 
    100234.2, 100327.6, 100536.6, 100814.6, 101129.7, 101459.9, 101803.6,
  100588.3, 100622.5, 100594.8, 100548.6, 100504.4, 100468, 100455.6, 
    100523.5, 100538, 100551.6, 100722.7, 100964.1, 101276.1, 101612.1, 
    101944.2,
  100657.7, 100701.4, 100720.4, 100701.3, 100664.2, 100647.8, 100667.3, 
    100707.8, 100733.6, 100772.3, 100937.6, 101171.4, 101453.1, 101774.2, 
    102069.3,
  101630.1, 101557.7, 101447.6, 101315.9, 101172.7, 101074.2, 101021.3, 
    101056.8, 101147, 100914.8, 101043.6, 101389.6, 101311.2, 101039.7, 
    101030.5,
  101605.5, 101530.5, 101412.4, 101269.6, 101082.7, 100780.6, 100929.3, 
    100906.1, 100954.1, 101113, 101203.4, 101319.6, 101400.7, 99610.41, 
    100412.6,
  101599.2, 101537.1, 101420.2, 101285.1, 100975.6, 97442.48, 100722.3, 
    100928.9, 100913.1, 100957, 101054.5, 101190.5, 101325.5, 101464.8, 
    101607.8,
  101591.6, 101549.3, 101444.2, 101287.9, 101140.2, 100797.6, 97075.26, 
    100604.5, 100845.2, 100888.1, 100953.9, 101060.9, 101231, 101436.8, 
    101620.8,
  101573.2, 101574.2, 101497.5, 101355, 101204.9, 101062.2, 100843.5, 
    94789.48, 94034.33, 100521.5, 100840, 100930.6, 101142.4, 101307.2, 
    101574.9,
  101550.9, 101565.1, 101493, 101380.1, 101220.8, 101100.8, 101027.1, 
    100891.1, 100661.9, 100713.9, 100718.3, 100835.2, 101066.9, 101276.4, 
    101534.1,
  101518.8, 101552.9, 101491.2, 101374.3, 101230.5, 101102.9, 101020.6, 
    101005.8, 100876.7, 100672.9, 100669.5, 100829.1, 101032.6, 101265.8, 
    101521.6,
  101500.6, 101511, 101414.9, 101300, 101161.7, 101054.7, 100990.6, 100963.4, 
    100880.9, 100766.9, 100731.5, 100868.3, 101067.1, 101315.7, 101585.7,
  101470.1, 101454.7, 101348.7, 101217.4, 101112, 101013.5, 100955.9, 
    101014.8, 100969.5, 100843.1, 100813.4, 100947.8, 101140.7, 101410.6, 
    101703.7,
  101421.3, 101317.2, 101183.9, 101101.1, 100997.2, 100925.5, 100918.4, 
    100967, 100959.1, 100876.3, 100897, 101045.2, 101254.9, 101545.3, 101805.4,
  102874.6, 102880.3, 102879, 102793, 102666.3, 102482.2, 102237, 102052.9, 
    101886, 101411, 101426.3, 101648.9, 101484.3, 101036.2, 100896.1,
  102843, 102844.2, 102794.3, 102675.2, 102489.9, 102075.2, 102090.3, 
    101777.3, 101586.7, 101539.5, 101499.9, 101516.8, 101497.7, 99578.39, 
    100236.1,
  102771.6, 102774.8, 102662.2, 102540.1, 102162.3, 98563.86, 101558.6, 
    101739, 101487.6, 101373.5, 101339.9, 101372.1, 101370.4, 101389.7, 
    101389.2,
  102675.9, 102633.7, 102503.1, 102295, 102032.6, 101557.7, 97721.52, 
    100934.1, 101152.3, 101217, 101245, 101242.5, 101284.2, 101326.9, 101401.7,
  102569.2, 102505.9, 102340.9, 102087.9, 101785.7, 101467.9, 101071.7, 
    95105.04, 94305.59, 100816.9, 101183.4, 101140.1, 101196.5, 101243.3, 
    101400.3,
  102489.5, 102369.4, 102123.5, 101849.9, 101504.8, 101228.7, 101026.8, 
    100861.5, 100745.6, 101050.8, 101106.1, 101100.1, 101111.9, 101209.2, 
    101381.6,
  102394.5, 102217.1, 101944.4, 101675.9, 101351.5, 101112.7, 100989.3, 
    100961.6, 100973.3, 101048.4, 101090.2, 101092.3, 101075.1, 101202.4, 
    101379.5,
  102276.9, 102065.4, 101772.8, 101511.8, 101195.4, 101071.2, 101013.7, 
    100861.5, 100885.7, 101067.5, 101118, 101101, 101109.1, 101244, 101420,
  102184.9, 101953.2, 101683.2, 101446.4, 101197.4, 101132.3, 101071.5, 
    100966.7, 101017.9, 101110.8, 101126.5, 101146.6, 101187.9, 101335.9, 
    101512.1,
  102105, 101843.5, 101584.7, 101381.3, 101162.8, 101133.6, 101129.8, 
    100957.6, 101014.1, 101084, 101152, 101217.3, 101286.1, 101445, 101591.6,
  102796.4, 102876, 102889.3, 102776, 102651.6, 102474.8, 102238.1, 102035.6, 
    101826.7, 101210.1, 100995.3, 101047.7, 100820.9, 100490.2, 100491.2,
  102851, 102840.9, 102763.6, 102613.6, 102438.6, 102016.6, 102111, 101771.3, 
    101516.4, 101300, 101000.4, 100833.1, 100778.1, 99047.38, 99890.6,
  102831.1, 102787.4, 102631.3, 102490.6, 102132.7, 98615.88, 101721.8, 
    101888.9, 101599, 101293, 100971.2, 100886.8, 100926.7, 101079.1, 101220.3,
  102790.1, 102707.4, 102547.9, 102382.9, 102224.5, 101844.4, 98128.26, 
    101422.7, 101463, 101413.4, 101234.2, 101190.2, 101257.7, 101374.4, 
    101451.7,
  102793.4, 102701.9, 102567.3, 102416.6, 102254.7, 102154.5, 101866.8, 
    95699.83, 94907.25, 101409.2, 101549.2, 101431.5, 101444.1, 101444.7, 
    101574.3,
  102794, 102699.1, 102572.7, 102461.7, 102262.6, 102162.9, 102092.7, 
    101929.2, 101650.9, 101783.5, 101708.6, 101616.9, 101573.8, 101567.9, 
    101659.2,
  102811.6, 102744.4, 102621.6, 102497.5, 102335.4, 102208.8, 102074.4, 
    102064.9, 102021.9, 101913.4, 101803.5, 101731.5, 101638.8, 101652.8, 
    101765,
  102858, 102771.7, 102634.2, 102503, 102308.7, 102188.2, 102089.8, 101975.1, 
    101930.7, 101941.2, 101893.1, 101813.8, 101758.6, 101817.2, 101892,
  102915.6, 102828.2, 102690.5, 102534.9, 102371.4, 102205.8, 102063, 
    101988.9, 101963.7, 101941.1, 101915.4, 101885.3, 101856.2, 101912, 
    101987.3,
  102948.9, 102820.4, 102668.3, 102488.9, 102283.6, 102128.1, 102007, 101857, 
    101761.8, 101787.2, 101866.4, 101921.4, 101940.9, 102003.5, 102055.3,
  102911.3, 103039.9, 103157.6, 103134.1, 103101.3, 102945.2, 102704.1, 
    102515.6, 102401.1, 101941.6, 101796, 101783.1, 101311.1, 100624.1, 
    100452.3,
  103014.7, 103128.2, 103196.8, 103169.1, 103081.1, 102666, 102734.7, 
    102359.1, 102164, 102221.8, 102109.4, 101921.5, 101608.6, 99468.09, 
    100028.6,
  103085.6, 103219.1, 103204.5, 103187, 102876.5, 99370.75, 102430.8, 
    102618.5, 102398.4, 102272.5, 102154, 102034.7, 101854.2, 101688.5, 
    101512.8,
  103143.8, 103207.5, 103186.1, 103121.8, 103047.8, 102617.2, 98829.99, 
    102017.9, 101995.3, 102186.2, 102184.1, 102092.2, 101995.5, 101926.4, 
    101844.7,
  103206.1, 103241.7, 103217.6, 103128.1, 103024.5, 102864.1, 102500.1, 
    96325.79, 95485.45, 101757.5, 102201.1, 102107.9, 102107.6, 102021.5, 
    102055.2,
  103206.1, 103236.5, 103205.9, 103158.7, 103017.9, 102846.3, 102658.6, 
    102358.4, 101929.5, 101952.5, 102067.4, 102087.9, 102119.7, 102134.3, 
    102153.5,
  103233.6, 103288.1, 103245.8, 103174.2, 103056.3, 102885.6, 102655.2, 
    102428.4, 102170.6, 101921, 101904.8, 102013.5, 102076.5, 102166.9, 
    102225.4,
  103252.7, 103287, 103255.8, 103179.1, 103029.5, 102863.4, 102662.9, 
    102378.8, 102047.5, 101815.2, 101736.6, 101858.1, 101974.6, 102131.6, 
    102231.8,
  103276.6, 103319.1, 103288.3, 103178, 103043.5, 102854.8, 102641.2, 102398, 
    102087.5, 101771.4, 101608.4, 101669.9, 101813.6, 102013.2, 102172,
  103278.3, 103276.6, 103227.4, 103123.7, 102948.8, 102769.3, 102575.9, 
    102290.6, 101953.8, 101616.1, 101455.8, 101476.5, 101607.3, 101833.2, 
    102045.1,
  103320.2, 103526, 103662.4, 103640.8, 103617.7, 103522.3, 103368, 103284.7, 
    103302.6, 102902.6, 102848.7, 102980.8, 102724.4, 102178.8, 101974.2,
  103442.1, 103598.3, 103692, 103692.2, 103667.2, 103390.8, 103480.5, 
    103229.6, 103115.3, 103238.7, 103185.1, 103138.7, 103001.7, 100989.7, 
    101656.3,
  103536.3, 103691.5, 103726.9, 103780.1, 103593.1, 100142.2, 103374.5, 
    103507.6, 103296.1, 103213.2, 103193.4, 103196.9, 103144.2, 103113.2, 
    103032,
  103597.2, 103700.5, 103758.1, 103794.3, 103818.9, 103498.2, 99757.32, 
    103147.3, 103135.3, 103149.7, 103129.6, 103175.9, 103169.2, 103193.6, 
    103161.5,
  103652.3, 103742.4, 103803.8, 103815, 103814.2, 103773.8, 103508.3, 
    97386.36, 96602.5, 102924.4, 103078.5, 103040.8, 103136.5, 103114.9, 
    103157,
  103672.6, 103755.3, 103786.3, 103820, 103778.4, 103715.6, 103650.4, 
    103458.8, 103145.8, 103153.7, 102997.7, 102895.2, 102948.7, 103005.7, 
    103060.8,
  103664.8, 103745.7, 103783.6, 103777.9, 103745.7, 103673.7, 103554.5, 
    103481.2, 103338, 103124.6, 102925.7, 102798.8, 102756.5, 102811, 102889,
  103631.8, 103678.8, 103693.5, 103702.6, 103624.8, 103540.5, 103438.4, 
    103299.1, 103146.2, 103003.2, 102831.3, 102681.8, 102577.2, 102596.6, 
    102664,
  103561.4, 103587.9, 103572.6, 103552.1, 103482.9, 103399.8, 103271.3, 
    103169.1, 103037.6, 102860.3, 102677.7, 102531.7, 102413.3, 102363.6, 
    102415,
  103442.2, 103423.3, 103382.8, 103352.2, 103250.9, 103153.3, 103037, 
    102894.8, 102740.6, 102574.6, 102460.2, 102330.7, 102224.1, 102141.5, 
    102146.6,
  103828.5, 104071.9, 104310, 104431, 104549.6, 104569.9, 104562, 104590.3, 
    104573.3, 104181.3, 104157.2, 104363.8, 104128, 103584.5, 103321.3,
  103944.8, 104149, 104345.8, 104449.5, 104524.7, 104370.5, 104549, 104383.9, 
    104270.5, 104285.3, 104239.8, 104212.1, 104148.6, 102105.2, 102671.5,
  104055.7, 104257.4, 104398.3, 104508, 104393.8, 100918.4, 104269.7, 
    104510.3, 104334.1, 104116.9, 104002.6, 103963.3, 103904.7, 103846.1, 
    103740.3,
  104116.7, 104278, 104375.3, 104430.1, 104469.5, 104207.6, 100432.8, 
    103819.9, 103944.5, 103942.8, 103787, 103662.7, 103602.2, 103549, 103485.9,
  104151.8, 104268.2, 104335, 104345, 104317.6, 104249.9, 103990.2, 97889.24, 
    96999.2, 103326.8, 103533.9, 103332.2, 103253.6, 103162.3, 103124.9,
  104119.3, 104194.9, 104183.7, 104171.2, 104069.2, 103979.1, 103852, 
    103615.7, 103286.2, 103320.1, 103157.5, 102982.2, 102864.8, 102735.6, 
    102673.6,
  104039.2, 104071.3, 104014.2, 103942.2, 103821.5, 103673, 103488.1, 
    103335.5, 103145.2, 102893.9, 102701.4, 102548.3, 102397.5, 102272.8, 
    102169.7,
  103889.6, 103845.8, 103733.4, 103621.1, 103442.4, 103260.9, 103056, 
    102826.6, 102594.3, 102420.2, 102236.2, 102048.9, 101894.4, 101771.7, 
    101679.5,
  103696.2, 103602.3, 103452.2, 103274.3, 103069.8, 102842.1, 102583.7, 
    102358.4, 102137.1, 101898.9, 101690, 101515.2, 101371.2, 101265.9, 
    101193.3,
  103387.4, 103217.6, 103012.5, 102799.9, 102536.9, 102282, 102036.9, 
    101777.4, 101532.9, 101293.3, 101142.5, 100994.6, 100877.3, 100809.2, 
    100780,
  104518.3, 104716.7, 104920.6, 105073.6, 105202, 105248.4, 105194.4, 
    105153.7, 104997.7, 104413.2, 104178.4, 104116.4, 103637.1, 102838.8, 
    102349.1,
  104465.5, 104624.2, 104802.9, 104952.3, 105029.7, 104881.1, 105017.2, 
    104811.3, 104562.6, 104382.5, 104090.7, 103791.4, 103456.7, 101243.5, 
    101491,
  104368.1, 104548.5, 104699.8, 104861.1, 104790.8, 101281.5, 104515.1, 
    104774.7, 104539.6, 104125.1, 103766.9, 103441.2, 103082.7, 102741.3, 
    102336,
  104240.4, 104412.9, 104547.7, 104658.2, 104731.7, 104483.7, 100682.8, 
    103848.2, 103797.8, 103689.7, 103421.2, 103057.7, 102733.5, 102381.6, 
    101983,
  104118, 104283.1, 104402.5, 104473.1, 104504.9, 104468, 104165, 98033.19, 
    96979.96, 103012.9, 103080, 102665.9, 102357.1, 101955.7, 101603,
  103975.7, 104126.5, 104209, 104271.6, 104216.5, 104144.3, 103993.8, 
    103667.2, 103222, 103053.8, 102709.2, 102340.2, 101990.5, 101563, 101169.5,
  103829.4, 103960.7, 104019, 104034.9, 103974.7, 103835.2, 103613.4, 
    103375.5, 103046, 102655.7, 102357.3, 102013.9, 101607.4, 101178.5, 
    100739.3,
  103681.5, 103757.3, 103774.5, 103753.2, 103630.5, 103454.1, 103201.3, 
    102893.4, 102581.3, 102352.1, 102046.5, 101673.6, 101257.2, 100812, 
    100344.6,
  103525, 103566.2, 103541.2, 103459.1, 103313.1, 103089.8, 102821.3, 
    102557.5, 102324.4, 102050.7, 101698.1, 101322.1, 100898.1, 100427.6, 
    99936.55,
  103347.4, 103312.8, 103232.4, 103116.7, 102903, 102665.1, 102414.9, 
    102199.7, 101972.9, 101686.6, 101369.8, 100986.5, 100535.7, 100054, 
    99571.75,
  104041.6, 104119.7, 104253.2, 104374.4, 104544.2, 104667.7, 104731.2, 
    104805.5, 104797.7, 104374.5, 104297.7, 104402.6, 104056.8, 103409.9, 
    103061.4,
  103917.3, 103958.1, 104079.8, 104216.1, 104316.7, 104283.7, 104540.1, 
    104516, 104448.9, 104443, 104309.7, 104184.6, 104004.8, 101941.5, 102382.4,
  103727.1, 103793.9, 103892, 104040.5, 104047.3, 100616.5, 104021.7, 
    104413.4, 104292.1, 104156, 104023.4, 103898.9, 103762, 103626.8, 103426.5,
  103534.8, 103582, 103654.5, 103741.9, 103914.2, 103783.5, 100141.5, 
    103592.1, 103876.2, 103871.4, 103744.9, 103583.6, 103501.1, 103404.1, 
    103227.2,
  103305.7, 103359.6, 103419.4, 103496.6, 103582.1, 103742, 103611.7, 
    97680.62, 96705.26, 103208.5, 103475.2, 103299.7, 103243.4, 103110.5, 
    103009.7,
  103093.4, 103138.1, 103171.6, 103249.2, 103289.9, 103348.2, 103438.8, 
    103308.1, 103177.4, 103317.5, 103163.6, 103036, 102949.2, 102821.4, 
    102720.3,
  102873, 102907.7, 102931.3, 102988.9, 103045, 103078.3, 103081.2, 103113.5, 
    103027.4, 102863.1, 102771, 102674.8, 102572.7, 102458.2, 102347.2,
  102663, 102682.5, 102696.6, 102747.5, 102766.9, 102787.4, 102767.9, 
    102689.6, 102605.6, 102530.9, 102422.5, 102311.1, 102207.8, 102102.8, 
    102004.6,
  102475.7, 102494.2, 102493, 102512.6, 102532.6, 102531.5, 102487.7, 
    102434.2, 102319.4, 102169.8, 102044.9, 101939.2, 101841.2, 101742.2, 
    101634.5,
  102276.7, 102302.6, 102318.2, 102334, 102311.7, 102280.8, 102208, 102091.5, 
    101952.8, 101809.9, 101721.5, 101621.6, 101516.6, 101420.9, 101323,
  104208, 104081.4, 103992, 103864.2, 103761.3, 103648.1, 103532.9, 103477.5, 
    103459.1, 103099.4, 103132.4, 103379.6, 103189.4, 102694.2, 102430,
  104034.5, 103873.1, 103775.4, 103637.2, 103508.9, 103223.1, 103368.7, 
    103254, 103193.2, 103222.5, 103188.7, 103189.2, 103132.9, 101132.8, 
    101649.5,
  103808.1, 103662.9, 103539.2, 103413.7, 103186.4, 99686.29, 102951.9, 
    103232.5, 103128.6, 103039, 102962.8, 102939.6, 102873, 102793.5, 102657.6,
  103605, 103455.4, 103314.7, 103171.8, 103073.5, 102829.5, 99134.01, 
    102619.3, 102838.9, 102829.6, 102748.9, 102686.6, 102632.3, 102578.5, 
    102455.6,
  103398.1, 103265.5, 103125.2, 102982.5, 102885, 102816.1, 102647.4, 
    96715.71, 95903.22, 102382.5, 102591, 102502.3, 102484.5, 102417, 102369.4,
  103205.6, 103057.4, 102900.4, 102783.9, 102666.8, 102612, 102592.9, 
    102497.9, 102355.1, 102500.1, 102415, 102365, 102372.8, 102309.6, 102215.7,
  102984.2, 102848, 102697.7, 102599, 102519.5, 102471.5, 102421.6, 102413.5, 
    102362.8, 102279.2, 102263.7, 102296, 102267.9, 102186.8, 102034.4,
  102773.6, 102640.4, 102508.4, 102437.3, 102356.3, 102333.8, 102289.4, 
    102227.4, 102189, 102214.2, 102238.8, 102233.8, 102183.6, 102065.9, 
    101885.9,
  102556.8, 102460.5, 102365.6, 102313.4, 102272.5, 102245.1, 102190.7, 
    102169.6, 102145.9, 102150.7, 102162.4, 102160.8, 102079.8, 101940.6, 
    101714,
  102392, 102294.9, 102231.8, 102201.9, 102158.6, 102129.4, 102091.9, 
    102063.8, 102059.7, 102070.1, 102073.9, 102042.1, 101957.7, 101803, 
    101567.1,
  104790.1, 104682.9, 104582.4, 104407, 104220.9, 103977.5, 103679.3, 
    103460.7, 103260.9, 102705.9, 102632, 102767.9, 102547.2, 102056.3, 101872,
  104644.3, 104519.5, 104404.1, 104224.4, 104002.9, 103534.9, 103556.8, 
    103200.5, 102971.5, 102888.8, 102761.4, 102665.4, 102574.4, 100601.8, 
    101175,
  104486.2, 104379.2, 104235, 104075.9, 103697.2, 100118.2, 103092.1, 
    103259.2, 102993.1, 102767.7, 102603.5, 102526.5, 102415.2, 102333.4, 
    102214.8,
  104335.3, 104219.2, 104069.7, 103864.4, 103655.1, 103206.5, 99383.4, 
    102552.7, 102631.6, 102616.7, 102464.9, 102352.7, 102249.5, 102160.3, 
    102037,
  104166.8, 104064, 103906.3, 103697.3, 103494.4, 103257.9, 102888.7, 
    96832.9, 95940.96, 102172.1, 102320, 102161.3, 102075.9, 101951.9, 101871,
  104000.6, 103879.6, 103698.2, 103519.4, 103282.1, 103078.7, 102867.4, 
    102585.2, 102248.9, 102265.9, 102119.3, 101969.3, 101873.1, 101750.3, 
    101701.3,
  103807.5, 103702.9, 103532.4, 103350.2, 103144.5, 102905.9, 102674, 102479, 
    102276.2, 102044.6, 101897.5, 101764.3, 101648.6, 101578.9, 101540.7,
  103623.8, 103499, 103326.4, 103152.4, 102916.1, 102693.2, 102451.7, 
    102197.7, 101978.1, 101828.9, 101677.4, 101548.7, 101486.4, 101486.8, 
    101429.2,
  103417.1, 103312, 103145.4, 102950.1, 102722.1, 102473.3, 102199, 101985.4, 
    101779.3, 101586.1, 101437.7, 101414.8, 101438.3, 101414.3, 101345.9,
  103213.3, 103062.1, 102877.1, 102689.4, 102428.4, 102172.8, 101907.5, 
    101658.7, 101438.9, 101287.6, 101319.3, 101408.3, 101408.5, 101383.2, 
    101279.1,
  105038.2, 104918, 104844.2, 104735.6, 104643.8, 104481.5, 104268.9, 
    104099.4, 103872.2, 103258, 103033.8, 102996.7, 102566.2, 101821.2, 
    101381.6,
  104823.5, 104693.2, 104612.7, 104526.6, 104401.3, 104056, 104100.4, 
    103810.4, 103546.3, 103359.9, 103082, 102817.6, 102511.1, 100360.1, 
    100648.2,
  104555.3, 104442.3, 104350.8, 104294.1, 104065.1, 100551.4, 103593.9, 
    103812, 103512.3, 103176.9, 102865.5, 102586.9, 102264.4, 101951, 101571.7,
  104269, 104161.4, 104071, 103985.7, 103918, 103596.7, 99844.81, 102971.3, 
    103004.5, 102904.1, 102645.1, 102305.8, 101987.9, 101674.8, 101339,
  103913.7, 103846.4, 103772.1, 103707.3, 103640.3, 103550.6, 103257.1, 
    97256.7, 96249.91, 102313.6, 102382.4, 102002.5, 101692.6, 101352.2, 
    101145.5,
  103569.1, 103521.6, 103445.9, 103409.2, 103316.3, 103231.5, 103117, 102833, 
    102479.7, 102407.3, 102083.2, 101721.6, 101383.9, 101084.2, 100946.5,
  103215.6, 103191.9, 103137.3, 103099.1, 103033.1, 102921.6, 102773.3, 
    102632.6, 102386.9, 102063.3, 101748.3, 101408.5, 101073.2, 100868.2, 
    100794.6,
  102938.5, 102892, 102828.9, 102785.8, 102690.4, 102590.2, 102432, 102214.4, 
    101978.2, 101742.4, 101430.8, 101098.5, 100839, 100771.6, 100809.6,
  102639.2, 102589.1, 102525.3, 102457.5, 102366.5, 102243.4, 102075.3, 
    101909.6, 101694.7, 101408.5, 101108.3, 100830.5, 100706.8, 100813.4, 
    100894.9,
  102289.7, 102221.9, 102150.6, 102086.3, 101982.5, 101857.2, 101698.3, 
    101505, 101278.1, 101024.9, 100815.5, 100642.9, 100751.4, 100916.5, 
    100948.2,
  104547.3, 104416.7, 104313.3, 104158.8, 104057.5, 103912.2, 103728.7, 
    103567.2, 103391.4, 102844, 102688.1, 102716.9, 102323.4, 101613.2, 
    101178.5,
  104205.3, 104050, 103945.4, 103823, 103697.4, 103348.3, 103413.4, 103192.5, 
    102990.6, 102861.8, 102649.2, 102464.8, 102215.4, 100121, 100458.4,
  103787.6, 103638.3, 103521.2, 103434.5, 103209.6, 99692.86, 102745.9, 
    103056.5, 102794.4, 102589.3, 102364.7, 102177.4, 101949, 101714, 101410.4,
  103371, 103240.9, 103131.5, 103017.1, 102946.2, 102647.1, 98952.56, 
    102149.4, 102358.3, 102284.4, 102116.9, 101895.6, 101707.8, 101493.8, 
    101214.4,
  102909.1, 102818.7, 102727, 102637, 102573.3, 102496.6, 102238.8, 96350.95, 
    95403.64, 101682.9, 101858.4, 101618.9, 101452.2, 101217.8, 101026.6,
  102469.3, 102406.1, 102310.8, 102268.8, 102178.6, 102128.1, 102069.3, 
    101870.5, 101662.3, 101740.2, 101556.8, 101371.9, 101195, 100984.7, 
    100818.3,
  102034.3, 101999.4, 101922, 101884.2, 101833.1, 101773.7, 101695.3, 
    101666.8, 101542.8, 101374.2, 101248.6, 101092.6, 100906.7, 100727, 
    100625.4,
  101708.6, 101656.4, 101573.8, 101552.8, 101492.2, 101450.6, 101371.5, 
    101265.6, 101165.3, 101085.7, 100955.8, 100800.2, 100643.8, 100501.7, 
    100496,
  101322.3, 101273.3, 101210.9, 101167.7, 101109.9, 101056, 100989.9, 
    100948.4, 100861.6, 100741.4, 100622.1, 100498.4, 100364.7, 100295.2, 
    100334.7,
  100868.6, 100808.5, 100749.2, 100718.3, 100672.1, 100621.5, 100562.8, 
    100486.4, 100413.5, 100324.6, 100272, 100190.3, 100105.5, 100113.6, 
    100193.5,
  103042.5, 103053.4, 103082, 103050.8, 103048.7, 102997.7, 102904.7, 
    102854.4, 102760.3, 102283.3, 102199.4, 102314.3, 102023, 101433, 101108.6,
  102636.5, 102604.9, 102628.9, 102610.9, 102585, 102377.3, 102519.8, 
    102380.2, 102273.5, 102228.5, 102085.7, 102001.1, 101876.9, 99876.31, 
    100309.9,
  102141.9, 102097.3, 102091.2, 102116.4, 102022.4, 98623.49, 101715.9, 
    102137.7, 101938.1, 101827.1, 101707.2, 101635.7, 101527.8, 101413.6, 
    101238.2,
  101656.5, 101620.9, 101596.3, 101586.5, 101601, 101424.1, 97877.58, 
    101147.3, 101502.3, 101471.5, 101400.1, 101279.6, 101230.6, 101145.9, 
    101002.1,
  101154.7, 101129.7, 101108.1, 101107.7, 101123.5, 101157.8, 100998.3, 
    95304.26, 94399.48, 100781.7, 101079, 100950.2, 100940.5, 100849.8, 
    100785.2,
  100704.5, 100683.3, 100653.7, 100676.9, 100669.7, 100704.9, 100750.1, 
    100639.4, 100571.2, 100806.9, 100751.9, 100717, 100690.6, 100621.9, 
    100535.5,
  100299.4, 100277.5, 100236.3, 100241.9, 100260.3, 100286.2, 100314.7, 
    100417.9, 100432.7, 100405.8, 100435.2, 100432.9, 100390.8, 100330.7, 
    100242.2,
  100086.3, 100038.6, 99956.92, 99928.62, 99895.37, 99926.18, 99957.36, 
    99969.45, 100018, 100102.5, 100130.3, 100127, 100108.9, 100061.6, 99988.34,
  99938.02, 99880.28, 99779.02, 99687.3, 99609.95, 99593.2, 99613.74, 
    99696.15, 99747.19, 99772.75, 99800.59, 99816.73, 99801.08, 99768.27, 
    99703.13,
  99890.44, 99791.55, 99655.91, 99533.21, 99427.16, 99362.02, 99324.38, 
    99307, 99344.91, 99399.7, 99472.25, 99500.66, 99499.35, 99478.03, 99416.65,
  101673.6, 101727.5, 101822.6, 101897.7, 102023.1, 102111.8, 102174.5, 
    102250.6, 102306.5, 101979.1, 102005.3, 102217.4, 101994.9, 101463.6, 
    101178.6,
  101333.6, 101376.4, 101471.4, 101557.3, 101625.9, 101556.6, 101801.4, 
    101815.8, 101823.6, 101915.9, 101871.1, 101864.6, 101814.5, 99866.88, 
    100332,
  100918.8, 100965, 101067.7, 101181.1, 101193.2, 97880.38, 101121.4, 
    101582.1, 101487.9, 101467.3, 101467.5, 101446.7, 101407.9, 101331.7, 
    101250.4,
  100559.6, 100568.3, 100640.8, 100698.7, 100828.1, 100713.7, 97252.46, 
    100610.2, 101037.3, 101075.6, 101081.3, 101023.4, 101031.6, 101002, 100948,
  100287.9, 100259.9, 100273.7, 100330.9, 100395.5, 100547.7, 100459.6, 
    94837.89, 93887.41, 100333.9, 100678.4, 100594.3, 100625.8, 100584.8, 
    100598.7,
  100231.1, 100160.3, 100093.2, 100085.5, 100052.4, 100075.2, 100175.3, 
    100117.5, 100085.6, 100368.8, 100321.2, 100312.4, 100329.4, 100312, 
    100308.8,
  100239, 100189.9, 100139.2, 100112.9, 100097.2, 100047.4, 99992.48, 100032, 
    100001, 99951.93, 99997.41, 100008.4, 100002.9, 100000.8, 99999.3,
  100267.8, 100192.1, 100093.8, 100042.9, 99952.7, 99892.91, 99818.95, 
    99729.18, 99703.06, 99751.97, 99749.25, 99737.62, 99731.93, 99713.09, 
    99703.57,
  100352.9, 100268.9, 100153.3, 100067, 99975.84, 99872.03, 99769.07, 
    99722.77, 99637.95, 99547.96, 99498.28, 99481.88, 99474.38, 99464.84, 
    99452.64,
  100493, 100379.7, 100243.2, 100103.8, 99982.3, 99908.3, 99862.54, 99700.8, 
    99485.43, 99332.98, 99283.05, 99254.3, 99231.52, 99210.2, 99194.79,
  101316.2, 101332.2, 101402.6, 101461.9, 101575.5, 101668.6, 101741.6, 
    101846.1, 101942.9, 101671.2, 101777, 102095.9, 101970.8, 101575, 101389.4,
  100964.5, 100986.7, 101047.1, 101121.5, 101184.8, 101115.5, 101369.9, 
    101412.5, 101461.2, 101593.5, 101628.3, 101728.7, 101762.8, 99915.49, 
    100483.5,
  100584.7, 100582, 100642.2, 100744.1, 100763.2, 97410.82, 100730.4, 
    101135.9, 101106.5, 101157.4, 101208.4, 101290.8, 101346, 101372.2, 
    101373.9,
  100358.2, 100266.8, 100241.3, 100236.4, 100353.8, 100319.3, 96828.44, 
    100295, 100689.7, 100749.8, 100807, 100839.3, 100916.3, 100988.9, 101030.7,
  100332.5, 100271.3, 100197, 100122.9, 100067.8, 100159.9, 100135.6, 
    94429.14, 93602.18, 100081.4, 100429.3, 100407, 100498.5, 100521.5, 100623,
  100376.6, 100290.4, 100213.8, 100140.1, 100033.6, 99961.58, 100024.2, 
    99994.57, 99957.16, 100220.8, 100180.1, 100168.7, 100191, 100200.7, 
    100242.2,
  100432.8, 100344.7, 100268.5, 100213.4, 100158.6, 100076.5, 99983.57, 
    100004.5, 99962.62, 99937.65, 99971.01, 99986.65, 99979.44, 99965.39, 
    99959.83,
  100512.8, 100410.4, 100315, 100245.5, 100152.6, 100095.1, 100058.3, 
    99972.8, 99943.43, 99985.33, 99944.27, 99909.38, 99887.38, 99861.62, 
    99838.34,
  100561.5, 100492.6, 100411.7, 100337.9, 100279.2, 100190.4, 100107.8, 
    100072.1, 100005, 99919.47, 99808.41, 99753.93, 99700.98, 99644.05, 
    99587.47,
  100625.5, 100538.5, 100464.9, 100368.8, 100295.5, 100224.7, 100173.5, 
    100061.1, 99943.75, 99839.08, 99758.77, 99671.92, 99567.98, 99479.2, 
    99357.45,
  100915.6, 100923.8, 100975, 101030.8, 101132.8, 101209.3, 101268.2, 
    101368.1, 101477.9, 101267.4, 101434.6, 101826.8, 101774.8, 101466.7, 
    101396.3,
  100616.6, 100628.7, 100678.9, 100735.1, 100792.8, 100713.1, 100949.3, 
    101010.6, 101090.5, 101258, 101364.5, 101529.7, 101640.8, 99858.49, 
    100550.5,
  100289.4, 100242.6, 100300.8, 100385.1, 100441.1, 97098.8, 100451.8, 
    100798, 100799.4, 100894.8, 101004.5, 101144.2, 101278.4, 101382.3, 
    101472.8,
  100082.5, 99995.67, 99977.59, 99966.04, 100059.3, 100044.5, 96515.27, 
    100035.8, 100414.7, 100497.4, 100621.7, 100728.2, 100886.2, 101047.7, 
    101178.8,
  99942.47, 99887.98, 99876.62, 99901.03, 99892.57, 99956.05, 99921.38, 
    94155.7, 93399.55, 99887.39, 100236.5, 100290.4, 100443.9, 100558.5, 
    100746.9,
  99903.91, 99818.62, 99782.41, 99784.86, 99811.5, 99811.29, 99824.29, 
    99767.8, 99695.66, 99940.34, 99958.3, 100017.6, 100117.2, 100218.3, 
    100340.3,
  99937.19, 99855.11, 99811.44, 99839.55, 99840.59, 99824.21, 99800.5, 
    99802.73, 99760.1, 99733.15, 99771.97, 99818.07, 99873.89, 99943.55, 
    100036.8,
  100037.4, 99968.65, 99936.21, 99966.4, 99960.49, 99931.8, 99907.55, 
    99860.67, 99848.46, 99876.51, 99827.34, 99817.19, 99831, 99865.16, 
    99920.47,
  100224.2, 100172.3, 100148, 100182.5, 100198.8, 100155.4, 100084.1, 
    100024.8, 99944.21, 99852.65, 99732.6, 99728.7, 99730.59, 99773.15, 
    99818.82,
  100435.7, 100359.6, 100332, 100348.8, 100339.1, 100285.3, 100233.6, 
    100105.3, 99984.18, 99877.99, 99821.77, 99798.84, 99750.88, 99755.93, 
    99765.8,
  100117.6, 100122.7, 100181.6, 100260, 100385, 100494.3, 100569.8, 100692.3, 
    100828.3, 100631.2, 100806.5, 101211.1, 101185.3, 100928.1, 100921.3,
  99824.75, 99816.73, 99865.04, 99948.07, 100046.4, 99997.8, 100285.7, 
    100398.4, 100509, 100710.5, 100848.8, 101013.1, 101140.9, 99387.05, 
    100134.6,
  99559.73, 99496.7, 99516.67, 99592.94, 99693.49, 96378.05, 99766.23, 
    100200.5, 100295, 100433.8, 100585.4, 100750, 100913.1, 101036.3, 101176.2,
  99440.47, 99340.39, 99256.76, 99194.43, 99292.37, 99308.42, 95864.62, 
    99451.1, 99922.48, 100110.4, 100304, 100451.4, 100646.3, 100837.6, 
    101002.6,
  99421.53, 99398.3, 99318.59, 99212.66, 99112.43, 99211.14, 99216.92, 
    93577.45, 92899.3, 99449.48, 99951.57, 100083.2, 100334.3, 100482.9, 
    100735.5,
  99405.72, 99445.21, 99424.95, 99375.47, 99242.83, 99153.66, 99209.08, 
    99168.94, 99144.98, 99475.85, 99605.36, 99774.87, 99982.93, 100193.3, 
    100400.4,
  99405.03, 99534.53, 99556.3, 99543.16, 99514.91, 99455.35, 99366.67, 
    99362.95, 99385.29, 99341.51, 99404, 99551.84, 99716.24, 99896.93, 
    100070.9,
  99421.76, 99565.48, 99608.66, 99647.85, 99627.12, 99640.09, 99639.86, 
    99601.91, 99576.12, 99562.22, 99464.41, 99487.42, 99578.19, 99712.8, 
    99855.62,
  99406.21, 99587.59, 99653.95, 99708.78, 99733.76, 99752.28, 99719.34, 
    99719.31, 99689.91, 99647.73, 99570.91, 99611.95, 99606.96, 99662.94, 
    99733.22,
  99414, 99614.88, 99715.84, 99764.52, 99772.42, 99822.92, 99818.05, 
    99763.34, 99703.39, 99676.3, 99685.51, 99731.07, 99730.84, 99740.66, 
    99735.35,
  99140.16, 99258.92, 99400.43, 99517.55, 99653.15, 99799.41, 99902.68, 
    100033, 100157, 99948.17, 100105.7, 100478.1, 100420.6, 100140.4, 100091.2,
  98839, 98971.55, 99144.13, 99270.8, 99387.91, 99362.08, 99638.42, 99737.5, 
    99856.75, 100037.7, 100145.5, 100293.9, 100384.8, 98634.61, 99368.34,
  98502.59, 98706.02, 98896.62, 99029.02, 99052.38, 95797.71, 99162.05, 
    99525.59, 99598.21, 99754.11, 99890.62, 100040.4, 100181.9, 100294.5, 
    100408,
  98280.23, 98513.98, 98748.35, 98856.17, 98938.39, 98847.36, 95367.04, 
    98912.1, 99330.38, 99485.73, 99663.94, 99791.15, 99969.47, 100147.3, 
    100313.8,
  98223.2, 98542.23, 98790.73, 98895.9, 98859.04, 98876.87, 98814.09, 
    93100.03, 92438.28, 98966.41, 99395.77, 99519.78, 99734.75, 99871, 
    100119.1,
  98286.48, 98591.77, 98812.75, 98918.11, 98903.52, 98839.98, 98935.91, 
    98943.73, 98961.98, 99207.24, 99200.34, 99299.66, 99490.33, 99683.46, 
    99913.25,
  98290.13, 98602.19, 98862.9, 98987.26, 99059.05, 99074.25, 99118.51, 
    99301.51, 99355.87, 99299.2, 99224.52, 99199.38, 99283.31, 99462.86, 
    99691.62,
  98418.55, 98703, 98889.66, 98941.03, 98938.83, 99024.76, 99152.48, 
    99248.49, 99338.98, 99356.62, 99289.16, 99168.33, 99148.1, 99293.99, 
    99527.42,
  98689.48, 98943.94, 99031.58, 99049.51, 99025.66, 99089.99, 99205, 
    99343.33, 99430.13, 99410.02, 99322.21, 99210.65, 99048.25, 99132.09, 
    99353.91,
  99211.08, 99266.25, 99308.41, 99326.1, 99367.47, 99423.73, 99441.12, 
    99426.95, 99415.49, 99422.8, 99388.54, 99290.39, 99047.05, 99033.08, 
    99241.77,
  98101.26, 98221.14, 98433.01, 98684.23, 99000, 99314.68, 99562.99, 
    99813.76, 100027.8, 99884.82, 100094.9, 100499.5, 100464.6, 100144.9, 
    100054.7,
  97946.26, 98050.83, 98258.2, 98512.23, 98779.84, 98956.1, 99370.89, 
    99595.97, 99797.52, 100040.9, 100202, 100388.4, 100524.1, 98750.98, 
    99496.78,
  97710.31, 97879.75, 98124.34, 98404.59, 98566.02, 95485.41, 99022.2, 
    99501.42, 99668.62, 99851.35, 100020.4, 100194.6, 100381.8, 100516.6, 
    100632.5,
  97570.8, 97733.26, 98029.45, 98312.84, 98637.93, 98607.38, 95265.9, 
    98945.52, 99434.28, 99653.52, 99846.42, 99993.5, 100200.7, 100384.9, 
    100559.4,
  97455.85, 97746.02, 98055.7, 98329.27, 98598.7, 98843.59, 98788.8, 
    93125.64, 92539.81, 99125.52, 99629.25, 99762.27, 99998.58, 100145.1, 
    100372.4,
  97648.48, 97934.74, 98206.02, 98430.12, 98583.28, 98678.62, 98848.72, 
    98858.69, 98857.52, 99257.12, 99408.02, 99563.93, 99766.31, 99944.17, 
    100139.6,
  97846.49, 98112.55, 98374.34, 98561.78, 98698.02, 98732.14, 98708.56, 
    98843.19, 99047.41, 99175.23, 99349.31, 99506.91, 99627.08, 99756.44, 
    99909.73,
  98094.65, 98399.59, 98672.92, 98825.04, 98855.18, 98787.68, 98660.35, 
    98612.72, 98836.16, 99132.36, 99359.03, 99519.65, 99653.44, 99732.12, 
    99794.69,
  98650.11, 98875.78, 99033.85, 99111.61, 99097.31, 98938.29, 98565.44, 
    98517.48, 98763.77, 99057.08, 99320.45, 99513.88, 99647.7, 99723.06, 
    99754.53,
  99137.2, 99246.46, 99334.84, 99387.7, 99325.48, 99218.13, 99009.54, 
    98792.59, 98891.2, 99096.59, 99365.91, 99533.75, 99626.97, 99677.12, 
    99682.4,
  98336.3, 98348.3, 98407.49, 98499.08, 98671.57, 98878.44, 99112.63, 
    99399.73, 99690.29, 99635.85, 99938.94, 100405.1, 100387.4, 100033.2, 
    99852,
  98238.12, 98255.85, 98290.65, 98393.51, 98509.89, 98584.52, 98962.91, 
    99215.45, 99497.91, 99835.14, 100081.6, 100312.9, 100464.9, 98632.11, 
    99282.18,
  98132, 98171.28, 98228.23, 98339.93, 98359.24, 95221.07, 98708.41, 
    99193.94, 99430.01, 99715.59, 99964.35, 100203.5, 100394.2, 100480.4, 
    100489.4,
  98034.77, 98033.23, 98131.67, 98258.98, 98463.8, 98370.57, 95068.89, 
    98792.57, 99350.23, 99638.42, 99889.07, 100078, 100305.1, 100452.4, 
    100502.9,
  98083.34, 98164.65, 98236.3, 98360.32, 98498.73, 98711.7, 98632.26, 
    93080.68, 92571.27, 99272.44, 99813.26, 99970.3, 100205.5, 100336.6, 
    100488.9,
  98356.77, 98408.09, 98465.42, 98550.02, 98611.76, 98721.47, 98898.91, 
    98935.96, 98934.55, 99429.55, 99645.64, 99860.66, 100089.5, 100266.5, 
    100424.9,
  98652.3, 98723.36, 98770.08, 98837.92, 98902.18, 98949.9, 98962.2, 
    99085.91, 99189.16, 99282.05, 99500.6, 99732.16, 99954.39, 100163.1, 
    100343.2,
  99045.41, 99135.89, 99158.77, 99233.16, 99235.87, 99268.09, 99263.94, 
    99173.3, 99096.84, 99157.92, 99348.12, 99582.14, 99828.54, 100059.1, 
    100272.8,
  99354.65, 99421.73, 99455.29, 99511.05, 99537.49, 99516.33, 99426.48, 
    99384.54, 99282.83, 99169.56, 99197.63, 99426.07, 99686.48, 99952.26, 
    100189.1,
  99624.33, 99661.8, 99699.62, 99743.95, 99704, 99662.34, 99554.55, 99353.48, 
    99131.76, 98983.07, 99077.73, 99293.38, 99578.19, 99881.95, 100146.4,
  98904.36, 98960.69, 99047.53, 99150.88, 99295.38, 99429.59, 99607.53, 
    99834.73, 100074.2, 99975.79, 100274.3, 100805.2, 100906.2, 100745.2, 
    100799,
  98806.1, 98844.84, 98894.3, 99014.02, 99108.63, 99143.87, 99448.37, 99614, 
    99828.24, 100117.5, 100347.1, 100652, 100898.8, 99289.39, 100127.4,
  98614.44, 98686.41, 98797.05, 98905.05, 98890.7, 95673.4, 99137.68, 
    99560.98, 99720.05, 99951.78, 100176.8, 100463.2, 100760.8, 100995.2, 
    101223.9,
  98587.76, 98538.23, 98549.3, 98657.61, 98902.31, 98759.52, 95393.23, 
    98987.69, 99491.33, 99759.08, 100038.9, 100288.4, 100627.5, 100943.6, 
    101201.2,
  98768.05, 98690.55, 98589.06, 98576.03, 98665.54, 98926.63, 98821.27, 
    93245.96, 92720, 99327.5, 99909.23, 100147.6, 100510.9, 100787.1, 101121.5,
  99054.7, 98986.53, 98863.17, 98725.81, 98659.41, 98740.66, 98919.13, 
    98911.55, 98902.78, 99454.18, 99733.54, 100046.6, 100412.8, 100737, 
    101063.6,
  99264.55, 99260.21, 99242.4, 99193.18, 99091.46, 99008.61, 98939.04, 
    99085.42, 99234.92, 99346.1, 99620.41, 99970.66, 100333, 100679.2, 
    101007.1,
  99481.54, 99477.45, 99496.17, 99493.7, 99448.23, 99430.25, 99356.98, 
    99133.65, 99121.39, 99314.95, 99597.29, 99928.36, 100303, 100659.7, 
    101000.7,
  99593.98, 99649.45, 99713.05, 99773.45, 99783.3, 99720.93, 99651.23, 
    99620.27, 99484.56, 99451.45, 99616.48, 99932.47, 100295.2, 100659.4, 
    100998.1,
  99722.96, 99846.13, 99906.32, 99997.02, 99983.27, 99965.95, 99873.24, 
    99714.52, 99600.67, 99562.23, 99703.3, 99982.03, 100317.9, 100679.3, 
    101003,
  99058.35, 99042.12, 99069.75, 99019.22, 98965.16, 98915.14, 98888.56, 
    98935.34, 99067.8, 98938.67, 99266.91, 99841.95, 99992.37, 99931.21, 
    100126.9,
  99019.67, 99004.35, 99062.71, 99057.92, 99003.48, 98798.3, 98985.91, 
    98969.73, 99084.22, 99343.62, 99614.63, 99958.72, 100231.3, 98729.44, 
    99722.58,
  99009.18, 98905.74, 99056.52, 99076.8, 98961.95, 95574.34, 98948.84, 
    99188.85, 99320.08, 99485.03, 99734.05, 100054.6, 100393.7, 100679.4, 
    101022.2,
  99132.27, 98879.82, 98912.5, 99033.59, 99166.53, 98900.03, 95427.08, 
    99005.26, 99358.66, 99597.23, 99875.85, 100161.6, 100528, 100909.7, 
    101226.3,
  99409.54, 99141.91, 98919.11, 98942.54, 99114.56, 99266.9, 99106.57, 
    93332.97, 92899.09, 99532.78, 100028.8, 100280.1, 100643.2, 100950.6, 
    101340.1,
  99547.69, 99446.13, 99188.61, 99012.16, 99065.25, 99198.09, 99405.39, 
    99391.25, 99328.23, 99854.6, 100098.6, 100399.6, 100743.9, 101087.5, 
    101427.3,
  99673.48, 99650.55, 99582.26, 99356.11, 99214.17, 99296.23, 99366.2, 
    99610.17, 99828.82, 99948, 100180.5, 100496.5, 100807.7, 101143.7, 
    101465.2,
  99797.26, 99839.59, 99826.68, 99778.8, 99574.7, 99511.01, 99536.95, 
    99556.77, 99705.38, 99976.16, 100255.6, 100556.6, 100872.2, 101203.8, 
    101534.4,
  100007.3, 100036.8, 100069.6, 100080, 100021, 99904.1, 99834.07, 99857.79, 
    99900.12, 100063.3, 100296.8, 100593.4, 100899.8, 101227.1, 101563.8,
  100310.5, 100309.2, 100316.4, 100336.9, 100261.8, 100189.7, 100068.9, 
    99937.23, 99882.05, 100006, 100293.7, 100600.1, 100915.4, 101263, 101611.7,
  99252.1, 99067.85, 98953.34, 98817.25, 98704.61, 98670, 98652.6, 98749.96, 
    98959.76, 98877.42, 99183.61, 99712.84, 99823.09, 99670.59, 99735.35,
  99267.94, 99001.43, 98835.7, 98679.13, 98546.3, 98311.01, 98530.55, 
    98569.75, 98759.93, 99060.76, 99356.88, 99661.55, 99922.77, 98304.35, 
    99178.19,
  99305.24, 98994.62, 98797.4, 98657.63, 98447.84, 95041.2, 98380.09, 
    98637.55, 98885.59, 99085.61, 99349.49, 99631.1, 99933.84, 100154.3, 
    100366.8,
  99445.8, 99054.94, 98799.61, 98662.23, 98675.85, 98391.03, 94888.93, 
    98546.69, 98879.8, 99134.11, 99425.05, 99659.73, 99962.91, 100227.9, 
    100459.6,
  99565.75, 99244.1, 98947.47, 98761.41, 98744.39, 98827.23, 98644.2, 
    92785.29, 92435.61, 99068.97, 99559.91, 99739.28, 100044, 100230.8, 
    100548.3,
  99745.12, 99428.23, 99123.15, 98904.57, 98832.35, 98848.27, 99027.29, 
    99000.85, 98922.84, 99402.95, 99628.63, 99870.16, 100143.9, 100387.8, 
    100661.7,
  99939.64, 99720.56, 99415.71, 99167.12, 99013.97, 99024.25, 99036.23, 
    99251.37, 99430.84, 99548.9, 99764.96, 100034.2, 100280.5, 100557, 
    100842.8,
  100161.7, 99997.92, 99752.89, 99515.23, 99288.37, 99224.95, 99285.3, 
    99336.79, 99481.78, 99709.19, 99971.11, 100225.4, 100518.1, 100840.9, 
    101159.1,
  100441.4, 100320.3, 100128.5, 99953.58, 99737.26, 99592.5, 99561.66, 
    99690.23, 99839.49, 100006.6, 100224.8, 100500.3, 100819.6, 101126.3, 
    101409.2,
  100745.5, 100654.9, 100493.3, 100308.9, 100101.5, 99965.16, 99907.55, 
    99933.3, 100061.2, 100224.5, 100509.5, 100803.2, 101097, 101397.1, 
    101646.4,
  98851.69, 98643.27, 98503.3, 98453.24, 98443.98, 98479.84, 98798.52, 
    99252.91, 99623.51, 99569.07, 99844.84, 100312.4, 100366.3, 100179.4, 
    100235.8,
  98771.82, 98607.28, 98535.14, 98506.91, 98433.57, 98214.27, 98697.99, 
    99172.9, 99529.38, 99879.66, 100138.8, 100398.7, 100612.3, 98944.84, 
    99801.14,
  98776.97, 98580.34, 98552.09, 98518.98, 98338.75, 94967.66, 98622.41, 
    99238.37, 99650.37, 99934.87, 100198.1, 100454.2, 100706.9, 100903.1, 
    101070.8,
  98881.63, 98661.59, 98604.88, 98577.9, 98634.93, 98402.59, 95174.41, 
    99107.48, 99671.02, 99995.02, 100285, 100514.8, 100773.8, 100990.4, 
    101180.3,
  99051.32, 98869.22, 98779.23, 98798.43, 98846.95, 99045.26, 98970.66, 
    93397.38, 93085.69, 99913.84, 100399.6, 100590.4, 100829.4, 100979.9, 
    101207.6,
  99305.15, 99120.66, 99023.05, 99045.63, 99095.98, 99254.56, 99531.44, 
    99623.39, 99686.81, 100242.3, 100468.2, 100688.2, 100881.3, 101048.9, 
    101214.4,
  99585.27, 99433.81, 99323.39, 99332.55, 99415.38, 99547.89, 99713.62, 
    100005.1, 100232.7, 100374.5, 100574.2, 100774.7, 100924.5, 101072.8, 
    101192.2,
  99925.88, 99774.27, 99647.7, 99618.8, 99648.36, 99793.48, 99950.13, 
    100115.3, 100293.8, 100509, 100703.6, 100848.4, 100983.4, 101107.1, 
    101257.4,
  100306.8, 100160.9, 100052.4, 100031.5, 100030.2, 100101.2, 100229.1, 
    100430.3, 100589.5, 100706.9, 100820.2, 100937.5, 101068, 101220.7, 
    101360.2,
  100684.9, 100547.2, 100433.3, 100381.3, 100351.1, 100407.1, 100486.7, 
    100576.9, 100694.7, 100793.2, 100947.3, 101090, 101237, 101394.8, 101515.8,
  99336.01, 99292.65, 99296.56, 99389.95, 99619.47, 99811.76, 99934.55, 
    100042.2, 100181.8, 99947.05, 100023.1, 100290.6, 100169.8, 99835.93, 
    99743.12,
  99458.22, 99420.68, 99428.64, 99504.98, 99626.46, 99600.8, 99932.94, 
    100104.3, 100184.8, 100249.3, 100229.3, 100238.8, 100295.2, 98582.34, 
    99342.48,
  99631.01, 99583.61, 99607.52, 99670.19, 99635.55, 96419.27, 100020.6, 
    100315.7, 100389, 100354.6, 100290.6, 100233.4, 100309.6, 100475.9, 
    100629.9,
  99919.18, 99852.1, 99876.59, 99938.98, 100097.1, 99939.31, 96506.38, 
    100253.3, 100489.9, 100494.8, 100430.2, 100310.1, 100362.6, 100583.8, 
    100796.5,
  100213.8, 100179.8, 100187.5, 100247.1, 100382.2, 100504.1, 100384.5, 
    94369.85, 93829.8, 100469, 100612.5, 100466.2, 100491.5, 100631.1, 
    100945.2,
  100450.8, 100410.6, 100423.7, 100463.7, 100533.7, 100637, 100766.3, 100739, 
    100625.4, 100835.9, 100796.8, 100708.6, 100709, 100862.5, 101114.2,
  100616.1, 100610.1, 100609.5, 100652, 100700.1, 100780.5, 100848, 100969.3, 
    101027, 101026.5, 101012.8, 100986.1, 100982.6, 101106.3, 101298.1,
  100765.4, 100770.1, 100751.4, 100781.9, 100804.4, 100894.7, 100982, 101075, 
    101137.2, 101204.5, 101238.2, 101256, 101292.1, 101397.6, 101546,
  100924.9, 100958, 100985, 101034.4, 101066, 101088.6, 101148, 101245.6, 
    101307.8, 101349.3, 101391.9, 101441.6, 101498.1, 101588.8, 101701.5,
  101127.3, 101143.1, 101179.6, 101236.2, 101235, 101262.6, 101289.9, 
    101316.5, 101351.6, 101373.2, 101466.9, 101546.8, 101622.8, 101726.1, 
    101818.8,
  100789.3, 100827.7, 100912.1, 100974.2, 101044.3, 101048.8, 100982.9, 
    100888.4, 100726.4, 100191.8, 100011.4, 100009.5, 99700.41, 99289.42, 
    99264.91,
  100951.6, 100965.4, 101030.7, 101089.4, 101128.5, 100956.7, 101104.8, 
    101015.2, 100856.6, 100704.9, 100494.7, 100314.3, 100114.4, 98233.87, 
    98975.14,
  101067.9, 101088.5, 101154, 101199.8, 101089, 97630.54, 101134.8, 101249.4, 
    101122.6, 100922.9, 100718.2, 100558.6, 100440.9, 100384.2, 100345.5,
  101138.7, 101156.4, 101222.3, 101279, 101354.2, 101116.4, 97403.62, 
    101060.3, 101120.9, 101078.9, 100911.8, 100745.4, 100652.6, 100638.9, 
    100634,
  101275.1, 101317.5, 101348.6, 101409.2, 101463.5, 101479.1, 101286.5, 
    95073.16, 94393.1, 100972, 101062.9, 100866.8, 100830.9, 100780, 100845.4,
  101336, 101369.5, 101396.1, 101441.6, 101475.7, 101529.9, 101576.5, 
    101488.6, 101255.2, 101305.2, 101137.9, 100960.6, 100909.9, 100950.2, 
    101003.5,
  101336.7, 101390.8, 101420.4, 101473, 101511.4, 101581.8, 101616.2, 
    101684.4, 101636.5, 101475.4, 101254, 101064.3, 100968, 101060.8, 101143.8,
  101332, 101388.8, 101401.1, 101452.3, 101489.5, 101604.8, 101683.6, 
    101735.5, 101704.2, 101618.1, 101438.9, 101228.6, 101126, 101205.6, 101312,
  101381.3, 101467.9, 101520.1, 101589.2, 101643.8, 101683.8, 101750, 
    101835.1, 101839.5, 101756.6, 101624, 101460.9, 101343.2, 101368.9, 
    101447.3,
  101476.1, 101547.3, 101600.6, 101674.8, 101688, 101709.6, 101763.6, 
    101795.4, 101815.4, 101781.4, 101747.8, 101650.5, 101545.1, 101540.6, 
    101574,
  101692.4, 101622.3, 101560.3, 101415.2, 101292.6, 101126.6, 100878.2, 
    100655.3, 100380.2, 99715.3, 99530.26, 99836.68, 99988.98, 99973.04, 
    100130,
  101668.4, 101629.4, 101564.8, 101448.5, 101304.9, 100902.2, 100948, 100586, 
    100222.3, 99902.46, 99599.38, 99665.44, 99997.99, 98547.39, 99573.86,
  101586.2, 101603.4, 101576.2, 101500.8, 101193.9, 97576.3, 100754.6, 
    100826, 100453.1, 99988.45, 99605.89, 99633.83, 99995.41, 100392.2, 
    100765.5,
  101484.7, 101476.4, 101501.4, 101471.4, 101438.5, 100979.1, 97142.5, 
    100392.3, 100262.4, 100136.4, 99827.66, 99809.62, 100128.7, 100546.5, 
    100914.1,
  101397.5, 101441.1, 101480.1, 101446.1, 101459.3, 101350.8, 101021.4, 
    94670.55, 93879.62, 100172, 100171.6, 100088.2, 100344.9, 100597.7, 
    101014.7,
  101216.6, 101280, 101339.9, 101389.4, 101388.1, 101390.4, 101365.1, 
    101112.9, 100723.3, 100654.1, 100480.7, 100419.5, 100583.2, 100799.4, 
    101108.4,
  100989.6, 101075.2, 101142.5, 101239.8, 101334.5, 101405, 101396.9, 101393, 
    101240.8, 100985, 100776.8, 100750.9, 100817, 100977.7, 101187.6,
  100816.3, 100901.7, 100958.2, 101093, 101189.3, 101377, 101491.5, 101465.9, 
    101354.4, 101242.5, 101118.2, 101043.7, 101088.9, 101202.7, 101357.9,
  100678.4, 100804.6, 100898.8, 101068, 101216.7, 101398.7, 101532, 101638.6, 
    101614.4, 101508.5, 101394.4, 101324.3, 101321.7, 101377.4, 101463.1,
  100524.5, 100674.9, 100819.8, 101023.4, 101190.4, 101359.7, 101526.8, 
    101632.8, 101660.1, 101631.5, 101617, 101557.2, 101521, 101552.6, 101583.5,
  101030.3, 101046.8, 101039.3, 100944.1, 100860, 100734.8, 100549.2, 
    100454.4, 100452.1, 100175.8, 100365.8, 100766.6, 100692.1, 100379.1, 
    100347.2,
  100791.8, 100836.3, 100834, 100747, 100637.8, 100262.1, 100368.2, 100196.4, 
    100136.1, 100277.9, 100459.7, 100712.1, 100858.7, 99123.54, 99916.79,
  100486.9, 100593.2, 100604.1, 100559.4, 100268.6, 96729.73, 99872.95, 
    100124.8, 100059.6, 100152.9, 100335.5, 100622.5, 100884.3, 101051, 
    101200.7,
  100273.5, 100364.6, 100353.5, 100246.5, 100130.4, 99770.25, 96153.69, 
    99669.45, 99936.67, 99999.3, 100250, 100565.2, 100910.8, 101177.6, 
    101357.2,
  100154.7, 100246.8, 100227.1, 100095.9, 100042.6, 100059.1, 99887.91, 
    93793.68, 93144.84, 99813.32, 100279.3, 100606.1, 100977.5, 101203.5, 
    101471.6,
  100087.6, 100177.5, 100147.7, 100088.5, 100037, 100120.3, 100093.8, 
    99983.32, 99796.66, 100117.8, 100391.6, 100758.9, 101097.4, 101360.6, 
    101590.9,
  100090, 100218.1, 100198.7, 100169.1, 100168.2, 100205.4, 100150.7, 
    100195.2, 100238, 100355.9, 100621.8, 100967.8, 101254.2, 101509.7, 
    101728.6,
  100182.3, 100306.7, 100317.6, 100358.1, 100385, 100416.3, 100396.6, 100393, 
    100459.3, 100655.4, 100921, 101205.2, 101463.7, 101705.2, 101921.4,
  100325.3, 100458.4, 100553.6, 100670.6, 100740, 100758.7, 100750.1, 
    100795.3, 100873.1, 101019.9, 101222.8, 101456.9, 101671.1, 101884.4, 
    102067.9,
  100536.2, 100689.4, 100853.4, 100982.6, 101035.5, 101076.3, 101083.2, 
    101101.4, 101175.9, 101291.1, 101497.2, 101690.1, 101870.9, 102054, 
    102185.7,
  99915.42, 100124.5, 100392, 100658.6, 100923.1, 101114.9, 101225.3, 
    101290.3, 101342, 101009.5, 101070.9, 101320.6, 101120.2, 100664.9, 
    100510.6,
  99721.41, 99866.35, 100094.5, 100371.6, 100629.1, 100664.2, 100958.8, 
    101010.6, 101023.2, 101055.9, 101095, 101156.2, 101111.1, 99194.38, 
    99867.02,
  99650.04, 99797.12, 99956.51, 100206.2, 100336, 97073.24, 100572.6, 
    100846.6, 100848.7, 100883.1, 100955, 101050.7, 101044.6, 101052.5, 
    101039.3,
  99676.22, 99772.95, 99877.41, 100039.3, 100270.8, 100163.5, 96638.78, 
    100361.9, 100711.3, 100846.4, 100996.9, 101037.7, 101048.1, 101064, 
    101081.9,
  99616.69, 99667.34, 99755.04, 99900.45, 100230.6, 100430.6, 100307.4, 
    94473.02, 93943.81, 100779, 101093, 101078.1, 101096.6, 101068.7, 101119.3,
  99738.12, 99765.87, 99832.98, 99962.8, 100186.4, 100369.1, 100531.3, 
    100596.3, 100674.5, 101079.7, 101158.3, 101183.3, 101182.1, 101178.9, 
    101183.7,
  99959.25, 99975.96, 100014.8, 100149.1, 100312.4, 100494.9, 100686.1, 
    100972.1, 101156.1, 101241.7, 101313.5, 101358.6, 101356.5, 101365.5, 
    101352.6,
  100273.6, 100294.3, 100319.9, 100410.8, 100525.4, 100733.4, 100942.6, 
    101137.2, 101302.5, 101453.5, 101524.8, 101549.8, 101546.8, 101532.9, 
    101514.7,
  100684.5, 100727.8, 100777, 100884.4, 101006.8, 101155.7, 101324.7, 
    101511.3, 101634.8, 101701.9, 101739.6, 101748.3, 101730.7, 101696.7, 
    101655.5,
  101193.2, 101235.3, 101311.1, 101378.9, 101435.6, 101545.8, 101650.7, 
    101736.6, 101822.2, 101866.2, 101935.2, 101944.2, 101912.1, 101870.2, 
    101804.8,
  99852, 99972.51, 100176.5, 100467.2, 100835.3, 101183.7, 101456.2, 
    101701.5, 101899.5, 101689.6, 101820.8, 102116.7, 101969.9, 101524.5, 
    101343.6,
  99781.43, 99837.91, 100003.8, 100306.9, 100656.9, 100873.9, 101348.2, 
    101587, 101734.1, 101903.1, 101950.9, 101989.5, 101947.5, 99980.57, 
    100584.8,
  99643.7, 99783.04, 99916.09, 100226.2, 100440.3, 97362.97, 101064.8, 
    101573.6, 101700.5, 101786.8, 101806.7, 101807.5, 101750.7, 101675.9, 
    101579.8,
  99644.51, 99671.79, 99863.13, 100155, 100566.5, 100559.5, 97279.59, 
    101139.5, 101568.2, 101656.1, 101671.8, 101623.5, 101575.9, 101505.5, 
    101418,
  99712.09, 99780.61, 99941.07, 100247.2, 100622.5, 100951.5, 100917.1, 
    95154.13, 94513.38, 101279.1, 101578.7, 101510.7, 101476.1, 101394.7, 
    101357,
  99936.27, 100021.7, 100166.3, 100432.8, 100688.2, 100934.3, 101190.6, 
    101198.1, 101197.3, 101499.1, 101499.9, 101476.2, 101421.4, 101341, 
    101282.7,
  100169.8, 100285.8, 100418, 100611.8, 100808.3, 101009.8, 101208.1, 
    101435.7, 101525.8, 101506.3, 101514.1, 101465.5, 101397.2, 101338.7, 
    101278.3,
  100417.3, 100532.5, 100624.9, 100788, 100938.3, 101161.1, 101344.4, 
    101481.1, 101561.6, 101625.1, 101570, 101494.9, 101420.1, 101357.6, 
    101306.4,
  100712.8, 100827.1, 100929.4, 101089, 101242, 101409.9, 101552.5, 101684.7, 
    101720.1, 101690.5, 101640.3, 101568.6, 101487, 101420.3, 101362,
  101136.7, 101231.2, 101344.3, 101448.7, 101518.5, 101626.2, 101692.1, 
    101726, 101751.8, 101730.2, 101727.9, 101665.3, 101580.2, 101509.9, 
    101444.7,
  99924.36, 99973.17, 100032.8, 100125.6, 100301.2, 100544.8, 100800.8, 
    101084, 101405.7, 101291.2, 101506.7, 101818.1, 101652.2, 101118.5, 
    100853.9,
  99818.73, 99883.5, 99964.41, 100100.8, 100306.1, 100401.8, 100834.3, 
    101122.7, 101369.1, 101605.9, 101723.5, 101776.9, 101724.9, 99698.72, 
    100243.7,
  99688.64, 99877.88, 99977.02, 100174.3, 100234.7, 97087.33, 100825.4, 
    101294.6, 101474, 101582.8, 101647, 101673.6, 101625.4, 101526.7, 101373.4,
  99659.52, 99856.63, 100004.9, 100214, 100501.1, 100424.7, 97133.67, 
    101011.4, 101428.7, 101543.5, 101598.3, 101560.3, 101520.2, 101412.4, 
    101287.2,
  99758.68, 99923.77, 100080.4, 100322, 100612.1, 100899.5, 100816.5, 
    95031.75, 94398.46, 101170.6, 101486.4, 101444.3, 101409.6, 101327.2, 
    101289.5,
  99917.11, 100050.2, 100201, 100449.7, 100675, 100885.2, 101127.7, 101127, 
    101096.1, 101391.2, 101416.3, 101420.8, 101386.5, 101325.6, 101267.9,
  100123.4, 100255.2, 100393, 100588.9, 100780.5, 100952, 101112.9, 101318.6, 
    101434.5, 101431.7, 101457.7, 101431.9, 101375.4, 101334.6, 101285.6,
  100362.2, 100457.9, 100546.1, 100684.8, 100808.9, 100983.9, 101161.8, 
    101305.1, 101410.9, 101503.4, 101494.2, 101461, 101416.4, 101375.4, 
    101337.6,
  100584.2, 100664.6, 100727.6, 100841.5, 100954.4, 101102.1, 101260, 
    101433.3, 101528.8, 101550.1, 101551.5, 101523.4, 101475.3, 101437.5, 
    101402,
  100918.4, 100954.3, 101010.1, 101078.4, 101136.2, 101236.4, 101341.6, 
    101426.6, 101500.6, 101531.1, 101593.9, 101590.7, 101556.2, 101525.6, 
    101492.7,
  100423.6, 100451.9, 100480.5, 100501, 100532.4, 100542.7, 100492.2, 
    100481.8, 100549.7, 100342.8, 100593.7, 101063, 101094.9, 100826.4, 
    100744.3,
  100395.3, 100405.2, 100407.4, 100456.3, 100520.1, 100414.6, 100560.2, 
    100567.2, 100644, 100842.4, 101040.2, 101259.8, 101371, 99505.62, 100192.8,
  100327.6, 100418, 100476.7, 100551.8, 100482.2, 97115.67, 100625.7, 
    100872.4, 100996.7, 101103.2, 101255, 101387.8, 101471.8, 101474.5, 
    101377.6,
  100336.1, 100399.7, 100500.9, 100594.5, 100760.9, 100546.5, 97062.64, 
    100835.4, 101157.8, 101308.4, 101418.8, 101456.2, 101488, 101450.7, 
    101354.9,
  100448.4, 100514.6, 100596.3, 100726.4, 100868.5, 101035.5, 100871.7, 
    94927.38, 94398.14, 101222.2, 101530.2, 101492.5, 101516.3, 101468.2, 
    101435,
  100562.1, 100630.9, 100711.9, 100858.8, 100975.2, 101102.6, 101266.6, 
    101229.1, 101152.8, 101507.9, 101565.2, 101593.3, 101589.1, 101546.4, 
    101499.7,
  100643.7, 100747.8, 100843.8, 100973.5, 101094, 101211.7, 101332.1, 101506, 
    101615.9, 101619.1, 101670, 101686.8, 101682.9, 101663.6, 101618.1,
  100698.8, 100823.5, 100918.4, 101033.2, 101131.8, 101304.8, 101470.7, 
    101580.7, 101655.6, 101753.2, 101789.2, 101798, 101796.6, 101780.4, 
    101758.8,
  100684.7, 100822.7, 100939.6, 101092.8, 101252.9, 101443.3, 101621.7, 
    101793.6, 101878.6, 101907.6, 101916.8, 101922.7, 101921.6, 101914.7, 
    101901.1,
  100762.1, 100896, 101043.1, 101221.7, 101399.5, 101611.7, 101767.8, 
    101879.6, 101945.6, 101982.2, 102050.9, 102064.6, 102069.3, 102071.8, 
    102058,
  101586.9, 101627.8, 101671.8, 101657.1, 101629.4, 101525.7, 101356.9, 
    101238.5, 101153.3, 100785.7, 100800.1, 101011.8, 100839.6, 100405.4, 
    100247.5,
  101662.1, 101686.8, 101734.4, 101756.6, 101724.3, 101445.5, 101563.7, 
    101399.5, 101283.2, 101262, 101225.7, 101214.8, 101154.2, 99205.45, 
    99876.51,
  101677.8, 101772.9, 101831, 101866.6, 101663.8, 98156.95, 101586.5, 
    101731.6, 101637.2, 101509.6, 101420.7, 101380.1, 101323.2, 101271.5, 
    101184,
  101643.5, 101739.8, 101848.2, 101905, 101950.7, 101618.7, 97919.55, 
    101575.1, 101683.1, 101713.4, 101619.7, 101521.4, 101471.1, 101403.4, 
    101327.2,
  101627, 101749.6, 101887.3, 101961.9, 102025.8, 102025, 101752.9, 95540.44, 
    94959.12, 101681.3, 101864.6, 101716, 101682.6, 101574.8, 101573,
  101636.3, 101791.7, 101915.5, 102033.8, 102070, 102086, 102127.3, 102023.6, 
    101850.1, 102042.2, 102014.9, 101921.6, 101877.5, 101805.6, 101776,
  101643, 101823.9, 101977.2, 102080.5, 102134.9, 102221.2, 102256, 102308.6, 
    102316.5, 102247.5, 102188.2, 102143.9, 102080.6, 102029.4, 101983.7,
  101677.4, 101879.8, 102014.7, 102116.8, 102208.9, 102314.6, 102399.3, 
    102425.1, 102402.2, 102405.9, 102372.7, 102325.1, 102281, 102235.7, 
    102202.3,
  101724.1, 101947.2, 102107.6, 102292.4, 102433.6, 102543.8, 102605.2, 
    102643.8, 102643.6, 102606.3, 102557.7, 102513.7, 102464.1, 102418.7, 
    102380,
  101774.9, 102061.4, 102331.2, 102548, 102649, 102735.4, 102760.2, 102759.6, 
    102743.6, 102712.4, 102723.4, 102694, 102644, 102598.3, 102541.1,
  101910.9, 102035.5, 102190.2, 102301.7, 102414.1, 102478.7, 102494.3, 
    102512.4, 102472.1, 102071.4, 102052, 102209.4, 101914.1, 101343.8, 
    101071.4,
  102161.4, 102257.5, 102369.2, 102475.9, 102541.5, 102409.8, 102625.9, 
    102548.7, 102467.9, 102442.3, 102357.9, 102272.6, 102099, 100008.1, 
    100573.1,
  102319.8, 102438.8, 102511, 102591, 102448.5, 98931.6, 102526, 102750.5, 
    102674.3, 102557.2, 102414.5, 102325.4, 102165.9, 102039.5, 101887.3,
  102369.8, 102456.1, 102525.8, 102580.8, 102609.4, 102378.8, 98626.05, 
    102447.4, 102572.3, 102623, 102511.3, 102366.7, 102234.8, 102112, 102027.7,
  102383.2, 102470.6, 102539.1, 102611.5, 102660.8, 102659.5, 102474.3, 
    96225.42, 95565.39, 102435.8, 102607.2, 102446.5, 102348.3, 102195.3, 
    102193.8,
  102386.1, 102493, 102573.1, 102662.7, 102717.1, 102746.2, 102757.9, 
    102685.8, 102529.9, 102699.1, 102675.6, 102564.8, 102484.3, 102379.2, 
    102343.9,
  102390.6, 102524.4, 102616.6, 102679.5, 102753.5, 102816.9, 102858, 
    102897.2, 102886.7, 102809.9, 102746.9, 102699.2, 102627.2, 102573, 
    102536.9,
  102430.5, 102525.4, 102622.6, 102701.7, 102770.5, 102847.3, 102901.9, 
    102915.8, 102888.9, 102889.6, 102861.1, 102816.4, 102782.3, 102745.7, 
    102725.6,
  102462.9, 102581.9, 102734.5, 102874.8, 102974.6, 103012.5, 103022.8, 
    103031, 103023, 102984.1, 102943.4, 102910.5, 102879, 102857.8, 102840.5,
  102543.7, 102756.5, 102955.9, 103078.8, 103116.7, 103122.9, 103090.3, 
    103032.1, 103008.7, 102984.5, 103012.6, 102994.3, 102964, 102934.1, 
    102893.8,
  101501.5, 101490.3, 101523.8, 101584.9, 101707.6, 101872.3, 102039.6, 
    102229.9, 102407.3, 102213, 102402, 102750.4, 102618.9, 102183.6, 102023.5,
  101860.5, 101855.6, 101898, 101987, 102061.4, 102036.2, 102337.3, 102461.6, 
    102545.6, 102704, 102765.6, 102836.6, 102800.7, 100799.6, 101430.6,
  102125.6, 102167.2, 102201.6, 102304.1, 102191.8, 98776.62, 102476.1, 
    102737.1, 102801.1, 102821.2, 102831.5, 102824.8, 102766, 102718.7, 
    102652.1,
  102193.6, 102254.5, 102338, 102438.4, 102527, 102311.4, 98620.15, 102563, 
    102821.3, 102890.8, 102871, 102786.9, 102727, 102669.3, 102652.6,
  102220.8, 102289.7, 102374.8, 102479.1, 102574.6, 102674.1, 102537.4, 
    96320.02, 95646.94, 102686.8, 102909.7, 102777.9, 102704.9, 102627.8, 
    102705.6,
  102270.7, 102347.5, 102434.7, 102541.2, 102607.4, 102647.4, 102739.1, 
    102737.5, 102679.3, 102930.9, 102931.2, 102854.9, 102799.1, 102752.3, 
    102763.9,
  102268.4, 102354.9, 102446.1, 102526.5, 102611.4, 102725.6, 102812.2, 
    102929.5, 103014.1, 103017.4, 103003, 102960.5, 102900, 102856.5, 102829.5,
  102217.1, 102262.8, 102341.2, 102430, 102496, 102662.8, 102846.5, 102957.6, 
    103022.3, 103076.6, 103067, 103028.2, 102977, 102914.5, 102851.8,
  102191, 102244.6, 102343.7, 102491.7, 102604.7, 102750.3, 102907.8, 
    103046.1, 103113, 103118.4, 103086.4, 103028.6, 102943.8, 102842.3, 
    102730.4,
  102248.1, 102368.8, 102473.3, 102586.3, 102675.4, 102806.7, 102957, 
    103035.3, 103092.7, 103071.6, 103061.8, 102971, 102835.9, 102677.6, 
    102506.3,
  101290.9, 101057, 100857.2, 100701.7, 100646.2, 100650.4, 100686.3, 
    100792.5, 100937, 100789, 101066.8, 101524.2, 101555.7, 101366, 101408.4,
  101611.3, 101437.6, 101255.8, 101196.9, 101124.8, 100995.4, 101194.4, 
    101262.1, 101360.4, 101562.4, 101707.8, 101913.3, 102014.4, 100263.6, 
    101108.6,
  101836.8, 101764.9, 101660.1, 101657, 101399.4, 98055.21, 101607.5, 
    101847.8, 101899.7, 101978.1, 102086.5, 102220.9, 102335, 102436.2, 102534,
  101938.2, 101923.3, 101937.7, 101934.1, 102003.5, 101653.3, 98106.53, 
    101893.9, 102192.4, 102301, 102369.9, 102408.5, 102517, 102618.6, 102694,
  102020.1, 102055.1, 102106.9, 102155.8, 102210.8, 102297.4, 102033.6, 
    95871.72, 95297.28, 102261.2, 102544.7, 102517.5, 102579.4, 102606.8, 
    102727.6,
  102103.1, 102137, 102198.5, 102265.7, 102305.1, 102325.2, 102432.4, 
    102341.9, 102251.3, 102556.1, 102602, 102599.8, 102633.2, 102662.9, 
    102721.5,
  102090.2, 102151.9, 102267.6, 102314.6, 102388.7, 102448.6, 102482.9, 
    102579, 102636.9, 102603.5, 102604.4, 102614.2, 102620, 102648.9, 102679,
  101880.6, 102083.6, 102167.1, 102250.1, 102271.6, 102410.4, 102508.6, 
    102520.8, 102497, 102510.2, 102492.3, 102484.5, 102504.1, 102561.6, 
    102629.3,
  101648.3, 101887.3, 102001.4, 102165.8, 102330.8, 102469, 102478.2, 102488, 
    102417.4, 102315.5, 102223.2, 102185.6, 102193.2, 102269.5, 102385.1,
  101641.5, 101843.1, 102039, 102286.3, 102404.9, 102498.3, 102452.9, 
    102306.8, 102113.2, 101929.8, 101832.8, 101762.3, 101761.7, 101880, 
    102066.5,
  101814.8, 101525.5, 101206.4, 100903.4, 100677.5, 100474.9, 100252.6, 
    100175.2, 100187.8, 99930.71, 100085.4, 100501.5, 100547.4, 100392.7, 
    100468,
  101976.9, 101741.8, 101449.9, 101208.6, 100973.7, 100621.9, 100663.6, 
    100456.5, 100402.9, 100456.3, 100535.6, 100708.8, 100859.6, 99242.69, 
    100112.1,
  102054.5, 101905.8, 101719.3, 101537.7, 101122.8, 97681.36, 100973.5, 
    101026.8, 100882.1, 100831.1, 100849.9, 100967.2, 101130.3, 101298.7, 
    101481.4,
  102102.9, 101970.8, 101898.7, 101751.6, 101669.8, 101195.4, 97545.28, 
    101094, 101253.8, 101298.9, 101275.5, 101318.8, 101461.3, 101650.7, 101788,
  102133.9, 102054.9, 101973.8, 101907.7, 101851.1, 101818.2, 101443.4, 
    95286.99, 94763.75, 101466, 101688.7, 101648.3, 101753.3, 101836.6, 
    102024.9,
  102050.9, 102002.4, 101994.3, 101942.4, 101914, 101875.5, 101909.3, 
    101788.3, 101621.5, 101892.5, 101926.7, 101904.2, 101991.4, 102071.5, 
    102222.1,
  101876.8, 101842, 101928.7, 101887.6, 101893.4, 101889.1, 101862, 101922.7, 
    101997.3, 101969.3, 101997.4, 102062.3, 102127.8, 102209.2, 102324.4,
  101702.4, 101686, 101818.9, 101863.2, 101834, 101802.6, 101782.9, 101726.7, 
    101719, 101802.2, 101905.2, 101995.9, 102131.3, 102277.6, 102411.1,
  101730.6, 101763.7, 101876.6, 101943.5, 101944.2, 101866.2, 101738.5, 
    101655.1, 101596.3, 101570.8, 101638.3, 101812.6, 102001.9, 102180.2, 
    102377.7,
  101938, 102007.2, 102051.3, 102036.4, 101933.7, 101826.5, 101686.2, 
    101543.3, 101424.9, 101336.8, 101346.6, 101479.4, 101721.4, 101998, 
    102265.2,
  102477.1, 102308.9, 102107.3, 101925.8, 101739.5, 101575.2, 101308.4, 
    101147, 101141.3, 100819.5, 100890.4, 101185.8, 101109, 100812.1, 100751.1,
  102448.4, 102308.3, 102136.4, 102021.3, 101833.6, 101499.2, 101544.7, 
    101267.9, 101113.6, 101092.1, 101081.6, 101144.6, 101228, 99483.91, 
    100231.8,
  102355, 102264.3, 102124, 102102, 101814.8, 98270.16, 101596.4, 101674.1, 
    101471, 101304.7, 101182.1, 101168.3, 101217.2, 101291, 101377,
  102233.6, 102164.7, 102054.9, 102060.2, 102072, 101703, 97954.63, 101495.1, 
    101606.4, 101605.7, 101470.3, 101353.1, 101329.4, 101356.7, 101421.3,
  102107.2, 102060.4, 101981.8, 101977, 102063.9, 102036.2, 101792.6, 
    95608.48, 94986.61, 101614.5, 101757.2, 101576.7, 101530.2, 101441.9, 
    101501.7,
  101947.4, 101904.8, 101881.8, 101932.6, 101980.8, 101972.7, 102033.1, 
    101938.7, 101792.6, 101985.8, 101912.5, 101794.5, 101710, 101633.4, 
    101617.4,
  101792.7, 101796.5, 101838.3, 101937.2, 101963.6, 101980.7, 102002, 
    102043.4, 102094.9, 102069.9, 102018.4, 101970.4, 101892.9, 101829.7, 
    101793.2,
  101700.7, 101729.6, 101835, 101978.9, 101978, 102001.2, 102044.2, 102021.4, 
    101995.9, 102007.7, 102033.4, 102062.2, 102050.1, 102038.3, 102028.9,
  101689.2, 101737.8, 101882.9, 102002.7, 102060.7, 102068.4, 102066.9, 
    102070.8, 102090.8, 102062.2, 102025.5, 102072.5, 102124.2, 102160.3, 
    102184,
  101706.3, 101785.8, 101957.6, 102042.9, 102067.6, 102083.9, 102077, 
    102031.4, 102037.8, 102042.4, 102038.4, 102056.2, 102142.9, 102237.6, 
    102297.6,
  102434.1, 102542.3, 102614.5, 102647.2, 102679.6, 102654.2, 102521.6, 
    102369.4, 102221.7, 101793.6, 101812.1, 102024.1, 101804.2, 101313.8, 
    101113.1,
  102288.8, 102410.5, 102514.4, 102556.8, 102600.9, 102451.4, 102605.5, 
    102446.1, 102296.8, 102181.3, 102072.1, 102015.7, 101981.6, 100070.7, 
    100688.6,
  102073.6, 102256.6, 102397.8, 102469.8, 102418, 98953.48, 102442.5, 
    102650.7, 102509.3, 102380, 102219.5, 102115.2, 102020.9, 101974.7, 
    101903.4,
  101824.5, 102043.1, 102218.1, 102331.4, 102417.5, 102292.1, 98564.12, 
    102293.6, 102488.2, 102500.5, 102400.8, 102271.8, 102172.8, 102072.7, 
    101970.5,
  101591.4, 101826.7, 102030.8, 102193.1, 102309.4, 102402.2, 102298.2, 
    96247.2, 95513.33, 102360.2, 102540.8, 102414.1, 102323.5, 102185.1, 
    102092.2,
  101388.1, 101622.1, 101851.1, 102042.2, 102173.1, 102294.9, 102391.5, 
    102378.4, 102295.8, 102602.5, 102599.8, 102541.2, 102459.4, 102332.2, 
    102205.7,
  101211.4, 101451.9, 101693.8, 101926.2, 102084.7, 102217.9, 102373.2, 
    102495, 102597.3, 102630, 102649.7, 102630.6, 102558.6, 102453.4, 102307.4,
  101078.8, 101322.6, 101568.3, 101825.9, 101981.2, 102132, 102346.3, 102447, 
    102548.9, 102633, 102688, 102698, 102648.1, 102551.9, 102405.2,
  100988.2, 101235.5, 101488.8, 101778.3, 101974.2, 102141.2, 102341.3, 
    102507.9, 102636.8, 102695, 102724.8, 102747.2, 102720.5, 102643.9, 
    102503.2,
  100940.3, 101187.8, 101464.8, 101764.2, 101970.6, 102156.5, 102343.7, 
    102478.8, 102609.7, 102674.8, 102739.2, 102799.3, 102798, 102755.4, 
    102644.7,
  101862.5, 101925.9, 102004, 102157.6, 102356.4, 102532.6, 102602.4, 
    102632.8, 102576.3, 102178.1, 102185, 102398.9, 102229, 101746.3, 101532.1,
  101777.5, 101861.4, 101968.8, 102131, 102317.1, 102358, 102606.9, 102612.3, 
    102573, 102578.5, 102492.5, 102462.1, 102409.8, 100458.3, 101068.1,
  101626, 101788.4, 101916.6, 102089, 102176.3, 98855.5, 102444.3, 102757.2, 
    102718.9, 102669.8, 102630, 102603.5, 102561.2, 102507.1, 102368.3,
  101431, 101608.5, 101807.7, 101988.4, 102229.2, 102139.7, 98586.31, 
    102355.9, 102644.4, 102716.4, 102715.2, 102696.1, 102697.4, 102651.3, 
    102538.9,
  101249.4, 101417.7, 101627.8, 101863.3, 102108.1, 102339.5, 102254.9, 
    96335.49, 95596.53, 102447.3, 102803.1, 102755, 102777.5, 102697.2, 
    102656.5,
  101060.2, 101234.1, 101441.7, 101701.8, 101958.7, 102179.3, 102356, 
    102363.1, 102264.3, 102609.2, 102776.8, 102819.6, 102854.8, 102782.2, 
    102696.5,
  100869.9, 101060.5, 101263, 101536.2, 101823.6, 102082.9, 102248.5, 
    102415.6, 102522.7, 102614.3, 102786.3, 102875.1, 102892.8, 102834, 102697,
  100717.6, 100917.4, 101104.1, 101391.6, 101666.6, 101932.1, 102157.8, 
    102347.2, 102527, 102687.4, 102832.3, 102936.9, 102962.4, 102894, 102736.7,
  100648.1, 100823.1, 101005.4, 101291.3, 101579.4, 101857.2, 102112.4, 
    102388.8, 102605.7, 102743.5, 102883.5, 102991.1, 103021.5, 102963.1, 
    102798.3,
  100666.8, 100818.7, 101000.9, 101270.2, 101544.2, 101820.2, 102095.6, 
    102380.8, 102607.9, 102741.1, 102920.5, 103052, 103109.2, 103069.2, 
    102923.4,
  101588.4, 101585.4, 101620.9, 101640.2, 101660.4, 101673, 101652.1, 
    101685.2, 101760.2, 101512.7, 101676.3, 102037.1, 101952.5, 101598.2, 
    101458.2,
  101493.1, 101500.6, 101597, 101664.9, 101730.6, 101597.7, 101773, 101721.5, 
    101757.6, 101874.2, 101971.4, 102085.1, 102172.1, 100286.8, 101008.4,
  101386.3, 101445.8, 101587.7, 101690.2, 101657.9, 98202.57, 101766.5, 
    101937.9, 101954, 101983.2, 102061.2, 102162.2, 102282.6, 102315.3, 
    102299.3,
  101259.8, 101357.1, 101553, 101672.5, 101811.1, 101611.9, 97985.54, 
    101722.5, 101990.9, 102091.5, 102199, 102301.4, 102413.6, 102469.7, 
    102457.6,
  101150.3, 101270.7, 101473, 101648.5, 101785.2, 101902.8, 101760.7, 
    95767.13, 95170.82, 102020.3, 102362.8, 102413.7, 102518.4, 102515, 
    102547.9,
  101071.6, 101201.6, 101429, 101608, 101780.9, 101864.9, 102009.5, 101944.6, 
    101824.7, 102282, 102422.7, 102534.9, 102613.5, 102605.4, 102564.4,
  100994.4, 101128.7, 101379.4, 101559.8, 101766.3, 101887.2, 101971.5, 
    102090.7, 102226.7, 102341.6, 102505.7, 102633.9, 102679.1, 102648.9, 
    102560.2,
  100958.2, 101111.4, 101352, 101535.6, 101714.7, 101863.7, 102019.7, 
    102082.6, 102216.5, 102427.2, 102613.9, 102728, 102765.5, 102705.3, 
    102603.2,
  100925.4, 101076.8, 101307.3, 101529.3, 101697.3, 101883.1, 102060.5, 
    102232.1, 102417.4, 102559.9, 102718.7, 102814.6, 102838.2, 102769, 
    102659.3,
  100929.9, 101046.1, 101263.4, 101499, 101689.4, 101894.8, 102107.4, 
    102274.6, 102454.8, 102587.2, 102798.8, 102903.7, 102928.4, 102863.2, 
    102749.1,
  101522.8, 101524.9, 101603.1, 101708.8, 101855.7, 101934.3, 101855.2, 
    101739.7, 101657.5, 101267.5, 101326.2, 101629.9, 101540.4, 101226.3, 
    101179.5,
  101322.7, 101330.3, 101470.1, 101610.8, 101798.6, 101685.1, 101875.1, 
    101697.9, 101624.8, 101615.8, 101625.7, 101699.5, 101761, 99960.4, 
    100723.2,
  101099.7, 101184.1, 101354.7, 101578.8, 101641.8, 98221.16, 101671.2, 
    101816.8, 101718.7, 101700.4, 101701.9, 101760.1, 101867.1, 101932.6, 
    102027.2,
  100915.4, 101055.5, 101290.3, 101556.8, 101709.3, 101571.2, 97865.04, 
    101573.8, 101778.9, 101806.3, 101842, 101887.6, 101987, 102112.5, 102191.4,
  100796, 100992.7, 101281.8, 101568.8, 101738.3, 101775.3, 101672.2, 
    95593.84, 94996.94, 101776.6, 102039.3, 102062.1, 102152.5, 102205.5, 
    102324,
  100748.5, 101016.8, 101322, 101582.7, 101691.8, 101763.3, 101808.9, 
    101789.7, 101716.3, 102081.6, 102165, 102240, 102311.6, 102368.8, 102434.6,
  100781, 101089.9, 101395.2, 101614.1, 101714.8, 101780.1, 101836.9, 
    101980.2, 102124.8, 102192.1, 102302.1, 102390.4, 102440.9, 102477.5, 
    102509.4,
  100892.9, 101179.5, 101464.7, 101608.6, 101677.8, 101812, 101965.6, 
    102041.8, 102175.4, 102325.3, 102452.2, 102521.7, 102574.6, 102589.7, 
    102609.3,
  101026.3, 101309.2, 101542.1, 101661.1, 101811.3, 101966.1, 102106.9, 
    102251.9, 102402.2, 102499.4, 102587.4, 102646.7, 102675.3, 102682.1, 
    102689.4,
  101176, 101421.3, 101632.8, 101802, 101954, 102096.9, 102238.1, 102352.8, 
    102471.8, 102554.9, 102685.7, 102749.5, 102777.9, 102788, 102782.3,
  101513.7, 101430.7, 101355, 101275.9, 101219, 101205.9, 101267.4, 101365.9, 
    101487.3, 101269.4, 101423.7, 101789.9, 101741.9, 101446.4, 101405.3,
  101409.8, 101291.8, 101222, 101122.3, 101071.2, 101017.4, 101317.8, 
    101384.4, 101472.9, 101579.8, 101637.3, 101754.7, 101836.6, 100051.9, 
    100832.5,
  101339.4, 101231, 101159.6, 101102.6, 101010, 97744.6, 101291.7, 101565.1, 
    101573.4, 101616.6, 101637.4, 101683, 101788.4, 101883.7, 102013,
  101336.7, 101252.1, 101214.4, 101190.6, 101247.6, 101099.1, 97555.92, 
    101326.2, 101642.1, 101669.1, 101661.9, 101642.7, 101746.4, 101904.2, 
    102075.9,
  101452.1, 101410, 101391.5, 101432.3, 101465.7, 101484.2, 101321.6, 
    95377.35, 94701.55, 101519.2, 101706.7, 101651.7, 101754.6, 101879.4, 
    102124.8,
  101631.4, 101627.4, 101606.3, 101609.2, 101601.4, 101596.4, 101619.2, 
    101579.8, 101508, 101760.5, 101746, 101751.2, 101847.8, 102007, 102209.5,
  101832.6, 101827.8, 101799.1, 101794.9, 101783.6, 101795.6, 101794.3, 
    101853, 101882.4, 101852.5, 101872.2, 101908.6, 102002.4, 102161.6, 
    102345.7,
  102038.1, 102015.7, 101967.7, 101937.4, 101908.5, 101948.9, 101987.6, 
    101968.3, 101990.8, 102032.5, 102058.1, 102116.8, 102233.6, 102389.7, 
    102571.6,
  102218.5, 102221.6, 102196.9, 102201.7, 102197.4, 102214.1, 102218.2, 
    102244.8, 102250, 102250.3, 102283.3, 102362.3, 102472.1, 102612.4, 
    102766.1,
  102390.7, 102398.6, 102394.1, 102406.8, 102391.3, 102387.9, 102398.8, 
    102388.2, 102400.7, 102409.4, 102494.7, 102584.4, 102694.6, 102825.8, 
    102941.4,
  102995, 102890.4, 102770.2, 102607.6, 102415, 102257.3, 102100.7, 101944.3, 
    101785.3, 101283.7, 101203.3, 101347.4, 101111.6, 100747, 100720.5,
  103041.1, 102901.4, 102779.8, 102618.4, 102424.8, 102047.2, 102156.2, 
    101927.1, 101744.8, 101635.9, 101486, 101395.5, 101306.3, 99437.46, 
    100224.2,
  103041.8, 102921, 102792.8, 102687.1, 102341.9, 98667.38, 101952.4, 
    102094.6, 101888.5, 101719.5, 101550, 101476.3, 101426.2, 101447.3, 
    101515.1,
  103062, 102939.7, 102804, 102693, 102541.6, 102126.1, 98206.48, 101729.2, 
    101818, 101768.2, 101619.6, 101534.3, 101531.7, 101588.6, 101685,
  103115.7, 103015.9, 102875.7, 102750.7, 102632.2, 102465.6, 102093.6, 
    95761.34, 94963.41, 101562.4, 101685, 101578.5, 101610.6, 101653.1, 101836,
  103167.6, 103071.5, 102944.6, 102809.2, 102649.1, 102541.6, 102382.3, 
    102133.7, 101805.8, 101805.9, 101700.2, 101648.2, 101699.3, 101794.2, 
    101942.9,
  103218.5, 103154, 103043.4, 102934.8, 102770.8, 102667.1, 102499.9, 
    102340.8, 102129.6, 101901.5, 101782.6, 101766.2, 101810, 101930.3, 
    102062.9,
  103265.7, 103209.9, 103119.5, 103051.8, 102891.7, 102772.9, 102633.2, 
    102435.8, 102250.3, 102093.5, 101966.9, 101949.1, 102004.9, 102124.9, 
    102263.8,
  103312, 103276.6, 103219.1, 103190.4, 103111.1, 102982.2, 102804.5, 
    102658.4, 102498.9, 102356.9, 102247.3, 102228.3, 102273.1, 102374.9, 
    102493.1,
  103357.8, 103300, 103252.8, 103252.1, 103182, 103073.9, 102934.5, 102775.7, 
    102649.5, 102538.1, 102516.2, 102509.7, 102541.3, 102618.9, 102688.5,
  102993.3, 102893.6, 102819.4, 102699.9, 102574.2, 102449, 102239.4, 
    102065.3, 101910.5, 101356.9, 101272.2, 101376.9, 101106.2, 100631, 
    100474.5,
  102950.8, 102826.1, 102763.5, 102666.4, 102545.8, 102151, 102290.9, 
    101969.1, 101750, 101610.1, 101450.4, 101305, 101178.5, 99223.28, 99933.62,
  102890.1, 102765.7, 102724.7, 102672.1, 102393.3, 98795.66, 102013.3, 
    102201.7, 101924.4, 101660.6, 101429.6, 101296.5, 101179.5, 101175.5, 
    101177.9,
  102811, 102669.1, 102649.4, 102599.6, 102587.8, 102159.3, 98339.7, 
    101745.9, 101778.6, 101707, 101511.7, 101363.5, 101294.2, 101309.2, 
    101390.2,
  102725, 102603.6, 102592.5, 102574.1, 102585.4, 102527.9, 102174.1, 
    95848.83, 95120.89, 101603.3, 101699.4, 101516.9, 101496.6, 101478.6, 
    101644.3,
  102615, 102468.6, 102459.3, 102523.6, 102518.6, 102529.3, 102473.5, 
    102246.8, 101912.5, 101969.7, 101864.9, 101760.8, 101733, 101750.1, 101856,
  102495.1, 102377.7, 102327.2, 102467.4, 102517.6, 102570.3, 102510, 
    102485.8, 102367.5, 102175.7, 102067.2, 102020.7, 101994.9, 102037.7, 
    102112.1,
  102383.9, 102219.6, 102146.1, 102318.8, 102443.7, 102556.1, 102584.9, 
    102494.5, 102406.3, 102357.8, 102296.4, 102267.8, 102271.8, 102313.7, 
    102388.2,
  102270.2, 102099, 102014.2, 102137, 102376.2, 102552, 102639.6, 102667.7, 
    102642.8, 102574.2, 102521.3, 102512.1, 102522.8, 102565.3, 102618.1,
  102145.1, 101924.2, 101787.4, 101873.1, 102190.2, 102460.7, 102623.1, 
    102646.3, 102668.4, 102659.5, 102705.6, 102712.7, 102727.3, 102754.7, 
    102781.6,
  100784.8, 100619.3, 100791.2, 101068.8, 101226.3, 101339.8, 101268.6, 
    101227.3, 101121, 100661.1, 100658.5, 100930.5, 100860.7, 100522.3, 
    100430.6,
  100717.3, 100580.4, 100808.4, 101097.3, 101280.9, 101145.7, 101358.7, 
    101168.3, 100991.4, 100900.3, 100837.5, 100860.6, 100933.5, 99134.29, 
    99893.66,
  100671.7, 100582.6, 100844.6, 101171, 101154.8, 97799.48, 101188.7, 
    101386.2, 101219.8, 101022.7, 100897.6, 100917.7, 100987.6, 101101.3, 
    101119.3,
  100652.4, 100592.2, 100863.1, 101166.6, 101373.2, 101167.4, 97555.37, 
    101132.9, 101191.9, 101200.5, 101110, 101077.2, 101127.3, 101192.5, 
    101224.9,
  100662.5, 100646.4, 100894.3, 101229.5, 101439.1, 101565.4, 101354.7, 
    95193.13, 94676.02, 101191.2, 101361, 101248.5, 101283.8, 101249, 101334.6,
  100681.4, 100703.2, 100899.7, 101295, 101502, 101666.2, 101762.2, 101685.6, 
    101457.8, 101633.5, 101580.7, 101509, 101498.7, 101482.2, 101498.3,
  100715.5, 100789.2, 100966, 101386.2, 101640.7, 101855.2, 101901.9, 102007, 
    102014, 101912.7, 101836.6, 101802.5, 101755.7, 101744.7, 101722.5,
  100791.7, 100894.8, 101055.6, 101459.7, 101711.3, 101979.7, 102121.5, 
    102146, 102137.2, 102158.3, 102127, 102088.3, 102047.1, 102011.4, 101971.4,
  100888.3, 101016.2, 101205.4, 101589, 101898.5, 102180.4, 102332.5, 
    102437.8, 102473.1, 102444.3, 102406.3, 102365.4, 102320.3, 102261.1, 
    102190.5,
  101003.8, 101127.3, 101334.4, 101701.1, 102040.4, 102332.4, 102519.9, 
    102590, 102626.4, 102620.8, 102661.4, 102630.1, 102586, 102522.6, 102444.4,
  101131.3, 101248.4, 101319.2, 101301.3, 101275, 101197, 101041.9, 100955.8, 
    100951.9, 100590.8, 100693.3, 101038.4, 100978.4, 100690.9, 100663.4,
  101356.8, 101438, 101454.4, 101438.6, 101373.6, 101053, 101200.3, 100948.1, 
    100830.6, 100897.6, 100954.8, 101057.7, 101160.5, 99337.79, 100131.5,
  101564.2, 101643.1, 101629.7, 101613.4, 101305, 97832.73, 101082.3, 
    101276.5, 101121.6, 100975.8, 100953.6, 101039.6, 101146.6, 101257.2, 
    101329.5,
  101708.1, 101756.1, 101797, 101720.3, 101678, 101225.5, 97514.8, 100939.3, 
    100997.6, 101047.5, 100965.5, 100988.9, 101088.4, 101221.9, 101341.2,
  101888.2, 101925.9, 101970, 101933.4, 101857, 101762.1, 101369.6, 95125.34, 
    94435.27, 100866.4, 101022.3, 100905.8, 100988.5, 101052.5, 101249.3,
  102081.6, 102132.6, 102148.5, 102141, 102055.1, 101941.2, 101841.3, 
    101575.8, 101200.8, 101202.6, 101041.6, 100938.2, 100943.5, 100994.6, 
    101131.2,
  102275.1, 102340.4, 102351.4, 102348, 102295.8, 102222.8, 102045.9, 
    101926.4, 101730.5, 101422.2, 101144.7, 100996.8, 100929.4, 100958.4, 
    101039.3,
  102479.1, 102546.2, 102566.8, 102563.4, 102502.7, 102446.9, 102311.4, 
    102102.9, 101875, 101668.1, 101395.1, 101146.3, 101005.6, 100977, 101021.8,
  102714.3, 102805.8, 102856.4, 102881, 102846.9, 102749.7, 102586.1, 
    102431.4, 102222.6, 101968.7, 101702.7, 101413.9, 101181.9, 101070.6, 
    101057.6,
  102974.3, 103080.4, 103143.5, 103145.7, 103074.2, 102981.5, 102832.1, 
    102631.6, 102435.1, 102214.2, 102023, 101766.6, 101483.8, 101289.6, 
    101194.6,
  101960.2, 101882.1, 101798.4, 101624, 101521.4, 101410.7, 101241.8, 
    101153.7, 101141.1, 100756.9, 100792.4, 100993, 100739.6, 100295.6, 
    100144.7,
  102047, 101950.4, 101840.3, 101679.9, 101517.6, 101144.2, 101305.5, 101034, 
    100906.8, 101019.6, 101047.2, 101065.1, 100980.6, 99034, 99704.4,
  102088, 102026.5, 101925.6, 101812.9, 101421.1, 97868.3, 101026.8, 
    101279.4, 101074.1, 100996.1, 101032, 101094.3, 101081.4, 101070.5, 
    101021.2,
  102128.6, 102052.5, 101983.1, 101876.9, 101731.5, 101241.9, 97437.67, 
    100817.7, 100934.1, 100981.5, 100991.2, 101089, 101143.1, 101188.3, 
    101205.3,
  102242.6, 102174.2, 102095.1, 101986.7, 101862.9, 101703.6, 101264, 
    94993.97, 94232.23, 100747.7, 100990.8, 101040.1, 101181.4, 101218.9, 
    101339.3,
  102367.4, 102300.1, 102199.6, 102103.2, 101935.1, 101798.7, 101636.1, 
    101335, 100976.9, 100981.5, 100943, 101019.2, 101162.3, 101271.1, 101389.3,
  102507.4, 102473, 102364.6, 102258.2, 102117.9, 101971, 101739.4, 101590.8, 
    101387.6, 101103, 100951.3, 101019.9, 101116.8, 101260.5, 101395.8,
  102678.4, 102646, 102566.4, 102448.9, 102285.6, 102120.2, 101913.9, 
    101660.1, 101427.8, 101248.1, 101048.1, 100997.3, 101092.1, 101226.2, 
    101380.4,
  102854.6, 102858.2, 102803.8, 102731, 102583.1, 102366.6, 102097.2, 
    101889.4, 101672, 101431.9, 101219.9, 101040.4, 101055, 101175.8, 101312.4,
  103068.3, 103057.5, 103020.4, 102937.7, 102761.5, 102560, 102322.1, 
    102021.4, 101798.8, 101561.9, 101390.3, 101187.8, 101053.2, 101115.5, 
    101238.3,
  101794.4, 101803, 101802.1, 101736, 101716.1, 101686.7, 101574.7, 101518.4, 
    101466.3, 101059.9, 101125.1, 101401, 101229.1, 100770.2, 100576.8,
  101852.8, 101850.9, 101837, 101768.2, 101693.8, 101429.5, 101605.4, 
    101397.4, 101271.3, 101285.1, 101290, 101342.8, 101311.9, 99352.42, 
    99965.08,
  101852.9, 101910.2, 101896.3, 101870.1, 101578.6, 98006.1, 101298.7, 
    101542.3, 101318.6, 101215.5, 101183.4, 101251.3, 101238.7, 101215.4, 
    101100.8,
  101863.6, 101893.7, 101906.2, 101893.1, 101792.4, 101449.4, 97544.16, 
    101050.5, 101203.3, 101165.2, 101116.6, 101149.5, 101166.3, 101150.1, 
    101035.4,
  101958.7, 101979.9, 101973.5, 101942.7, 101869.6, 101734.7, 101401.9, 
    95071.4, 94260.88, 100906.9, 101084.6, 101073, 101109.4, 101055.7, 100990,
  102090.7, 102097.2, 102061.1, 102004.9, 101885, 101797.8, 101617.3, 
    101386.1, 101075.7, 101097.9, 101005.6, 101026.4, 101075.9, 101038.3, 
    100935.1,
  102225.1, 102245.4, 102203.6, 102134, 102016.2, 101877, 101670.8, 101525.2, 
    101333.4, 101085.6, 100966.7, 101031.3, 101067.1, 101042.7, 100936.9,
  102394.7, 102399.6, 102374, 102301, 102169.6, 102015.2, 101783.5, 101544.7, 
    101340.9, 101160.4, 101026.6, 101027.6, 101079.1, 101074.2, 100999.6,
  102543.7, 102591, 102583, 102536, 102425, 102214.2, 101953.2, 101728.1, 
    101518.1, 101281.5, 101103.4, 101024.1, 101090.8, 101098.5, 101052.8,
  102723.1, 102767.2, 102765.3, 102712.7, 102563.5, 102391.3, 102161.1, 
    101879.1, 101651, 101419.6, 101232.6, 101087.1, 101080.3, 101138, 101120.3,
  101878.3, 101892.4, 101894.5, 101875.5, 101876.3, 101850, 101789.6, 
    101793.2, 101795.4, 101425.1, 101493.8, 101791.2, 101668.8, 101261.3, 
    101130.5,
  102054.4, 102042.8, 102006.8, 101960.6, 101902.1, 101686.5, 101863.7, 
    101734, 101660, 101683.2, 101672.3, 101722.4, 101731.3, 99830.93, 100503.6,
  102150.1, 102143.5, 102119.3, 102072.4, 101816.6, 98227.12, 101631.6, 
    101859.3, 101701.1, 101616.1, 101546.7, 101580.1, 101615, 101657.3, 
    101673.7,
  102100.2, 102113.4, 102133.9, 102117.8, 102015.4, 101702.5, 97798.24, 
    101396.4, 101562.3, 101529.3, 101451.6, 101429.8, 101463.6, 101541.6, 
    101580.8,
  102139.5, 102168.7, 102150, 102149.8, 102079.8, 101966.8, 101667.3, 
    95348.98, 94539.79, 101253.1, 101417.4, 101341.1, 101361.2, 101367, 
    101453.4,
  102201.7, 102210, 102177.8, 102152.8, 102063, 101999.6, 101862.5, 101664.7, 
    101396.8, 101456.6, 101347.4, 101273.2, 101269, 101279.4, 101317.6,
  102233.7, 102252.2, 102221.3, 102187.3, 102112.2, 102041.7, 101887.8, 
    101770.5, 101618.9, 101438.2, 101312.6, 101236.4, 101201, 101190.7, 
    101182.6,
  102273.2, 102272.2, 102241.5, 102201.7, 102124.3, 102046.5, 101902.1, 
    101714.9, 101570.2, 101446.8, 101322.3, 101204.8, 101133.9, 101092.8, 
    101042.2,
  102268.1, 102304.6, 102284.5, 102249.5, 102188, 102051.6, 101892.4, 
    101736.2, 101589.9, 101433.5, 101299.8, 101160.4, 101048, 100963, 100873.2,
  102261, 102272, 102247.2, 102204, 102077.9, 101951.9, 101814.3, 101621.8, 
    101487.2, 101350.5, 101267.5, 101123.5, 100975.8, 100869, 100749.2,
  102316.9, 102321.1, 102323.6, 102298.4, 102292.6, 102241.7, 102164.5, 
    102126.4, 102048.2, 101588.9, 101556.4, 101751.9, 101495.5, 100996.5, 
    100793.6,
  102420.4, 102381.9, 102340.8, 102285.9, 102209, 101962.8, 102120.1, 
    101950.9, 101861, 101858.1, 101797.3, 101755.8, 101696.3, 99694.81, 
    100316.1,
  102395.2, 102357, 102300.9, 102238, 102000.5, 98420.38, 101727.5, 101992.4, 
    101853, 101709.5, 101630.8, 101619.7, 101606.5, 101594.3, 101572,
  102219, 102140.9, 102047.8, 101968.3, 101888.6, 101593.1, 97800.76, 
    101203.5, 101449.8, 101477, 101430.7, 101374.6, 101409.4, 101451.3, 101503,
  102097.5, 101972.5, 101810.9, 101696.5, 101588.3, 101496.6, 101257.8, 
    95175.62, 94284.15, 100820.8, 101147.9, 101064, 101140.3, 101166.5, 
    101310.7,
  101961.9, 101767, 101574.8, 101437.3, 101284, 101200, 101110.6, 100921.8, 
    100686.7, 100841.9, 100795.6, 100769.9, 100835.5, 100913.8, 101053.3,
  101762.6, 101570.4, 101390.2, 101272.4, 101125, 100993.6, 100869.2, 100774, 
    100655.6, 100517.8, 100489.8, 100497.8, 100532, 100625.9, 100783.2,
  101581.3, 101410.5, 101279.7, 101119.5, 100960.8, 100822.3, 100669.8, 
    100473.7, 100313.8, 100236.4, 100191.4, 100198.5, 100269.6, 100379.7, 
    100564.8,
  101463, 101355.2, 101220.2, 101070.6, 100945.4, 100750.2, 100545.8, 
    100318.2, 100102.8, 99926.14, 99862.53, 99886.95, 99989.45, 100136, 
    100336.9,
  101419.5, 101288.5, 101149.6, 100997.5, 100818.2, 100626.7, 100426.2, 
    100105.7, 99818.39, 99604.1, 99558.98, 99591.7, 99719.71, 99930.47, 
    100170.8,
  102573.1, 102452.2, 102311.4, 102168, 102085, 102024.8, 102014.6, 102068.4, 
    102099.8, 101739.7, 101816.2, 102115, 101989.4, 101562.3, 101415.1,
  102527.9, 102377.4, 102200.7, 102034.9, 101888.1, 101639.2, 101840, 
    101780.7, 101794.9, 101905.7, 101919.2, 101972.7, 101996, 100102.6, 
    100733.4,
  102417.9, 102253, 102033.9, 101842.2, 101550.4, 98087.77, 101347.6, 
    101708.2, 101604.1, 101573.4, 101601.3, 101654.3, 101689.4, 101715.6, 
    101731.5,
  102276.5, 102056.6, 101780, 101559.1, 101413.7, 101156.8, 97565.23, 101014, 
    101363.8, 101436.6, 101387.5, 101347.8, 101378.1, 101417.3, 101452.6,
  102112.1, 101828, 101559.6, 101357.2, 101349.3, 101317.8, 101133.4, 
    95172.78, 94312.09, 100910.3, 101218.4, 101076.8, 101095.6, 101040.8, 
    101120.3,
  101852.1, 101558.9, 101322.9, 101286, 101233.7, 101230.1, 101197, 101035.7, 
    100895.2, 101088.7, 100984.4, 100891.5, 100846.2, 100771.8, 100775,
  101605, 101375.9, 101280.4, 101238.3, 101182.5, 101120.8, 101094, 101122.6, 
    101018.5, 100820, 100709, 100604.3, 100513.6, 100451.2, 100434.7,
  101457.2, 101331.4, 101231.2, 101191.1, 101129, 101175.6, 101139.6, 
    100956.3, 100777.5, 100605, 100397.3, 100216.4, 100108.4, 100058.2, 
    100065.8,
  101428.5, 101326.6, 101280.7, 101269.5, 101308.1, 101256.1, 101113.4, 
    100916.8, 100628.9, 100294.6, 100042.7, 99860.57, 99745.89, 99702.35, 
    99712.34,
  101441.6, 101366.6, 101331, 101356.2, 101328.9, 101254.8, 101071.7, 
    100743.9, 100404.2, 100076.1, 99817.3, 99595.04, 99477.29, 99454.16, 
    99471.2,
  103096.3, 103029.8, 102918.4, 102719, 102504.8, 102271.1, 102073.9, 
    102014.1, 101974.1, 101542.2, 101513.7, 101702.9, 101479.3, 100963.8, 
    100753.7,
  102980.9, 102873.2, 102713.1, 102501.5, 102253.4, 101855.5, 101954.9, 
    101837.4, 101744.5, 101787.5, 101710, 101669.8, 101596.2, 99641.89, 
    100233.9,
  102760.3, 102654.1, 102447.8, 102254.9, 101907.3, 98397.59, 101647, 
    101986.3, 101800.4, 101698, 101607.3, 101565.6, 101503.8, 101460, 101386.3,
  102558.5, 102394, 102168.5, 101985.8, 101883.3, 101709.6, 98025.77, 
    101373.7, 101650, 101694.6, 101581.1, 101470.8, 101430.1, 101387.9, 
    101350.8,
  102327.3, 102141.8, 101954.3, 101901.4, 102073.4, 102040.2, 101760.5, 
    95576.6, 94687.64, 101295.2, 101520.4, 101322.7, 101291, 101188.3, 
    101204.7,
  102079.9, 101894.4, 101819.5, 102037.6, 102020.9, 102065.8, 102007.4, 
    101741.9, 101514.4, 101605, 101419, 101259.7, 101176.1, 101068.6, 101035,
  101856.8, 101806.1, 101976.3, 102035.7, 102024.2, 102021.6, 101950.8, 
    101891.6, 101697.8, 101431.3, 101283.5, 101152.3, 101031.2, 100919.8, 
    100858.5,
  101793.5, 101952.6, 101953.1, 101993.4, 101990.5, 101988.3, 101858.1, 
    101621.2, 101420.9, 101286, 101124.8, 100975.8, 100839.5, 100702, 100606.1,
  101894.6, 101993.4, 102073.9, 102108.3, 102081.8, 101944.7, 101755, 
    101566.1, 101331, 101104.1, 100947, 100804.8, 100621.4, 100431, 100286.4,
  101988.1, 102099, 102136.6, 102105.2, 101986.8, 101843.8, 101627.8, 
    101355.8, 101126.2, 100988.2, 100851.8, 100665.1, 100419.8, 100189.1, 
    100023.5,
  102899.8, 103061.4, 103223, 103306.5, 103361, 103331, 103221.9, 103161.7, 
    103128.2, 102727, 102746.2, 102958.6, 102707.6, 102088.7, 101775.2,
  102803.3, 102932.6, 103061.1, 103138.9, 103132.2, 102912.2, 103052.4, 
    102927.5, 102874.7, 102976.7, 102941.8, 102904, 102773.3, 100666.5, 
    101124.3,
  102640.7, 102783.4, 102870.1, 102942.4, 102803.8, 99338.18, 102617.6, 
    103041.4, 102934.2, 102868.4, 102783.7, 102748.6, 102605.3, 102462.7, 
    102260.5,
  102478.4, 102576.1, 102634.5, 102667, 102662.1, 102463.1, 98830.02, 
    102367.7, 102708.8, 102768.3, 102675.1, 102537.4, 102441.5, 102305.4, 
    102112.7,
  102303.5, 102372.4, 102413, 102413.9, 102528.7, 102558.3, 102451.1, 
    96426.16, 95552.62, 102243.5, 102533.2, 102332.4, 102249, 102048.4, 
    101941.6,
  102149.7, 102177.8, 102180.6, 102264, 102329.5, 102450.9, 102508.2, 
    102389.1, 102305.7, 102490.4, 102345.9, 102175.7, 102043.1, 101850, 
    101717.4,
  101942.6, 101967.3, 102018.2, 102129.9, 102218.6, 102284.4, 102403.1, 
    102522.1, 102449.8, 102253.2, 102127.4, 101979.1, 101807.1, 101636.5, 
    101469.1,
  101750.4, 101779.5, 101873.1, 102008.1, 102130.5, 102330.6, 102388.8, 
    102302.1, 102197.3, 102106.5, 101953.7, 101792.9, 101636.3, 101451.4, 
    101255.2,
  101478.2, 101625.3, 101804.9, 102002.7, 102198.7, 102295.3, 102311.2, 
    102265.5, 102113.9, 101917.1, 101788.6, 101660.6, 101465.4, 101245.6, 
    101017.7,
  101399.7, 101560.1, 101783.5, 102036.9, 102198.8, 102262.1, 102235.1, 
    102067.3, 101917.3, 101809.5, 101708, 101533.4, 101308.3, 101056.1, 
    100796.4,
  101241.6, 101374.2, 101564.4, 101786.9, 102040.8, 102277.1, 102508.2, 
    102768.7, 102980.8, 102774.1, 102943.7, 103278.9, 103167.7, 102773.3, 
    102617.8,
  101209.9, 101314.7, 101483, 101716.6, 101929.1, 102030.6, 102428.5, 
    102593.8, 102759.5, 102957.6, 103047.8, 103148.8, 103195.5, 101276.4, 
    101886.6,
  101123.2, 101250.6, 101413.2, 101654.7, 101731.5, 98556.63, 102098.1, 
    102591.7, 102651.1, 102748, 102834.6, 102937.3, 102975.8, 102975.3, 
    102952.8,
  101004.6, 101110.7, 101286.4, 101494.1, 101754.7, 101653.9, 98304.05, 
    101959.5, 102441.5, 102563.2, 102651.5, 102685.1, 102757.6, 102783.2, 
    102757.5,
  100874.2, 100970.8, 101124.7, 101338.7, 101584.7, 101826.6, 101748.2, 
    96050.26, 95366.6, 101980.1, 102412.3, 102407.4, 102486.9, 102490.7, 
    102512.5,
  100760.7, 100830.8, 100954.8, 101152.9, 101382.6, 101573.5, 101802.6, 
    101763.2, 101764.6, 102123.1, 102191, 102228.9, 102293.4, 102282.3, 
    102300.2,
  100645, 100721.5, 100839.1, 100994.4, 101217.2, 101397.4, 101558.6, 
    101763.4, 101904.1, 101944.7, 102038.9, 102098.1, 102118.5, 102111.9, 
    102077.6,
  100546.4, 100630.4, 100722, 100866.9, 101015.5, 101208.9, 101380, 101515.4, 
    101687.4, 101867.8, 101969.9, 102008.4, 102016.4, 101964.2, 101878.5,
  100468.5, 100576.6, 100667.7, 100786, 100917.7, 101083.5, 101303.3, 
    101538.8, 101718.6, 101818.5, 101902.9, 101924.2, 101878.8, 101760, 
    101605.3,
  100458.9, 100511.2, 100600.4, 100712.4, 100873.3, 101131.4, 101397.5, 
    101592.5, 101748.3, 101824.2, 101885.5, 101841.3, 101720.6, 101538.7, 
    101325,
  100144.7, 100066.2, 100019, 100011, 100073.8, 100144.7, 100249.9, 100405.8, 
    100593.5, 100463.5, 100740.6, 101254.5, 101350.4, 101201.7, 101263,
  99958.05, 99868.05, 99813.88, 99808.32, 99834.05, 99798.5, 100085.8, 
    100224.2, 100393.3, 100639.6, 100848.9, 101136.2, 101372.6, 99744.09, 
    100561.1,
  99759.93, 99682.14, 99641.36, 99636.18, 99588.66, 96335.98, 99813.62, 
    100190.9, 100343.7, 100535.7, 100744.1, 100985, 101240.1, 101403, 101588.3,
  99646.67, 99571.98, 99523.55, 99502.38, 99624.27, 99477.45, 96115.05, 
    99798.2, 100240.4, 100451.1, 100654.4, 100834.6, 101083.7, 101316.1, 
    101496.3,
  99613.5, 99539.33, 99474.55, 99506.48, 99607.18, 99772.2, 99667.76, 
    94028.91, 93503.78, 100123.1, 100599.7, 100716.2, 100931, 101073.3, 
    101280.6,
  99614.07, 99557.77, 99505.66, 99553.45, 99641.71, 99749.34, 99938.5, 
    99914.55, 99903.06, 100332.1, 100476.9, 100619.6, 100790.6, 100930.5, 
    101073,
  99662.62, 99601.98, 99587.6, 99636.2, 99763.59, 99871.59, 99983.58, 
    100190.6, 100313.6, 100347.2, 100461.8, 100591.3, 100693.6, 100794.3, 
    100887.2,
  99787.33, 99749.42, 99721.03, 99776.76, 99874.38, 100022.8, 100122.3, 
    100185.5, 100274.1, 100406.7, 100510, 100613.4, 100753.8, 100865.2, 
    100952.5,
  100004.3, 99972.62, 99983.42, 100034.5, 100127.6, 100231, 100336.5, 
    100476.6, 100590.1, 100689.4, 100789.4, 100897.6, 100980.6, 101023.8, 
    101028.5,
  100413.9, 100338.7, 100341.8, 100389.9, 100449.5, 100555.5, 100649.5, 
    100727.9, 100806.3, 100890, 100995.2, 101041.5, 101041.4, 101016.7, 
    100956.1,
  99718.15, 99544.93, 99386.27, 99254.33, 99151.25, 99079.59, 99033.12, 
    99051.94, 99101.71, 98839.81, 98937.69, 99223.94, 99083.79, 98698.29, 
    98564.96,
  99586.02, 99387.12, 99217.08, 99061.09, 98916.18, 98655.88, 98808.72, 
    98777.59, 98800.88, 98892.52, 98962.64, 99054.09, 99100.66, 97304.24, 
    97951.45,
  99519.84, 99330.91, 99139.87, 98987.45, 98700.44, 95250.13, 98437.59, 
    98636.88, 98621.94, 98684.96, 98768.86, 98870.46, 98962.3, 99005.02, 
    99026.72,
  99543.36, 99326.98, 99135.8, 98981.81, 98804.53, 98447.43, 94795.49, 
    98244.2, 98507.28, 98574.52, 98651.85, 98733.23, 98839.67, 98935.88, 
    99004.72,
  99612.8, 99440.51, 99271.69, 99110.98, 98943.03, 98761.86, 98469, 92553.81, 
    91902.12, 98333.32, 98622.27, 98655.82, 98761.45, 98809.05, 98944.25,
  99728.93, 99557.35, 99409.68, 99276.14, 99106.25, 98951.95, 98806.37, 
    98659.31, 98460.52, 98628.48, 98642.97, 98686.32, 98782.9, 98857.85, 
    98966.5,
  99875.9, 99735.62, 99605.55, 99502.14, 99384.52, 99256.45, 99100.58, 
    99015.1, 98930.94, 98860.95, 98861.91, 98893.84, 98931.48, 98986.92, 
    99054.59,
  100021.2, 99898.45, 99788.1, 99713.84, 99612.76, 99531.77, 99416.05, 
    99320.52, 99267.22, 99260.44, 99256.53, 99269.73, 99298.32, 99324.2, 
    99345.41,
  100121.3, 100048.7, 99989.24, 99964.14, 99915.6, 99830.69, 99750.09, 
    99716.78, 99679.15, 99653.88, 99642.59, 99638.16, 99625.88, 99616.07, 
    99593.48,
  100176.7, 100080, 100043, 100060.3, 100026.1, 99986.16, 99933.95, 99886.84, 
    99885.52, 99858.3, 99878.63, 99863.48, 99818.54, 99768.43, 99691.63,
  100345.3, 100349.6, 100344.3, 100302.4, 100252.2, 100121.8, 99954.83, 
    99804.43, 99627.25, 99094.61, 98975.74, 99086.52, 98835.13, 98373.87, 
    98213.29,
  100247.3, 100220.9, 100193.8, 100155.3, 100084, 99763.16, 99871.62, 
    99627.35, 99390.28, 99251.01, 99043.01, 98914.98, 98789.01, 96888.3, 
    97458.66,
  100084.6, 100071.2, 100034.5, 100044.3, 99856.62, 96372.05, 99512.57, 
    99680.38, 99399.4, 99206.36, 98968.92, 98837.63, 98692.59, 98601.48, 
    98486.73,
  99884.62, 99857.59, 99831.89, 99851.55, 99861.2, 99606.99, 95855.62, 
    99210.91, 99328.14, 99240.58, 99029.88, 98846.99, 98698.16, 98578.19, 
    98445.62,
  99645.6, 99655.91, 99664.03, 99706.85, 99780.41, 99776.52, 99545.99, 
    93408.88, 92605.99, 99068.01, 99134.05, 98920.9, 98776.85, 98589.57, 
    98470.22,
  99367.05, 99395.67, 99432.59, 99532.59, 99660.22, 99776.72, 99761.06, 
    99602.73, 99376.04, 99406.02, 99247.44, 99054.52, 98880.36, 98682.77, 
    98510.15,
  99062.37, 99142.97, 99211.62, 99409.9, 99691.26, 99821.96, 99820.59, 
    99811.56, 99715.32, 99545.5, 99379.89, 99213.3, 99024.25, 98830.42, 
    98622.69,
  98809.99, 98885.04, 99020.38, 99397.95, 99743.43, 99890.12, 99894.65, 
    99818.32, 99715.71, 99623.27, 99478.31, 99313.38, 99147.07, 98966.62, 
    98772.2,
  98696.07, 98852.63, 99091.67, 99575.16, 99855.05, 99999.58, 99969.59, 
    99940.53, 99828.59, 99698.62, 99548.95, 99414.37, 99253.37, 99083.89, 
    98893.84,
  98833.62, 98995.58, 99263.87, 99721.43, 99954.37, 100076.8, 100045.2, 
    99949.04, 99835.95, 99715.32, 99615.77, 99495.17, 99352.02, 99208.23, 
    99043.34,
  99604.79, 99669.52, 99771.48, 99907.05, 100073.8, 100218, 100361.2, 
    100541.2, 100694.1, 100484.1, 100640, 100963.4, 100825.7, 100378.5, 
    100171.9,
  99679.02, 99723.1, 99799.55, 99933.74, 100055, 100066.2, 100354.1, 
    100446.8, 100561.8, 100721, 100771.6, 100829.5, 100832.9, 98913.57, 
    99474.18,
  99664.61, 99763.02, 99846.4, 99983.12, 99963.34, 96723.54, 100112.9, 
    100459.7, 100464.7, 100524.3, 100588.4, 100651.5, 100646.3, 100613.7, 
    100546,
  99590.88, 99703.26, 99821.65, 99937.45, 100050.2, 99906.94, 96405.45, 
    99950.85, 100370.4, 100487.4, 100518.6, 100501.8, 100527.2, 100490.7, 
    100425.2,
  99487.64, 99625.45, 99737.3, 99855.75, 99954.07, 100015.8, 99897.9, 
    94136.86, 93465.88, 100170.7, 100526.3, 100437.1, 100455, 100355.4, 
    100331.7,
  99450.9, 99600.1, 99737.16, 99905.05, 100016.8, 100104.8, 100278.9, 
    100247.1, 100280.4, 100567.5, 100500.2, 100425.4, 100371.5, 100271.9, 
    100211.1,
  99709.87, 99888.94, 100072, 100259.3, 100409.8, 100511.3, 100587.8, 
    100693.8, 100630.8, 100491.8, 100436.4, 100361.3, 100277, 100202.3, 100098,
  100068.1, 100209.5, 100324.9, 100486.9, 100582.7, 100678.9, 100670.3, 
    100608.9, 100555.1, 100520, 100406.4, 100296.4, 100211.5, 100118.1, 
    100004.5,
  100474, 100594.6, 100691.8, 100814.5, 100885.7, 100866.4, 100811.3, 
    100749.6, 100608.9, 100436.3, 100295.4, 100183.4, 100068.4, 99983.34, 
    99885.11,
  100805.4, 100861.8, 100927.5, 100964.4, 100922.8, 100878.7, 100778.8, 
    100599.3, 100432.4, 100255.5, 100117.1, 99975.63, 99860.24, 99800.84, 
    99733.23,
  99173.34, 98975.45, 98718.85, 98462.74, 98324.17, 98393.62, 98588.52, 
    98821.27, 99100.14, 99065.85, 99433.98, 99972.32, 100103.9, 100018.8, 
    100145.7,
  99425.1, 99250.73, 99045.34, 98905.49, 98762.72, 98658.5, 98901.53, 
    99065.88, 99279.55, 99557.53, 99811.03, 100103.5, 100356.6, 98778.18, 
    99650.55,
  99647.46, 99544.47, 99420.17, 99354.98, 99096.95, 95879.43, 99275.27, 
    99506.33, 99621.23, 99791.9, 100011.3, 100249, 100479.2, 100662.3, 
    100869.2,
  99825.1, 99763.27, 99747.46, 99695.2, 99740.02, 99402.09, 96017.16, 
    99635.36, 100004, 100142.6, 100323.4, 100471.3, 100701.2, 100878.5, 
    101027.4,
  99960.44, 99966.95, 99984.84, 99986.49, 99979.23, 100033.8, 99785.63, 
    94044.05, 93586.66, 100269.6, 100637.4, 100726, 100900.4, 101007.6, 
    101171.6,
  100208.3, 100212.6, 100251.8, 100297.2, 100269.2, 100233.6, 100285.6, 
    100189.9, 100235.9, 100672.7, 100782.7, 100882.7, 101004.5, 101093.1, 
    101206.7,
  100383, 100432.7, 100479.3, 100533.6, 100562.5, 100586.6, 100570.7, 
    100703.1, 100780.4, 100757.6, 100823.8, 100895.5, 100944.9, 101004.3, 
    101072.3,
  100388.9, 100438.9, 100473.4, 100530.8, 100564, 100613.2, 100626.3, 
    100591.1, 100600.7, 100674.7, 100700.5, 100706.3, 100727.4, 100748.8, 
    100810.2,
  100309.9, 100356.7, 100396.6, 100439.8, 100515.3, 100549.9, 100550, 100575, 
    100548.4, 100469.3, 100405.9, 100365, 100338.5, 100343, 100408.4,
  100138.4, 100144.5, 100164.9, 100235.2, 100267.5, 100279.7, 100262.5, 
    100199.2, 100116.4, 100040.5, 100002.3, 99941.75, 99901.84, 99912.72, 
    99980.91,
  99628.99, 99280.81, 98792.82, 98169.91, 97688.3, 97585.23, 97618.05, 
    97756.98, 97953.55, 97916.98, 98292.29, 98869.37, 99022.64, 98907.68, 
    99003.14,
  99658.59, 99338.11, 98903.89, 98404.97, 97862.47, 97449.17, 97606.41, 
    97731.09, 97926.77, 98267.2, 98586.37, 98954.81, 99219.62, 97706.02, 
    98583.61,
  99685.2, 99442.78, 99095.33, 98692.53, 98036.1, 94509.45, 97642.54, 
    97868.02, 98114.55, 98361.47, 98666.88, 98987.8, 99302.75, 99522.92, 
    99773.42,
  99699.66, 99524.8, 99282.97, 98947.37, 98594.66, 97904.73, 94396.41, 
    97827.02, 98187.62, 98438.17, 98743.39, 99014, 99332.12, 99625.31, 99901.6,
  99702.46, 99634.4, 99470.4, 99239.68, 98890.6, 98617.48, 98051.92, 
    92445.16, 92058.91, 98419.14, 98870.19, 99076.34, 99384.73, 99628.44, 
    99978.96,
  99603.48, 99597.41, 99526.23, 99458.88, 99254.47, 98992.16, 98843.98, 
    98566.48, 98422.28, 98830.09, 98995.38, 99215.75, 99487.02, 99767.95, 
    100102,
  99486.68, 99542.46, 99545.45, 99533.73, 99483.69, 99367.37, 99207.56, 
    99204.32, 99163.43, 99125.53, 99229.19, 99422.38, 99644.23, 99922.01, 
    100238.8,
  99254.53, 99294.92, 99316.93, 99395.7, 99481.91, 99548.98, 99504.42, 
    99384.08, 99317.62, 99398.98, 99496.34, 99649.52, 99865.72, 100137.5, 
    100457.9,
  99041.54, 99083.34, 99122.25, 99197.07, 99321.8, 99485.05, 99603.37, 
    99709.05, 99740.48, 99715.3, 99763.23, 99896.24, 100092.7, 100352.4, 
    100643,
  98761.51, 98749.85, 98762.46, 98849.41, 98982.41, 99245.55, 99490.27, 
    99627.16, 99711.61, 99790.62, 99933.72, 100085.5, 100284.8, 100541.1, 
    100786.9,
  99749.81, 99709.17, 99638.67, 99439.08, 99177.74, 98826.91, 98666.93, 
    98701.38, 98791.39, 98528.92, 98686.41, 99068.88, 99068.83, 98811.47, 
    98764.91,
  99609.87, 99564.35, 99506.28, 99309.78, 99052.8, 98492.97, 98664.09, 
    98698.77, 98740.72, 98823.66, 98962.48, 99139.53, 99254.06, 97565.2, 
    98316.09,
  99412.02, 99407.96, 99388.47, 99258.62, 98907.69, 95276.77, 98456.09, 
    98730.18, 98789.87, 98893.52, 99033.19, 99192.8, 99336.95, 99440.46, 
    99518.62,
  99269.59, 99264.38, 99278.27, 99185.44, 99037.35, 98545.91, 94879.89, 
    98504.04, 98766.79, 98938.59, 99119.02, 99246.2, 99391.34, 99552.8, 
    99656.8,
  99164.68, 99146.68, 99202.38, 99169.2, 99077.38, 98839.12, 98461.37, 
    92859.91, 92421.44, 98842.75, 99206.55, 99314.23, 99481.83, 99596.32, 
    99770.85,
  99142.52, 99090.25, 99109.05, 99116.62, 99079.93, 98932.78, 98719.12, 
    98725.28, 98663.41, 99119.7, 99246.48, 99418.25, 99568.5, 99728.12, 
    99889.33,
  99151.55, 99080.72, 99053.5, 99093.8, 99091.79, 99059.81, 98870.91, 
    98896.65, 99071.26, 99206.84, 99334.5, 99521.81, 99669.98, 99856.2, 100058,
  99219.38, 99098.79, 98994.23, 98977.18, 99000.95, 99105.88, 99029.88, 
    98964.46, 99044.45, 99234.55, 99421.59, 99607.04, 99798.22, 100021.3, 
    100270.9,
  99354.97, 99194.66, 99025.1, 98935.98, 98947.66, 99087.47, 99120.97, 
    99152.64, 99230.41, 99331.6, 99483.36, 99682.39, 99907.9, 100166.3, 
    100439.7,
  99598.9, 99409.62, 99162.64, 98938.77, 98861.4, 99033.36, 99175.59, 
    99205.68, 99247.16, 99322.61, 99514.39, 99729.41, 99983.98, 100284.2, 
    100570.7,
  100239.9, 100064.4, 99898.19, 99760.26, 99619.79, 99532.1, 99438.38, 
    99425.12, 99457.43, 99149.86, 99225.01, 99503.94, 99417.86, 99140.75, 
    99147.92,
  100267.4, 100040.1, 99858.73, 99714.73, 99575.52, 99327.98, 99464.23, 
    99446.73, 99479.52, 99473.55, 99491.45, 99547.02, 99613.12, 97902.93, 
    98697.06,
  100306.2, 100039, 99830.62, 99709.47, 99457.76, 96011, 99288.86, 99527.98, 
    99494.55, 99488.72, 99521.34, 99580.91, 99693.44, 99805.52, 99931.07,
  100363.3, 100086, 99817.1, 99681.35, 99544.43, 99271.75, 95625.64, 
    99222.24, 99464.4, 99477.21, 99566.45, 99640.61, 99765.32, 99932.27, 
    100069.9,
  100389.6, 100166.5, 99873.86, 99677.97, 99529.3, 99437.57, 99225.75, 
    93439.75, 92801.37, 99300.2, 99616.86, 99713.68, 99855.05, 99987.67, 
    100181.8,
  100440.5, 100210.5, 99902.73, 99675.09, 99470.51, 99381.84, 99264.04, 
    99279.24, 99187, 99497.64, 99637.68, 99793.41, 99942.2, 100098.8, 100273.2,
  100472.1, 100261, 99954.3, 99700.19, 99466.27, 99347.32, 99258.48, 
    99331.34, 99420.27, 99533.88, 99689.66, 99869.39, 100021.5, 100203.9, 
    100508.7,
  100541.6, 100324.7, 99991.12, 99703.99, 99363.73, 99285.79, 99269.56, 
    99337.61, 99420.31, 99574.92, 99761.78, 99955.52, 100157.9, 100490, 
    100824.9,
  100618.1, 100414.2, 100113.6, 99834.21, 99428.6, 99310.9, 99301.18, 
    99410.68, 99520.72, 99676.33, 99862.97, 100088.9, 100397.4, 100756.8, 
    101060.3,
  100724.4, 100529.7, 100233.5, 99903.95, 99448.98, 99347.18, 99373.87, 
    99469.47, 99579.84, 99732.62, 99972.5, 100275.3, 100622.2, 100966.5, 
    101249.4,
  100733.2, 100595.3, 100434.8, 100289.3, 100081.2, 99834.8, 99755.99, 
    99699.46, 99569.23, 99094.99, 98994.99, 99070.63, 98776.02, 98227.48, 
    97982.35,
  100762.2, 100573.6, 100414.6, 100289.9, 100086.8, 99663.1, 99812.2, 
    99712.12, 99554.48, 99471.88, 99339.23, 99267.66, 99146.18, 97254.51, 
    97868.75,
  100808.6, 100573.2, 100411.1, 100330.5, 100003.7, 96432.97, 99636.4, 
    99838.62, 99692.72, 99556.56, 99468.72, 99430.99, 99416.2, 99410.31, 
    99390.1,
  100883.8, 100619.4, 100418, 100317.8, 100195.8, 99777.41, 96048.68, 
    99549.76, 99689.37, 99662.89, 99630.12, 99614.56, 99657.75, 99734.63, 
    99784.63,
  100977.3, 100738, 100504.9, 100370.2, 100218.8, 100087.8, 99768.13, 
    93815.21, 93188.87, 99624.8, 99834.2, 99827.45, 99927.88, 99991.83, 
    100164.2,
  101095.5, 100852.6, 100600, 100423, 100254.7, 100144.4, 100043.2, 99950.71, 
    99794.55, 100005.1, 100055.7, 100108.3, 100231.8, 100345.2, 100508.8,
  101213.2, 101026.5, 100763.9, 100538.5, 100364.1, 100291.3, 100201.5, 
    100220.6, 100254.6, 100265.6, 100317.9, 100422.9, 100554.1, 100709.1, 
    100864.2,
  101355.7, 101192.4, 100965.2, 100713.3, 100474.9, 100422.8, 100387.9, 
    100395.6, 100426.8, 100513.5, 100620.2, 100764.2, 100936.2, 101095.4, 
    101227.4,
  101495, 101384.2, 101190.1, 100991.8, 100708.1, 100592.7, 100573.2, 
    100635.5, 100710, 100806.2, 100929.1, 101089.7, 101248.5, 101381.9, 
    101489.7,
  101640.7, 101537.2, 101368.6, 101196.9, 100917.6, 100724.1, 100708.8, 
    100768.7, 100857.5, 100980.9, 101185.1, 101367.3, 101524.3, 101657.6, 
    101734.5,
  101889.1, 101750.5, 101578.8, 101345.3, 101168.2, 101036.1, 100844.5, 
    100672.8, 100479.7, 99918.52, 99758.91, 99748.3, 99376.19, 98806.06, 
    98591.52,
  101941.8, 101791.9, 101644.1, 101455, 101255.2, 100893.3, 101032.3, 
    100778.7, 100577.3, 100421.2, 100191.8, 99963.15, 99641.3, 97624.3, 
    98173.98,
  101972.8, 101835.3, 101720.1, 101607.6, 101226, 97703.26, 100950.9, 
    101113.9, 100901.6, 100689.9, 100457.2, 100250.6, 100007.9, 99798.18, 
    99606.74,
  101998.7, 101869.1, 101773.8, 101680, 101558.4, 101105.5, 97365.34, 
    100863.5, 100941.2, 100922.6, 100766.4, 100561.1, 100391.7, 100214.4, 
    100049.1,
  101998.4, 101921.5, 101839.4, 101777.2, 101665.9, 101547.1, 101189.7, 
    95035.88, 94411.24, 100940.2, 101078.6, 100885.8, 100775.2, 100600.3, 
    100537.5,
  101980.9, 101923.3, 101831.9, 101801.6, 101731.7, 101643.4, 101573.2, 
    101407.6, 101173.3, 101336.7, 101282.6, 101165.6, 101076.2, 100956.2, 
    100872.1,
  101937.5, 101947.4, 101845.4, 101796, 101775.1, 101759, 101661.6, 101657.5, 
    101624.4, 101538.2, 101461.4, 101395.9, 101303.2, 101221.5, 101129.2,
  101883.7, 101896.4, 101849.9, 101773.6, 101696.9, 101751.6, 101746.5, 
    101701.1, 101653.9, 101648.4, 101608.7, 101544.8, 101476.2, 101397.1, 
    101310.1,
  101807.1, 101856.8, 101833.3, 101802.3, 101708.1, 101678.7, 101713.7, 
    101752.5, 101775.1, 101747.4, 101703, 101651.1, 101586.4, 101510.8, 
    101411.6,
  101734.4, 101751.2, 101734.5, 101717.4, 101627.2, 101567.4, 101623.2, 
    101642.5, 101672.4, 101674.7, 101716.5, 101708, 101659.9, 101597.8, 
    101489.3,
  102163.1, 102092.1, 102009.6, 101894.9, 101801, 101709.4, 101543.6, 
    101457.4, 101331.4, 100806.9, 100702.3, 100765, 100428.7, 99858.77, 
    99620.54,
  102018.9, 101920.5, 101818.8, 101714.5, 101592.9, 101254.8, 101428, 101185, 
    101046.2, 101026.1, 100904.6, 100815.7, 100624.6, 98611.18, 99161.39,
  101883, 101770, 101656.9, 101581.7, 101329.2, 97838.8, 100905.3, 101286.4, 
    101036.2, 100883.4, 100803.8, 100780.5, 100692.4, 100591.3, 100471,
  101766.8, 101626.1, 101494, 101386, 101297.5, 100947.8, 97207.39, 100423, 
    100718.6, 100762.8, 100709, 100683.6, 100713.7, 100669.7, 100602.2,
  101662.7, 101525.5, 101384.2, 101254.2, 101173, 101023.4, 100738.6, 
    94658.74, 93736.16, 100209.3, 100565.7, 100526, 100667.5, 100669.3, 
    100723.6,
  101582.6, 101422.6, 101252, 101114.2, 100945.9, 100827.9, 100674.6, 
    100380.9, 100107.9, 100289.8, 100300.5, 100356.5, 100538.5, 100651.5, 
    100734.2,
  101527.7, 101366, 101201.6, 101025.1, 100869.7, 100651.6, 100423.4, 100243, 
    100072, 99948.88, 100001.1, 100146.8, 100368.2, 100566.4, 100691,
  101520.7, 101328.1, 101149.3, 100957.9, 100728.9, 100478.4, 100175.8, 
    99820.48, 99631.16, 99628.61, 99734.02, 99922.55, 100212.8, 100460.8, 
    100631.2,
  101540, 101373.6, 101207.7, 100987.1, 100766.1, 100416.4, 100022.2, 
    99638.88, 99414.4, 99348.87, 99480.64, 99759.73, 100086.6, 100361.3, 
    100541.8,
  101591.4, 101391.4, 101220.1, 100999.7, 100728.1, 100353.5, 99926.03, 
    99416.66, 99148.18, 99119.88, 99344.82, 99685.03, 100015.9, 100288.3, 
    100457,
  101657, 101472.5, 101274.5, 101022, 100782.8, 100494.4, 100163.6, 99906.59, 
    99683.83, 99105.18, 99037.57, 99274.81, 99146.79, 98818.51, 98821.62,
  101724.7, 101520.8, 101325.5, 101090.1, 100792.3, 100192.5, 100235.1, 
    99741.81, 99397.54, 99257.63, 99129.38, 99128.84, 99142.38, 97362.22, 
    98155.25,
  101786.9, 101587.3, 101395.7, 101218, 100712.6, 97031.34, 99821.85, 
    99987.37, 99552.23, 99232.87, 99047.67, 99017.08, 99005.9, 99097.33, 
    99263.02,
  101850.6, 101651, 101492, 101265.7, 100996.4, 100324.3, 96374.01, 99285.25, 
    99239.05, 99164.4, 99037.41, 98934.17, 98912.55, 99065.58, 99294.47,
  101917.6, 101756.8, 101618.9, 101390.5, 101109.1, 100734.4, 100084.3, 
    93727.1, 92784.12, 98941.44, 99112.43, 98939.63, 98942.84, 99094.54, 
    99406.36,
  101959.9, 101824.6, 101681.3, 101491.7, 101171.1, 100808.1, 100425.9, 
    99885.48, 99356.2, 99307.59, 99219.16, 99109.55, 99142.59, 99322.4, 
    99541.03,
  101991.7, 101911.7, 101785.8, 101603, 101358.3, 100982.9, 100530.2, 
    100164.3, 99817.88, 99513.64, 99412.6, 99358.41, 99401.88, 99575.44, 
    99727.7,
  101994, 101926.6, 101833.4, 101687.9, 101422.4, 101114.2, 100744.8, 
    100320.7, 99981.18, 99775.76, 99669.03, 99634.48, 99706.01, 99846.89, 
    99966.73,
  101979.9, 101956.1, 101901.1, 101801.9, 101601.5, 101285.5, 100939, 
    100634.2, 100356.4, 100104.3, 99957.28, 99926.01, 99973.6, 100063.7, 
    100130.6,
  101942, 101894.5, 101836.1, 101737.7, 101565.2, 101362, 101121.3, 100805.5, 
    100559.7, 100365.7, 100282.3, 100223.6, 100219.2, 100245, 100253.9,
  102326.8, 102224.4, 102110.1, 101919.7, 101756.7, 101567.4, 101324, 101141, 
    100941.5, 100331.8, 100201.1, 100309.1, 100058.6, 99508.04, 99277.77,
  102219.1, 102105.2, 101989.6, 101843.8, 101665.7, 101215, 101356.6, 
    101021.1, 100811.2, 100701.8, 100512.5, 100358.8, 100184.6, 98168.05, 
    98725.2,
  102063.1, 101950.1, 101820.8, 101740.9, 101414.3, 97921.68, 100944.6, 
    101262.3, 101030.4, 100768.8, 100560.5, 100406.6, 100227.2, 100091.2, 
    99929.68,
  101900.9, 101772, 101640.1, 101523.1, 101422.7, 101052.5, 97336.37, 
    100560.7, 100694.1, 100773.2, 100631.4, 100454.9, 100309, 100159.8, 
    100033.8,
  101706.8, 101584.9, 101452.2, 101331.6, 101225.9, 101134.9, 100867.2, 
    94849.33, 94044.93, 100404.6, 100668.8, 100496, 100418.2, 100240.3, 
    100162.7,
  101499.8, 101362.2, 101198.3, 101097.8, 100966.4, 100876.5, 100824.5, 
    100645.5, 100408.3, 100604.9, 100572.4, 100504.3, 100457.8, 100352.6, 
    100263.1,
  101275.1, 101131.6, 100964.1, 100847.1, 100743.5, 100648.1, 100542.9, 
    100539, 100512.9, 100431.1, 100423.6, 100457.2, 100438.9, 100400.6, 100331,
  101052.9, 100872.7, 100687.9, 100571.2, 100428.4, 100334.5, 100253.4, 
    100150.3, 100101.6, 100158.4, 100254.2, 100335.7, 100382.5, 100380.4, 
    100340.1,
  100831.6, 100644.8, 100465, 100315.6, 100183.2, 100062.4, 99959.11, 
    99922.22, 99912.92, 99921.45, 100029.3, 100199.1, 100297.7, 100327.2, 
    100298.3,
  100620.2, 100390, 100196.4, 100043.2, 99881.65, 99752.86, 99657.94, 
    99566.17, 99531.73, 99598.3, 99833.2, 100067.9, 100201.3, 100256.2, 
    100225.6,
  101018.9, 100754.7, 100509.8, 100285.5, 100156.8, 100066, 99984.39, 
    99975.69, 100017.5, 99763.44, 99913.73, 100267.6, 100217, 99882.55, 
    99782.63,
  100937.5, 100633.7, 100377.3, 100130.4, 99963.35, 99665.53, 99807.94, 
    99670.88, 99650.79, 99741.48, 99852.88, 100003.2, 100134.2, 98377.96, 
    99063.98,
  100864.2, 100564.9, 100297.5, 100069.7, 99748.23, 96372.34, 99425.54, 
    99613.94, 99500.84, 99479.61, 99533.98, 99682.08, 99845.37, 99977.53, 
    100078.8,
  100814.2, 100517.8, 100249.7, 100004.8, 99819.09, 99465.83, 95854.77, 
    99064.92, 99246.73, 99264.59, 99279.29, 99363.82, 99552.49, 99765.24, 
    99942.08,
  100786.2, 100509.7, 100245.6, 100008.8, 99820.76, 99653.97, 99341.14, 
    93524.52, 92732.95, 98838.71, 99047.31, 99053.6, 99233.66, 99465.58, 
    99756.18,
  100770.5, 100502.8, 100244.5, 100031.2, 99805.71, 99647.74, 99465.11, 
    99233.49, 98942.67, 98963.41, 98830.91, 98805.58, 98965.77, 99238.12, 
    99596.93,
  100769.6, 100533.3, 100293.1, 100095.2, 99899.88, 99695.84, 99481.64, 
    99305.39, 99081.16, 98827.99, 98654.52, 98601.86, 98755.21, 99108.8, 
    99528.49,
  100793.9, 100561.2, 100341.9, 100168, 99952.86, 99762.96, 99531.97, 
    99294.91, 99058.62, 98842.13, 98607.13, 98530.6, 98771.86, 99223.94, 
    99602.98,
  100819.9, 100615.8, 100430.6, 100285.9, 100099.6, 99881.69, 99648.54, 
    99438.41, 99200.8, 98960.71, 98773.31, 98798.84, 99143.93, 99466.59, 
    99735.27,
  100829.4, 100613, 100444.1, 100326.9, 100154.1, 99974.91, 99773.97, 
    99545.69, 99341.46, 99165.05, 99113.8, 99245.86, 99472.19, 99696.32, 
    99878.84,
  101164.9, 100942.8, 100734.9, 100534.1, 100402.7, 100268, 100140.7, 
    99998.65, 99868.95, 99401.41, 99368.71, 99584.41, 99520.69, 99286.52, 
    99309.2,
  101122.8, 100877.5, 100677.1, 100492.9, 100362.9, 100025, 100190.9, 
    99933.62, 99772.8, 99705.38, 99589.89, 99523.13, 99533.22, 97825.34, 
    98559.54,
  101053.6, 100809.9, 100615.6, 100472.7, 100217.2, 96818.66, 99922.05, 
    100144.5, 99956.29, 99772.02, 99577.2, 99455.42, 99386.95, 99447.02, 
    99541.53,
  100950.4, 100714, 100529.9, 100382.5, 100311.4, 100022.6, 96369.07, 
    99679.14, 99783.12, 99797.88, 99582.39, 99370.24, 99251.58, 99264.66, 
    99378.16,
  100830.6, 100609.4, 100432.9, 100298.9, 100239.7, 100212.4, 100004.8, 
    94022.12, 93281.91, 99553.68, 99578.48, 99273.5, 99125.1, 99053.95, 
    99187.7,
  100687.9, 100461.6, 100274.1, 100165.5, 100079.9, 100074.3, 100101.8, 
    99972.66, 99755.8, 99821.41, 99563.45, 99248.85, 99016.19, 98927.27, 
    98998.06,
  100540.7, 100331.4, 100132.9, 100011.3, 99938.31, 99930.53, 99932.26, 
    100019, 100011.8, 99860.13, 99639.23, 99377.23, 99109.96, 98984.16, 
    99093.49,
  100402.4, 100167.8, 99941.62, 99810.96, 99709.89, 99724.83, 99760.26, 
    99798.61, 99827.91, 99856.28, 99780.97, 99646.14, 99528.43, 99472.82, 
    99515.12,
  100276, 100036.1, 99809.2, 99639.23, 99539.52, 99532.98, 99571.2, 99681.39, 
    99779.21, 99817.45, 99812.7, 99784.9, 99735.4, 99730.71, 99765.25,
  100146.4, 99864.02, 99618.2, 99430.02, 99306.25, 99301.17, 99361.16, 
    99415.28, 99503.05, 99603.47, 99734.13, 99808.19, 99841.64, 99880.14, 
    99896.62,
  100475.5, 100156.2, 99877.51, 99649.2, 99565.97, 99583.12, 99622.38, 
    99733.62, 99845.58, 99539.59, 99585.15, 99787.21, 99531.85, 99057.68, 
    98940.45,
  100489.2, 100125.8, 99849.9, 99611.38, 99486.87, 99309.33, 99562.84, 
    99582.66, 99673.59, 99780.01, 99786.2, 99771.79, 99682.86, 97777.17, 
    98400.09,
  100494.2, 100114.9, 99835.29, 99612.73, 99335.22, 96027.43, 99253.66, 
    99587.02, 99636.62, 99661.62, 99687.04, 99689.14, 99643.91, 99568.97, 
    99518.39,
  100484.1, 100107.8, 99817.4, 99583.98, 99427.27, 99144.46, 95618.81, 
    99091.96, 99440.06, 99537.48, 99578.82, 99561.15, 99543.93, 99484.67, 
    99475.74,
  100480.1, 100117.3, 99833.98, 99599.9, 99427.42, 99301.91, 99113.7, 
    93426.14, 92742.66, 99039.34, 99404.74, 99396.18, 99422.93, 99356.65, 
    99374.68,
  100476.1, 100107.3, 99819.47, 99607.77, 99405.75, 99271.2, 99172.45, 
    99080.19, 98964.21, 99189.22, 99238.46, 99272.77, 99314.59, 99276, 
    99248.76,
  100464.8, 100123, 99835.59, 99645.06, 99460.43, 99288.59, 99138.96, 
    99075.97, 99036.9, 99025.8, 99087.32, 99157.66, 99204.11, 99190.95, 99139,
  100439.5, 100100.2, 99815.25, 99667.88, 99484.36, 99319.91, 99148.48, 
    99010.55, 98936.35, 98949.51, 98989.04, 99041.59, 99097.38, 99155.92, 
    99146.55,
  100406.8, 100092.8, 99852.13, 99736.26, 99593.95, 99415.11, 99238.45, 
    99108.7, 98985.98, 98906.85, 98893.38, 98913.41, 98956.75, 99041.71, 
    99117.84,
  100353.6, 100031.6, 99820.07, 99743.3, 99648.55, 99504.57, 99348.91, 
    99171.45, 99029.67, 98902.6, 98847.23, 98812.14, 98818.74, 98911.5, 
    99031.14,
  100815, 100516.5, 100256.7, 100045.2, 99865.19, 99687.63, 99523.85, 
    99419.33, 99402.66, 99124.03, 99275.55, 99591.68, 99460, 99043.52, 
    98850.77,
  100833.6, 100507.9, 100271, 100089.5, 99905.95, 99486.11, 99580.57, 
    99323.32, 99275.43, 99323.7, 99398.06, 99503.23, 99571.48, 97736.17, 
    98340.09,
  100838.1, 100522, 100298.2, 100170.5, 99862.41, 96346.3, 99393.7, 99491.86, 
    99343.54, 99294.42, 99285.2, 99352.54, 99429.91, 99519.83, 99494.84,
  100823.7, 100544, 100331.4, 100215, 100107.7, 99701.76, 95924.55, 99176.17, 
    99356.84, 99357.62, 99260.58, 99211.17, 99253.12, 99373.69, 99456.99,
  100820.3, 100589, 100394, 100308.5, 100216.7, 100066.5, 99701.66, 93634.68, 
    92864.22, 99164.31, 99282.02, 99117.09, 99073.95, 99101.7, 99283.37,
  100817.6, 100615.8, 100444.2, 100392.5, 100289, 100189.6, 100002.2, 
    99796.11, 99526.34, 99541.98, 99362.16, 99185.2, 99061.81, 98981.91, 
    99071.02,
  100823.1, 100680.9, 100542.8, 100518.1, 100461.9, 100321.7, 100156.5, 
    100029, 99856.5, 99653.55, 99477.78, 99296.24, 99102.77, 98982.73, 98915.4,
  100846.6, 100742, 100640.8, 100652.1, 100552.1, 100453.2, 100273.1, 
    100097.6, 99934.31, 99799.69, 99628.89, 99423.47, 99210.34, 99007.72, 
    98885.8,
  100914.5, 100847.1, 100820.3, 100846.1, 100760, 100602.4, 100416.5, 
    100256.7, 100074.7, 99881.96, 99712.84, 99529.15, 99312.18, 99079.13, 
    98888.15,
  101010.2, 100937.2, 100927.1, 100935.8, 100824.9, 100705.7, 100522.7, 
    100301, 100104.8, 99918.98, 99778.77, 99604.08, 99384.16, 99165.95, 
    98927.91,
  101161.4, 101084.7, 100946.8, 100747.1, 100582.1, 100436.4, 100250.5, 
    100078, 99880.43, 99271.27, 99110.43, 99179.99, 98938.35, 98574.35, 
    98456.34,
  101225.4, 101110.9, 101011.5, 100850.6, 100675.7, 100308.1, 100446.4, 
    100153.5, 99971.92, 99824.39, 99561.51, 99346.99, 99173.44, 97298.11, 
    97923.45,
  101248.1, 101124.7, 101024.7, 100962.9, 100619.8, 97048.16, 100267.4, 
    100481.4, 100226.6, 100010, 99761.61, 99540.4, 99291.65, 99184.25, 
    99073.59,
  101273.7, 101145.2, 101035.5, 100966.3, 100850.9, 100469.9, 96615.33, 
    100003.1, 100111.7, 100100, 99908.81, 99675.12, 99445.84, 99246.95, 
    99132.95,
  101280.1, 101160.9, 101044.1, 100960.9, 100841.7, 100742.8, 100431, 
    94177.78, 93333.22, 99868.52, 100003, 99763.05, 99581.7, 99294.16, 
    99156.06,
  101282.5, 101144.2, 101004.7, 100922.8, 100776.3, 100692.1, 100550.5, 
    100312.4, 100036.8, 100104.6, 99976.52, 99802.56, 99625.59, 99418.19, 
    99179.38,
  101282.7, 101150.5, 100995.2, 100896.9, 100787.2, 100637.8, 100452.8, 
    100318.9, 100159.6, 99989.59, 99890.07, 99785.06, 99643.44, 99433.56, 
    99219.05,
  101302.5, 101140.2, 100961.8, 100868.7, 100702.4, 100541.4, 100335, 
    100117.1, 99942.94, 99855.04, 99785.55, 99720.45, 99629.32, 99459.9, 
    99262.19,
  101339.3, 101173.9, 101002.1, 100872.7, 100706.1, 100481.5, 100249.9, 
    100052.8, 99868.98, 99729.11, 99670.39, 99655.47, 99589.22, 99476.41, 
    99246.89,
  101392.3, 101174.9, 100978.4, 100807.2, 100595.3, 100385.3, 100152.4, 
    99887.36, 99689.92, 99576.47, 99571.98, 99579.91, 99549.19, 99478.59, 
    99294.3,
  100532.8, 100311.6, 100093.8, 99935.43, 99837.3, 99888.18, 100043.1, 
    100234, 100327.2, 99976.94, 99955.71, 100071.3, 99647.29, 99031.26, 
    98759.79,
  100387.9, 100114.4, 99891.88, 99733.23, 99649.9, 99568.93, 99972.3, 
    100090.9, 100182.5, 100293.2, 100255.5, 100204.8, 99986.2, 97919.91, 
    98416.81,
  100249.9, 99972.52, 99736.58, 99620.54, 99448.57, 96153.6, 99643.81, 
    100101.9, 100143, 100210.9, 100233.8, 100251.5, 100142.5, 99985.29, 
    99736.2,
  100142.9, 99890.7, 99644.52, 99546.5, 99495.04, 99345.32, 95848.87, 
    99550.61, 99986.4, 100093.9, 100184.6, 100221.5, 100224, 100106.1, 
    99942.02,
  100081.4, 99849.71, 99604.8, 99528.09, 99498.69, 99481.22, 99405.5, 
    93619.49, 92951.55, 99659.98, 100058.1, 100148.5, 100251.1, 100156.8, 
    100075.4,
  100073.5, 99839.84, 99610.98, 99523.63, 99440.41, 99470.55, 99492.55, 
    99493.78, 99476.76, 99798.38, 99913.01, 100075.5, 100220.8, 100222.4, 
    100139.5,
  100103.7, 99911.76, 99686.52, 99587.12, 99537.11, 99529.98, 99480.26, 
    99582.09, 99641.65, 99684.81, 99813.35, 100009.1, 100181.1, 100229.6, 
    100178.2,
  100184.1, 99997.3, 99781.19, 99675.5, 99510.77, 99465.66, 99462.02, 
    99466.08, 99524.43, 99637.27, 99755.18, 99949.62, 100156.3, 100238.4, 
    100203.8,
  100302.8, 100136.4, 99931.76, 99753.48, 99579.78, 99440.45, 99384.82, 
    99432.8, 99508.58, 99580.7, 99707.84, 99923.09, 100142.9, 100233.8, 
    100209.8,
  100435.8, 100257.2, 100030.1, 99806.41, 99547.79, 99381.07, 99325.55, 
    99312.88, 99411.2, 99521.43, 99721.03, 99951.33, 100158.1, 100245.8, 
    100222.6,
  100042.1, 99843.7, 99663.52, 99520.59, 99383.73, 99224.8, 99157.98, 
    99287.7, 99553.8, 99469.96, 99727.72, 100077, 99858.16, 99318.34, 99081.52,
  99983.04, 99736.91, 99534.47, 99370.73, 99172.22, 98875.58, 99052.34, 
    99217.07, 99505.92, 99831.58, 100022.5, 100131.7, 100016.4, 98015.77, 
    98593.77,
  99949.59, 99682.92, 99455.39, 99294.77, 98991.68, 95555.12, 99021.44, 
    99419.65, 99723.52, 99941.88, 100104.6, 100173.3, 100110.9, 99929.38, 
    99793.61,
  99960.95, 99709.32, 99477.59, 99334.65, 99259.23, 99022.02, 95487.15, 
    99342.36, 99815.83, 100055.8, 100193.4, 100209.5, 100147, 100009.9, 
    99913.45,
  100018.4, 99766.12, 99535.86, 99452.44, 99361.97, 99410.95, 99185.84, 
    93550.28, 93032.58, 99888.13, 100264, 100275.6, 100234.2, 100053.6, 
    100022.6,
  100134.4, 99871.83, 99627.85, 99501.23, 99417.57, 99443.57, 99499.82, 
    99542.98, 99605.16, 100146.7, 100274.1, 100348.4, 100298.4, 100173.6, 
    100094.9,
  100279.5, 100044.1, 99774.38, 99599.92, 99509.57, 99493.48, 99466.77, 
    99822.27, 100072.9, 100220.2, 100353.2, 100432.9, 100372.4, 100275.9, 
    100202.6,
  100475.8, 100284.6, 100025.8, 99807.95, 99609.9, 99612.45, 99693.69, 
    99881.83, 100090.4, 100337.4, 100467.8, 100524.1, 100482.1, 100410.8, 
    100365.6,
  100678.4, 100539.5, 100361.9, 100178.5, 100006.5, 99956.37, 100028.9, 
    100229.9, 100393.7, 100512.5, 100605.6, 100655.6, 100624.6, 100557.9, 
    100504.8,
  100888.5, 100770.5, 100607.7, 100455, 100313.9, 100285.3, 100334, 100406.1, 
    100518.2, 100623.9, 100751.6, 100805.1, 100790.4, 100729.1, 100659.1,
  100660.2, 100484.8, 100301.6, 100095.1, 99744.18, 99433.34, 99281.87, 
    99369.56, 99458.31, 99035.3, 99235.7, 99734.87, 99866.98, 99739.97, 
    99784.02,
  100636.7, 100460.3, 100299.4, 100076.8, 99683.41, 99122.26, 99201.33, 
    99271.98, 99362.91, 99404.37, 99617.53, 99899.87, 100153.4, 98512.91, 
    99321.3,
  100643, 100481.4, 100349, 100186.1, 99673.49, 95976.7, 99141.09, 99333.26, 
    99473.39, 99562.11, 99797.3, 100050.4, 100293.5, 100444.2, 100537,
  100669.1, 100543.4, 100446.5, 100293.9, 100062.9, 99558.91, 95814.96, 
    99423.2, 99618.73, 99795.65, 100011, 100180.2, 100358.2, 100489.8, 
    100598.7,
  100718.6, 100630, 100569.7, 100481.3, 100277.6, 100158, 99722.92, 93730.13, 
    93281.52, 99887.66, 100234.2, 100262.4, 100376.5, 100399.7, 100577.6,
  100808.1, 100713.7, 100666.4, 100635.1, 100492.2, 100370.2, 100332.9, 
    100159.2, 99991.84, 100302.4, 100317.3, 100321.4, 100333.3, 100376.7, 
    100512.2,
  100926.6, 100844.8, 100800.7, 100787.2, 100713.7, 100624.6, 100491.4, 
    100519.7, 100507.4, 100391, 100321.1, 100277.2, 100252.1, 100318.7, 
    100446.9,
  101093.2, 101038, 100970.7, 100945, 100866, 100790.6, 100688.2, 100543, 
    100421.1, 100378.7, 100272.8, 100204.5, 100209, 100323.6, 100457.5,
  101240.2, 101229.1, 101200.9, 101136.1, 101057.5, 100963.3, 100814.9, 
    100712.9, 100578.5, 100405.4, 100256.2, 100213.4, 100262.4, 100387.4, 
    100488.9,
  101392.4, 101389.9, 101330.2, 101285.5, 101187.9, 101096.3, 100962.6, 
    100759.2, 100580.1, 100431.7, 100381.3, 100366.2, 100408.3, 100494.7, 
    100542.2,
  101300.9, 101361.6, 101303.3, 101079.8, 100700.1, 100265.2, 99773.6, 
    99282.45, 98999.77, 98566.04, 98636.91, 98867.38, 98745.48, 98509.42, 
    98575.08,
  101313.5, 101387.3, 101308, 101111.5, 100735.8, 100102.7, 99971.18, 
    99465.13, 99135.13, 99021.12, 98947.04, 98962.75, 99007.96, 97389.71, 
    98227.61,
  101341.9, 101401.1, 101352.6, 101228.6, 100731.6, 97014.12, 100051.2, 
    99960.57, 99700.93, 99519.59, 99432.61, 99407.41, 99452.09, 99542.84, 
    99618.9,
  101417.1, 101433.6, 101422, 101280.9, 101102.6, 100512.6, 96679.07, 
    100028.6, 100021.7, 100016.7, 99942.16, 99892.66, 99909.09, 99935.16, 
    99951.54,
  101508.2, 101508.7, 101503.7, 101395.9, 101223.4, 101063.4, 100585.5, 
    94438.13, 93867.71, 100286.4, 100440, 100339.5, 100338.5, 100283.9, 
    100316.7,
  101618.7, 101591.6, 101544.9, 101474, 101312.7, 101146.7, 101074, 100863.6, 
    100597.1, 100742.4, 100706.3, 100646.4, 100631, 100604.4, 100596.5,
  101756.9, 101729.6, 101669.9, 101560.1, 101428.7, 101267.6, 101072.9, 
    101048.4, 101030.9, 100922.6, 100859.8, 100845.7, 100812.3, 100789.1, 
    100763.7,
  101897.3, 101866, 101797.9, 101677.4, 101464, 101291, 101109, 100951.6, 
    100868.1, 100893.5, 100901.7, 100895.4, 100889.3, 100885.9, 100858.7,
  102016.1, 102007, 101954.1, 101818.3, 101615.3, 101369, 101090.5, 100930.3, 
    100867.8, 100836.1, 100822.9, 100843.1, 100872.1, 100870, 100850.1,
  102124, 102113.7, 102035.5, 101913.7, 101712.6, 101488.1, 101205.8, 
    100914.4, 100736.1, 100665.7, 100698, 100738.2, 100787.3, 100827.2, 
    100839.3,
  102668.8, 102515.7, 102351.1, 102124.8, 101882.7, 101628.9, 101329.8, 
    100987.2, 100619.8, 99905.87, 99662.17, 99816.96, 99654.98, 99203.61, 
    99044.73,
  102649.4, 102491.4, 102345.9, 102166.3, 101910.3, 101432, 101442.4, 101059, 
    100712.2, 100422.3, 100057.3, 99857.95, 99896.32, 98011.88, 98688.66,
  102610.8, 102467.6, 102337.5, 102226.4, 101841.4, 98171.23, 101236.1, 
    101305.9, 100953.4, 100621.7, 100288.4, 99967.12, 99897.92, 100001.2, 
    99982.63,
  102574.5, 102448.7, 102332.1, 102209.8, 102034.9, 101569, 97634.19, 
    100843.7, 100838.9, 100735.3, 100496.5, 100169.3, 99869.98, 99982.94, 
    100076.2,
  102526.8, 102438.7, 102325.3, 102207, 102036.8, 101850.5, 101432.1, 
    95149.9, 94250.5, 100615.2, 100653, 100376.5, 100119.6, 99963.55, 100100.7,
  102465.6, 102393.1, 102277.7, 102164.2, 101987.9, 101808.2, 101587.5, 
    101267.4, 100880.5, 100889, 100750.9, 100526.1, 100271.1, 100094, 100096.4,
  102388.1, 102342.4, 102228, 102131.3, 101995.3, 101792.3, 101540.3, 
    101305.6, 101049.4, 100872.6, 100766.7, 100637.4, 100433.1, 100242.1, 
    100161.5,
  102290.4, 102210.1, 102117.4, 102053.1, 101919, 101754.4, 101516.5, 
    101200.7, 100939.5, 100817.8, 100768, 100670.1, 100543.4, 100382.5, 
    100287.1,
  102113.7, 102062.9, 102018.6, 101978.9, 101909, 101747.5, 101519.9, 
    101228.4, 100971.7, 100782.4, 100732.3, 100689.6, 100599.7, 100478.8, 
    100374.4,
  101910.9, 101876.5, 101868.2, 101880, 101807.3, 101713.1, 101521.8, 101203, 
    100916, 100703.4, 100683.3, 100665.4, 100606.8, 100533.9, 100452.9,
  102480.1, 102345.6, 102218.4, 102056.2, 101929.1, 101759.6, 101527.2, 
    101354.8, 101197.4, 100596.6, 100421, 100407.8, 100094.4, 99348.5, 
    98901.69,
  102255.9, 102103, 101985.3, 101836, 101708, 101313.3, 101431.6, 101207.7, 
    101043.3, 100889.5, 100659.1, 100466.6, 100291.8, 98195.65, 98571.84,
  102036.6, 101901.5, 101778, 101675.6, 101400.3, 97917.67, 100990.3, 
    101294.5, 101112.1, 100913.1, 100677, 100492.3, 100362.2, 100252, 99967.73,
  101846.4, 101728.7, 101609.8, 101471.5, 101334.5, 100981.2, 97340.35, 
    100794.1, 100982.4, 100891.2, 100720.5, 100502.7, 100396.9, 100347.5, 
    100220,
  101690.9, 101580, 101466.5, 101322.6, 101220.7, 101110, 100994.8, 94996.91, 
    94227.94, 100676.3, 100731.9, 100520.6, 100376.7, 100319, 100318.7,
  101573.5, 101453.1, 101335, 101218.8, 101118.5, 101131.3, 101200.1, 
    101077.2, 100850.5, 100892.5, 100719.4, 100529.8, 100331.2, 100243.7, 
    100235.6,
  101482.9, 101375.5, 101279.4, 101193.9, 101169.7, 101235, 101214.4, 101159, 
    101066.2, 100838, 100707, 100549, 100324.6, 100169.4, 100082.7,
  101423.5, 101317.8, 101251.6, 101214.5, 101243, 101278.7, 101222, 101052.3, 
    100915.3, 100797.3, 100698.1, 100552.7, 100339, 100164.7, 100012,
  101374.1, 101328, 101299.9, 101331.3, 101372.9, 101347.3, 101238.4, 
    101073.9, 100908.7, 100774.7, 100688.3, 100563.2, 100359.5, 100175.4, 
    100022.8,
  101361.6, 101340.3, 101338.8, 101366.5, 101379.6, 101375.3, 101253.5, 
    101020.6, 100824.4, 100709.7, 100680.9, 100565.7, 100378.3, 100202.6, 
    100074.9,
  101715.8, 101619.2, 101509.1, 101361, 101229.3, 101097.3, 100981.3, 
    100921.2, 100963, 100677.7, 100749.2, 100915.4, 100616.6, 99981.49, 
    99588.8,
  101673.1, 101559, 101467.2, 101343.3, 101223.4, 100884.1, 101042.7, 
    100899.3, 100913.4, 100998.3, 100955.5, 100883.4, 100694.1, 98639.79, 
    99058.79,
  101651.6, 101572.4, 101489.9, 101429.9, 101161.2, 97668.13, 100882, 
    101154.8, 101067.3, 101014, 100908.6, 100813.4, 100620, 100427, 100175.5,
  101650, 101599, 101537.7, 101506.8, 101422.4, 101084.8, 97317.83, 100780.2, 
    100976.4, 100995.2, 100867.7, 100724.8, 100532.1, 100334, 100111.7,
  101646.3, 101646.5, 101612.6, 101592.9, 101537.1, 101451.5, 101117.4, 
    94991.81, 94181.02, 100684.3, 100817.5, 100631.4, 100434, 100199.5, 
    100013.9,
  101624.7, 101644.6, 101611.2, 101609.4, 101521.1, 101460.7, 101338.2, 
    101089.9, 100808.8, 100882.5, 100719.4, 100540, 100324.9, 100086.8, 
    99905.42,
  101580, 101603, 101564.3, 101585.2, 101556.8, 101471.2, 101325.6, 101175.2, 
    100973.1, 100766.7, 100613.3, 100440, 100208.9, 99978.69, 99823.97,
  101535.3, 101511.2, 101455.3, 101481.1, 101471.2, 101459.3, 101314.6, 
    101071.4, 100846.9, 100709, 100543.1, 100351.7, 100122.5, 99927.75, 
    99820.34,
  101490.2, 101450.4, 101395.6, 101393.3, 101443.8, 101468, 101333.5, 
    101124.6, 100873.4, 100671.4, 100483, 100293.3, 100083.3, 99945.7, 
    99863.92,
  101459.9, 101379.2, 101310.8, 101283.2, 101365.8, 101460.2, 101342.9, 
    101075.7, 100824.8, 100621.2, 100467.1, 100301.1, 100135.1, 100045.2, 
    99980.63,
  101954.4, 101947.6, 101882.8, 101761.1, 101650.9, 101560.1, 101430.3, 
    101331.4, 101196.3, 100694.1, 100640.5, 100817.7, 100597.3, 100131.8, 
    99926.66,
  101936.7, 101882.1, 101805.4, 101683.6, 101557.3, 101254.4, 101450.6, 
    101212.8, 101039.5, 100968.1, 100843.5, 100774, 100675, 98721.66, 99259.05,
  101851.7, 101783.7, 101684.6, 101598.8, 101324.5, 97896.49, 101133.4, 
    101389.3, 101151.9, 100929, 100731.4, 100636.1, 100496.1, 100401.5, 
    100243.7,
  101737.4, 101668, 101565.6, 101448.1, 101369.6, 101151.6, 97483.35, 
    100824.8, 100895.8, 100840.9, 100629.3, 100466.5, 100300.4, 100153.3, 
    99967.55,
  101648.2, 101582.9, 101487.9, 101341, 101301.2, 101352.4, 101174.8, 
    95058.34, 94222.48, 100505, 100547.4, 100312.6, 100124.4, 99914.4, 
    99756.49,
  101583.6, 101520.5, 101412.6, 101273.1, 101266.1, 101337.3, 101332.5, 
    101098.5, 100733.8, 100689.3, 100455.5, 100209.4, 99968.98, 99723.79, 
    99524.2,
  101546.2, 101513, 101422.4, 101288.5, 101342.9, 101384.7, 101294.1, 
    101153.8, 100919.7, 100657.2, 100411.5, 100132.8, 99816.02, 99523.97, 
    99251.69,
  101527.8, 101515.2, 101454.9, 101347.7, 101389.1, 101419.2, 101297.3, 
    101069.4, 100870, 100697, 100443, 100129.7, 99767.49, 99411.98, 99061.11,
  101513.2, 101544.2, 101545.8, 101480.7, 101544.5, 101486, 101331.7, 
    101150.6, 100992.4, 100794.7, 100557.7, 100244.6, 99859.65, 99467.01, 
    99093.58,
  101506, 101536.4, 101565, 101558.2, 101610.7, 101520.8, 101368.1, 101162.7, 
    101033.6, 100887.6, 100724.6, 100446.6, 100084.4, 99714.72, 99339.08,
  101929.5, 101920.3, 101879.2, 101793.6, 101719, 101658.5, 101607.9, 
    101581.5, 101492.2, 100980.5, 100868.1, 100961.1, 100687.2, 100179.3, 
    99986.33,
  101919.8, 101912.5, 101889.5, 101816.4, 101731.4, 101476.8, 101696.4, 
    101485.1, 101307.1, 101189.1, 101014.2, 100858.7, 100694, 98729.49, 
    99323.62,
  101927.9, 101952, 101936.5, 101918.2, 101673, 98258.18, 101509.5, 101681.8, 
    101460.2, 101201.3, 100926.6, 100742.4, 100535.1, 100418.1, 100319,
  101934.8, 101984.2, 101995.4, 101975, 101945.4, 101631.9, 97886.84, 
    101238.7, 101188.8, 101144.8, 100874.2, 100612.3, 100380.9, 100215.2, 
    100128.7,
  101952, 102014.2, 102047.6, 102054, 102055.5, 101972.1, 101673.3, 95500.23, 
    94702.64, 100886.2, 100843.9, 100473.3, 100199.6, 99942.75, 99886.34,
  101932.8, 102033.3, 102067.6, 102108.9, 102073.1, 101997.4, 101902.7, 
    101660.2, 101281.6, 101152.7, 100806.7, 100405.8, 100051.7, 99743.14, 
    99577.85,
  101894.7, 102046.9, 102094.8, 102144.2, 102141.4, 102049.2, 101912.3, 
    101792.5, 101552, 101185.3, 100805, 100408.4, 100000.7, 99649.16, 99395.49,
  101874.2, 102041.1, 102095.9, 102161.5, 102127.5, 102065.9, 101956.7, 
    101767.9, 101509.5, 101224.7, 100875.8, 100474.5, 100052.2, 99661.1, 
    99351.98,
  101823.4, 101998.2, 102107.5, 102166.4, 102170, 102085.6, 101983.8, 
    101858.5, 101636.2, 101317.7, 100970.5, 100575.2, 100134.4, 99716.09, 
    99355.65,
  101774.1, 101910.6, 102046.3, 102101.5, 102109.1, 102061.2, 101982.9, 
    101835.4, 101629.7, 101350.3, 101063.7, 100694.9, 100246.9, 99806.58, 
    99410.66,
  102885.8, 102894, 102884.5, 102897.7, 102890.1, 102825.7, 102727.7, 
    102652.4, 102515.6, 101989.8, 101863.2, 101928.4, 101565.2, 100915, 
    100622.5,
  102888.4, 102890.2, 102891, 102880.4, 102849.1, 102604.7, 102739.8, 
    102530.4, 102370.2, 102277.9, 102104, 101937.2, 101700.5, 99602.21, 
    100059.2,
  102790.5, 102820.9, 102857.8, 102878, 102687, 99184.15, 102466.2, 102686.4, 
    102498.8, 102267.6, 102058.2, 101893.5, 101664.2, 101450.4, 101180.9,
  102613.5, 102668.4, 102725.9, 102764.3, 102762.9, 102495.8, 98740.24, 
    102113.2, 102193.5, 102200.3, 102011.5, 101803.6, 101594.5, 101372.6, 
    101108.4,
  102432.5, 102514.6, 102569.5, 102621.1, 102628.6, 102623.5, 102407.1, 
    96303.18, 95462.02, 101805.5, 101938.8, 101685.8, 101487.5, 101220.3, 
    101001.7,
  102294.8, 102349, 102378.6, 102435.3, 102432.8, 102432, 102404.9, 102219.2, 
    101930.8, 101977.8, 101782.2, 101563.2, 101342.6, 101086.5, 100827.1,
  102190.4, 102223.6, 102234.6, 102258.1, 102261.3, 102242.8, 102164.8, 
    102116.4, 101980.2, 101757.2, 101570, 101398.7, 101172, 100930.9, 100627.6,
  102095, 102098.6, 102065, 102086, 102046.3, 102009.2, 101922.9, 101786.8, 
    101632.3, 101518.5, 101374.3, 101213.9, 101020.6, 100779.7, 100469.1,
  102029.9, 102013.8, 101971.6, 101927.9, 101862.1, 101780.7, 101670.4, 
    101583.1, 101465.4, 101311.4, 101175.1, 101050, 100876.8, 100629.1, 
    100315.6,
  101991.6, 101905.2, 101801, 101716.1, 101603.7, 101497.4, 101410.8, 
    101286.8, 101178, 101066.7, 101011.8, 100916.6, 100752.3, 100504.9, 
    100202.7,
  102917.3, 102837.7, 102775.4, 102710.2, 102713.8, 102725.9, 102707.6, 
    102710, 102665.6, 102200.4, 102156.6, 102322.5, 102107.6, 101577.5, 
    101342.3,
  102672.1, 102573.4, 102528.6, 102492.8, 102505.8, 102329.9, 102566.8, 
    102444.8, 102352.5, 102320.5, 102232.3, 102191.3, 102151.7, 100204.6, 
    100783.2,
  102444.7, 102358.6, 102330, 102322.8, 102262.8, 98909.93, 102114.6, 
    102424.1, 102276.3, 102125.9, 102013.3, 101966.9, 101931.6, 101917.4, 
    101857,
  102272.4, 102204.5, 102182.2, 102187.2, 102194.3, 102018.3, 98398.41, 
    101700.1, 101859, 101836.5, 101755.8, 101666.9, 101641.9, 101642.4, 
    101656.3,
  102161.2, 102140.1, 102126.8, 102096.6, 102091.9, 102039, 101831.1, 
    95936.28, 95084.24, 101279.8, 101482.8, 101344.3, 101315.5, 101264.6, 
    101312.6,
  102117.2, 102084, 102036.3, 102011.9, 101900.9, 101823.6, 101713.8, 
    101517.7, 101254.4, 101324.7, 101187.9, 101070.3, 100999, 100939.9, 100948,
  102040.6, 102012.8, 101954.7, 101891.2, 101795.1, 101651, 101491.8, 
    101373.9, 101237, 101069.2, 100927.9, 100805.6, 100684.7, 100611.7, 
    100583.7,
  101940.1, 101897.3, 101824.5, 101743.5, 101588.1, 101458.6, 101309.5, 
    101185.6, 101043.5, 100905.9, 100742.5, 100598.9, 100480.7, 100402.9, 
    100364.7,
  101841.6, 101813.5, 101733, 101624.3, 101505, 101382.9, 101278.1, 101161.4, 
    100969, 100781.9, 100642.4, 100499.9, 100337.7, 100232.8, 100162.8,
  101780.9, 101725.4, 101607.6, 101525.1, 101403.7, 101381.5, 101258.5, 
    101058.8, 100881.1, 100715.1, 100555.1, 100342.5, 100137.4, 100026.3, 
    99951.62,
  101899.8, 101851.3, 101781.4, 101687.6, 101632.9, 101571.2, 101514.2, 
    101534.5, 101579.2, 101224.6, 101264.6, 101465.5, 101265, 100780.9, 
    100569.9,
  101860.8, 101776.1, 101703.1, 101625.9, 101577.7, 101328.8, 101521.3, 
    101403.7, 101369.3, 101422.6, 101362.3, 101329.9, 101279.8, 99399.9, 
    99977.28,
  101832.4, 101760.3, 101690.8, 101648.2, 101462.3, 98097.89, 101241.1, 
    101532.8, 101412.6, 101303.2, 101205.4, 101148.1, 101074.7, 101042.2, 
    101003.9,
  101855, 101790.9, 101738.3, 101680.1, 101619.6, 101351.1, 97736.43, 
    101052.5, 101275.4, 101283.3, 101166.2, 101046.4, 100981, 100933, 100885.3,
  101921.9, 101879.8, 101839.3, 101779.9, 101739.5, 101654.6, 101396.6, 
    95443.89, 94641.66, 101042.4, 101239.8, 101104.1, 101093, 101017.6, 
    100986.1,
  101997.3, 101968.6, 101920.4, 101892.6, 101801.5, 101765.1, 101670.3, 
    101465.9, 101244.6, 101387.7, 101282.1, 101178.9, 101109.5, 101010.9, 
    100967.4,
  102064.1, 102075.8, 102053.9, 102039.5, 102000.2, 101900.1, 101799, 101734, 
    101589.5, 101387.4, 101256.6, 101136.9, 101014.6, 100905.8, 100818.3,
  102142.1, 102163.3, 102169.1, 102181.6, 102118.1, 102049.1, 101901.5, 
    101686.1, 101493.2, 101352.9, 101198.4, 101039.8, 100887.2, 100750.1, 
    100632.8,
  102225.1, 102287.9, 102331.6, 102341.5, 102279.4, 102151.6, 101973.1, 
    101779.5, 101540.3, 101299.6, 101099.7, 100926.6, 100739.2, 100580.6, 
    100426.4,
  102324.2, 102360.7, 102391.1, 102379.5, 102279.3, 102178.6, 101991.2, 
    101716.3, 101450.7, 101213.3, 101020.2, 100815.2, 100603.9, 100430.8, 
    100268.2,
  102620.5, 102538.4, 102425.5, 102286.1, 102183.8, 102117.2, 101965.1, 
    101839.3, 101676.3, 101110.6, 100955.6, 101002.2, 100663.6, 100109.2, 
    99862.08,
  102762.8, 102676.7, 102586.6, 102457.1, 102321.3, 101986.7, 102167.4, 
    101881.8, 101685.2, 101559.8, 101334.7, 101143.2, 100902.4, 98872.55, 
    99385.46,
  102845.5, 102787.2, 102714.2, 102657.3, 102323.2, 98808.26, 102001.6, 
    102224.1, 101965.9, 101714.4, 101459.7, 101283, 101047.6, 100863.1, 
    100607.1,
  102892.9, 102837.9, 102784.5, 102736.1, 102638.7, 102229.3, 98402.62, 
    101762.9, 101808.8, 101771.9, 101549.4, 101360.7, 101176.5, 101008.4, 
    100783.7,
  102900.1, 102866.4, 102816.7, 102781.7, 102704.4, 102602.3, 102237.8, 
    95988.6, 95170.7, 101570.1, 101625.1, 101391, 101240.4, 101058.5, 100969.6,
  102862.9, 102820.5, 102765.9, 102757.2, 102672.2, 102581, 102459.1, 
    102172.9, 101822.5, 101818.2, 101625.3, 101420, 101252.3, 101095.7, 
    100999.2,
  102810.8, 102773, 102719.9, 102720.5, 102680.1, 102576.8, 102426.8, 
    102297.2, 102100.4, 101826.6, 101619.4, 101433.3, 101239.2, 101085.6, 
    100971.5,
  102744.3, 102672.1, 102613.8, 102627.6, 102560.4, 102505.9, 102393.5, 
    102194.3, 101981.9, 101805.2, 101622.3, 101427.6, 101242.3, 101073.3, 
    100938.8,
  102678.2, 102599.7, 102561.4, 102544.8, 102500.6, 102436.7, 102340.7, 
    102217.7, 102031.4, 101796.3, 101612.9, 101431.6, 101236.4, 101059, 
    100912.2,
  102588.9, 102480.4, 102395, 102359.1, 102302, 102294.4, 102267.8, 102121.1, 
    101935.8, 101734.6, 101593, 101419.5, 101226.4, 101056, 100896.2,
  102935.2, 102935.3, 102907.9, 102796.9, 102699.8, 102559.8, 102375.4, 
    102315.8, 102263.7, 101760.6, 101682.1, 101770.6, 101406.4, 100742.3, 
    100393,
  102764.9, 102742.6, 102716.4, 102634.6, 102506.6, 102128, 102298.9, 
    102048.7, 101977.8, 102019.4, 101918.3, 101815.1, 101620.3, 99539.59, 
    99992.23,
  102557.8, 102543.4, 102494.8, 102451.2, 102180.9, 98715.37, 101792.3, 
    102159.5, 102009.2, 101919.4, 101856, 101799.6, 101649.7, 101513.4, 
    101270.3,
  102343.2, 102336.4, 102279.1, 102190, 102091.7, 101775, 98082.53, 101397.2, 
    101701.9, 101821.9, 101799.8, 101732.4, 101651.6, 101523.7, 101360.9,
  102163.3, 102159.8, 102090.1, 101987.8, 101880.4, 101773.3, 101538.4, 
    95615.09, 94805.85, 101356.6, 101719.9, 101647.2, 101624.2, 101484.1, 
    101402.6,
  102004.1, 101990.1, 101891.7, 101799.9, 101640.6, 101528.6, 101448.4, 
    101296.5, 101196, 101533.1, 101582.6, 101584.4, 101554.5, 101454.7, 101360,
  101865.2, 101857.2, 101757.4, 101653.9, 101489.9, 101342, 101235.5, 
    101261.7, 101409.3, 101443.5, 101486.5, 101504.4, 101461.2, 101398.5, 
    101302.3,
  101754.2, 101740.3, 101633.5, 101507, 101297.7, 101184.8, 101074.8, 
    101071.4, 101241.8, 101388.7, 101425.2, 101404.2, 101371.5, 101328.1, 
    101247.1,
  101665.9, 101656.2, 101559.9, 101390.4, 101218.8, 101097.3, 100998.6, 
    101118.5, 101304.8, 101320.5, 101330.4, 101315.9, 101278.6, 101234.7, 
    101171.7,
  101616.5, 101550.5, 101428.9, 101280.2, 101148.5, 101057.3, 101007.2, 
    101094.7, 101203.8, 101238.9, 101302.2, 101257.7, 101186.3, 101144.8, 
    101087.4,
  100951.2, 100869.8, 100791.2, 100698.4, 100648.7, 100602.4, 100526.3, 
    100482.6, 100455.7, 100106.8, 100206.1, 100573, 100576.6, 100301.2, 
    100163.8,
  100865.3, 100741.9, 100635.9, 100524.2, 100447.4, 100220.6, 100426.6, 
    100268.7, 100187.8, 100199.6, 100225.5, 100388.7, 100616.2, 98934.71, 
    99644.1,
  100804.6, 100684.6, 100572.1, 100481.2, 100288, 96994.54, 100154.3, 
    100412.3, 100255.8, 100116.8, 100080.8, 100252.5, 100548, 100783.5, 100858,
  100793.1, 100685.9, 100592.2, 100512.6, 100472.9, 100207.6, 96636.22, 
    99951.47, 100143.4, 100128.3, 100074.7, 100261.5, 100616.8, 100854.7, 
    100937.2,
  100810.8, 100745.4, 100686.3, 100627, 100633, 100534.9, 100305.1, 94403.77, 
    93685.2, 99994.33, 100276.8, 100444.7, 100717.9, 100862.6, 101008.8,
  100857.1, 100822.4, 100774.7, 100787.8, 100723, 100723, 100658.6, 100497.3, 
    100330.4, 100429, 100485.3, 100632.8, 100825.5, 100951, 101059,
  100902.7, 100924.4, 100923.8, 100940, 100939.7, 100888.4, 100852.9, 
    100843.5, 100780.5, 100668.3, 100686.9, 100793.1, 100886.1, 100983.5, 
    101065.2,
  100984.2, 101031.6, 101050.6, 101090.4, 101067.8, 101074.2, 101009, 
    100940.2, 100886.8, 100877.3, 100862.1, 100876.3, 100913.2, 100974.2, 
    101045.2,
  101095.4, 101161.4, 101245.7, 101283.5, 101296.8, 101246, 101191.8, 
    101154.6, 101068.8, 100979.1, 100930.1, 100907, 100896.6, 100912.9, 
    100953.4,
  101261.5, 101313.3, 101389.6, 101444.5, 101443.3, 101419.9, 101344.5, 
    101219.9, 101124.1, 101029.3, 100989.5, 100935.2, 100891.3, 100880.5, 
    100878.6,
  101215.4, 101110, 100972.7, 100796.9, 100688.7, 100598.3, 100400.7, 
    100207.5, 99987.09, 99384.48, 99196.94, 99278.75, 99127.03, 98864.66, 
    98924.62,
  101357.1, 101244.5, 101143.1, 100962, 100804, 100491.4, 100624.2, 100301.2, 
    100053.9, 99787.52, 99453.96, 99173.59, 99167.27, 97508.64, 98363.6,
  101460, 101369.7, 101298.8, 101182, 100831.4, 97305.16, 100510.5, 100626.3, 
    100328.7, 99955.02, 99504.94, 99157.65, 99085.88, 99272.99, 99520.46,
  101547.8, 101482.1, 101442.9, 101328.4, 101199.3, 100759.9, 96963.42, 
    100287.7, 100252.5, 100102.1, 99737.82, 99332.47, 99251.45, 99475.1, 
    99687.7,
  101635.4, 101606.1, 101582.3, 101480.9, 101367.8, 101193.3, 100816.2, 
    94604.46, 93843.66, 100133.5, 100103.4, 99773.01, 99660.98, 99698.85, 
    99872.48,
  101708.8, 101716.6, 101682.6, 101608.3, 101459.9, 101308, 101144.8, 
    100877.2, 100539, 100553.2, 100367.4, 100158.2, 100073.3, 100074.9, 
    100153.9,
  101779, 101834.8, 101799.1, 101743.4, 101617.2, 101441.6, 101228.9, 
    101087.5, 100926.7, 100741.7, 100580.4, 100473.3, 100389.8, 100366.2, 
    100378.5,
  101894, 101946.6, 101902.1, 101841.3, 101678.1, 101531.5, 101333.8, 
    101114.9, 100935.6, 100833.2, 100726.3, 100634.3, 100590.3, 100580.8, 
    100575,
  102020.5, 102066.3, 102037.4, 101941.7, 101806.9, 101635.5, 101419.6, 
    101236.8, 101069, 100925.7, 100818.6, 100751.9, 100701.5, 100677.8, 
    100665.5,
  102168.7, 102145.7, 102077.8, 101961.4, 101815.9, 101673.3, 101488.7, 
    101247.1, 101068.5, 100925.2, 100846.8, 100785.4, 100775.6, 100768.8, 
    100741.6,
  102182, 102020, 101799.1, 101556.7, 101379.1, 101225.4, 101045.7, 100875.5, 
    100693.5, 100111.1, 99906.78, 99880.07, 99539.02, 99098.16, 98969.47,
  102172.2, 101951.5, 101740.9, 101517.7, 101331.4, 100940.4, 101066.7, 
    100767.4, 100540.8, 100349.6, 100027.3, 99697.73, 99458.93, 97602.05, 
    98277.55,
  102154, 101920.5, 101695.9, 101532.2, 101192.5, 97650.47, 100770.2, 
    100924.8, 100651.5, 100362.8, 99948.88, 99571.12, 99208.12, 99189.25, 
    99272.78,
  102138.5, 101909.2, 101689.1, 101501.7, 101344.2, 100949.7, 97133.11, 
    100448.5, 100461.7, 100357.2, 100010.3, 99575.23, 99148.69, 99072.09, 
    99211.75,
  102125.7, 101923.5, 101709.7, 101525.9, 101377.3, 101227.6, 100879, 
    94687.91, 93895.2, 100210, 100151.2, 99754.3, 99367.28, 99138.85, 99279.85,
  102123.9, 101923.4, 101716.6, 101544.5, 101362.4, 101221.9, 101083.6, 
    100837.2, 100534.9, 100537.2, 100296.5, 100005.6, 99768.7, 99556.6, 
    99522.19,
  102122.7, 101952.4, 101757.3, 101609.3, 101437.8, 101282.6, 101101.2, 
    100988.4, 100872.5, 100670.3, 100451, 100231.3, 100012.5, 99881.89, 
    99806.45,
  102129.1, 101963.4, 101788.8, 101637, 101448, 101319.9, 101165.8, 100991.2, 
    100868.2, 100772.8, 100620.9, 100449.4, 100262.9, 100104.2, 99969.59,
  102148.3, 102014.3, 101873.7, 101735.6, 101585.4, 101423.1, 101250.9, 
    101122.5, 101016.8, 100900, 100765.6, 100620, 100447, 100268, 100070.5,
  102163, 102022.9, 101886.5, 101770.5, 101619.1, 101491.3, 101354, 101181.4, 
    101061.5, 100956.6, 100892.3, 100786.1, 100623.7, 100430.3, 100171.6,
  101819.2, 101827.6, 101814.2, 101693.9, 101540.7, 101419.3, 101261.1, 
    101118.6, 100966.8, 100428.1, 100273, 100298, 99892.34, 99235.83, 98921.89,
  101798.2, 101824.8, 101830, 101737.8, 101575.6, 101220.7, 101348, 101060, 
    100849.8, 100735.6, 100546, 100357.2, 100136.4, 98116.73, 98645.57,
  101770.7, 101830.8, 101841.8, 101834.9, 101524.9, 97963.41, 101151, 
    101310.5, 101089.2, 100801.5, 100547.4, 100356.3, 100145.9, 100005.2, 
    99902.7,
  101753.8, 101835.8, 101862.3, 101846.2, 101774.2, 101356, 97551.16, 100869, 
    100841.2, 100802.3, 100558.4, 100328.1, 100139.6, 99971.65, 99967.8,
  101758.5, 101880.1, 101916.5, 101918.7, 101845.7, 101732.7, 101356.7, 
    95134.77, 94345.61, 100585.3, 100587.9, 100267.6, 100099, 99909.55, 
    99905.87,
  101773.1, 101911, 101946.3, 101966.6, 101874.2, 101753.1, 101629.6, 
    101342.9, 100942.7, 100866.4, 100572.8, 100245, 100023.2, 99914.88, 
    99856.56,
  101802.2, 101958.5, 102035.4, 102063.4, 101991.2, 101854.9, 101655.5, 
    101502.6, 101264.4, 100927.4, 100577, 100203.2, 99879.43, 99760.88, 
    99781.53,
  101841.8, 102007, 102088.9, 102109.8, 102021.1, 101911.1, 101737.8, 101508, 
    101246.2, 100980.3, 100632.5, 100209.7, 99805.05, 99612.09, 99611.45,
  101875.7, 102065.4, 102174.9, 102200.5, 102150.3, 102022.2, 101821.4, 
    101644.9, 101404.8, 101097.9, 100733.3, 100298, 99824.54, 99479.03, 
    99417.27,
  101925.9, 102088.2, 102198.6, 102221.1, 102162.8, 102080.7, 101920.4, 
    101700.1, 101466.9, 101183.3, 100885.6, 100469.3, 99999.53, 99571.11, 
    99310.03,
  101037.1, 101361.9, 101656.1, 101734.9, 101750.5, 101648.9, 101457.3, 
    101259.7, 101060.4, 100495.5, 100338.3, 100381, 99984.49, 99223.11, 
    98800.73,
  101196.9, 101541, 101714.9, 101790.4, 101733.4, 101402.4, 101457.8, 
    101095.2, 100809.8, 100684, 100515.7, 100384.7, 100168.1, 98096.54, 
    98426.68,
  101438.2, 101686.8, 101809.5, 101892.2, 101641.3, 98090.86, 101171.4, 
    101304.7, 101011.2, 100686.3, 100414.9, 100307, 100172.1, 100042.1, 
    99692.51,
  101639.4, 101774.5, 101901.3, 101909.8, 101882.3, 101428.7, 97601.46, 
    100736.4, 100667.5, 100590.4, 100333.2, 100176.4, 100124.3, 100079.5, 
    99863.88,
  101782.2, 101909.8, 101989.9, 102004.7, 101936.9, 101763, 101346.5, 
    95107.65, 94270.71, 100349.4, 100289.1, 100024.4, 100056.8, 100040.8, 
    100014,
  101900.2, 102004.2, 102059.1, 102072, 101964.4, 101801.8, 101607.4, 
    101245.7, 100786.1, 100622.8, 100257.4, 99969.67, 99975.34, 100050.7, 
    100057,
  101980.7, 102095.1, 102164.3, 102174.5, 102078.7, 101894.7, 101654.4, 
    101435.2, 101140, 100725.5, 100321.3, 100021.7, 99921.98, 100032.4, 
    100084.4,
  102033.5, 102164.8, 102234.9, 102228.4, 102115.9, 101978.9, 101759.8, 
    101466.7, 101156.4, 100840.7, 100482.6, 100151.8, 99991.32, 100066, 100115,
  102080.4, 102241.3, 102318.3, 102319.4, 102231.4, 102089.3, 101877.4, 
    101645.9, 101376.1, 101031.8, 100673.2, 100338.8, 100097, 100083.4, 100152,
  102126.9, 102273.6, 102337, 102316.3, 102236, 102155.5, 101992.1, 101739.5, 
    101478.1, 101175.8, 100874.2, 100549.5, 100249.7, 100109.1, 100163.7,
  101449.8, 101577.4, 101634, 101612.6, 101538.2, 101435.3, 101295.3, 
    101170.4, 101017.4, 100494.3, 100370.8, 100488.5, 100234.9, 99695.25, 
    99376.9,
  101707.7, 101759.3, 101738.2, 101682, 101540.2, 101206, 101307.1, 101051.7, 
    100827, 100669.9, 100489.2, 100367.7, 100257.1, 98301.84, 98740.15,
  101862.6, 101870.8, 101847.6, 101804.9, 101473.5, 97932.66, 101080.8, 
    101227.4, 100975.7, 100677.6, 100425.8, 100305.8, 100201, 100117.3, 
    99822.2,
  101975.3, 101965.6, 101930.3, 101864.5, 101765.5, 101332.5, 97519.21, 
    100795.1, 100766.9, 100676.9, 100438.2, 100292, 100195.8, 100079.2, 
    99741.62,
  102050.2, 102066.2, 102029.9, 101964.2, 101855.1, 101713.2, 101318.8, 
    95132.78, 94352.87, 100503.5, 100505.1, 100297.1, 100223.3, 100033.6, 
    99784.95,
  102100.1, 102127.3, 102101.7, 102052.6, 101919.6, 101780.9, 101607.4, 
    101302.3, 100907, 100794, 100553.9, 100355.7, 100257.8, 100087.8, 99837.57,
  102104.1, 102159, 102170.5, 102140.1, 102027.2, 101878.2, 101670.9, 101489, 
    101257.1, 100928.5, 100646.1, 100430.2, 100302.1, 100161.6, 99944.63,
  102068, 102147.7, 102192.2, 102182, 102064.7, 101962.5, 101777, 101527, 
    101282, 101043.8, 100789.2, 100534.9, 100371.7, 100249.7, 100073.3,
  102000.1, 102109.1, 102206, 102216.5, 102119.9, 102043.6, 101873.9, 
    101682.8, 101472.7, 101213.7, 100952.2, 100676.9, 100472.2, 100349.5, 
    100207.2,
  101914.4, 102018.4, 102138.9, 102169.1, 102105.1, 102086.6, 101966.5, 
    101755.3, 101546.8, 101321.7, 101113.2, 100860.4, 100607.1, 100457.3, 
    100367.1,
  102058.3, 102060.5, 101978.2, 101853.1, 101727, 101631, 101510, 101412.1, 
    101271.8, 100785.1, 100660.3, 100774, 100524.3, 100070.5, 99891.38,
  102089.4, 102065.2, 102018.6, 101912.3, 101765.1, 101450.3, 101562.6, 
    101338.4, 101162.4, 101052.8, 100857.5, 100725.1, 100611.7, 98678.81, 
    99259.67,
  102074.6, 102078.2, 102042.7, 102020.6, 101705.8, 98164.38, 101372.7, 
    101512.2, 101294.2, 101072.8, 100824.9, 100661, 100506.6, 100427.2, 
    100301.6,
  102060.4, 102087.1, 102063, 102041.4, 101958.2, 101582, 97740.53, 101125.6, 
    101144, 101070.9, 100814.9, 100599.5, 100429.6, 100303, 100139.9,
  102025.8, 102104.8, 102100.8, 102089.5, 102006.7, 101895.2, 101541.7, 
    95377.13, 94593.67, 100865.2, 100841.8, 100551.1, 100369.8, 100178.9, 
    100033.5,
  101976.1, 102083.8, 102104.6, 102119.2, 102026.5, 101921.1, 101762.1, 
    101508.6, 101174.6, 101116.2, 100852.7, 100552.9, 100337.1, 100112.2, 
    99922.29,
  101915.2, 102062.4, 102116.4, 102157.9, 102085.5, 101978.1, 101786.4, 
    101642.3, 101443.6, 101178.2, 100889.9, 100588.5, 100321.8, 100089.3, 
    99884.12,
  101878.9, 102036.1, 102082.6, 102163.8, 102095.5, 102024.7, 101842.9, 
    101644.4, 101440.1, 101248.2, 100976.5, 100654.7, 100357.5, 100107.2, 
    99894.34,
  101838.8, 101960, 102081.6, 102187.7, 102153.5, 102090.5, 101933.9, 
    101760.8, 101565.6, 101342.8, 101079.8, 100754.4, 100423.4, 100161.6, 
    99947.23,
  101819, 101923.9, 102029.7, 102139.4, 102151, 102132, 102011.7, 101816.9, 
    101634.2, 101421.5, 101213.5, 100891.1, 100530.4, 100262.9, 100060.7,
  102310.7, 102367.8, 102339.7, 102253, 102170.1, 102064.2, 101937.8, 
    101834.8, 101704.5, 101207.4, 101091.6, 101125.1, 100758.5, 100173.1, 
    99917.84,
  102345.1, 102345.2, 102351.2, 102278.7, 102171.8, 101849.2, 101971.4, 
    101740, 101585.9, 101502.1, 101327.7, 101132.4, 100890.7, 98859.03, 
    99370.86,
  102329, 102360.8, 102352.4, 102342.5, 102075.4, 98514.95, 101750.4, 
    101912.6, 101725.2, 101543.7, 101325.5, 101119.5, 100873.8, 100685.7, 
    100492.1,
  102296.4, 102351.1, 102371.5, 102348.9, 102277.5, 101913.1, 98084.62, 
    101497.4, 101556, 101541.5, 101324.8, 101087.9, 100828.1, 100627.6, 
    100457.6,
  102308.2, 102393.3, 102404, 102393.1, 102315.5, 102199.9, 101869.3, 
    95722.78, 94927.41, 101303.4, 101332.6, 101039.8, 100769, 100534.6, 
    100390.8,
  102341.1, 102413.5, 102410.6, 102424, 102321.3, 102210.7, 102081.8, 101852, 
    101540.1, 101538.1, 101300.2, 100997.3, 100685.9, 100456.9, 100292.6,
  102380.9, 102440.2, 102442.8, 102464.1, 102382.5, 102250.2, 102086, 
    101967.6, 101786.7, 101540.6, 101274.1, 100951.2, 100611.6, 100397.2, 
    100225.5,
  102429.4, 102441.9, 102433.4, 102461.7, 102366.5, 102267.1, 102105.3, 
    101919, 101732.1, 101532.9, 101269.6, 100915, 100578.3, 100377.6, 100227.9,
  102457.7, 102457.9, 102434.1, 102452.2, 102377.8, 102267.8, 102128.1, 
    101985.6, 101805.1, 101560.8, 101283.6, 100908.1, 100573.9, 100395.3, 
    100262.1,
  102500.8, 102431.1, 102375, 102333.1, 102254, 102189.9, 102116.3, 101958.1, 
    101799.5, 101569.9, 101322.5, 100933.3, 100608.6, 100440.2, 100325.5,
  102430.6, 102406.4, 102362.3, 102267.4, 102192.2, 102095.2, 101987.1, 
    101928.2, 101856.3, 101412.1, 101382.5, 101535.2, 101239.6, 100634.2, 
    100328.2,
  102443.3, 102367, 102310.2, 102220.3, 102111, 101813.5, 101966, 101775.9, 
    101678.8, 101675.4, 101576, 101509, 101344.5, 99300.91, 99793.88,
  102393.6, 102315.5, 102213.2, 102158.8, 101901.1, 98394.14, 101612.1, 
    101874.6, 101712.4, 101610.1, 101498.8, 101429.5, 101272.4, 101117.4, 
    100926.8,
  102327.1, 102240.9, 102114, 102016.3, 101913.3, 101608.5, 97862.5, 
    101262.7, 101461, 101508.1, 101419.8, 101314.6, 101178.1, 101029.9, 100871,
  102284.9, 102145.1, 101995.2, 101871, 101758.5, 101657.2, 101411, 95426.94, 
    94625.76, 101102.8, 101318.6, 101178, 101057, 100891.4, 100790.9,
  102187.3, 102001.9, 101834, 101700.1, 101556, 101458, 101369.8, 101221.7, 
    101052.1, 101231.6, 101150.3, 101044.4, 100906.4, 100756.8, 100669.3,
  102086.4, 101904.3, 101735.3, 101596.5, 101460.3, 101309.8, 101168.1, 
    101125.2, 101094.4, 101040.2, 100980.9, 100892.4, 100736.9, 100612.8, 
    100532.3,
  102022.5, 101841.6, 101665.2, 101501.2, 101318.4, 101155.3, 101003.9, 
    100876.5, 100855.7, 100889, 100848.1, 100735.1, 100588.8, 100476.7, 
    100397.2,
  102000.5, 101836, 101663.4, 101477.2, 101288.3, 101085.3, 100914.6, 100866, 
    100867.5, 100820.3, 100724.1, 100582.1, 100427.1, 100330.4, 100265.3,
  102021.1, 101826.2, 101635.8, 101467, 101265.3, 101072.1, 100938.9, 
    100843.7, 100818.2, 100727.6, 100617, 100429.8, 100260.5, 100177.8, 100120,
  101732.1, 101736.1, 101740, 101720.7, 101721.3, 101682.3, 101639.4, 
    101655.5, 101685.4, 101360.2, 101447.2, 101738, 101591.9, 101132.3, 
    100892.1,
  101659.6, 101605, 101562, 101516, 101463.7, 101249.9, 101417.2, 101360, 
    101380.2, 101488.5, 101530.9, 101639.9, 101694.9, 99806.32, 100416.8,
  101589.7, 101489.9, 101401.7, 101344.8, 101128.8, 97689.5, 100888.3, 
    101163.1, 101087.3, 101168.8, 101297.7, 101454.4, 101600.8, 101675.3, 
    101648.6,
  101507.4, 101398.1, 101300.4, 101205, 101110.3, 100793.1, 97144.42, 100499, 
    100835.6, 100905, 101063.1, 101241, 101469.4, 101613.2, 101677,
  101486.5, 101376.6, 101287.1, 101182.2, 101073.6, 100956.5, 100675.2, 
    94773.78, 93972.67, 100402.7, 100813.7, 101013.9, 101317.7, 101498.8, 
    101657.1,
  101511.8, 101400.1, 101294.8, 101183.8, 100987.1, 100848.9, 100742.4, 
    100559.6, 100409, 100653, 100651.5, 100859.4, 101172.2, 101417.8, 101589.6,
  101558.4, 101455.9, 101327.6, 101174.4, 100945.3, 100714.2, 100538.3, 
    100495.4, 100421.8, 100407.4, 100533.5, 100748, 101058.3, 101337.6, 
    101519.1,
  101601.3, 101471.1, 101314.5, 101121.1, 100829.9, 100587.4, 100378, 
    100247.2, 100225, 100306.7, 100443.6, 100664.6, 100987.8, 101271.5, 
    101465.4,
  101648.5, 101523.2, 101361.7, 101144.9, 100855.1, 100530.9, 100283, 
    100215.5, 100248, 100242.9, 100368.6, 100622.1, 100936.3, 101218.1, 
    101413.3,
  101725.1, 101553.5, 101369.5, 101136.9, 100823.8, 100494.2, 100225.2, 
    100030.7, 100097.4, 100192.9, 100349.5, 100604.1, 100904.4, 101186.1, 
    101383.1,
  101504.5, 101462.9, 101418.2, 101372.8, 101345.6, 101311.7, 101300.7, 
    101349.3, 101438, 101190.8, 101350.7, 101705.7, 101655.8, 101311, 101152.6,
  101489.7, 101399.7, 101341.2, 101279.6, 101236.7, 101039.1, 101244.4, 
    101182.9, 101234.1, 101388.9, 101501.7, 101640.7, 101768.4, 99974.41, 
    100653.1,
  101368.3, 101264.2, 101178.8, 101125, 100989, 97599.8, 100926.5, 101221.5, 
    101152.2, 101213.1, 101364.6, 101529.8, 101704.3, 101834.8, 101882.9,
  101245.8, 101119.6, 101000.7, 100924.6, 100901.4, 100724.4, 97158.04, 
    100734.4, 101081.5, 101099.5, 101212.4, 101394.3, 101619, 101824.7, 
    101939.1,
  101131.3, 100991.9, 100880.4, 100803.8, 100825, 100794.4, 100656.9, 
    94878.2, 94216.48, 100814.6, 101105.3, 101267.9, 101534.9, 101765, 
    101975.8,
  101050.4, 100905.3, 100789.8, 100784.8, 100714.5, 100666.3, 100651.5, 
    100624.3, 100600.1, 100984.9, 101017, 101185, 101472.7, 101773.6, 101973.7,
  101001.6, 100865.1, 100775.8, 100734.7, 100635.9, 100529.1, 100442.2, 
    100510.9, 100671, 100867, 101001, 101140.3, 101455.8, 101792.1, 101986.8,
  100983.2, 100844.2, 100742.5, 100648.1, 100487.1, 100371.1, 100292.8, 
    100301.8, 100482.7, 100822.1, 100984.4, 101138, 101496.9, 101841.7, 
    102037.7,
  101004.2, 100861.3, 100733.9, 100580.8, 100388.9, 100245.8, 100200.7, 
    100276.2, 100501, 100811.5, 100980.1, 101195.4, 101581.8, 101907.3, 
    102098.4,
  101050.6, 100874.7, 100706.5, 100530.2, 100326.5, 100204.2, 100187.2, 
    100257, 100547.3, 100800.4, 101006.7, 101319.9, 101703.6, 102002.7, 
    102165.6,
  100781.7, 100775.6, 100802, 100830.6, 100931.7, 100993, 101036.4, 101091.8, 
    101108.1, 100830.2, 100994.1, 101364.3, 101307.7, 100982.2, 100846.2,
  100690.5, 100652.6, 100652.6, 100655.9, 100704, 100637.6, 100929.4, 
    100982.7, 101034.9, 101136.5, 101234.5, 101406, 101522.2, 99737.03, 
    100425.1,
  100644.4, 100571.5, 100541.6, 100513.1, 100420.1, 97134.23, 100505.8, 
    100934.2, 101028.7, 101114.6, 101237.7, 101413.3, 101580.9, 101671.5, 
    101704.7,
  100572.8, 100484.8, 100441.6, 100403.1, 100417.3, 100246.4, 96762.59, 
    100424.8, 100927.7, 101077.6, 101242.6, 101396.6, 101597.6, 101745.2, 
    101825,
  100508.3, 100431.9, 100400.3, 100402.4, 100453.8, 100502.7, 100265.8, 
    94674.02, 94186.16, 100795.9, 101245.1, 101397.1, 101618, 101737.9, 
    101909.9,
  100477.2, 100382.2, 100329.6, 100384.9, 100416.1, 100471.8, 100507.7, 
    100438.5, 100494.9, 100991.4, 101190.8, 101411.5, 101626.2, 101793, 
    101935.2,
  100453.2, 100373, 100344.2, 100335.2, 100383.8, 100450.2, 100454.2, 
    100589.9, 100822.5, 100977.7, 101202.6, 101441.8, 101646.7, 101822.4, 
    101914.6,
  100486.9, 100409.7, 100352.4, 100298.5, 100282.3, 100412.5, 100463.2, 
    100543.7, 100757.8, 101025.1, 101263.9, 101487.5, 101700, 101865.5, 
    101921.9,
  100546.5, 100461.6, 100384.4, 100306, 100302.9, 100404.6, 100512.2, 
    100708.1, 100922.6, 101124.6, 101337.9, 101562.2, 101761.6, 101891.3, 
    101948.5,
  100650.6, 100546.3, 100454.8, 100374.9, 100367.3, 100467.2, 100599.6, 
    100763.4, 100976.8, 101183, 101433.4, 101657.5, 101837.3, 101949.6, 
    101960.3,
  100763.4, 100793.4, 100788.5, 100754.8, 100705.2, 100689, 100732.8, 
    100848.2, 100924.5, 100630.2, 100751.7, 100932.6, 100621.4, 100039.2, 
    99699.1,
  100767.9, 100723.2, 100703.1, 100646.4, 100593, 100427.6, 100686.4, 
    100778.2, 100855.2, 100927.6, 101010.4, 101009.2, 100877.3, 98894.06, 
    99397.94,
  100692.2, 100627.4, 100584.4, 100549.4, 100407, 97056.89, 100441.7, 
    100793.9, 100880.1, 100940.6, 101042.5, 101083.5, 101025.5, 100927.9, 
    100745.4,
  100618, 100546.1, 100485.3, 100461.5, 100434.9, 100225.8, 96722.55, 
    100411.1, 100792.2, 100931.8, 101079.1, 101138.2, 101140.2, 101096.5, 
    101020,
  100539.2, 100465.2, 100399.7, 100379.7, 100432.3, 100443.7, 100261.2, 
    94648.28, 94134.31, 100718.6, 101124.1, 101211.7, 101265.9, 101224.8, 
    101249.5,
  100506.7, 100396.2, 100361.6, 100335.7, 100400.1, 100487.8, 100522.6, 
    100455.4, 100472.1, 100939.4, 101141.7, 101294.1, 101372.7, 101399.9, 
    101416.2,
  100447.8, 100364.5, 100366.7, 100364.1, 100413.5, 100526.8, 100566.2, 
    100606.7, 100788, 100978.7, 101202, 101392, 101495.6, 101559.6, 101592.2,
  100459, 100383.1, 100372.4, 100352.5, 100384.4, 100528.4, 100563.1, 
    100578.6, 100766.1, 101055.6, 101289, 101492.5, 101624.7, 101704.7, 
    101762.5,
  100511.1, 100446.7, 100401.1, 100390.6, 100461.6, 100547.9, 100577.9, 
    100718.5, 100935.5, 101186.5, 101401.1, 101610.8, 101737.9, 101827.7, 
    101887.2,
  100637.6, 100571.5, 100533.7, 100508.5, 100529.2, 100587.1, 100659.4, 
    100811.3, 101050.8, 101272.3, 101514.5, 101708.8, 101841.4, 101942.5, 
    102002.6,
  101198.6, 101249.6, 101248.2, 101253.6, 101262.4, 101256.8, 101231.1, 
    101221.1, 101223.4, 100880.9, 100961.1, 101204.4, 100978, 100407.3, 
    100010.6,
  101194.5, 101174.9, 101186.9, 101155.7, 101140, 100950.7, 101128.9, 
    101075.6, 101076.1, 101106.3, 101137.6, 101157, 101058.4, 99036, 99438.2,
  101145.1, 101111.3, 101077.3, 101047.8, 100911.1, 97537.73, 100812.8, 
    101025.9, 101042.9, 101071.4, 101119.2, 101098.5, 100975.2, 100791.4, 
    100571.8,
  101077.6, 101021.5, 100953.1, 100920.8, 100892.9, 100713.4, 97105.95, 
    100685.7, 101022.3, 101050.8, 101093.9, 100996.1, 100881.3, 100718, 
    100655.1,
  101001.5, 100922.6, 100865.1, 100820.4, 100833.6, 100866.1, 100712.3, 
    94916.98, 94282.88, 100787.2, 101045.7, 100913.8, 100818.6, 100703.7, 
    100808.5,
  100941.5, 100857, 100819.2, 100829.1, 100827.1, 100828.6, 100823.6, 
    100806.8, 100720.3, 101008.6, 100970.6, 100879.5, 100827.9, 100844.2, 
    100952.9,
  100896.2, 100844.1, 100846.8, 100867.3, 100862.6, 100882.1, 100811.8, 
    100917.3, 101020.4, 101035.5, 100980.9, 100946.2, 100963.9, 101043.1, 
    101162.4,
  100901.7, 100871.3, 100881.8, 100869.4, 100878.1, 100895.9, 100885.7, 
    100969.3, 101081.2, 101127.6, 101124.6, 101144.2, 101218.7, 101325.4, 
    101438.6,
  100933.8, 100914.1, 100933.8, 100953.4, 100965.6, 100983.8, 101026.5, 
    101171.4, 101282.6, 101314.9, 101340.2, 101399.2, 101479.3, 101573, 
    101653.3,
  101020.6, 100990.1, 101005.4, 101021.2, 101045.7, 101099.8, 101200, 
    101320.5, 101428.6, 101472, 101568, 101649.5, 101722.8, 101807.3, 101868,
  101202.2, 101280.7, 101390.4, 101451.9, 101508.7, 101537, 101550.7, 
    101596.7, 101656.5, 101345.6, 101420.6, 101690.1, 101562.1, 101197.7, 
    101061.3,
  101319, 101382.7, 101432.8, 101426.4, 101433, 101251.3, 101463.9, 101426.8, 
    101447, 101516.7, 101529, 101589.1, 101632.2, 99823.18, 100465.1,
  101401.7, 101404.3, 101406, 101399.4, 101265.9, 97878.16, 101110.5, 
    101357.1, 101283.8, 101333, 101372, 101458.5, 101532.2, 101586.7, 101569.4,
  101413.4, 101410.8, 101355.8, 101313.4, 101270.9, 101064.6, 97451.43, 
    100900.8, 101206.1, 101243.8, 101300.1, 101349.2, 101437.7, 101501.2, 
    101498,
  101380.5, 101336.2, 101280.8, 101254, 101281.4, 101253.2, 101035.6, 
    95153.67, 94422.91, 100908, 101206.7, 101244.2, 101325.9, 101341.3, 
    101396.9,
  101328.8, 101289.6, 101253.9, 101279.2, 101195.6, 101145.3, 101108, 
    101014.9, 100875.3, 101066.6, 101074.8, 101138.8, 101191.3, 101239.9, 
    101299.2,
  101302.5, 101270.8, 101283.3, 101230.5, 101142.2, 101052.4, 100956.4, 
    100986.8, 100981, 100971.7, 100992.6, 101033.5, 101073.8, 101164, 101269.5,
  101309.5, 101307.7, 101272.4, 101168.7, 101033.4, 100961.3, 100931.4, 
    100880.2, 100849.7, 100837.2, 100888.5, 100962.4, 101078.5, 101228.8, 
    101381.8,
  101354, 101359.8, 101289.2, 101167.3, 101062.4, 100989.2, 100898.4, 
    100834.3, 100743.6, 100793.4, 100902.3, 101053.3, 101214.5, 101380.8, 
    101499.6,
  101439, 101408, 101339.7, 101222.7, 101086.2, 100979.9, 100886.5, 100816, 
    100825.3, 100901.1, 101083.4, 101257.1, 101414.6, 101555.2, 101652.9,
  101184.3, 101406.8, 101600.7, 101760, 101899.8, 101940.7, 101902.8, 
    101911.1, 101903.3, 101504.7, 101523.5, 101738.1, 101548, 101162.1, 
    101011.5,
  101096.3, 101302.6, 101534.2, 101713.6, 101815.9, 101659.5, 101880.5, 
    101756.1, 101719.2, 101739.5, 101673.1, 101694.6, 101698.8, 99859.62, 
    100527.5,
  101013.5, 101262, 101478.8, 101639.3, 101617.3, 98277.12, 101511.2, 
    101811.1, 101661.4, 101626.8, 101577.8, 101596.4, 101635.2, 101704, 101697,
  100951, 101253.6, 101426.5, 101573.8, 101596.3, 101462.3, 97866.43, 
    101304.6, 101570.1, 101551.8, 101514.3, 101503.8, 101558, 101661.4, 
    101719.9,
  101025.5, 101259.4, 101398.9, 101488.6, 101606.2, 101597.3, 101429, 
    95546.48, 94774.73, 101248.1, 101467.2, 101449.2, 101503.7, 101587.4, 
    101721,
  101100, 101290.7, 101368.6, 101479.7, 101454.3, 101474.9, 101446, 101359, 
    101248.9, 101451.7, 101402.5, 101432.9, 101470.4, 101570.7, 101685.7,
  101198.4, 101326, 101375.4, 101414.6, 101377.4, 101319.5, 101277.6, 
    101340.2, 101355.4, 101374.6, 101414.3, 101439.4, 101480.7, 101565.8, 
    101655.8,
  101297.3, 101343.9, 101352.1, 101309.1, 101177.4, 101138.6, 101148.5, 
    101176.6, 101241.1, 101354.1, 101412.1, 101448, 101495.1, 101557.4, 
    101625.4,
  101351.4, 101341.1, 101290.8, 101169.9, 101045.7, 101010.1, 101070.7, 
    101181, 101253.2, 101309.7, 101369.7, 101424.5, 101453.4, 101510.5, 
    101561.3,
  101363.7, 101292.5, 101211.1, 101048.6, 100906.8, 100926.9, 101007.1, 
    101089.8, 101168.8, 101221.2, 101300.1, 101375.3, 101420.1, 101489.3, 
    101540.3,
  100125.6, 100123.8, 100167.3, 100205.2, 100291.1, 100381.9, 100514, 
    100695.5, 100904.6, 100767.9, 101038, 101474.3, 101476.7, 101221.6, 
    101166.9,
  99892.7, 99850.91, 99880.05, 99929.31, 100015.1, 100034.3, 100385, 
    100539.4, 100737.8, 100995.6, 101217.1, 101458, 101625.2, 99907.09, 
    100647.9,
  99632.46, 99581.59, 99620.45, 99720.76, 99764.83, 96758.48, 100182.6, 
    100634.1, 100786.9, 101035.3, 101271.2, 101505.3, 101644.8, 101754.8, 
    101820.8,
  99414.69, 99351.25, 99431.15, 99604.07, 99840.08, 99873.26, 96796.83, 
    100479.3, 101001.7, 101199.5, 101400.4, 101540.4, 101690.1, 101792.2, 
    101855.1,
  99318.1, 99319.45, 99497.76, 99770.98, 100098.9, 100380.6, 100388.9, 
    94906.98, 94435.12, 101086.1, 101496.4, 101585.1, 101706.8, 101761.3, 
    101897.6,
  99682.98, 99730.4, 99909.59, 100158.5, 100368, 100640.8, 100861.4, 
    100902.2, 101022.4, 101430, 101529.4, 101615.9, 101703.4, 101788.8, 
    101893.7,
  100167.5, 100234.4, 100364.9, 100528.1, 100729, 100882.6, 101068.5, 
    101298.2, 101434.8, 101494, 101589.1, 101619.5, 101678.7, 101794.1, 101905,
  100527.5, 100606.8, 100718, 100833.1, 100958.2, 101109.2, 101238, 101332.6, 
    101471.9, 101603.7, 101643.3, 101661.7, 101741.5, 101847.7, 101951.4,
  100805.1, 100885.1, 100965.8, 101051.6, 101161.2, 101277.1, 101416.2, 
    101559.3, 101636.8, 101671.4, 101714.6, 101766.8, 101827.2, 101913.4, 
    101991.6,
  100977.1, 101034, 101112, 101191.5, 101300.7, 101419.6, 101516.2, 101580.3, 
    101640.1, 101673.6, 101758.3, 101829.8, 101888.5, 101958.8, 101989.5,
  101608.9, 101409, 101157.7, 100861.7, 100621.3, 100452.1, 100351.5, 100292, 
    100263.8, 99925.76, 99951.53, 100185.7, 100039.3, 99710.74, 99673.91,
  101507, 101187, 100860.7, 100516.6, 100249.4, 99918.66, 100054.6, 99979.9, 
    99924.66, 99917.49, 99888.18, 99908.11, 99949.71, 98287.91, 99069.94,
  101333.6, 100978.3, 100604.6, 100251.3, 99909.52, 96566.76, 99792.02, 
    100011.2, 99903.75, 99852.97, 99783.58, 99774.59, 99841.29, 99978.74, 
    100208.9,
  101242.6, 100880.6, 100490, 100196.8, 100018.2, 99781.43, 96434.88, 
    99904.04, 100087.3, 100042.5, 99937.59, 99883.79, 99933, 100135.4, 
    100387.3,
  101244.2, 100956.8, 100650.3, 100462.6, 100337.6, 100321.8, 100135.1, 
    94366.67, 93812.78, 100117.9, 100257.6, 100168.1, 100236.5, 100372.2, 
    100651.6,
  101362.6, 101185.4, 100984.1, 100833.7, 100729.3, 100728.2, 100728.2, 
    100613.8, 100490.6, 100642.7, 100609.1, 100585.5, 100644.8, 100758.5, 
    100944.6,
  101472.9, 101401.2, 101295.7, 101210.5, 101133.8, 101080.5, 101050.8, 
    101069.1, 101029.6, 100941.3, 100920.3, 100937.8, 100982.5, 101076.2, 
    101201.9,
  101608, 101597.2, 101545.1, 101485.1, 101411.2, 101374.2, 101315.1, 
    101243.8, 101206.4, 101203.7, 101194.1, 101214.6, 101262.5, 101337.2, 
    101416.7,
  101685.2, 101740.2, 101736.5, 101712.2, 101674.1, 101620.9, 101557.9, 
    101522.4, 101459.4, 101405.4, 101392.3, 101420.1, 101457.7, 101497.2, 
    101518.7,
  101771.8, 101834.1, 101852.1, 101832.5, 101796, 101765.4, 101717.6, 
    101634.5, 101583.1, 101544.7, 101586.7, 101612.1, 101631.9, 101644.2, 
    101620.7,
  101479.8, 101626.3, 101796.5, 101895.2, 101918.6, 101887.6, 101867.8, 
    101805.6, 101686.5, 101155.3, 101008.6, 101043, 100692.2, 100127.9, 
    99897.57,
  101331.3, 101479.9, 101686, 101816.4, 101865.8, 101700.4, 101910, 101727, 
    101593.1, 101456.2, 101206.8, 100947.5, 100691.4, 98694.35, 99200.38,
  101180.9, 101387.2, 101622.6, 101808.1, 101745.4, 98393.71, 101699.5, 
    101899.5, 101705.7, 101470.8, 101183.8, 100867.4, 100540.5, 100313.8, 
    100190.7,
  101038.5, 101342.3, 101613.2, 101820.4, 101915, 101701.8, 98063.83, 
    101483.9, 101596.6, 101500.4, 101195.4, 100802.8, 100424.9, 100119.5, 
    100059,
  101247.7, 101524, 101745.2, 101908.6, 101998.3, 102000.4, 101786.1, 
    95792.65, 94994.87, 101269.3, 101258.1, 100804.8, 100384.2, 99974.18, 
    100001.3,
  101576.2, 101735, 101875, 102001.8, 102014.5, 102022.4, 101981.9, 101805.9, 
    101566.6, 101567.9, 101290.7, 100885.3, 100458.5, 100072.1, 100057.8,
  101742.6, 101895.9, 102001.9, 102076.1, 102084.6, 102044.2, 101961.6, 
    101919.1, 101778.1, 101580, 101328.6, 100978.9, 100610.6, 100352.4, 
    100319.1,
  101876.5, 101972.3, 102053.3, 102095.9, 102064.4, 102029.6, 101941.4, 
    101817.1, 101721.7, 101603, 101385.1, 101074.3, 100817.4, 100681.3, 
    100639.2,
  101897.4, 102017.3, 102100.7, 102088.5, 102047.9, 101977.2, 101891.9, 
    101839.7, 101744.8, 101606.6, 101419.7, 101171.1, 100981.9, 100893, 
    100878.8,
  101957, 102052, 102052.6, 102015.8, 101940.2, 101877.8, 101810.6, 101735.3, 
    101664.8, 101559.6, 101440.4, 101259.6, 101131.6, 101089.2, 101095.6,
  101595.9, 101229.4, 100836, 100468.8, 100234.6, 100148, 100273.8, 100514, 
    100819.5, 100766.8, 101095.4, 101550.9, 101506.4, 101100.2, 100880.7,
  101496.4, 101055, 100627.7, 100278.2, 100031.6, 99876.52, 100190.9, 
    100437.2, 100752.3, 101099.9, 101361, 101580.8, 101632.7, 99757, 100253.7,
  101430.7, 100976, 100565, 100250.2, 99947.68, 96693.96, 100142, 100611.4, 
    100926.9, 101217.9, 101438.2, 101584.4, 101581.5, 101473.7, 101259.3,
  101489.7, 101082.6, 100747.5, 100468, 100371.3, 100110.9, 96941.76, 
    100684.2, 101174.5, 101386.1, 101542.2, 101549.3, 101477.5, 101276.4, 
    100993.1,
  101668.5, 101411.3, 101163.9, 100977.2, 100871.4, 100928.9, 100726.2, 
    95102.84, 94663.11, 101255.5, 101589.2, 101475.6, 101333.2, 101005, 
    100704.9,
  101797.5, 101672.2, 101514.7, 101389.9, 101251, 101232.3, 101344.3, 
    101257.5, 101239.3, 101573.9, 101550.2, 101408.2, 101174.9, 100816.6, 
    100630.5,
  101853.6, 101815.4, 101730.2, 101647.6, 101580.2, 101530.3, 101493.1, 
    101606.7, 101660.1, 101582.9, 101503.7, 101312.1, 101057.5, 100809.6, 
    100705,
  101860.6, 101860.1, 101827.3, 101766.5, 101682.6, 101672, 101655.5, 
    101594.4, 101585.7, 101572.5, 101449, 101217.7, 101063.6, 100940, 100855.6,
  101829.1, 101835.2, 101828.5, 101776, 101720.9, 101684.4, 101657.6, 
    101683.3, 101655.1, 101558.4, 101369.4, 101199.8, 101109, 101038.7, 
    101011.8,
  101808.8, 101762.9, 101727.9, 101698.3, 101659, 101667.5, 101646.3, 101597, 
    101556.4, 101481.7, 101347.3, 101259, 101218.9, 101195.9, 101186.2,
  102627.4, 102579.5, 102527.9, 102443.2, 102200.8, 101823, 101424.7, 
    100956.9, 100504.6, 99839.8, 99736.05, 99954.95, 99916.12, 99683.07, 
    99675.6,
  102501.1, 102464.6, 102486.2, 102422.8, 102188.7, 101618.4, 101576.9, 
    101077.2, 100654.8, 100380.2, 100257.4, 100321.7, 100368.7, 98694.68, 
    99442.49,
  102386.1, 102402.9, 102453.1, 102444.8, 102099.3, 98456.71, 101469.3, 
    101480.4, 101113.4, 100834.8, 100700.4, 100718.5, 100759.9, 100799.4, 
    100808.2,
  102269, 102324.1, 102434.3, 102418.8, 102302.6, 101834.6, 98030.23, 
    101314.6, 101292.8, 101206.6, 101075.4, 101023, 101016.4, 101038, 101004,
  102173.8, 102292.6, 102397.1, 102421.6, 102345.9, 102173.6, 101817.5, 
    95681.36, 94983.41, 101233.6, 101313.1, 101177.1, 101122, 101029.2, 
    100985.5,
  102148.5, 102247.5, 102324.5, 102389.4, 102317, 102228.8, 102125, 101924.2, 
    101576.8, 101587.3, 101417.8, 101286, 101175.2, 101085.8, 101048.2,
  102132, 102163.2, 102193.4, 102266.2, 102272.8, 102237.2, 102125.3, 
    102061.2, 101933.5, 101694.4, 101498.9, 101364.8, 101252, 101178.4, 
    101144.4,
  102074.1, 102044.3, 102024.1, 102090.4, 102120, 102163.4, 102151.8, 102056, 
    101900.1, 101744.5, 101577.9, 101441.9, 101348.1, 101290.5, 101269.4,
  102019.1, 101970.7, 101930.8, 101932.2, 101987.4, 102074.6, 102095.9, 
    102078.2, 101997.1, 101804.2, 101644.7, 101543.3, 101459.5, 101417.5, 
    101382.5,
  102000.9, 101918.1, 101851.3, 101808.1, 101847.3, 101964.8, 102071.7, 
    102026.6, 101923.8, 101768.2, 101709.5, 101652, 101577.4, 101540, 101506.5,
  102259.2, 102336.5, 102383.7, 102464.1, 102673.7, 102753.6, 102679.4, 
    102553.1, 102356.1, 101711, 101475.5, 101457.1, 101041.6, 100365.4, 
    100006.1,
  102263.3, 102297.5, 102368.7, 102517.5, 102697.7, 102529.6, 102742.1, 
    102494.5, 102292.2, 102057.5, 101768.9, 101560.9, 101289.7, 99244.57, 
    99657.34,
  102287.6, 102378.9, 102463.1, 102616.2, 102578.2, 99186.85, 102481.2, 
    102651.2, 102392.5, 102137.2, 101834.8, 101627.7, 101400.4, 101205.2, 
    100921.8,
  102374.1, 102405.3, 102513.2, 102676.6, 102734.7, 102544.6, 98837.55, 
    102255.2, 102319.2, 102173.1, 101911.3, 101677.6, 101475.2, 101297.8, 
    101085.7,
  102422.8, 102479.6, 102563.4, 102664.5, 102766.4, 102765.1, 102582.2, 
    96494.87, 95716.64, 102013, 101985, 101736.5, 101560.8, 101370.7, 101235,
  102477.6, 102521, 102521.8, 102627.3, 102646.2, 102721.8, 102721.7, 
    102586.9, 102305.2, 102262.1, 102017.9, 101794.9, 101615.7, 101452.8, 
    101301.1,
  102524.4, 102561.3, 102541.3, 102528.1, 102511.8, 102569.1, 102598.9, 
    102644.5, 102528, 102294.8, 102066, 101851.9, 101672, 101513.8, 101355.5,
  102550, 102589.8, 102565.1, 102523.6, 102421.1, 102451.9, 102535.4, 
    102579.2, 102465.4, 102317.9, 102110.7, 101914.2, 101742.6, 101577.2, 
    101408.3,
  102649, 102673.8, 102629.8, 102540.4, 102457.7, 102467.9, 102577.2, 
    102627.6, 102524.9, 102352.9, 102162.7, 101984.1, 101819.2, 101649.9, 
    101476,
  102725.1, 102720.4, 102634.7, 102537.4, 102482.2, 102532.9, 102646.4, 
    102610.6, 102483, 102330.4, 102202.8, 102055.4, 101903, 101748.7, 101582.8,
  101833, 101970.3, 102120.3, 102248.6, 102396.9, 102488.8, 102456.4, 
    102410.6, 102312, 101793.9, 101636.4, 101635.6, 101261, 100630.1, 100303.9,
  102035.4, 102151, 102319.2, 102421.3, 102537.6, 102352, 102577.3, 102386.5, 
    102265.5, 102115.4, 101889.5, 101663.5, 101410.1, 99384.85, 99838.89,
  102200.7, 102386.9, 102478.5, 102596.9, 102473.3, 99110.44, 102404.7, 
    102552.1, 102402.8, 102184.4, 101893.9, 101665, 101415.3, 101248.5, 
    101003.1,
  102372.7, 102546.1, 102624.4, 102710.7, 102723.1, 102482.6, 98773.98, 
    102214.2, 102237.7, 102191.3, 101916.9, 101665.2, 101431.1, 101257.4, 
    101060.1,
  102571, 102703.2, 102775.7, 102790.5, 102821.2, 102787.9, 102539.8, 
    96445.09, 95705.38, 101978.4, 101961.9, 101674.4, 101471.6, 101263.5, 
    101127.3,
  102688.5, 102808.8, 102842.5, 102855.9, 102797.1, 102784.7, 102746.2, 
    102578.5, 102243.2, 102211.4, 101969.4, 101720.6, 101517.6, 101316.3, 
    101161.6,
  102835.9, 102960.5, 102993.2, 102975.9, 102923.1, 102852.9, 102738.8, 
    102633.2, 102462.7, 102233.8, 101994.5, 101774.5, 101567.7, 101380, 
    101197.5,
  102971.9, 103072.8, 103106.6, 103090.4, 103018.4, 102944.3, 102820.2, 
    102626.1, 102409.2, 102245.3, 102038.4, 101829.2, 101634.8, 101454.8, 
    101257.6,
  103081.4, 103182.9, 103222.6, 103211.2, 103157.9, 103040, 102854.8, 
    102671.9, 102481.3, 102284.7, 102090.6, 101892.3, 101700.5, 101526.3, 
    101315.8,
  103191.6, 103289.8, 103310.9, 103295.9, 103221, 103100.4, 102910.2, 
    102690.3, 102488.4, 102286.9, 102148.4, 101961.3, 101773.1, 101598.6, 
    101382.2,
  102378.7, 102533.3, 102641, 102658.9, 102650.9, 102591.4, 102508.7, 
    102420.9, 102270.1, 101728.3, 101566.9, 101588.8, 101232.2, 100634.9, 
    100333.6,
  102562.6, 102680.5, 102745.9, 102750.6, 102684.9, 102428.9, 102552.3, 
    102318.9, 102133.9, 101999.6, 101792.9, 101587.4, 101366.7, 99356.46, 
    99814.4,
  102686.9, 102820.5, 102854.4, 102870.3, 102622.5, 99134.75, 102324.9, 
    102486.7, 102270.8, 102018.4, 101764.2, 101567.6, 101345.4, 101171.3, 
    100933.5,
  102769.8, 102892.9, 102940.6, 102919.4, 102848.3, 102482.1, 98689.25, 
    101991.1, 102018.7, 101998.7, 101748.2, 101524.4, 101309.1, 101122.2, 
    100896.9,
  102843.5, 102982.3, 103014.8, 102981.5, 102880.9, 102740.8, 102397, 
    96307.66, 95506.45, 101721.6, 101744.3, 101469.1, 101259.1, 101024.1, 
    100840.8,
  102908.5, 103038, 103070.6, 103036.9, 102882, 102725, 102552.3, 102296.7, 
    101956.1, 101935.2, 101697.1, 101439.4, 101204.5, 100963.9, 100754.2,
  102980.9, 103134.6, 103152.1, 103077.8, 102924.3, 102737.1, 102530, 
    102387.3, 102182.1, 101925.1, 101682.3, 101427.3, 101166.1, 100934.9, 
    100709.9,
  103061.1, 103183.7, 103184.1, 103096.1, 102925.5, 102746.6, 102544.6, 
    102324.8, 102107.6, 101922.2, 101698.9, 101432.8, 101183.5, 100951.3, 
    100731.9,
  103160.2, 103250.3, 103235.8, 103136.9, 102987.4, 102784.6, 102583.4, 
    102399.4, 102189.5, 101959.9, 101731.2, 101482.1, 101233.7, 101008.6, 
    100792.7,
  103243.3, 103282, 103240.3, 103141.8, 102996.5, 102808.3, 102614.3, 
    102387.3, 102166.4, 101950.6, 101779.5, 101555.3, 101323.5, 101111.8, 
    100906.5,
  102545.3, 102625.7, 102651.2, 102601.7, 102535.5, 102438.8, 102322.2, 
    102220.7, 102098.2, 101613.5, 101523.3, 101610.2, 101284.3, 100687.3, 
    100407.2,
  102689.2, 102724.3, 102715, 102639.9, 102524.4, 102193.9, 102327.1, 
    102080.5, 101923.9, 101850.4, 101693.2, 101539.8, 101326.9, 99316.32, 
    99790.8,
  102762.4, 102809.8, 102767.3, 102707.3, 102425.2, 98894.34, 102043, 
    102208.3, 102007.3, 101831.7, 101627.5, 101437.6, 101207.8, 101034.5, 
    100842.6,
  102808.4, 102854.1, 102797.8, 102705.6, 102576.9, 102202.9, 98410.48, 
    101716.9, 101810.7, 101773.1, 101565.7, 101331.2, 101118.9, 100949.9, 
    100773.9,
  102860.1, 102889.5, 102833.2, 102739.1, 102590.9, 102429.6, 102090.1, 
    96032.2, 95217.23, 101489.6, 101517.2, 101243, 101051.5, 100875.7, 
    100754.5,
  102886.3, 102911, 102841.1, 102738.6, 102548.3, 102392, 102222, 101976.9, 
    101648.9, 101655.6, 101422.6, 101188, 101014.5, 100854.9, 100709.7,
  102908, 102930.6, 102850.8, 102737.7, 102565.8, 102363.7, 102152.3, 
    101993.4, 101793.4, 101560.4, 101343.8, 101148.6, 100978.2, 100828.2, 
    100669.4,
  102933, 102915.8, 102824.4, 102694.2, 102508, 102317.1, 102089.7, 101844.1, 
    101631.3, 101468, 101280.9, 101110.9, 100960.6, 100807.2, 100645.2,
  102965.8, 102918, 102807.1, 102679.3, 102520.8, 102286.6, 102034.1, 101808, 
    101600, 101389.7, 101214.2, 101069.5, 100925.9, 100784.2, 100623.2,
  102981.1, 102881.7, 102743.5, 102621.3, 102441.4, 102220.8, 101962.7, 
    101681.3, 101446, 101249.8, 101135.1, 101022.7, 100894, 100769.2, 100616.7,
  102739.4, 102803.9, 102785.6, 102696, 102591.6, 102456.5, 102310.8, 
    102202.3, 102095.1, 101622.5, 101590.9, 101749.5, 101507.2, 100990.6, 
    100755,
  102827.7, 102825.4, 102777.6, 102676.7, 102529.8, 102164.8, 102290.9, 
    102022.3, 101866.8, 101826.2, 101742.1, 101690.3, 101597.1, 99667.88, 
    100217.5,
  102843.3, 102848.2, 102758.8, 102667.2, 102360.8, 98842.12, 101899.6, 
    102105.2, 101873.7, 101709.4, 101610, 101584, 101512, 101463.5, 101343.9,
  102835.9, 102819.2, 102711.7, 102570, 102425.3, 102019, 98253.02, 101427, 
    101549, 101560, 101473.2, 101419.8, 101389.6, 101372.6, 101314.6,
  102835.5, 102786.9, 102657.9, 102504, 102336.7, 102138.1, 101758.1, 
    95761.35, 94883.77, 101118.8, 101322.9, 101240.8, 101239, 101215.6, 
    101234.5,
  102790.9, 102722.8, 102563.9, 102415.5, 102194.3, 101996.9, 101769.3, 
    101463.5, 101135.2, 101195.9, 101093, 101046.2, 101052.6, 101060.6, 
    101094.8,
  102746.4, 102668.3, 102506.2, 102351, 102149.3, 101890.1, 101623.1, 
    101413.5, 101191.5, 100987.6, 100887.7, 100857, 100851.5, 100881.6, 
    100923.3,
  102713.9, 102601.3, 102436.7, 102277.5, 102055.6, 101813, 101536.1, 
    101245.3, 101015.6, 100876.9, 100764.1, 100695.4, 100688.3, 100719.3, 
    100770.2,
  102706.8, 102580.5, 102433.3, 102273.7, 102070.2, 101792.6, 101505.6, 
    101255.8, 101018.9, 100816.3, 100675.2, 100599.9, 100562.8, 100569.9, 
    100614,
  102716.8, 102552.4, 102399.1, 102247.1, 102044, 101792.2, 101524.6, 
    101236.8, 100989.2, 100778.3, 100658.2, 100558.8, 100494.2, 100480.8, 
    100498.5,
  102197.2, 102317.1, 102352, 102277.3, 102161, 102027.9, 101877.3, 101781.4, 
    101703.3, 101268.9, 101286.1, 101546.2, 101420.9, 101053, 100899,
  102314.2, 102356.9, 102312.4, 102194, 102044.4, 101695.4, 101810.5, 
    101580.7, 101453.5, 101427.5, 101385.9, 101438.2, 101504.9, 99724.75, 
    100390.6,
  102352.7, 102356.5, 102244.2, 102148.5, 101847.9, 98380.82, 101438.4, 
    101608.8, 101399.5, 101287.2, 101245.7, 101294.9, 101406.8, 101505.2, 
    101543.6,
  102350, 102304.4, 102188.9, 102057.5, 101913.6, 101535.9, 97814.47, 
    101063.8, 101206.1, 101196.2, 101152, 101171, 101286.1, 101445, 101551.5,
  102353.8, 102277.1, 102173, 102039, 101874.5, 101669.4, 101336.9, 95409.26, 
    94594.52, 100873, 101068.6, 101054.4, 101178.8, 101323.4, 101527.5,
  102315.6, 102255.9, 102151.6, 102008.5, 101764.5, 101563.8, 101359.6, 
    101136.2, 100901.3, 101016.7, 100955.3, 100965.5, 101069.4, 101251.3, 
    101459.5,
  102313.5, 102277, 102180.8, 102002.5, 101761.7, 101482.8, 101236.9, 
    101094.4, 100990.3, 100905.5, 100861.4, 100889.1, 100983.8, 101179.3, 
    101395.6,
  102337.3, 102280.8, 102178.1, 101969, 101688.4, 101413.9, 101142.2, 
    100913.9, 100819.4, 100828.3, 100795.9, 100828.4, 100929.8, 101135.6, 
    101365.8,
  102375.3, 102325.8, 102222.4, 102020.1, 101747.8, 101419.5, 101105.4, 
    100886.1, 100774.8, 100752.6, 100732.6, 100790.6, 100910, 101119.4, 
    101350.7,
  102417, 102338.6, 102222, 102020.3, 101729.8, 101436.1, 101123.3, 100835.9, 
    100671.6, 100638.4, 100695.7, 100765.4, 100930.2, 101144, 101366.1,
  101463.9, 101510.6, 101502.7, 101430.9, 101366.5, 101287.7, 101197.1, 
    101183.2, 101216.3, 100906.8, 101026.6, 101369.9, 101317, 100971.5, 
    100816.5,
  101600.9, 101564.3, 101508.9, 101415.9, 101309.3, 100984.9, 101164, 
    101066.6, 101077.2, 101144.1, 101206.3, 101353.4, 101482.9, 99731.84, 
    100406,
  101639.7, 101584.6, 101498.5, 101408.9, 101116, 97678.57, 100791, 101041.7, 
    101013.2, 101096.9, 101171.3, 101331.5, 101514.8, 101609.4, 101624.1,
  101650.6, 101586.2, 101487.5, 101339.7, 101148.2, 100798.6, 97138.27, 
    100625.9, 100940.7, 101034.7, 101168.8, 101321.4, 101526.7, 101687.4, 
    101748.6,
  101667.2, 101603.9, 101486, 101292.4, 101092.6, 100885.2, 100649.7, 
    94860.59, 94341.12, 100818.5, 101201.4, 101346.1, 101570.7, 101706.1, 
    101839.8,
  101680.6, 101618.9, 101473.6, 101282.8, 101023.9, 100849.4, 100724.9, 
    100722.9, 100676, 101064.3, 101213.8, 101409.4, 101617.4, 101796.2, 
    101913.1,
  101713, 101660.9, 101512.4, 101320.6, 101104.5, 100914.8, 100784.1, 
    100845.7, 101003.2, 101141.3, 101292.9, 101489.4, 101682, 101869.4, 
    101995.1,
  101759.7, 101704.4, 101569.6, 101398.1, 101198.4, 101048.8, 100959.1, 
    100970.3, 101085.1, 101251.1, 101392.6, 101576.6, 101779, 101969.4, 
    102114.4,
  101836, 101794.9, 101681.4, 101532, 101382.1, 101247.4, 101168.7, 101206.3, 
    101293.7, 101386.8, 101510.3, 101690.7, 101888.7, 102073.1, 102211.9,
  101924, 101876.4, 101786.7, 101657.2, 101514.8, 101419.8, 101368.2, 
    101363.1, 101404.2, 101465.1, 101631.3, 101820.6, 102017.9, 102196.3, 
    102326.1,
  101312.4, 101355.5, 101349.5, 101294.5, 101245.3, 101189.4, 101130.8, 
    101160.5, 101208.1, 100926.8, 101063.5, 101387.3, 101252.7, 100801.9, 
    100519.9,
  101341.6, 101325.7, 101315.5, 101242.1, 101171.1, 100891.9, 101073.8, 
    101053.6, 101116.6, 101210.6, 101306.1, 101434.8, 101436.2, 99557.81, 
    100081.8,
  101308.2, 101301.8, 101267.7, 101211.6, 100986.6, 97581.09, 100830.6, 
    101059.8, 101143.9, 101230.4, 101322.4, 101451.5, 101482.6, 101445.3, 
    101250.9,
  101267.4, 101295.6, 101246.7, 101170.8, 101044.4, 100817, 97192.12, 
    100859.1, 101113.1, 101237.5, 101381.5, 101479, 101522.8, 101485, 101334.2,
  101282.9, 101313.2, 101263.1, 101152.5, 101061.9, 100999.1, 100872.9, 
    95116.43, 94628.09, 101109.4, 101454.1, 101517.8, 101551.5, 101475.9, 
    101421.2,
  101317, 101356.7, 101302.7, 101214.6, 101094.8, 101041.5, 101053.8, 
    101089.3, 101017.4, 101395.7, 101506.1, 101592.8, 101597.6, 101566.4, 
    101512,
  101368.6, 101436.5, 101386.3, 101323.9, 101245, 101213.8, 101197.9, 
    101314.3, 101442.2, 101523.4, 101611.9, 101673.7, 101688.6, 101695.1, 
    101675,
  101464.8, 101522.1, 101495.1, 101449.3, 101383.6, 101371, 101390.2, 
    101436.2, 101521.5, 101658, 101756.2, 101818.9, 101863.6, 101880, 101873.9,
  101579.3, 101626.4, 101617.6, 101592, 101573.4, 101569.7, 101592.8, 
    101686.6, 101782.8, 101872, 101946, 102017.2, 102049.1, 102069, 102050.6,
  101703.1, 101737.1, 101739.7, 101733.9, 101724.2, 101748.4, 101799.7, 
    101851.7, 101923.8, 102004.1, 102138.2, 102222.4, 102260, 102292.5, 102268,
  100584.6, 100766.2, 100936.7, 101082.4, 101240.6, 101345.9, 101396.4, 
    101475.2, 101512.3, 101176.1, 101229.3, 101535.7, 101366.2, 100875.7, 
    100573.7,
  100686.9, 100855.5, 101021.3, 101148.5, 101237.5, 101127.9, 101364, 
    101386.9, 101436.3, 101502.7, 101500.5, 101585, 101546.3, 99638.54, 
    100117.3,
  100770.9, 100962.6, 101091.4, 101202.4, 101131, 97799.85, 101121, 101396.9, 
    101417, 101497, 101517.8, 101576.1, 101560.7, 101480.2, 101259,
  100860.4, 101052.9, 101128.6, 101206.6, 101217.9, 101063.3, 97465.11, 
    101076.2, 101392.7, 101454, 101516.7, 101539.9, 101533.2, 101444.6, 
    101248.2,
  100980.1, 101133.1, 101182.8, 101203.7, 101225.2, 101240.2, 101089.1, 
    95349.53, 94737.65, 101215.1, 101494.9, 101499.4, 101470.9, 101333.4, 
    101217.7,
  101109.8, 101217.2, 101223.9, 101231.2, 101155.3, 101181, 101220.6, 101207, 
    101110.2, 101408.1, 101438.7, 101449.1, 101392.7, 101270.5, 101193.3,
  101242.4, 101305.2, 101308.7, 101289.9, 101264.2, 101244.1, 101249.3, 
    101343.4, 101381, 101391.7, 101417.8, 101402.8, 101315.3, 101257.7, 
    101241.5,
  101357.2, 101394.1, 101378.1, 101346.1, 101300.8, 101313.1, 101322.8, 
    101319.9, 101320.8, 101354.9, 101357.4, 101341.4, 101319.3, 101333.2, 
    101360.2,
  101484.9, 101507.5, 101486, 101451, 101423.6, 101391.7, 101371.4, 101395.2, 
    101392.4, 101361.8, 101348.7, 101364.2, 101386.5, 101435.5, 101482.9,
  101637.7, 101642.9, 101618.7, 101564.9, 101499.6, 101475.9, 101466.3, 
    101441.8, 101401.5, 101371.4, 101426.5, 101470.4, 101517.1, 101585.6, 
    101640.8,
  99784.87, 99978.18, 100173.3, 100477.2, 100802.9, 101098.9, 101370.5, 
    101584.5, 101747.9, 101488.9, 101593, 101841.3, 101625.4, 101152.5, 
    100864.9,
  99882.52, 100080.4, 100322.7, 100653.7, 100948, 101118, 101488.6, 101670.8, 
    101775.4, 101877.7, 101878.3, 101923.8, 101849.3, 99891.12, 100352.3,
  100059, 100279.6, 100524.7, 100825.1, 100931.1, 97921.99, 101442.1, 101820, 
    101865.6, 101934, 101953.7, 101918.4, 101843.6, 101722.2, 101460.7,
  100301.1, 100517.3, 100726.6, 100961, 101175.8, 101105.3, 97816.82, 
    101478.3, 101846.7, 101920.3, 101926, 101876.1, 101802.3, 101648, 101372.2,
  100586.9, 100760.7, 100930.3, 101114, 101302.7, 101480.7, 101351.4, 
    95775.01, 95137.41, 101638.5, 101886.8, 101832.2, 101742.9, 101514.3, 
    101331.1,
  100852.1, 100976, 101078, 101226, 101306.9, 101459.4, 101604.5, 101574.5, 
    101552.2, 101812.1, 101834.7, 101798.5, 101651.7, 101442.7, 101298.6,
  101069.4, 101152.7, 101221.7, 101296.2, 101390.5, 101466.5, 101562.9, 
    101725.9, 101794.8, 101808.9, 101836.2, 101749.9, 101559.3, 101418.9, 
    101367.8,
  101190.8, 101232.3, 101281.8, 101332.2, 101362.5, 101468.5, 101571.8, 
    101654.7, 101773.4, 101849.7, 101801.1, 101668.3, 101530.1, 101489.8, 
    101495.9,
  101247.4, 101283.1, 101308.9, 101345.5, 101405.8, 101476, 101579.8, 
    101718.9, 101820.4, 101799.2, 101733.2, 101622.6, 101581, 101596.4, 
    101632.2,
  101296.2, 101269.5, 101271.4, 101304.1, 101349.6, 101451.9, 101572.1, 
    101658, 101715.2, 101695.5, 101665.6, 101653.9, 101673, 101741.7, 101816.2,
  99731.52, 99891.48, 100076.9, 100314.5, 100573.1, 100858, 101200.4, 
    101488.7, 101759, 101628, 101865.1, 102204.2, 102092, 101677.7, 101480,
  99728.07, 99909.41, 100128.7, 100440.5, 100732.3, 100940.1, 101400.3, 
    101673.8, 101865.8, 102096.3, 102238.6, 102342.6, 102337.3, 100418.9, 
    100995.6,
  99741.09, 99963.86, 100242.2, 100593.1, 100741.7, 97939.48, 101533.4, 
    101933.4, 102134.2, 102257.6, 102348.2, 102378.6, 102349.4, 102285.4, 
    102130.8,
  99794.8, 100051, 100377.7, 100705, 101046.6, 101052, 98035.19, 101790.4, 
    102220.4, 102323, 102367.9, 102352.3, 102291, 102167.4, 102039.9,
  99919.41, 100200.9, 100542.1, 100893.7, 101234.4, 101623.4, 101542.2, 
    96093.52, 95571.13, 102115.8, 102369.6, 102289.4, 102174, 101992.8, 
    101925.8,
  100109, 100388.8, 100710.4, 101078, 101382.2, 101714.7, 101967.6, 101954.2, 
    102022, 102336.8, 102358.3, 102219.6, 102042.4, 101886.7, 101824.6,
  100374.4, 100635.9, 100940.9, 101266.3, 101582.1, 101844.6, 102040.1, 
    102288.9, 102406.5, 102408.3, 102330.5, 102150.9, 101988.3, 101880.1, 
    101850,
  100669.8, 100897.6, 101170.3, 101450.6, 101723.6, 101967.2, 102164.2, 
    102292.7, 102388, 102415, 102290.2, 102118.2, 102019.1, 101962.5, 101959.2,
  100958.9, 101184.7, 101426.9, 101671.1, 101898.5, 102115, 102305.6, 
    102452.3, 102519.1, 102412.3, 102274.3, 102140.8, 102072.5, 102050.2, 
    102050.4,
  101183, 101369.2, 101590.4, 101815.8, 102025.4, 102224.5, 102395.4, 
    102460.3, 102458, 102362.6, 102257.7, 102173.1, 102151.4, 102157.2, 
    102177.6,
  99498.84, 99540.32, 99690.33, 99911.15, 100177.7, 100435.4, 100699, 
    100991.4, 101303.4, 101290.6, 101641.5, 102119.7, 102142.9, 101853.2, 
    101701.5,
  99416.8, 99465.38, 99643.88, 99911.36, 100188.5, 100360.5, 100779.7, 
    101088.6, 101363.7, 101696, 101964.5, 102232.4, 102354.5, 100597.8, 
    101250.7,
  99454.24, 99553.34, 99754.52, 100047.6, 100191.4, 97389.22, 100920, 
    101355.1, 101620.6, 101864.8, 102092.5, 102302.5, 102422.4, 102482.5, 
    102451.5,
  99645.58, 99756.89, 99977.18, 100223.8, 100539.1, 100538.1, 97604.85, 
    101321.4, 101812.3, 102033.6, 102205.7, 102337.1, 102431.8, 102459.1, 
    102432.8,
  99883.91, 100042.9, 100260.7, 100530.7, 100813.6, 101176.7, 101068.6, 
    95778.59, 95353.21, 101886.8, 102297.6, 102324.5, 102358.8, 102287, 
    102287.7,
  100135.6, 100322, 100526.2, 100816.1, 101051.3, 101327.5, 101537, 101499.9, 
    101617.8, 102157.8, 102239.8, 102262.3, 102203.4, 102116, 102085.6,
  100353.2, 100582, 100822.2, 101079.5, 101345, 101575.6, 101739.3, 102010.7, 
    102179.4, 102189.7, 102204.1, 102168.5, 102087.1, 102044.2, 102046.5,
  100572.8, 100830.6, 101073.6, 101342.1, 101553.6, 101783.4, 101936.7, 
    102024.7, 102112.5, 102198.8, 102180.1, 102151, 102108.2, 102098.1, 
    102117.8,
  100812.1, 101106.8, 101402.6, 101663.3, 101875.3, 102040.2, 102171.6, 
    102284.6, 102307.5, 102257, 102230.6, 102193.7, 102155.6, 102147.7, 
    102151.7,
  101088.8, 101377.4, 101647.8, 101883.8, 102078.4, 102231.7, 102317.2, 
    102322.2, 102314.8, 102284.2, 102299.1, 102264, 102226.5, 102237.5, 
    102266.5,
  100085.2, 100252.1, 100392.1, 100534.5, 100526.9, 100552.3, 100575.1, 
    100613.8, 100703.3, 100607.2, 100936.1, 101490.8, 101660.2, 101486.9, 
    101462.5,
  99837.4, 100043, 100260.1, 100453.3, 100512.7, 100464.5, 100670.9, 
    100671.7, 100727, 100931.8, 101195, 101529.7, 101838.8, 100269.2, 101044.4,
  99583.05, 99854.16, 100141.8, 100395.8, 100423.2, 97317.74, 100583.8, 
    100787.1, 100827.7, 100954.1, 101233.6, 101551.9, 101886.3, 102072.9, 
    102259.3,
  99487.93, 99753.48, 100068.7, 100302.8, 100531.6, 100391.9, 97119.81, 
    100541.5, 100870.5, 101021.9, 101289.6, 101593.7, 101942.3, 102189.7, 
    102356.9,
  99647.86, 99857.3, 100104.9, 100340.2, 100528.6, 100713.7, 100575.7, 95100, 
    94601.23, 100930, 101397.3, 101661.9, 101983, 102180.7, 102375.9,
  99931.93, 100077.6, 100235.4, 100435.4, 100562.9, 100696.4, 100823.5, 
    100769.9, 100779.4, 101265.3, 101491.6, 101775.2, 102049.9, 102225.2, 
    102344.9,
  100271.8, 100364.1, 100470.7, 100610, 100731.7, 100850.9, 100954.2, 
    101178.8, 101359.8, 101471.8, 101685.7, 101918, 102074.2, 102184.8, 
    102252.5,
  100623.2, 100683.9, 100759.1, 100867.2, 100971.2, 101105.6, 101230.5, 
    101343, 101498.5, 101693, 101860.5, 101986.9, 102092.8, 102172.7, 102220.8,
  100977.3, 101051.1, 101128.2, 101221.3, 101321.4, 101427.5, 101543.1, 
    101686.3, 101801.1, 101879.5, 101965.2, 102047.5, 102111.5, 102168.4, 
    102177.1,
  101295.9, 101361.4, 101436.2, 101517.8, 101603.6, 101703.7, 101793.7, 
    101855.1, 101911.7, 101965.3, 102063.6, 102133, 102199.5, 102246.3, 
    102221.6,
  100281.9, 100398.7, 100434.2, 100493.5, 100458, 100391.4, 100417.3, 
    100509.5, 100686.2, 100502.1, 100695.2, 101081.3, 101144, 100953.5, 
    100959.6,
  100365.1, 100445.3, 100467.3, 100481.6, 100338, 100108.2, 100286.9, 
    100388.9, 100527.5, 100714.9, 100914.1, 101151.5, 101354.7, 99800.48, 
    100588.6,
  100470.2, 100503.7, 100485.9, 100452.4, 100140.1, 96855.13, 100087.9, 
    100366.5, 100541.4, 100696, 100916.5, 101172.6, 101445.5, 101613.4, 
    101824.3,
  100550.3, 100538.9, 100507, 100375.7, 100283.6, 99891.65, 96655.41, 
    100097.8, 100483.6, 100670.7, 100944.6, 101207.8, 101529.4, 101803, 
    102008.4,
  100633, 100600.1, 100526.8, 100423.3, 100273.9, 100308.7, 100029, 94661.88, 
    94225.52, 100501.9, 101006.6, 101266.5, 101596.8, 101841.1, 102117.6,
  100726.4, 100689.4, 100596.2, 100511.7, 100377.8, 100339.4, 100459.8, 
    100372.7, 100298.5, 100785.5, 101037.9, 101357.5, 101676.5, 101956.7, 
    102202.9,
  100850.4, 100810.6, 100737.9, 100640.7, 100561.5, 100507.2, 100505.3, 
    100673.4, 100805.7, 100905, 101148.8, 101472.9, 101780.8, 102056.1, 
    102266.6,
  101017.7, 100994.1, 100933.1, 100869.7, 100793.3, 100774.8, 100788.4, 
    100796.9, 100894.9, 101114.5, 101373.1, 101653.8, 101927.1, 102174.4, 
    102372.1,
  101274.7, 101275.8, 101252.4, 101217.2, 101186.8, 101158.7, 101173.8, 
    101261.9, 101358.4, 101462.9, 101638, 101859.3, 102077.9, 102277.9, 
    102435.6,
  101555.4, 101557.8, 101554.5, 101535.3, 101515.5, 101516, 101526.2, 
    101532.8, 101589.6, 101691.6, 101881.9, 102054.1, 102216.3, 102371.9, 
    102494.8,
  100870.9, 100800.7, 100735.2, 100731.2, 100781, 100861, 100939.9, 101079.4, 
    101236.3, 101086.4, 101146.4, 101393.4, 101308.4, 101085.1, 101062.1,
  100825.7, 100698.7, 100615.4, 100617.6, 100619.6, 100600.5, 100879.5, 
    100982.3, 101121.9, 101365.4, 101399.2, 101449.4, 101487.2, 99893.2, 
    100640.5,
  100701.2, 100515.7, 100412.6, 100407.3, 100384.5, 97252.24, 100637, 
    101027.7, 101184.6, 101357.4, 101410.7, 101469.2, 101551.8, 101654.2, 
    101794.3,
  100590.2, 100349.1, 100183.4, 100102.9, 100270.5, 100195.5, 97044.02, 
    100624.8, 101087.5, 101337.1, 101434.1, 101476.7, 101574.9, 101742.4, 
    101922.5,
  100507.8, 100204.1, 99935.44, 99800.12, 99932.91, 100318.4, 100295.7, 
    95090.31, 94688.66, 101053.1, 101438.4, 101493.9, 101597.8, 101736.7, 
    101997.5,
  100488.7, 100119.1, 99761.2, 99542.89, 99644.96, 100059.7, 100479.5, 
    100577.1, 100662.1, 101247, 101364.4, 101496.1, 101628.5, 101803.2, 
    102060.5,
  100553.1, 100158.3, 99775.06, 99536.68, 99627.58, 100017.7, 100377.3, 
    100810.7, 101077.8, 101205.7, 101332.4, 101502.1, 101654, 101848.6, 
    102094.3,
  100711.3, 100336.1, 99953.31, 99715.39, 99765.62, 100113.8, 100429.7, 
    100659.2, 100880, 101161, 101341.1, 101520.1, 101712.8, 101925.2, 102185.7,
  100948.6, 100632.8, 100309.5, 100106.3, 100127.4, 100327, 100564.5, 
    100856.5, 101072.3, 101235.9, 101385.4, 101579.3, 101782.5, 102016.1, 
    102266.3,
  101215.8, 100967.9, 100696.3, 100511.7, 100481.4, 100603.8, 100762.8, 
    100913.7, 101070.9, 101254.8, 101469.8, 101677.4, 101893.7, 102144.7, 
    102358.9,
  101538.9, 101510.4, 101470.2, 101415.4, 101379.1, 101327.8, 101271.7, 
    101237.8, 101190.2, 100857.3, 100882.5, 101112.5, 100943.4, 100581.6, 
    100484.9,
  101450, 101364.8, 101301.8, 101234.8, 101173.5, 100992.3, 101171.4, 
    101104.1, 101046, 101090.6, 101079.9, 101090.7, 101079.1, 99362.9, 
    100059.2,
  101276.9, 101159, 101067.1, 101003.5, 100870.1, 97574.2, 100821.9, 
    101092.1, 101040.6, 101038.9, 101051, 101038, 101085.4, 101139.3, 101248.2,
  101089.3, 100924.4, 100791.3, 100709.5, 100730.1, 100586.5, 97187.71, 
    100636.3, 100916.5, 100992.6, 101037, 100998, 101086.9, 101228.3, 101415.9,
  100869.7, 100667, 100492, 100422.9, 100449.6, 100599.1, 100538.4, 95047.64, 
    94478.2, 100732.5, 101033, 100987, 101117.2, 101278.7, 101568.7,
  100660, 100404.2, 100182, 100108.3, 100156.9, 100339.2, 100604.6, 100651.3, 
    100582.8, 100958.8, 100973, 101015.6, 101183.4, 101406.8, 101677,
  100486.8, 100182.1, 99915.42, 99842.87, 99958.57, 100184, 100458.7, 
    100773.6, 100901.2, 100955.3, 100971.4, 101085.4, 101267.5, 101494.1, 
    101758.2,
  100405.2, 100066.2, 99777.13, 99684.27, 99828.88, 100134.6, 100437.8, 
    100650.3, 100780.3, 100965.2, 101033.4, 101172.4, 101374, 101607, 101888.4,
  100442.7, 100131.4, 99868.57, 99805.91, 99963.35, 100229.9, 100503.5, 
    100745.6, 100923.1, 101037.6, 101126.6, 101281.6, 101482, 101730.8, 
    102001.2,
  100589.2, 100340.1, 100145.2, 100088.7, 100197.9, 100405.4, 100623.4, 
    100791.4, 100956.8, 101069.3, 101226.7, 101394.4, 101596.1, 101859.9, 
    102101.9,
  101536.8, 101595, 101651.8, 101697.7, 101768.9, 101794.5, 101813, 101836.1, 
    101848.9, 101491, 101487.6, 101632.9, 101364, 100796.5, 100469.2,
  101464.8, 101495.7, 101533.9, 101565.4, 101584, 101446.9, 101665.7, 
    101624.4, 101588.2, 101618.8, 101564.2, 101522.6, 101417.1, 99498.52, 
    99951.44,
  101432.1, 101435.6, 101426.2, 101428.5, 101313.9, 98050.13, 101229, 
    101538.2, 101444.6, 101424.9, 101383.8, 101367.3, 101297.5, 101218.9, 
    101056.5,
  101371.2, 101299, 101221.9, 101164.7, 101157.4, 100985.6, 97541.16, 
    100923.6, 101236.8, 101242.8, 101228.6, 101194.4, 101178.5, 101137.4, 
    101068.6,
  101184.8, 101056.6, 100928.9, 100847.6, 100840.3, 100908.9, 100820, 
    95263.77, 94535.41, 100845.7, 101098.6, 101075.5, 101076, 101043, 101102.4,
  100966.5, 100783.3, 100608.5, 100514.5, 100483.9, 100567.4, 100737.2, 
    100763.7, 100762.6, 101033.4, 101018.8, 101011.8, 100997.1, 101044.2, 
    101141.2,
  100760.6, 100554.2, 100375.7, 100254.7, 100247, 100332.2, 100489, 100731.1, 
    100871.1, 100881.1, 100908, 100900.1, 100946.8, 101064.6, 101236.2,
  100641.7, 100442.2, 100237, 100097.1, 100065.1, 100193.9, 100369, 100535.4, 
    100673.7, 100781.1, 100786.3, 100837.7, 100975.3, 101168.5, 101419.7,
  100620.5, 100436.4, 100257.8, 100145.6, 100146.1, 100227.6, 100382.7, 
    100560.1, 100653.9, 100678, 100723.8, 100885.9, 101089.3, 101346.7, 
    101596.5,
  100674.2, 100506.5, 100350.3, 100254.9, 100243.4, 100326.9, 100438.3, 
    100514.1, 100556.3, 100595.3, 100787.4, 101024.4, 101271.3, 101540.4, 
    101763.1,
  100524.3, 100731.4, 100935, 101139.3, 101342, 101502.1, 101676.1, 101855.2, 
    101988.6, 101746.2, 101896.1, 102168.3, 101989.8, 101411.2, 101014.7,
  100529.4, 100727.6, 100921.6, 101129.1, 101306.6, 101362.6, 101690.6, 
    101810.6, 101934.9, 102086.4, 102140.6, 102167.1, 102065.3, 100097.2, 
    100424.4,
  100647.7, 100841.9, 101006.7, 101187.3, 101206.2, 98168.18, 101502.4, 
    101902.6, 101943.3, 102025.2, 102078, 102084.4, 102019.6, 101836.3, 
    101503.6,
  100938.5, 101013.9, 101118.8, 101230.8, 101356.5, 101233.5, 97965.94, 
    101429.9, 101872.4, 101964.3, 102030.3, 101989.3, 101972.2, 101824.4, 
    101534.8,
  101132.1, 101147.2, 101181.2, 101244, 101319.2, 101442.3, 101329.5, 
    95872.95, 95229.05, 101599.6, 101941.3, 101919.2, 101957.2, 101809.3, 
    101658.9,
  101139.8, 101121.6, 101113.1, 101146.2, 101170.1, 101246, 101379, 101372.5, 
    101408.3, 101780.6, 101839, 101948.8, 101988.8, 101867.4, 101739.6,
  101066.8, 101024.3, 100993.6, 100994.6, 101025.1, 101072.1, 101156, 
    101377.2, 101557.6, 101666.6, 101802.5, 101956.6, 101986.1, 101922.1, 
    101886.8,
  100953.7, 100887.2, 100820.7, 100805, 100794.1, 100855.4, 100955.7, 
    101090.2, 101317.1, 101574.9, 101764.9, 101938.9, 102005.6, 102005.9, 
    102053.3,
  100845.4, 100750.8, 100667, 100622.1, 100632.5, 100678.6, 100799.5, 101020, 
    101265.1, 101504.4, 101727, 101935.4, 102011.6, 102093.5, 102193.5,
  100731.8, 100566.5, 100448.9, 100424.8, 100473, 100550.5, 100691.4, 
    100887.2, 101155, 101419.5, 101703.8, 101924.4, 102032.4, 102197.9, 
    102327.3,
  100310.5, 100026.7, 99920.98, 99953.88, 100034.6, 100207.8, 100533.8, 
    100878.9, 101208.2, 101180.4, 101525.9, 101957.6, 101896.6, 101469, 
    101215.4,
  100283.8, 100006.5, 99962.85, 100069.2, 100181.4, 100266.9, 100716, 
    101020.2, 101295.5, 101630.1, 101895.9, 102092.6, 102132.7, 100249.5, 
    100764,
  100350.6, 100084, 100060.3, 100220.9, 100256.4, 97364.22, 100841.5, 
    101242.4, 101541.5, 101811.1, 102029.6, 102175.5, 102213, 102127.6, 
    101945.2,
  100533.5, 100213, 100186.9, 100325.9, 100584, 100522.7, 97535.45, 101190.1, 
    101720.8, 101955.4, 102148.1, 102210.9, 102265.7, 102173.5, 102050.9,
  100791, 100432.6, 100336.7, 100500, 100709.5, 101024.3, 101005.7, 95774.62, 
    95384.93, 101835.8, 102230.3, 102263.4, 102310.2, 102221.7, 102202.8,
  101024, 100747, 100559.2, 100694, 100858.5, 101093.6, 101387, 101440.4, 
    101555.2, 102090.6, 102235.8, 102347.4, 102353.9, 102330.7, 102312.7,
  101140.4, 101003.5, 100837, 100897.8, 101048, 101265.1, 101469.6, 101768.4, 
    102006.4, 102141.7, 102296.6, 102417.1, 102432.9, 102467.9, 102480.2,
  101188.5, 101176.8, 101052.6, 101084.1, 101176.1, 101364, 101557.9, 
    101724.4, 101930.5, 102194.9, 102364.3, 102479, 102541.8, 102605.8, 
    102640.5,
  101182.6, 101216.3, 101193, 101202.4, 101287.5, 101439.5, 101627.5, 
    101866.6, 102087.5, 102277.5, 102409.6, 102551.3, 102626.9, 102713.1, 
    102750.3,
  101124.8, 101146.7, 101184.5, 101229, 101314.6, 101459.2, 101647.1, 
    101843.3, 102049.7, 102244.6, 102445.2, 102614.7, 102712.3, 102819.3, 
    102864.9,
  101630.9, 101345.1, 100934.2, 100604, 100380.8, 100376.3, 100438.9, 
    100574.3, 100771.2, 100651.7, 100928.5, 101357.5, 101371.3, 101096.4, 
    101004,
  101642.1, 101369, 101026.7, 100798.7, 100618.6, 100467.5, 100729.5, 
    100859.2, 101020.9, 101229.3, 101417.1, 101617, 101705.9, 99981.74, 
    100673.6,
  101607.6, 101413.9, 101144.7, 101033.1, 100779, 97644.89, 100981, 101256.5, 
    101419.4, 101544.1, 101686.2, 101830.1, 101925.4, 101966.7, 101956.5,
  101565.6, 101446.4, 101236.6, 101175.1, 101233, 100973.5, 97761.55, 
    101328.4, 101644.5, 101797.4, 101919.3, 101991.9, 102079.9, 102130.1, 
    102126.1,
  101514.7, 101464.6, 101291.2, 101304.3, 101381.3, 101554.3, 101335.5, 
    95817.59, 95386.42, 101816.6, 102137.4, 102166.5, 102262.4, 102276.7, 
    102326.5,
  101459.8, 101440.4, 101277.5, 101354.3, 101423, 101557.1, 101694.3, 
    101669.2, 101683.7, 102135.6, 102237.2, 102343.4, 102412, 102457.6, 
    102476.5,
  101415.4, 101418.4, 101272.9, 101334.3, 101483.1, 101648.3, 101740.8, 
    102001.3, 102197.7, 102281.7, 102387.2, 102498.4, 102565.3, 102612.4, 
    102611.5,
  101390.9, 101382.3, 101229.4, 101281, 101445.2, 101665.1, 101856.7, 
    102030.5, 102189.4, 102393.1, 102530.7, 102636.1, 102704.3, 102730.2, 
    102713.2,
  101354.2, 101375.9, 101240.3, 101257.5, 101447.9, 101682.6, 101924.9, 
    102192.2, 102401.7, 102553.1, 102653.9, 102757.9, 102799.5, 102814.1, 
    102771.4,
  101331.4, 101336.8, 101232.5, 101204.6, 101406.6, 101683.9, 101989.2, 
    102233.1, 102430.2, 102562.7, 102742.8, 102844.9, 102897, 102908.2, 
    102854.3,
  101343.5, 101402.8, 101476.3, 101523.1, 101580.6, 101570.3, 101561.9, 
    101583.4, 101615.9, 101339.3, 101465.4, 101748, 101645.1, 101289.6, 
    101157.4,
  101278.5, 101313.8, 101397, 101466.1, 101543.6, 101463.5, 101692.3, 
    101693.8, 101728.6, 101824.8, 101875.3, 101975.7, 101984.9, 100207.9, 
    100863.7,
  101169.4, 101200.2, 101277.5, 101398.2, 101395.7, 98308.05, 101671.3, 
    101939.8, 101968.5, 102004.6, 102066.8, 102144.8, 102201.1, 102220.5, 
    102180.8,
  100985.9, 101023, 101112.8, 101243, 101451.4, 101352.5, 98147.23, 101721.2, 
    102043.6, 102140.7, 102224.4, 102291.7, 102358.1, 102389.8, 102344.7,
  100784.5, 100823.8, 100921.7, 101104.2, 101350.6, 101618.3, 101562.3, 
    96090.59, 95535.07, 102019.1, 102357.1, 102430.7, 102504.4, 102503.7, 
    102515.8,
  100633.5, 100646.7, 100709.6, 100928.6, 101194.7, 101493.2, 101759.1, 
    101758.8, 101761.7, 102267.6, 102406.4, 102541.6, 102601.2, 102619, 
    102581.5,
  100666.8, 100608.4, 100593.3, 100797.8, 101124.2, 101448.3, 101685.3, 
    101984.6, 102192.4, 102335.7, 102489.7, 102625.4, 102668.4, 102671.5, 
    102619.8,
  100830.1, 100697.1, 100601.4, 100730.1, 101052.8, 101420.7, 101698.4, 
    101916.4, 102137.9, 102393.3, 102575.9, 102677.4, 102715.5, 102678.5, 
    102608.7,
  100974.8, 100858.5, 100759.5, 100849.5, 101135.4, 101460.6, 101742.4, 
    102039, 102291.3, 102504, 102641.4, 102733.5, 102738.9, 102688.3, 102604.1,
  101077.8, 100991.2, 100901, 100982.7, 101203.2, 101506.5, 101799.9, 
    102075.6, 102317.5, 102508.9, 102686.8, 102778, 102777.7, 102722.3, 
    102640.3,
  101478, 101580.9, 101633.9, 101641.1, 101612.7, 101610.3, 101631.1, 
    101692.7, 101743.6, 101428.7, 101565.5, 101884.5, 101777.3, 101411.5, 
    101247.8,
  101624, 101688.5, 101720.6, 101704.3, 101611.8, 101434.6, 101651.7, 
    101584.3, 101619.4, 101730.8, 101780.9, 101926.7, 102005, 100225, 100857.4,
  101724.1, 101762.4, 101757.6, 101745.5, 101555.7, 98216.69, 101392.5, 
    101688.4, 101604.2, 101649, 101746.4, 101909.9, 102030, 102098.9, 102095.3,
  101756.8, 101768.8, 101731.3, 101681.6, 101629.4, 101374.4, 97854.8, 
    101170.8, 101519.1, 101627.6, 101721.4, 101869.2, 102042.1, 102156.9, 
    102176,
  101758, 101723.4, 101648.6, 101577.6, 101505.3, 101479.9, 101273.3, 
    95669.16, 94961.65, 101308.2, 101718.5, 101842.1, 102044, 102146.6, 
    102248.6,
  101665.1, 101584.1, 101440.7, 101339.1, 101219.5, 101189.1, 101237.1, 
    101160, 101121.1, 101524.3, 101650.1, 101825.1, 102039.4, 102175.4, 
    102277.2,
  101505.9, 101374, 101190.9, 101031.4, 100902.3, 100861, 100911.6, 101119.2, 
    101272.1, 101379, 101583.2, 101821.3, 102031, 102187.4, 102277.5,
  101316.3, 101127.1, 100867.4, 100618.4, 100412, 100431.1, 100572.9, 
    100753.8, 100987.8, 101284.6, 101553.5, 101813.5, 102045, 102194.8, 
    102280.5,
  101141.8, 100890.5, 100573.1, 100224.5, 99962.23, 100025, 100282.2, 
    100634.2, 100953.9, 101253.6, 101559.3, 101853.6, 102065.2, 102200.3, 
    102277.7,
  100994, 100682.4, 100336.9, 99827.92, 99550.27, 99717, 100089, 100505.1, 
    100901.5, 101259.3, 101623.7, 101919.4, 102098, 102240.8, 102298.5,
  99950.98, 100070.1, 100199.4, 100342.3, 100519.3, 100681.1, 100812.8, 
    100922.8, 100985.9, 100717.7, 100840.4, 101150.5, 101091.2, 100824, 
    100747.9,
  100050.3, 100191, 100356.1, 100545.6, 100706.3, 100759.9, 101028.3, 
    101040.2, 101086.9, 101165.7, 101147, 101169.3, 101204.6, 99537.02, 
    100222.6,
  100389.4, 100507.3, 100636.9, 100778.5, 100728.8, 97604.99, 100966.4, 
    101233.4, 101127, 101134.3, 101145.4, 101161.7, 101190.6, 101263.5, 
    101335.1,
  100733.7, 100822.9, 100907.8, 100996.9, 101049.6, 100867.5, 97425.6, 
    100876.8, 101201.2, 101251.3, 101190.3, 101127.5, 101146.5, 101224.5, 
    101334.3,
  100959.1, 101019.1, 101054.5, 101095.5, 101119.5, 101171, 100992.7, 
    95317.49, 94544.19, 100912.9, 101202.6, 101096.9, 101096.1, 101128.2, 
    101298,
  101073.3, 101087.3, 101061.5, 101058.4, 101011, 101007.6, 101021.4, 
    100930.2, 100874.8, 101154.5, 101145.5, 101107.9, 101078.5, 101108.9, 
    101269.9,
  101074.2, 101059.1, 101000.3, 100943.2, 100863, 100784.4, 100722.1, 100776, 
    100819.8, 100865.2, 100990.5, 101053, 101056.3, 101128.9, 101277.1,
  101040.2, 100992.7, 100888.5, 100774.8, 100624.1, 100491.5, 100381.5, 
    100341.5, 100450.6, 100672.6, 100853.7, 100951.3, 101033.4, 101157.2, 
    101353,
  100998.4, 100911.8, 100770.1, 100629, 100421.5, 100200.6, 100043.5, 
    100051.8, 100189.5, 100409.7, 100669.4, 100859.6, 101006.3, 101209.5, 
    101407.6,
  100938.1, 100789.5, 100645.6, 100508.8, 100247.2, 100024.1, 99886.62, 
    99901.07, 100059.8, 100320.4, 100622.9, 100843, 101057.2, 101297.7, 
    101455.4,
  100641.7, 100469.6, 100307.9, 100128, 100001.4, 99899.73, 99819.97, 
    99800.4, 99833.71, 99581.11, 99682.06, 99976.55, 99872.99, 99568.47, 
    99537.22,
  100505, 100220.2, 99997.21, 99810.05, 99649.8, 99416.02, 99544, 99518.91, 
    99550.71, 99689.34, 99784.98, 99908.25, 99937.49, 98272.73, 98933.01,
  100524.6, 100197.6, 99908.45, 99675.14, 99384.16, 96182.72, 99241.2, 
    99485.16, 99449.77, 99581.41, 99724.73, 99873.55, 99954.83, 99971, 
    100054.4,
  100690.9, 100429.5, 100154.6, 99890.01, 99698.74, 99310.04, 95961.77, 
    99281.3, 99572.81, 99659.34, 99807.8, 99913.59, 100035.6, 100095.5, 
    100157.2,
  100778.1, 100601.8, 100406.8, 100201.5, 100028, 99890.27, 99502.3, 93935.4, 
    93402.2, 99663.23, 100007.6, 100060.9, 100175.2, 100172, 100290.6,
  100853.7, 100714.4, 100542.5, 100372.3, 100172.4, 100060.7, 99984.05, 
    99810.1, 99717.4, 100087, 100164.6, 100251, 100310.7, 100316.9, 100368.9,
  100879.5, 100780.2, 100657, 100505, 100365.1, 100213.4, 100100.9, 100151.1, 
    100171.9, 100180.9, 100269.6, 100375.9, 100398.3, 100399.6, 100434,
  100909.5, 100827.7, 100716.8, 100578.7, 100411, 100293.2, 100188.5, 
    100095.3, 100108.9, 100240.7, 100356.8, 100440.5, 100486.2, 100503.8, 
    100587.8,
  100915.9, 100865.9, 100788, 100677.2, 100538.2, 100384.4, 100261.3, 
    100230.3, 100225.3, 100260.7, 100385.8, 100515.9, 100580.4, 100658.6, 
    100780.1,
  100936.9, 100891.5, 100851.6, 100752.8, 100619.2, 100504.1, 100385.4, 
    100283, 100274.5, 100337.1, 100498.1, 100628.4, 100707.1, 100833.1, 
    100927.8,
  101039.3, 101161.2, 101298.1, 101403.7, 101462.8, 101450.4, 101393.5, 
    101316.3, 101167.3, 100650.2, 100489.2, 100534.1, 100189.1, 99579.97, 
    99258.83,
  101315.4, 101373.5, 101436.4, 101477.2, 101434, 101206, 101346.9, 101112.7, 
    100879, 100733.4, 100473.7, 100266.4, 100029.8, 98103.91, 98482.46,
  101474.4, 101507.7, 101516.4, 101529.5, 101332.6, 97951.36, 100976.9, 
    101158.3, 100849.6, 100589.5, 100273.2, 99994.98, 99706.49, 99521.41, 
    99397.93,
  101530.7, 101529.6, 101529.6, 101502.2, 101433.6, 101111.3, 97461.34, 
    100547.2, 100641.6, 100480.1, 100136.8, 99772.2, 99507.11, 99372.67, 
    99326.43,
  101534.2, 101520.8, 101513.9, 101460.5, 101402.8, 101268.4, 100948.3, 
    95079.91, 94224.22, 100255.7, 100137.1, 99727.17, 99455.81, 99303.81, 
    99353.57,
  101484, 101476.4, 101450.1, 101419.8, 101277, 101182.6, 101074.9, 100858.6, 
    100603.3, 100549.3, 100206, 99916.59, 99685.77, 99546.11, 99565.13,
  101427.5, 101428.3, 101426.3, 101358.5, 101256.1, 101120.2, 101015.5, 
    100989.8, 100818.7, 100553.7, 100329.8, 100169.1, 100012.7, 99940.36, 
    99944.05,
  101372.6, 101410.5, 101392.3, 101311.7, 101180.4, 101095.6, 101010.8, 
    100887.4, 100767.5, 100643.4, 100468.5, 100377.2, 100314.4, 100280.4, 
    100291.7,
  101380.1, 101434.6, 101384.3, 101305.8, 101211.8, 101112.7, 101026.8, 
    100984.6, 100876.8, 100724.7, 100621.9, 100570.4, 100544.6, 100539.4, 
    100550,
  101430.9, 101447, 101389.1, 101312.7, 101210.2, 101133.3, 101053.3, 
    100950.4, 100870.1, 100785.5, 100757.2, 100743.3, 100743.5, 100760.4, 
    100776.2,
  99768.73, 99802.19, 99884.43, 100012.5, 100192.3, 100400.1, 100683.6, 
    100971.3, 101239.6, 101132.4, 101368.4, 101706.9, 101548.1, 101027.5, 
    100710.9,
  99969.32, 99851.24, 99945.44, 100119.5, 100271.1, 100403.3, 100781.5, 
    101008.9, 101231.2, 101496, 101631.1, 101740.6, 101681.1, 99764.4, 
    100166.2,
  100420.5, 100211.5, 100193.1, 100341.8, 100312, 97413.94, 100824.4, 
    101245.1, 101377.5, 101555.8, 101663.5, 101720.4, 101655.8, 101516.3, 
    101260,
  100781.7, 100657.5, 100585.9, 100599.8, 100728.6, 100548, 97466.95, 
    101035.4, 101506, 101626.9, 101692.3, 101676.1, 101645.5, 101474.3, 
    101250.9,
  101062.2, 100989.3, 100945, 100930.3, 100996.2, 101137.2, 100950.6, 
    95520.34, 94966.63, 101391.3, 101691.2, 101658, 101624.3, 101431.5, 
    101299.6,
  101257.5, 101228.7, 101195.1, 101201.1, 101184.1, 101252, 101380, 101275.2, 
    101285.2, 101664.5, 101639.8, 101673.1, 101612, 101483.2, 101371.4,
  101397.9, 101406.2, 101400.3, 101391.5, 101415.7, 101425.8, 101461, 
    101624.4, 101672.1, 101613.7, 101644.5, 101663, 101603.3, 101521.8, 
    101449.9,
  101490.1, 101533.5, 101523, 101520.4, 101503.8, 101551.9, 101574.5, 
    101562.3, 101603.4, 101666.1, 101676.4, 101677.9, 101631.8, 101574.9, 
    101553,
  101583.3, 101619.1, 101609.2, 101612.2, 101612.7, 101629.9, 101660.5, 
    101724.5, 101730.2, 101700.5, 101694.9, 101710.8, 101658.6, 101619.4, 
    101602.7,
  101663.2, 101659.2, 101644.7, 101640.6, 101640.9, 101655.8, 101675.6, 
    101663.9, 101664.7, 101696.8, 101733.3, 101742.1, 101707.1, 101699.8, 
    101689.9,
  100729.6, 100635.7, 100559.2, 100518.2, 100510.6, 100465.3, 100536.8, 
    100724, 100899.6, 100745.8, 100990.8, 101438.4, 101522.8, 101350.6, 
    101298.1,
  100826.1, 100640.8, 100507.7, 100495.7, 100418.9, 100277.2, 100509.2, 
    100593.2, 100742.2, 100952, 101135, 101412.8, 101653.8, 100089, 100792.9,
  100926.7, 100701.4, 100489.5, 100438.1, 100289.1, 97168.02, 100321.4, 
    100665.3, 100739.7, 100888.3, 101089.7, 101378.8, 101655.6, 101831.6, 
    101955.9,
  101027.8, 100799.3, 100559.9, 100342.8, 100362.4, 100069.6, 96939.6, 
    100246.3, 100669.9, 100873.1, 101093.3, 101345.5, 101661.7, 101890.7, 
    101996,
  101148.8, 100934.5, 100691.7, 100450.5, 100293.9, 100353.5, 100130, 
    94962.39, 94430.73, 100593.4, 101136.8, 101350.2, 101670.7, 101866.5, 
    102052.9,
  101258.8, 101084.8, 100834.4, 100597, 100353.6, 100255.2, 100355.4, 
    100232.8, 100238.6, 100847, 101121.7, 101406, 101709.3, 101929.4, 102094.6,
  101363.1, 101222.4, 101023.9, 100786.9, 100563, 100398.3, 100339.8, 
    100547.8, 100756.4, 100904.5, 101175, 101492.4, 101763.2, 101982.8, 
    102127.9,
  101455.4, 101352.5, 101171.2, 100975.4, 100735.8, 100586.3, 100478.8, 
    100503.3, 100715.2, 101028.6, 101327.8, 101606.1, 101850.7, 102048.2, 
    102203.8,
  101523.9, 101468.8, 101348, 101198, 101008.4, 100856.5, 100784.4, 100884.8, 
    101054.8, 101258.6, 101504.8, 101744.2, 101941.4, 102114.4, 102245.4,
  101571.2, 101526.5, 101470.3, 101362.2, 101250.2, 101152.8, 101094.2, 
    101122.2, 101250.8, 101442, 101691.7, 101885.4, 102035.6, 102184.6, 
    102300.4,
  101191.1, 101077.6, 100924.2, 100802.1, 100704.6, 100625.3, 100678.9, 
    100829.9, 100966.6, 100757.4, 100920.7, 101257.3, 101216, 100982.1, 
    100976.9,
  101409.5, 101272.1, 101116.7, 100988.9, 100777, 100613.8, 100754.8, 
    100748.4, 100853.5, 100992.1, 101065.3, 101204.4, 101301.5, 99733.41, 
    100456.8,
  101563.3, 101464.9, 101308.9, 101203.2, 100881.5, 97565.78, 100716.9, 
    100885.7, 100870.7, 100936, 101002.6, 101121, 101252.6, 101359.7, 101505.4,
  101694.8, 101576.6, 101470.2, 101309, 101231.3, 100842.1, 97346.47, 
    100565.6, 100848.4, 100936.9, 100993.6, 101052.1, 101185.8, 101344, 
    101515.3,
  101764.1, 101689.9, 101570.6, 101445.8, 101294, 101251.9, 100921.9, 
    95262.53, 94615.13, 100676.2, 100972.9, 100990.9, 101106.5, 101241.7, 
    101477.2,
  101767.1, 101715.4, 101606.7, 101485.3, 101315.3, 101199.1, 101137.9, 
    100957.1, 100745.1, 101018.9, 100966.7, 100972.6, 101051.8, 101194.7, 
    101437.2,
  101722.7, 101698.7, 101632.8, 101493.7, 101336.3, 101178.5, 101034.4, 
    101026.2, 101016.8, 100920.4, 100913.2, 100943.9, 101002.8, 101151.8, 
    101396.1,
  101636.1, 101636, 101581.3, 101453.6, 101263.9, 101107.1, 100932.5, 
    100747.8, 100671.9, 100721.7, 100785.3, 100852.6, 100962.6, 101140.5, 
    101409.3,
  101530.3, 101578.1, 101561.5, 101436.8, 101261.5, 101060.3, 100834.3, 
    100682.3, 100599.7, 100561.8, 100613.1, 100734.8, 100910.8, 101150.8, 
    101443.2,
  101441.6, 101502.5, 101500.1, 101393.3, 101230.2, 101043.5, 100808, 
    100540.8, 100389.3, 100357.9, 100476.9, 100647.8, 100881.5, 101171.1, 
    101473.3,
  100062.1, 99795.45, 99658.91, 99739.14, 99866.6, 100061.9, 100279.7, 
    100523.7, 100737.3, 100635.9, 100880.6, 101278.4, 101264.4, 101024.6, 
    100979.6,
  100536.3, 100249.6, 100004.9, 99950.02, 99977.09, 100036.9, 100360.9, 
    100539.5, 100720.6, 100926.5, 101089.5, 101284.3, 101400.1, 99822.05, 
    100489.4,
  100974.2, 100699.2, 100468.7, 100299.4, 100075.6, 97139.49, 100399.6, 
    100736.8, 100867.6, 100995.1, 101130.7, 101281, 101417.7, 101485.9, 
    101538.1,
  101338.2, 101114.9, 100905.5, 100708.9, 100597.9, 100277.2, 97188.24, 
    100617.5, 101001.8, 101161.6, 101251.9, 101321.8, 101415.3, 101510.8, 
    101554.9,
  101585.1, 101454.6, 101296.3, 101111.9, 100968, 100932.6, 100604.9, 
    95318.4, 94891.87, 101111.6, 101393.8, 101389.2, 101443.3, 101458.6, 
    101547.2,
  101717.9, 101666, 101563.7, 101468, 101302.8, 101230.7, 101223.3, 101058.4, 
    101038, 101452.7, 101486.1, 101496, 101491, 101483.1, 101508.5,
  101771.3, 101750.4, 101736.4, 101691.5, 101622.4, 101545.9, 101496.6, 
    101604.2, 101640.7, 101564.6, 101567.5, 101591.9, 101565.9, 101541.9, 
    101489,
  101752, 101747.5, 101747.1, 101802.4, 101758.8, 101743, 101699.3, 101605.8, 
    101584.2, 101650.3, 101658.6, 101639.4, 101614.2, 101587.7, 101547.7,
  101662.9, 101690.9, 101726.1, 101803.9, 101840.9, 101830.5, 101820.2, 
    101851.4, 101821.9, 101741.9, 101684.9, 101660.2, 101629.8, 101593.1, 
    101539,
  101556.7, 101568.4, 101618.6, 101711.1, 101791.7, 101836, 101813.4, 
    101745.4, 101687, 101649.6, 101653.8, 101618, 101563.1, 101525.9, 101489.9,
  99569.21, 99431.12, 99570.66, 99815.08, 99968.28, 100002.9, 100107.6, 
    100288.7, 100516.3, 100463.4, 100785.3, 101251.7, 101326.2, 101151.8, 
    101143.4,
  99768.34, 99454.27, 99545.59, 99771.43, 99862.57, 99822.52, 100075.4, 
    100253, 100463.2, 100733.4, 100991.9, 101273, 101479.6, 99976.55, 100695.2,
  100073.6, 99699.89, 99633.35, 99786.44, 99731.19, 96725.53, 99982.36, 
    100355.4, 100566.2, 100742.9, 100992.3, 101251.1, 101493, 101638.8, 
    101751.4,
  100415.7, 100001.9, 99794.61, 99783.47, 99871.14, 99632.79, 96637.77, 
    100042.3, 100527.3, 100754.5, 100997.2, 101214.6, 101472.4, 101658.4, 
    101781.6,
  100739, 100375.3, 100076.2, 99933.37, 99878.87, 100005.7, 99831.9, 
    94830.52, 94461.4, 100537.2, 101011.8, 101188.1, 101436.7, 101604.6, 
    101778.4,
  100995.7, 100734, 100415.3, 100185.6, 99980.74, 99963.45, 100152.2, 
    100102.1, 100173.6, 100729.6, 100941.1, 101169.6, 101401.8, 101596, 
    101762.6,
  101204.5, 101023.8, 100776.1, 100526.9, 100297.6, 100142.3, 100184.7, 
    100434.5, 100637.4, 100740.2, 100935.3, 101170.4, 101390.8, 101590.1, 
    101749.4,
  101370.8, 101237.4, 101061.4, 100864.7, 100637.6, 100427.7, 100350.7, 
    100368.9, 100515.3, 100757.2, 100982.2, 101201.5, 101413.4, 101614.3, 
    101780.6,
  101490.4, 101399.8, 101281.6, 101167.8, 101002.8, 100822.9, 100679.8, 
    100716.5, 100809.7, 100928.1, 101094.3, 101301.1, 101493.5, 101680.6, 
    101835.2,
  101564.4, 101468.4, 101408.3, 101325.1, 101251, 101149.3, 101019.9, 
    100916.2, 100936.6, 101043.1, 101239.5, 101413.6, 101581.9, 101758.1, 
    101895.6,
  100882.2, 100569.7, 100520, 100668, 100861.4, 100937.5, 101021, 101001.1, 
    100838.6, 100517.3, 100795.1, 101235.8, 101291.8, 101052.3, 101008.3,
  100833.6, 100464.9, 100377.3, 100546.2, 100711.6, 100719.1, 100959.4, 
    100926.3, 100786.6, 100844.2, 101070.1, 101350, 101538.4, 99989.77, 
    100720.9,
  100875.8, 100472.3, 100327.9, 100490.1, 100538.8, 97448.47, 100762.8, 
    100979.7, 100924.8, 100904.2, 101143.8, 101403.6, 101663.7, 101801.4, 
    101906.1,
  100965.8, 100580, 100387.3, 100417.1, 100648.6, 100436.1, 97247.5, 
    100543.8, 100781.6, 100932.3, 101192.8, 101436.6, 101721.5, 101912.7, 
    102035.3,
  101092, 100755.5, 100516, 100454.6, 100540.7, 100752.7, 100516.8, 95188.45, 
    94675.66, 100751.8, 101226.1, 101455.3, 101743.9, 101922.5, 102098.7,
  101213, 100940.6, 100639.9, 100493.4, 100449.6, 100519.8, 100740, 100620.1, 
    100528.5, 100978.8, 101180.5, 101449.8, 101717.2, 101929, 102100,
  101328.1, 101106.2, 100831.2, 100599.7, 100446.7, 100455.8, 100535.9, 
    100807.4, 100967.9, 100987.1, 101139.6, 101397.9, 101652.9, 101871, 
    102041.6,
  101425.9, 101240.1, 100990, 100740.6, 100486.3, 100351.8, 100433.1, 
    100525.9, 100679.3, 100910.9, 101096.2, 101312, 101556.5, 101780.3, 
    101971.7,
  101488.2, 101364.3, 101161.8, 100934.9, 100674.2, 100409.1, 100318.6, 
    100510.6, 100711.3, 100869, 101033.1, 101232.8, 101449.8, 101664.8, 101855,
  101507.3, 101430.5, 101273.6, 101081.4, 100847.3, 100589.6, 100321.6, 
    100323.4, 100485.9, 100691.4, 100934.2, 101132.4, 101332.2, 101540.4, 
    101729.5,
  101951.6, 101806.6, 101631.8, 101548.9, 101550.3, 101558.9, 101534.5, 
    101546.6, 101440.5, 100939.4, 100821, 101087.8, 100967.6, 100613.5, 
    100442.3,
  101855.8, 101643.6, 101431.3, 101354.6, 101310.6, 101220.4, 101417.6, 
    101400.1, 101271.8, 101218.9, 101134.5, 101227.4, 101236.3, 99568.5, 
    100197.7,
  101746.5, 101497.2, 101267.5, 101185.4, 101081.3, 97862.98, 101134.6, 
    101380.7, 101309.5, 101214.9, 101210.2, 101314.7, 101416.2, 101459.7, 
    101432.6,
  101659.9, 101404.8, 101186.5, 101046.8, 101118.6, 100872, 97546.36, 
    100852.4, 101068.5, 101130.5, 101271.4, 101399, 101535.3, 101606.1, 101627,
  101596.9, 101385.9, 101128.9, 101029.9, 101021.2, 101159.2, 100897.9, 
    95333.2, 94736.14, 100896.3, 101336.6, 101473.7, 101634.4, 101675.6, 
    101783.5,
  101568.1, 101399.4, 101117, 100995.6, 100974.7, 101004.2, 101138.5, 
    100920.6, 100710, 101129.8, 101329.1, 101535.2, 101699.8, 101794.9, 
    101893.6,
  101566.3, 101447.4, 101176.7, 100994.4, 101002, 101020.5, 101030.4, 101082, 
    101071.4, 101116.9, 101342, 101570.9, 101751.4, 101877.8, 101992,
  101603.6, 101502.1, 101254.7, 101032.6, 100941.4, 100978.1, 101031, 
    100915.1, 100895.6, 101097.6, 101358.6, 101580.6, 101788.8, 101940.1, 
    102085.4,
  101644.5, 101587.5, 101402.7, 101180.4, 101014.3, 100964.6, 100984.5, 
    101013.4, 101030.6, 101156, 101367.4, 101592.5, 101799.4, 101961.7, 
    102105.1,
  101684.9, 101649.3, 101528.3, 101351.4, 101121.4, 100996.2, 100961.9, 
    100915.4, 100954.7, 101110.5, 101367.7, 101586.3, 101783.6, 101954.3, 
    102098.1,
  102276.5, 102341.9, 102326.4, 102289.6, 102240.3, 102118, 102027.3, 
    101942.6, 101814, 101286, 101149.3, 101156.9, 100907.2, 100569, 100484.4,
  102230, 102270.5, 102270.2, 102241, 102142.1, 101893.7, 102023.5, 101841.6, 
    101686.2, 101606.6, 101419.9, 101258.2, 101160.2, 99492.55, 100184.6,
  102174.7, 102192.4, 102179.3, 102160.7, 102011.8, 98591.86, 101760.1, 
    101944.3, 101768.3, 101598, 101431, 101303.1, 101292.7, 101365.4, 101411.1,
  102123, 102094.3, 102079.9, 102035.4, 102014.8, 101759.8, 98166.34, 
    101430.8, 101621, 101583.1, 101449.7, 101354.6, 101384.3, 101507.4, 
    101615.1,
  102032.2, 102001, 101965.7, 101937.6, 101888.8, 101891.5, 101646.5, 
    95933.95, 95124.55, 101376.7, 101497, 101413.1, 101458.9, 101576.1, 
    101765.7,
  101934.6, 101900, 101833.6, 101768.9, 101675.8, 101643.8, 101696.5, 
    101575.8, 101457.2, 101664.4, 101536.8, 101483, 101503.5, 101671.5, 
    101843.1,
  101850.1, 101788.8, 101682.1, 101573.7, 101482.7, 101454.2, 101452.5, 
    101601.9, 101666.8, 101574.3, 101556.1, 101498.7, 101526.8, 101713.1, 
    101896.5,
  101761.2, 101638.2, 101494.6, 101362.4, 101216.7, 101204.8, 101248.5, 
    101299.6, 101387.6, 101489.4, 101516.7, 101480.4, 101546.5, 101745.4, 
    101956.7,
  101652.4, 101509.2, 101366.5, 101227.7, 101058.7, 100998.9, 101050.5, 
    101200.4, 101337.7, 101390.2, 101436.9, 101463.7, 101544.5, 101757.2, 
    101971.1,
  101575.8, 101387, 101270.4, 101117.2, 100867, 100746.2, 100822.2, 100936.4, 
    101091.2, 101205.9, 101354.8, 101424.2, 101534.2, 101765.3, 101974.5,
  102345.6, 102452.4, 102473.4, 102481.4, 102450.4, 102387.9, 102300.5, 
    102163.2, 101958.1, 101424.7, 101280.8, 101348.3, 101092.4, 100646.4, 
    100436.6,
  102371.5, 102480.1, 102535.6, 102547.8, 102487.5, 102310.9, 102429.8, 
    102243.2, 102080, 101921.5, 101667.2, 101556.1, 101433.2, 99667.96, 
    100244.8,
  102333.3, 102455.9, 102536.4, 102578.7, 102453.3, 99071.81, 102358.7, 
    102513.8, 102306.1, 102117.2, 101877.2, 101713, 101654.1, 101601.8, 
    101514.1,
  102285.6, 102389.6, 102475.4, 102529.9, 102542.1, 102384.6, 98741.38, 
    102168.3, 102321, 102306.6, 102089.9, 101918.7, 101797.8, 101790.2, 
    101736.5,
  102335.6, 102352.5, 102394.4, 102450.1, 102489.6, 102551, 102402.2, 
    96570.4, 95820.41, 102180.1, 102296.8, 102092.6, 101945.6, 101892.9, 
    101913.2,
  102317.1, 102311.2, 102293.2, 102313.4, 102330.8, 102383.1, 102457.4, 
    102403.5, 102287.5, 102469.9, 102384.9, 102246.6, 102060.5, 102025, 
    102031.7,
  102202.7, 102177.9, 102152.4, 102151.5, 102169.7, 102208.7, 102256.3, 
    102397.4, 102445.8, 102429.1, 102415.4, 102337.9, 102162.6, 102100.7, 
    102125.9,
  102090.7, 102035.8, 101966.6, 101936.2, 101917.9, 101960.9, 102029.6, 
    102087.2, 102181.8, 102314, 102359.4, 102330.2, 102247.2, 102165.7, 
    102213.4,
  102015.3, 101918.2, 101810.7, 101715.3, 101678.4, 101694, 101773.6, 
    101914.8, 102054.9, 102146.3, 102239.1, 102285.7, 102262, 102206.7, 
    102248.2,
  101952.7, 101777.5, 101598.8, 101466, 101411.2, 101422.5, 101500.3, 
    101594.5, 101741, 101885.7, 102079.5, 102180.3, 102221.4, 102226.6, 102266 ;

 scalar_axis = 0 ;

 sftlf =
  0.5159525, 0.045606, 0.3841295, 0, 0.09859309, 0.3330989, 0.003261217, 0, 
    0.03607289, 0.7158654, 0.6944581, 0.4642971, 0.7396766, 0.6573148, 1,
  0.001847372, 0, 0, 0, 0.5296907, 0.5066301, 0, 0, 0, 0.1899712, 0.5492381, 
    0.118482, 0.0927158, 0.843343, 1,
  0, 0, 0, 0, 0.3371468, 0.8556198, 0.1306061, 0, 0, 0, 0.02473423, 
    6.294356e-05, 0.005740512, 0.06632636, 0.5030367,
  0, 0, 0, 0, 0, 0.2586107, 0.8765578, 0.2410029, 0, 0, 0, 0, 0, 0.04698182, 
    0.2655103,
  0, 0, 0, 0, 0, 0, 0.144052, 0.8812297, 0.6102951, 0.3213011, 0.03357667, 0, 
    0, 0.005859504, 0,
  0, 0, 0, 0, 0, 0, 0, 0.03178087, 0.2700712, 0.3195445, 0.3046227, 0, 0, 0, 
    0.0009363425,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01283686, 0, 0, 0, 0, 0.04670987,
  0, 0, 0, 0, 0, 0, 0, 0.01840907, 0.1205428, 0.4131123, 0.2665586, 0, 
    0.02034558, 0.008879703, 0.0442122 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.141347, 0.07456003, 0.2762221, 0, 0.2154952, 0.5089986, 0.007178012, 0, 
    0.1467785, 25.31165, 20.60715, 2.120196, 15.979, 48.81725, 63.64272,
  0.001503375, 0, 0, 0, 0.8848332, 11.68672, 0, 0, 0, 0.4694104, 0.9680001, 
    0.09868675, 1.334438, 150.908, 101.0153,
  0, 0, 0, 0, 8.803595, 280.9762, 7.478715, 0, 0, 0, 0.0046135, 0, 
    0.00845787, 0.9458157, 6.678408,
  0, 0, 0, 0, 0, 12.95772, 307.1121, 15.76765, 0, 0, 0, 0, 0.001950179, 
    0.08926713, 2.882818,
  0, 0, 0, 0, 0, 0, 9.245329, 485.3841, 540.1508, 15.00115, 0.01623012, 0, 0, 
    0.06344586, 0.01027276,
  0, 0, 0, 0, 0, 0, 0, 1.278773, 12.13823, 0.8518202, 0.2699268, 0, 0, 
    0.01012854, 0.01599434,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05785002, 0, 0, 0, 0, 0.2725836,
  0, 0, 0, 0, 0, 0, 0, 0.3482242, 1.154397, 3.605569, 0.8750445, 0, 0.158783, 
    0.02233585, 0.6264485 ;
}
