netcdf atmos.1980-1981.aliq.06 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:19 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.06.nc reduced/atmos.1980-1981.aliq.06.nc\n",
			"Mon Aug 25 14:40:42 2025: cdo -O -s -select,month=6 merged_output.nc monthly_nc_files/all_years.6.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.171193e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002102946, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.406456e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0005630884, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.536484e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002303574, 0, 0, 0.0003734573, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008678528, 0.0003892796, 0.0008556678, 0, 
    0, 0, 0, 0, 0, 0, -5.195371e-06, -2.199852e-05, 1.33398e-06, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.000742732, 0, 8.977097e-05, -2.783366e-06, 
    -6.425088e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.622653e-05, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, -3.746482e-06, 2.721147e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.227532e-05, -1.034185e-05, 
    2.553835e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 3.430411e-06, 0, 0.0009568257, 0, 0, 0.00288872, 
    2.879459e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -2.002385e-06, 0, 0, 0, 0, 0, 0, 0, 0, -8.092668e-06, 0.006371549, 
    0.00074921, 0.004358876, -3.246882e-06, 0, 0, 0, 0, 2.894262e-05, 
    -7.950248e-06, -2.726876e-05, 3.582692e-05, 1.79661e-05, 0, 0, 
    -7.033881e-07, 0.0006919198, 6.72864e-05, 0,
  0, 0, 0, 0, 0, 0, -1.230499e-05, 0.001525508, 0, 0.0005339765, 
    0.0003088727, 0.0002238412, -5.165744e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0005302972, -5.1049e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -2.247889e-05, 0.0002485114, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.508483e-05, 0, -1.068438e-06, -5.569397e-05, -8.163322e-06, 
    0, -2.57509e-05, 0, 0.0003300051, 0.0008055291, -4.357067e-05, 
    0.0004674318, 1.565624e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 4.817576e-05, 0, 0, 0, -8.684445e-06, 0, 1.007286e-05, 1.096211e-06, 
    0.001984987, 0, -2.442739e-11, 0.005263955, -3.559056e-06, 1.296357e-05, 
    -9.314459e-07, 0, -3.532664e-05, 0, 0, 0, 0, 0, 1.186832e-05, 
    0.0003370769, 0, 0, 0, 0,
  -2.551894e-06, 0, 0, 0, 0, 0, 0, 0, 0, -4.781859e-05, 0.009888076, 
    0.00122029, 0.01089039, 0.001628543, -2.903688e-06, 0.00109497, 
    -1.259217e-05, 0, 0.0004196631, -4.09419e-05, 0.0001213032, 0.0004492466, 
    0.001509752, 9.167794e-06, 0.000426853, -2.873622e-05, 0.001315498, 
    0.000308495, 0.0004375288,
  0, 0, 0, 0, 0, 0, 0.001127918, 0.003926818, 0, 0.001028856, 0.001684226, 
    0.001441947, -5.252958e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006704045, 
    9.618536e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -6.118441e-05, 0.00041589, 0.0001284354, 
    -8.447724e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.567809e-08, 0, 4.114292e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.541885e-07, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000220416, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.001504789, 0, 0.0008691188, 0.0002500225, -5.943493e-05, 0, 
    2.675046e-05, -3.669267e-06, 0.003082738, 0.002368959, -5.906778e-05, 
    0.002440971, 0.0001231739, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 7.93279e-05, -3.777035e-06, 0, 0, 5.688198e-05, 0, 3.074501e-05, 
    0.0002561661, 0.002264448, 0, 0.000647849, 0.01005241, -4.086201e-06, 
    0.0009094456, -4.935152e-06, 6.570405e-06, -1.709484e-05, 0, 0, 0, 0, 0, 
    0.001526416, 0.001492395, 0, 0, 0, 0,
  -1.28985e-05, 0, 0, 0, 0, 0, 0, 0, 0, -4.552579e-05, 0.01395857, 
    0.002535556, 0.02105077, 0.003570749, -2.342717e-05, 0.002060616, 
    -7.251409e-05, -2.99125e-05, 0.0006705938, -5.625244e-05, 0.0004995379, 
    0.003123851, 0.005914791, 3.667118e-05, 0.001635083, 0.0009186276, 
    0.002723379, 0.001924624, 0.001061971,
  0, 0, 0, 0, 0, -4.523368e-06, 0.005296267, 0.0078215, 0, 0.003206443, 
    0.00293403, 0.00766473, 0.002524501, 0, 0, 0, 0, 0, 0, 0, 0, 0.001440515, 
    0.001080876, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0001062716, 0.003256653, 0.000952834, 0.0004409293, 
    -3.537503e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.102299e-05, -3.530639e-08, 0.0007619441, 
    0, 0, 0, 0, 0, 0, 0, 0, -1.857715e-05, 1.941943e-05, -1.186215e-05, 
    8.847512e-06, -2.52019e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.429309e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.909807e-05, -6.517223e-06, 0, 
    0, 0, 4.258817e-05, -2.382211e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.869625e-06, 0.001107982, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.002400339, 9.08835e-06, 0.002083541, 0.0007937691, 
    -2.363134e-05, 0, 0.000612536, -5.719167e-06, 0.005710593, 0.004562792, 
    0.0001102939, 0.003666335, 0.0009577465, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0001160145, -1.157047e-05, 0, 0, 0.0002219554, 0, -4.316318e-05, 
    0.0005952763, 0.002562009, 2.483836e-06, 0.001458697, 0.02190699, 
    0.0002336282, 0.001194948, -1.451903e-05, 0.0002684599, 2.899665e-05, 0, 
    0, 0, 0, -3.384745e-09, 0.003053786, 0.003310948, 0, -5.950134e-06, 0, 0,
  -1.786929e-05, 0, 0, 0, 0, 0, 0, -7.713586e-06, -9.206666e-06, 
    0.0009544626, 0.02026557, 0.008048557, 0.03362794, 0.007549801, 
    0.001544768, 0.003015632, -0.0002016458, -8.089953e-05, 0.001094485, 
    -9.120073e-05, 0.004835841, 0.01125636, 0.01075038, 0.0001132624, 
    0.002800456, 0.001121075, 0.004407872, 0.007546599, 0.00245106,
  0, 0, 0, 0, 0, -4.2847e-05, 0.009109744, 0.01207492, -1.067153e-05, 
    0.00837573, 0.007394536, 0.01955789, 0.007294177, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002975009, 0.003569657, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -0.0002399381, 0.008740885, 0.002247422, 0.004076225, 
    0.002550481, -2.803348e-06, 0, 0, 0, -5.622454e-06, 0, 0, 0, 0, 0, 0, 0, 
    -8.25106e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -6.851652e-06, 0.0008548247, 0.001515965, 
    0.001915282, 0.0006475989, 0.0001186654, 0, 0, 0, 0, 0, 0, 0.0001871467, 
    0.002250536, -6.724121e-05, 0.0009424026, -1.771933e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001339757, 0, 0, 0, 0, 0, 0, 0, 
    0.0007183905, 0.0008671766, 4.585681e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -2.697295e-07, 2.276662e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -8.561324e-06, 0.001264289, 0, 0, 0, 0, 0.0003998092, 0, 
    -1.048478e-05, 0.001658016,
  0, 0, 0, 2.694347e-05, -1.069066e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002805016, 0.0001939005, 0.0003660694, -4.781928e-05, -3.071555e-05, 
    0.001342421, -2.979576e-05, 0, 0, 0, 0, 0.0004043798, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.150706e-05, 0.003012583, 0, 0, 0, 
    0, -2.063313e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.003450436, 0.0001928229, 0.003723523, 0.002109757, 
    0.0005750505, 0, 0.001536925, 0.002089864, 0.01228145, 0.009689319, 
    8.783529e-05, 0.008746195, 0.002700984, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 9.479901e-05, -7.380415e-05, 0, 0, 0.0009566686, -1.258377e-05, 
    0.001904946, 0.001319497, 0.002539934, 0.0001716519, 0.003159055, 
    0.04017132, 0.000448488, 0.003894842, -3.051784e-05, 0.0003126002, 
    0.001062174, 0, 0, 0, 0, -1.5216e-05, 0.004795987, 0.005230624, 0, 
    -2.211221e-05, -8.073053e-06, 0,
  0.0001784983, 0, -1.026377e-06, 0, 0, -9.999791e-06, 4.589777e-05, 
    0.0001587559, 0.0001378398, 0.003645491, 0.0238621, 0.01856651, 
    0.04912184, 0.01416398, 0.002430547, 0.007771592, 0.0003007424, 
    -0.0002449178, 0.001956668, 0.0001847343, 0.009945451, 0.02318206, 
    0.01587473, 0.002000356, 0.005277283, 0.001798961, 0.008851251, 
    0.01896522, 0.002845486,
  0, 0, 0, 0, 0, 2.532904e-05, 0.01267984, 0.01605238, 0.0006499996, 
    0.02184418, 0.01367051, 0.03133325, 0.0152001, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.005138481, 0.00971485, -8.00581e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.912826e-05, -0.0003003807, 0.01582352, 0.003873987, 
    0.01330825, 0.01103155, 7.41782e-06, 0, -2.686893e-06, 0.001089482, 
    -1.967099e-05, 0, 0, 0, 0, -1.555785e-05, 3.243746e-07, 0, 0.0005876576, 
    0, 0, 0, 0,
  0, 3.963477e-06, -6.125656e-07, 0, 0, 0, 0, 0, 0.0002712384, 0.0006928657, 
    0.005734147, 0.006048746, 0.005018118, 0.00395474, 0.003673024, 
    -1.992706e-05, 0, -1.714769e-06, 0, 0, 0, 0.001925346, 0.006019815, 
    -7.764385e-05, 0.002656304, 0.007014059, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001926403, -9.590203e-05, 0.000703902, 
    0.001224965, 0, -1.81734e-05, -9.620874e-07, 0, 0, 0, 0.0002043012, 
    0.002401869, 0.002304468, 0.001445199, 0.0009446337, 0.00113576, 
    -4.491578e-07, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.814485e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005221962, 
    0, 0, -1.043502e-05, 0, 0, -7.303741e-06, 0.0008036988, 0,
  0, 0, 0, 0.0003694767, 0.003392402, -3.067094e-06, -4.297588e-06, 0, 0, 0, 
    -1.570406e-05, 0, 0, 0, 0, 0.0002564281, 0, 0, 0.0002671218, 
    8.655028e-05, 0.00673949, 0.0006475483, 0, 0.0001483789, 0, 0.002542383, 
    0.002420344, 0.0008975122, 0.002529085,
  0, 0, 0, 0.0003135863, -7.700036e-07, 0, 0, 0, 0, 0, 5.748809e-06, 
    -1.026772e-06, 0, 0, 0.005251176, 0.006773027, 0.003197072, 0.00111173, 
    0.001613614, 0.003710283, 0.002135964, -5.068294e-07, 0, 0, 0, 
    0.001733668, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002296147, 0.006621686, 
    0.0002460501, -9.680804e-06, -7.481379e-06, 4.0035e-05, -9.778091e-07, 0, 
    0, 0.000464453, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.009112999, 0.00461571, 0.00909544, 0.004966216, 0.00429878, 
    -9.747264e-05, 0.005744685, 0.004518969, 0.02610767, 0.01819832, 
    0.0005411529, 0.01641724, 0.006908323, 0.0001416062, 0, 0, 0, 
    -1.330684e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 6.864336e-05, -0.0001662979, 0, 0, 0.00181625, -3.430671e-05, 
    0.006753427, 0.002423449, 0.002816647, 0.0006501816, 0.006719923, 
    0.06823082, 0.008367917, 0.01248155, -6.454311e-05, 0.001200264, 
    0.004046759, 0, 0, 2.290462e-05, 0, -3.584065e-05, 0.008475663, 
    0.008312561, -5.024966e-05, 3.176499e-05, 3.136825e-06, -2.71486e-05,
  0.002600215, 6.514273e-05, 0.0002076556, 0, -1.206854e-06, 0.0003319134, 
    0.001659689, 0.001407038, 0.001216056, 0.01248994, 0.02806821, 
    0.04735884, 0.06917706, 0.02697301, 0.005650532, 0.01331957, 0.006773489, 
    0.001568881, 0.006267276, 0.001074396, 0.01850775, 0.04186111, 
    0.02317737, 0.007297812, 0.009212329, 0.004991434, 0.01260806, 
    0.05117419, 0.004121501,
  0, 0, 0, 7.248931e-06, -3.228316e-09, 6.506803e-05, 0.01933227, 0.02932558, 
    0.002872705, 0.0376834, 0.0323555, 0.05240482, 0.03419129, 1.985106e-07, 
    0.0002195388, -1.603282e-05, 0, 4.0693e-05, 9.957701e-05, -4.019375e-09, 
    -2.99064e-07, 0.008579977, 0.02289464, 0.001430299, 0, -9.206754e-05, 
    -1.951564e-05, 0, 0,
  0, -1.187192e-05, 0, 0, 0, 0, 0.0005006811, 0.00040292, 0.02624629, 
    0.010593, 0.03159853, 0.02933933, 0.0004398026, 0, -6.153688e-06, 
    0.002010046, 0.0003790388, 0, -1.548185e-06, 0, 0, 0.0005414615, 
    0.000198675, 2.739576e-05, 0.0008946251, 0, 0, 0, 0,
  -4.004611e-06, 0.000799407, 0.0007468596, 0, 0, 0, -1.758884e-06, 
    -1.820243e-09, 0.001801113, 0.004537364, 0.01250708, 0.01340413, 
    0.02123138, 0.01312421, 0.006800865, 0.002154049, 0, -1.985446e-05, 
    -2.750726e-09, 0, 0, 0.003669226, 0.01232134, 0.004213824, 0.008229953, 
    0.01027688, -6.575781e-08, -2.041203e-05, 0,
  0, 0, 0, 0, 0, -1.16849e-06, 0, -3.336702e-05, 0, 0.002094829, 0.002441353, 
    0.00424742, 0.004222119, 0.00363101, 0.0001009137, 0.002000834, 
    -3.075779e-06, 0, 0, 0, 0.003410422, 0.005463097, 0.007148621, 
    0.003104955, 0.004242441, 0.002329906, 0.000219561, 0.00102312, 0,
  0, 0, 0, -1.650057e-06, 0, 0, 0, 0, 0.0001438408, 0, 0, 0, 0.0003520765, 0, 
    0, 0, 0, 0, 0, 0, -5.774547e-05, 6.382781e-05, 0, -2.050712e-06, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002327711, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -6.308172e-06, 0, 0, 0.0004942449, 0.001653363, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003732354, 0, -1.436528e-05, 0, 0.0001146335, -1.103655e-05, 
    0.001245623, 0, 3.086729e-05, 0.0001773837, 0, 0, 0.001471539, 
    0.001810835, -4.31085e-06,
  -4.155764e-08, 0, -1.167144e-06, 0.001236471, 0.006267666, 5.032549e-05, 
    0.0005977851, -2.153796e-06, 0, 0, 0.001261115, 0, -1.473223e-06, 
    -6.42754e-07, -9.775784e-06, 0.002857185, 0.0006699657, 0.0002821773, 
    0.00276526, 0.002452064, 0.01464955, 0.006760249, -3.077763e-05, 
    0.003576166, -1.42272e-05, 0.00560829, 0.006885601, 0.003236416, 
    0.003668553,
  0, 0, 0.0001667843, 0.001583568, -1.264736e-05, -1.554746e-05, 0, 0, 0, 
    0.0001299554, 0.0005278281, 0.0003144706, 0, 0.0001361662, 0.009241381, 
    0.02013439, 0.01132351, 0.01005103, 0.01567667, 0.008725167, 0.006377217, 
    -6.627071e-05, 0, 0, 0, 0.004048995, -3.036944e-05, 0, 0,
  0, 0, 0, 0, 6.881604e-09, 0, 0, 0, -6.838254e-06, -1.255749e-05, 0, 0, 0, 
    0.001746253, 0.01075819, 0.005462386, 0.00461557, -3.127724e-05, 
    0.0003413364, 0.001183033, 0, 0, 0.0002352907, 4.164584e-05, 0, 0, 0, 
    -6.729059e-10, 0,
  0, 8.356008e-09, 0, 0, 0.013808, 0.01177178, 0.01352212, 0.01190795, 
    0.01611152, 6.568721e-05, 0.01352581, 0.009272758, 0.05103309, 0.0310056, 
    0.009436266, 0.03454382, 0.01928916, 0.0003703315, 3.466486e-06, 
    -2.89844e-08, 5.485232e-10, 7.45986e-08, -7.832534e-07, -6.450837e-06, 
    -3.867641e-11, -2.667892e-05, -1.027475e-11, -3.148687e-10, 1.415158e-06,
  -3.094762e-06, 0.003095708, 0.0003094412, -6.952458e-06, 0, 0.006454619, 
    0.0006846657, 0.01226834, 0.01032156, 0.01040754, 0.007006478, 
    0.02113828, 0.1119915, 0.03086797, 0.02891621, 0.0003558696, 0.004615984, 
    0.00598876, -5.178996e-07, -1.989839e-06, 0.001114279, 1.888529e-05, 
    0.001425778, 0.03387206, 0.01822618, 0.000138099, 9.063203e-05, 
    0.002791101, 2.614083e-05,
  0.009165992, 0.0001769551, 0.0002754912, -1.504133e-08, -1.920862e-05, 
    0.002353766, 0.01235861, 0.02401966, 0.01905287, 0.04123417, 0.04019789, 
    0.08904409, 0.1088389, 0.04255337, 0.01446255, 0.02491829, 0.02809934, 
    0.01325172, 0.01504909, 0.006224941, 0.03409411, 0.07664825, 0.06434414, 
    0.01548519, 0.01463967, 0.01029567, 0.01753862, 0.07621354, 0.009493352,
  -6.177848e-07, 0, 0, 5.786093e-05, 1.352418e-06, 0.007509127, 0.03215427, 
    0.1077718, 0.01905534, 0.06849083, 0.06487449, 0.07164147, 0.04580056, 
    0.0002884796, 0.0001018628, 0.001611153, -2.039054e-05, 0.00261401, 
    0.003004499, 4.482733e-05, 0.0006321049, 0.01768014, 0.03510291, 
    0.006836913, -3.000224e-07, 1.663259e-05, -6.276343e-05, 0, 0.0006643804,
  0, -6.416773e-05, 0, 0, -1.199801e-08, -1.628527e-06, 0.004942433, 
    0.003923525, 0.05774356, 0.03435761, 0.05643308, 0.04683463, 0.005241357, 
    0.000189635, 0.0001651924, 0.003431049, 0.001114294, 0.001494862, 
    -3.280752e-05, 0, 0, 0.005170768, 0.001450587, 0.001641187, 0.003422883, 
    0.000397413, -9.06501e-06, 0, -7.581598e-12,
  -1.636708e-07, 0.004599484, 0.001771324, -2.590847e-13, 0.0003098213, 
    -1.644212e-05, 3.814262e-05, 5.177957e-05, 0.00328213, 0.006886925, 
    0.02099293, 0.02960241, 0.04336242, 0.02777693, 0.01329964, 0.002912525, 
    8.034788e-05, 9.493521e-05, 0.0004695713, 0, 0, 0.009292857, 0.01945645, 
    0.008436215, 0.01338954, 0.01624568, 0.0005343659, -3.693828e-05, 
    -5.063283e-06,
  -4.630855e-06, -5.749325e-06, 0.001371373, -3.294981e-05, 2.106634e-06, 
    0.0003799633, -1.54359e-06, -8.969941e-05, 0.0006326903, 0.004850264, 
    0.004228243, 0.008101463, 0.01352674, 0.006679395, 0.001403156, 
    0.003406956, -7.161299e-06, -2.055863e-06, 0.0006788562, -2.117385e-05, 
    0.008052219, 0.009234929, 0.01133475, 0.009207888, 0.005763085, 
    0.005955168, 0.005932487, 0.00273489, -2.249867e-06,
  0, -3.747641e-06, 9.509175e-05, -3.144643e-05, 0, -1.844873e-06, 0, 0, 
    0.0004577705, 0, 0, -1.793615e-06, 0.00119152, 6.630094e-05, 
    -1.756199e-05, 0, -2.663874e-05, 0, 0, -6.109159e-06, 0.0009878565, 
    0.001910155, -0.000210629, -3.067309e-06, 0.001872441, 0, -5.137253e-10, 
    0, 0,
  0, 0, 0, 0, 0, -4.460503e-05, 0, 0.001823122, 0, 0, -4.155643e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -8.543058e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001159981, 
    -7.050269e-06, 0, 0, -7.311527e-06, 0.001355232, 0.0004938677, 0, 0, 0, 
    0, 0, 0, 0, 0,
  -2.992444e-05, 0.002460955, -7.645578e-06, 0.001562531, 0.002029476, 
    0.000402743, 0.0001828979, 0.001496291, 0.0002669922, 0.0003735848, 0, 0, 
    0.0001046889, -8.122637e-06, 0.001364386, -1.035716e-06, 0.0001056856, 
    -6.544406e-06, 0.001000319, 0.0007128025, 0.002316982, 6.271443e-05, 
    0.001698015, 0.001006925, -2.528596e-06, 0, 0.005620386, 0.002381946, 
    0.0002908675,
  6.343373e-05, 0, 0.0004255668, 0.001583441, 0.01472739, 0.003689396, 
    0.002490229, 0.0007796268, 0.0004344865, 1.005033e-11, 0.002050871, 
    -4.75983e-05, 0.001116208, 0.001014488, 0.0008275529, 0.01239618, 
    0.006689831, 0.007148894, 0.01190981, 0.01433801, 0.02334089, 0.02198751, 
    0.003980986, 0.01190461, 9.554509e-05, 0.01141537, 0.01507543, 
    0.00538992, 0.00553109,
  -5.035219e-06, 0, 0.001297302, 0.004685367, -6.647845e-05, 5.60799e-05, 
    -1.430722e-07, 0, -3.443157e-09, 0.001908344, 0.002652133, 0.00393272, 
    3.703446e-05, 0.007612532, 0.01827542, 0.03561539, 0.02208247, 
    0.02468027, 0.04419513, 0.02677996, 0.00992428, 0.0004068377, 
    -6.344168e-08, 0.0004029504, 5.62165e-05, 0.009472212, 0.00193687, 
    -1.363335e-05, -1.873128e-06,
  -6.752956e-10, 0.0001552894, -1.374523e-09, -5.239782e-10, 9.780306e-06, 
    5.133765e-06, -5.115806e-06, -2.407283e-08, 0.0001863891, -4.289905e-05, 
    1.597186e-07, 1.023209e-05, 1.170576e-05, 0.004256655, 0.0200689, 
    0.01742752, 0.01853665, 0.003600765, 0.002624778, 0.006692849, 
    1.930407e-05, 1.568835e-07, 6.033643e-05, 0.0005384331, 1.052073e-05, 
    -1.208256e-11, -1.319299e-07, 4.181057e-05, 2.047991e-06,
  0, 8.636654e-06, 0, -9.12246e-08, 0.0202118, 0.01843179, 0.02917121, 
    0.05909222, 0.05945282, 0.01733937, 0.02566784, 0.04097663, 0.1176497, 
    0.1355338, 0.1030832, 0.1324401, 0.07295451, 0.003506589, 0.004354395, 
    -2.746432e-05, 3.575314e-05, 0.0001370719, -1.237593e-07, 0.001456663, 
    0.0001235375, -3.31835e-05, 1.378038e-05, 7.411538e-06, 0.001217154,
  0.001555762, 0.009663431, 0.002271663, -1.380737e-05, -1.902586e-05, 
    0.01135978, 0.03350063, 0.0767093, 0.05285776, 0.06573235, 0.1222269, 
    0.1748721, 0.2811428, 0.1395193, 0.1646583, 0.05600218, 0.01395412, 
    0.01583234, 0.0003584309, 5.931332e-05, 0.008155623, 0.01828671, 
    0.02373384, 0.1044102, 0.05493404, 0.002329869, 0.002018143, 0.01983993, 
    0.01746684,
  0.03610371, 0.004965425, 0.0007990247, -7.354563e-06, 0.004316649, 
    0.1150421, 0.2251554, 0.508709, 0.3945862, 0.3015647, 0.2186195, 
    0.2687762, 0.3410273, 0.1868594, 0.1107855, 0.1179845, 0.1079553, 
    0.04940706, 0.03929134, 0.02481627, 0.08791558, 0.2224136, 0.1862592, 
    0.08809052, 0.04519596, 0.0164238, 0.0341715, 0.1537232, 0.03792594,
  0.004000092, 0.0001357113, 1.006723e-05, 0.00348817, 0.008866834, 
    0.0547806, 0.1083899, 0.2731764, 0.1971861, 0.2202746, 0.2185834, 
    0.1818898, 0.1264929, 0.01435943, 0.0006841801, 0.007995457, 0.003123283, 
    0.009694556, 0.01712709, 0.00296936, 0.01783618, 0.0829688, 0.07520693, 
    0.02243223, 0.0004087309, 0.0002023739, -5.926027e-05, 0.0001881232, 
    0.002254519,
  0.0008933598, 0.0006648883, -7.579021e-06, -1.56905e-07, 0.000168593, 
    -2.497533e-05, 0.03840818, 0.006842926, 0.102188, 0.1662296, 0.2260637, 
    0.1673707, 0.09599026, 0.03504319, 0.01410334, 0.01262829, 0.008797533, 
    0.004394183, 0.0003791954, -1.526382e-06, 0, 0.04265796, 0.02770037, 
    0.006101067, 0.009559225, 0.0006108973, 0.0004379742, -4.251e-06, 
    -6.79989e-06,
  0.002961414, 0.01653049, 0.003145472, 0.0001269385, 0.0008928149, 
    0.001285589, 0.001753582, 0.01112066, 0.01681244, 0.01263333, 0.05467737, 
    0.09972273, 0.1638709, 0.08384759, 0.03381483, 0.01513169, 0.005919962, 
    0.003056623, 0.001357144, -4.038217e-05, -1.915631e-05, 0.01739193, 
    0.02870307, 0.01759225, 0.02094681, 0.02800289, 0.004534383, 
    -3.754312e-05, -9.888398e-06,
  0.0002534325, 3.131378e-05, 0.01217353, 0.002334456, 0.0005868633, 
    0.001225984, -5.618178e-05, 0.0007677729, 0.002686293, 0.01049544, 
    0.0102337, 0.009855358, 0.02132039, 0.01280214, 0.002736335, 0.008085615, 
    0.002232273, 0.001891279, 0.002185388, 5.014362e-05, 0.01639193, 
    0.01482794, 0.01716956, 0.01625574, 0.0126181, 0.01439366, 0.0168598, 
    0.009124337, 0.0004515399,
  -8.579984e-06, 0.001261232, 0.000169156, 0.001067194, 2.95368e-05, 
    0.000780624, -4.370246e-05, -9.942516e-09, 0.00164969, 0, 0.000895102, 
    0.0002967125, 0.004516476, 0.0007950506, -7.424831e-05, 0, 0.0003988482, 
    0.0006551255, 0, -3.042198e-05, 0.004648111, 0.004271191, 0.002306144, 
    3.152666e-05, 0.004810027, -9.044008e-05, 0.0002120122, 5.754276e-06, 
    -2.675483e-05,
  0, 0, 0, 0, 0, 0.001359328, -4.995926e-05, 0.002495302, 0.0005520037, 0, 
    -1.246693e-06, 0, 0, 0, 0, 0, 0, 0, -4.639214e-06, -4.424308e-06, 
    -0.0002589387, 7.907455e-05, 0, 0, -1.83012e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -2.655955e-06, 0, -6.433085e-07, 0.0001397973, 0, 3.271451e-05, 0, 0, 
    9.173725e-05, 5.058232e-05, -1.88007e-05, -0.0001108662, 0.0002001067, 
    -2.947192e-05, -7.36615e-06, 0, 2.38167e-05, 0.003343713, 0.002320826, 
    -2.220292e-05, 0.001748552, -8.977393e-06, 0, 0, 0, 0, 0,
  -0.0001154914, 0.005294361, 0.000378617, 0.001837207, 0.003344813, 
    0.001352044, 0.001393093, 0.00190116, 0.001838028, 0.002241823, 
    0.0008532473, 0.002153685, 0.001766645, 0.002303476, 0.002637761, 
    -2.383061e-05, 0.001083181, 0.002005741, 0.003828482, 0.004487661, 
    0.005568756, 0.001056793, 0.002050648, 0.002920788, 0.001365177, 
    -4.535072e-05, 0.01204853, 0.008497481, 0.0009272464,
  0.00198638, -0.0002035226, 0.006389925, 0.004572855, 0.0231701, 0.01411073, 
    0.005207099, 0.00357931, 0.003841814, 0.001570734, 0.007984854, 
    0.002171876, 0.002206485, 0.005484303, 0.004655308, 0.0253781, 0.0206609, 
    0.01889038, 0.03105068, 0.03316962, 0.03770052, 0.04750938, 0.01383591, 
    0.02226136, 0.001646653, 0.01973363, 0.02809358, 0.01292959, 0.007038986,
  0.003607049, 0.0001733227, 0.002389345, 0.007042609, 0.000262293, 
    0.0008821451, -1.678745e-06, -2.213081e-08, -6.539142e-06, 0.001333869, 
    0.01341647, 0.02234103, 0.001175359, 0.01327199, 0.03217334, 0.06754201, 
    0.04528562, 0.05723258, 0.08629726, 0.05122264, 0.01553665, 0.00823533, 
    0.0004111068, 0.00397956, 0.0060582, 0.02065095, 0.009470556, 
    0.001006408, 0.002652659,
  0.006612001, 0.001303965, 3.327062e-05, 2.116307e-06, 0.006616096, 
    -5.743294e-05, 0.000396443, -9.419231e-06, -0.0001090198, -5.205139e-05, 
    9.318172e-06, 3.522041e-06, 6.786e-05, 0.00316747, 0.05440306, 0.0776976, 
    0.06470253, 0.03275818, 0.02691935, 0.02113479, 0.0008692994, 
    1.447616e-05, 0.0005985461, 0.03037917, 0.0006617376, 0.0001898723, 
    0.004695707, 0.0004770347, 0.003621416,
  0.0009164797, 0.01452831, 0.0003269614, 1.019663e-05, 0.04166686, 
    0.04928944, 0.04455503, 0.08190793, 0.08550492, 0.01382337, 0.03012415, 
    0.02313387, 0.1088131, 0.1206173, 0.09456503, 0.1241694, 0.06038015, 
    0.004519949, 0.01244866, 0.0003082869, 0.001934322, 0.007223248, 
    0.004608553, 0.01826333, 0.003100181, 0.00225849, -2.659772e-05, 
    0.004847004, 0.001686966,
  0.08627836, 0.167485, 0.2038454, 0.003017943, 0.00200669, 0.06373584, 
    0.1899942, 0.1551999, 0.2326912, 0.2771334, 0.09472834, 0.1470191, 
    0.2490177, 0.116453, 0.1348373, 0.02682274, 0.01689185, 0.01309297, 
    2.221999e-05, 0.00124945, 0.02803127, 0.04018011, 0.06610195, 0.2605864, 
    0.1220452, 0.0278825, 0.012814, 0.08038587, 0.0712441,
  0.1914195, 0.1103836, 0.04915594, -1.026044e-05, 0.02149672, 0.1590078, 
    0.2478727, 0.3924251, 0.3555948, 0.2231066, 0.1783792, 0.2265985, 
    0.2692975, 0.1634047, 0.1070928, 0.1678826, 0.121776, 0.06079703, 
    0.06148716, 0.03357606, 0.08448452, 0.2113955, 0.3266224, 0.1739055, 
    0.1350662, 0.0907557, 0.05961214, 0.2373103, 0.2283227,
  0.07761826, 0.003156261, 0.01878332, 0.001888756, 0.005638511, 0.05343251, 
    0.1075988, 0.2297177, 0.1536862, 0.1727426, 0.1840105, 0.1495496, 
    0.1163146, 0.06566087, 0.0493648, 0.05171616, 0.05147861, 0.05578707, 
    0.060126, 0.03674843, 0.01414641, 0.1052008, 0.1688046, 0.2397923, 
    0.08063465, 0.02219664, 0.004732005, 0.01836925, 0.03545997,
  0.02168529, 0.01998637, 0.005831478, 0.0005378199, 0.0001017874, 
    -6.57401e-06, 0.03613917, 0.01331946, 0.1650125, 0.1710576, 0.2893403, 
    0.2289398, 0.1740361, 0.1286294, 0.1417413, 0.1058292, 0.07025184, 
    0.02894441, 0.004824925, 0.006758746, -3.819716e-05, 0.1002745, 0.146895, 
    0.169105, 0.1664204, 0.05283216, 0.005870077, 0.004142163, 0.002762764,
  0.006947326, 0.04068837, 0.008679461, 0.000917068, 0.007985631, 0.01070591, 
    0.007427699, 0.02919948, 0.06528269, 0.0311827, 0.101586, 0.1654907, 
    0.2567797, 0.1808441, 0.1012623, 0.1257353, 0.07314599, 0.03752586, 
    0.01239782, 1.326287e-05, 0.0001080266, 0.04118831, 0.1059496, 
    0.05389071, 0.07497464, 0.07071941, 0.02854102, 0.01316916, 0.005962305,
  0.009343309, 0.0001797926, 0.02289693, 0.005004456, 0.001321412, 
    0.006647079, 0.003347048, 0.002324021, 0.007604854, 0.0207008, 
    0.02070118, 0.01863888, 0.03786216, 0.05292616, 0.02799708, 0.0260352, 
    0.01406198, 0.02794449, 0.01158687, 0.002436664, 0.02997145, 0.0240301, 
    0.03364775, 0.02276951, 0.02845929, 0.03406849, 0.02766028, 0.02812505, 
    0.01968983,
  -5.104858e-05, 0.004184382, 0.002045307, 0.003332939, 0.0003568042, 
    0.0007488749, 0.001229479, 5.621234e-05, 0.002043124, -1.971716e-05, 
    0.002115583, 0.002576184, 0.008027902, 0.007234506, 0.003857283, 
    1.98169e-06, 0.004444737, 0.001602302, -9.139809e-05, 0.001282225, 
    0.01208621, 0.01172386, 0.008127142, 0.002639626, 0.007343732, 
    0.002248987, 0.002270749, 0.003583841, 0.0006014656,
  -1.989662e-05, 0, 0, 0, 0.001403101, 0.001845681, -7.272191e-05, 
    0.003534951, 0.001366428, 0, 0.0002013872, 0, 0, 0, 0, 0, 0.0006773873, 
    -1.364052e-05, -8.722619e-06, -0.0001668912, 0.003688711, 0.0004582191, 
    0, 0, 0.001302731, 0.001299507, 0, -9.817068e-05, -0.0001538094,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.086893e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.78995e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  2.792961e-06, 0, -1.826563e-06, -1.301365e-05, 8.507282e-05, 0.0005596649, 
    0, 0.0003843581, -4.752761e-05, 0, 0.0009421736, 0.001344334, 
    0.0005019034, -0.0001752969, 0.0005876801, -4.112997e-05, 0.001087274, 0, 
    0.003325368, 0.006670793, 0.008374691, 0.005375728, 0.005485085, 
    0.002497588, 0.0004102475, -1.646566e-05, -6.657897e-06, 0, 0,
  0.003855977, 0.008783452, 0.003766047, 0.00325339, 0.005670888, 
    0.005106787, 0.00389842, 0.006483917, 0.00777618, 0.004789727, 
    0.003972463, 0.008354248, 0.007877841, 0.005345823, 0.008123439, 
    0.001617974, 0.01057954, 0.00891698, 0.01082553, 0.0131665, 0.01299172, 
    0.01257342, 0.007906456, 0.006601739, 0.004481177, 0.001214851, 
    0.02226668, 0.03307448, 0.003562596,
  0.006392963, 0.001908586, 0.01434842, 0.02418792, 0.03421647, 0.02183021, 
    0.01330622, 0.01529679, 0.01724149, 0.008185223, 0.01252709, 0.008008205, 
    0.004489703, 0.01820371, 0.01832546, 0.05024801, 0.037051, 0.0459885, 
    0.0580607, 0.05891952, 0.06507183, 0.08588968, 0.0340147, 0.04902854, 
    0.007643984, 0.03632247, 0.04789443, 0.03238047, 0.01414161,
  0.006318895, 0.0007055238, 0.003390371, 0.01377627, 0.00590447, 0.02278492, 
    0.001335241, -4.927924e-05, 0.000377468, 0.001519894, 0.03290403, 
    0.05253833, 0.01431007, 0.03488198, 0.07672378, 0.09499823, 0.08876599, 
    0.1226134, 0.1932015, 0.1624953, 0.09724906, 0.02620544, 0.02167126, 
    0.03931097, 0.03744674, 0.03075709, 0.0498946, 0.01619551, 0.00436339,
  0.0001958438, 3.01898e-05, 3.532061e-05, 1.176801e-06, 0.002324833, 
    -4.401224e-06, 2.333487e-05, -4.481635e-07, -8.88721e-05, 0.0001013365, 
    -8.721878e-06, 3.55413e-06, 1.868727e-05, 0.002444701, 0.04842637, 
    0.06872944, 0.09098314, 0.04048929, 0.06157867, 0.02665677, 0.0004771236, 
    -1.037575e-05, 4.036225e-05, 0.004156727, 0.001801491, 0.004904923, 
    0.004582644, 1.980886e-05, 0.005972472,
  3.981361e-05, 0.0001189778, 1.904102e-05, -3.329227e-06, 0.03264026, 
    0.03724987, 0.03645626, 0.07007255, 0.07257295, 0.01129506, 0.02378689, 
    0.01464764, 0.09846232, 0.1022108, 0.07334377, 0.09982846, 0.04322827, 
    0.0006088733, 0.002924226, 6.465465e-05, 3.203034e-05, 0.003227313, 
    0.009496854, 0.0117095, 0.001735817, 0.0003041809, -3.521816e-05, 
    7.279473e-05, 7.65618e-05,
  0.04155938, 0.1337344, 0.1085765, 0.0007391826, 0.0006594657, 0.02992842, 
    0.1101289, 0.09348738, 0.1979205, 0.23845, 0.05952178, 0.1181625, 
    0.2311082, 0.09280741, 0.1014641, 0.0138675, 0.01823688, 0.01190365, 
    1.006823e-05, 0.0001248628, 0.008770672, 0.02283325, 0.0708245, 
    0.2340552, 0.08750039, 0.01343638, 0.01019349, 0.0434866, 0.02133915,
  0.1412608, 0.08622771, 0.0480131, 0.007303428, 0.01469341, 0.1142043, 
    0.1720803, 0.2594207, 0.3115357, 0.1711856, 0.1457623, 0.1961037, 
    0.2245968, 0.1241172, 0.08098958, 0.1268949, 0.09072552, 0.0375244, 
    0.0434485, 0.01788917, 0.06712188, 0.1793635, 0.288302, 0.1222725, 
    0.08765013, 0.06058744, 0.04079445, 0.2091685, 0.1726458,
  0.1017658, 0.0201322, 0.01961386, 0.00144714, 0.002106498, 0.0564624, 
    0.1120732, 0.2054486, 0.1301242, 0.145401, 0.1598261, 0.1237517, 
    0.09424758, 0.04097387, 0.03414002, 0.04214271, 0.05166399, 0.06728031, 
    0.06178363, 0.01479494, 0.007983682, 0.08400805, 0.1396347, 0.1881879, 
    0.05849448, 0.01263354, 0.003783535, 0.01782916, 0.03478222,
  0.0602832, 0.08290966, 0.01147589, 0.01501343, 0.002648095, 0.0014721, 
    0.03562991, 0.05027001, 0.2592817, 0.1468655, 0.2746119, 0.2150766, 
    0.1454734, 0.1083434, 0.1420937, 0.1110821, 0.1047522, 0.03314155, 
    0.02322238, 0.01930405, 0.01059734, 0.1063239, 0.1061609, 0.1444732, 
    0.1750697, 0.1086686, 0.04611742, 0.006514495, 0.008003818,
  0.04332988, 0.09320546, 0.02563265, 0.0137619, 0.06161983, 0.03858673, 
    0.0175178, 0.1232302, 0.1668183, 0.0873719, 0.1282425, 0.1677407, 
    0.280605, 0.2094111, 0.1374486, 0.2327785, 0.2105073, 0.1104822, 
    0.03325566, 0.003680052, 0.001092136, 0.113813, 0.1112914, 0.08215037, 
    0.1671053, 0.1546721, 0.09597901, 0.08283511, 0.0454501,
  0.0399594, 0.001899633, 0.0403356, 0.01900349, 0.03160057, 0.01732808, 
    0.01181218, 0.01228145, 0.01794974, 0.06803068, 0.06848767, 0.08568308, 
    0.06672094, 0.06775881, 0.06493718, 0.09042235, 0.1045203, 0.1440228, 
    0.07476953, 0.004589683, 0.04294488, 0.0821825, 0.08282591, 0.05770601, 
    0.08925262, 0.1123411, 0.1224791, 0.111922, 0.08621908,
  0.01723569, 0.007064107, 0.004698283, 0.00580683, 0.003079905, 0.00184855, 
    0.01067605, 0.0004953687, 0.005161296, 0.0005728986, 0.006225583, 
    0.01370595, 0.01461473, 0.02057414, 0.01563597, 0.00852043, 0.03445575, 
    0.02463265, 0.001363583, 0.00352031, 0.02974499, 0.03544037, 0.02629457, 
    0.00924981, 0.02958138, 0.01102836, 0.01679633, 0.03177229, 0.0314998,
  0.005969089, 0.002716527, -2.114314e-06, 1.500217e-05, 0.003799079, 
    0.002226724, 0.0006124569, 0.004571003, 0.007639687, 0.001700453, 
    0.0003898371, -1.129087e-09, -4.153447e-06, 0, -1.705562e-07, 
    -1.278894e-06, 0.0006879761, 0.01447683, 0.01393087, 0.009259463, 
    0.01987145, 0.001109893, -4.051781e-05, -1.972843e-05, 0.002384235, 
    0.00322207, -6.482827e-07, 0.001513003, 0.01025358,
  -9.172585e-07, -7.573411e-06, 0, 0, 0, 0, 0, -1.11143e-05, 7.182722e-07, 
    -3.15952e-08, 1.032912e-06, -5.193862e-05, -1.855876e-05, 0, 0, 
    3.270207e-06, -3.061486e-06, -1.879721e-10, 0, 0, 3.625255e-09, 
    1.861206e-05, 0, 0, 0, 0, 0, -2.224502e-07, 7.339267e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.255574e-05, 0, 0, 0, 0, 0, 0, -1.87331e-05, 4.757197e-06, 
    0.0005962481, 0, 0, 0, -2.169413e-06, -2.567656e-05, 0, 0, 0, 0, 
    0.001077597, 9.170875e-05, 0, 0, 0,
  0.001132533, 0.003177258, 0.001196131, 0.002132907, 0.0004285698, 
    0.002274065, 0.0002634856, 0.003425937, -0.0001013469, -2.785992e-07, 
    0.0009404821, 0.00594915, 0.002994195, 0.0001478257, 0.001706544, 
    0.002174987, 0.003473727, 0.0001581252, 0.01210147, 0.01425566, 
    0.0166107, 0.01647791, 0.0211174, 0.006187439, 0.003452384, 0.001211767, 
    0.001095619, 0.0008038571, -4.287955e-05,
  0.02047989, 0.01673126, 0.009986974, 0.00519944, 0.01331299, 0.008883377, 
    0.009442572, 0.01450511, 0.01449029, 0.01261942, 0.00951633, 0.01833786, 
    0.02231328, 0.0104993, 0.01503365, 0.01057668, 0.04330908, 0.03891183, 
    0.03437136, 0.03563331, 0.04006211, 0.04327264, 0.03849221, 0.01677063, 
    0.02316898, 0.01603538, 0.04927748, 0.06470127, 0.02149865,
  0.06192763, 0.03222286, 0.03445097, 0.04624058, 0.05036692, 0.04661987, 
    0.03660345, 0.03733529, 0.03784896, 0.01316401, 0.03042639, 0.0256547, 
    0.01260248, 0.03507757, 0.03902368, 0.08024656, 0.0998218, 0.09821285, 
    0.1215013, 0.1172015, 0.1410444, 0.1612016, 0.08812991, 0.0886078, 
    0.0805434, 0.1005138, 0.1211477, 0.1016396, 0.08067843,
  0.02664656, 0.01820771, 0.006000012, 0.03349657, 0.02860915, 0.03473257, 
    0.009955428, 0.000589401, 0.005802637, 0.01035679, 0.04144732, 
    0.05276153, 0.02233662, 0.04768525, 0.08288938, 0.1096379, 0.1198406, 
    0.1436151, 0.2269838, 0.1888837, 0.07634898, 0.04426614, 0.02864368, 
    0.0539493, 0.03960824, 0.06254944, 0.09706551, 0.07436232, 0.0303168,
  0.0001369849, 6.865398e-06, 0.0001372506, 2.445483e-07, 0.001188022, 
    0.0006200227, -2.558717e-05, 1.897436e-06, 0.001072792, -1.047748e-05, 
    0.0005563793, 7.053604e-06, -2.16434e-05, 0.005636674, 0.04665456, 
    0.05974027, 0.07736137, 0.03419778, 0.03039604, 0.01789727, 0.0003139688, 
    5.004895e-06, 2.362334e-06, 0.0001440164, 0.0002807464, 0.006934641, 
    0.008561375, 0.00154071, 0.003433348,
  7.70806e-06, 1.884814e-05, 4.119689e-06, -5.791668e-06, 0.03257029, 
    0.02817391, 0.02790834, 0.05852848, 0.07095025, 0.01570436, 0.02369311, 
    0.01589091, 0.0901426, 0.08487296, 0.06066183, 0.08472043, 0.03921976, 
    0.0003001193, 9.885224e-05, 3.310011e-05, 7.589164e-07, 2.495036e-05, 
    0.004890111, 0.005356785, -2.280688e-05, -1.875492e-05, 1.093512e-05, 
    9.260584e-06, 9.502885e-06,
  0.01223908, 0.104356, 0.06355061, 0.0003152182, 0.0007815792, 0.02764752, 
    0.0785704, 0.07845204, 0.1568725, 0.2119519, 0.0468497, 0.1035852, 
    0.2141566, 0.08309156, 0.08355932, 0.01334111, 0.01943533, 0.01293269, 
    9.781777e-06, 0.001165665, 0.001890187, 0.01343122, 0.08127626, 
    0.1902346, 0.06913398, 0.01744141, 0.01168778, 0.02189534, 0.00722601,
  0.1299741, 0.08758377, 0.04834229, 0.0008552513, 0.01741246, 0.06349738, 
    0.1353367, 0.145908, 0.2719003, 0.1398194, 0.1198361, 0.1784026, 
    0.1990883, 0.105001, 0.07415044, 0.1018871, 0.08569135, 0.02879612, 
    0.03830298, 0.01632144, 0.06373259, 0.1731003, 0.256716, 0.1027375, 
    0.06620485, 0.03796976, 0.03190666, 0.1786998, 0.1534019,
  0.1048426, 0.02564083, 0.008655581, 0.001254424, 0.004721734, 0.0551219, 
    0.1049725, 0.1962361, 0.1186927, 0.118376, 0.1234001, 0.113039, 0.08162, 
    0.03563228, 0.02816504, 0.02893732, 0.03214185, 0.05182838, 0.04722449, 
    0.002774886, 0.00876838, 0.0666831, 0.1372594, 0.1693429, 0.05279318, 
    0.007524216, 0.003166383, 0.01540466, 0.02908798,
  0.05460945, 0.07447891, 0.007508602, 0.01195536, 0.002059631, 0.005489809, 
    0.02749088, 0.07685746, 0.2798647, 0.126728, 0.2543454, 0.1950131, 
    0.1260475, 0.1072868, 0.125582, 0.09616379, 0.08751576, 0.04091701, 
    0.03164381, 0.01560427, 0.0468912, 0.07909628, 0.07460092, 0.125191, 
    0.1540442, 0.08536817, 0.02344728, 0.0103453, 0.01313636,
  0.1047983, 0.1266125, 0.04768096, 0.06473818, 0.07341994, 0.05556734, 
    0.03052443, 0.2136292, 0.2063603, 0.1426357, 0.151216, 0.1700551, 
    0.2722274, 0.2068477, 0.121757, 0.2153041, 0.2242781, 0.1321922, 
    0.04600467, 0.01641329, 0.01705626, 0.1013779, 0.08716689, 0.08474328, 
    0.134485, 0.1345213, 0.1014757, 0.09324098, 0.06196966,
  0.09834541, 0.0579647, 0.1173072, 0.09670796, 0.1090616, 0.1106337, 
    0.07134574, 0.02896622, 0.06473047, 0.1177275, 0.1386356, 0.173726, 
    0.1078968, 0.1007491, 0.1131603, 0.1616177, 0.2120798, 0.2181072, 
    0.1313982, 0.02849413, 0.1315696, 0.1111999, 0.08822479, 0.08507735, 
    0.1258975, 0.1772755, 0.1890689, 0.1659708, 0.1780902,
  0.1216251, 0.05180568, 0.03422623, 0.06033385, 0.05417068, 0.06004834, 
    0.05666799, 0.05339549, 0.05964067, 0.03215214, 0.06284048, 0.06241322, 
    0.05162626, 0.1157441, 0.08008549, 0.05913715, 0.06511223, 0.059491, 
    0.02993406, 0.07867783, 0.09459554, 0.1097335, 0.07485568, 0.04679753, 
    0.07445557, 0.03919129, 0.06108882, 0.147164, 0.1172082,
  0.07321643, 0.06890607, 0.01997236, 0.018998, 0.0317334, 0.03113342, 
    0.03449848, 0.01981772, 0.04750044, 0.05235383, 0.03862946, 0.05223604, 
    0.01717759, 0.0158964, 0.01544427, 0.02111111, 0.02926029, 0.03811378, 
    0.0299589, 0.05725769, 0.06330349, 0.01546447, 0.003884112, -0.001341583, 
    0.01312856, 0.003860184, -2.083462e-05, 0.01423078, 0.04701324,
  0.01401579, 0.01860292, 0.009983006, 0.004759009, -0.000159548, 
    -3.684371e-06, -0.0004897203, 0.001982987, 9.447051e-05, 0.005962224, 
    0.0105415, 0.009404113, 0.008845788, 0.007721889, 0.005251731, 
    0.003833793, 0.0001707303, 7.473529e-05, 4.819228e-05, -1.340225e-05, 
    -0.0001319692, 0.001702623, -8.460083e-06, -6.125695e-05, -2.427522e-05, 
    -4.759307e-06, -3.295399e-05, 0.002658901, 0.01013856,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.002694257, 0.0001244202, 0, 0, 0, -0.0001035055, 0.001193862, 0, 0, 
    -9.764664e-06, -5.326626e-07, 0, -3.74662e-05, 8.600084e-06, 0.005179434, 
    0.001151335, -4.035875e-06, 0.0004962659, 0.002023027, 0.002236143, 
    0.0003154006, 0.001942162, -3.315589e-05, 0.00279488, 0.002902434, 
    0.002495453, 0.0002723642, 0, 0.0003432884,
  0.02083531, 0.01212856, 0.01244659, 0.01407599, 0.00759731, 0.01141631, 
    0.00377031, 0.01185758, 0.003914685, 0.002965271, 0.008187798, 
    0.01290965, 0.0164851, 0.01521269, 0.03005714, 0.01743174, 0.009438949, 
    0.007666117, 0.03294839, 0.03095369, 0.03192091, 0.03443806, 0.04619725, 
    0.02830228, 0.02310058, 0.01444477, 0.009308103, 0.007905983, 0.00872697,
  0.1097524, 0.09859306, 0.07572483, 0.05341629, 0.05865663, 0.07242591, 
    0.04389419, 0.06198841, 0.03995203, 0.03873546, 0.03620399, 0.06057895, 
    0.06282526, 0.03750797, 0.05922905, 0.05886083, 0.1181118, 0.1168297, 
    0.1054512, 0.1142249, 0.1029631, 0.09352034, 0.08672719, 0.03713791, 
    0.08022836, 0.08302215, 0.09568328, 0.1479863, 0.09285215,
  0.1329326, 0.08777383, 0.077876, 0.1062869, 0.1173534, 0.1016876, 
    0.08347173, 0.08948763, 0.09233205, 0.05076799, 0.07232486, 0.05650318, 
    0.0617188, 0.1072117, 0.08158602, 0.1021443, 0.121838, 0.1273799, 
    0.1402432, 0.1402062, 0.1613834, 0.1882381, 0.1409135, 0.1266908, 
    0.1075315, 0.1401156, 0.1488785, 0.140115, 0.1315112,
  0.03130793, 0.01744793, 0.01241414, 0.03155175, 0.01841157, 0.02806611, 
    0.01106174, 0.002473043, 0.01387189, 0.02257992, 0.06451476, 0.06790652, 
    0.02668577, 0.046034, 0.1043006, 0.1383096, 0.1269488, 0.1359734, 
    0.2062757, 0.189901, 0.04753936, 0.04095794, 0.03892585, 0.02942774, 
    0.03872668, 0.05490046, 0.09139136, 0.04927823, 0.02503931,
  -8.55788e-07, -1.701183e-05, 0.002259007, -6.965305e-09, 0.001676578, 
    0.004292319, -3.66649e-07, -2.28521e-06, 0.01116252, 0.0005790135, 
    0.001684737, 0.00168001, -3.687868e-05, 0.01601984, 0.05086981, 
    0.05745203, 0.05181894, 0.03460366, 0.02486226, 0.009623502, 
    9.647077e-05, 4.716621e-08, 9.359263e-08, 0.0002835683, 0.000467577, 
    0.003566645, 0.008008303, 0.0122535, 0.001032282,
  4.032866e-06, 4.86514e-06, 3.788798e-06, -3.438079e-05, 0.04045669, 
    0.02572714, 0.0243612, 0.04020112, 0.0639616, 0.02814043, 0.02179624, 
    0.01657165, 0.09100497, 0.07344247, 0.05633198, 0.06596551, 0.03328946, 
    0.0003462984, 5.690151e-05, 4.839529e-05, 2.18173e-08, 6.918827e-07, 
    0.001711741, 0.00133298, -2.137267e-05, 4.694634e-05, 1.186146e-06, 
    1.790232e-05, 3.264443e-06,
  0.008434105, 0.07762358, 0.0372609, 0.0005281472, 0.0006229469, 0.02712918, 
    0.05529941, 0.06226446, 0.119157, 0.1821109, 0.03410865, 0.08154202, 
    0.1933144, 0.0660575, 0.07649355, 0.008966688, 0.02740686, 0.01245601, 
    3.107392e-06, 0.0004803232, 2.929372e-06, 0.006049726, 0.0561363, 
    0.1469355, 0.05803912, 0.02808008, 0.02010691, 0.01588622, 0.003037507,
  0.1120348, 0.09627859, 0.05637695, -4.354843e-05, 0.01393434, 0.04009078, 
    0.1155356, 0.07303212, 0.2221619, 0.1111329, 0.1050108, 0.147181, 
    0.1688429, 0.09721918, 0.06953626, 0.06957698, 0.07821892, 0.01811165, 
    0.03801134, 0.01454055, 0.05909682, 0.1520995, 0.2010116, 0.07062432, 
    0.05080676, 0.02206838, 0.02698455, 0.1567558, 0.1242017,
  0.0918266, 0.01702999, 0.0042098, 0.0003324016, 0.007521354, 0.06018271, 
    0.1040741, 0.1732876, 0.1098362, 0.10545, 0.1115007, 0.102546, 
    0.06047439, 0.02350608, 0.02373322, 0.01727508, 0.01236008, 0.01750936, 
    0.04163761, 0.0003507872, 0.006135487, 0.05276147, 0.1165856, 0.1437511, 
    0.04168572, 0.007755765, 0.002792284, 0.01769269, 0.03113808,
  0.04537351, 0.06865066, 0.006123972, 0.006958066, 0.0004880413, 
    0.005787536, 0.02603842, 0.07556847, 0.2676369, 0.1117745, 0.2382654, 
    0.1870074, 0.11347, 0.1068085, 0.1056865, 0.08639799, 0.07397107, 
    0.03700447, 0.0291248, 0.01116286, 0.02927073, 0.05677515, 0.05028939, 
    0.1060864, 0.1421869, 0.06542509, 0.009420157, 0.01524499, 0.004719274,
  0.1009934, 0.1122971, 0.04736442, 0.07858627, 0.06766176, 0.0499296, 
    0.0669951, 0.1999319, 0.196125, 0.1485123, 0.1627986, 0.1570811, 
    0.249412, 0.188696, 0.1218977, 0.202536, 0.2019173, 0.1135743, 
    0.04381204, 0.04935346, 0.08387531, 0.0799061, 0.06766581, 0.0732767, 
    0.1111531, 0.1244468, 0.08827198, 0.06356159, 0.05898659,
  0.102964, 0.1536439, 0.1192731, 0.08209069, 0.1272293, 0.09937166, 
    0.08374052, 0.06960018, 0.1508142, 0.1828138, 0.1845973, 0.2278716, 
    0.1311818, 0.1281839, 0.1509833, 0.2091479, 0.2134985, 0.2221004, 
    0.1318105, 0.06025364, 0.1685283, 0.08584687, 0.0794079, 0.09616759, 
    0.1479984, 0.185902, 0.184779, 0.1524249, 0.1606477,
  0.1588442, 0.0802632, 0.1088011, 0.09604114, 0.09183151, 0.1008498, 
    0.13288, 0.113957, 0.1210104, 0.06785975, 0.1519483, 0.163606, 0.104106, 
    0.1671662, 0.13575, 0.125623, 0.1190678, 0.1424405, 0.08312527, 
    0.1088741, 0.0988104, 0.1200708, 0.1033227, 0.1033374, 0.1399952, 
    0.09006274, 0.1342334, 0.1909696, 0.1716764,
  0.1622275, 0.1564721, 0.1188147, 0.09415279, 0.1282789, 0.1326918, 
    0.08175859, 0.07462662, 0.109458, 0.09632039, 0.1208136, 0.09394805, 
    0.09678215, 0.0307256, 0.06029146, 0.06779227, 0.08327741, 0.1065582, 
    0.1482595, 0.1410085, 0.1332245, 0.08730797, 0.04502315, -0.00307579, 
    0.09561327, 0.005905824, 0.001456208, 0.1048157, 0.1319011,
  0.0440222, 0.06914793, 0.07224488, 0.03553089, 0.02122048, 0.03509118, 
    0.04595453, 0.07455046, 0.07839934, 0.07465211, 0.09860007, 0.08364737, 
    0.05582526, 0.03674163, 0.03586511, 0.04394914, 0.05106592, 0.03056878, 
    0.02068494, 0.01340454, 0.02370059, 0.04331927, 0.0377856, 0.02302679, 
    0.01119941, 1.520431e-05, -0.0005346542, 0.0146618, 0.03534221,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.14494e-07, -2.178985e-06, 0, 
    -0.0001632166, 0.002009742, 0, 0, 0, 0, 0, -1.753743e-05, 0, 0, 0, 0, 0,
  0.008632009, 0.00535702, 0.002108613, 0.0001570322, -3.375707e-06, 
    -0.0001858099, 0.01262389, -7.107874e-05, 0, -0.0001963384, 
    -1.259755e-05, -3.29849e-05, -0.0002604565, 0.002584138, 0.01965749, 
    0.0131628, 0.008601999, 0.007807675, 0.006612693, 0.009118497, 
    0.01159791, 0.01558345, 0.01180512, 0.0172122, 0.009105443, 0.004457472, 
    0.00587954, 0.006499887, 0.003479803,
  0.05907223, 0.05160637, 0.06816836, 0.07631024, 0.06517612, 0.05738157, 
    0.0764067, 0.07004791, 0.08298507, 0.03198369, 0.03498803, 0.04612011, 
    0.05514669, 0.08185479, 0.08672073, 0.08246405, 0.06548546, 0.06125845, 
    0.1013041, 0.1050262, 0.09320531, 0.09940657, 0.0974554, 0.07151465, 
    0.0779922, 0.06337038, 0.04611807, 0.03601641, 0.05778924,
  0.1449395, 0.1241588, 0.1486554, 0.1310958, 0.1266845, 0.1363225, 
    0.1153263, 0.1201975, 0.09540095, 0.1160188, 0.09307157, 0.145264, 
    0.1235602, 0.152888, 0.1994387, 0.1545212, 0.1827399, 0.1763374, 
    0.1819707, 0.1628405, 0.1657821, 0.1422501, 0.115632, 0.08104298, 
    0.09321012, 0.1512441, 0.1763796, 0.2001455, 0.1182192,
  0.1395447, 0.1030312, 0.1070242, 0.1314025, 0.1233297, 0.1087254, 
    0.08816044, 0.09967628, 0.1060581, 0.06519315, 0.09535012, 0.09928411, 
    0.1004907, 0.1682424, 0.1254772, 0.1464369, 0.1481084, 0.1368379, 
    0.1498869, 0.1384988, 0.1436953, 0.2051032, 0.1483878, 0.1624054, 
    0.103337, 0.1426624, 0.1493816, 0.1341455, 0.1346263,
  0.02937311, 0.01077297, 0.02785873, 0.027092, 0.01566293, 0.01190622, 
    0.002262738, 0.003891643, 0.0156574, 0.02987768, 0.05503892, 0.06526396, 
    0.03301106, 0.04397482, 0.1152847, 0.1468049, 0.1039817, 0.132162, 
    0.1887917, 0.1779673, 0.03248203, 0.030926, 0.03050648, 0.02841796, 
    0.0401745, 0.05215936, 0.0723106, 0.03388567, 0.01919624,
  7.957171e-07, -1.296049e-05, 0.002035298, 9.533433e-07, 0.007283609, 
    0.000940282, 0.0005768876, -0.0001397751, 0.009101826, 0.005101627, 
    0.003802598, 0.00652031, 0.000324515, 0.04176914, 0.05507118, 0.06012256, 
    0.03215412, 0.02538635, 0.01968417, 0.008845164, 7.751206e-05, 
    -6.377072e-07, 8.7704e-08, 0.001434769, 0.0004254431, 0.0004400873, 
    0.006720566, 0.01671194, 0.004303857,
  2.738796e-06, 7.678154e-07, 3.977864e-06, 0.0004964995, 0.04622579, 
    0.02246014, 0.02341163, 0.02233234, 0.05802641, 0.02083725, 0.01832563, 
    0.01823488, 0.08655149, 0.05717077, 0.05186858, 0.0624903, 0.02840983, 
    0.0003473721, 4.769269e-05, 3.847231e-07, 3.058704e-09, 6.519398e-08, 
    0.004620228, -5.960985e-05, 2.436278e-06, 0.0004210147, 4.396349e-06, 
    0.000342035, 2.326848e-06,
  0.007037901, 0.0621459, 0.03177296, 0.002118937, 0.0009969862, 0.02403811, 
    0.03874115, 0.04648376, 0.08380426, 0.1275271, 0.02102054, 0.05098366, 
    0.1565828, 0.05145445, 0.05954864, 0.007323614, 0.03028632, 0.01197419, 
    2.420397e-05, 8.796212e-06, 3.838428e-06, 0.002427938, 0.0364931, 
    0.1210598, 0.0510917, 0.04589312, 0.02637707, 0.01585517, 0.002299894,
  0.08338294, 0.08577474, 0.09406229, -3.554554e-05, 0.009742448, 0.02609443, 
    0.09210517, 0.036126, 0.1524587, 0.09664975, 0.08019214, 0.116606, 
    0.1439222, 0.08262402, 0.06576984, 0.04492753, 0.06902227, 0.009211304, 
    0.03931, 0.01456938, 0.06177368, 0.1321443, 0.1548305, 0.04830026, 
    0.04409183, 0.01583739, 0.02866997, 0.14186, 0.1044168,
  0.06438324, 0.01408046, 0.001742265, 0.0001840429, 0.00601637, 0.06675531, 
    0.1007421, 0.1461087, 0.09597618, 0.09935302, 0.09732057, 0.09172412, 
    0.04300156, 0.01519504, 0.01857063, 0.01199307, 0.005841919, 0.004291579, 
    0.03215714, -5.257674e-05, 0.005240863, 0.04936855, 0.08137299, 
    0.1095699, 0.02997789, 0.00433265, 0.001206101, 0.02138515, 0.03836651,
  0.02652375, 0.06456235, 0.007517634, 0.004169717, -0.0001562291, 
    0.004509964, 0.02123318, 0.06437238, 0.2525602, 0.09638095, 0.2135553, 
    0.1728045, 0.1056902, 0.1001306, 0.09559642, 0.07406478, 0.06052219, 
    0.02572747, 0.01523575, 0.006541084, 0.01050363, 0.03654315, 0.0350436, 
    0.07496486, 0.1293098, 0.05880914, 0.002620434, 0.01415633, 0.008008374,
  0.08329631, 0.1045106, 0.03696825, 0.05276953, 0.06235651, 0.04913459, 
    0.1201189, 0.1673277, 0.1774157, 0.1210893, 0.1633446, 0.1452606, 
    0.2273964, 0.1787703, 0.1272057, 0.1976428, 0.186839, 0.09531356, 
    0.03842338, 0.05346416, 0.07923493, 0.07840244, 0.0587841, 0.06177794, 
    0.09738107, 0.1224485, 0.07807542, 0.05492472, 0.0587846,
  0.08988255, 0.1363014, 0.1135767, 0.06992521, 0.1091339, 0.08378896, 
    0.09224831, 0.1214961, 0.187089, 0.1950634, 0.1676157, 0.2260877, 
    0.1279725, 0.1241164, 0.1379029, 0.2103958, 0.2224934, 0.2028378, 
    0.1237837, 0.08354822, 0.1624123, 0.07216437, 0.08369119, 0.09299088, 
    0.1420825, 0.1844791, 0.1663857, 0.1371612, 0.1373498,
  0.1768979, 0.09234378, 0.1037795, 0.1023999, 0.1073681, 0.122866, 
    0.1360978, 0.1300298, 0.139397, 0.119525, 0.1773774, 0.2118973, 
    0.1490592, 0.1698877, 0.1302095, 0.1734956, 0.1612148, 0.1957811, 
    0.1416146, 0.1135229, 0.09684706, 0.1285939, 0.1316773, 0.1537178, 
    0.1921252, 0.1583727, 0.1502378, 0.2033554, 0.1654029,
  0.2033343, 0.1782511, 0.1645972, 0.103211, 0.154632, 0.2032724, 0.1234465, 
    0.1060687, 0.1414789, 0.1158943, 0.1090167, 0.09926471, 0.1004145, 
    0.05816668, 0.1129029, 0.1630025, 0.1410594, 0.1670236, 0.167058, 
    0.1955196, 0.1659611, 0.1481184, 0.1294612, 0.04864677, 0.1358811, 
    0.03134567, 0.001944995, 0.1544872, 0.1701181,
  0.1280032, 0.1413112, 0.1141867, 0.07235768, 0.09374116, 0.1693863, 
    0.1886399, 0.1885555, 0.1758854, 0.1465925, 0.1785018, 0.1764134, 
    0.1587035, 0.11319, 0.1423301, 0.1211591, 0.07644, 0.04926666, 
    0.08618713, 0.08715498, 0.06629759, 0.06978844, 0.06990661, 0.05397977, 
    0.07092354, 0.008864474, 0.01110062, 0.03711724, 0.1318926,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.948085e-07, 0.0003344404, 
    0.0001089079, 0.002761609, 0.003812298, 0.0001363745, 3.640494e-06, 
    -8.915282e-07, 0, 3.674492e-05, 7.460485e-05, 4.068484e-05, 0, 0, 0, 0,
  0.01685115, 0.01946981, 0.01771565, 0.005055591, -0.0002970931, 
    -0.001514658, 0.03204903, -7.07267e-05, -0.0003567371, -0.0005735426, 
    4.30668e-05, 0.0001046711, -0.0004826578, 0.03145483, 0.0428934, 
    0.03978264, 0.03452581, 0.03550456, 0.04586878, 0.08663465, 0.04736537, 
    0.05699155, 0.06079917, 0.04288556, 0.06152175, 0.02516407, 0.03999266, 
    0.02202721, 0.01732875,
  0.1118987, 0.1049279, 0.1185655, 0.1108751, 0.09922337, 0.1003952, 
    0.137832, 0.1236462, 0.1486658, 0.1298298, 0.1308676, 0.1646046, 
    0.1311831, 0.1879242, 0.1947589, 0.1510752, 0.1633087, 0.1310056, 
    0.1746552, 0.1890031, 0.185882, 0.1583851, 0.1750006, 0.121086, 
    0.1513451, 0.09765001, 0.0928743, 0.1126285, 0.1155416,
  0.1660806, 0.1423416, 0.1680363, 0.1617154, 0.1432296, 0.1648576, 
    0.1453382, 0.152598, 0.1368462, 0.1799435, 0.1559648, 0.2002799, 
    0.1963551, 0.2573825, 0.2624287, 0.1863809, 0.204089, 0.1976513, 
    0.2194836, 0.2161661, 0.2186724, 0.1755771, 0.1475175, 0.1108468, 
    0.13209, 0.1622529, 0.1971613, 0.2206969, 0.1368741,
  0.1278007, 0.08672077, 0.1028515, 0.126732, 0.1229383, 0.09967302, 
    0.08515367, 0.09785879, 0.1194775, 0.07590386, 0.09719927, 0.1232758, 
    0.127751, 0.1722634, 0.1434366, 0.1464016, 0.1474499, 0.1563434, 
    0.1435884, 0.1468418, 0.1364663, 0.20738, 0.1631419, 0.1679885, 
    0.09472926, 0.1316354, 0.1355825, 0.1232233, 0.1252215,
  0.03124187, 0.004094027, 0.02762324, 0.02783112, 0.008831222, 0.008498766, 
    0.0007684534, 0.005884079, 0.02540573, 0.01853101, 0.05237034, 0.0670779, 
    0.03417788, 0.04694984, 0.08491617, 0.1422691, 0.09287453, 0.124933, 
    0.1813056, 0.1754538, 0.02420896, 0.02405743, 0.02196079, 0.02738974, 
    0.03636663, 0.0506836, 0.05324464, 0.03181626, 0.02420234,
  9.051153e-08, 6.229943e-07, 0.0006681934, 1.425999e-05, 0.006392373, 
    0.01912325, 0.004779208, 0.00254662, 0.005509012, 0.001844654, 
    0.002270425, 0.005616322, 0.001927748, 0.04336708, 0.05997828, 
    0.05103143, 0.02151419, 0.01831817, 0.01743898, 0.01631968, 3.130047e-05, 
    -7.251487e-07, 3.924526e-08, 0.004440411, 0.0004063422, 2.284817e-05, 
    0.004944918, 0.009551033, 0.001304295,
  1.616582e-05, 4.167477e-06, 3.498844e-06, 0.003201101, 0.05228287, 
    0.02022043, 0.02341399, 0.0221555, 0.0583556, 0.02224882, 0.01525979, 
    0.02283467, 0.08882116, 0.05151983, 0.05731969, 0.0575272, 0.02226273, 
    0.000868974, 0.001307373, 7.636912e-09, -1.065546e-08, 7.262071e-08, 
    0.006298341, 0.0001331065, -1.618305e-07, 1.374961e-05, 0.0007438347, 
    -6.177254e-05, 1.029513e-06,
  0.007172228, 0.04471869, 0.03015316, 0.004700452, 0.001301347, 0.02315019, 
    0.0232465, 0.04505728, 0.05210415, 0.0776482, 0.01897906, 0.0375182, 
    0.1365106, 0.05185982, 0.04589648, 0.007053433, 0.03282871, 0.01312277, 
    1.926267e-05, 0.000378938, 1.580968e-06, 0.0001525346, 0.03115414, 
    0.1129547, 0.05484845, 0.06355492, 0.04423526, 0.01248525, 0.003697535,
  0.05662934, 0.07371691, 0.0910636, -2.021878e-05, 0.00520353, 0.02048613, 
    0.07414036, 0.02069028, 0.103746, 0.07718156, 0.0698004, 0.1022613, 
    0.1319449, 0.06813731, 0.06008727, 0.03677, 0.06977602, 0.005355314, 
    0.0419616, 0.01475547, 0.06641234, 0.1216474, 0.1241385, 0.03879807, 
    0.04506097, 0.01763132, 0.03801713, 0.1402822, 0.0800743,
  0.03649167, 0.01262533, 0.0003669278, 6.432092e-05, 0.001763577, 
    0.07080119, 0.08519213, 0.1170136, 0.07444105, 0.1000332, 0.1006749, 
    0.08359291, 0.03243827, 0.01116488, 0.01687105, 0.01718866, 0.003276282, 
    0.002329286, 0.01661073, 5.238676e-07, 0.002832817, 0.04608449, 
    0.0608708, 0.08525403, 0.01617376, 0.001400116, 0.004012994, 0.02639141, 
    0.03110324,
  0.0200434, 0.06613552, 0.007979695, 0.005366046, -2.68972e-05, 0.003081244, 
    0.01768168, 0.06327773, 0.2579399, 0.09184624, 0.2003147, 0.1579432, 
    0.09717721, 0.07812852, 0.08100417, 0.06624778, 0.06173972, 0.01801019, 
    0.006556363, 0.003734799, 0.002088619, 0.02179418, 0.0294846, 0.04690545, 
    0.1144389, 0.03914241, 0.001406986, 0.009730551, 0.009942412,
  0.07486952, 0.1005872, 0.02824198, 0.04595242, 0.06376317, 0.04815407, 
    0.168252, 0.1352294, 0.1518565, 0.1073289, 0.1569155, 0.127256, 0.207934, 
    0.1683631, 0.1171544, 0.1800173, 0.1832266, 0.07930902, 0.02941229, 
    0.05465717, 0.0646479, 0.0812903, 0.05033021, 0.05518976, 0.09095209, 
    0.1102625, 0.05531214, 0.05111105, 0.03556844,
  0.09425761, 0.1220527, 0.1007533, 0.06676342, 0.08472264, 0.07339583, 
    0.08676416, 0.1095407, 0.1871028, 0.1831984, 0.1631967, 0.2145488, 
    0.1153421, 0.1111301, 0.1175176, 0.2052758, 0.2230799, 0.2081194, 
    0.1209493, 0.07782622, 0.1548969, 0.06602059, 0.08292335, 0.09354337, 
    0.1342475, 0.1779262, 0.1635132, 0.1274309, 0.1431141,
  0.147933, 0.07965653, 0.09281068, 0.09400129, 0.09814654, 0.142397, 
    0.1331902, 0.1386137, 0.1746083, 0.1296413, 0.1637046, 0.2132125, 
    0.150508, 0.1544437, 0.1178247, 0.1683534, 0.1944436, 0.2083132, 
    0.1292566, 0.1178908, 0.08836883, 0.1191101, 0.1292151, 0.1821092, 
    0.1983803, 0.1911436, 0.146004, 0.2148646, 0.1672043,
  0.199905, 0.161668, 0.1661327, 0.09887616, 0.147442, 0.2122298, 0.1355787, 
    0.1177663, 0.137021, 0.1130328, 0.1212061, 0.09620051, 0.108826, 
    0.06218082, 0.1212082, 0.1527823, 0.1457634, 0.1924111, 0.1647905, 
    0.1909177, 0.181755, 0.1486441, 0.1264181, 0.08487037, 0.136241, 
    0.07873017, 0.01453838, 0.1729529, 0.1854952,
  0.1484333, 0.186916, 0.1363027, 0.1204547, 0.1482347, 0.2335933, 0.2328289, 
    0.2260816, 0.18954, 0.1648985, 0.1830395, 0.1935308, 0.206938, 0.1772783, 
    0.2242841, 0.1968053, 0.1351957, 0.09699643, 0.1280043, 0.1184682, 
    0.09955864, 0.115648, 0.08722843, 0.04557999, 0.1018046, 0.040835, 
    0.03906737, 0.07235324, 0.1529058,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001722708, 0.005760387, 
    0.007406279, 0.0126069, 0.005368571, 0.004361722, 0.0006543408, 
    0.0007824122, 1.633018e-06, 0.001879409, 0.03896289, 0.03860477, 
    0.007675647, 0.01399477, 0.002798518, 0,
  0.04218625, 0.04962423, 0.05308948, 0.02348199, 0.0008514166, 0.008070635, 
    0.05862632, 0.002607028, 0.000685835, 0.00112198, 0.002420834, 
    0.0004221615, 0.01851545, 0.1203598, 0.1730654, 0.1277109, 0.130914, 
    0.104016, 0.1377273, 0.157825, 0.1097547, 0.11523, 0.1171081, 0.102553, 
    0.1398565, 0.09085002, 0.1293396, 0.1531709, 0.07673392,
  0.1637736, 0.1699139, 0.184202, 0.1553054, 0.1552388, 0.1455417, 0.1510792, 
    0.1561182, 0.1981937, 0.2076885, 0.2143623, 0.2400422, 0.2294399, 
    0.2302658, 0.26881, 0.2225031, 0.2029782, 0.1692551, 0.2058221, 
    0.2464521, 0.2300843, 0.1900192, 0.2444118, 0.1765404, 0.2244107, 
    0.1553381, 0.1301502, 0.1589527, 0.163677,
  0.1816983, 0.1630774, 0.1830028, 0.154125, 0.1536802, 0.1626861, 0.1582419, 
    0.1593131, 0.1603615, 0.1874139, 0.1742321, 0.2021324, 0.1993075, 
    0.2489596, 0.2245073, 0.1527702, 0.2231967, 0.2072679, 0.2138883, 
    0.2229454, 0.2379851, 0.1795608, 0.1670582, 0.134321, 0.1291527, 
    0.1836607, 0.2187466, 0.2287477, 0.155763,
  0.1079681, 0.07762811, 0.09186879, 0.1152221, 0.1179853, 0.09057213, 
    0.09022921, 0.1054985, 0.1196643, 0.08733141, 0.1065343, 0.1153063, 
    0.1151965, 0.1611343, 0.1393605, 0.1464079, 0.1333936, 0.1479876, 
    0.1566691, 0.1547281, 0.1208496, 0.1936919, 0.168649, 0.1759783, 
    0.07822862, 0.1203249, 0.1266784, 0.1163787, 0.104994,
  0.03872447, 0.00233988, 0.02504887, 0.0275499, 0.009447903, 0.01123378, 
    0.003993235, 0.01098181, 0.02868806, 0.01223749, 0.04447192, 0.07211922, 
    0.03418873, 0.05285577, 0.06558256, 0.1353186, 0.08201151, 0.1218273, 
    0.1649874, 0.1591453, 0.02443155, 0.02272258, 0.02139498, 0.01881921, 
    0.03013691, 0.05233027, 0.04541761, 0.03265169, 0.03270039,
  -6.00906e-07, -1.134723e-06, 0.0004911856, 0.000118183, 0.006124334, 
    0.02344608, 0.006226411, 0.001192856, 0.006540957, 0.000747951, 
    0.001912573, 0.001625621, -5.402271e-05, 0.04267326, 0.06101528, 
    0.04955578, 0.016762, 0.01870447, 0.01878065, 0.01828565, 1.106257e-05, 
    1.504148e-07, 3.493553e-09, 0.006971348, 0.0003850514, 1.340912e-05, 
    0.00202147, 0.0002802304, 3.544096e-05,
  3.279261e-05, 9.011114e-06, 2.447244e-06, 0.004518205, 0.05345491, 
    0.02857473, 0.0234473, 0.01958153, 0.05496681, 0.02020936, 0.02986297, 
    0.01601389, 0.09514101, 0.05101236, 0.05738198, 0.05199368, 0.03011536, 
    0.002288393, 0.0001948548, 2.16375e-08, -4.772589e-09, 2.003014e-07, 
    0.0035424, 0.001376977, 4.124176e-05, 3.213157e-05, 0.003136716, 
    -4.121702e-07, 4.956074e-07,
  0.001807556, 0.04145161, 0.02908352, 0.006438105, 0.003240815, 0.02236678, 
    0.02157782, 0.04665248, 0.03704147, 0.04922997, 0.02463935, 0.04060635, 
    0.1328349, 0.04792269, 0.041256, 0.008107865, 0.03316122, 0.01000575, 
    0.0006387245, 0.00594581, 3.442901e-05, 0.0003364905, 0.02668461, 
    0.1169125, 0.06866375, 0.08132301, 0.06684332, 0.02341953, 0.004786497,
  0.03724613, 0.0601318, 0.08544453, 0.0001597469, 0.001470415, 0.01976682, 
    0.06907484, 0.01841685, 0.07181666, 0.06342614, 0.06042433, 0.09317761, 
    0.1195378, 0.06711899, 0.06126566, 0.03686773, 0.0765873, 0.01042497, 
    0.05612619, 0.01828253, 0.07004086, 0.115845, 0.1047381, 0.03493191, 
    0.04722991, 0.01762303, 0.03090069, 0.134236, 0.06033789,
  0.04004138, 0.01436116, -7.253363e-05, 0.0009431404, 0.001767125, 
    0.0631118, 0.08641551, 0.0886239, 0.07888144, 0.1047532, 0.09095193, 
    0.07393301, 0.02512856, 0.008869041, 0.01522484, 0.01526183, 0.001854085, 
    0.000670129, 0.003357302, 0.0002806, 0.001736698, 0.04413443, 0.04678056, 
    0.06627549, 0.009573752, 0.006582462, 0.02277117, 0.02065285, 0.02920792,
  0.01380825, 0.07010613, 0.01012514, 0.01108082, -2.333647e-05, 0.002974759, 
    0.02475362, 0.0743178, 0.2629125, 0.08563372, 0.1979234, 0.1466976, 
    0.1015392, 0.06501542, 0.07773753, 0.05472061, 0.06105055, 0.01733242, 
    0.006453975, 0.001498684, 0.00123939, 0.01658335, 0.02971794, 0.03341214, 
    0.107946, 0.03024738, 0.0001511061, 0.0005092978, 0.01136359,
  0.06503284, 0.09940659, 0.0248171, 0.04834014, 0.06645069, 0.03318161, 
    0.1680605, 0.1056547, 0.1243343, 0.1102439, 0.1449785, 0.1095209, 
    0.1858075, 0.1625338, 0.1036931, 0.1810436, 0.1721127, 0.06352083, 
    0.02298672, 0.04481966, 0.056247, 0.07678846, 0.04617919, 0.04450434, 
    0.09005812, 0.107891, 0.06014618, 0.05095377, 0.02833192,
  0.09605582, 0.1122131, 0.09502207, 0.06210245, 0.07088356, 0.06412116, 
    0.08293944, 0.09892616, 0.1858363, 0.1686156, 0.1617057, 0.2058144, 
    0.1034732, 0.1071725, 0.1078816, 0.1984202, 0.2133104, 0.2104487, 
    0.129862, 0.07235975, 0.1534758, 0.06627934, 0.08608477, 0.08823857, 
    0.1294559, 0.1840689, 0.1584699, 0.1377544, 0.1450938,
  0.1352866, 0.06951799, 0.08377272, 0.08960681, 0.09874289, 0.1433541, 
    0.123658, 0.1285437, 0.1755833, 0.1251347, 0.1512858, 0.1991403, 
    0.1492749, 0.1448098, 0.1071578, 0.1642393, 0.1903353, 0.2109461, 
    0.1233653, 0.1029855, 0.07464246, 0.1062731, 0.1288614, 0.1918468, 
    0.1894324, 0.2169674, 0.1500048, 0.2216549, 0.16496,
  0.1879192, 0.1475169, 0.161315, 0.08368637, 0.1412759, 0.2086756, 
    0.1357923, 0.1291923, 0.1214632, 0.1117716, 0.1215053, 0.1057366, 
    0.1078284, 0.05343845, 0.114421, 0.132839, 0.1332262, 0.1722816, 
    0.1565612, 0.1777437, 0.1771039, 0.1402439, 0.1336136, 0.09698159, 
    0.1152388, 0.1801797, 0.05889672, 0.1616871, 0.2031296,
  0.1384604, 0.1691241, 0.1251727, 0.1347881, 0.1641884, 0.2450962, 
    0.2258933, 0.2207799, 0.1856966, 0.1529962, 0.1544029, 0.1789974, 
    0.2018682, 0.1945595, 0.2448136, 0.2109714, 0.1433628, 0.1044101, 
    0.1484348, 0.1505489, 0.1472847, 0.1620148, 0.1420251, 0.08706575, 
    0.1233196, 0.05891674, 0.07753901, 0.07975227, 0.1459952,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.358788e-05, 0.01417667, 0.0552721, 
    0.04756778, 0.05290637, 0.02868539, 0.01039821, 0.002386144, 0.002316389, 
    0.0007912758, 0.01283687, 0.1833582, 0.1272644, 0.06165918, 0.04944117, 
    0.003504156, 0,
  0.09561408, 0.1545134, 0.139877, 0.08875389, 0.005637394, 0.0240904, 
    0.09920998, 0.02300475, 0.003287934, 0.008061749, 0.01693068, 
    0.007601053, 0.07342906, 0.2063983, 0.1964873, 0.1558133, 0.1726864, 
    0.1871389, 0.1794132, 0.1951349, 0.1775938, 0.2051415, 0.1743664, 
    0.1722241, 0.237315, 0.1671455, 0.2273321, 0.2116857, 0.1503443,
  0.1864105, 0.2042574, 0.2469907, 0.2047035, 0.222477, 0.1928379, 0.1793417, 
    0.1855455, 0.2356453, 0.274217, 0.240816, 0.2851996, 0.2409573, 
    0.2269794, 0.2741715, 0.2312063, 0.2108364, 0.1855201, 0.211035, 
    0.2329277, 0.232549, 0.1983678, 0.2509934, 0.1983118, 0.2509349, 
    0.2100499, 0.198391, 0.1877559, 0.1967854,
  0.1901014, 0.1739551, 0.1909865, 0.149468, 0.14555, 0.158101, 0.1609835, 
    0.1742137, 0.1782238, 0.1923052, 0.1863803, 0.1955791, 0.1880774, 
    0.2339779, 0.2210168, 0.1352749, 0.2140794, 0.213772, 0.2167445, 
    0.2056178, 0.2089634, 0.1864465, 0.1668411, 0.1397035, 0.1345917, 
    0.1814662, 0.2314456, 0.2334711, 0.1750996,
  0.09406412, 0.08065011, 0.07677637, 0.1081592, 0.1164508, 0.08369817, 
    0.08401343, 0.09412564, 0.1115684, 0.09371409, 0.1111739, 0.1088962, 
    0.1076995, 0.1557799, 0.134575, 0.1271188, 0.1416678, 0.1384838, 
    0.1526991, 0.1622256, 0.1181622, 0.1799056, 0.1659891, 0.190111, 
    0.07324798, 0.1187294, 0.1239636, 0.1051699, 0.09596786,
  0.03933605, 0.002133084, 0.02468214, 0.03247532, 0.01022615, 0.01380883, 
    0.008775651, 0.01294391, 0.03315991, 0.0151193, 0.03729645, 0.06516566, 
    0.03526326, 0.04837099, 0.05394323, 0.1252095, 0.08618265, 0.1107166, 
    0.1601262, 0.1647989, 0.02435218, 0.03167163, 0.0201456, 0.01672692, 
    0.02678426, 0.05109913, 0.03845398, 0.0322521, 0.03412197,
  5.391301e-05, 6.103052e-08, 0.0005375885, 8.647906e-05, 0.009402777, 
    0.02053528, 0.00320899, 0.0006553058, 0.007946742, 0.003238288, 
    0.005595911, 0.009401095, 0.001280124, 0.04415671, 0.06513596, 
    0.04632225, 0.01809585, 0.021248, 0.0155374, 0.02121441, 2.641847e-05, 
    -4.518847e-07, -3.898577e-10, 0.01701248, 0.0003581217, 8.204262e-06, 
    2.862479e-06, 0.0006884746, 0.002694933,
  9.98622e-06, 5.624103e-06, 1.499726e-05, 0.005118657, 0.04749185, 
    0.03740554, 0.02411046, 0.02112668, 0.05112503, 0.02219976, 0.04410102, 
    0.01266604, 0.09810975, 0.05204674, 0.0607008, 0.05773689, 0.04131819, 
    0.003796816, 0.000251445, 4.737194e-08, 4.913471e-09, 3.028042e-07, 
    0.0001929871, 0.001683911, 0.0001697294, 0.0006449078, 0.009374787, 
    -4.680535e-08, 2.394203e-07,
  0.002758763, 0.04437212, 0.02958883, 0.01205533, 0.003474845, 0.01799656, 
    0.02028824, 0.03562883, 0.03553129, 0.04019587, 0.02581985, 0.03668606, 
    0.1251474, 0.05498321, 0.0397962, 0.008564238, 0.03154062, 0.007486401, 
    0.002254894, 0.006750023, 0.002789211, 2.986818e-06, 0.03068849, 
    0.1241288, 0.09048441, 0.09080458, 0.0770195, 0.007978609, 0.005356606,
  0.02970057, 0.05375747, 0.07869399, 0.006618788, 0.001288975, 0.02156251, 
    0.05945064, 0.0273182, 0.05529268, 0.06494572, 0.05405223, 0.08741331, 
    0.1181616, 0.0689503, 0.05146104, 0.04581477, 0.08474462, 0.02613727, 
    0.07324233, 0.02528799, 0.06709506, 0.1139095, 0.09807345, 0.03630346, 
    0.04058861, 0.02266189, 0.03354523, 0.129818, 0.05718397,
  0.06992589, 0.02167803, -0.000191672, 0.0003631113, 0.0005172915, 
    0.05329903, 0.09578974, 0.08846092, 0.0779829, 0.1026985, 0.09699106, 
    0.06959331, 0.02358336, 0.006234071, 0.00965459, 0.01473324, 0.002708048, 
    7.383795e-06, 0.01037493, 0.01220982, 0.003249379, 0.0466007, 0.03789981, 
    0.05472516, 0.007676463, 0.01444557, 0.01828124, 0.0162484, 0.02480746,
  0.01334175, 0.07123172, 0.01142334, 0.01441792, -0.0002122599, 0.004659319, 
    0.01760905, 0.08133665, 0.2711155, 0.0774002, 0.199901, 0.1516556, 
    0.1048738, 0.05462617, 0.07614498, 0.04872743, 0.04988332, 0.01303687, 
    0.006996097, 0.0008227363, 0.003961448, 0.01903338, 0.02416288, 
    0.02955728, 0.09241137, 0.02807202, -0.0003331953, 6.341656e-06, 
    0.01482639,
  0.05786688, 0.09489688, 0.02277841, 0.04953187, 0.06257685, 0.02243169, 
    0.1633039, 0.08251394, 0.1004726, 0.1176362, 0.1404681, 0.09732296, 
    0.1686896, 0.1583438, 0.09791909, 0.182353, 0.1539151, 0.04408591, 
    0.02244284, 0.03691255, 0.06076416, 0.07323363, 0.04635892, 0.0406067, 
    0.09158593, 0.1050609, 0.0557007, 0.04451995, 0.01963644,
  0.09020372, 0.1019743, 0.09375741, 0.05796504, 0.06386244, 0.0592277, 
    0.08762019, 0.09952234, 0.1813073, 0.1632399, 0.1691211, 0.1910619, 
    0.09708823, 0.1107174, 0.1052978, 0.1969209, 0.2019905, 0.2023798, 
    0.1177906, 0.06811978, 0.1579776, 0.06692983, 0.07861929, 0.08645141, 
    0.1290328, 0.1947632, 0.1486921, 0.1254073, 0.1234301,
  0.1298524, 0.06406058, 0.07449745, 0.08597176, 0.09285326, 0.1523963, 
    0.1241861, 0.1164931, 0.1682343, 0.1317365, 0.1408846, 0.1795924, 
    0.1458983, 0.1266468, 0.09765776, 0.1638014, 0.2002514, 0.2245324, 
    0.1213812, 0.08998124, 0.06852446, 0.0917712, 0.1333277, 0.2098669, 
    0.180344, 0.243953, 0.15826, 0.2159995, 0.1624857,
  0.1852656, 0.1407475, 0.1581209, 0.08075748, 0.1373938, 0.2143348, 
    0.1397092, 0.1362527, 0.1102352, 0.1152169, 0.114128, 0.1021901, 
    0.1080724, 0.05588465, 0.1118564, 0.1143539, 0.1227445, 0.1607885, 
    0.1563915, 0.1714686, 0.1646844, 0.1352894, 0.1377424, 0.1131772, 
    0.1100425, 0.2840912, 0.1074009, 0.1595034, 0.2002535,
  0.132932, 0.1675085, 0.1341851, 0.1521674, 0.1675836, 0.2559909, 0.2468792, 
    0.2260388, 0.1807616, 0.1515575, 0.1481552, 0.1698677, 0.1838677, 
    0.1891162, 0.2434215, 0.2109644, 0.1452268, 0.1087991, 0.1480446, 
    0.1691615, 0.1591915, 0.1748189, 0.1708481, 0.1098591, 0.1215064, 
    0.08827736, 0.1088506, 0.08261315, 0.1439143,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005900447, 0.07914361, 0.08975123, 
    0.1105896, 0.1320651, 0.1060618, 0.04858137, 0.02468555, 0.006096557, 
    0.004481892, 0.06239768, 0.2725258, 0.2379109, 0.1725181, 0.1231346, 
    0.03598095, 9.969653e-05,
  0.1435688, 0.2323566, 0.251947, 0.1914632, 0.02145921, 0.06063207, 
    0.1524162, 0.05130417, 0.03385397, 0.03207766, 0.04313251, 0.03262303, 
    0.1478572, 0.2314337, 0.2166342, 0.1753111, 0.1745627, 0.2270225, 
    0.2191106, 0.2800964, 0.2588252, 0.2556108, 0.2041929, 0.2953309, 
    0.2999744, 0.2209544, 0.2628456, 0.2665052, 0.2192011,
  0.1966706, 0.2484947, 0.2662725, 0.2449152, 0.279334, 0.2503565, 0.2047735, 
    0.1986051, 0.2536618, 0.3285509, 0.2474934, 0.278346, 0.2253988, 
    0.218152, 0.2521947, 0.2425339, 0.2221291, 0.1851985, 0.2008392, 
    0.2097984, 0.2280136, 0.2266806, 0.2849891, 0.2181264, 0.2674207, 
    0.2556408, 0.2331525, 0.2106124, 0.2225088,
  0.1845995, 0.1632761, 0.1860233, 0.1511188, 0.1451158, 0.153246, 0.1606096, 
    0.1881758, 0.1809197, 0.2028915, 0.1912708, 0.1850405, 0.1856543, 
    0.2139139, 0.2156028, 0.1034255, 0.212125, 0.1936281, 0.2054363, 
    0.2031359, 0.2104954, 0.1896524, 0.1405692, 0.1328552, 0.1240213, 
    0.1873744, 0.2298735, 0.2394439, 0.172249,
  0.08084316, 0.08870965, 0.06911177, 0.1110526, 0.1167941, 0.08690552, 
    0.08841685, 0.104697, 0.1008241, 0.08681015, 0.1152804, 0.1104953, 
    0.1068877, 0.136775, 0.1284394, 0.114673, 0.1320784, 0.1431254, 
    0.1524647, 0.1595474, 0.1132371, 0.1517005, 0.1559433, 0.2013565, 
    0.06694264, 0.1104088, 0.1197534, 0.09006477, 0.09122285,
  0.045663, 0.003639275, 0.02160454, 0.03427158, 0.01478771, 0.014503, 
    0.01205824, 0.0185889, 0.02681731, 0.01501762, 0.02972017, 0.05718572, 
    0.02895681, 0.0422264, 0.05221145, 0.1240679, 0.07761815, 0.09904481, 
    0.1475979, 0.1761063, 0.0295711, 0.02926623, 0.01896813, 0.01982834, 
    0.02293602, 0.05317911, 0.03955118, 0.03924299, 0.04409464,
  1.922703e-07, 2.395502e-08, 0.0004372651, 5.12168e-05, 0.01949817, 
    0.02181721, 0.00331712, 0.001737111, 0.005031025, 0.003641545, 
    0.007474528, 0.001292297, 0.005674713, 0.04226604, 0.04601804, 
    0.04325534, 0.02570708, 0.023734, 0.01316806, 0.02365042, 0.0001749739, 
    -8.75991e-07, 2.04814e-09, 0.01849348, 0.0003197955, 6.818337e-06, 
    -0.0001219711, 0.0002051107, 0.004158498,
  6.161753e-06, -2.76864e-06, 1.786184e-05, 0.005982968, 0.04347312, 
    0.03645035, 0.02717916, 0.03030619, 0.04259561, 0.01833362, 0.04949495, 
    0.01618992, 0.1059471, 0.05362644, 0.0631392, 0.06787399, 0.04728355, 
    0.002278047, 0.000282758, -5.159408e-07, 4.819255e-08, 7.510451e-07, 
    4.216665e-06, 0.0006604559, 0.0001650937, 2.067822e-05, 0.001395122, 
    1.182806e-07, 2.910964e-07,
  0.0270045, 0.04083231, 0.03037202, 0.01766724, 0.004108141, 0.0119182, 
    0.02486321, 0.03643516, 0.03460391, 0.03813378, 0.02953096, 0.04169562, 
    0.1298185, 0.0761025, 0.0367869, 0.01379311, 0.02848753, 0.005317911, 
    0.01196676, 0.01491405, 0.02433193, 0.0001552613, 0.03507484, 0.1326008, 
    0.09955405, 0.08149142, 0.0809281, 0.01013028, 0.003820488,
  0.02872885, 0.03811308, 0.04995688, 0.08173966, 0.002564398, 0.01051868, 
    0.06232492, 0.03604351, 0.05550309, 0.07642286, 0.06053739, 0.08988405, 
    0.1163585, 0.08064167, 0.05499098, 0.05348631, 0.07793905, 0.03263292, 
    0.09001531, 0.03099482, 0.07563513, 0.1206285, 0.09945714, 0.04453315, 
    0.04523263, 0.02639266, 0.04306106, 0.1260298, 0.05812595,
  0.08916333, 0.02506957, 0.0002434685, -3.078601e-05, 0.0004888849, 
    0.04426003, 0.1135561, 0.1316199, 0.09602173, 0.118336, 0.109055, 
    0.07525818, 0.02639633, 0.005140139, 0.007458893, 0.01138123, 
    0.002258742, 1.74012e-05, 0.01439845, 0.001929738, 0.005840757, 
    0.05227533, 0.03360102, 0.05198452, 0.007169801, 0.01408597, 0.01640304, 
    0.01639805, 0.02274788,
  0.009908276, 0.05380156, 0.003501372, 0.007907783, 0.002440242, 
    0.001638262, 0.01714274, 0.07933066, 0.2703767, 0.07123126, 0.1978595, 
    0.1599835, 0.1023327, 0.04789796, 0.08099927, 0.04723791, 0.04016789, 
    0.01081382, 0.00273938, 0.000280719, 0.005957784, 0.01398281, 0.02097334, 
    0.02384825, 0.08491026, 0.02671324, -0.0001483273, 9.620153e-06, 
    0.01151215,
  0.05297801, 0.08559796, 0.02318583, 0.05233881, 0.05767224, 0.02017507, 
    0.1646072, 0.06547582, 0.08078811, 0.1212691, 0.1377197, 0.08221814, 
    0.1563304, 0.148633, 0.09318393, 0.1761677, 0.1374165, 0.04751525, 
    0.02158677, 0.02992419, 0.07032908, 0.06037422, 0.05445432, 0.03741547, 
    0.08821292, 0.1002237, 0.05319101, 0.03221081, 0.01652579,
  0.08084758, 0.1085937, 0.102744, 0.05992267, 0.07051499, 0.06613477, 
    0.1021925, 0.09835194, 0.1782299, 0.1599929, 0.1617108, 0.1826693, 
    0.09131682, 0.1196955, 0.1124573, 0.1982037, 0.2211685, 0.1968006, 
    0.1236907, 0.07061215, 0.151416, 0.07256491, 0.07706235, 0.08316585, 
    0.1275488, 0.1825946, 0.1402972, 0.114316, 0.1133346,
  0.1385927, 0.07681172, 0.06829704, 0.08709101, 0.09042503, 0.1563892, 
    0.1311118, 0.1178578, 0.1665484, 0.1401772, 0.1320086, 0.1633214, 
    0.1492651, 0.1202777, 0.09338912, 0.1801693, 0.212503, 0.245125, 
    0.1313738, 0.08371495, 0.07102428, 0.0879574, 0.1521319, 0.2145856, 
    0.1730013, 0.25657, 0.1905697, 0.2279529, 0.160403,
  0.1837746, 0.1360109, 0.1634791, 0.07972956, 0.1401377, 0.2362434, 
    0.1610375, 0.1421344, 0.103468, 0.1264967, 0.1073915, 0.1130694, 
    0.1269092, 0.0724286, 0.116836, 0.09883323, 0.1153948, 0.1463728, 
    0.1599297, 0.161871, 0.1691527, 0.1376119, 0.1396682, 0.1294855, 
    0.09530658, 0.3176176, 0.2553545, 0.1606666, 0.1937539,
  0.136529, 0.1852838, 0.1529761, 0.1575304, 0.1630919, 0.2616325, 0.2352436, 
    0.2048085, 0.1775841, 0.1494713, 0.1643028, 0.1743733, 0.1777119, 
    0.1925443, 0.2473541, 0.2039261, 0.1488148, 0.1084912, 0.1433517, 
    0.1772899, 0.173356, 0.1818165, 0.1841452, 0.1160661, 0.1208388, 
    0.1119092, 0.1135246, 0.08820374, 0.163472,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001038164, -9.522424e-05, 
    -8.663206e-05, -7.803989e-05, -6.944771e-05, -6.085554e-05, 
    -5.226337e-05, 2.878378e-05, 2.019161e-05, 1.159944e-05, 3.007261e-06, 
    -5.584914e-06, -1.417709e-05, -2.276926e-05, 0,
  6.024103e-05, -1.834097e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.214482e-05, 
    0.001115164, 0.1365593, 0.1651776, 0.1919234, 0.1669611, 0.1638435, 
    0.1303946, 0.05600888, 0.02435666, 0.0226381, 0.1354666, 0.3330185, 
    0.3217731, 0.2259566, 0.2130984, 0.06013103, 0.001474798,
  0.1529079, 0.2781278, 0.2643954, 0.2726429, 0.04245873, 0.1161307, 
    0.2187285, 0.09720863, 0.0793547, 0.07422113, 0.09024781, 0.1056615, 
    0.1827848, 0.2278676, 0.2054275, 0.1951305, 0.1995413, 0.2506287, 
    0.2355845, 0.2889914, 0.302036, 0.3103786, 0.2628626, 0.3329265, 
    0.3148519, 0.2234155, 0.2519036, 0.3020672, 0.2583914,
  0.1971812, 0.2793487, 0.276308, 0.2515375, 0.3051436, 0.2643588, 0.2178466, 
    0.2114592, 0.260377, 0.3387677, 0.2504198, 0.2615659, 0.2343897, 
    0.2195043, 0.2328147, 0.2266857, 0.2190564, 0.1954959, 0.2214745, 
    0.2165479, 0.2277572, 0.2490308, 0.2847259, 0.2347762, 0.2639967, 
    0.2573938, 0.2386308, 0.2215782, 0.2181424,
  0.1819565, 0.1555217, 0.1804525, 0.1485121, 0.1499702, 0.1522302, 
    0.1588451, 0.197695, 0.1853883, 0.1985564, 0.1834572, 0.1824607, 
    0.1712311, 0.2046902, 0.2168217, 0.1292379, 0.212307, 0.1777556, 
    0.2044913, 0.2070943, 0.1940093, 0.1910905, 0.1389763, 0.1249584, 
    0.11801, 0.1661845, 0.214163, 0.2297682, 0.1729381,
  0.0739824, 0.09912644, 0.07997297, 0.1211827, 0.1276229, 0.09005825, 
    0.08713789, 0.1015698, 0.113664, 0.09111414, 0.1282643, 0.1075042, 
    0.1053526, 0.1314312, 0.1345757, 0.1058837, 0.1245515, 0.1479761, 
    0.1466388, 0.1441828, 0.1054335, 0.1419606, 0.1562657, 0.2134594, 
    0.06550785, 0.09731936, 0.1119125, 0.08837893, 0.1011007,
  0.03814028, 0.005554047, 0.02164408, 0.04057847, 0.02323358, 0.01582592, 
    0.01502217, 0.02005343, 0.03233248, 0.01702687, 0.02355536, 0.05243375, 
    0.03066659, 0.04006431, 0.05172516, 0.1307373, 0.06311461, 0.08721583, 
    0.1371553, 0.1902246, 0.0358352, 0.03095606, 0.01907101, 0.01860355, 
    0.01982409, 0.06513487, 0.03934488, 0.03728876, 0.04536297,
  9.303165e-08, 2.604936e-08, 0.0004647024, 0.0001078242, 0.02879983, 
    0.02627917, 0.001720164, 0.005414894, 0.003329738, 0.002522034, 
    0.008656939, -4.948741e-05, 0.008475519, 0.04975473, 0.03887663, 
    0.03697748, 0.03178342, 0.03021253, 0.01177054, 0.02615243, 0.0007263968, 
    -2.2856e-05, 4.429929e-08, 0.01409269, 0.0003985242, 9.477915e-06, 
    0.0002001356, 0.0004291877, 0.006931406,
  2.903654e-06, 2.368607e-05, 1.613845e-06, 0.01210019, 0.05098293, 
    0.03655143, 0.03252139, 0.03508037, 0.04555815, 0.01764905, 0.05514557, 
    0.02758414, 0.1177697, 0.0690048, 0.07001851, 0.07335512, 0.05874015, 
    0.005272286, 0.001142469, -1.674839e-06, 2.075498e-07, 1.144326e-06, 
    0.0002346522, 0.001286955, 0.0002415968, 1.306033e-05, 1.499834e-05, 
    5.495856e-07, 1.478071e-06,
  0.04407182, 0.05087601, 0.03707907, 0.01908592, 0.002298639, 0.01436931, 
    0.03558636, 0.03940652, 0.0424997, 0.04163143, 0.0545268, 0.05559144, 
    0.1548968, 0.09467545, 0.03861804, 0.01978026, 0.02788943, 0.007083197, 
    0.01140383, 0.01805833, 0.007242798, 0.001037536, 0.03733145, 0.155871, 
    0.1090485, 0.08382018, 0.08228265, 0.01409565, 0.006117197,
  0.0299615, 0.02331774, 0.0240168, 0.2580581, 0.002288363, 0.01391638, 
    0.06822893, 0.04090839, 0.08911971, 0.1058549, 0.0934242, 0.1087265, 
    0.1365227, 0.09145035, 0.06876749, 0.05994637, 0.07350498, 0.04576997, 
    0.09752132, 0.03821, 0.08284903, 0.1368577, 0.1167598, 0.05565438, 
    0.06063341, 0.04003024, 0.05653841, 0.1454321, 0.07402738,
  0.0421927, 0.01998132, 0.0001019905, -3.114977e-05, -1.529161e-05, 
    0.02599417, 0.1224008, 0.1636458, 0.1496638, 0.1437341, 0.1374875, 
    0.08392198, 0.03593713, 0.006306999, 0.01003668, 0.009255781, 
    0.002414911, 0.0002024049, 0.01550534, 0.0002120745, 0.006198796, 
    0.05993522, 0.04002659, 0.05512506, 0.007983564, 0.01503714, 0.02243766, 
    0.01996122, 0.02191726,
  0.003522573, 0.03874001, 0.003054834, 0.004102206, 0.0005325063, 
    9.06331e-05, 0.0148859, 0.09074216, 0.2653806, 0.06984462, 0.1988698, 
    0.1786856, 0.1055195, 0.04975054, 0.08733094, 0.05144875, 0.04116678, 
    0.01232682, 0.002570155, 9.03389e-05, 0.007363939, 0.01331132, 
    0.02471368, 0.02774341, 0.09051459, 0.02573609, 0.0002640077, 
    1.851614e-05, 0.004636895,
  0.05434339, 0.0747582, 0.02681232, 0.05552964, 0.04812161, 0.01487312, 
    0.1596884, 0.05445031, 0.0700651, 0.1113585, 0.137277, 0.07027168, 
    0.1459683, 0.1447503, 0.08784534, 0.1698394, 0.1313514, 0.04959564, 
    0.02721886, 0.02576436, 0.07070023, 0.05100834, 0.05140214, 0.04338065, 
    0.0877251, 0.1115389, 0.05181539, 0.03096927, 0.01949231,
  0.089543, 0.1100472, 0.1238615, 0.06420949, 0.07934694, 0.06514095, 
    0.1058798, 0.09704983, 0.174475, 0.1597041, 0.1684296, 0.1791284, 
    0.1034745, 0.1342951, 0.123653, 0.1950769, 0.1940277, 0.1788229, 
    0.1336437, 0.07788429, 0.1639469, 0.08444919, 0.08345918, 0.09169886, 
    0.1367383, 0.1739061, 0.1380353, 0.1137287, 0.1003837,
  0.1391273, 0.06548336, 0.07000852, 0.08566169, 0.09572634, 0.1743999, 
    0.1320364, 0.1219476, 0.1677458, 0.1456621, 0.1293687, 0.1601702, 
    0.1435914, 0.1158119, 0.1071705, 0.1888018, 0.2238274, 0.2592558, 
    0.119343, 0.08514781, 0.08619013, 0.08108007, 0.161906, 0.213866, 
    0.1966408, 0.2845098, 0.2101648, 0.2248198, 0.150505,
  0.1676506, 0.1201338, 0.1693185, 0.09701463, 0.1404094, 0.2343791, 
    0.1861529, 0.1341651, 0.09667358, 0.1378175, 0.1031917, 0.1335283, 
    0.122832, 0.1118376, 0.1123988, 0.09396229, 0.1055002, 0.1447432, 
    0.1640033, 0.1611792, 0.1709032, 0.1403027, 0.1561828, 0.1313399, 
    0.0716761, 0.3186438, 0.294462, 0.1645704, 0.2023464,
  0.1234392, 0.1871141, 0.1669874, 0.1808793, 0.1720871, 0.2531525, 
    0.2489707, 0.2245923, 0.200559, 0.1873835, 0.1597632, 0.1742647, 
    0.1864662, 0.2186003, 0.2689466, 0.2064243, 0.1561673, 0.1423308, 
    0.151212, 0.2070116, 0.1839774, 0.1990088, 0.2040047, 0.124049, 0.125984, 
    0.1101217, 0.1149092, 0.114387, 0.1479683,
  0, 0, 0, 0, 0, 0, 0, -7.604075e-05, -5.026422e-05, -2.44877e-05, 
    1.288826e-06, 2.706535e-05, 5.284188e-05, 7.86184e-05, -0.0003753903, 
    -0.0003667981, -0.000358206, -0.0003496138, -0.0003410216, -0.0003324294, 
    -0.0003238373, 0.0001151351, 8.076644e-05, 4.639774e-05, 1.202904e-05, 
    -2.233965e-05, -5.670835e-05, -9.107705e-05, 0,
  -0.000951823, 0.0002880678, -1.022431e-05, 0, 0, -1.707552e-06, 
    -9.76271e-06, 0, 0, 0, -0.0003347971, 0.0008382877, 0.005961027, 
    0.1815204, 0.1993517, 0.2061861, 0.2004479, 0.189143, 0.1905208, 
    0.1525397, 0.07523263, 0.07771572, 0.197061, 0.3395751, 0.3199232, 
    0.2504911, 0.2764216, 0.134265, 0.02132137,
  0.1486197, 0.2770699, 0.2690283, 0.3013566, 0.0822515, 0.1652577, 
    0.2763813, 0.1634509, 0.126987, 0.1354407, 0.1288459, 0.1495516, 
    0.2098434, 0.2427509, 0.2096416, 0.1856397, 0.1935865, 0.2550701, 
    0.2786321, 0.3190219, 0.2958433, 0.327699, 0.2634373, 0.3454728, 
    0.3134388, 0.2104636, 0.23438, 0.2892735, 0.2519397,
  0.2187125, 0.2910094, 0.286402, 0.2676567, 0.3002118, 0.270364, 0.2237219, 
    0.2042123, 0.2637169, 0.358407, 0.2588623, 0.2710584, 0.2204698, 
    0.2023136, 0.2263543, 0.2169608, 0.2156579, 0.2039471, 0.2177805, 
    0.2055682, 0.2357991, 0.2192381, 0.2833074, 0.2409369, 0.2689124, 
    0.2402006, 0.2237548, 0.1992033, 0.2071254,
  0.1890578, 0.1567839, 0.1844741, 0.1431655, 0.1546633, 0.1458955, 
    0.1588894, 0.1992962, 0.1771341, 0.1841934, 0.1991673, 0.1905524, 
    0.170929, 0.1985092, 0.1954822, 0.1374251, 0.2159986, 0.1701726, 
    0.1954394, 0.1813667, 0.1939886, 0.1955473, 0.1461002, 0.1207019, 
    0.1202486, 0.1588911, 0.1950758, 0.210014, 0.1802895,
  0.06852502, 0.1112175, 0.08547297, 0.1316887, 0.1373561, 0.09756084, 
    0.08756395, 0.1024357, 0.1166188, 0.1018374, 0.1508695, 0.1254461, 
    0.09986117, 0.1363586, 0.142517, 0.1039739, 0.1253791, 0.1264258, 
    0.1428456, 0.1289956, 0.1025425, 0.1387456, 0.1579576, 0.2163499, 
    0.06479413, 0.09627329, 0.1166136, 0.08549614, 0.08938104,
  0.04212712, 0.004788905, 0.0261616, 0.0521134, 0.03145016, 0.02267637, 
    0.01766069, 0.02702864, 0.03489015, 0.01582031, 0.02226857, 0.03987977, 
    0.02783635, 0.04452346, 0.05416943, 0.1347408, 0.0677295, 0.08330001, 
    0.129211, 0.2021692, 0.05243476, 0.03266502, 0.02293492, 0.01272043, 
    0.02617595, 0.07989898, 0.05072208, 0.04225914, 0.03771874,
  1.071407e-07, 5.208752e-08, 0.0006078638, -1.734508e-05, 0.04610048, 
    0.02969018, 0.004637894, 0.02838887, 0.002193865, 0.003891818, 
    0.01193975, 0.0005062523, 0.012252, 0.06353664, 0.04083655, 0.03751141, 
    0.03378254, 0.04021556, 0.01672489, 0.02445716, 0.007923704, 
    -3.467012e-05, 6.734511e-08, 0.002049345, 0.002274775, 3.419191e-05, 
    0.001190256, 0.0005176236, 0.009283578,
  3.101174e-06, 7.047965e-05, 5.160408e-06, 0.01349581, 0.0584207, 0.0437924, 
    0.02894164, 0.03811187, 0.05765057, 0.02496266, 0.05225721, 0.02783306, 
    0.1299059, 0.08465865, 0.07391827, 0.08308018, 0.06738383, 0.00542672, 
    0.001784874, 1.444293e-07, -5.349705e-09, 6.337041e-07, 0.0003655192, 
    0.00310411, 0.0002905496, 1.910961e-05, 8.687918e-05, 7.011554e-05, 
    -1.250864e-06,
  0.0348955, 0.07731769, 0.06558009, 0.01630569, 0.001731993, 0.01524035, 
    0.03650827, 0.0446514, 0.05418113, 0.04937633, 0.06170382, 0.06231773, 
    0.1802253, 0.09708227, 0.04468817, 0.02118162, 0.02811015, 0.01667512, 
    0.01740091, 0.02134825, 0.005169368, 0.002651707, 0.05144576, 0.1943893, 
    0.1183493, 0.0852958, 0.08708277, 0.01634609, 0.009715112,
  0.03231825, 0.01813387, 0.01476712, 0.3093855, 0.001753733, 0.02282936, 
    0.07733691, 0.04091631, 0.1108103, 0.1130611, 0.1221924, 0.1265345, 
    0.1498069, 0.09307659, 0.06868931, 0.05875729, 0.07885776, 0.04829236, 
    0.09364306, 0.03878241, 0.08584915, 0.1445812, 0.1400214, 0.06980962, 
    0.07328913, 0.05734945, 0.0786826, 0.1681006, 0.09316546,
  0.01881025, 0.009439868, 7.660635e-06, -6.268733e-06, -2.48416e-07, 
    0.01448437, 0.1456062, 0.1366131, 0.1917249, 0.1622705, 0.1437481, 
    0.08657566, 0.04163047, 0.005623891, 0.01347231, 0.008798181, 0.00393762, 
    3.30498e-05, 0.008388388, 0.0001746573, 0.007475464, 0.06708349, 
    0.04423078, 0.05969326, 0.00752461, 0.0124211, 0.02048875, 0.0189417, 
    0.02259495,
  0.0006325567, 0.02926118, 0.001011336, 0.0004986578, 5.081203e-05, 
    -7.074106e-05, 0.01174001, 0.1026915, 0.2704392, 0.06383312, 0.196697, 
    0.1703028, 0.11692, 0.06468487, 0.09517694, 0.04434443, 0.05122654, 
    0.01242483, 0.005272631, 6.899155e-06, 0.003749813, 0.01427877, 
    0.0322744, 0.04147004, 0.1198099, 0.02670008, 0.001982846, 9.317287e-05, 
    0.0008305238,
  0.06146808, 0.05351647, 0.02715367, 0.05975033, 0.04620329, 0.007621282, 
    0.1423768, 0.05105279, 0.05376938, 0.09602876, 0.1444394, 0.06967928, 
    0.1444702, 0.1442354, 0.0952546, 0.1739431, 0.1281638, 0.05119119, 
    0.03046773, 0.02116308, 0.04666082, 0.04837165, 0.05942476, 0.06331089, 
    0.09430224, 0.1256487, 0.05614373, 0.03162356, 0.0181297,
  0.1004327, 0.1274025, 0.1317883, 0.07399631, 0.09219337, 0.07234477, 
    0.09219207, 0.09959925, 0.163253, 0.1467672, 0.1732242, 0.1728474, 
    0.09239517, 0.1400469, 0.1559707, 0.2130883, 0.203387, 0.1815056, 
    0.1582405, 0.08229022, 0.1574247, 0.09322105, 0.09679605, 0.1022729, 
    0.141939, 0.1703449, 0.1380886, 0.1139257, 0.0974451,
  0.1390262, 0.06647106, 0.07453346, 0.1173733, 0.1053161, 0.1967023, 
    0.1340853, 0.1160188, 0.163808, 0.1346799, 0.119517, 0.164797, 0.157746, 
    0.1457203, 0.1476084, 0.2031864, 0.2435594, 0.2869726, 0.1211012, 
    0.08267821, 0.07900423, 0.08889138, 0.1709597, 0.2430274, 0.2185712, 
    0.2936259, 0.2089039, 0.2020754, 0.147157,
  0.1702607, 0.1117168, 0.1898941, 0.0927379, 0.1433556, 0.2347769, 0.173281, 
    0.1310603, 0.09413359, 0.1532409, 0.1147499, 0.1428537, 0.1073646, 
    0.0987239, 0.0915705, 0.08136865, 0.1029151, 0.1520598, 0.1606661, 
    0.1513952, 0.1681595, 0.1472828, 0.1666984, 0.1362998, 0.04459662, 
    0.328339, 0.3083252, 0.1718666, 0.1802961,
  0.1145665, 0.1691506, 0.1609301, 0.1864577, 0.1992927, 0.2550941, 
    0.2291383, 0.2239448, 0.2035056, 0.2084256, 0.1701319, 0.1684518, 
    0.1851583, 0.2347241, 0.2917084, 0.2180579, 0.1870746, 0.1581855, 
    0.144492, 0.2572633, 0.2487443, 0.2351879, 0.2329816, 0.1303764, 
    0.1293814, 0.1168472, 0.1134016, 0.09348749, 0.1413083,
  5.368079e-07, 1.725998e-07, -1.916084e-07, -5.558165e-07, -9.200247e-07, 
    -1.284233e-06, -1.648441e-06, -0.0001981455, -0.0001309775, 
    -6.380957e-05, 3.358398e-06, 7.052636e-05, 0.0001376943, 0.0002048623, 
    -0.000764931, -0.0007384217, -0.0007119124, -0.0006854031, -0.0006588938, 
    -0.0006323846, -0.0006058753, 0.0003097511, 0.0002164381, 0.000123125, 
    2.981199e-05, -6.350106e-05, -0.0001568141, -0.0002501272, 8.281744e-07,
  0.01163819, 0.003767408, -0.0001790118, 0, 0, -0.0005703578, -0.0003345808, 
    -2.047966e-05, -1.433485e-07, 0.0003910089, 0.004874893, 0.00116615, 
    0.0159754, 0.214705, 0.2266869, 0.2192116, 0.2141437, 0.2173992, 
    0.2020208, 0.2176675, 0.1540704, 0.1537868, 0.2243134, 0.353897, 
    0.315504, 0.2410577, 0.2675128, 0.2177356, 0.03712843,
  0.1557521, 0.2949919, 0.269731, 0.3121399, 0.1528224, 0.2077645, 0.3090032, 
    0.2110054, 0.1836965, 0.1856647, 0.1857476, 0.1784337, 0.2298434, 
    0.2743035, 0.2296193, 0.1803271, 0.2080867, 0.2963893, 0.2801885, 
    0.3248003, 0.3082867, 0.3354982, 0.2660869, 0.3507524, 0.3106323, 
    0.1856479, 0.2276273, 0.2869618, 0.2180476,
  0.2391433, 0.2953082, 0.3084752, 0.2878553, 0.310446, 0.2938536, 0.2483767, 
    0.2131146, 0.2432112, 0.3465125, 0.2814971, 0.2742511, 0.2524704, 
    0.2098209, 0.2492453, 0.2171412, 0.1893232, 0.2068031, 0.213254, 
    0.1988215, 0.2361178, 0.2117096, 0.3008175, 0.2441261, 0.2578296, 
    0.2175792, 0.2376704, 0.1884661, 0.2182395,
  0.1803423, 0.1573103, 0.1764792, 0.1521203, 0.1736843, 0.166329, 0.1559521, 
    0.2215755, 0.1810354, 0.1965057, 0.2223125, 0.1996026, 0.179555, 
    0.1956593, 0.1904113, 0.1211326, 0.2134354, 0.1764361, 0.1925074, 
    0.1755015, 0.1812687, 0.2166197, 0.1439761, 0.1155254, 0.1248586, 
    0.1541986, 0.1850969, 0.2081209, 0.1868547,
  0.07868938, 0.1262129, 0.08837803, 0.1334568, 0.1449448, 0.1045296, 
    0.08462933, 0.1080482, 0.1206653, 0.1083544, 0.167492, 0.1331607, 
    0.1030768, 0.1403856, 0.1348953, 0.1049099, 0.126762, 0.1248026, 
    0.1350619, 0.1135904, 0.1085153, 0.1362515, 0.1637029, 0.2146447, 
    0.07306536, 0.09971611, 0.1229255, 0.08845122, 0.08782268,
  0.04885885, 0.008068403, 0.03133205, 0.06567448, 0.03408743, 0.02808117, 
    0.01839456, 0.02963476, 0.03595886, 0.01887918, 0.03365741, 0.03686428, 
    0.02557302, 0.05082464, 0.06246749, 0.1330031, 0.0764517, 0.0844181, 
    0.1314935, 0.2034103, 0.05891536, 0.0310304, 0.02850936, 0.004507124, 
    0.02767868, 0.1003886, 0.05352238, 0.04859565, 0.04385085,
  1.425008e-07, 1.505126e-08, 0.001212656, -1.692305e-05, 0.04799538, 
    0.01906161, 0.003836684, 0.04457283, 0.001406946, 0.01152275, 
    0.009384482, 0.001101744, 0.01918397, 0.07155582, 0.04482567, 0.02990519, 
    0.03193276, 0.05020056, 0.03369711, 0.02958978, 0.01772395, 4.723699e-05, 
    2.637899e-08, 2.096947e-05, 0.004230052, 0.0002347015, 0.004558626, 
    0.002652634, 0.001357818,
  1.842562e-05, 3.013033e-05, 1.432496e-05, 0.0148292, 0.06296898, 
    0.04030404, 0.02247385, 0.03841116, 0.0539609, 0.01815575, 0.04926164, 
    0.02295759, 0.1090055, 0.07893553, 0.07011965, 0.07980362, 0.06873437, 
    0.01071952, 0.002802093, -1.575209e-08, 1.025642e-06, 5.200651e-07, 
    0.0003115591, 0.004568634, 0.0002578849, 4.474646e-05, 0.0003225137, 
    0.0005896876, 3.60459e-05,
  0.0289722, 0.1028103, 0.0696741, 0.01474967, 0.001613123, 0.01412168, 
    0.03413731, 0.04090849, 0.05063161, 0.05464888, 0.05985255, 0.04289673, 
    0.1413847, 0.08390551, 0.03865965, 0.02281922, 0.02687167, 0.01074512, 
    0.01626399, 0.01387073, 0.006495108, 0.01338952, 0.04641071, 0.2373293, 
    0.1323553, 0.07547943, 0.08271386, 0.01378413, 0.01834697,
  0.02578347, 0.01210793, 0.008988531, 0.2142042, 0.002113731, 0.01465246, 
    0.07893914, 0.02916079, 0.04848925, 0.07659902, 0.07697001, 0.08463599, 
    0.1165283, 0.07536374, 0.05341767, 0.04519479, 0.06263767, 0.05187205, 
    0.09700507, 0.03839925, 0.07984539, 0.1206872, 0.1380169, 0.07034374, 
    0.0679647, 0.06791968, 0.0725258, 0.1437602, 0.105301,
  0.01679934, 0.001670735, 4.094294e-06, 1.121721e-07, 5.67099e-06, 
    0.002452538, 0.1283892, 0.07341203, 0.2120718, 0.1344683, 0.1162958, 
    0.07007954, 0.03114701, 0.006833247, 0.01606432, 0.008449304, 
    0.004048119, -8.934594e-05, 0.001162932, 0.0002738546, 0.004314717, 
    0.05945302, 0.03550314, 0.0501924, 0.006924307, 0.009359717, 0.01163534, 
    0.0107361, 0.01849292,
  0.0003023827, 0.01459625, 3.723273e-05, 2.895311e-06, -1.175685e-05, 
    -1.28706e-05, 0.009485736, 0.1219934, 0.2888244, 0.05747198, 0.1600833, 
    0.1486541, 0.1204649, 0.06383631, 0.09810709, 0.04434142, 0.05657962, 
    0.01047618, 0.008232968, 1.205291e-06, 0.001833347, 0.01388338, 
    0.03221311, 0.04988225, 0.1343861, 0.02774509, 0.0030147, 0.0002997163, 
    0.0006479856,
  0.07563746, 0.04954095, 0.03061321, 0.06333093, 0.035105, 0.006850813, 
    0.126118, 0.04401238, 0.03178406, 0.08392653, 0.1740597, 0.07303373, 
    0.1420065, 0.1475948, 0.1039109, 0.1947847, 0.1451439, 0.05983955, 
    0.03422128, 0.02173679, 0.02751858, 0.04885606, 0.07155771, 0.06915956, 
    0.09695151, 0.1355831, 0.07199411, 0.0338002, 0.028822,
  0.1005349, 0.1280226, 0.1452629, 0.09632327, 0.07115781, 0.07880089, 
    0.09368038, 0.1056808, 0.1479982, 0.1471845, 0.1836789, 0.1711415, 
    0.1047208, 0.1424488, 0.199345, 0.2245884, 0.2141839, 0.1867962, 
    0.1750878, 0.1028607, 0.152593, 0.09783784, 0.1127167, 0.1047768, 
    0.1532313, 0.1792573, 0.1425436, 0.1122315, 0.1073617,
  0.1500717, 0.06895237, 0.07782418, 0.1220387, 0.1294403, 0.1876855, 
    0.1390014, 0.1487448, 0.1817497, 0.1469966, 0.1264179, 0.1983242, 
    0.1584102, 0.1534784, 0.1459018, 0.1872256, 0.2523046, 0.3072457, 
    0.1236928, 0.08553417, 0.0899518, 0.1012063, 0.1796812, 0.2549922, 
    0.2015965, 0.2947999, 0.2243201, 0.2258761, 0.1661365,
  0.187085, 0.1201923, 0.1941532, 0.1087265, 0.1513016, 0.2341195, 0.2147982, 
    0.1197769, 0.09308705, 0.1482253, 0.1047582, 0.1653684, 0.1840972, 
    0.1194835, 0.09399652, 0.1101827, 0.1302787, 0.1568548, 0.1645977, 
    0.1567064, 0.1867592, 0.1479839, 0.1697188, 0.132914, 0.04572947, 
    0.3343267, 0.3176549, 0.166793, 0.1886149,
  0.1750282, 0.1778867, 0.1775933, 0.2028597, 0.2322555, 0.2529662, 
    0.2165262, 0.2019307, 0.2153715, 0.2167332, 0.1388994, 0.172132, 
    0.1810027, 0.2773918, 0.2797631, 0.2207436, 0.2366826, 0.2551526, 
    0.2062855, 0.2612549, 0.2951276, 0.2572206, 0.2649629, 0.1548163, 
    0.1270459, 0.1126435, 0.1030128, 0.1446557, 0.2138034,
  0.001152415, 0.0006428289, 0.0001332425, -0.0003763439, -0.0008859303, 
    -0.001395517, -0.001905103, -0.0006127742, -0.000392595, -0.0001724158, 
    4.776339e-05, 0.0002679426, 0.0004881218, 0.000708301, -0.002355323, 
    -0.001812823, -0.001270323, -0.0007278225, -0.0001853225, 0.0003571776, 
    0.0008996776, -0.0009092604, -0.001162353, -0.001415446, -0.001668539, 
    -0.001921632, -0.002174725, -0.002427818, 0.001560084,
  0.03121779, 0.008555475, 0.0002000662, 0, -0.0002416821, 0.001719433, 
    0.003363715, -0.001590731, 0.0004259922, 0.007662481, 0.00936624, 
    0.006993625, 0.03556192, 0.2269151, 0.2231742, 0.2215777, 0.1918569, 
    0.2303767, 0.2069233, 0.2306295, 0.23608, 0.2440673, 0.240187, 0.3681071, 
    0.3101707, 0.1934495, 0.2601966, 0.2295816, 0.07989848,
  0.1595715, 0.3095069, 0.2882236, 0.3218044, 0.2259613, 0.2397142, 0.349614, 
    0.3188863, 0.2496462, 0.213289, 0.2021256, 0.1883464, 0.2379601, 
    0.2929222, 0.2402841, 0.2007657, 0.2231297, 0.3105329, 0.3124273, 
    0.3428435, 0.3182523, 0.347939, 0.297611, 0.3529484, 0.3058694, 
    0.1746807, 0.2249955, 0.2996546, 0.2110982,
  0.2655142, 0.2923715, 0.3094258, 0.3086167, 0.3243489, 0.3114331, 
    0.3015773, 0.2642027, 0.2693432, 0.3873627, 0.2973729, 0.2845672, 
    0.2669036, 0.1896501, 0.2358151, 0.1974042, 0.226776, 0.2050427, 
    0.2228017, 0.2228928, 0.2636613, 0.2568942, 0.2907738, 0.2268436, 
    0.243398, 0.2403561, 0.2569024, 0.2287402, 0.2838154,
  0.1980622, 0.1638837, 0.2098191, 0.1703372, 0.1916517, 0.1725544, 
    0.1697561, 0.2172637, 0.2058456, 0.2102567, 0.2263487, 0.2051572, 
    0.1813941, 0.1859068, 0.199596, 0.1404058, 0.2032848, 0.2018486, 
    0.1953747, 0.1679332, 0.1676002, 0.2077546, 0.1407584, 0.1255427, 
    0.1286395, 0.1591782, 0.1855561, 0.1959292, 0.1917056,
  0.09954944, 0.1417632, 0.1036525, 0.1315688, 0.1555928, 0.1120368, 
    0.1013022, 0.1147418, 0.1324218, 0.1195482, 0.1641011, 0.135051, 
    0.1161714, 0.1523156, 0.1421053, 0.1170584, 0.1389933, 0.1272171, 
    0.1294775, 0.1059706, 0.117824, 0.1256049, 0.1585217, 0.2121013, 
    0.09333554, 0.1096435, 0.1337626, 0.0987906, 0.09783956,
  0.05976294, 0.01349237, 0.03820156, 0.06673993, 0.03747161, 0.03520645, 
    0.02656436, 0.03762148, 0.03731722, 0.02879889, 0.03514584, 0.04379397, 
    0.023338, 0.05798204, 0.07308269, 0.1358761, 0.08090607, 0.09237176, 
    0.1381411, 0.2242083, 0.07337755, 0.04017369, 0.04339254, 0.004325045, 
    0.0440532, 0.1123878, 0.06051278, 0.05483004, 0.05254053,
  1.104011e-07, -5.774617e-06, 0.00200091, 0.002811234, 0.04030528, 
    0.01564785, 0.004190312, 0.0586628, 0.0009472262, 0.01231625, 
    0.004788448, 0.0004324306, 0.02795212, 0.07451756, 0.04575091, 0.0241634, 
    0.02992843, 0.05577201, 0.05444742, 0.04488231, 0.02139986, 0.0009675385, 
    -3.101671e-07, 9.287942e-06, 0.01008545, 0.0006026392, 0.01210477, 
    0.004098348, 0.001560811,
  3.301589e-06, -4.276254e-06, 3.676669e-05, 0.0180993, 0.06559305, 
    0.04072855, 0.01915351, 0.04250463, 0.05031729, 0.01393142, 0.04810791, 
    0.02637171, 0.1039348, 0.06594519, 0.06833886, 0.07485065, 0.07589214, 
    0.01692947, 0.004523485, 2.022863e-05, 1.411351e-06, 4.129361e-07, 
    7.060356e-05, 0.007274925, 0.0004410919, 0.0002255354, 0.002053545, 
    0.0006641423, 2.052713e-05,
  0.01540731, 0.07118928, 0.05584427, 0.01345741, 0.001520555, 0.0125048, 
    0.03269805, 0.03125734, 0.04031174, 0.04751994, 0.05343153, 0.03183084, 
    0.1106132, 0.07768948, 0.03738102, 0.02039808, 0.02744669, 0.009047785, 
    0.008755783, 0.005167771, 0.00399111, 0.009060916, 0.03233451, 0.238393, 
    0.1484607, 0.06836418, 0.093235, 0.01437619, 0.01040598,
  0.01984405, 0.01141855, 0.01038187, 0.1233862, 0.004453873, 0.00772444, 
    0.08258359, 0.02803541, 0.03098503, 0.0604427, 0.04955768, 0.06495228, 
    0.1024647, 0.06076938, 0.04885674, 0.04493923, 0.04848289, 0.05540165, 
    0.0960636, 0.04015856, 0.07444413, 0.09956185, 0.1166816, 0.06833201, 
    0.06230441, 0.07276182, 0.06526512, 0.1158355, 0.06897421,
  0.008901387, 5.99833e-05, 2.512225e-06, 1.104356e-07, 3.86609e-06, 
    0.0001455292, 0.1209435, 0.06276789, 0.1822758, 0.1339434, 0.1087863, 
    0.05664222, 0.02498424, 0.008062779, 0.01650975, 0.008424301, 
    0.003194845, 1.44898e-05, 3.697992e-05, 0.0003968499, 0.001734811, 
    0.05728719, 0.02664325, 0.02650747, 0.009296648, 0.004588032, 
    0.004743812, 0.001535487, 0.007529292,
  0.0002914482, 0.002018073, 5.70499e-06, 4.446276e-06, -8.556801e-06, 
    -4.78685e-07, 0.006543782, 0.187442, 0.3185549, 0.0549379, 0.1306794, 
    0.1384149, 0.11201, 0.05239592, 0.08431077, 0.03523817, 0.05865456, 
    0.0112662, 0.008157228, 7.976854e-07, 3.834541e-05, 0.01194547, 
    0.0359764, 0.04122797, 0.1096586, 0.02676824, 0.005933509, 0.001198166, 
    0.0004209805,
  0.08169389, 0.05116424, 0.03178084, 0.06524438, 0.0212773, 0.006160484, 
    0.1062093, 0.0405161, 0.01954484, 0.0740555, 0.1895447, 0.08275069, 
    0.1425654, 0.1385944, 0.1147804, 0.1843195, 0.1500669, 0.06776525, 
    0.03659403, 0.02332437, 0.01829661, 0.0470546, 0.07755642, 0.06059721, 
    0.09908693, 0.1377078, 0.06827036, 0.03608203, 0.03565392,
  0.1141791, 0.1369492, 0.1607825, 0.09804334, 0.06034458, 0.06771316, 
    0.06487383, 0.09851696, 0.1364306, 0.1456238, 0.1969532, 0.187941, 
    0.1021997, 0.1449506, 0.2205174, 0.2558205, 0.2442024, 0.219208, 
    0.1739298, 0.1319746, 0.1649719, 0.09582155, 0.1184019, 0.1293028, 
    0.1645877, 0.1977177, 0.1489841, 0.1485114, 0.1180289,
  0.1531247, 0.07845138, 0.09470212, 0.1221227, 0.1368608, 0.1897914, 
    0.1535381, 0.1463182, 0.2037628, 0.1640837, 0.1388877, 0.2415083, 
    0.1785834, 0.1646257, 0.1603289, 0.197241, 0.2632397, 0.3528753, 
    0.1464543, 0.09533663, 0.1097945, 0.1144478, 0.1878411, 0.2685199, 
    0.1845421, 0.2950473, 0.2350004, 0.2186143, 0.1683139,
  0.1938587, 0.1204881, 0.1867071, 0.09962621, 0.1931026, 0.2602632, 
    0.2011677, 0.1293986, 0.1222183, 0.1625973, 0.1132446, 0.1489131, 
    0.1432494, 0.1291295, 0.1239092, 0.1174577, 0.1387721, 0.1602213, 
    0.1617125, 0.1476302, 0.1858432, 0.1524964, 0.188732, 0.1608194, 
    0.0447083, 0.3225552, 0.3040428, 0.168276, 0.2094982,
  0.1700744, 0.2271174, 0.2286521, 0.2048837, 0.1798283, 0.2012765, 
    0.1826456, 0.1916059, 0.1634427, 0.1705523, 0.112909, 0.1291226, 
    0.1713921, 0.2158453, 0.2792341, 0.2492678, 0.2196826, 0.2348593, 
    0.2066689, 0.2623079, 0.2627006, 0.2307086, 0.2890704, 0.1621119, 
    0.1417501, 0.1214754, 0.1250866, 0.1398431, 0.2072535,
  0.0253783, 0.02193014, 0.01848198, 0.01503382, 0.01158565, 0.008137492, 
    0.004689331, 0.006334284, 0.007418212, 0.008502138, 0.009586065, 
    0.01066999, 0.01175392, 0.01283785, 0.01124097, 0.01655561, 0.02187024, 
    0.02718487, 0.03249951, 0.03781414, 0.04312877, 0.05176188, 0.04881148, 
    0.04586109, 0.04291069, 0.03996029, 0.03700989, 0.03405949, 0.02813683,
  0.06936412, 0.01487099, 0.004953799, -0.0001478566, 0.004512099, 
    0.01122791, 0.01633328, 0.0173448, 0.004014511, 0.01459065, 0.008926352, 
    0.03849886, 0.06561556, 0.2266181, 0.2190876, 0.2252659, 0.1918977, 
    0.221317, 0.212781, 0.2164935, 0.2529761, 0.3045513, 0.2460426, 
    0.3791951, 0.2995474, 0.1757776, 0.2538093, 0.2211389, 0.1203248,
  0.1757193, 0.2898429, 0.3090376, 0.3365758, 0.2702934, 0.2523805, 
    0.3759159, 0.4205623, 0.3144407, 0.2156802, 0.2189659, 0.2009371, 
    0.2426404, 0.319338, 0.274464, 0.2270255, 0.2368813, 0.2812237, 0.310156, 
    0.3457466, 0.3131462, 0.3107247, 0.2799284, 0.3800275, 0.3029919, 
    0.1365132, 0.2111143, 0.2902106, 0.2068722,
  0.3017669, 0.3368199, 0.3604162, 0.3309407, 0.3596496, 0.370726, 0.3097371, 
    0.2805877, 0.3099336, 0.3807784, 0.2959422, 0.2969543, 0.2649813, 
    0.2106161, 0.2669898, 0.2513306, 0.2405641, 0.2121185, 0.2478686, 
    0.2866355, 0.3120623, 0.253658, 0.3029713, 0.2308372, 0.2506946, 
    0.2506816, 0.2515727, 0.2039081, 0.2760314,
  0.224416, 0.2035743, 0.2472959, 0.199479, 0.2107342, 0.1724294, 0.1773023, 
    0.2290129, 0.2069226, 0.2323386, 0.2245748, 0.1959303, 0.1906884, 
    0.1874859, 0.2044047, 0.1637597, 0.2369016, 0.194255, 0.2092796, 
    0.1811993, 0.1925068, 0.2128097, 0.1588978, 0.1346944, 0.1333017, 
    0.166567, 0.1844463, 0.2107131, 0.1890482,
  0.1395142, 0.165775, 0.1330715, 0.138882, 0.1843413, 0.1241457, 0.1275605, 
    0.1347149, 0.1514183, 0.132132, 0.179908, 0.1460851, 0.1371577, 
    0.1691832, 0.1620197, 0.1230684, 0.1664595, 0.1286576, 0.1390176, 
    0.1190635, 0.1507932, 0.1272835, 0.1601495, 0.2176872, 0.1096298, 
    0.128833, 0.1435269, 0.1085234, 0.1234548,
  0.07675244, 0.0201672, 0.05657787, 0.06623218, 0.0463047, 0.04148106, 
    0.03444862, 0.05542405, 0.04241434, 0.03297694, 0.03478188, 0.04531612, 
    0.03451537, 0.06861697, 0.08905268, 0.1480476, 0.08702622, 0.104036, 
    0.1458533, 0.2344866, 0.08958971, 0.04779251, 0.05936199, 0.005146791, 
    0.05984917, 0.1291625, 0.06830022, 0.0653927, 0.06299166,
  1.537072e-07, -5.699314e-06, 0.01460431, 0.006641349, 0.05099361, 
    0.01616588, 0.007923717, 0.07810781, 0.00518701, 0.01373332, 0.0033715, 
    -2.110701e-05, 0.03066498, 0.06458428, 0.06286489, 0.01535872, 
    0.03128763, 0.06687969, 0.07084035, 0.07311713, 0.02701318, 0.002691034, 
    7.391075e-06, 9.083215e-06, 0.02607752, 0.002624656, 0.03044386, 
    0.009005168, 0.005637384,
  2.259105e-06, -2.245009e-05, 0.0001377556, 0.05252822, 0.07009304, 
    0.04763223, 0.02194456, 0.0433395, 0.05027846, 0.01161333, 0.0504365, 
    0.0328548, 0.1120884, 0.0649301, 0.06316984, 0.0736884, 0.08500639, 
    0.02098269, 0.009898285, 6.110232e-05, 8.168578e-07, 1.757129e-07, 
    5.673714e-06, 0.009146214, 0.001031896, 0.0070407, 0.0099897, 
    0.0008010686, 1.281447e-05,
  0.007819382, 0.0718478, 0.05895743, 0.01197098, 0.001805089, 0.01146241, 
    0.03412767, 0.02892386, 0.03637297, 0.04888386, 0.05518902, 0.02422656, 
    0.09726305, 0.07216142, 0.04011892, 0.02472618, 0.03211596, 0.0146378, 
    0.01412074, 0.001956732, 0.001460337, 0.002492079, 0.03604645, 0.2526806, 
    0.1695473, 0.06267491, 0.1023043, 0.01749595, 0.006749067,
  0.01780479, 0.006787268, 0.007110797, 0.05348846, 0.002425977, 0.006977234, 
    0.09040573, 0.02412664, 0.0238569, 0.05170191, 0.03122266, 0.06109681, 
    0.09215792, 0.05633915, 0.04792953, 0.04258751, 0.04743191, 0.06551114, 
    0.09727594, 0.03672023, 0.07678777, 0.08904018, 0.1082999, 0.06681934, 
    0.05902781, 0.07619494, 0.05563774, 0.1027939, 0.06115482,
  0.001197728, 1.756233e-05, 1.646429e-06, 6.882274e-08, 9.095871e-07, 
    -4.498533e-05, 0.1132282, 0.06095913, 0.1835285, 0.1287003, 0.1037677, 
    0.05446128, 0.02555403, 0.0143629, 0.01868148, 0.01633838, 0.002602508, 
    9.675271e-05, -6.606115e-07, 0.0004062345, 0.000712745, 0.05399645, 
    0.02330993, 0.02990677, 0.01397896, 0.00947931, 9.918452e-05, 
    0.0003486986, 0.007083148,
  0.0002829299, 9.109078e-05, 1.911496e-06, 2.246442e-06, -8.136371e-06, 
    2.095061e-08, 0.004607441, 0.2347731, 0.3247347, 0.05464887, 0.1200998, 
    0.1335416, 0.09701848, 0.04671443, 0.07074039, 0.05360752, 0.04926528, 
    0.01701365, 0.007232059, 4.817342e-07, -6.901019e-05, 0.01136994, 
    0.03634366, 0.03656067, 0.1021406, 0.02476496, 0.01087908, 0.002732453, 
    0.0002669514,
  0.07182501, 0.04825643, 0.03097098, 0.06376272, 0.01000036, 0.002335483, 
    0.0861252, 0.03533518, 0.01512764, 0.07266904, 0.1922413, 0.08597182, 
    0.140452, 0.1263742, 0.1194057, 0.1691549, 0.1747943, 0.08261631, 
    0.04028281, 0.03527942, 0.01170253, 0.04070213, 0.08047783, 0.05335509, 
    0.07933449, 0.1372892, 0.06480521, 0.0447272, 0.03537336,
  0.162607, 0.1707302, 0.1933376, 0.08651786, 0.07079373, 0.06327072, 
    0.06036536, 0.1065493, 0.1372315, 0.1670385, 0.2142014, 0.2149193, 
    0.1127688, 0.1817193, 0.2397158, 0.2415153, 0.2584152, 0.2362743, 
    0.1780528, 0.1536986, 0.1479254, 0.09577422, 0.1193331, 0.1507185, 
    0.1837882, 0.203058, 0.1493543, 0.1572696, 0.1366897,
  0.1612795, 0.09589522, 0.1032194, 0.1438919, 0.1692068, 0.2201197, 
    0.1786002, 0.1528707, 0.1869048, 0.1637763, 0.1788038, 0.2674208, 
    0.2279618, 0.1939568, 0.1807723, 0.2295624, 0.3062069, 0.4059152, 
    0.1641769, 0.09987147, 0.1169896, 0.1400024, 0.1884188, 0.2936788, 
    0.2082292, 0.2997227, 0.2600086, 0.2298012, 0.1657902,
  0.2399083, 0.1513659, 0.2036805, 0.125715, 0.1894406, 0.2582642, 0.2403965, 
    0.1669666, 0.1944566, 0.2107083, 0.1163933, 0.1509666, 0.1492165, 
    0.1315504, 0.1607463, 0.1326765, 0.1307068, 0.1699183, 0.1672115, 
    0.1556626, 0.1975209, 0.1735119, 0.1917572, 0.1760581, 0.07280126, 
    0.3007462, 0.2920891, 0.1795517, 0.2398239,
  0.1868486, 0.2439066, 0.1993356, 0.2056136, 0.2061515, 0.2473172, 
    0.1991963, 0.1879414, 0.1751047, 0.1917808, 0.1469823, 0.2125815, 
    0.2589685, 0.2799028, 0.3122865, 0.3112893, 0.3086978, 0.3042148, 
    0.2805011, 0.293458, 0.313584, 0.2692172, 0.295027, 0.1658422, 0.1713042, 
    0.1426789, 0.1576526, 0.1401314, 0.2021281,
  0.07457809, 0.07222106, 0.06986403, 0.06750701, 0.06514999, 0.06279296, 
    0.06043594, 0.07588242, 0.07935046, 0.08281851, 0.08628655, 0.08975459, 
    0.09322264, 0.09669068, 0.08492063, 0.08865254, 0.09238444, 0.09611635, 
    0.09984826, 0.1035802, 0.1073121, 0.1021692, 0.09732626, 0.09248334, 
    0.08764041, 0.08279749, 0.07795457, 0.07311164, 0.07646371,
  0.0952231, 0.04832619, 0.00907582, 0.002553397, 0.006405715, 0.0177973, 
    0.02907633, 0.03283221, 0.03902893, 0.01605588, 0.02025024, 0.07477183, 
    0.1158674, 0.226049, 0.2228781, 0.1930545, 0.167549, 0.2144007, 
    0.2149081, 0.2257436, 0.2777268, 0.3350531, 0.264631, 0.3775033, 
    0.2993652, 0.1523705, 0.2715825, 0.2150941, 0.1603681,
  0.1738398, 0.2851045, 0.3491489, 0.3275098, 0.3085654, 0.2579193, 
    0.3998772, 0.478035, 0.3362766, 0.2290141, 0.2230924, 0.2124518, 
    0.2370347, 0.3284739, 0.2391366, 0.2152404, 0.2328506, 0.2867888, 
    0.3203333, 0.32312, 0.3138772, 0.281514, 0.2510852, 0.3695471, 0.2879975, 
    0.118403, 0.1981871, 0.2679335, 0.2006436,
  0.2900654, 0.3269998, 0.3353704, 0.2962281, 0.3299427, 0.3400118, 
    0.2951547, 0.2364571, 0.3145263, 0.3592225, 0.3087188, 0.3101479, 
    0.2956552, 0.2286741, 0.3063533, 0.2722941, 0.2464969, 0.2380289, 
    0.2654136, 0.2833001, 0.2872616, 0.2927886, 0.3119281, 0.2623023, 
    0.2582534, 0.245479, 0.2761685, 0.2524403, 0.2711985,
  0.2431236, 0.2348778, 0.2879372, 0.2231821, 0.2313849, 0.1927911, 
    0.1976772, 0.2472563, 0.2078855, 0.2551672, 0.2515675, 0.218234, 
    0.1934081, 0.1926581, 0.2313668, 0.1679758, 0.2505469, 0.2392044, 
    0.2418626, 0.211645, 0.2056931, 0.2275192, 0.1755368, 0.1498242, 
    0.1263846, 0.1715495, 0.195408, 0.2177081, 0.199167,
  0.1429503, 0.187042, 0.1479458, 0.1512239, 0.1953811, 0.1642567, 0.1583968, 
    0.159354, 0.1786276, 0.1544749, 0.1976345, 0.155011, 0.1401518, 
    0.1878747, 0.1950437, 0.1345535, 0.1844589, 0.1467718, 0.1538661, 
    0.12294, 0.1777839, 0.146333, 0.168209, 0.2281647, 0.1172592, 0.1406119, 
    0.1483783, 0.1219238, 0.1467427,
  0.08311862, 0.02716192, 0.06736559, 0.06386358, 0.03830619, 0.05306571, 
    0.04671789, 0.06027188, 0.05491811, 0.04918759, 0.03173778, 0.03521964, 
    0.05547849, 0.08074433, 0.09915006, 0.1494558, 0.09494812, 0.1049119, 
    0.1506082, 0.2325859, 0.1114972, 0.05993557, 0.06816003, 0.005809508, 
    0.07664984, 0.1233579, 0.08222942, 0.07175466, 0.07746772,
  2.489047e-05, 3.829756e-06, 0.01886628, 0.02088646, 0.06490592, 0.01874371, 
    0.01291775, 0.1020755, 0.02070595, 0.01647392, 0.006142986, 0.008235432, 
    0.02807719, 0.06518919, 0.09746584, 0.01960355, 0.03046346, 0.08238465, 
    0.08446442, 0.08593436, 0.04720728, 0.01128019, 0.0003584133, 
    0.000176902, 0.05533679, 0.006984936, 0.0497024, 0.02901676, 0.008164673,
  1.043998e-06, 0.0001277948, 0.000342135, 0.08358796, 0.08338799, 0.0531104, 
    0.02688839, 0.04441797, 0.0521835, 0.01254456, 0.06539471, 0.05204304, 
    0.1174, 0.07032295, 0.06025286, 0.07468288, 0.08153646, 0.02369631, 
    0.01660631, 0.002800171, 4.184771e-05, 1.298156e-07, 1.34302e-06, 
    0.01109697, 0.01099981, 0.09671139, 0.03127193, 0.001260981, 1.709068e-05,
  0.003252843, 0.0843155, 0.06551322, 0.01455559, 0.003686005, 0.01227677, 
    0.03570385, 0.02648672, 0.03726137, 0.05238417, 0.05668858, 0.01990665, 
    0.09039202, 0.06430417, 0.0408461, 0.03051266, 0.03980269, 0.0238518, 
    0.0193205, 0.001179714, 0.0009245246, 0.00173693, 0.03100062, 0.2587223, 
    0.1805363, 0.05006242, 0.1050506, 0.02170134, 0.005547544,
  0.01740468, 0.004882885, 0.003671488, 0.01669315, 0.000601012, 0.006964397, 
    0.08528528, 0.02286358, 0.01956845, 0.0396542, 0.02304213, 0.05620231, 
    0.08680025, 0.06339225, 0.05152829, 0.04903396, 0.04994264, 0.08004999, 
    0.1020126, 0.04315326, 0.08432783, 0.08425612, 0.1131926, 0.07333124, 
    0.05829667, 0.07712371, 0.05116229, 0.09562073, 0.06028503,
  6.697726e-05, 3.049057e-06, 9.604028e-07, 3.423786e-08, 1.903848e-07, 
    -1.620221e-06, 0.09015102, 0.06082858, 0.1915761, 0.1337471, 0.09647822, 
    0.05456327, 0.02757904, 0.0254844, 0.03006757, 0.02548217, 0.003490088, 
    0.0003176959, 1.891671e-06, 0.001498208, 0.0003709663, 0.05021657, 
    0.02012323, 0.0294915, 0.01842684, 0.02056178, 2.099818e-06, 
    5.532485e-05, 0.004356946,
  0.0003037991, 1.464331e-05, 1.067175e-06, 1.384248e-06, -6.085712e-06, 
    8.625813e-08, 0.003571828, 0.2042642, 0.3103985, 0.05420887, 0.1160867, 
    0.1297933, 0.09036077, 0.05127902, 0.07688085, 0.05100681, 0.05090302, 
    0.02170383, 0.006324694, 1.21276e-06, -5.69794e-06, 0.01056214, 
    0.04551677, 0.03686495, 0.09334117, 0.02832289, 0.01853153, 0.004049147, 
    0.000567784,
  0.04986769, 0.04994235, 0.02939964, 0.06560308, 0.005367421, 0.001037161, 
    0.06657337, 0.02021346, 0.006702513, 0.0516196, 0.2048644, 0.08637349, 
    0.1394513, 0.1216004, 0.1233848, 0.1678589, 0.1727003, 0.07409876, 
    0.04401151, 0.04961815, 0.0110349, 0.03335688, 0.07726957, 0.0554882, 
    0.08160976, 0.1392461, 0.06290588, 0.04001245, 0.03500571,
  0.1433699, 0.1814079, 0.1984355, 0.08040947, 0.05646271, 0.05897889, 
    0.04717975, 0.115294, 0.1485961, 0.1758325, 0.2213653, 0.2190845, 
    0.1047163, 0.1798962, 0.2184445, 0.2807698, 0.2751367, 0.2331677, 
    0.1807135, 0.1783656, 0.1484238, 0.08270191, 0.1081511, 0.1739773, 
    0.1938566, 0.1997314, 0.1597586, 0.1708942, 0.1253204,
  0.1599769, 0.1225735, 0.1168258, 0.1550345, 0.2561238, 0.2474409, 
    0.1986835, 0.1594305, 0.227288, 0.1684421, 0.2138322, 0.3011999, 
    0.2065184, 0.2117121, 0.2445201, 0.231784, 0.3354446, 0.4322588, 
    0.162968, 0.1118434, 0.1271, 0.1464588, 0.1856598, 0.2937071, 0.1897516, 
    0.3022166, 0.2602451, 0.2641987, 0.1854511,
  0.2752711, 0.214351, 0.2184815, 0.1218083, 0.2141753, 0.2660519, 0.2705936, 
    0.1752285, 0.1766341, 0.1870592, 0.1526083, 0.1785208, 0.1589116, 
    0.1532375, 0.1330875, 0.1694067, 0.1510767, 0.1798772, 0.1632281, 
    0.1758973, 0.2054561, 0.1876005, 0.1920821, 0.1454578, 0.06481355, 
    0.2789942, 0.2778041, 0.1872793, 0.285403,
  0.1788011, 0.247308, 0.2016894, 0.227861, 0.2313088, 0.2078823, 0.1881623, 
    0.1997496, 0.1853501, 0.2007402, 0.2020633, 0.2258753, 0.2762646, 
    0.3127582, 0.3134578, 0.3046858, 0.262855, 0.2402626, 0.2038715, 
    0.2748801, 0.3048337, 0.3213281, 0.3244256, 0.2036657, 0.1504682, 
    0.1523896, 0.1515678, 0.1363529, 0.2038496,
  0.1079489, 0.1063224, 0.1046959, 0.1030693, 0.1014428, 0.09981621, 
    0.09818967, 0.1109358, 0.1163907, 0.1218457, 0.1273006, 0.1327555, 
    0.1382105, 0.1436654, 0.1429438, 0.1455709, 0.148198, 0.1508251, 
    0.1534522, 0.1560793, 0.1587064, 0.1521868, 0.1457313, 0.1392758, 
    0.1328203, 0.1263648, 0.1199093, 0.1134539, 0.1092502,
  0.1135766, 0.09725294, 0.02824293, 0.008749545, 0.009909773, 0.03341394, 
    0.06225954, 0.06100531, 0.04457226, 0.01569688, 0.05036396, 0.1000921, 
    0.1580376, 0.2201546, 0.2156698, 0.1584459, 0.1667389, 0.1971117, 
    0.2125894, 0.2183755, 0.2985083, 0.3476931, 0.2952413, 0.3767394, 
    0.2919398, 0.1414213, 0.2734858, 0.1991302, 0.1876617,
  0.183533, 0.2901521, 0.3638712, 0.3185736, 0.3490898, 0.2638068, 0.4225169, 
    0.4751192, 0.3307786, 0.2400606, 0.2306772, 0.2302048, 0.2302082, 
    0.3240762, 0.2316546, 0.1837022, 0.2337049, 0.2679463, 0.3043199, 
    0.2940393, 0.3173409, 0.2850304, 0.2505197, 0.3550381, 0.2633152, 
    0.1409342, 0.2070464, 0.2926578, 0.1935502,
  0.2450653, 0.346398, 0.346506, 0.297048, 0.3462526, 0.2962402, 0.3228641, 
    0.2544627, 0.307531, 0.3568047, 0.2938561, 0.3173918, 0.2925259, 
    0.2507659, 0.288468, 0.2388314, 0.2570945, 0.2210819, 0.2673718, 
    0.2717093, 0.2932928, 0.2982785, 0.3046117, 0.2924767, 0.2405123, 
    0.2449657, 0.2783748, 0.2672837, 0.262685,
  0.2671052, 0.2417088, 0.2924874, 0.2547852, 0.2525798, 0.2085501, 
    0.1998844, 0.2689503, 0.2390145, 0.2739104, 0.255311, 0.2305103, 
    0.2457496, 0.2155653, 0.2625827, 0.1843089, 0.2622182, 0.2871273, 
    0.2916019, 0.2469574, 0.2226225, 0.2376055, 0.1958302, 0.1581274, 
    0.1347482, 0.1812844, 0.2046679, 0.2326694, 0.2355562,
  0.1669775, 0.2068722, 0.1757325, 0.1844488, 0.2066773, 0.1828176, 
    0.1698792, 0.18571, 0.1902065, 0.1891665, 0.2115676, 0.1839757, 
    0.1450929, 0.1948379, 0.2194391, 0.15098, 0.1858574, 0.157984, 0.1662018, 
    0.1379341, 0.1917385, 0.1510155, 0.1980574, 0.244625, 0.1347934, 
    0.1580266, 0.1670197, 0.1523865, 0.1669034,
  0.09397131, 0.041907, 0.06868751, 0.06269678, 0.03907512, 0.06463248, 
    0.06559915, 0.0835672, 0.07059149, 0.06546482, 0.02961079, 0.02711541, 
    0.05602447, 0.08551013, 0.09512374, 0.1391006, 0.09709415, 0.1070755, 
    0.1450264, 0.2243593, 0.1228907, 0.07481764, 0.06863422, 0.004978077, 
    0.09251863, 0.1147828, 0.09624174, 0.07580911, 0.08028272,
  0.006089401, -1.868172e-06, 0.0649491, 0.03200047, 0.06026312, 0.03835398, 
    0.03903702, 0.09041514, 0.02824332, 0.02084208, 0.003528234, 0.01238836, 
    0.02905346, 0.05352765, 0.1167174, 0.0230429, 0.04370542, 0.08678454, 
    0.08127194, 0.09220826, 0.06726265, 0.02185681, 0.001212025, 
    0.0008746557, 0.06263219, 0.02831278, 0.04612104, 0.05544717, 0.01173693,
  -1.970037e-07, 0.0001586215, 0.001117603, 0.1223182, 0.08040655, 
    0.05918488, 0.03303576, 0.04942497, 0.0523685, 0.01898262, 0.08662485, 
    0.07720956, 0.1185574, 0.066139, 0.05163014, 0.06388066, 0.07891849, 
    0.02294573, 0.02159334, 0.01140574, 0.0001895709, -3.965179e-07, 
    2.972735e-07, 0.01110614, 0.006231119, 0.02090259, 0.04402398, 
    0.005656413, 0.001232545,
  0.002198596, 0.08812749, 0.08730454, 0.01935054, 0.01062707, 0.01527185, 
    0.03459922, 0.02328814, 0.04306892, 0.06153749, 0.05981169, 0.01688306, 
    0.0727934, 0.05221575, 0.03645256, 0.02908802, 0.03863814, 0.03094756, 
    0.01979577, 0.002321149, 0.0003292069, 0.001681293, 0.02390882, 
    0.2566374, 0.1858222, 0.03949481, 0.09117137, 0.02007816, 0.003530943,
  0.0170942, 0.003086356, 0.001835827, 0.004479253, 0.0003042953, 
    0.007748158, 0.07447996, 0.02119351, 0.01503499, 0.03273175, 0.01873012, 
    0.04860336, 0.08010844, 0.06103611, 0.05531424, 0.05692597, 0.05372738, 
    0.08626065, 0.1009116, 0.04737628, 0.08655638, 0.081075, 0.119002, 
    0.08350671, 0.05568799, 0.08454838, 0.06030218, 0.08430689, 0.05153783,
  1.21356e-05, 1.694908e-06, 5.021103e-07, 2.644077e-08, 6.57358e-08, 
    -1.373301e-06, 0.07385625, 0.05718881, 0.1897151, 0.1283436, 0.08837667, 
    0.04986034, 0.02969313, 0.03076966, 0.03574378, 0.03458012, 0.01654458, 
    0.004370399, 1.663369e-06, 0.002978029, 9.364111e-05, 0.04851208, 
    0.0168662, 0.01873951, 0.02814465, 0.02815414, 0.001600762, 1.016954e-06, 
    0.002318742,
  0.0002805835, 6.257703e-06, 5.059441e-07, 1.018504e-06, -1.624142e-06, 
    7.132822e-08, 0.001892583, 0.1424849, 0.3146089, 0.04944177, 0.1159906, 
    0.1344785, 0.08047009, 0.05027534, 0.09024178, 0.0444142, 0.07558469, 
    0.0351572, 0.004729541, 3.375502e-05, 2.363619e-06, 0.01338334, 
    0.04749675, 0.04157958, 0.07794519, 0.03759981, 0.04029875, 0.004504044, 
    0.001314634,
  0.03918199, 0.03490965, 0.028259, 0.06750216, 0.002047169, 0.0002901161, 
    0.05073565, 0.008979652, 0.00253676, 0.0360691, 0.2144111, 0.08154446, 
    0.1309717, 0.1232281, 0.1060753, 0.1963166, 0.1658291, 0.07739614, 
    0.0422556, 0.05246057, 0.0047072, 0.02960153, 0.06983174, 0.05221122, 
    0.09404399, 0.1534949, 0.08035514, 0.05492756, 0.0308516,
  0.1307776, 0.2085755, 0.1889172, 0.09969057, 0.04626201, 0.03691593, 
    0.02997975, 0.1190749, 0.1508936, 0.1476802, 0.2277112, 0.2318139, 
    0.09973238, 0.1695657, 0.2205693, 0.3099049, 0.2649541, 0.2282681, 
    0.1675892, 0.1797576, 0.1456473, 0.07172272, 0.1017018, 0.1858084, 
    0.1862674, 0.2047096, 0.1694242, 0.1726781, 0.1242819,
  0.1712913, 0.1187599, 0.1351658, 0.1666287, 0.2723398, 0.2654632, 
    0.1798302, 0.1548285, 0.2378472, 0.1782279, 0.2234819, 0.2915397, 
    0.2116359, 0.2248238, 0.2457297, 0.2265164, 0.3490992, 0.4373622, 
    0.177866, 0.1207576, 0.1184072, 0.1231421, 0.1674659, 0.2763539, 
    0.1697919, 0.2945161, 0.2611738, 0.2672548, 0.1791618,
  0.2754192, 0.1688623, 0.2403384, 0.1182356, 0.225001, 0.2968943, 0.234548, 
    0.1761851, 0.1372788, 0.1652379, 0.1652804, 0.1475643, 0.1625418, 
    0.1315278, 0.09512974, 0.1030762, 0.1277723, 0.1801058, 0.1314406, 
    0.1717884, 0.1838032, 0.1961546, 0.207876, 0.1255868, 0.0612267, 
    0.3057041, 0.284201, 0.1887082, 0.2867728,
  0.1631091, 0.2205642, 0.1915822, 0.1939796, 0.1761969, 0.1717432, 
    0.1590902, 0.173685, 0.142647, 0.1354066, 0.158308, 0.1513291, 0.1716759, 
    0.2696725, 0.2934749, 0.2554534, 0.2366325, 0.1966137, 0.1721261, 
    0.2062212, 0.2479367, 0.2834505, 0.3676309, 0.205774, 0.1567738, 
    0.1485323, 0.1765283, 0.1464871, 0.1945325,
  0.1333422, 0.1322241, 0.1311059, 0.1299877, 0.1288695, 0.1277514, 
    0.1266332, 0.1607573, 0.167433, 0.1741087, 0.1807844, 0.1874602, 
    0.1941359, 0.2008116, 0.1929935, 0.1951208, 0.1972481, 0.1993754, 
    0.2015027, 0.20363, 0.2057573, 0.1909003, 0.1832155, 0.1755307, 
    0.1678458, 0.160161, 0.1524762, 0.1447913, 0.1342368,
  0.1329883, 0.1195185, 0.09021607, 0.01874488, 0.02160902, 0.06924929, 
    0.1096124, 0.0901161, 0.03760284, 0.01659985, 0.0586741, 0.1196236, 
    0.191938, 0.199801, 0.2260256, 0.1565001, 0.1545932, 0.1820316, 
    0.2144383, 0.2136516, 0.3311415, 0.3704467, 0.3488247, 0.3659469, 
    0.2761079, 0.146941, 0.2651308, 0.1847941, 0.2135268,
  0.2054067, 0.2644287, 0.3192752, 0.3029809, 0.353932, 0.2754441, 0.4063676, 
    0.4575696, 0.3204007, 0.2449342, 0.2382596, 0.2379436, 0.2335685, 
    0.3115418, 0.2694376, 0.2115366, 0.2292718, 0.2900446, 0.3479253, 
    0.3096863, 0.3380426, 0.2885509, 0.2442555, 0.3632362, 0.2553765, 
    0.1480478, 0.24874, 0.3294655, 0.216737,
  0.3217999, 0.4174325, 0.3614547, 0.3222666, 0.3810371, 0.3158298, 0.359196, 
    0.2973276, 0.3417836, 0.3949925, 0.3472425, 0.3344528, 0.3468275, 
    0.2915013, 0.2924901, 0.2683313, 0.2745726, 0.2259813, 0.296769, 
    0.3130342, 0.3270628, 0.2980721, 0.363498, 0.3167098, 0.2527776, 
    0.2880176, 0.2913498, 0.2827274, 0.3174551,
  0.29855, 0.2730667, 0.306633, 0.2536209, 0.2682516, 0.2235107, 0.2196707, 
    0.2861574, 0.2510996, 0.3071086, 0.2795554, 0.2584748, 0.2482684, 
    0.2629319, 0.3102239, 0.2334817, 0.2756469, 0.3170688, 0.3299277, 
    0.2657833, 0.2591438, 0.2709499, 0.2302036, 0.1803887, 0.1413493, 
    0.2121169, 0.2416636, 0.2805365, 0.2799062,
  0.2288786, 0.2199242, 0.2051976, 0.2152827, 0.2411237, 0.204416, 0.1744477, 
    0.2007147, 0.2138929, 0.205556, 0.2233025, 0.1922659, 0.1484158, 
    0.1979253, 0.2395822, 0.1565316, 0.1964067, 0.174687, 0.2125289, 
    0.1860226, 0.1827472, 0.172065, 0.2260768, 0.2661422, 0.1525135, 
    0.1823267, 0.1982452, 0.1804292, 0.1868619,
  0.1350604, 0.06209732, 0.05337127, 0.07938035, 0.06142025, 0.103947, 
    0.07984334, 0.1085916, 0.1003303, 0.1071415, 0.01364823, 0.03615911, 
    0.04198132, 0.08283564, 0.09109364, 0.1421014, 0.1098128, 0.1234189, 
    0.1432798, 0.2079468, 0.1444525, 0.08934608, 0.09568596, 0.005537709, 
    0.1073299, 0.1314726, 0.09301192, 0.06873541, 0.09319055,
  0.02430541, -1.25821e-05, 0.01223156, 0.03473865, 0.06354894, 0.05119444, 
    0.07096583, 0.109374, 0.09909293, 0.03899311, 0.001036703, 0.01333174, 
    0.053079, 0.05310224, 0.1365045, 0.02979371, 0.07832622, 0.1001899, 
    0.09221109, 0.09630045, 0.1052191, 0.06504361, 0.0102878, 0.001878353, 
    0.06212021, 0.07074397, 0.03911274, 0.06341214, 0.0765378,
  1.119047e-06, -2.898765e-05, 0.002888652, 0.14073, 0.07371454, 0.05616, 
    0.03364202, 0.0550229, 0.05257129, 0.0321273, 0.1058986, 0.09290623, 
    0.1254489, 0.05806259, 0.04377247, 0.05330264, 0.06464811, 0.02341298, 
    0.02002533, 0.01996664, 0.002121398, 0.0001413448, 3.534515e-07, 
    0.01663916, 0.006228455, 0.001129897, 0.04215702, 0.01709785, 0.01006094,
  0.003192812, 0.09742216, 0.08476494, 0.01510482, 0.01921417, 0.0190462, 
    0.0304944, 0.02298963, 0.04970364, 0.08095209, 0.04516743, 0.01457778, 
    0.06166251, 0.03886237, 0.03237464, 0.02508695, 0.03388439, 0.02852715, 
    0.02053957, 0.007281328, 0.001428064, 0.001904225, 0.01521622, 0.2486617, 
    0.1844703, 0.03192149, 0.07546549, 0.0221164, 0.002301815,
  0.01645808, 0.001737168, 0.0008713559, 0.001026775, 0.0001892395, 
    0.0109017, 0.06490857, 0.01988153, 0.01837914, 0.02734742, 0.01904235, 
    0.04059725, 0.0649095, 0.05418003, 0.05331817, 0.05624842, 0.06150489, 
    0.09653202, 0.1032789, 0.05159105, 0.08478643, 0.08047156, 0.1158804, 
    0.08748376, 0.04830221, 0.09416736, 0.08513831, 0.08030021, 0.04463816,
  2.06765e-06, 1.143042e-06, 2.045922e-07, 2.500573e-08, 4.078509e-08, 
    -3.333158e-05, 0.06066481, 0.05154355, 0.1950437, 0.1205915, 0.07581732, 
    0.04354, 0.02570116, 0.02585228, 0.03053998, 0.02961056, 0.04955891, 
    0.0202149, 0.0003820028, 0.004037564, 0.0002364364, 0.04463148, 
    0.01662355, 0.01239134, 0.02718786, 0.04557363, 0.02020265, 1.725617e-06, 
    0.001438127,
  0.0002068793, 3.232464e-06, 1.906223e-07, 8.355413e-07, 2.908073e-07, 
    4.91218e-08, 0.001013185, 0.09848853, 0.31089, 0.04732632, 0.1129772, 
    0.1507371, 0.06918959, 0.04883845, 0.09487431, 0.05393051, 0.08760047, 
    0.05564097, 0.01916091, 0.0001099255, 2.027209e-06, 0.01355435, 
    0.04232439, 0.04450986, 0.06494468, 0.04583478, 0.08139049, 0.01979659, 
    0.001723443,
  0.02668444, 0.02414716, 0.0237284, 0.07036014, 0.0007542329, 4.366507e-05, 
    0.03629309, 0.005055185, 0.001373141, 0.02893575, 0.2103344, 0.08804677, 
    0.131052, 0.1273151, 0.1321317, 0.2185036, 0.1853848, 0.09168489, 
    0.05882356, 0.05522817, 0.003237722, 0.02772396, 0.06253339, 0.05432609, 
    0.1112788, 0.1794549, 0.1358018, 0.09627222, 0.03436403,
  0.1230794, 0.2030264, 0.1814619, 0.08097343, 0.03331729, 0.02421991, 
    0.02005255, 0.1442095, 0.1472559, 0.1202786, 0.2300152, 0.2260116, 
    0.08509694, 0.1593818, 0.2673683, 0.3352852, 0.2948721, 0.2739244, 
    0.1757377, 0.1676601, 0.1307274, 0.07180807, 0.09598529, 0.1708551, 
    0.1726845, 0.221768, 0.1859846, 0.1780374, 0.1542173,
  0.1884268, 0.1558942, 0.1495867, 0.1625549, 0.2541527, 0.2549743, 
    0.1837226, 0.1789317, 0.2222916, 0.1660322, 0.2314776, 0.2722557, 
    0.2113516, 0.2550014, 0.27462, 0.2443279, 0.3599297, 0.4587293, 
    0.2137043, 0.08829612, 0.1014725, 0.1049583, 0.1387164, 0.2421197, 
    0.1804263, 0.2606928, 0.300078, 0.3057167, 0.1894208,
  0.26634, 0.1756622, 0.2690572, 0.1371786, 0.2597778, 0.2720998, 0.225602, 
    0.1611213, 0.1443951, 0.2017899, 0.1955555, 0.1531326, 0.1381592, 
    0.1358768, 0.1103166, 0.100668, 0.1671603, 0.1565952, 0.1337107, 
    0.1718508, 0.1787079, 0.1918131, 0.2636951, 0.1694484, 0.07413722, 
    0.3337092, 0.2750899, 0.1988031, 0.3053184,
  0.2272687, 0.2710271, 0.2379163, 0.1816679, 0.1675702, 0.2194812, 0.166804, 
    0.1852842, 0.1863527, 0.1861065, 0.1761318, 0.1555873, 0.169358, 
    0.2489181, 0.2784957, 0.2954634, 0.2997503, 0.2529944, 0.252628, 
    0.2674604, 0.2905105, 0.3176885, 0.3224093, 0.2192926, 0.1385014, 
    0.1690778, 0.1706065, 0.1524542, 0.23226,
  0.1601758, 0.1597049, 0.1592341, 0.1587632, 0.1582923, 0.1578215, 
    0.1573506, 0.1998958, 0.2080208, 0.2161458, 0.2242708, 0.2323958, 
    0.2405208, 0.2486458, 0.2523148, 0.2531218, 0.2539288, 0.2547358, 
    0.2555428, 0.2563498, 0.2571568, 0.2251519, 0.2166907, 0.2082296, 
    0.1997685, 0.1913074, 0.1828462, 0.1743851, 0.1605525,
  0.1525485, 0.1498038, 0.1415656, 0.04556727, 0.03936291, 0.1136732, 
    0.1458565, 0.1146159, 0.02417567, 0.03018715, 0.07043757, 0.1308649, 
    0.2096755, 0.1806175, 0.2212099, 0.1828167, 0.1537097, 0.1782057, 
    0.2181759, 0.2222019, 0.3973727, 0.3966293, 0.4045227, 0.3336704, 
    0.2831646, 0.1788033, 0.2417257, 0.1718265, 0.2235495,
  0.2422669, 0.2830902, 0.3052142, 0.2717457, 0.3504555, 0.2962692, 
    0.3961815, 0.4608056, 0.3124938, 0.2462648, 0.2410179, 0.2453337, 
    0.2473012, 0.293483, 0.2996435, 0.2412605, 0.2452962, 0.3279693, 
    0.3353773, 0.3587745, 0.3442121, 0.3025575, 0.2498766, 0.3570184, 
    0.2661113, 0.1829908, 0.2656462, 0.3474667, 0.2276139,
  0.3950022, 0.4271667, 0.3829147, 0.3691247, 0.4297117, 0.3743159, 
    0.4474019, 0.3775258, 0.4286946, 0.4634376, 0.4266521, 0.3974221, 
    0.4049402, 0.3747375, 0.3631867, 0.3068298, 0.2957598, 0.2397584, 
    0.3806996, 0.3373606, 0.3003529, 0.3037256, 0.3754215, 0.3684389, 
    0.3541215, 0.306385, 0.3152586, 0.3164552, 0.3475579,
  0.3115736, 0.2590107, 0.3268482, 0.2588188, 0.252502, 0.2358353, 0.258992, 
    0.3080399, 0.2550176, 0.2602634, 0.3013883, 0.3119876, 0.2583237, 
    0.3084226, 0.3265889, 0.323568, 0.3360299, 0.3751726, 0.3632421, 
    0.3157399, 0.3028364, 0.2821508, 0.2649754, 0.2179639, 0.1681379, 
    0.2232524, 0.2844969, 0.3341876, 0.3160931,
  0.2161821, 0.2244782, 0.1896897, 0.2201115, 0.2468937, 0.2005744, 
    0.1747529, 0.2094843, 0.2160129, 0.1992487, 0.2010211, 0.1732959, 
    0.1378357, 0.1770544, 0.2591992, 0.1729059, 0.1917244, 0.1899026, 
    0.2428186, 0.2380655, 0.2215115, 0.2138433, 0.2238236, 0.2970915, 
    0.1975101, 0.168804, 0.1919156, 0.2493125, 0.2223038,
  0.1501595, 0.09157433, 0.03411119, 0.109303, 0.09391235, 0.1523569, 
    0.1281588, 0.1514879, 0.1550539, 0.1459663, 0.01035138, 0.01848919, 
    0.02896904, 0.09095061, 0.1393751, 0.1604654, 0.1334719, 0.13496, 
    0.162658, 0.2212077, 0.1413424, 0.1098527, 0.1252748, 0.008044044, 
    0.09478336, 0.1611624, 0.1152644, 0.09906314, 0.132898,
  0.137548, -0.0001141147, 0.002204802, 0.05601013, 0.0812321, 0.04848737, 
    0.09466058, 0.1638679, 0.1069047, 0.02700355, 0.0001930398, 0.006762418, 
    0.1210531, 0.1058417, 0.1375286, 0.04514845, 0.09279072, 0.1109534, 
    0.1118265, 0.09693265, 0.1379564, 0.1146509, 0.03478646, 0.0002494465, 
    0.07034751, 0.05277489, 0.05277531, 0.1150537, 0.2160732,
  0.0004431101, -3.791009e-06, 0.008015375, 0.1352212, 0.06719346, 
    0.05108177, 0.04320778, 0.06036128, 0.05080402, 0.04228326, 0.1274778, 
    0.0942132, 0.130477, 0.05085439, 0.03926378, 0.05050981, 0.05471484, 
    0.02374885, 0.02339353, 0.03484342, 0.02056119, 0.01114894, 3.172583e-06, 
    0.03101295, 0.009913483, 0.0001100021, 0.05236477, 0.04023407, 0.03466509,
  0.007959946, 0.1113171, 0.08096057, 0.01194252, 0.02766426, 0.02504386, 
    0.02916376, 0.02548438, 0.0590027, 0.1011042, 0.03420903, 0.01480296, 
    0.04868228, 0.0314462, 0.0298521, 0.02382114, 0.02766903, 0.02375664, 
    0.01778776, 0.01442245, 0.01449179, 0.00643972, 0.00801385, 0.2378437, 
    0.1790382, 0.02961194, 0.06489989, 0.02430585, 0.009999198,
  0.01582953, 0.002156459, 0.0004123046, 6.113293e-05, 9.335377e-05, 
    0.01517535, 0.05819277, 0.02216759, 0.01579021, 0.02527339, 0.02251245, 
    0.03722246, 0.05465617, 0.04730712, 0.05065948, 0.05075432, 0.06575584, 
    0.09992655, 0.107885, 0.05801412, 0.0807997, 0.07106708, 0.1215917, 
    0.08468238, 0.04113229, 0.09363591, 0.09649865, 0.07412521, 0.03912596,
  1.499818e-06, 9.107461e-07, 9.811303e-08, 2.209958e-08, 3.429891e-08, 
    -0.0001594024, 0.0470609, 0.04566931, 0.1930524, 0.1103774, 0.06401915, 
    0.04163379, 0.02749514, 0.02766179, 0.03074431, 0.03067335, 0.06068052, 
    0.07173283, 0.01899334, 0.006632905, 0.001997754, 0.04484056, 0.02096818, 
    0.01017795, 0.0335593, 0.07023479, 0.06360479, 0.0001808388, 0.0008966943,
  0.0001185043, 2.109581e-06, 5.27348e-08, 7.043288e-07, 2.947973e-07, 
    3.774684e-08, 0.0007139921, 0.08267656, 0.321882, 0.04375917, 0.110952, 
    0.1594152, 0.06311297, 0.05067531, 0.1012098, 0.06789535, 0.1245519, 
    0.08937281, 0.07536258, 0.001013885, 1.523838e-06, 0.01391894, 
    0.04439176, 0.0461963, 0.05428489, 0.04713631, 0.1027818, 0.0582415, 
    0.003202325,
  0.01975426, 0.0166772, 0.01101377, 0.07191241, -0.0001653371, 5.201723e-07, 
    0.03108053, 0.002900947, 0.0008292954, 0.02801501, 0.2164524, 0.107078, 
    0.1474009, 0.1460208, 0.2032213, 0.2504637, 0.210991, 0.1244395, 
    0.09931359, 0.04928019, 0.00301244, 0.0288877, 0.05726042, 0.0498483, 
    0.1286321, 0.2030111, 0.1520048, 0.1266664, 0.04986329,
  0.1205587, 0.184827, 0.1617224, 0.04939826, 0.01961981, 0.011503, 
    0.01735652, 0.1372891, 0.1351442, 0.09978488, 0.2098546, 0.2198571, 
    0.0935875, 0.1713711, 0.3012984, 0.3809502, 0.3715512, 0.3100985, 
    0.2003039, 0.1522414, 0.111825, 0.05056682, 0.08559629, 0.1737266, 
    0.1613624, 0.2222503, 0.2294362, 0.2158814, 0.1572115,
  0.1979807, 0.1309903, 0.09329453, 0.1635028, 0.230215, 0.2183079, 0.134776, 
    0.19959, 0.1939855, 0.1501813, 0.1982057, 0.2783974, 0.2134168, 
    0.2600186, 0.3223987, 0.2719806, 0.3275365, 0.4718073, 0.2168726, 
    0.05809069, 0.07574359, 0.08927059, 0.1178009, 0.2185454, 0.1781478, 
    0.2139026, 0.3755705, 0.3566289, 0.2491654,
  0.2979337, 0.213263, 0.2942494, 0.1882679, 0.284537, 0.2549888, 0.2305626, 
    0.1745007, 0.1406249, 0.1692374, 0.189946, 0.158201, 0.1170452, 
    0.1487596, 0.1573834, 0.1652129, 0.2075534, 0.1545109, 0.1218353, 
    0.1811157, 0.1932472, 0.2181466, 0.273303, 0.2173513, 0.0825647, 
    0.3349323, 0.2685515, 0.2078086, 0.3275303,
  0.2999279, 0.3103579, 0.2752548, 0.2181787, 0.2174208, 0.2817996, 
    0.2361875, 0.2411862, 0.2987545, 0.2584473, 0.1748005, 0.2187085, 
    0.2208459, 0.2704653, 0.3065603, 0.3551411, 0.3478225, 0.3986602, 
    0.3203629, 0.3649449, 0.3398953, 0.3259682, 0.291109, 0.2205927, 
    0.1718796, 0.1785747, 0.1507749, 0.1652131, 0.2691881,
  0.1825961, 0.1825614, 0.1825266, 0.1824919, 0.1824572, 0.1824225, 
    0.1823877, 0.2331667, 0.2421895, 0.2512123, 0.2602351, 0.2692579, 
    0.2782807, 0.2873036, 0.2894949, 0.2891946, 0.2888944, 0.2885941, 
    0.2882938, 0.2879935, 0.2876932, 0.2518138, 0.243126, 0.2344382, 
    0.2257504, 0.2170627, 0.2083749, 0.1996871, 0.1826239,
  0.1711527, 0.1674391, 0.1637707, 0.09556073, 0.05860289, 0.1491325, 
    0.1507294, 0.1351825, 0.01947927, 0.0340263, 0.06887453, 0.1303969, 
    0.2276, 0.1278274, 0.2149237, 0.1855505, 0.1618301, 0.1761132, 0.2278742, 
    0.2301092, 0.424208, 0.4178719, 0.4269412, 0.2960956, 0.278648, 
    0.2018766, 0.2047036, 0.1553204, 0.228474,
  0.2672042, 0.2744851, 0.3058797, 0.2424767, 0.3623685, 0.3070356, 
    0.3341994, 0.4475312, 0.3075299, 0.2557831, 0.2416971, 0.2377671, 
    0.2562695, 0.274128, 0.3013467, 0.3288279, 0.3199453, 0.3641948, 
    0.3572396, 0.3721635, 0.3317495, 0.3393998, 0.2616402, 0.3615065, 
    0.2760639, 0.2268283, 0.2996128, 0.3698232, 0.2329386,
  0.4180703, 0.4008158, 0.3531178, 0.3732622, 0.4260439, 0.4405574, 
    0.5217137, 0.4641136, 0.4723462, 0.5240833, 0.4771897, 0.4697684, 
    0.409826, 0.4315754, 0.4267073, 0.3482729, 0.3394794, 0.3256963, 
    0.3918956, 0.3345469, 0.3080357, 0.2971055, 0.3263948, 0.3819271, 
    0.3853222, 0.3612244, 0.3610695, 0.39477, 0.3681213,
  0.3394374, 0.2990223, 0.3316811, 0.2451084, 0.2640879, 0.2347373, 
    0.2726286, 0.2900016, 0.2591934, 0.2528074, 0.3171899, 0.3088763, 
    0.2415844, 0.3170684, 0.3425432, 0.405471, 0.3875949, 0.3814606, 
    0.3823912, 0.3499243, 0.3196777, 0.2766539, 0.251478, 0.247891, 
    0.1767396, 0.2249569, 0.3970111, 0.3511823, 0.3471731,
  0.2003365, 0.2021535, 0.1433398, 0.189702, 0.2019067, 0.1796419, 0.1958197, 
    0.2587042, 0.2282599, 0.1870585, 0.1844441, 0.1581367, 0.1097082, 
    0.1510385, 0.3041, 0.1947872, 0.2116012, 0.1960108, 0.2227567, 0.199692, 
    0.2438044, 0.2419401, 0.2098208, 0.3506488, 0.1646103, 0.1477522, 
    0.2151672, 0.2410223, 0.2432538,
  0.1925732, 0.05420316, 0.0250319, 0.1047334, 0.1145684, 0.151331, 0.180567, 
    0.1983333, 0.151288, 0.1028023, 0.006324015, 0.01147372, 0.02528749, 
    0.06327415, 0.1310766, 0.1353477, 0.111536, 0.09467432, 0.1436592, 
    0.2004251, 0.1600748, 0.1289861, 0.126386, 0.008161636, 0.1139828, 
    0.1399937, 0.1009577, 0.1377657, 0.1380538,
  0.2241319, -0.0001685142, 0.0006602102, 0.03509411, 0.09423237, 0.07052405, 
    0.1040533, 0.1625488, 0.1219815, 0.02367424, 8.876062e-05, 0.006327786, 
    0.1127112, 0.169489, 0.1496178, 0.08193235, 0.08220457, 0.1335075, 
    0.09108233, 0.1157037, 0.1494782, 0.1848492, 0.1970088, 5.786153e-06, 
    0.07640949, 0.04790365, 0.06186178, 0.1700951, 0.2174172,
  0.0487786, 6.333614e-07, 0.003900046, 0.1045566, 0.0638407, 0.05528792, 
    0.07071167, 0.08112517, 0.08175584, 0.06753717, 0.1164482, 0.09724002, 
    0.1354149, 0.05055531, 0.04649574, 0.06297529, 0.05904737, 0.04509804, 
    0.05337982, 0.07590421, 0.1201611, 0.1362454, -5.491883e-05, 0.07427032, 
    0.002877494, 6.544818e-06, 0.08773817, 0.06306776, 0.1640725,
  0.02958514, 0.1060328, 0.06803539, 0.01474216, 0.04069395, 0.05748372, 
    0.03436626, 0.03342252, 0.05700415, 0.1079925, 0.03800976, 0.02041812, 
    0.04553286, 0.03218573, 0.03098424, 0.0339218, 0.026427, 0.02344044, 
    0.01931735, 0.01724166, 0.02495243, 0.03200103, 0.002990012, 0.223982, 
    0.1577788, 0.03149699, 0.06033517, 0.03016858, 0.02494986,
  0.01265214, 0.002652589, 0.0001920512, -0.000176108, 3.73244e-05, 
    0.02247203, 0.05398222, 0.03119983, 0.008339603, 0.02951641, 0.0255513, 
    0.03781064, 0.0526009, 0.04421354, 0.04943129, 0.04968707, 0.06830113, 
    0.1101018, 0.1139265, 0.07294133, 0.07593833, 0.06638061, 0.1222432, 
    0.07438301, 0.04346187, 0.08720618, 0.1111945, 0.08145879, 0.02959457,
  1.151433e-06, 7.611625e-07, 4.789782e-08, 2.143296e-08, 3.130366e-08, 
    0.001722234, 0.03271591, 0.03436793, 0.1870753, 0.1054947, 0.05622425, 
    0.04898921, 0.03638571, 0.04229023, 0.04283943, 0.0428068, 0.06275232, 
    0.1257782, 0.08300672, 0.01804571, 0.003211503, 0.04585771, 0.02690732, 
    0.009367675, 0.04186799, 0.07371235, 0.1423903, 0.008275094, 0.0005033946,
  4.262067e-05, 1.596238e-06, -6.60431e-07, 6.202358e-07, 2.59766e-07, 
    3.24809e-08, 0.0002381711, 0.07514752, 0.3242494, 0.04444292, 0.1232914, 
    0.1833107, 0.08230165, 0.07154528, 0.1249345, 0.09567059, 0.1617614, 
    0.1241749, 0.2082206, 0.03199577, 1.071417e-06, 0.01496805, 0.03646125, 
    0.05152721, 0.07330512, 0.06517088, 0.1290503, 0.1335681, 0.002150608,
  0.01588931, 0.01222501, 0.005874654, 0.07389535, -0.0002471827, 
    -2.416775e-05, 0.02806995, 0.0003008795, 0.0002148874, 0.01985538, 
    0.2246432, 0.1303057, 0.1789377, 0.1989921, 0.2956348, 0.2912804, 
    0.2703214, 0.1867143, 0.1754297, 0.05669728, 0.003345254, 0.03214716, 
    0.04306781, 0.03779409, 0.1548523, 0.2441858, 0.2069997, 0.2168395, 
    0.08606062,
  0.1184684, 0.1689289, 0.1346362, 0.03315812, 0.01089337, 0.006951808, 
    0.02272883, 0.1359181, 0.1193816, 0.07365256, 0.1786654, 0.2096174, 
    0.1279, 0.2023232, 0.3758351, 0.4652181, 0.4343528, 0.331722, 0.2562709, 
    0.141459, 0.08823417, 0.04667009, 0.0760925, 0.1814245, 0.1538454, 
    0.230903, 0.2444588, 0.2627166, 0.1757233,
  0.1833016, 0.09906927, 0.06444291, 0.1092094, 0.203925, 0.1635697, 
    0.1019009, 0.1301768, 0.1651066, 0.1202386, 0.1882772, 0.2501583, 
    0.1951109, 0.2533484, 0.3155134, 0.2801076, 0.3190084, 0.4576413, 
    0.2087136, 0.0405664, 0.05124611, 0.07239374, 0.1089637, 0.1989865, 
    0.1869601, 0.1912395, 0.4460247, 0.3917037, 0.2652405,
  0.310666, 0.291186, 0.3265212, 0.218893, 0.3208241, 0.288202, 0.2442426, 
    0.148824, 0.1301133, 0.1557284, 0.1589486, 0.1589404, 0.1262544, 
    0.1632171, 0.1530888, 0.1666681, 0.2397112, 0.1683078, 0.09380059, 
    0.1889559, 0.239448, 0.2622643, 0.2508939, 0.2297932, 0.1178252, 
    0.302651, 0.2677603, 0.2211255, 0.3715897,
  0.321005, 0.3646842, 0.3036268, 0.2826752, 0.3404171, 0.3256177, 0.3354833, 
    0.2751664, 0.30669, 0.2907445, 0.2601817, 0.2312247, 0.2939284, 0.339421, 
    0.3933774, 0.4046303, 0.4255366, 0.4170989, 0.3571997, 0.4222604, 
    0.3880771, 0.3417492, 0.2782469, 0.2631598, 0.1956854, 0.2041741, 
    0.1717501, 0.2067949, 0.3129643,
  0.2031624, 0.2036224, 0.2040824, 0.2045424, 0.2050024, 0.2054624, 
    0.2059224, 0.2496105, 0.2583155, 0.2670205, 0.2757254, 0.2844304, 
    0.2931353, 0.3018403, 0.3041553, 0.3035341, 0.3029128, 0.3022915, 
    0.3016702, 0.3010489, 0.3004276, 0.2693865, 0.2608429, 0.2522992, 
    0.2437555, 0.2352118, 0.2266681, 0.2181244, 0.2027944,
  0.186087, 0.1837318, 0.1928406, 0.1255793, 0.08529739, 0.1818153, 
    0.1761079, 0.1464569, 0.02250666, 0.04507936, 0.07430319, 0.1356297, 
    0.2405232, 0.07574593, 0.2028795, 0.1867025, 0.1584861, 0.1878312, 
    0.2309851, 0.2488837, 0.437624, 0.4264065, 0.4072827, 0.2770367, 
    0.2530331, 0.2144777, 0.1800536, 0.1375654, 0.2394946,
  0.2344815, 0.2301316, 0.3008238, 0.1969505, 0.3642249, 0.3154255, 
    0.2614364, 0.4442332, 0.2901083, 0.2682937, 0.2426496, 0.2300839, 
    0.2743876, 0.270555, 0.3348853, 0.3824996, 0.41081, 0.4114219, 0.3712879, 
    0.3778283, 0.3730592, 0.3618437, 0.256433, 0.3574487, 0.2814119, 
    0.2522796, 0.3704797, 0.3644258, 0.2382312,
  0.4450542, 0.3785048, 0.3190389, 0.3177177, 0.3609883, 0.4124388, 
    0.4929899, 0.4215502, 0.4199562, 0.4643969, 0.4159398, 0.4485995, 
    0.4229321, 0.4118074, 0.4163652, 0.377697, 0.3975037, 0.4114634, 
    0.3657211, 0.3195144, 0.3131232, 0.2636991, 0.3007216, 0.3476515, 
    0.3682245, 0.4032736, 0.4041712, 0.4225177, 0.4125252,
  0.3370187, 0.314737, 0.315358, 0.258099, 0.2611874, 0.2323195, 0.285605, 
    0.246658, 0.2661003, 0.2620683, 0.2491068, 0.2591896, 0.2121475, 
    0.2875147, 0.3368241, 0.344217, 0.3939056, 0.4070375, 0.3649795, 
    0.3408304, 0.3068724, 0.2886504, 0.2295809, 0.2635654, 0.1584117, 
    0.2765109, 0.3703033, 0.2985365, 0.3016583,
  0.1704543, 0.1457692, 0.09454647, 0.137242, 0.1982873, 0.1505993, 
    0.2259314, 0.2528131, 0.2099931, 0.1515857, 0.1552037, 0.1180337, 
    0.06740646, 0.1287712, 0.3783015, 0.1395189, 0.1688302, 0.1973335, 
    0.2067591, 0.1526399, 0.1971807, 0.2033568, 0.2270772, 0.3894912, 
    0.1152416, 0.1194513, 0.1981658, 0.2069853, 0.2016407,
  0.1958786, 0.04928253, 0.02569233, 0.06348851, 0.1050217, 0.1290988, 
    0.1357916, 0.1524082, 0.09877881, 0.05541301, 0.002604175, 0.004355555, 
    0.02118652, 0.03427939, 0.07108, 0.09814581, 0.07219958, 0.06731347, 
    0.1101715, 0.1633171, 0.1446639, 0.1099341, 0.1419488, 0.01528371, 
    0.09041372, 0.09707889, 0.0830289, 0.09333991, 0.1086748,
  0.2033767, 0.007789381, 9.892264e-05, 0.07294103, 0.06202325, 0.03607655, 
    0.05169595, 0.1097172, 0.1374497, 0.01797192, 7.316627e-05, 0.004496156, 
    0.0345709, 0.1184967, 0.1383932, 0.08373987, 0.1132757, 0.1108703, 
    0.08563891, 0.08639851, 0.09275001, 0.1888766, 0.3515112, 0.0006254535, 
    0.1034397, 0.03812167, 0.05456632, 0.07656787, 0.1141553,
  0.2632903, 0.0001164973, 0.003610623, 0.0836058, 0.06009457, 0.05985161, 
    0.04883248, 0.1060749, 0.06726769, 0.06489407, 0.0892074, 0.08086964, 
    0.1364379, 0.06273656, 0.05668054, 0.07797378, 0.06022728, 0.08268306, 
    0.07142818, 0.06888232, 0.1244975, 0.3615345, 0.07715897, 0.06509517, 
    0.0006464004, -1.569939e-06, 0.05841913, 0.0663333, 0.3036404,
  0.0959072, 0.05889651, 0.03547458, 0.02243023, 0.06878063, 0.08794594, 
    0.1026345, 0.07229789, 0.03704134, 0.07900815, 0.07781295, 0.06216218, 
    0.08013877, 0.06648608, 0.04807194, 0.07516391, 0.05170373, 0.0490934, 
    0.04836415, 0.04134118, 0.04432424, 0.09257136, 0.01464735, 0.185138, 
    0.1116515, 0.0405609, 0.07219541, 0.0777384, 0.05511855,
  0.008094466, 0.002130053, 9.661892e-05, -0.0001376009, 8.620409e-07, 
    0.02496672, 0.05070145, 0.03488158, 0.004583021, 0.06709906, 0.02733967, 
    0.04720593, 0.05721393, 0.05096997, 0.05032311, 0.05548005, 0.06725152, 
    0.150565, 0.1581389, 0.1491084, 0.09571382, 0.08037437, 0.1283226, 
    0.08060215, 0.06130724, 0.09630908, 0.1484264, 0.09494164, 0.0165615,
  9.408018e-07, 6.943194e-07, 2.933142e-08, 2.173823e-08, 2.907155e-08, 
    0.01699241, 0.02429191, 0.02913046, 0.1623234, 0.1036641, 0.05843428, 
    0.06183888, 0.04048781, 0.04531121, 0.0549919, 0.05837248, 0.05579782, 
    0.1469405, 0.2646873, 0.03564021, 0.005752335, 0.05366147, 0.04159676, 
    0.01134969, 0.04615464, 0.06122338, 0.2087932, 0.01470546, 0.000203972,
  2.599023e-05, 8.981387e-07, -5.440104e-05, 5.604909e-07, 2.270865e-07, 
    2.944083e-08, 0.0001980403, 0.08520782, 0.3252419, 0.04692969, 0.1732514, 
    0.1957623, 0.1029638, 0.1153256, 0.1731851, 0.1164639, 0.1627432, 
    0.1850936, 0.3703045, 0.1296412, 7.159018e-07, 0.02547794, 0.02513046, 
    0.06620597, 0.07120014, 0.1370716, 0.1196572, 0.32807, 0.002547095,
  0.009928381, 0.01136496, 0.002992593, 0.08929653, -0.0002999751, 
    -7.091274e-06, 0.02394593, 3.028365e-05, 2.413983e-05, 0.01876818, 
    0.2249809, 0.1455848, 0.2647529, 0.3360629, 0.4014692, 0.3830284, 
    0.3150153, 0.3230328, 0.3165312, 0.05999842, 0.003698273, 0.04905272, 
    0.03591193, 0.03775999, 0.1858343, 0.2670338, 0.2980942, 0.3424233, 
    0.1120845,
  0.1038624, 0.1340163, 0.1214445, 0.02139041, 0.009534535, 0.004752954, 
    0.02234453, 0.1253034, 0.09750593, 0.05843607, 0.1510864, 0.1859133, 
    0.1748737, 0.2523799, 0.4141138, 0.5588726, 0.4906377, 0.3606571, 
    0.3179532, 0.1189771, 0.07757127, 0.0364252, 0.06891803, 0.1558721, 
    0.1416431, 0.2542388, 0.2710611, 0.2965978, 0.1850075,
  0.1529704, 0.07236551, 0.05075698, 0.08371069, 0.1808757, 0.1120549, 
    0.08537151, 0.08776011, 0.1402283, 0.09381132, 0.168431, 0.2358974, 
    0.1890489, 0.2476673, 0.3652073, 0.4049504, 0.2962604, 0.4278789, 
    0.1795591, 0.03048846, 0.03130205, 0.05867825, 0.1044989, 0.1796888, 
    0.2238878, 0.1754693, 0.4613044, 0.4334182, 0.2972124,
  0.3492722, 0.3176369, 0.3619075, 0.2906905, 0.3103686, 0.3272581, 
    0.2434113, 0.148467, 0.1184135, 0.1530807, 0.1337841, 0.1606018, 
    0.1262181, 0.1783891, 0.1842468, 0.2221162, 0.2862487, 0.1543183, 
    0.08218911, 0.2052563, 0.274235, 0.3642542, 0.2552374, 0.2959087, 
    0.1066121, 0.2807938, 0.2778076, 0.2549801, 0.4324665,
  0.3246173, 0.3907718, 0.3609409, 0.3801282, 0.4638688, 0.4065013, 
    0.4090127, 0.4176889, 0.3842889, 0.3498137, 0.2923563, 0.2897663, 
    0.3234462, 0.3847162, 0.4866787, 0.4444129, 0.4647708, 0.3914208, 
    0.3693486, 0.4538562, 0.4433004, 0.3721897, 0.2949319, 0.3148404, 
    0.2213238, 0.2258009, 0.1841255, 0.2301229, 0.3463756,
  0.2293641, 0.2295009, 0.2296378, 0.2297746, 0.2299114, 0.2300482, 0.230185, 
    0.2529372, 0.2608358, 0.2687344, 0.276633, 0.2845316, 0.2924301, 
    0.3003287, 0.3020762, 0.2994696, 0.2968631, 0.2942566, 0.2916501, 
    0.2890435, 0.286437, 0.2662929, 0.260864, 0.2554351, 0.2500063, 
    0.2445774, 0.2391485, 0.2337196, 0.2292547,
  0.1872083, 0.2110775, 0.2095165, 0.1545115, 0.1052858, 0.1955229, 
    0.2069643, 0.1775827, 0.01903127, 0.04434732, 0.08529958, 0.1443583, 
    0.2536536, 0.03638289, 0.2032638, 0.1920067, 0.1667173, 0.1916665, 
    0.2326606, 0.2457548, 0.4392479, 0.4133363, 0.3777765, 0.2526359, 
    0.2454372, 0.2165743, 0.1520698, 0.1418803, 0.2398885,
  0.2143646, 0.1825303, 0.2666759, 0.148437, 0.3268836, 0.3084071, 0.1754741, 
    0.4205186, 0.2788044, 0.2657008, 0.2482189, 0.2261018, 0.27101, 
    0.2555678, 0.3335582, 0.396912, 0.4373763, 0.4549836, 0.3845759, 
    0.3681403, 0.3939239, 0.3676118, 0.2593637, 0.3545671, 0.2947503, 
    0.2624871, 0.4706663, 0.4232674, 0.2608462,
  0.4412266, 0.329819, 0.2572284, 0.2677408, 0.3022293, 0.3169533, 0.4327511, 
    0.3162607, 0.3343869, 0.3840888, 0.3724347, 0.4063843, 0.38931, 
    0.3603926, 0.4364391, 0.3839648, 0.4121469, 0.3946378, 0.3603778, 
    0.2869211, 0.2897584, 0.2313041, 0.2679343, 0.294504, 0.3521545, 
    0.4265209, 0.4630135, 0.4231884, 0.4453866,
  0.3095002, 0.2918099, 0.2962895, 0.2547652, 0.2651513, 0.2605942, 
    0.2572048, 0.2275531, 0.2523776, 0.2481846, 0.2043431, 0.2251133, 
    0.1971011, 0.2353037, 0.2971767, 0.3009428, 0.3781056, 0.3889093, 
    0.351976, 0.3095316, 0.2757816, 0.2849006, 0.2101108, 0.2585336, 
    0.1297009, 0.2560629, 0.3425059, 0.2936136, 0.2851425,
  0.1428077, 0.1083894, 0.07573735, 0.09957756, 0.1571123, 0.1324485, 
    0.1952727, 0.2216791, 0.1950085, 0.1136723, 0.1354969, 0.09537312, 
    0.03880778, 0.09968276, 0.4317192, 0.1042333, 0.1375139, 0.1763131, 
    0.1685169, 0.1217123, 0.18039, 0.1476535, 0.1567246, 0.4159998, 
    0.07956198, 0.08449879, 0.1514919, 0.1736479, 0.1699433,
  0.0949219, 0.04811495, 0.01962922, 0.04367866, 0.09389237, 0.09824298, 
    0.06416088, 0.07175487, 0.05450375, 0.02203793, 0.001331661, 0.001488065, 
    0.01874575, 0.02231874, 0.04669595, 0.08010317, 0.05763435, 0.06126148, 
    0.0956526, 0.123761, 0.09561822, 0.06316434, 0.1084374, 0.02069774, 
    0.07200915, 0.06934484, 0.06893352, 0.05806673, 0.05850274,
  0.09338824, 0.0114406, -0.0001439566, 0.07496146, 0.02032898, 0.007834194, 
    0.01813088, 0.0624541, 0.0624412, 0.02104462, 3.807204e-05, 0.002216327, 
    0.01632648, 0.06467807, 0.1171734, 0.07412512, 0.09041804, 0.09736013, 
    0.03675813, 0.03519195, 0.03135432, 0.06645691, 0.2167227, 0.001987675, 
    0.1320558, 0.02581266, 0.02370794, 0.02371185, 0.05582627,
  0.3407067, 0.005758358, 0.001931947, 0.07174826, 0.04179727, 0.02523481, 
    0.0194859, 0.05058203, 0.02227832, 0.03903345, 0.04836761, 0.0297242, 
    0.1120052, 0.05572678, 0.03846464, 0.0374255, 0.0221898, 0.01960327, 
    0.0233549, 0.01187174, 0.0285246, 0.1357839, 0.3187024, 0.0149711, 
    7.174278e-05, 2.647469e-06, 0.005758351, 0.01823792, 0.1068876,
  0.2845843, 0.03227454, 0.01381008, 0.02293812, 0.05596528, 0.02486336, 
    0.03732451, 0.05811694, 0.02989842, 0.04664082, 0.06889541, 0.1553416, 
    0.05164869, 0.02492563, 0.0281739, 0.01973248, 0.04812137, 0.03933593, 
    0.03906749, 0.03593542, 0.09266448, 0.207717, 0.06570952, 0.1330517, 
    0.05859645, 0.03280254, 0.04336441, 0.05553187, 0.09524556,
  0.003652046, 0.001368649, 6.337568e-05, 0.0003894351, 1.641369e-06, 
    0.007303516, 0.04719694, 0.007187922, 0.0009144681, 0.02702961, 0.030411, 
    0.09830029, 0.04804143, 0.03276138, 0.03520446, 0.03689911, 0.04378822, 
    0.09439235, 0.09850709, 0.1728922, 0.119919, 0.08224173, 0.1483116, 
    0.06164842, 0.05373637, 0.06613591, 0.1523555, 0.233525, 0.009288074,
  8.115811e-07, 6.385557e-07, 2.357209e-08, 1.543123e-08, 2.79132e-08, 
    0.1692015, 0.02474564, 0.02805895, 0.140001, 0.1010209, 0.09118444, 
    0.02984121, 0.01131459, 0.0161207, 0.02800865, 0.0583299, 0.0157321, 
    0.06590317, 0.3345006, 0.2996814, 0.03159418, 0.06538555, 0.02025223, 
    0.001860102, 0.01402801, 0.01342519, 0.07066333, 0.1690386, 0.0001048664,
  3.190446e-05, -2.382236e-06, -8.129101e-05, 4.984084e-07, 2.040295e-07, 
    2.747757e-08, -0.0001507331, 0.08833945, 0.3092909, 0.05151299, 
    0.1805216, 0.234443, 0.1119023, 0.1508954, 0.2484798, 0.1464574, 
    0.1131694, 0.111613, 0.2134369, 0.2815177, 4.496055e-07, 0.02419204, 
    0.02171461, 0.1106328, 0.07348217, 0.09091662, 0.05666856, 0.1753286, 
    0.004902353,
  0.009875213, 0.01211887, 0.001989009, 0.1111911, 0.0003468901, 
    -2.055619e-06, 0.02051058, -4.036727e-05, -5.922722e-06, 0.01677126, 
    0.218765, 0.1858045, 0.3533123, 0.4891083, 0.4194607, 0.4238486, 
    0.3772414, 0.4871168, 0.4293646, 0.05393182, 0.003853683, 0.05685995, 
    0.02825644, 0.02950844, 0.2398814, 0.2909284, 0.2940474, 0.3668967, 
    0.1462266,
  0.09452831, 0.1076065, 0.1038916, 0.0163273, 0.009749431, 0.003343282, 
    0.01716362, 0.1240854, 0.08229791, 0.05689104, 0.1340153, 0.1598154, 
    0.3378048, 0.3666132, 0.5163578, 0.6223532, 0.5107781, 0.4112264, 0.3831, 
    0.107811, 0.07248294, 0.03239518, 0.05193046, 0.1433315, 0.1321712, 
    0.2629602, 0.2864258, 0.3487651, 0.1690597,
  0.1443823, 0.05005425, 0.04120405, 0.06937575, 0.1451198, 0.07623319, 
    0.06684737, 0.06348734, 0.1209112, 0.07708725, 0.1544784, 0.2277722, 
    0.1791712, 0.2320359, 0.3927275, 0.4618121, 0.2761577, 0.4089341, 
    0.1751584, 0.02125536, 0.02116946, 0.04726772, 0.09212092, 0.1796567, 
    0.2857578, 0.1920442, 0.4912903, 0.4011467, 0.2427166,
  0.4306831, 0.3612118, 0.3207586, 0.4276203, 0.3027166, 0.3524965, 
    0.2530301, 0.1441644, 0.103428, 0.1225386, 0.1202063, 0.1339131, 
    0.09985629, 0.1740579, 0.2078868, 0.2818192, 0.2419145, 0.1607461, 
    0.1449792, 0.1833795, 0.3330975, 0.4224748, 0.1981712, 0.3250291, 
    0.1135705, 0.2738245, 0.268436, 0.2439449, 0.456103,
  0.3971133, 0.4234252, 0.3951856, 0.5332549, 0.6224815, 0.5529883, 0.501097, 
    0.5102348, 0.4488781, 0.417457, 0.323691, 0.3855898, 0.4333472, 
    0.5280954, 0.5194553, 0.4545692, 0.4434281, 0.350574, 0.3827162, 
    0.482825, 0.4308975, 0.3596256, 0.2867432, 0.3264246, 0.2583577, 
    0.1924768, 0.1709816, 0.2568299, 0.4883512,
  0.2204048, 0.2209765, 0.2215482, 0.2221198, 0.2226915, 0.2232632, 
    0.2238349, 0.2468678, 0.2551709, 0.2634741, 0.2717772, 0.2800804, 
    0.2883836, 0.2966867, 0.2890561, 0.2849194, 0.2807826, 0.2766459, 
    0.2725092, 0.2683724, 0.2642357, 0.2599997, 0.2552616, 0.2505235, 
    0.2457854, 0.2410473, 0.2363091, 0.231571, 0.2199475,
  0.1964178, 0.2405339, 0.195101, 0.1621264, 0.1170409, 0.1846446, 0.2179714, 
    0.1847302, 0.01817356, 0.04448907, 0.09346567, 0.1206463, 0.2591142, 
    0.01865682, 0.204584, 0.2108084, 0.2026991, 0.1924963, 0.2319511, 
    0.2630532, 0.4449276, 0.4086088, 0.3479742, 0.2362149, 0.2382991, 
    0.23762, 0.1443955, 0.1705912, 0.2342396,
  0.2001368, 0.151701, 0.2321628, 0.1071356, 0.2677943, 0.2964597, 0.1073985, 
    0.398409, 0.2677816, 0.2534686, 0.2467571, 0.2333903, 0.2380376, 
    0.2330652, 0.3462091, 0.3979631, 0.4329364, 0.4670916, 0.3607255, 
    0.3745488, 0.400435, 0.3815535, 0.2737026, 0.3647448, 0.3083186, 
    0.3172194, 0.5043018, 0.4637677, 0.2775534,
  0.4404792, 0.2804722, 0.1868796, 0.2208421, 0.2846729, 0.2565239, 
    0.3633927, 0.2580856, 0.2588884, 0.3137603, 0.3169799, 0.3583247, 
    0.3665461, 0.3713271, 0.3964268, 0.3640747, 0.3971664, 0.3843608, 
    0.3415965, 0.2675584, 0.2385375, 0.1994879, 0.2426779, 0.2475553, 
    0.3263602, 0.4315215, 0.4746612, 0.4294572, 0.4467663,
  0.2728249, 0.2543713, 0.2842311, 0.237338, 0.2477151, 0.2594621, 0.2572907, 
    0.2036952, 0.2348911, 0.2330816, 0.1760964, 0.1992013, 0.1700383, 
    0.22056, 0.2787863, 0.2605145, 0.3311811, 0.3565505, 0.3503426, 
    0.2810296, 0.2377385, 0.2324412, 0.1691989, 0.2413419, 0.09136276, 
    0.1922763, 0.3055899, 0.2912561, 0.2696902,
  0.126162, 0.07470843, 0.057276, 0.06457777, 0.1094422, 0.1028581, 
    0.1516502, 0.1838523, 0.1550536, 0.07947443, 0.1007188, 0.06458414, 
    0.01921856, 0.07504995, 0.3996954, 0.08607017, 0.1220667, 0.1427148, 
    0.1318379, 0.1082076, 0.1598309, 0.1195624, 0.1123753, 0.41606, 
    0.06238145, 0.06421649, 0.1285023, 0.1531484, 0.1322901,
  0.0443462, 0.05692683, 0.01439304, 0.0329113, 0.05533498, 0.05319829, 
    0.02768985, 0.04144892, 0.03760193, 0.01325114, 0.001329881, 
    0.0002853074, 0.02037362, 0.01350715, 0.03543893, 0.07305133, 0.04759786, 
    0.05494965, 0.06831388, 0.08704659, 0.06998818, 0.02826861, 0.05702535, 
    0.03015145, 0.06396003, 0.04926737, 0.04596209, 0.03205708, 0.03525261,
  0.06333267, 0.01401142, -3.218678e-05, 0.02606916, 0.001439654, 
    0.001343473, 0.003432727, 0.03823572, 0.02738297, 0.004560424, 
    -2.654608e-05, 0.0008287643, 0.009340469, 0.03810926, 0.07311878, 
    0.03029003, 0.04583856, 0.05660773, 0.01608702, 0.02336543, 0.01070182, 
    0.02277162, 0.07252401, 0.01334067, 0.1134157, 0.0283806, 0.005096265, 
    0.005543463, 0.01730208,
  0.152653, 0.01540946, 0.002075227, 0.08421907, 0.02045672, 0.006949376, 
    0.005062357, 0.01118364, 0.007823418, 0.007733232, 0.02748803, 
    0.01027098, 0.08725062, 0.01998567, 0.0139282, 0.01764542, 0.005030205, 
    0.003482975, 0.002959555, 0.001921587, 0.007257598, 0.04011366, 
    0.2707856, 0.00276807, 8.321074e-06, 2.39598e-06, -0.002933802, 
    0.004600234, 0.03867115,
  0.2073293, 0.02036729, 0.006922557, 0.01995766, 0.02258316, 0.003676792, 
    0.005546846, 0.01012528, 0.03616832, 0.02707797, 0.01096467, 0.02832465, 
    0.03719334, 0.0105441, 0.01225619, 0.004459105, 0.01564661, 0.009572409, 
    0.01262142, 0.01334991, 0.04654421, 0.1261609, 0.4255518, 0.09497499, 
    0.02974303, 0.01096419, 0.02360864, 0.01136979, 0.04527763,
  0.002131559, 0.00060215, 3.196808e-05, 0.001445818, -8.349778e-06, 
    0.0005527233, 0.04806869, 0.0006737888, -0.000835084, 0.006079944, 
    0.007552328, 0.0307449, 0.0252455, 0.01388555, 0.01438645, 0.01334402, 
    0.01971355, 0.04328925, 0.05483989, 0.05234316, 0.04388288, 0.05519844, 
    0.1423661, 0.04791779, 0.0132933, 0.03206366, 0.06881607, 0.1727081, 
    0.005574404,
  7.348808e-07, 5.944094e-07, 2.185095e-08, 1.377364e-08, 2.725766e-08, 
    0.1195047, 0.0181966, 0.02116466, 0.1314845, 0.08030592, 0.03907702, 
    0.01572504, 0.001337633, 0.002238058, 0.003981228, 0.008498433, 
    0.008122195, 0.02598256, 0.1623579, 0.2792456, 0.07950812, 0.05089213, 
    0.002392935, -0.0004433439, 0.001520585, 0.001140633, 0.02196334, 
    0.07458529, 2.823208e-05,
  2.388466e-05, -6.816229e-05, 7.427278e-05, 4.095835e-07, 1.894741e-07, 
    2.623481e-08, -0.0004501493, 0.08650999, 0.3025956, 0.04519916, 
    0.1781406, 0.2882075, 0.1958527, 0.1539718, 0.1643801, 0.08098264, 
    0.07576829, 0.05216489, 0.08446345, 0.2491616, 3.721814e-07, 0.02093387, 
    0.02372302, 0.05666366, 0.05207883, 0.04033279, 0.03180854, 0.06894431, 
    0.009904681,
  0.007609141, 0.01333991, 0.001232602, 0.1364433, 8.536356e-05, 
    -3.353895e-07, 0.01849539, -3.603219e-05, -3.472718e-05, 0.01390897, 
    0.2012546, 0.2118707, 0.3703581, 0.4777792, 0.4253421, 0.3592912, 
    0.4652069, 0.4867997, 0.4082727, 0.05070883, 0.003495775, 0.05505484, 
    0.0270048, 0.05479192, 0.2446204, 0.3143317, 0.2474121, 0.2675624, 
    0.1557302,
  0.07980078, 0.09286644, 0.0831499, 0.01090334, 0.005600959, 0.001838683, 
    0.01229751, 0.1210902, 0.07088916, 0.05162332, 0.1294464, 0.1645141, 
    0.4911617, 0.4664265, 0.5633639, 0.6113706, 0.5341434, 0.4903489, 
    0.3853113, 0.1022518, 0.06315724, 0.02203167, 0.04445311, 0.1336467, 
    0.127158, 0.2712349, 0.3233504, 0.3516261, 0.1541631,
  0.1780808, 0.03875171, 0.03276027, 0.06618346, 0.1182565, 0.06270352, 
    0.05143847, 0.04789935, 0.10281, 0.06862243, 0.1481083, 0.2215228, 
    0.169766, 0.2230086, 0.4064125, 0.4247568, 0.2574905, 0.3901107, 
    0.1661543, 0.0168876, 0.01260614, 0.04467967, 0.101281, 0.1586707, 
    0.2958218, 0.182671, 0.4584862, 0.3497429, 0.2085257,
  0.5065663, 0.3758985, 0.2732035, 0.4582064, 0.2761698, 0.3123763, 
    0.2260615, 0.12786, 0.07823573, 0.09477291, 0.0996179, 0.09354636, 
    0.06430764, 0.2017725, 0.2404144, 0.3046935, 0.2021968, 0.1616979, 
    0.1939831, 0.2063644, 0.2815061, 0.3963176, 0.1473668, 0.3122513, 
    0.2658419, 0.2362355, 0.2089095, 0.2314799, 0.5197221,
  0.5743877, 0.4489464, 0.4115858, 0.5265635, 0.582142, 0.5552349, 0.4985339, 
    0.4538673, 0.3843246, 0.387138, 0.3779694, 0.4464433, 0.474283, 
    0.5199554, 0.5365005, 0.5144385, 0.4688405, 0.4254467, 0.4295818, 
    0.4773951, 0.4095707, 0.3571805, 0.3059573, 0.3651946, 0.2751584, 
    0.1753194, 0.1562469, 0.3423693, 0.5790804,
  0.1448265, 0.1426884, 0.1405503, 0.1384122, 0.1362741, 0.134136, 0.1319979, 
    0.1352451, 0.1477369, 0.1602287, 0.1727206, 0.1852124, 0.1977042, 
    0.210196, 0.2411707, 0.2375199, 0.2338692, 0.2302184, 0.2265676, 
    0.2229168, 0.2192661, 0.2071156, 0.2004126, 0.1937097, 0.1870068, 
    0.1803038, 0.1736009, 0.1668979, 0.146537,
  0.1996718, 0.2506925, 0.1452294, 0.1426634, 0.09990519, 0.1487875, 
    0.2039436, 0.1674874, 0.008292524, 0.00598809, 0.03451353, 0.1146392, 
    0.2592866, 0.006080892, 0.2211622, 0.2636903, 0.2941202, 0.2327538, 
    0.2345079, 0.2959825, 0.4436722, 0.4314774, 0.298871, 0.1849851, 
    0.2186381, 0.2406078, 0.1752295, 0.1855665, 0.2112621,
  0.1953638, 0.1291667, 0.195245, 0.07136355, 0.2048109, 0.2747698, 
    0.07078717, 0.3470705, 0.253036, 0.2315641, 0.2355531, 0.2323147, 
    0.1936058, 0.1976951, 0.3655636, 0.4238964, 0.4341792, 0.4454531, 
    0.3448201, 0.3526266, 0.3793253, 0.3800089, 0.2702008, 0.355296, 
    0.2985033, 0.3822629, 0.5572173, 0.4874802, 0.2946275,
  0.403029, 0.2163656, 0.1392529, 0.1728806, 0.2368817, 0.2109467, 0.304911, 
    0.211851, 0.2159846, 0.2594356, 0.25675, 0.289919, 0.3421296, 0.3515477, 
    0.3204969, 0.3395061, 0.3831917, 0.3443372, 0.3123449, 0.2348167, 
    0.1964554, 0.1747567, 0.2211918, 0.2067007, 0.2815257, 0.4198067, 
    0.4418635, 0.3955721, 0.4115174,
  0.2368656, 0.2136456, 0.2579701, 0.2166993, 0.223753, 0.2516012, 0.2409783, 
    0.1692868, 0.2097951, 0.2000397, 0.1468893, 0.1706506, 0.1278506, 
    0.1910363, 0.25642, 0.2302357, 0.2717594, 0.3215091, 0.3265141, 
    0.2621962, 0.2067644, 0.2090635, 0.1179333, 0.2066405, 0.05965816, 
    0.1320563, 0.2525314, 0.2666903, 0.2465701,
  0.09386659, 0.04775476, 0.03852067, 0.03919315, 0.0690636, 0.07444577, 
    0.1137281, 0.1409559, 0.1106964, 0.05094204, 0.07325979, 0.03860349, 
    0.008731865, 0.05160738, 0.3463818, 0.07360164, 0.1052698, 0.1133735, 
    0.101533, 0.1033377, 0.1236278, 0.09044078, 0.08031195, 0.4071816, 
    0.04553784, 0.04607104, 0.1001219, 0.116796, 0.1018709,
  0.02083353, 0.02929845, 0.01423485, 0.01975096, 0.02719637, 0.02835019, 
    0.01445231, 0.03034532, 0.02781487, 0.004639582, 0.0005828447, 
    0.0001865567, 0.02670602, 0.007736902, 0.02388053, 0.057969, 0.03850543, 
    0.04435362, 0.04093382, 0.05392286, 0.0363983, 0.01164623, 0.02640347, 
    0.02999153, 0.05429087, 0.02440276, 0.02621443, 0.01474555, 0.01974234,
  0.03398736, 0.01467405, 9.120551e-05, 0.009494059, -0.002497375, 
    0.0006002667, 0.001105371, 0.02641381, 0.0143319, 0.001250896, 
    -5.748984e-05, 0.0002716436, 0.00640268, 0.02201891, 0.03602558, 
    0.0106161, 0.01610386, 0.02392866, 0.006732144, 0.01662426, 0.004095046, 
    0.008701155, 0.02843773, 0.02420294, 0.08661023, 0.04150177, 0.001546405, 
    0.002433861, 0.006018818,
  0.0684756, 0.006078518, 0.0009972339, 0.0825307, 0.008685028, 0.001434607, 
    0.0008956699, 0.003020741, 0.003099954, 0.0004103866, 0.01577175, 
    0.004765634, 0.05175446, 0.005168396, 0.002912581, 0.005503382, 
    0.001121837, 0.0008145801, 0.0008670558, 0.0008329983, 0.003231438, 
    0.01475777, 0.1213957, 0.0008928566, -6.073086e-06, 2.383723e-06, 
    -0.0008553822, 0.001707585, 0.0167928,
  0.06669857, 0.01357167, 0.00548694, 0.01307893, 0.003809027, 0.001021534, 
    0.001464274, 0.003904215, 0.0377859, 0.0157113, 0.001802183, 0.007622612, 
    0.02313441, 0.003138147, 0.004739851, 0.0006295043, 0.005680777, 
    0.001230213, 0.0019961, 0.001325766, 0.007480091, 0.03068985, 0.1881269, 
    0.08300191, 0.02635887, 0.004300554, 0.015029, 0.001710167, 0.008342765,
  0.00157178, 0.0004808218, 9.915036e-06, 0.001751376, 4.688858e-06, 
    1.851369e-05, 0.03279053, 8.942604e-05, -0.0005865679, 0.001794834, 
    0.002760252, 0.01418262, 0.01301068, 0.005688542, 0.004417209, 
    0.003315005, 0.008323225, 0.01617941, 0.02943028, 0.0179147, 0.01351842, 
    0.02180632, 0.1612538, 0.03982633, 0.003286709, 0.01091647, 0.01900014, 
    0.06398164, 0.004408899,
  6.879863e-07, 5.534716e-07, 2.147417e-08, 1.209509e-08, 2.6425e-08, 
    0.03987246, 0.009690481, 0.01095459, 0.1166797, 0.03714455, 0.01723576, 
    0.009582398, 0.0001232099, 0.0001892593, 0.0006599522, 0.002098397, 
    0.004438612, 0.01008306, 0.07303604, 0.1455119, 0.07080314, 0.04331835, 
    0.000591868, -0.0009058563, 0.0001435248, 0.0002308636, 0.008265289, 
    0.03001571, 7.958923e-06,
  1.291269e-05, -3.743015e-05, -4.051169e-05, 1.434441e-08, 1.791029e-07, 
    2.543693e-08, -0.0004622716, 0.07731147, 0.2894174, 0.03619975, 
    0.1997935, 0.2736917, 0.1870903, 0.08490495, 0.08541851, 0.0385158, 
    0.04955498, 0.02081917, 0.0382318, 0.151423, 3.471781e-07, 0.01540459, 
    0.02522777, 0.02687984, 0.02818294, 0.02171552, 0.01016246, 0.02342816, 
    0.01876038,
  0.006192601, 0.007513217, 0.0003594512, 0.1420616, -2.288482e-05, 
    1.051717e-07, 0.01650187, -6.138758e-05, -5.375201e-05, 0.0109031, 
    0.1922706, 0.2039307, 0.3391392, 0.4254182, 0.3718725, 0.3024882, 
    0.4164622, 0.322557, 0.271811, 0.04572559, 0.003517456, 0.04889117, 
    0.02129347, 0.06010067, 0.1708069, 0.2510583, 0.1767259, 0.1708508, 
    0.1529802,
  0.09174879, 0.08363553, 0.06128699, 0.005774301, 0.002220414, 0.0008308017, 
    0.009636935, 0.1167414, 0.06256308, 0.05108386, 0.1281576, 0.1618989, 
    0.5739975, 0.5110174, 0.5576299, 0.5314896, 0.528035, 0.5264883, 
    0.3396323, 0.09701066, 0.0471065, 0.01209926, 0.04551718, 0.1207932, 
    0.1270852, 0.2779827, 0.3256107, 0.3037232, 0.1622605,
  0.1893398, 0.02865905, 0.02595983, 0.05846807, 0.09850841, 0.05327193, 
    0.04250406, 0.03767841, 0.08905005, 0.06335516, 0.1394931, 0.2011195, 
    0.1494088, 0.2155055, 0.4145698, 0.4226491, 0.23489, 0.3520754, 
    0.1448807, 0.01137036, 0.009638863, 0.04597011, 0.1015086, 0.1271779, 
    0.2967534, 0.160656, 0.3866521, 0.3072715, 0.1764675,
  0.5334518, 0.341872, 0.2267382, 0.3898956, 0.2826244, 0.3029618, 0.1812114, 
    0.1119526, 0.05641665, 0.07607223, 0.08150987, 0.06592707, 0.04355547, 
    0.2097112, 0.2478999, 0.2853519, 0.1615332, 0.1714421, 0.212413, 
    0.1956421, 0.2120802, 0.3294397, 0.1118612, 0.2794381, 0.3166059, 
    0.2060152, 0.1621613, 0.2236514, 0.5719494,
  0.6304767, 0.4017226, 0.372167, 0.459232, 0.5217249, 0.5034855, 0.4777702, 
    0.4579702, 0.3600436, 0.4081027, 0.4204795, 0.4133648, 0.4366206, 
    0.4547481, 0.5069945, 0.4897301, 0.4330645, 0.4420978, 0.4422775, 
    0.4083652, 0.3703081, 0.3163918, 0.2447828, 0.3611401, 0.2414836, 
    0.1404066, 0.1448698, 0.4131806, 0.5952799,
  0.05159587, 0.04950647, 0.04741706, 0.04532766, 0.04323824, 0.04114884, 
    0.03905943, 0.04251825, 0.05382301, 0.06512778, 0.07643253, 0.08773729, 
    0.09904206, 0.1103468, 0.1344336, 0.1335112, 0.1325889, 0.1316665, 
    0.1307441, 0.1298218, 0.1288994, 0.1222483, 0.1139553, 0.1056623, 
    0.09736931, 0.08907631, 0.08078332, 0.07249033, 0.0532674,
  0.2002286, 0.2024932, 0.1030594, 0.08018649, 0.05976154, 0.09668175, 
    0.1451145, 0.1296429, 0.01187103, 0.005260209, 0.004277024, 0.06980506, 
    0.2504118, 0.0002125569, 0.2720828, 0.3042109, 0.3789022, 0.262859, 
    0.2112928, 0.3113349, 0.466538, 0.4615952, 0.2161707, 0.1400232, 
    0.1961745, 0.287725, 0.2035817, 0.1768955, 0.2032003,
  0.1995018, 0.1169055, 0.1688207, 0.04228005, 0.1530347, 0.2506688, 
    0.04474461, 0.2774983, 0.2316133, 0.1981838, 0.216243, 0.2302341, 
    0.1535487, 0.1655783, 0.3840595, 0.4000316, 0.4121087, 0.4344535, 
    0.3140591, 0.3138459, 0.371646, 0.3496878, 0.2790894, 0.3415956, 
    0.2884046, 0.4082936, 0.5514072, 0.4952655, 0.2986901,
  0.3545823, 0.1546985, 0.1014357, 0.1261357, 0.1857904, 0.1563354, 
    0.2439748, 0.1686709, 0.1661417, 0.1964841, 0.1936902, 0.2276783, 
    0.2946255, 0.2923872, 0.2724486, 0.2943772, 0.342918, 0.2946432, 
    0.2694283, 0.1934331, 0.1550756, 0.1400688, 0.1916858, 0.1643953, 
    0.2346648, 0.3820306, 0.3956499, 0.3402935, 0.3605752,
  0.1929518, 0.165381, 0.2135168, 0.1786034, 0.1909772, 0.2174284, 0.2190881, 
    0.1348604, 0.1694067, 0.165523, 0.1112318, 0.1284913, 0.08743153, 
    0.1412325, 0.2137629, 0.1815086, 0.2013656, 0.2757004, 0.2726863, 
    0.2195088, 0.1644256, 0.1697902, 0.07940406, 0.16912, 0.0402301, 
    0.08666757, 0.2045613, 0.2289971, 0.2007402,
  0.06427565, 0.02702564, 0.02540278, 0.02255438, 0.04111354, 0.04611175, 
    0.07529959, 0.104721, 0.07242897, 0.03077818, 0.04685606, 0.02349539, 
    0.00377253, 0.0335453, 0.2857355, 0.06049897, 0.08028521, 0.08355336, 
    0.07534853, 0.08804846, 0.09091386, 0.06064752, 0.05746597, 0.3848694, 
    0.03010198, 0.03407147, 0.07319485, 0.07643334, 0.08001179,
  0.009998694, 0.01705766, 0.01245754, 0.01046645, 0.01209221, 0.01460704, 
    0.00770695, 0.02295357, 0.01937478, 0.002355526, 0.0002046436, 
    0.0001844852, 0.0277376, 0.004901593, 0.01635516, 0.04356922, 0.03063195, 
    0.0300148, 0.02637886, 0.02785737, 0.01757664, 0.004425993, 0.01198488, 
    0.01565652, 0.03858095, 0.01202541, 0.01187374, 0.006471537, 0.01005464,
  0.02095405, 0.01638852, 2.466035e-05, 0.005236565, -0.002354528, 
    0.0003418582, 0.0005485588, 0.01478423, 0.007383372, 0.0006260167, 
    -6.784376e-05, 0.000116741, 0.004264333, 0.009379266, 0.01434744, 
    0.004158913, 0.007290914, 0.01104684, 0.002958131, 0.008735285, 
    0.001512319, 0.004735436, 0.01502576, 0.01499085, 0.07073206, 0.05196102, 
    0.0007861426, 0.001242658, 0.003031057,
  0.03873579, 0.002310046, 0.00041761, 0.06654251, 0.003206992, 0.0004128342, 
    0.0002780464, 0.001287034, 0.0009725206, -0.0002046303, 0.009684731, 
    0.001970287, 0.02562558, 0.001192906, 0.001287372, 0.001677769, 
    0.0002915782, 0.0004260105, 0.0004452233, 0.0004734461, 0.001857593, 
    0.007645567, 0.06897814, 0.0006015393, -2.023901e-05, -4.352207e-07, 
    -0.0006051577, 0.0008471789, 0.009141795,
  0.03197736, 0.01334534, 0.004900947, 0.007970991, 0.0005739827, 
    0.0005601393, 0.0007423381, 0.001960673, 0.03568462, 0.01343685, 
    0.0006820272, 0.003798741, 0.01283165, 0.001349329, 0.001510318, 
    0.000239593, 0.002104887, 0.000512165, 0.0008407381, 0.0003610958, 
    0.002731089, 0.0115547, 0.08569683, 0.08206303, 0.02992221, 0.001610635, 
    0.01166646, 0.0007709675, 0.002792173,
  0.001087626, 0.00040226, 2.331595e-06, 0.001230841, 1.116185e-07, 
    4.98507e-06, 0.01582523, 2.968509e-05, -0.000255084, 0.000888648, 
    0.001153744, 0.007057416, 0.006734475, 0.003207985, 0.001383888, 
    0.0007786876, 0.002880893, 0.005300395, 0.01407649, 0.009387866, 
    0.00604621, 0.01050843, 0.1486298, 0.03807323, 0.001111478, 0.003712778, 
    0.007456469, 0.03165041, 0.006739728,
  6.543138e-07, 5.237954e-07, 2.152201e-08, 4.193174e-09, 2.6175e-08, 
    0.01776322, 0.003012308, 0.002310438, 0.09201054, 0.01324682, 0.00623773, 
    0.006069001, 4.84265e-05, 4.166154e-05, 0.0001884368, 0.001027794, 
    0.002434838, 0.004830604, 0.03775463, 0.07932277, 0.06876901, 0.03615179, 
    0.0002748235, -0.0008840229, 3.934496e-05, 0.0001167144, 0.004011457, 
    0.01497412, 2.117962e-06,
  5.790963e-06, -1.168921e-05, 2.315008e-05, -1.095774e-06, 1.679907e-07, 
    2.487161e-08, -0.0004249999, 0.06908636, 0.2690715, 0.02614671, 
    0.1855051, 0.1816562, 0.1250852, 0.02807411, 0.04878773, 0.01712999, 
    0.02417309, 0.009189129, 0.02218134, 0.09329672, 3.184207e-07, 
    0.01085616, 0.02121228, 0.01433974, 0.01544274, 0.00887587, 0.003773252, 
    0.01203501, 0.01798073,
  0.004826299, 0.002882471, -3.753869e-05, 0.1404251, -9.60121e-05, 
    2.870918e-07, 0.01361007, -5.082997e-05, -4.728249e-05, 0.008096172, 
    0.1781812, 0.2085148, 0.3144751, 0.3579357, 0.3227484, 0.2593425, 
    0.3500939, 0.1980808, 0.178465, 0.03854708, 0.003992275, 0.03724375, 
    0.01547636, 0.05421243, 0.1233238, 0.1779077, 0.120128, 0.1104641, 
    0.1089421,
  0.0866008, 0.07794214, 0.04007529, 0.003645656, 0.0009856077, 0.0001149406, 
    0.007406229, 0.1065728, 0.05246474, 0.0464372, 0.1266278, 0.1485508, 
    0.5804456, 0.4879901, 0.499402, 0.4388623, 0.4482178, 0.4716325, 
    0.2807218, 0.08853487, 0.03527423, 0.006405622, 0.03942608, 0.1054406, 
    0.1285301, 0.2914721, 0.2943254, 0.2448632, 0.1503994,
  0.1827071, 0.02238376, 0.01856859, 0.04545118, 0.07673453, 0.04241642, 
    0.03423891, 0.0281552, 0.07608641, 0.05561381, 0.1308746, 0.167284, 
    0.1328855, 0.1945658, 0.4015345, 0.4091176, 0.2074794, 0.3034901, 
    0.1131208, 0.009250669, 0.007200901, 0.03865782, 0.09981717, 0.1006599, 
    0.2670111, 0.1404341, 0.3059713, 0.242609, 0.1717848,
  0.5251313, 0.303094, 0.1881294, 0.3321705, 0.248683, 0.3002865, 0.1865822, 
    0.08742719, 0.04216132, 0.059787, 0.06578111, 0.05064769, 0.02948041, 
    0.1855314, 0.2266148, 0.2785708, 0.1110558, 0.1488004, 0.2167534, 
    0.1524992, 0.1637405, 0.2737556, 0.08401895, 0.2545912, 0.3482175, 
    0.1772636, 0.1237127, 0.2259855, 0.5928895,
  0.5767016, 0.3345184, 0.2960731, 0.4154871, 0.4734629, 0.4909334, 
    0.4639511, 0.438167, 0.3480734, 0.3796732, 0.3649985, 0.3511827, 
    0.3700159, 0.4211943, 0.4615979, 0.4328146, 0.3937874, 0.4006068, 
    0.3826366, 0.3028522, 0.3259257, 0.2551057, 0.1819017, 0.307421, 
    0.2102102, 0.1076785, 0.1248116, 0.4084972, 0.552393,
  0.01187622, 0.01048053, 0.009084838, 0.007689146, 0.006293454, 0.004897761, 
    0.003502069, -0.002246648, 0.005205844, 0.01265834, 0.02011083, 
    0.02756332, 0.03501581, 0.04246831, 0.06166835, 0.06190859, 0.06214882, 
    0.06238906, 0.0626293, 0.06286953, 0.06310977, 0.05183589, 0.04553885, 
    0.03924181, 0.03294478, 0.02664774, 0.0203507, 0.01405367, 0.01299278,
  0.205489, 0.1243365, 0.05364404, 0.01979239, 0.01136744, 0.04324077, 
    0.0735834, 0.07459228, 0.01992681, 0.006938693, 0.01295394, 0.02975417, 
    0.1586848, -0.0009808999, 0.2980961, 0.3637823, 0.4061413, 0.2827476, 
    0.1816911, 0.3218268, 0.4896896, 0.4952596, 0.1610078, 0.1036859, 
    0.183339, 0.3720261, 0.2200493, 0.1550592, 0.2254129,
  0.2133633, 0.1012634, 0.1387348, 0.02856058, 0.118285, 0.22409, 0.03468746, 
    0.2060164, 0.2025888, 0.1720448, 0.2029455, 0.2247105, 0.1231134, 
    0.147737, 0.387649, 0.38498, 0.3742959, 0.3954132, 0.2649817, 0.2631216, 
    0.3279051, 0.3022555, 0.2621129, 0.3319862, 0.2737694, 0.4088261, 
    0.5066426, 0.4705487, 0.2853871,
  0.2891974, 0.1068841, 0.07345232, 0.09085843, 0.1372619, 0.1108229, 
    0.187957, 0.1304432, 0.1253668, 0.1396845, 0.1355915, 0.1768241, 
    0.2283173, 0.2247086, 0.2083005, 0.2303256, 0.2835565, 0.2350673, 
    0.2226264, 0.145618, 0.1181098, 0.09890492, 0.1501092, 0.1229672, 
    0.1888212, 0.3214078, 0.3204162, 0.280413, 0.2926607,
  0.1531022, 0.1259593, 0.1638842, 0.1454304, 0.1581726, 0.1725864, 
    0.1830131, 0.105127, 0.1275106, 0.1321172, 0.07327046, 0.08735588, 
    0.05294324, 0.08772171, 0.157571, 0.1189818, 0.1423295, 0.2092124, 
    0.2000562, 0.1537932, 0.1168391, 0.1183041, 0.04867758, 0.1461275, 
    0.02734825, 0.05334746, 0.1507823, 0.1874681, 0.1565501,
  0.04104387, 0.01509139, 0.01579053, 0.01309616, 0.0235183, 0.02509765, 
    0.04832772, 0.07077701, 0.04509103, 0.01608269, 0.02625458, 0.0139406, 
    0.001905315, 0.01733692, 0.2281132, 0.04180108, 0.0492605, 0.0532282, 
    0.04789714, 0.06170686, 0.06253705, 0.03848632, 0.03763129, 0.3553512, 
    0.02149733, 0.02164036, 0.04765617, 0.04988829, 0.05462601,
  0.005937182, 0.01125625, 0.01059144, 0.005543022, 0.005241043, 0.007054543, 
    0.004177243, 0.01495422, 0.01320202, 0.001695074, 6.304409e-05, 
    0.0007353139, 0.02493714, 0.003101175, 0.008920287, 0.02923218, 
    0.02022288, 0.01613965, 0.015588, 0.0131581, 0.007938528, 0.002302606, 
    0.006069279, 0.008367474, 0.02928404, 0.005966738, 0.004612065, 
    0.002812795, 0.004434126,
  0.01345113, 0.01571285, 5.440398e-05, 0.003505831, -0.00177133, 
    0.0001734705, 0.0003332502, 0.006068994, 0.003183565, 0.0003967603, 
    -5.368473e-05, 4.412271e-05, 0.00227367, 0.004119642, 0.005780553, 
    0.002381129, 0.003574879, 0.004890824, 0.00123039, 0.004131783, 
    0.0008116669, 0.00311868, 0.009770211, 0.01004939, 0.05618508, 
    0.05661029, 0.0005332172, 0.0008002135, 0.001942122,
  0.02564551, 0.001220309, 0.0002438513, 0.04797776, 0.001130113, 
    0.0002145531, 0.0001239452, 0.0007982008, 0.0004210772, -5.251002e-05, 
    0.00586616, 0.0006964209, 0.01100958, 0.0004429714, 0.0007373174, 
    0.0005700642, 0.0001719829, 0.0002800143, 0.0002811741, 0.0003205159, 
    0.001245732, 0.004856776, 0.04486623, 0.001222318, -1.149956e-05, 
    -3.75375e-07, -0.000265017, 0.0005119145, 0.005921399,
  0.01945177, 0.01512278, 0.003357421, 0.005109309, 0.000304004, 
    0.0003670641, 0.0004814869, 0.001063243, 0.02768759, 0.01470654, 
    0.0003933485, 0.002319387, 0.005852737, 0.0005596408, 0.0005229226, 
    0.0001462497, 0.000803565, 0.0003245309, 0.0005206917, 0.0002034776, 
    0.001494934, 0.006278916, 0.0513423, 0.0686219, 0.03446087, 0.0005866271, 
    0.006667537, 0.0004693022, 0.001583661,
  0.0007902353, 0.0009479398, 2.794949e-07, 0.001039694, 5.921844e-07, 
    2.361789e-06, 0.006745859, 1.697496e-05, -8.747212e-05, 0.0005550632, 
    0.0005647022, 0.003292939, 0.00281737, 0.001697591, 0.0004894831, 
    0.0002539991, 0.000898699, 0.001856459, 0.00617341, 0.005227387, 
    0.00315455, 0.004860768, 0.1236787, 0.03852033, 0.0004122357, 
    0.001306367, 0.003566002, 0.01608242, 0.005774489,
  6.302923e-07, 5.073767e-07, 2.173239e-08, 2.709676e-09, 2.599061e-08, 
    0.0100393, 0.0001638336, 0.0006037147, 0.0715949, 0.003803048, 
    0.002142728, 0.003132757, 2.961338e-05, 2.496481e-05, 0.000113486, 
    0.0006540833, 0.001350383, 0.00282612, 0.0233001, 0.04945549, 0.04648063, 
    0.02850413, 0.0001587016, -0.0008005956, 2.141514e-05, 7.520162e-05, 
    0.002411006, 0.009366293, 1.251622e-06,
  9.251165e-07, -6.128181e-06, 2.271392e-05, -9.794792e-07, 1.603596e-07, 
    2.445285e-08, -0.0003914304, 0.06153126, 0.246334, 0.01612664, 0.1311502, 
    0.09973609, 0.05372671, 0.008902071, 0.02769552, 0.00664447, 0.01050969, 
    0.005440214, 0.01402083, 0.05966769, 2.930858e-07, 0.009054335, 
    0.01601057, 0.006812859, 0.006276278, 0.00417595, 0.002118667, 
    0.007827649, 0.01520189,
  0.003088829, 0.001259469, -6.65126e-05, 0.1293213, -8.636371e-05, 
    2.463061e-07, 0.01121194, -3.473573e-05, -4.020605e-05, 0.005504583, 
    0.1516552, 0.1791115, 0.2651526, 0.2950972, 0.2634886, 0.2038669, 
    0.2721785, 0.1244294, 0.1145903, 0.03322173, 0.00319878, 0.02640526, 
    0.01268681, 0.06700106, 0.08212823, 0.1146687, 0.07352423, 0.065935, 
    0.07799879,
  0.07013594, 0.06560083, 0.02586388, 0.002232397, 0.0005886016, 
    3.635084e-05, 0.006137845, 0.09471744, 0.04421055, 0.04030764, 0.1143467, 
    0.126965, 0.4958321, 0.4144083, 0.3927101, 0.3480147, 0.3490513, 
    0.3533585, 0.2093496, 0.07802013, 0.02582038, 0.003562984, 0.03257527, 
    0.08824747, 0.1264988, 0.2683139, 0.2352175, 0.17108, 0.1172869,
  0.1997957, 0.01731613, 0.01114618, 0.03497639, 0.0575217, 0.03207197, 
    0.02902213, 0.02204515, 0.06555051, 0.04469615, 0.117282, 0.1333818, 
    0.1134676, 0.1612662, 0.3447468, 0.3418404, 0.1757624, 0.2607779, 
    0.08182476, 0.007235427, 0.00497197, 0.02743814, 0.08810259, 0.07764461, 
    0.2186543, 0.1184516, 0.2082069, 0.1563843, 0.1364127,
  0.4482673, 0.2429868, 0.1551974, 0.2727355, 0.2095111, 0.282857, 0.1739724, 
    0.08046162, 0.03526386, 0.04710731, 0.04728207, 0.03764543, 0.01949723, 
    0.1621757, 0.2009156, 0.2981701, 0.0713367, 0.1261218, 0.1998593, 
    0.1312818, 0.1298148, 0.2298103, 0.06142121, 0.2219547, 0.3109533, 
    0.1483674, 0.1009528, 0.2100793, 0.5491872,
  0.5002718, 0.2932014, 0.2457987, 0.3788669, 0.4189859, 0.4275268, 0.408703, 
    0.3787845, 0.3104758, 0.3240489, 0.3012394, 0.2850632, 0.2974643, 
    0.354881, 0.3770077, 0.3395886, 0.330088, 0.3243049, 0.3046488, 
    0.2156415, 0.2430235, 0.1925451, 0.1355888, 0.2574722, 0.1824908, 
    0.08798413, 0.1060361, 0.3911901, 0.4760444,
  0.004640122, 0.00443754, 0.004234958, 0.004032376, 0.003829793, 
    0.003627211, 0.003424629, 0.001301511, 0.004058764, 0.006816017, 
    0.00957327, 0.01233052, 0.01508778, 0.01784503, 0.02451495, 0.02478543, 
    0.02505591, 0.02532639, 0.02559687, 0.02586735, 0.02613784, 0.01719383, 
    0.01436868, 0.01154353, 0.008718378, 0.005893226, 0.003068074, 
    0.0002429223, 0.004802188,
  0.1665531, 0.07786223, 0.027105, 0.0137185, 0.0029773, 0.01100405, 
    0.01279142, 0.01604953, 0.005749984, 0.004345212, 0.005519833, 
    0.01381133, 0.09684673, -0.000636037, 0.3080034, 0.3879181, 0.3972487, 
    0.3131012, 0.1610572, 0.394033, 0.5058459, 0.516193, 0.1290483, 
    0.08081655, 0.1873081, 0.3980148, 0.2482877, 0.1304784, 0.18642,
  0.2128334, 0.08262611, 0.110055, 0.02200497, 0.1001085, 0.1974936, 
    0.02951508, 0.163605, 0.1778601, 0.1510616, 0.1983053, 0.2327499, 
    0.1051282, 0.1297559, 0.379321, 0.3548304, 0.3319443, 0.3675543, 
    0.2264093, 0.2345456, 0.3021316, 0.2696268, 0.2584552, 0.321611, 
    0.2527386, 0.3756772, 0.4497554, 0.4138217, 0.2526986,
  0.2487393, 0.07804418, 0.05823204, 0.0726455, 0.1094063, 0.0867682, 
    0.1520795, 0.104537, 0.09927787, 0.10627, 0.1053578, 0.140208, 0.1804902, 
    0.1841017, 0.1624868, 0.1846008, 0.2379789, 0.1945482, 0.182327, 
    0.1147579, 0.09300372, 0.0746361, 0.1195234, 0.09673954, 0.1548929, 
    0.2810131, 0.2677827, 0.2369053, 0.2484804,
  0.1295394, 0.1041009, 0.1339858, 0.1231649, 0.13474, 0.143151, 0.1525232, 
    0.08148355, 0.09914035, 0.1050203, 0.05215217, 0.06140079, 0.03628344, 
    0.05456398, 0.115734, 0.08074217, 0.09757219, 0.1494516, 0.1447376, 
    0.105393, 0.08537526, 0.08330745, 0.03317852, 0.1368007, 0.01927139, 
    0.03581529, 0.1140788, 0.1544068, 0.1342101,
  0.02641192, 0.009541733, 0.01021079, 0.008675532, 0.01301005, 0.01558089, 
    0.03273967, 0.04599185, 0.02641375, 0.009356542, 0.01459647, 0.008641751, 
    0.001304705, 0.008781853, 0.1879033, 0.02652453, 0.03055249, 0.03287216, 
    0.02782618, 0.04036827, 0.04409937, 0.02334702, 0.02457146, 0.3321902, 
    0.01676102, 0.01198018, 0.03034711, 0.03489732, 0.03711728,
  0.004331294, 0.007982085, 0.009166721, 0.003451418, 0.00329472, 
    0.004172492, 0.003114765, 0.009055377, 0.01019736, 0.001355563, 
    2.23382e-05, 0.001919911, 0.02226943, 0.002147861, 0.004837801, 
    0.01574246, 0.01133626, 0.008469433, 0.008840488, 0.008212882, 
    0.004273844, 0.001647831, 0.003724368, 0.005811087, 0.02341898, 
    0.003539494, 0.002582117, 0.001726032, 0.002471435,
  0.009828812, 0.01353814, -4.790392e-05, 0.002642774, -0.00127903, 
    0.0001090202, 0.0002350706, 0.002855887, 0.001516584, 0.0002945016, 
    -3.477562e-05, 6.153331e-05, 0.001288982, 0.002279531, 0.002886861, 
    0.001340511, 0.002218518, 0.002862737, 0.0006961508, 0.002101158, 
    0.0005532754, 0.002331704, 0.007205606, 0.007762068, 0.04909464, 
    0.05342193, 0.0004078996, 0.0005938979, 0.001420694,
  0.01915108, 0.000850256, 0.0001919432, 0.03376081, 0.0005373003, 
    0.0001537369, 8.024171e-05, 0.000583519, 0.0002435471, -3.942999e-05, 
    0.00390908, 0.0003123634, 0.004988001, 0.0002358432, 0.0003959532, 
    0.0003154193, 0.0001307209, 0.0002082396, 0.0002045605, 0.0002362246, 
    0.0009401617, 0.003548446, 0.03320344, 0.001942558, -4.462769e-06, 
    -1.156004e-06, -0.0001634464, 0.000360513, 0.004378472,
  0.01369994, 0.01419498, 0.002618093, 0.003395961, 0.0002075563, 
    0.0002721474, 0.0003582881, 0.0006098418, 0.02422824, 0.02326482, 
    0.0002686852, 0.001559993, 0.002779566, 0.0002931042, 0.0002659019, 
    0.0001056015, 0.0003888312, 0.0002340167, 0.0003756578, 0.0001429999, 
    0.001066577, 0.004250147, 0.03625318, 0.04775909, 0.03388174, 
    0.0002720221, 0.003095537, 0.0003359871, 0.001117385,
  0.0006098374, 0.0004898527, -4.708922e-07, 0.001980247, 2.018642e-07, 
    1.570609e-06, 0.004022913, 1.234475e-05, -8.563073e-05, 0.0003996787, 
    0.000371167, 0.001708771, 0.001144425, 0.0007762845, 0.0002380259, 
    0.0001239463, 0.0004110495, 0.0009761367, 0.002832043, 0.003174601, 
    0.001728769, 0.002343713, 0.1137653, 0.03688853, 0.0002331503, 
    0.0005135358, 0.001993741, 0.009287243, 0.005656529,
  6.105029e-07, 4.976914e-07, 2.205404e-08, 2.088921e-09, 2.583484e-08, 
    0.006758232, -0.0003240265, 0.0003165462, 0.06040253, 0.0007864822, 
    0.001173147, 0.001429087, 2.167002e-05, 1.778328e-05, 8.185994e-05, 
    0.0004772926, 0.0009320533, 0.0019639, 0.0167225, 0.03630773, 0.03264695, 
    0.02272336, 0.0001089588, -0.0009027176, 1.446453e-05, 5.585147e-05, 
    0.001697244, 0.006765248, 1.837963e-07,
  4.915315e-07, -4.264959e-06, 0.0002197552, -6.014747e-07, 1.569281e-07, 
    2.412689e-08, -0.0003666285, 0.05821361, 0.2268049, 0.01030225, 
    0.08178547, 0.05701654, 0.02865602, 0.004469268, 0.01748371, 0.004234883, 
    0.005305866, 0.003860422, 0.009365922, 0.04200189, 2.724856e-07, 
    0.01271604, 0.01297563, 0.002641922, 0.002916947, 0.002704454, 
    0.001526597, 0.005803532, 0.0128212,
  0.002240786, 0.000796431, -6.728375e-05, 0.124066, -7.479485e-05, 
    2.646632e-07, 0.009863052, -2.193408e-05, -3.411163e-05, 0.003886039, 
    0.1291141, 0.144887, 0.2261483, 0.2464741, 0.2155111, 0.1581708, 
    0.2049035, 0.08444061, 0.07663171, 0.03056032, 0.002681365, 0.02028274, 
    0.009840271, 0.04605239, 0.05184479, 0.06865456, 0.03937083, 0.03597561, 
    0.06213184,
  0.05581533, 0.05479457, 0.0177878, 0.001304872, 0.0003868128, 2.055764e-05, 
    0.005118689, 0.08767528, 0.03974552, 0.03621086, 0.1009579, 0.109365, 
    0.4146085, 0.3335642, 0.2979318, 0.2640638, 0.2660148, 0.2614546, 
    0.1471566, 0.07249171, 0.01966826, 0.002105569, 0.03034133, 0.07671507, 
    0.1279263, 0.2392435, 0.1668262, 0.1090237, 0.07823414,
  0.1776532, 0.0134407, 0.007516987, 0.02696794, 0.04637919, 0.02539252, 
    0.02898794, 0.0231058, 0.06251448, 0.03876328, 0.1050501, 0.1108837, 
    0.09532185, 0.1348228, 0.2684075, 0.2522106, 0.1505781, 0.2287936, 
    0.06378638, 0.006818797, 0.003531741, 0.01993601, 0.08278502, 0.06049347, 
    0.175904, 0.1051569, 0.1446773, 0.09964924, 0.0969788,
  0.3551989, 0.2002759, 0.131331, 0.2321473, 0.1705978, 0.2778695, 0.165353, 
    0.07903392, 0.03388325, 0.03943187, 0.03642172, 0.02971615, 0.01397463, 
    0.1388595, 0.1772171, 0.2930042, 0.04611187, 0.1086499, 0.1754174, 
    0.1377178, 0.106943, 0.2024367, 0.04520106, 0.1990227, 0.2684639, 
    0.1287363, 0.09166034, 0.1889972, 0.4598801,
  0.4149453, 0.247496, 0.2166142, 0.3220978, 0.324132, 0.3499325, 0.3459913, 
    0.3200245, 0.2609556, 0.2700472, 0.2474866, 0.2327294, 0.2453114, 
    0.2846219, 0.3097847, 0.2782703, 0.2737532, 0.2618352, 0.2522582, 
    0.1649073, 0.1968593, 0.1518993, 0.1102704, 0.2214035, 0.1624266, 
    0.0747574, 0.09297052, 0.3651594, 0.3998104,
  0.003059692, 0.003145799, 0.003231905, 0.003318012, 0.003404119, 
    0.003490226, 0.003576333, 0.001442755, 0.003315693, 0.005188631, 
    0.007061569, 0.008934507, 0.01080745, 0.01268038, 0.01533062, 0.01508733, 
    0.01484403, 0.01460074, 0.01435744, 0.01411415, 0.01387085, 0.008535612, 
    0.006819864, 0.005104115, 0.003388366, 0.001672616, -4.313255e-05, 
    -0.001758882, 0.002990806,
  0.1272504, 0.04453463, 0.01716991, 0.01039083, 0.002094779, 0.006544206, 
    0.006013313, 0.003623033, 0.005783634, 0.0008784309, 0.002124216, 
    0.01188434, 0.08598991, 0.0004061498, 0.3804179, 0.3064502, 0.3617271, 
    0.3491199, 0.1594227, 0.4568298, 0.4906465, 0.5428125, 0.1231262, 
    0.07283366, 0.1463145, 0.3802632, 0.2263498, 0.1200072, 0.1204923,
  0.2185735, 0.08294852, 0.0921607, 0.01942223, 0.08992494, 0.1774462, 
    0.0257516, 0.1474303, 0.1669688, 0.1453122, 0.1966519, 0.2360803, 
    0.1003902, 0.1207679, 0.3596141, 0.3370607, 0.3126123, 0.3417317, 
    0.2080228, 0.2275116, 0.2869225, 0.2525771, 0.2441517, 0.3035753, 
    0.2334987, 0.3359036, 0.3961601, 0.3707286, 0.2280673,
  0.2272438, 0.06555989, 0.05090754, 0.06365674, 0.09307145, 0.07502826, 
    0.1338293, 0.09167464, 0.08508056, 0.08815768, 0.08955552, 0.1194234, 
    0.1508431, 0.1560421, 0.133321, 0.1588376, 0.2085185, 0.1662897, 0.15483, 
    0.09908637, 0.07825945, 0.06220677, 0.1024456, 0.08202218, 0.1344005, 
    0.2587412, 0.243329, 0.2119073, 0.2280403,
  0.1119228, 0.08957747, 0.1142805, 0.1023954, 0.1151438, 0.1216716, 
    0.1290458, 0.06755246, 0.08156738, 0.08845343, 0.04160554, 0.04896697, 
    0.02880538, 0.04092579, 0.0884603, 0.06209791, 0.07462086, 0.1157865, 
    0.1109929, 0.07800841, 0.06535091, 0.06272262, 0.02631706, 0.1696946, 
    0.01481469, 0.02860728, 0.09612995, 0.1288109, 0.1151588,
  0.01896084, 0.007213573, 0.007218475, 0.006660981, 0.009175831, 0.01156116, 
    0.02381303, 0.03322419, 0.01926989, 0.006759045, 0.009718496, 
    0.006015076, 0.001063401, 0.005476916, 0.1743471, 0.01819832, 0.02088856, 
    0.02240611, 0.01958168, 0.03086512, 0.03297043, 0.01721133, 0.0171928, 
    0.3368458, 0.01191875, 0.007736596, 0.02213265, 0.02769772, 0.02679796,
  0.003593613, 0.006167821, 0.01005535, 0.002275344, 0.002609455, 
    0.002731598, 0.002427565, 0.005364669, 0.007127375, 0.001158506, 
    -9.223116e-06, 0.005188984, 0.02649734, 0.001654584, 0.003321147, 
    0.008222788, 0.006067463, 0.005140819, 0.006060645, 0.004896308, 
    0.002924791, 0.001382094, 0.002804441, 0.004633296, 0.02799233, 
    0.002646094, 0.001854017, 0.001365134, 0.001814043,
  0.008077988, 0.01158187, -0.0001256908, 0.002201052, -0.001180419, 
    8.949157e-05, 0.0001933728, 0.001870177, 0.001039249, 0.0002440201, 
    -2.607441e-05, 6.049989e-05, 0.0008006046, 0.001652633, 0.001991102, 
    0.0008915776, 0.001680798, 0.002097818, 0.0005174925, 0.001400913, 
    0.0004425149, 0.001952746, 0.005983207, 0.006590448, 0.05897354, 
    0.05759697, 0.0003427424, 0.0004948262, 0.001174228,
  0.01592727, 0.0006756005, 0.0001439314, 0.02797175, 0.0003238613, 
    0.0001267522, 6.685231e-05, 0.0004856894, 0.0001865207, -0.0004051369, 
    0.003035774, 0.0002074754, 0.003165672, 0.0001706112, 0.0002676933, 
    0.0002375089, 0.0001105346, 0.0001816483, 0.000169049, 0.0002041024, 
    0.0007947353, 0.002947231, 0.02738182, 0.008401677, -3.34093e-06, 
    -3.799594e-06, -0.0001434258, 0.0002951785, 0.00365461,
  0.01095435, 0.02625387, 0.004827514, 0.00313907, 0.0001726642, 
    0.0002238996, 0.0002934999, 0.0004613647, 0.04022697, 0.05899202, 
    0.0002113338, 0.001171739, 0.001780647, 0.000210794, 0.0001897293, 
    8.664602e-05, 0.0002836471, 0.0001967532, 0.0003060344, 0.0001182393, 
    0.0008168957, 0.003341982, 0.02903748, 0.07473364, 0.06979752, 
    0.0001884132, 0.001693679, 0.0002736197, 0.000885105,
  0.01320475, 0.0007908401, -9.431117e-05, 0.002223929, 1.992049e-07, 
    1.345858e-06, 0.02237441, 1.03175e-05, -0.001946307, 0.0003259881, 
    0.0002933087, 0.001116887, 0.0006748106, 0.0004360077, 0.0001645719, 
    9.099558e-05, 0.0002769832, 0.0006929411, 0.001819863, 0.002331403, 
    0.001157858, 0.001456389, 0.1735178, 0.04391916, 0.0001665902, 
    0.0003134091, 0.001383439, 0.006661479, 0.02759036,
  5.996192e-07, 4.936372e-07, 2.232347e-08, 2.085891e-09, 2.567332e-08, 
    0.005285915, -0.0004148663, 0.0002317761, 0.1420334, -0.0003062226, 
    0.0008485189, 0.0007845053, 1.810304e-05, 1.488609e-05, 6.770355e-05, 
    0.0003902318, 0.0007410108, 0.001577942, 0.01359419, 0.02985369, 
    0.02545313, 0.0206406, 8.672169e-05, -0.001642074, 1.181078e-05, 
    4.724906e-05, 0.001388259, 0.005534925, 1.249336e-07,
  4.308702e-07, -1.856716e-06, -2.794143e-06, -2.724375e-07, 1.582067e-07, 
    2.385336e-08, -0.0003601428, 0.06159914, 0.2327619, 0.009250592, 
    0.05350653, 0.03466958, 0.01684181, 0.002953181, 0.01004639, 0.002603792, 
    0.003385315, 0.003136369, 0.007196028, 0.03291225, 2.704567e-07, 
    0.04967294, 0.02872894, 0.001708182, 0.001798657, 0.002144675, 
    0.00123692, 0.004827218, 0.01062827,
  0.002120944, 0.0003942589, -0.0001266655, 0.1261869, -7.173081e-05, 
    2.933214e-07, 0.009738481, -1.540635e-05, -3.041479e-05, 0.003267054, 
    0.1350426, 0.1147606, 0.1804693, 0.1952522, 0.1684278, 0.1182108, 
    0.1603442, 0.06007098, 0.05805574, 0.02965281, 0.002911872, 0.02569102, 
    0.01598845, 0.03295236, 0.032553, 0.0414727, 0.02426498, 0.02185065, 
    0.05421384,
  0.04902452, 0.05793206, 0.0191314, 0.001324085, 0.0002906169, 1.345825e-05, 
    0.005453888, 0.08741625, 0.04433013, 0.04612397, 0.1199935, 0.1186112, 
    0.350662, 0.2804152, 0.2358207, 0.2082477, 0.2072875, 0.2011119, 
    0.1049334, 0.08391174, 0.01753781, 0.001726135, 0.04237979, 0.1001402, 
    0.1311624, 0.2006556, 0.1304257, 0.0768175, 0.05552875,
  0.1514112, 0.01503792, 0.006415742, 0.0335878, 0.05264177, 0.03479949, 
    0.05089413, 0.03682095, 0.08930448, 0.06048458, 0.1158183, 0.1090876, 
    0.08173279, 0.1296924, 0.2102175, 0.1994097, 0.1622606, 0.2210512, 
    0.06329492, 0.0109551, 0.007117011, 0.01520906, 0.072998, 0.04963347, 
    0.1450158, 0.09263843, 0.1097037, 0.0718045, 0.07283854,
  0.2946771, 0.1720544, 0.1209569, 0.1914507, 0.1393023, 0.2897874, 
    0.1712571, 0.09315428, 0.04120675, 0.04945304, 0.03186313, 0.02677771, 
    0.01186087, 0.1210937, 0.1686547, 0.2651948, 0.03392645, 0.09723135, 
    0.1678812, 0.1597531, 0.09244891, 0.185683, 0.03395353, 0.1876506, 
    0.2427967, 0.1175402, 0.09296799, 0.1669485, 0.3626364,
  0.3640577, 0.2075234, 0.1976617, 0.28016, 0.2690134, 0.306722, 0.2988209, 
    0.2826334, 0.2311657, 0.2299257, 0.2161837, 0.197594, 0.2051991, 
    0.2391291, 0.2589929, 0.2317706, 0.2364225, 0.2243876, 0.2223069, 
    0.1393241, 0.1671264, 0.1313871, 0.09552458, 0.2004746, 0.149576, 
    0.06879763, 0.09138416, 0.3448593, 0.3474061 ;

 average_DT = 730 ;

 average_T1 = 167 ;

 average_T2 = 897 ;

 climatology_bounds =
  167, 897 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
