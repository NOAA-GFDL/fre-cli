netcdf atmos_level_cmip.185001-185412.ps {
dimensions:
    time = UNLIMITED ; // (60 currently)
    bnds = 2 ;
    lat = 2 ;
    lon = 2 ;
variables:
    double average_DT(time) ;
        average_DT:long_name = "Length of average period" ;
        average_DT:units = "days" ;
        average_DT:missing_value = 1.e+20 ;
        average_DT:_FillValue = 1.e+20 ;
    double average_T1(time) ;
        average_T1:long_name = "Start time for average period" ;
        average_T1:units = "days since 1850-01-01 00:00:00" ;
        average_T1:missing_value = 1.e+20 ;
        average_T1:_FillValue = 1.e+20 ;
    double average_T2(time) ;
        average_T2:long_name = "End time for average period" ;
        average_T2:units = "days since 1850-01-01 00:00:00" ;
        average_T2:missing_value = 1.e+20 ;
        average_T2:_FillValue = 1.e+20 ;
    double bnds(bnds) ;
        bnds:long_name = "vertex number" ;
    double lat(lat) ;
        lat:long_name = "latitude" ;
        lat:units = "degrees_N" ;
        lat:axis = "Y" ;
        lat:bounds = "lat_bnds" ;
    double lat_bnds(lat, bnds) ;
        lat_bnds:long_name = "latitude bounds" ;
        lat_bnds:units = "degrees_N" ;
        lat_bnds:axis = "Y" ;
    double lon(lon) ;
        lon:long_name = "longitude" ;
        lon:units = "degrees_E" ;
        lon:axis = "X" ;
        lon:bounds = "lon_bnds" ;
    double lon_bnds(lon, bnds) ;
        lon_bnds:long_name = "longitude bounds" ;
        lon_bnds:units = "degrees_E" ;
        lon_bnds:axis = "X" ;
    float ps(time, lat, lon) ;
        ps:long_name = "Surface Air Pressure" ;
        ps:units = "Pa" ;
        ps:missing_value = 1.e+20f ;
        ps:_FillValue = 1.e+20f ;
        ps:cell_methods = "time: mean" ;
        ps:cell_measures = "area: area" ;
        ps:time_avg_info = "average_T1,average_T2,average_DT" ;
        ps:standard_name = "surface_air_pressure" ;
        ps:interp_method = "conserve_order2" ;
    double time(time) ;
        time:long_name = "time" ;
        time:units = "days since 1850-01-01 00:00:00" ;
        time:axis = "T" ;
        time:calendar_type = "NOLEAP" ;
        time:calendar = "noleap" ;
        time:bounds = "time_bnds" ;
    double time_bnds(time, bnds) ;
        time_bnds:long_name = "time axis boundaries" ;
        time_bnds:units = "days since 1850-01-01 00:00:00" ;
        time_bnds:missing_value = 1.e+20 ;
        time_bnds:_FillValue = 1.e+20 ;

// global attributes:
        :filename = "atmos_level_cmip.185001-185412.ps.nc" ;
        :title = "ESM4_historical_D1" ;
        :associated_files = "area: 18540101.grid_spec.nc" ;
        :grid_type = "regular" ;
        :grid_tile = "N/A" ;
        :history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 18540101.atmos_level_cmip --interp_method conserve_order2 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field ap,b,ap_bnds,b_bnds,lev_bnds,ps,cl,clw,cli,mc,pfull,phalf,tntrl,tntrs,tntrlcs,tntrscs,tntpbl,tntscp,tnhuspbl,tnhusscp,ec550aer,rsu,rsd,rsucs,rsdcs,rsuaf,rsdaf,rsucsaf,rsdcsaf,time_bnds --output_file out.nc" ;
        :code_version = "$Name: bronx-10_performance_z1l $" ;
        :external_variables = "area" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 
    30, 31, 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31, 31, 28, 31, 30, 
    31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 
    396, 424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 
    820, 850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 
    1215, 1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 
    1580, 1611, 1641, 1672, 1703, 1733, 1764, 1794 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365, 396, 
    424, 455, 485, 516, 546, 577, 608, 638, 669, 699, 730, 761, 789, 820, 
    850, 881, 911, 942, 973, 1003, 1034, 1064, 1095, 1126, 1154, 1185, 1215, 
    1246, 1276, 1307, 1338, 1368, 1399, 1429, 1460, 1491, 1519, 1550, 1580, 
    1611, 1641, 1672, 1703, 1733, 1764, 1794, 1825 ;

 bnds = 1, 2 ;

 lat = -89.5, -88.5 ;

 lat_bnds =
  -90, -89,
  -89, -88 ;

 lon = 0.625, 1.875 ;

 lon_bnds =
  0, 1.25,
  1.25, 2.5 ;

 ps = 
  69429.03, 69408.66, 69388.28, 69367.91, 69347.53, 69327.16, 69306.78, 
    69286.4, 69266.02, 69245.65, 69225.27, 69204.9, 69184.52, 69164.15, 
    69143.77, 69123.4, 69103.02, 69082.64, 69062.27, 69041.89, 69021.52, 
    69001.14, 68980.77, 68960.39, 68940.02, 68919.64, 68899.26, 68878.88, 
    68858.51, 68838.13, 68817.76, 68797.38, 68777.01, 68756.63, 68736.26, 
    68715.88, 68695.5, 68675.12, 68654.75, 68634.38, 68614, 68593.62, 
    68573.25, 68552.88, 68532.5, 68512.12, 68491.74, 68471.37, 68450.99, 
    68430.62, 68410.24, 68389.87, 68369.49, 68349.12, 68328.73, 68308.36, 
    68287.98, 68267.61, 68247.23, 68226.86, 68206.48, 68186.11, 68165.73, 
    68145.36, 68592.73, 68589.53, 68586.34, 68583.14, 68579.95, 68576.76, 
    68573.56, 68570.37, 68567.17, 68563.98, 68560.78, 68557.59, 68554.39, 
    68551.2, 68548, 68544.8, 68541.62, 68538.42, 68535.23, 68532.03, 
    68528.84, 68525.64, 68522.45, 68519.25, 68516.05, 68512.86, 68509.66, 
    68506.48, 68503.28, 68500.09, 68496.89, 68493.7, 68490.5, 68487.3, 
    68484.11, 68480.91, 68477.72, 68474.52, 68471.34, 68468.14, 68464.95, 
    68461.75, 68458.55, 68455.36, 68452.16, 68448.97, 68445.77, 68442.58, 
    68439.38, 68436.19, 68433, 68429.8, 68426.61, 68423.41, 68420.22, 
    68417.02, 68413.83, 68410.63, 68407.44, 68404.24, 68401.05, 68397.86, 
    68394.66, 68391.47, 68388.27, 68385.08, 68381.88, 68378.69, 68375.49, 
    68372.3, 68369.1, 68365.91, 67715.44, 67732.84, 67750.23, 67767.64, 
    67785.04, 67802.45, 67819.84, 67837.25, 67854.65, 67872.05, 67889.45, 
    67906.85, 67924.26, 67941.66, 67959.05, 67976.46, 67993.86, 68011.27, 
    68028.66, 68046.07, 68063.47, 68080.87, 68098.27, 68115.67, 68133.08, 
    68150.48, 68167.88, 68185.28, 68202.68, 68220.09, 68237.48, 68254.88, 
    68272.29, 68289.69, 68307.09, 68324.49, 68341.9, 68359.3, 68376.7, 
    68394.1, 68411.5, 68428.91, 68446.3, 68463.7, 68481.11, 68498.51, 
    68515.91, 68533.31, 68550.72, 68568.12, 68585.52, 68602.92, 68620.32, 
    68637.73, 68655.12, 68672.52, 68689.93, 68707.33, 68724.73, 68742.13, 
    68759.53, 68776.94, 68794.34, 68811.74, 68829.14, 68846.55, 68863.95, 
    68881.34, 68898.75, 68916.15, 68933.55, 68950.95, 69104.03, 69110.2, 
    69116.37, 69122.54, 69128.71, 69134.88, 69141.05, 69147.21, 69153.38, 
    69159.55, 69165.72, 69171.89, 69178.06, 69184.23, 69190.4, 69196.56, 
    69202.73, 69208.91, 69215.07, 69221.24, 69227.41, 69233.58, 69239.75, 
    69245.91, 69252.09, 69258.25, 69264.42, 69270.59, 69276.76, 69282.93, 
    69289.09, 69295.27 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 
    349.5, 380.5, 410, 439.5, 470, 500.5, 531, 561.5, 592.5, 623, 653.5, 684, 
    714.5, 745.5, 775, 804.5, 835, 865.5, 896, 926.5, 957.5, 988, 1018.5, 
    1049, 1079.5, 1110.5, 1140, 1169.5, 1200, 1230.5, 1261, 1291.5, 1322.5, 
    1353, 1383.5, 1414, 1444.5, 1475.5, 1505, 1534.5, 1565, 1595.5, 1626, 
    1656.5, 1687.5, 1718, 1748.5, 1779, 1809.5 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365,
  365, 396,
  396, 424,
  424, 455,
  455, 485,
  485, 516,
  516, 546,
  546, 577,
  577, 608,
  608, 638,
  638, 669,
  669, 699,
  699, 730,
  730, 761,
  761, 789,
  789, 820,
  820, 850,
  850, 881,
  881, 911,
  911, 942,
  942, 973,
  973, 1003,
  1003, 1034,
  1034, 1064,
  1064, 1095,
  1095, 1126,
  1126, 1154,
  1154, 1185,
  1185, 1215,
  1215, 1246,
  1246, 1276,
  1276, 1307,
  1307, 1338,
  1338, 1368,
  1368, 1399,
  1399, 1429,
  1429, 1460,
  1460, 1491,
  1491, 1519,
  1519, 1550,
  1550, 1580,
  1580, 1611,
  1611, 1641,
  1641, 1672,
  1672, 1703,
  1703, 1733,
  1733, 1764,
  1764, 1794,
  1794, 1825 ;
}