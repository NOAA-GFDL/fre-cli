netcdf atmos.1980-1981.alb_sfc.01 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:15 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.01.nc reduced/atmos.1980-1981.alb_sfc.01.nc\n",
			"Mon Aug 25 14:40:02 2025: cdo -O -s -select,month=1 merged_output.nc monthly_nc_files/all_years.1.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.23267, 76.23267, 76.23267, 76.23267, 76.23267, 76.23267, 76.23267, 
    76.23283, 76.23283, 76.23283, 76.23283, 76.23283, 76.23283, 76.23283, 
    76.22655, 76.22655, 76.22655, 76.22655, 76.22655, 76.22655, 76.22655, 
    76.24745, 76.24745, 76.24745, 76.24745, 76.24745, 76.24745, 76.24745, 
    76.23267,
  76.49063, 76.2739, 76.16951, 76.07027, 76.06326, 76.0631, 76.04036, 
    76.02043, 76.05639, 76.13631, 76.18135, 76.29651, 76.37398, 75.76569, 
    76.9165, 72.44071, 74.8634, 71.20247, 67.30618, 73.26184, 74.97375, 
    76.02705, 74.67429, 67.05026, 73.98146, 66.56528, 73.06624, 69.02693, 
    76.53729,
  39.97103, 42.6682, 44.53755, 64.21826, 72.20937, 72.37304, 50.66593, 
    72.71266, 72.61586, 71.8877, 72.55252, 72.91833, 67.9734, 43.1772, 
    6.316841, 6.134087, 6.385586, 6.609262, 6.361966, 31.15282, 28.50522, 
    28.47579, 57.97995, 61.37165, 61.25329, 36.83862, 29.81477, 6.501078, 
    9.452572,
  4.604814, 4.676425, 4.88024, 4.774986, 4.70841, 4.611859, 4.729652, 
    4.60995, 4.726584, 4.777658, 4.784083, 4.667452, 4.641747, 4.805507, 
    4.88038, 4.823759, 4.604949, 4.734746, 4.774827, 5.012154, 5.095692, 
    5.043339, 5.068858, 4.993554, 4.793861, 4.582891, 11.80887, 4.758969, 
    4.619605,
  4.181644, 4.29203, 4.240377, 4.365281, 4.331936, 4.303432, 4.333741, 
    4.219655, 4.246339, 4.268391, 4.408224, 4.381993, 4.472157, 4.457103, 
    4.408319, 4.423872, 4.26683, 4.349495, 4.334805, 4.36984, 4.372739, 
    4.351821, 4.36996, 8.624498, 4.864033, 4.402624, 4.31779, 4.220292, 
    4.268884,
  4.19315, 4.110131, 4.330577, 4.171401, 4.031809, 4.037183, 4.061778, 
    4.111396, 3.904371, 4.114984, 3.956092, 4.27564, 4.127986, 4.03132, 
    10.26554, 4.03397, 4.181191, 4.024014, 4.007151, 3.869534, 4.019423, 
    4.015054, 4.099564, 10.00854, 4.543853, 4.176139, 3.931249, 3.915059, 
    4.019889,
  4.002278, 4.055106, 12.60526, 3.835495, 4.003094, 4.030794, 3.793797, 
    3.98241, 3.812176, 4.084562, 10.31545, 15.91999, 10.38852, 3.900531, 
    4.041914, 3.860006, 3.833383, 3.652178, 3.628936, 3.837499, 4.184121, 
    4.16984, 3.951359, 4.626525, 9.637185, 3.736104, 3.763609, 3.94642, 
    4.003505,
  3.637431, 10.10725, 12.32863, 3.644678, 3.550663, 3.472622, 3.73898, 
    3.708578, 3.67863, 3.463841, 12.17498, 11.17589, 3.528108, 3.519952, 
    3.640141, 3.669344, 3.364697, 3.63422, 3.616143, 4.006081, 3.917354, 
    3.902304, 3.365593, 3.294021, 9.226721, 9.428365, 3.950979, 3.921249, 
    4.026099,
  3.402283, 6.494687, 8.727841, 9.370113, 3.341715, 3.321693, 3.478166, 
    3.410533, 3.525913, 3.263133, 4.596019, 3.289837, 4.356509, 3.561458, 
    3.446259, 3.489925, 3.390093, 3.768706, 3.592235, 3.989404, 3.660187, 
    3.752735, 3.485017, 8.749596, 8.551068, 8.945084, 3.742415, 3.562161, 
    3.732562,
  3.242565, 8.88798, 8.686348, 9.973007, 3.452828, 3.434671, 3.167229, 
    3.306105, 8.701897, 8.238229, 3.405158, 3.393892, 3.242504, 3.409903, 
    3.442074, 3.611695, 3.672125, 3.88739, 3.780538, 3.927022, 3.638591, 
    3.396252, 3.363677, 8.535877, 8.435765, 3.195887, 3.341912, 3.472915, 
    3.215913,
  10.18067, 10.25406, 10.58913, 9.625751, 14.27646, 3.462219, 5.420032, 
    3.563966, 3.456795, 3.501905, 4.116955, 3.423054, 3.32419, 3.538214, 
    3.642063, 3.58934, 3.819775, 3.586876, 3.85488, 3.518491, 3.498654, 
    3.592799, 8.591267, 7.262965, 3.595617, 3.721086, 3.329552, 3.759384, 
    9.009521,
  16.14083, 18.6687, 20.70445, 3.713118, 20.74915, 4.080397, 10.06667, 
    4.007038, 9.008829, 3.317509, 3.561971, 3.771078, 3.672481, 3.987378, 
    4.065104, 3.772914, 3.988953, 3.837881, 3.848425, 3.489404, 3.846314, 
    6.140777, 3.770617, 4.545951, 3.825474, 4.052248, 3.672032, 3.7641, 
    21.19227,
  20.48906, 16.26445, 17.19365, 16.614, 11.26028, 12.70199, 12.24097, 
    25.51131, 9.734715, 10.31121, 3.399524, 3.733083, 4.029523, 3.857799, 
    3.866054, 3.902126, 3.847343, 3.602057, 3.753562, 4.008671, 9.207573, 
    11.05214, 9.692469, 3.720354, 3.9571, 3.835543, 3.749384, 3.94968, 
    9.970427,
  5.777046, 4.174219, 5.486395, 21.59912, 1.618877, 12.08853, 22.05826, 
    13.98775, 10.45017, 23.61456, 11.16404, 3.598372, 3.995757, 4.116332, 
    3.913164, 3.77073, 3.530632, 3.539215, 3.53737, 11.28327, 21.37163, 
    18.62497, 16.01394, 4.823305, 3.517333, 3.467555, 3.608656, 3.533894, 
    4.869901,
  4.382843, 15.4181, 18.35289, 23.70248, 25.53226, 25.93858, 12.38102, 
    25.60696, 11.6648, 6.162197, 7.399197, 17.98231, 3.534197, 3.714916, 
    3.496224, 3.35418, 3.230659, 3.376678, 3.683931, 18.60765, 17.19287, 
    22.69472, 17.91301, 21.58281, 8.053755, 3.431259, 3.719141, 3.554709, 
    3.53227,
  3.182451, 13.19842, 9.963753, 14.51696, 13.98608, 14.89089, 15.30038, 
    15.69397, 12.94773, 13.23608, 11.35011, 20.72614, 21.59224, 17.33226, 
    2.292719, 19.75172, 18.21741, 9.211101, 20.85629, 13.01678, 14.92194, 
    21.52704, 25.92181, 21.60022, 2.318715, 5.825578, 3.04392, 3.010769, 
    3.157359,
  0.2291971, 0.2093325, 1.794062, 0.2354309, 1.202312, 2.970822, 2.57245, 
    2.555763, 2.463318, 2.390499, 1.640874, 1.384348, 2.465297, 3.075774, 
    3.047408, 3.295175, 2.816517, 3.135645, 3.215559, 3.319413, 2.739849, 
    3.048805, 2.885937, 2.84402, 3.00572, 2.61534, 2.674233, 3.028145, 
    0.2641115,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 average_DT = 732 ;

 average_T1 = 14.5 ;

 average_T2 = 746.5 ;

 climatology_bounds =
  14.5, 746.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
