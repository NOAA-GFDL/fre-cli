netcdf atmos.1980-1981.aliq.07 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:20 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.07.nc reduced/atmos.1980-1981.aliq.07.nc\n",
			"Mon Aug 25 14:40:45 2025: cdo -O -s -select,month=7 merged_output.nc monthly_nc_files/all_years.7.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.042865e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.14169e-05, 0.0002174616, 0, 0, 9.671025e-05, 
    2.206927e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.563109e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.290004e-05, 0, -8.717577e-07, 0, 0, 0, 
    0, 0, 0, 0, -6.191454e-05, -8.044475e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0002057924, 0.000278531, 0, 0, 0.003914091, 
    0.0009706871, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.674693e-05, 0.0007964445, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0003302352, 0, 0, 0, 0, 0, -7.08744e-05, 
    1.450145e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005650484, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002212147, 0.0001461699, -7.165509e-06, 
    -1.410502e-06, 0, 0.000295075, 0, -1.713409e-06, -5.506641e-06, 
    0.001348513, 0.001516916, -3.153511e-05, -3.301977e-06, -1.845552e-06, 0, 
    0, -1.568488e-06, 0,
  0, 0, 0, 0, 0, 0, 0.002031098, 0.000545153, -1.211383e-05, -1.229883e-05, 
    0.008935427, 0.002444368, -2.438964e-05, -3.74793e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.00032104, -3.233964e-06, -2.405073e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0004054964, 0.001762367, 0, 0, 5.992272e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001214283, 0, 0, -2.362696e-06, 0, -9.748767e-05, 
    -8.50537e-05, 8.05308e-06, -2.87564e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.714786e-05, -2.706246e-05, 
    0.001494696, -5.922289e-07, 0, 0, 0, 0, 0, 0, 0, -2.042299e-06, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001341, 0.0007947416, 0.001663189, 
    -1.957942e-05, 3.418433e-05, 0.001120231, -2.414499e-05, 0.000197568, 
    0.001265509, 0.003590584, 0.005677114, 0.0001130651, -3.301977e-06, 
    -8.978092e-06, -2.002543e-05, 0, 0.0002874371, 0.0009082346,
  0, 0, 0, 0, 0, 0, 0.006604519, 0.001330235, -2.951023e-05, 0.0002682989, 
    0.0122637, 0.005341358, 0.0004812803, 0.0002187607, 0, 0, 0, 0, 0, 0, 
    8.943747e-06, -1.785749e-05, 0, 0.0014205, -3.171126e-05, -8.631425e-05, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0005228667, 0.002602359, 0.0004385535, 
    -4.596034e-06, 2.603378e-05, 5.836523e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.85539e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.315446e-09, -6.286011e-05, 
    7.549522e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.376665e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.88984e-05, 0.001810766, -2.363412e-08, 0, 
    -3.239385e-05, 0, 0.0002446509, 0.0002146518, 0.001148935, 3.073598e-05, 
    -1.651882e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.277429e-05, 0, 0, 0, 0.0001760165, 0, -6.221958e-06, 
    -6.589696e-05, 0.0001108027, 0.004046161, -2.543085e-06, 0, 0, 0, 0, 0, 
    0, 0, 3.914754e-06, -4.36032e-06, 0, 0, 0, 0,
  3.802986e-08, 0, 0, -3.473799e-06, 0.0001015363, 0, 0, 0, 0, 0, 
    -8.338725e-06, 0.004232185, 0.002354499, 0.00235177, 0.0008051826, 
    0.0001902686, 0.002235902, 0.0004907572, 0.002124538, 0.004674288, 
    0.01146017, 0.01071759, 0.0001490593, 1.279115e-05, -1.959777e-05, 
    -4.387437e-05, 0.0002645866, 0.001067834, 0.002003494,
  0, 0, 0, 0, 0, 0.0004819388, 0.01456144, 0.001973583, 0.003242921, 
    0.0004315528, 0.0180464, 0.02043881, 0.002141035, 0.001946884, 0, 0, 0, 
    0, 0, 0, -3.201408e-05, 9.15803e-05, 0, 0.00371428, 0.0001310873, 
    0.0001428996, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0003377347, 0.0004510008, 0.004060395, 0.001374474, 
    0.0001505245, 0.0008798485, -4.049019e-05, 2.465592e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, -0.0001414457, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 7.618605e-06, 3.069614e-05, -1.443464e-06, 
    -5.717968e-05, 0.004177857, -2.452255e-05, 0, 0, 0, 0, 0, 0, 0, 
    -4.590036e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.100136e-05, 0, 3.531179e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002806922, 0, -6.002761e-06, 0, 
    -5.927074e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -0.000173413, 0.0033914, -1.894591e-05, 0, 0.0003415882, 
    0, 0.002477495, 0.007372499, 0.00378151, 0.0002464106, -1.865174e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -1.916143e-05, 1.070896e-05, 0, 1.060849e-06, 0.0008614543, 
    0.0001057378, 0.0004071752, 0.001024187, 0.001474513, 0.005949374, 
    -8.687126e-06, -1.2133e-05, 0, 0, 0, 0, 0, 0, 0.000286271, 0.001461406, 
    0, 0, 0, 0,
  2.66209e-07, 6.880243e-05, 0.0002293793, 8.536089e-06, 0.0009223546, 0, 0, 
    0, 0, -1.055622e-05, -2.640045e-05, 0.005946078, 0.006771182, 
    0.005820174, 0.00157749, 0.002593797, 0.003810497, 0.001827473, 
    0.005947665, 0.009452061, 0.01879018, 0.02123219, 0.001977218, 
    7.142073e-05, -8.580888e-05, 2.15542e-05, 0.0007698997, 0.005676501, 
    0.003588377,
  0, 0, 0, 0, 0, 0.001744475, 0.03552606, 0.005670489, 0.008907091, 
    0.0005525252, 0.03285544, 0.03250228, 0.005815929, 0.004826608, 
    -1.484502e-06, 0, 0, 0, 0, 0, -5.321267e-05, 3.896144e-05, -3.920994e-06, 
    0.006803628, 0.001115009, 9.931997e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001160163, 0.001803152, 0.007870058, 0.003111881, 
    0.002421064, 0.001492545, 0.002879168, 0.0003926068, 2.363508e-05, 0, 0, 
    0, 0, 0, -1.057266e-05, 0, 0.0003508579, 0.0004177338, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -4.95171e-06, 3.695745e-05, 0.0004255738, 
    0.0004678345, 0.0028191, 0.01087604, 0.0006164719, 0, 0, 0, 0, 0, 0, 0, 
    -4.648586e-05, 0, 7.120526e-05, -8.214992e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.340193e-07, 0.0001265152, -8.776909e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, -7.51314e-05, -7.868918e-05, -2.054234e-06, 
    0.0009947388, -3.025021e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.113492e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006117517, 0, 
    -2.281578e-06, 0.0001356163, 0, 0, 0, -8.040124e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006509593, 0.0009404657, 
    0.0001086226, -2.716591e-06, 0.0003078216, 0.0006400673, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.973069e-05, -7.310974e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -7.172145e-06, 0, 0.0003667988, 0.007991324, 0.0002234535, 0, 
    0.001212536, 0, 0.009607683, 0.01667215, 0.007375147, 0.0009190114, 
    -2.834656e-05, 0, 0, 0, 0, -1.726053e-07, 0, 0, 0, 0, 0, 0, 0,
  0, -1.452382e-05, 0, 0, 0, -2.183355e-05, 0.0004965828, -4.062229e-06, 
    -1.562539e-05, 0.002344878, 0.0005123473, 0.001979418, 0.004783015, 
    0.004967131, 0.009058979, -1.421398e-05, 0.0001214932, 0, 0, 0, 0, 0, 0, 
    0.001334428, 0.003125983, 0, -7.805151e-07, 0, 0,
  0.0003009647, 0.0008915986, 0.001024054, 0.0003750134, 0.002877127, 0, 
    -9.456273e-06, -6.337397e-05, -1.190184e-05, 4.50131e-05, 0.002430442, 
    0.009499371, 0.01291563, 0.01243127, 0.00300892, 0.00922688, 0.005613009, 
    0.003541067, 0.01415277, 0.01742123, 0.03176686, 0.04012796, 0.004376691, 
    0.0001231755, -0.0001737954, 0.00340592, 0.002397852, 0.01569436, 
    0.005690323,
  0, 0, 0, 0, 0, 0.007252417, 0.07359058, 0.01297813, 0.01987286, 
    0.002748789, 0.05157956, 0.04426027, 0.01406812, 0.007517328, 
    -2.36886e-06, 0, 0, 0, 0, 0, -7.116325e-05, 0.0001203893, -3.300871e-05, 
    0.00794055, 0.005192174, 0.0004110728, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.004629708, 0.005119617, 0.01554258, 0.006708182, 
    0.005580394, 0.004639178, 0.01305045, 0.005976119, 0.0008896057, 0, 0, 0, 
    0, 0, 5.040626e-05, 0.0001823883, 0.001651724, 0.00212872, -2.09078e-07, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.789595e-08, 0, -1.879142e-05, 0.001504803, 
    0.003837873, 0.006298817, 0.009442942, 0.01930915, 0.00595978, 
    -9.1222e-06, 0, 0, 0, 0, -1.640447e-06, 9.969297e-05, 0.0005683635, 
    0.001324518, 0.0004788945, 0.001979081, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.107116e-05, -5.169139e-05, 0.001885363, 
    0.0007958956, -1.043699e-05, 0, 1.1278e-05, 0, -9.778946e-06, 0, 0, 0, 
    0.002573316, 0.001772131, 0.001350754, 0.002822095, 0.0008085587, 
    2.583616e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.350323e-06, -6.980945e-07, 7.039635e-05, 
    -4.978662e-06, 0.0003467565, -7.620302e-06, 0, 0, 0, 0, 0, -8.413544e-07, 
    0, 0, -2.976361e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.64654e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.187965e-05, 0, 
    0, 0, 0, 0, 0, 0, 0.0001614072, 0.0001341614,
  0, 0, -1.197217e-07, -2.00977e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.714749e-05, 0.002298275, 0.0006521074, 0.000739628, 0.0003704757, 
    -1.396022e-05, 0, 0, 0.002156554, 0.002852474, 0.0001864331, 
    -6.650655e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009562567, 0.006288419, 
    0.00310885, 0.001750595, 0.002066448, 0.001039893, 0, 0, 0, 0, 0, 
    0.0005188785, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004248001, -3.142604e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -5.290869e-06, 0, 0.002997832, 0.0192877, 0.0007127417, 
    -1.151399e-05, 0.004192902, -1.226898e-05, 0.02278663, 0.03636467, 
    0.01528757, 0.001305192, 0.0003913852, 0, 0, 0, 0, -9.301289e-08, 0, 0, 
    0, 0, -2.446036e-10, 0, 0,
  0, 0.001086927, -4.053749e-06, 0, 0, -2.622903e-05, 0.0005042507, 
    2.95676e-05, 0.0001948784, 0.00420067, 0.002694808, 0.004986219, 
    0.01055675, 0.01143786, 0.01386278, -7.304799e-05, 0.001330993, 0, 0, 0, 
    0, 3.588004e-05, 0, 0.002758128, 0.00460267, -8.380637e-06, 
    -1.322668e-05, 0, 0,
  0.001624572, 0.002605075, 0.002344028, 0.003985788, 0.004889764, 0, 
    0.0005876389, 0.001605265, 0.0006144782, 0.001318303, 0.005048967, 
    0.01878406, 0.03067585, 0.02100133, 0.009599534, 0.01657227, 0.008382753, 
    0.007953994, 0.02468136, 0.02761712, 0.0604789, 0.06784558, 0.01614506, 
    0.0005095463, 0.0008448175, 0.01580267, 0.007335678, 0.0399208, 0.0123679,
  0, 0, 0, 5.065938e-07, -5.845307e-06, 0.01432447, 0.1083614, 0.02724765, 
    0.05608778, 0.006888941, 0.07883459, 0.07086243, 0.03094684, 0.02051022, 
    -7.476007e-06, 0, -1.934523e-05, 0, 0, 0, 0.002403128, 0.002141034, 
    -0.0001651559, 0.01470605, 0.006423547, 0.001135381, -1.361631e-05, 0, 0,
  0, 0, 0, 0, 0, -3.382936e-06, 0.01798551, 0.01004199, 0.03170244, 
    0.01429753, 0.01149302, 0.01341972, 0.02980011, 0.01706952, 0.00190772, 
    -2.707593e-06, 0, 0, 0, 0, 0.0002027742, 0.000780435, 0.008713607, 
    0.004982264, -9.066207e-07, -2.272608e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -3.762812e-06, 0, 0.002811561, 0.00570175, 0.01503225, 
    0.01397161, 0.02305653, 0.03246209, 0.02482844, 0.002219825, 
    0.0005637998, 0, 0, 0, -9.24807e-06, 0.001134434, 0.0015524, 0.005036299, 
    0.003340776, 0.003346708, 0, 0, 0,
  0, 2.061347e-06, 1.99889e-05, 0, 0, 0.0001547013, 0, -2.790271e-06, 
    -2.490407e-06, 0.0001116369, -8.315493e-05, 0.005436814, 0.007058877, 
    0.004513328, 0.0009900375, 0.0007023175, -6.460346e-07, 0.0009225652, 0, 
    0, 2.555996e-05, 0.004366495, 0.006071773, 0.003255639, 0.0101286, 
    0.00397719, 0.002470965, 0.0009923981, -2.514404e-06,
  0.0001342052, 1.342808e-06, -4.965572e-06, 0, 0, -6.505151e-05, 
    0.001168621, -2.060193e-05, 0, 4.161801e-05, 0.0005192992, 0.003909314, 
    0.003057671, 0.001422803, -1.297473e-06, -2.300558e-05, -3.718662e-09, 0, 
    0, 0, -7.898732e-05, 0, -6.492381e-05, 2.829024e-05, 0, -5.299964e-05, 0, 
    -2.207292e-10, 0,
  0, 0, 0, -1.763724e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.496457e-09, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.995591e-11, -5.74138e-10, 2.575797e-09, -6.768711e-10, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007460956, 0, 0, 0, 0, 0,
  8.813942e-05, -4.832367e-05, 0, -9.655412e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001341234, 0, 0, -5.930007e-06, 0, 0, 0.0008550425, 0.0004273214, 0, 
    1.287867e-05, 0, 0, -9.037097e-07, 0, 0.0018067, 0.0002372755,
  0, 0, -1.302795e-05, 0.0008329189, -1.004748e-05, -1.613083e-05, 0, 
    6.151332e-05, 0, 0, 0, 0, 0, 0.0004269457, 5.589493e-05, 0, 0.0001551441, 
    0.006861486, 0.001325416, 0.00875521, 0.00422202, 3.317712e-05, 
    0.0006393724, 0, 0.003225911, 0.004517945, 0.003070299, -0.0001022334, 
    -2.049948e-05,
  0, 0, 0, 0, 0, 0, 0, 0, -2.432174e-12, 0, 0, 0, 0, -2.110781e-06, 
    0.0108791, 0.02082366, 0.0114587, 0.004391385, 0.008365177, 0.002373931, 
    -1.303542e-05, 0, 0, 0, -2.464444e-05, 0.001208917, 0, 7.960683e-06, 0,
  0, 0, 0, -9.436186e-16, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002146822, 0.006584258, 
    0.0001577196, 0.00203273, 0.0003023605, -1.0369e-06, 0, 0, 0, 
    1.712505e-06, -2.221376e-10, 0.0002778529, 0, 0, 0, 9.60583e-08, 0,
  8.910928e-08, 0, 0, 0, 7.364197e-07, 0, 0.01146825, 0.03390461, 
    0.0009514007, -0.0002572888, 0.006912654, 0.003216957, 0.03651855, 
    0.06407318, 0.02887735, 0.002488381, 0.001897347, 0, 0, 0, -1.329025e-08, 
    1.443493e-08, -1.959051e-08, 0.0002096659, -6.727406e-08, 1.876302e-07, 
    7.920247e-09, 0, 0,
  -5.39801e-06, 0.002246014, -3.185392e-05, 9.938739e-08, -1.52117e-07, 
    0.0006789266, 0.001354216, 0.005483734, 0.002820433, 0.01969778, 
    0.01067369, 0.01461714, 0.02653721, 0.0308883, 0.02635444, 0.000422719, 
    0.001965287, 0, -2.938046e-05, -8.212532e-06, -5.74021e-08, 0.0008272784, 
    8.008527e-06, 0.01299693, 0.006052955, -0.0001001759, -3.939915e-05, 
    -3.286425e-10, -3.068914e-06,
  0.006651675, 0.00506688, 0.005893505, 0.01119093, 0.005740895, 
    4.199039e-05, 0.006654176, 0.007493297, 0.005203538, 0.008238588, 
    0.01315912, 0.04201819, 0.08934345, 0.05137691, 0.0292736, 0.03044757, 
    0.01303999, 0.01854827, 0.03903248, 0.041097, 0.1091787, 0.1002933, 
    0.04888634, 0.002190907, 0.006167803, 0.03217467, 0.0154721, 0.08113177, 
    0.0226282,
  0, 0, 0.0001419577, 0.001060367, 0.002304031, 0.07729661, 0.1635588, 
    0.1283728, 0.108424, 0.02825769, 0.1326261, 0.1112225, 0.07627457, 
    0.03923559, -2.160122e-05, -6.092153e-06, 0.0002788392, 0.003283786, 0, 
    -2.280464e-06, 0.0075294, 0.005796602, 0.0001653979, 0.02716236, 
    0.01115506, 0.002435572, -5.694148e-05, -7.138735e-07, 0,
  0, -3.087324e-07, 0, 6.037151e-07, -5.860164e-07, -8.094568e-05, 0.1060356, 
    0.01917016, 0.04162766, 0.08749091, 0.02603539, 0.0289721, 0.07479163, 
    0.03280514, 0.007947892, 0.0001503002, 0, 0, 0, 0, 0.0001286571, 
    0.006890347, 0.03968597, 0.01887384, 5.505677e-05, -2.330791e-05, 0, 0, 
    -4.304673e-05,
  0.0001382618, 3.436211e-06, -3.70105e-05, 0, 2.611734e-08, 2.472897e-05, 
    -1.279504e-05, 0.0001309441, 0.01301252, 0.02043656, 0.03843059, 
    0.02846799, 0.04133474, 0.06313003, 0.0418369, 0.005946877, 0.0008589436, 
    0, 0, 0, 0.0005922277, 0.002657581, 0.008420737, 0.006334969, 
    0.007183865, 0.007213855, 0.0001656738, 0, 0,
  0, 0.002490385, 0.001209971, 0.0005400336, -3.579367e-07, 0.0003426599, 
    -1.350303e-05, 0.0004595585, 0.001145843, 0.006593545, 0.005133559, 
    0.02508195, 0.0291125, 0.01488639, 0.004886124, 0.002295123, 0.002624078, 
    0.004151889, -1.311019e-05, 0, 0.004107319, 0.01140983, 0.01245848, 
    0.009993761, 0.02551407, 0.01189699, 0.006255579, 0.006837527, 
    0.0007304594,
  0.00227289, 0.002797447, -0.0001014591, 0, -4.525179e-05, -0.000155842, 
    0.002373523, 0.00106445, 0.001402219, 0.005215679, 0.003983235, 
    0.01250526, 0.0119764, 0.007569133, 0.0002841645, 0.0007183565, 
    0.0002398825, 0, 0, -3.735501e-06, 0.0006398535, -7.365835e-05, 
    0.003095913, 0.003871871, 0.0006155382, 0.001117721, 0.000934338, 
    -7.172301e-05, 0.000257994,
  0, -1.721551e-08, -2.141534e-07, -6.605409e-05, -3.963133e-05, 0, 0, 
    -1.310106e-06, 0.0013287, 0.000361806, 0, -1.213836e-05, 0, 
    -2.194041e-06, -1.178843e-05, 0, 0, 0, 0, 0, -6.07627e-05, 0, 
    -1.067229e-05, -1.334968e-09, 0, 0, 0, 0, -2.249507e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.575391e-10, 2.504508e-08, -3.5734e-09, 1.436236e-08, -2.041872e-11, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -8.308972e-06, 0, 0, 0, -6.26096e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, -2.399026e-05, 0.001831291, 0, 0, 0, 0, 0,
  0.001655562, 0.003953089, -1.34411e-06, 0.0006223925, 6.416717e-06, 
    9.527868e-06, -5.088737e-07, 0, -1.03913e-05, 1.147094e-05, 0, 0, 
    -1.651893e-06, 0.002382146, 0, 0, 3.501814e-06, 0, -5.748501e-05, 
    0.001293035, 0.001636283, -1.205631e-05, 0.001093006, 0.000438376, 0, 
    0.0005366502, 0, 0.003280474, 0.000303792,
  -3.062185e-05, 0.0001171097, -2.774235e-06, 0.003235605, 0.005052592, 
    -8.339203e-05, -4.145773e-05, 0.004348115, 1.341504e-05, -1.067076e-10, 
    0, -3.048607e-06, -2.419119e-07, 0.0042527, 0.001508145, 6.881854e-05, 
    0.002700349, 0.01734495, 0.009453045, 0.0284178, 0.01764, 0.001505417, 
    0.001202624, -4.061956e-06, 0.004654965, 0.005971954, 0.005321162, 
    0.0005678314, 0.002937641,
  0.001267885, 0, 0, -3.629683e-09, -8.524652e-05, -2.242337e-07, 
    0.0005330939, -1.049667e-09, -2.011948e-06, 7.630035e-08, 1.347384e-09, 
    -6.223316e-10, 0, -6.79548e-07, 0.02119687, 0.04632029, 0.0343285, 
    0.01649027, 0.02467354, 0.008119322, 0.0008320215, 0, 7.844537e-06, 0, 
    0.0004070526, 0.001911339, 7.362396e-06, 0.003974207, 1.582564e-05,
  2.769379e-06, 1.532077e-08, 0, 4.40767e-07, 1.278546e-10, 8.760138e-09, 
    2.941099e-07, 4.67178e-05, 5.993727e-07, 1.090618e-07, 3.8936e-07, 
    1.516317e-07, 0.001235574, 0.01611599, 0.006539126, 0.01318996, 
    0.006664777, 0.0002630148, 0.0005129638, 0, 4.926871e-08, 0.0003385563, 
    3.943108e-06, 0.001839662, -2.383113e-08, -1.405322e-08, 1.948979e-05, 
    1.68422e-06, -1.544689e-07,
  5.708597e-05, -3.244362e-08, -1.945391e-07, -1.432496e-10, 1.891979e-05, 
    2.330072e-06, 0.01911929, 0.06925245, 0.004280049, 0.002079401, 
    0.01067837, 0.01448574, 0.07661353, 0.1526504, 0.0935324, 0.002882918, 
    0.004873707, 4.572528e-09, 0, -7.759779e-07, -2.957424e-05, 0.0005630174, 
    4.145474e-06, 4.84936e-05, 0.0001367413, 0.0005008677, -1.33679e-06, 
    9.906134e-07, 4.089867e-10,
  4.803451e-05, 0.008298069, 0.003556645, 8.864271e-05, 1.951858e-06, 
    0.005346623, 0.009197464, 0.04738216, 0.02098211, 0.04408241, 0.138714, 
    0.189578, 0.1274351, 0.1256702, 0.1079396, 0.008338834, 0.004449231, 
    6.45687e-06, 0.000684322, 0.004482933, 0.0004530899, 0.01243693, 
    0.002534969, 0.03046601, 0.00953877, -0.0001909571, 0.0006863778, 
    6.051014e-05, 3.518265e-05,
  0.03507414, 0.02137944, 0.01820171, 0.017347, 0.00942058, 0.01034272, 
    0.1403853, 0.4755185, 0.3163919, 0.2862403, 0.2884165, 0.2665741, 
    0.2766127, 0.1996759, 0.1798421, 0.09219356, 0.02770792, 0.06327265, 
    0.1021316, 0.1088952, 0.2238213, 0.2064275, 0.1244337, 0.02492678, 
    0.01663965, 0.0508384, 0.02734219, 0.1330278, 0.04982948,
  7.145073e-06, 7.497082e-05, 0.003018631, 0.02415921, 0.1488185, 0.2226626, 
    0.3467355, 0.2037865, 0.407563, 0.1418154, 0.2939636, 0.2188496, 
    0.2672575, 0.07650203, 0.001347469, 0.000858288, 0.0008048999, 
    0.006276333, -2.215897e-06, 0.003298461, 0.07900404, 0.05635068, 
    0.01524654, 0.06807892, 0.01911158, 0.00815913, 7.484431e-06, 
    -1.071497e-06, 3.839234e-05,
  -1.402299e-11, -3.452368e-05, -1.692578e-09, 8.162933e-06, 0.0006159482, 
    0.001528254, 0.0855069, 0.03542106, 0.05973918, 0.1227659, 0.09245878, 
    0.1497235, 0.2527722, 0.1105756, 0.02566755, 0.009636817, 0.0002299446, 
    0.0001891538, -1.005565e-07, 7.580133e-05, 0.003422612, 0.0676586, 
    0.2291006, 0.08709215, 0.001580036, 6.761027e-05, 5.936694e-08, 
    -6.916898e-12, 0.001200552,
  0.0001073186, 0.001585272, 0.0001581021, -7.038567e-11, 1.276977e-07, 
    0.0005913541, 0.0003027614, 0.003853576, 0.06693913, 0.07462867, 
    0.1412001, 0.1110356, 0.1326359, 0.1169098, 0.08107898, 0.02931182, 
    0.005198834, 0.0004861745, 4.683342e-06, 0, 0.0006098609, 0.004890861, 
    0.01943904, 0.04281087, 0.02238409, 0.01181877, 0.00108658, 0.0003613764, 0,
  0.0005835337, 0.005984727, 0.002184806, 0.002665151, 3.760034e-05, 
    0.002439927, 0.0001937294, 0.005679505, 0.007370527, 0.0151464, 
    0.01961194, 0.06532647, 0.07863101, 0.04585911, 0.02690718, 0.007612301, 
    0.0071974, 0.01027498, 0.000973461, -4.20962e-06, 0.0104658, 0.02079579, 
    0.0199308, 0.01831521, 0.03792486, 0.02908697, 0.01605522, 0.01746776, 
    0.007152782,
  0.003155277, 0.004348753, 0.001958152, -5.118825e-06, 0.005634849, 
    0.005752666, 0.002512617, 0.009558599, 0.002669078, 0.01442576, 
    0.0119003, 0.02087671, 0.02510259, 0.01824756, 0.001487015, 0.001381606, 
    0.0005808946, 0, -4.104474e-05, 0.0001044498, 0.001212495, -0.0001660755, 
    0.006867419, 0.006868603, 0.003196628, 0.005056498, 0.005024679, 
    -0.0002156385, 0.008215768,
  0, -3.915803e-05, 0.0002152054, 0.00104985, 0.0002578562, -3.554713e-05, 
    7.057758e-05, 1.525234e-05, 0.002743996, 0.002116773, 3.638463e-06, 
    -2.12197e-05, -0.000163387, 1.455382e-05, 0.001115068, 0, 0, 0, 0, 0, 
    0.003554909, 0.0002534407, 0.0002359252, -1.491254e-05, 0, 0, 
    -1.583365e-06, -1.430629e-07, 0.0009580054,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 7.244054e-05, -1.04082e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -9.679101e-10, -5.089254e-08, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.400641e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -2.626045e-06, 0, 0, 0, 0, 0, -1.822016e-05, 0, -9.743692e-07, 0, 
    0.001007401, 0, 0.0003163591, -6.280727e-06, 0, 0, 0, 0, 0.0001944956, 
    0.003927839, 0.002291018, 0, 0.0004915371, -1.738005e-05, 0, -1.207506e-05,
  0.004788903, 0.009059186, 0.001346584, 0.003667003, 0.000134198, 
    0.002927016, 0.000602821, 0.0001961402, 0.001853818, 9.389681e-05, 
    1.214508e-05, 0.001517288, 0.001354277, 0.002508914, 0.0002393679, 
    -9.938448e-07, 0.0002458939, 3.010254e-05, 2.813068e-06, 0.003859356, 
    0.00675564, 0.0002151956, 0.004365857, 0.003199892, -2.009421e-05, 
    0.001656398, 4.310601e-06, 0.006886885, 0.002471224,
  0.005828133, 0.002665039, 0.002135252, 0.01148063, 0.0154343, 0.004259714, 
    0.004602168, 0.006849497, 0.0003331178, 2.090429e-06, 6.682814e-06, 
    -2.778631e-05, -1.530697e-05, 0.007670629, 0.007106963, 0.004185842, 
    0.01124558, 0.03460545, 0.02821187, 0.05105633, 0.04496748, 0.007863783, 
    0.005551655, 0.0008397257, 0.008642305, 0.006429264, 0.01065719, 
    0.005462546, 0.01077955,
  0.008672691, -1.375937e-06, 0.000375606, -8.959505e-08, -3.785461e-05, 
    -2.527836e-05, 0.004770546, 1.939133e-09, 1.898735e-05, 1.560792e-06, 
    4.016706e-06, 7.192319e-07, -1.210444e-08, -3.399436e-05, 0.04838613, 
    0.09459995, 0.07564158, 0.03812678, 0.06059981, 0.02374264, 0.003606681, 
    0.0001018925, 0.0001148161, 0.002732865, 0.002984298, 0.005486303, 
    0.0004376764, 0.01235612, 0.004077171,
  0.0001192083, 0.0007678564, 6.021565e-07, 2.207773e-07, -6.401683e-10, 
    -4.930973e-09, 0.002669323, 0.0009842897, 6.990565e-06, 1.346976e-06, 
    1.664481e-07, 1.086051e-06, 0.000736835, 0.04064226, 0.05673041, 
    0.06278337, 0.03573848, 0.01192611, 0.004994019, -3.341746e-06, 
    4.034966e-06, 0.004017833, 0.00284252, 0.005601242, 0.007614671, 
    -1.886871e-06, 0.002420345, 0.0003141085, 1.251704e-05,
  0.003647159, 0.003777598, 2.042984e-05, 2.984138e-06, 0.007810032, 
    0.0008964139, 0.0815233, 0.1364973, 0.008876456, 0.007945781, 0.01872878, 
    0.01652641, 0.1108343, 0.1736249, 0.1167991, 0.01888677, 0.005530469, 
    -2.200916e-07, 1.291365e-06, 0.0001402685, 4.548611e-05, 0.0120321, 
    0.002135442, 0.0201796, 0.01016324, 0.008095901, 0.0002053918, 
    0.01434222, 0.008096231,
  0.02429298, 0.1684594, 0.1825007, 0.009088731, 0.005855308, 0.06183746, 
    0.1971777, 0.3605706, 0.2312721, 0.3139062, 0.1682893, 0.2000023, 
    0.1476421, 0.1130748, 0.1012533, 0.008053499, 0.005151524, 4.150726e-06, 
    0.0005782729, 0.03118628, 0.03315915, 0.06002855, 0.06790195, 0.1235894, 
    0.05014904, 0.005646378, 0.01230174, 0.0590499, 0.01633343,
  0.2922158, 0.3377678, 0.2877882, 0.02855618, 0.03332871, 0.05303549, 
    0.2166793, 0.45044, 0.2736512, 0.2185354, 0.2094879, 0.20182, 0.2447332, 
    0.1712582, 0.2256881, 0.1292526, 0.04566692, 0.08525133, 0.1241229, 
    0.1306275, 0.2940974, 0.3001851, 0.3877894, 0.1564534, 0.07804964, 
    0.1364319, 0.09171156, 0.3035238, 0.3322824,
  0.00116377, 0.004107594, 0.003106149, 0.02251463, 0.1219658, 0.2286204, 
    0.3293077, 0.1623473, 0.3872202, 0.1113594, 0.2516027, 0.1745959, 
    0.2417271, 0.1320059, 0.1345406, 0.08829056, 0.02863204, 0.04971455, 
    0.001594009, 0.008099865, 0.05298038, 0.07254082, 0.06112275, 0.1152504, 
    0.1607387, 0.02182214, 0.001346528, 0.009446051, 0.001251092,
  0.0008037722, 0.0006173566, -1.215069e-09, 3.494052e-06, 0.007648748, 
    0.001933194, 0.06535042, 0.06578176, 0.1192202, 0.09880877, 0.07134447, 
    0.112611, 0.2716394, 0.2532273, 0.1438609, 0.02700405, 0.03947997, 
    0.01136488, 0.001798436, 0.003105948, 0.04694915, 0.1315576, 0.2641262, 
    0.2548881, 0.110984, 0.06367379, 0.0007217069, 0.001077053, 0.006221463,
  0.006026896, 0.007886974, 0.001271943, -6.425614e-08, -5.712026e-06, 
    0.001571365, 0.005736989, 0.0357402, 0.1106663, 0.1685139, 0.2379559, 
    0.1801392, 0.2353748, 0.2281887, 0.1744079, 0.1246133, 0.04885752, 
    0.04409197, 0.0179362, -8.420746e-06, 0.001496347, 0.08120784, 
    0.09293795, 0.1418988, 0.1512481, 0.1034946, 0.04219967, 0.01575326, 
    0.004164849,
  0.004789652, 0.01127206, 0.003258537, 0.007750347, 0.01536512, 0.01358046, 
    0.003504514, 0.009338576, 0.01374291, 0.03541286, 0.07945684, 0.1806821, 
    0.1558522, 0.1287375, 0.1311354, 0.09734234, 0.060629, 0.06307478, 
    0.03778145, 0.002124125, 0.01380826, 0.03795642, 0.03631165, 0.06076452, 
    0.08768018, 0.09419377, 0.07938744, 0.05411311, 0.02711997,
  0.004576619, 0.006868324, 0.006088446, 0.0002738221, 0.008986139, 
    0.008621179, 0.0123956, 0.04541197, 0.01154567, 0.02708365, 0.02848303, 
    0.04850394, 0.09047659, 0.08210651, 0.05608903, 0.02451814, 0.003334703, 
    -7.03658e-05, 0.001324333, 0.002709911, 0.004532669, 1.714285e-05, 
    0.01322027, 0.01035417, 0.03279787, 0.04066169, 0.03653245, 0.01528392, 
    0.01627695,
  -2.71159e-05, 0.001779318, 0.003280469, 0.004812398, 0.002907123, 
    0.000485532, 0.001883007, 0.002101545, 0.006256962, 0.008043229, 
    0.001352863, 0.000815912, 0.003599107, 0.01297812, 0.01470327, 
    0.001891373, -1.770319e-06, -4.959854e-09, -9.713571e-06, -5.535185e-07, 
    0.007153322, 0.001134695, 0.005313477, 0.00273633, -4.242378e-06, 0, 
    0.0002851218, 0.0004997056, 0.004471381,
  0, -3.13185e-07, 1.689302e-09, -0.0001714009, -1.175641e-05, 0, 0, 0, 
    -0.0002829951, 0.002457238, -6.944782e-05, 0, 0.0006612365, 
    -7.725492e-05, 1.18893e-09, -2.099207e-06, -1.446153e-06, 0, 0, 0, 0, 0, 
    0, -2.39016e-11, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.39855e-05, 0.001088511, 
    7.710509e-05, 0, 0, -5.1587e-07, 0, 0, 0.001237049, 0, -1.577744e-05, 0, 
    0, 0, 0, 0,
  -3.891027e-05, -2.612129e-07, -1.805557e-06, -1.436217e-05, 0, 0, 0, 
    -2.82579e-07, 0.0004987018, -4.826985e-05, 1.324242e-05, -8.024642e-05, 
    0, 0.002374047, 2.19031e-05, 0.001030604, 3.487838e-05, -1.850502e-05, 0, 
    -5.343647e-06, 0, 0.0003739401, 0.006746653, 0.007672711, -2.833116e-05, 
    0.0008339604, -2.116105e-05, 0, -2.730983e-05,
  0.01869279, 0.01775694, 0.003235077, 0.01030532, 0.002673938, 0.007228161, 
    0.002585596, 0.001421734, 0.006478776, 0.005660953, 0.00622792, 
    0.002095271, 0.003891883, 0.002851375, 0.00941828, -4.666909e-05, 
    0.002996044, 0.001414054, 0.004277316, 0.006477721, 0.0134061, 
    0.009179283, 0.01629511, 0.01086044, 0.0004531132, 0.002876729, 
    0.0007391346, 0.01137531, 0.01292534,
  0.01597201, 0.003038295, 0.006131168, 0.01666188, 0.02431298, 0.01595872, 
    0.01013901, 0.01121149, 0.005339283, 0.005843593, 0.00177404, 
    0.0004807478, -0.0001124332, 0.01264163, 0.02310897, 0.02079891, 
    0.03500167, 0.06038389, 0.06204773, 0.09122105, 0.07946281, 0.03084754, 
    0.02452083, 0.008047654, 0.01910073, 0.01267732, 0.01993518, 0.0195528, 
    0.02443035,
  0.003059743, 0.0007811545, 0.0009426296, 3.629416e-05, 0.000680354, 
    0.001535772, 0.008488985, -2.067966e-06, 0.00364446, 0.0002999617, 
    0.0004494278, 0.0007959896, -4.034178e-05, 0.001124126, 0.08177689, 
    0.1306605, 0.1385692, 0.1398022, 0.1553511, 0.1192917, 0.07687593, 
    0.03152527, 0.007756012, 0.0006873634, 0.00976475, 0.01814296, 
    0.009270286, 0.02546558, 0.008786133,
  2.806878e-06, 7.563363e-05, 2.077343e-06, 0.000111438, -1.023866e-08, 
    6.286524e-10, 0.0002950955, 0.0005066872, 6.855903e-07, 8.524673e-07, 
    1.667933e-07, 5.514636e-07, 6.104411e-06, 0.04586735, 0.05444035, 
    0.09063374, 0.04293602, 0.02167817, 0.009075576, 0.001601907, 
    5.81678e-05, 0.0001176212, 0.0003362849, 0.0008453806, 0.001062347, 
    0.003996654, 0.0002207021, 4.0878e-05, -5.169256e-05,
  0.000308761, 7.645146e-05, 1.630554e-05, 4.533581e-07, 0.003090667, 
    0.0001702715, 0.04571756, 0.1142662, 0.005408008, 0.004848415, 
    0.01325936, 0.01113597, 0.1001329, 0.1500693, 0.08856291, 0.01213388, 
    0.003225602, 2.619394e-06, 2.010493e-07, 7.315579e-06, 7.612221e-06, 
    0.0007110329, 0.0004282093, 0.0243363, 0.001833003, 0.00154654, 
    0.002383027, 0.01004128, 0.0002343762,
  0.005952525, 0.1180791, 0.09271559, 0.00551509, 0.001761368, 0.02829862, 
    0.103112, 0.2557841, 0.1807731, 0.2642516, 0.1142592, 0.1545534, 
    0.1172404, 0.09330467, 0.07673496, 0.00484087, 0.005153762, 4.695738e-05, 
    -5.929506e-05, 0.002135264, 0.004676096, 0.04378198, 0.02520452, 
    0.1113452, 0.03522805, 0.002809485, 0.005717548, 0.03126466, 0.01241596,
  0.2229537, 0.2971037, 0.2333977, 0.1287909, 0.02641724, 0.02100794, 
    0.1274696, 0.3349482, 0.2296862, 0.1171009, 0.1300296, 0.1581434, 
    0.2221532, 0.1420914, 0.1517913, 0.1039037, 0.02854664, 0.05655767, 
    0.08594871, 0.09734833, 0.2655271, 0.2469387, 0.3198085, 0.1022223, 
    0.05256096, 0.1008316, 0.07424997, 0.2660766, 0.2746395,
  0.00103858, 0.003699443, 0.004016267, 0.02151454, 0.1065581, 0.2065932, 
    0.333758, 0.1311155, 0.3832444, 0.09593821, 0.2255881, 0.1550765, 
    0.2171017, 0.1144914, 0.1004562, 0.06741463, 0.01173364, 0.02904779, 
    0.005347024, 0.009611671, 0.02978512, 0.04196545, 0.03842662, 0.0774978, 
    0.1166831, 0.01407573, 0.005365838, 0.007508355, 0.0008960462,
  0.0103876, 0.004169641, -1.932283e-08, 0.0007588549, 0.003447375, 
    0.0006542745, 0.07076985, 0.1726765, 0.1626796, 0.08909109, 0.0629653, 
    0.1013766, 0.230103, 0.2223751, 0.1282312, 0.1037753, 0.09262808, 
    0.009849538, 0.01062309, 0.001198633, 0.07586509, 0.1118588, 0.1913946, 
    0.2133192, 0.09167442, 0.06709392, 0.00486558, 0.0006678636, 0.01824205,
  0.06697293, 0.03567025, 0.004260977, 3.176019e-05, -2.52074e-05, 
    0.003467313, 0.01195295, 0.06203523, 0.1526155, 0.1821437, 0.2375278, 
    0.1369194, 0.2102201, 0.2398376, 0.1890692, 0.2066565, 0.1186219, 
    0.1030268, 0.01122058, 0.005619929, 0.02890974, 0.06857138, 0.07953122, 
    0.1212324, 0.1517022, 0.153804, 0.1118973, 0.06753749, 0.02916195,
  0.0856192, 0.04459083, 0.03116861, 0.03159756, 0.07270099, 0.08637735, 
    0.04096374, 0.01976641, 0.02895964, 0.120185, 0.1622267, 0.2100803, 
    0.1911308, 0.162296, 0.1847337, 0.162214, 0.1220809, 0.1270634, 
    0.1035658, 0.02719637, 0.08514163, 0.1171609, 0.08967903, 0.1060584, 
    0.1150547, 0.1267927, 0.1316549, 0.1439213, 0.1135144,
  0.07666456, 0.03016395, 0.06254471, 0.03296335, 0.06333482, 0.08100145, 
    0.07446125, 0.1034424, 0.06012383, 0.09625567, 0.1359282, 0.1505407, 
    0.1659516, 0.1295472, 0.09549021, 0.06415861, 0.02281378, 0.02116976, 
    0.00762266, 0.01211524, 0.02166056, 0.0309366, 0.03876378, 0.02631113, 
    0.06735048, 0.06529417, 0.05902918, 0.05669133, 0.0750733,
  0.01036475, 0.01662184, 0.03153756, 0.04491792, 0.01858655, 0.009847477, 
    0.01461727, 0.0295656, 0.03127725, 0.03867475, 0.02472759, 0.02500723, 
    0.02061469, 0.05643638, 0.02864799, 0.01549941, 0.006630086, 0.001676282, 
    0.002576259, 0.002499804, 0.01296072, 0.002987806, 0.01093674, 
    0.009148734, 0.005455581, 0, 0.001069964, 0.0101828, 0.01683957,
  0.0001861413, -4.197693e-05, 0.0006524652, 0.0006411755, -0.0001124185, 
    0.001235296, 0.0003449296, 0.003074939, 0.0001355998, 0.003183647, 
    0.001326065, -3.27067e-05, 0.000971546, 0.003406686, 0.004142717, 
    0.0007451845, -5.104042e-05, -2.871994e-05, -1.297241e-10, -1.690306e-09, 
    0, 1.380069e-08, -1.955286e-06, 4.071027e-06, -1.031087e-07, 0, 0, 
    -1.5554e-07, -1.639038e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.0002285478, -6.120805e-06, -3.285853e-07, 0, 0, 0, 0, 0, -1.159831e-05, 
    -5.768487e-06, -1.094013e-05, 0, 0, -6.07032e-05, 0.002214708, 
    0.001070206, -2.868519e-05, -6.357508e-05, -3.133341e-06, 0, 0.001449556, 
    0.002385753, 0, 0.0001099218, 0.001295185, 7.936209e-05, -1.614889e-06, 
    0, 0,
  0.0001049715, 0.001363053, 0.0003272569, 0.0004001087, 8.638324e-05, 0, 0, 
    0.000351867, 0.0004689807, 0.0004142833, 0.001287591, 0.002016513, 
    0.001687406, 0.006143374, 0.002529508, 0.003807365, 0.0008117257, 
    -6.428854e-05, 0, 0.0003507821, -3.681242e-05, 0.001534275, 0.01576376, 
    0.01788431, 0.0004037815, 0.003006403, 0.004773414, 0.0018721, 
    -6.005727e-05,
  0.03625989, 0.03967562, 0.0106475, 0.02222198, 0.01101394, 0.01374431, 
    0.003551475, 0.004543195, 0.01349167, 0.02589185, 0.02498285, 
    0.007995318, 0.006072138, 0.003341862, 0.01513505, 0.003215858, 
    0.006642748, 0.008102817, 0.01908396, 0.02210881, 0.04144467, 0.04587098, 
    0.05319234, 0.04043528, 0.007920194, 0.009251272, 0.004478123, 
    0.01994989, 0.03542637,
  0.05448879, 0.02711241, 0.01502461, 0.04315523, 0.0399519, 0.02891337, 
    0.0221111, 0.02079949, 0.02503581, 0.01437904, 0.01586283, 0.01511148, 
    0.01042144, 0.01964886, 0.03362191, 0.04760066, 0.07634605, 0.09925677, 
    0.09490681, 0.1555844, 0.1534222, 0.1074195, 0.1165539, 0.02563665, 
    0.05499818, 0.06168829, 0.05935199, 0.06688821, 0.09322605,
  0.007120916, 0.002580176, 0.001981245, 0.00251919, 0.003853765, 
    0.006589561, 0.009183267, -3.185608e-05, 0.00324098, 0.001861893, 
    0.01106584, 0.00719304, 0.003549245, 0.009556369, 0.09580146, 0.1461002, 
    0.1493303, 0.1483868, 0.2023519, 0.168504, 0.09970001, 0.04309483, 
    0.01861107, 0.005981605, 0.008913524, 0.03401254, 0.03046462, 0.05559396, 
    0.02494151,
  7.741098e-07, 2.761209e-05, 4.55076e-07, 0.002749888, -4.079726e-06, 
    5.385635e-08, 1.84923e-05, 0.0001955316, 5.650737e-07, 2.090008e-07, 
    1.925648e-07, 4.881543e-07, 0.00077603, 0.05496822, 0.05789319, 
    0.08208358, 0.05013674, 0.02052286, 0.00916952, 0.00086933, 6.276302e-06, 
    2.726961e-06, 4.5445e-05, 0.0003425725, 0.0001307839, 0.0004887341, 
    1.729441e-05, -7.705617e-06, 5.06183e-07,
  2.133515e-05, 8.474385e-06, 1.796549e-06, 2.745895e-07, 0.001728551, 
    0.0002328581, 0.03177154, 0.116604, 0.005015721, 0.008421052, 0.01275826, 
    0.002415972, 0.09470785, 0.1348109, 0.08069026, 0.01264921, 0.002790651, 
    1.840017e-06, 6.730314e-09, 5.024704e-07, 1.40668e-06, 0.0003628693, 
    0.003447382, 0.01935891, 2.956556e-05, 8.767046e-05, 9.864081e-05, 
    0.004418756, 4.668507e-05,
  0.002024156, 0.08760472, 0.04957256, 0.001865292, 0.0002852152, 0.02113688, 
    0.04747588, 0.1458612, 0.1575332, 0.2228346, 0.08860811, 0.132779, 
    0.1066259, 0.09133044, 0.06440579, 0.005815709, 0.004648235, 
    -3.078951e-05, -4.019049e-05, 0.001107516, 0.003089662, 0.01955993, 
    0.002757736, 0.1023889, 0.02958917, 0.004376092, 0.01029811, 0.01776002, 
    0.004135683,
  0.1909557, 0.2849854, 0.2151408, 0.103075, 0.02722879, 0.01573463, 
    0.09242983, 0.1836716, 0.2087933, 0.0777366, 0.08862029, 0.139454, 
    0.1946816, 0.1280557, 0.1080593, 0.08640077, 0.03073569, 0.05089594, 
    0.0738726, 0.09460969, 0.2532741, 0.224316, 0.2778684, 0.08396447, 
    0.05210308, 0.08719875, 0.06992662, 0.2447391, 0.2456013,
  0.0006533433, 0.0007403849, 0.003160218, 0.02289998, 0.1056729, 0.1971011, 
    0.3438934, 0.1052248, 0.360752, 0.07772521, 0.201992, 0.1410913, 
    0.1831202, 0.1069147, 0.06635962, 0.05384582, 0.004949418, 0.01739053, 
    0.006226509, 0.009946846, 0.02130874, 0.03662699, 0.03146274, 0.06636529, 
    0.07729004, 0.01161483, 0.006442092, 0.006314425, 0.001210132,
  0.01307095, 0.007363985, -1.439031e-08, 1.561053e-05, 0.0001849702, 
    0.0001226123, 0.058348, 0.1566578, 0.1624388, 0.0784485, 0.0560178, 
    0.08652145, 0.2206489, 0.2226149, 0.1189391, 0.0958184, 0.07061887, 
    0.006416942, 0.001759191, 6.791378e-05, 0.07786514, 0.1204117, 0.1445804, 
    0.1979645, 0.08315235, 0.03967024, 0.01086523, 2.633834e-05, 0.01677262,
  0.0753559, 0.04421911, 0.009212331, 0.0005278366, 0.0005509997, 
    0.005245182, 0.01820859, 0.09523802, 0.192154, 0.175576, 0.1982939, 
    0.1142533, 0.1871233, 0.2338516, 0.1836306, 0.1846531, 0.1251252, 
    0.101554, 0.004318243, 0.005399307, 0.05873369, 0.04609483, 0.07005545, 
    0.110629, 0.1385547, 0.1408339, 0.09237347, 0.05097032, 0.03856079,
  0.1152238, 0.1185271, 0.0787372, 0.1250953, 0.09363346, 0.1443778, 
    0.1016826, 0.06479101, 0.1305997, 0.191384, 0.1331513, 0.1885228, 
    0.1838621, 0.1180958, 0.1747446, 0.1848725, 0.143075, 0.1475227, 
    0.1297633, 0.07038649, 0.1022039, 0.1199001, 0.106637, 0.1429667, 
    0.1221351, 0.1331211, 0.1216761, 0.1467609, 0.108436,
  0.1308015, 0.1242735, 0.1081919, 0.08055386, 0.1083413, 0.1129065, 
    0.1541767, 0.1735944, 0.1403326, 0.1639499, 0.1740338, 0.2197254, 
    0.202273, 0.1742916, 0.108011, 0.1087762, 0.08232699, 0.09719053, 
    0.06717963, 0.09412516, 0.1390593, 0.1259414, 0.1439291, 0.08867499, 
    0.1276719, 0.1007868, 0.08614047, 0.1194211, 0.1750893,
  0.0762031, 0.1072462, 0.1238843, 0.1296473, 0.08466246, 0.06061094, 
    0.0561898, 0.09928937, 0.08745261, 0.1704201, 0.07870072, 0.05012554, 
    0.1288377, 0.1474559, 0.1137094, 0.1013059, 0.08780503, 0.05117037, 
    0.0336126, 0.02028027, 0.03092126, 0.02434759, 0.02269186, 0.02582805, 
    0.04670079, -0.0001635033, 0.002228904, 0.1285444, 0.09334105,
  0.006787708, 0.01127738, 0.04345261, 0.02371707, 0.009494793, 0.02244716, 
    0.01307991, 0.01839576, 0.01128008, 0.0302668, 0.04049652, 0.05888886, 
    0.04373957, 0.04602392, 0.02873666, 0.03572636, 0.037486, 0.03240993, 
    0.03328191, 0.01698378, 0.004139097, 0.001289778, 5.977227e-05, 
    -0.0007927126, 0.0006097749, 0.0001460848, -0.0003960604, -0.001743327, 
    0.02230146,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.019074e-05, 
    0.0002157805, 0, 0, 0, 0, 9.465223e-05, 0, 0, 0, 0, 0,
  0.001391773, 0.003163652, 0.002764266, 0.0002871641, -6.086822e-05, 0, 0, 
    0, -9.44147e-05, -1.153697e-05, -2.188027e-05, 0, 0.0006789069, 
    -9.541758e-05, 0.007775541, 0.005268224, 0.0005969689, 0.0005801353, 
    7.95918e-06, -1.234822e-06, 0.007150885, 0.005441534, -6.869399e-06, 
    0.001755975, 0.00715898, 0.003945215, 0.001776502, 0, 0,
  0.01420161, 0.02244752, 0.02936163, 0.0202827, 0.0009541807, 9.366311e-05, 
    0, 0.001396017, 0.001259029, 0.003620931, 0.009910146, 0.007670728, 
    0.004609447, 0.01043031, 0.01082814, 0.01352128, 0.004481331, 
    0.003285936, 0.0004671353, 0.002888364, 0.002707162, 0.009950046, 
    0.02042724, 0.02927092, 0.0121171, 0.01133107, 0.009108135, 0.009110078, 
    0.007736614,
  0.1112254, 0.1238512, 0.09728488, 0.1162191, 0.06684452, 0.04192353, 
    0.01295296, 0.01705248, 0.02779175, 0.04940732, 0.04155328, 0.02696682, 
    0.02370614, 0.005242182, 0.02702985, 0.01472388, 0.03123764, 0.04888729, 
    0.05108619, 0.07103461, 0.1029665, 0.09872659, 0.1247407, 0.09437521, 
    0.06953122, 0.08386459, 0.0616721, 0.05253252, 0.09597003,
  0.1339291, 0.086707, 0.0776886, 0.07142139, 0.08062802, 0.08584613, 
    0.08644684, 0.05899203, 0.0546827, 0.05563354, 0.05161377, 0.04025655, 
    0.02300741, 0.02653094, 0.04622721, 0.07061807, 0.09741044, 0.145804, 
    0.1310233, 0.1799047, 0.1925458, 0.1504193, 0.1535896, 0.07510392, 
    0.1253388, 0.1267369, 0.1152161, 0.14682, 0.1732728,
  0.008698632, 0.005452965, 0.005035922, 0.007512629, 0.008257197, 
    0.01002352, 0.009983596, 0.00154954, 0.001266015, 0.001551954, 
    0.02562642, 0.0165925, 0.009426071, 0.022197, 0.102088, 0.1500168, 
    0.1529088, 0.1343871, 0.1891516, 0.1368392, 0.08195908, 0.02647088, 
    0.007846175, 0.003841578, 0.01258493, 0.04475637, 0.03109462, 0.06460315, 
    0.02515414,
  1.233767e-07, 5.091444e-06, 3.584476e-07, 0.003110807, 1.259985e-05, 
    -8.300191e-06, -2.320779e-05, 0.0001085981, 3.006756e-06, 1.679666e-08, 
    8.564626e-08, -2.333656e-05, 0.007577017, 0.07457309, 0.06996416, 
    0.07885482, 0.0396171, 0.01431014, 0.004176339, 0.0006550546, 
    3.005388e-07, 1.53106e-07, 4.612818e-06, 2.458743e-06, 0.0001099735, 
    0.0003777248, -3.524746e-06, 0.0001463397, 4.308598e-07,
  3.08349e-06, 3.247373e-06, 1.170697e-06, -1.266812e-06, 0.001614519, 
    0.0001253887, 0.02779738, 0.122943, 0.01276483, 0.01183849, 0.01337435, 
    0.001309897, 0.09734432, 0.1309542, 0.07123654, 0.01151876, 0.002523297, 
    3.606118e-05, 2.603758e-08, 2.310929e-07, 1.322965e-06, 4.359329e-06, 
    0.001701949, 0.01119274, -1.681332e-05, 1.424535e-05, -2.210835e-06, 
    6.899465e-05, 8.155705e-06,
  0.0002489032, 0.07234312, 0.02488465, 0.0004317813, 0.0001834436, 
    0.01342048, 0.02291157, 0.06900422, 0.1192069, 0.168608, 0.06445839, 
    0.1077729, 0.1030396, 0.08348448, 0.05846383, 0.0108502, 0.003748948, 
    1.736661e-06, -5.761374e-05, 0.001319698, 0.001259779, 0.004385597, 
    0.002957378, 0.08973282, 0.02107741, 0.005873539, 0.006012227, 
    0.01205803, 0.0002895647,
  0.1491074, 0.2462372, 0.170936, 0.1013169, 0.03172446, 0.00991049, 
    0.0823735, 0.07416549, 0.1934104, 0.0589812, 0.06188224, 0.1208629, 
    0.1665462, 0.1127423, 0.08255444, 0.07443766, 0.03962399, 0.04694996, 
    0.06676307, 0.08869159, 0.2478132, 0.1921785, 0.2076942, 0.05988835, 
    0.04376452, 0.07450585, 0.06331047, 0.2260685, 0.2036149,
  0.002258607, 0.0002078908, 0.0005127246, 0.02841959, 0.1075565, 0.1848349, 
    0.343183, 0.09260201, 0.3268236, 0.05734321, 0.1836835, 0.1307608, 
    0.1403153, 0.1031521, 0.04478082, 0.04280676, 0.001421676, 0.01461733, 
    0.00484279, 0.009277805, 0.01835726, 0.02977863, 0.02034208, 0.05883897, 
    0.0429504, 0.0132412, 0.001390147, 0.006069991, 0.001563135,
  0.01301447, 0.006885455, 9.705642e-09, 2.685846e-06, 6.457164e-05, 
    0.0002446481, 0.05120853, 0.1416803, 0.1474632, 0.06676009, 0.04921141, 
    0.0692105, 0.2025983, 0.2089866, 0.116112, 0.1024927, 0.05905494, 
    0.003463143, 0.002594314, 3.213548e-05, 0.09580058, 0.115235, 0.101664, 
    0.1778511, 0.07191014, 0.02759331, 0.01817449, 9.390095e-05, 0.01423244,
  0.05408422, 0.03954889, 0.004412887, 0.001061074, 0.004986661, 0.006638233, 
    0.05365038, 0.1087749, 0.1793394, 0.1639178, 0.1812763, 0.1136027, 
    0.1774277, 0.2410034, 0.192254, 0.1580466, 0.1157945, 0.09068237, 
    0.001443938, 0.002985182, 0.05346997, 0.04128276, 0.06552431, 0.1046657, 
    0.1280713, 0.123972, 0.08302358, 0.0387695, 0.03303373,
  0.08609195, 0.1154708, 0.06375518, 0.1140286, 0.08060965, 0.133733, 
    0.07758661, 0.1255333, 0.1745589, 0.1541921, 0.1002548, 0.1722929, 
    0.1781325, 0.09050182, 0.1541216, 0.1673674, 0.1506355, 0.1685267, 
    0.1267494, 0.07185046, 0.07951145, 0.1026357, 0.1011704, 0.1463789, 
    0.1262295, 0.1318661, 0.1159727, 0.1200574, 0.09726032,
  0.1380864, 0.1398785, 0.109857, 0.09685852, 0.119106, 0.102255, 0.21261, 
    0.1956179, 0.1371135, 0.1334945, 0.1712754, 0.2053551, 0.2094815, 
    0.1692399, 0.108487, 0.1892644, 0.1498618, 0.2031674, 0.20823, 0.1486183, 
    0.1981634, 0.1667404, 0.1809036, 0.1277974, 0.1644375, 0.1438556, 
    0.116528, 0.1543709, 0.1886816,
  0.1522417, 0.1755022, 0.2195723, 0.1839605, 0.1344326, 0.139844, 0.1084607, 
    0.1380306, 0.1616138, 0.1965683, 0.1198592, 0.1278082, 0.1662336, 
    0.1601259, 0.1467677, 0.1756018, 0.1721777, 0.09817063, 0.129432, 
    0.1465973, 0.1485858, 0.08734933, 0.08967796, 0.05298062, 0.1525303, 
    0.003769531, 0.005381351, 0.2290895, 0.198829,
  0.06869899, 0.08839623, 0.1277029, 0.08482739, 0.0850964, 0.102115, 
    0.1099116, 0.1191306, 0.1151001, 0.1369617, 0.1365919, 0.1470574, 
    0.1559774, 0.1119215, 0.09331416, 0.1409695, 0.152198, 0.1524675, 
    0.1411935, 0.134535, 0.06940174, 0.08360711, 0.02840933, 0.01118037, 
    0.0476916, 0.005711109, -0.001266825, 0.05788716, 0.08650716,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001011072, 
    0.0005428356, 0, 0, 0, 0.0003325453, 0.002968938, 1.450068e-07, 0, 0, 0, 0,
  0.006513281, 0.01715452, 0.0275941, 0.01027596, -0.0001530756, 0, 
    -3.050905e-08, -3.670021e-06, -0.0002052042, 0.0002116038, -8.704302e-05, 
    -5.739292e-05, 0.002239401, 0.005610805, 0.02551527, 0.0146511, 
    0.002740532, 0.003801679, 0.001465564, -6.765651e-05, 0.01179313, 
    0.01517779, 0.0005252739, 0.007472302, 0.0121707, 0.01230964, 
    0.006077332, -0.0002622955, -7.47674e-05,
  0.01878605, 0.04457873, 0.09305923, 0.09437594, 0.05373613, 0.01483524, 
    0.003475056, 0.003566251, 0.006180609, 0.008934665, 0.03033287, 
    0.03147665, 0.05066619, 0.0409692, 0.03783346, 0.03859807, 0.03639552, 
    0.02858697, 0.006109246, 0.01313722, 0.03392177, 0.04397368, 0.05535965, 
    0.0742522, 0.04767316, 0.04022985, 0.04747984, 0.0411929, 0.01565348,
  0.1625336, 0.2148064, 0.1949374, 0.2036614, 0.1888619, 0.1421444, 
    0.08923347, 0.09724298, 0.07892191, 0.1118887, 0.1326853, 0.1231739, 
    0.1185659, 0.0589832, 0.08690591, 0.0853234, 0.074854, 0.1096851, 
    0.09755342, 0.1231056, 0.1734125, 0.1402434, 0.186957, 0.1632616, 
    0.1291759, 0.1680131, 0.1748572, 0.1260794, 0.1600566,
  0.1387161, 0.09058111, 0.07511889, 0.06876037, 0.0688739, 0.1075905, 
    0.1060473, 0.1000458, 0.08511472, 0.07306328, 0.07188927, 0.09614897, 
    0.07440878, 0.09813542, 0.0767211, 0.1270569, 0.1550779, 0.1832024, 
    0.1424186, 0.1912668, 0.2050523, 0.1564841, 0.1667091, 0.1363963, 
    0.1367694, 0.1121955, 0.1217875, 0.1703119, 0.1663107,
  0.01184396, 0.008888192, 0.006318704, 0.00794735, 0.01167026, 0.01577969, 
    0.008963875, 0.01256872, 0.0004664002, 0.003313355, 0.02465069, 
    0.02237974, 0.01971293, 0.02352473, 0.09331173, 0.1601714, 0.1461368, 
    0.1100298, 0.1480422, 0.101227, 0.05620491, 0.01900115, 0.001435812, 
    0.005626688, 0.01422188, 0.0444727, 0.03426087, 0.06559903, 0.02748802,
  1.165931e-07, 1.355934e-06, 1.552293e-07, 0.005195928, 0.002188462, 
    -6.646943e-07, -4.322152e-06, 3.425879e-05, 2.398424e-06, 4.611553e-08, 
    5.27134e-09, -9.09042e-05, 0.02190067, 0.08139525, 0.07102864, 
    0.07070516, 0.02074277, 0.004988275, 0.0007788822, 0.0001491225, 
    -7.15708e-07, -1.74292e-06, 7.177254e-07, -1.181136e-06, 0.0002711423, 
    0.00183087, -5.065035e-05, 0.003541526, 3.116647e-07,
  3.397705e-07, 1.950117e-06, 1.082101e-06, 7.054817e-05, 0.001255548, 
    5.256362e-05, 0.0309313, 0.1101021, 0.01314548, 0.01773639, 0.01529981, 
    0.002435135, 0.0972411, 0.1189266, 0.05273733, 0.00863425, 0.002585659, 
    9.722818e-06, 9.708347e-09, 1.515394e-07, 4.973619e-07, 1.861902e-07, 
    2.804854e-05, 0.0004975505, -2.55244e-06, 3.036652e-06, 3.569563e-07, 
    1.011669e-06, 3.764849e-07,
  0.0003403335, 0.0556118, 0.01252304, 0.0009584302, 0.0003335056, 
    0.009794448, 0.01389291, 0.02938898, 0.06988835, 0.1358786, 0.04893488, 
    0.08732595, 0.09513728, 0.06412382, 0.05156769, 0.009016472, 0.002635445, 
    2.253227e-05, -3.040247e-05, 0.0006973904, -2.993117e-05, 0.0005216501, 
    0.00560614, 0.07175846, 0.02943574, 0.008967289, 0.00438163, 0.003263169, 
    5.716729e-05,
  0.1133265, 0.192824, 0.1328283, 0.1241376, 0.03562164, 0.006258575, 
    0.06742638, 0.03357883, 0.1570345, 0.04257086, 0.03589142, 0.08994497, 
    0.1458865, 0.09214013, 0.06041381, 0.06701683, 0.04975758, 0.04864864, 
    0.0727928, 0.09404522, 0.2428331, 0.1708798, 0.1625931, 0.04375184, 
    0.03583838, 0.07071625, 0.05963897, 0.1958811, 0.1817297,
  0.001149336, 0.0006062215, 8.640157e-05, 0.02654026, 0.1213833, 0.1583523, 
    0.3620934, 0.08542274, 0.2950658, 0.03795164, 0.1829842, 0.127187, 
    0.09227495, 0.09294851, 0.03302576, 0.03270252, 0.00174947, 0.01058621, 
    0.00424926, 0.00669778, 0.01900263, 0.02367508, 0.01376795, 0.05078012, 
    0.02629657, 0.008386085, 0.0008901962, 0.00369956, 0.0006524481,
  0.01474083, 0.009314847, -3.836016e-11, 2.810185e-07, 0.0001852369, 
    0.0005290458, 0.04170775, 0.1304001, 0.1466043, 0.06005882, 0.04964661, 
    0.06207011, 0.1830659, 0.1818131, 0.1143321, 0.1085362, 0.05684609, 
    0.002688003, 0.008032305, 0.001266638, 0.0898671, 0.09500553, 0.07032529, 
    0.1551095, 0.05707265, 0.01966767, 0.01299002, 7.431552e-06, 0.01057527,
  0.04017732, 0.03396665, 0.003172864, 0.001867031, 0.01656091, 0.008548014, 
    0.0801231, 0.1035185, 0.1536598, 0.1561137, 0.1728487, 0.1217098, 
    0.1578705, 0.2275773, 0.2079611, 0.1304991, 0.1010302, 0.08445561, 
    0.000777362, 0.001134817, 0.03816565, 0.03464866, 0.05430762, 0.08978701, 
    0.1155379, 0.1124664, 0.07015849, 0.02795643, 0.02170187,
  0.07611278, 0.09216011, 0.04613603, 0.1021397, 0.07527728, 0.1213115, 
    0.06636935, 0.1521495, 0.1572979, 0.1377049, 0.08139125, 0.159382, 
    0.1603959, 0.08376779, 0.1366575, 0.1511641, 0.1422179, 0.1603325, 
    0.1298184, 0.07077946, 0.06328769, 0.09413292, 0.09053013, 0.1372404, 
    0.1228273, 0.1239996, 0.113436, 0.1156134, 0.08853857,
  0.1342268, 0.1308935, 0.1010609, 0.08406854, 0.1113547, 0.0837194, 
    0.1889377, 0.176805, 0.115965, 0.1193432, 0.1468949, 0.1795402, 
    0.1977173, 0.1574738, 0.1061876, 0.1929738, 0.171881, 0.2392713, 
    0.2789443, 0.1456345, 0.176517, 0.1515875, 0.1588951, 0.1320692, 
    0.1547641, 0.1504968, 0.1194194, 0.16873, 0.170654,
  0.1606581, 0.1699104, 0.1988812, 0.1706675, 0.1430734, 0.1487886, 
    0.1313922, 0.1451313, 0.1442245, 0.1643104, 0.1349786, 0.1212333, 
    0.1511872, 0.1518141, 0.1610867, 0.199336, 0.1847662, 0.1019222, 
    0.1198583, 0.1338235, 0.1479265, 0.12234, 0.1684163, 0.1118052, 
    0.1702168, 0.06075122, 0.01983649, 0.2277663, 0.2091737,
  0.09940183, 0.1232871, 0.1902998, 0.100703, 0.0886631, 0.1238763, 
    0.1749216, 0.1692764, 0.16703, 0.1617081, 0.1760107, 0.1790114, 
    0.1938676, 0.1544324, 0.1212914, 0.158597, 0.1796377, 0.1739752, 
    0.1773455, 0.1819579, 0.1496521, 0.1507057, 0.1370595, 0.05458431, 
    0.1665114, 0.04087148, 0.06513686, 0.08286831, 0.09679571,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.397549e-05, -9.760766e-06, 
    0.0001334786, 0.0008675585, 0.00383622, -2.848466e-05, -2.005667e-05, 
    -4.098374e-05, 0.001452118, 0.01135597, 0.006615304, 0.001489494, 
    0.004636579, -3.545139e-05, 0,
  0.03810383, 0.05773051, 0.08797365, 0.05947094, -0.0003568209, 
    -2.602928e-05, 0.0005313995, -2.383554e-05, -0.0003204912, 0.0004433683, 
    -6.689439e-05, -4.444391e-05, 0.004159315, 0.06654893, 0.07248869, 
    0.04036655, 0.03113328, 0.03482249, 0.02778358, 0.01987718, 0.03824682, 
    0.0455897, 0.05139767, 0.04230855, 0.04403611, 0.0262185, 0.01617679, 
    0.01495962, 0.02932236,
  0.08460352, 0.07974837, 0.1680789, 0.2043311, 0.1544467, 0.07016041, 
    0.04179538, 0.0376281, 0.05751099, 0.07166679, 0.1367764, 0.1708649, 
    0.1968642, 0.1376109, 0.1677386, 0.1221849, 0.1126571, 0.1003442, 
    0.04148785, 0.09324367, 0.1030509, 0.09674671, 0.1070815, 0.1371098, 
    0.1015736, 0.09676758, 0.1002089, 0.08598494, 0.08026385,
  0.2163226, 0.2681051, 0.2104183, 0.2029777, 0.187309, 0.1816761, 0.1239455, 
    0.1400361, 0.1683304, 0.1893618, 0.180716, 0.1972517, 0.2427044, 
    0.1670972, 0.1327114, 0.1245192, 0.1429388, 0.1429776, 0.1380284, 
    0.1652919, 0.2160823, 0.1939728, 0.2091906, 0.1978817, 0.154111, 
    0.1997995, 0.2154132, 0.1663605, 0.2144326,
  0.134618, 0.07455895, 0.05744048, 0.06051871, 0.06272345, 0.1082471, 
    0.09687835, 0.1042448, 0.09342545, 0.07479235, 0.07105336, 0.1069539, 
    0.08074769, 0.1295356, 0.1124921, 0.1397575, 0.1545906, 0.1889162, 
    0.1583763, 0.2025073, 0.2216446, 0.1626509, 0.1777464, 0.1658917, 
    0.1136856, 0.09675671, 0.1156492, 0.1505991, 0.1583987,
  0.01134823, 0.01325538, 0.006885564, 0.01202977, 0.01781419, 0.02461501, 
    0.008187292, 0.01244477, 0.0003196212, 0.00286163, 0.01824417, 
    0.01851201, 0.02196138, 0.02111578, 0.08313508, 0.1454237, 0.145444, 
    0.1066236, 0.1350715, 0.08685735, 0.04192747, 0.01051403, 0.003706674, 
    0.004374838, 0.0138867, 0.04383272, 0.03513439, 0.06109999, 0.02677833,
  6.848369e-08, 8.875615e-08, 4.797979e-08, 0.005918922, 0.005845471, 
    -1.105374e-06, -4.187083e-05, -0.0001344219, 3.285087e-06, 3.864773e-08, 
    3.956004e-10, -8.762838e-05, 0.0159334, 0.08592984, 0.06840864, 
    0.05735619, 0.0105141, 0.00388474, 0.0002709987, 5.661001e-07, 
    -3.121797e-07, -1.609616e-05, 3.658501e-07, 3.366258e-06, 0.001265004, 
    0.006027947, -9.687711e-05, 0.01166889, -8.758107e-07,
  7.919238e-08, 2.282292e-06, 1.924235e-06, 9.853919e-05, 0.001586745, 
    0.000155589, 0.02456263, 0.1045916, 0.01173986, 0.01682732, 0.01454657, 
    0.01954076, 0.09658065, 0.1215956, 0.0470891, 0.009374234, 0.006103034, 
    1.735148e-06, 1.204839e-09, 3.475387e-08, 8.784227e-08, 1.890349e-07, 
    1.552507e-06, 0.0002306286, -5.364891e-07, 7.46751e-07, 4.504993e-06, 
    9.711775e-07, 7.936541e-08,
  3.12323e-05, 0.03911825, 0.01353366, 0.001875573, 0.0006692763, 
    0.007854959, 0.01016443, 0.01554811, 0.05130034, 0.1286512, 0.04079225, 
    0.06667551, 0.09400177, 0.05731311, 0.0476848, 0.01261198, 0.001947619, 
    0.001160811, 0.001954906, 0.0002590465, -6.956529e-06, 9.219611e-05, 
    0.00672065, 0.05735401, 0.0422699, 0.0160153, 0.005808704, 0.001636207, 
    3.890364e-06,
  0.08764364, 0.1462291, 0.1125382, 0.139374, 0.03770574, 0.008510974, 
    0.0461095, 0.01688332, 0.1384724, 0.03337037, 0.02409424, 0.07466102, 
    0.1302543, 0.0904758, 0.05214705, 0.07124659, 0.06055243, 0.06342362, 
    0.07619609, 0.09589157, 0.236863, 0.1611243, 0.1347556, 0.03585712, 
    0.03488579, 0.06685811, 0.05811071, 0.177626, 0.1598907,
  0.003739719, 0.0001646999, 0.0001787591, 0.0270792, 0.122798, 0.1514347, 
    0.3549219, 0.08592768, 0.2840112, 0.0326945, 0.1886585, 0.1232298, 
    0.07066624, 0.08380071, 0.0201767, 0.02346789, 0.0001799658, 0.004594065, 
    0.001647959, 0.002709112, 0.02602049, 0.02013224, 0.01010745, 0.0475275, 
    0.01932239, 0.004309964, 0.005404803, 0.002111026, 0.003344546,
  0.03522673, 0.01167532, -2.946093e-11, 2.272862e-08, 0.0006093853, 
    0.001399328, 0.03421151, 0.1283917, 0.1443266, 0.0515634, 0.04942904, 
    0.05639829, 0.1656398, 0.1642604, 0.1054909, 0.08789573, 0.03465713, 
    0.001874033, 0.01327426, 0.001499898, 0.07521397, 0.06653121, 0.05169399, 
    0.130229, 0.04004297, 0.01077379, 0.01329694, -1.60165e-05, 0.01809802,
  0.03686091, 0.03689896, 0.00254678, 0.001880976, 0.02468909, 0.0115561, 
    0.08267074, 0.09594373, 0.1250381, 0.1361703, 0.1416023, 0.1151846, 
    0.1610754, 0.2058966, 0.1850488, 0.1105123, 0.1126007, 0.07170574, 
    0.00102655, 0.000202546, 0.03950686, 0.02697972, 0.04387949, 0.08222662, 
    0.1087857, 0.09000516, 0.05258444, 0.02041386, 0.01293821,
  0.06970421, 0.08662176, 0.0354039, 0.09185664, 0.07055568, 0.1048475, 
    0.06268947, 0.1577159, 0.1440695, 0.132509, 0.06992449, 0.1455017, 
    0.1565406, 0.08106403, 0.128521, 0.1402263, 0.1370793, 0.1501437, 
    0.1246736, 0.07095069, 0.05141843, 0.08424671, 0.0836622, 0.1293554, 
    0.1179333, 0.1183703, 0.1019977, 0.1231935, 0.07674795,
  0.1313552, 0.1262619, 0.09667134, 0.07697111, 0.09006853, 0.06603336, 
    0.1634168, 0.1606824, 0.1011317, 0.109054, 0.1249862, 0.1545442, 
    0.1850482, 0.1481751, 0.1128249, 0.204659, 0.1588318, 0.2462717, 0.27173, 
    0.125025, 0.1444904, 0.1202509, 0.1353089, 0.1426971, 0.1413463, 
    0.1446331, 0.1107599, 0.164158, 0.1551898,
  0.162119, 0.1638927, 0.1855555, 0.166913, 0.1312281, 0.1368574, 0.1383682, 
    0.1288826, 0.1133013, 0.1315663, 0.109042, 0.1115885, 0.1394745, 
    0.1350602, 0.1625191, 0.1889584, 0.1623287, 0.08922058, 0.1111456, 
    0.1233183, 0.1417045, 0.1298929, 0.1989384, 0.1580802, 0.1787048, 
    0.1871178, 0.108505, 0.2177349, 0.199257,
  0.0995303, 0.1291628, 0.1973924, 0.1100224, 0.08518183, 0.1316046, 
    0.175183, 0.1706661, 0.1550161, 0.1494979, 0.16603, 0.1848268, 0.1914083, 
    0.1531059, 0.1212922, 0.1577416, 0.1871902, 0.1539652, 0.1719587, 
    0.177806, 0.1522263, 0.153836, 0.1772776, 0.0886642, 0.211689, 0.1293435, 
    0.1377559, 0.08352627, 0.08807614,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.103322e-06, 0.002983405, 
    0.0142994, 0.01325393, 0.0105505, 0.008641879, -8.94387e-05, 
    -0.0002178518, 0.0007328084, 0.005510862, 0.03882567, 0.03857921, 
    0.02205606, 0.02665698, 0.0003090955, 0,
  0.08765777, 0.1421727, 0.1470089, 0.1174266, -0.001047291, -0.001113185, 
    0.01507308, -7.963431e-05, -0.0003193613, -0.0001321175, 0.0008126751, 
    0.0009550001, 0.03549021, 0.1839575, 0.1796139, 0.1270427, 0.1143209, 
    0.1114469, 0.09233734, 0.108672, 0.1293754, 0.1361202, 0.1277663, 
    0.1063562, 0.08361714, 0.03953933, 0.03236669, 0.03916972, 0.06847718,
  0.1416255, 0.1379777, 0.238464, 0.2313067, 0.1837639, 0.1176209, 
    0.09401216, 0.07777964, 0.08711959, 0.1315985, 0.1994272, 0.237936, 
    0.2579853, 0.2021425, 0.2246449, 0.1540604, 0.1878533, 0.1575559, 
    0.1139201, 0.1583467, 0.1907406, 0.1959376, 0.162776, 0.215648, 
    0.1809398, 0.1797709, 0.1796924, 0.1252188, 0.1511435,
  0.2417729, 0.2833835, 0.1994517, 0.1966328, 0.1904432, 0.1900322, 
    0.1400012, 0.1538678, 0.1983727, 0.213393, 0.2075405, 0.2287179, 
    0.2443722, 0.1486551, 0.1384177, 0.1654338, 0.1561397, 0.175982, 
    0.1617215, 0.182193, 0.2223778, 0.1923198, 0.2360191, 0.1990841, 
    0.1551975, 0.2041607, 0.2322379, 0.1837862, 0.2283788,
  0.1203434, 0.06740886, 0.04881593, 0.05960213, 0.06529465, 0.1075105, 
    0.09737962, 0.105753, 0.09078106, 0.07892568, 0.07744032, 0.1033599, 
    0.07199182, 0.1155405, 0.1087255, 0.1380514, 0.1477474, 0.1853583, 
    0.1666128, 0.1975834, 0.2193217, 0.1660394, 0.1877342, 0.1657119, 
    0.08520027, 0.08446986, 0.1035306, 0.1371283, 0.1447954,
  0.009814717, 0.02000131, 0.007737223, 0.01939131, 0.02629838, 0.03030188, 
    0.008698197, 0.00904142, -7.94282e-07, 0.001067527, 0.01309998, 
    0.007442999, 0.02000385, 0.02036571, 0.06762503, 0.1364913, 0.1380789, 
    0.09484373, 0.1322241, 0.08339955, 0.0467904, 0.007530613, 0.002272706, 
    0.0005806171, 0.01411114, 0.04275013, 0.03023162, 0.05498107, 0.02748518,
  5.635467e-09, -3.325238e-09, -3.374603e-08, 0.007750284, 0.007164254, 
    -5.299712e-07, 0.0003179551, 0.0003004283, -8.711768e-06, 2.680614e-08, 
    1.967035e-09, 0.002270567, 0.01383837, 0.08361031, 0.06585474, 
    0.05340442, 0.005582686, 0.004154888, 5.99474e-05, 3.132627e-07, 
    -6.873282e-08, -0.0001293095, 1.026286e-07, 1.433975e-05, 0.0008615184, 
    0.002899173, -8.574274e-05, 0.01329421, -3.222389e-05,
  5.421798e-09, 3.46565e-06, 4.150437e-06, 6.599528e-05, 0.00209965, 
    0.0006138312, 0.01693697, 0.09983052, 0.01587412, 0.008303882, 
    0.02006228, 0.03023652, 0.1077566, 0.1165715, 0.05326, 0.01228548, 
    0.009087538, 4.047665e-06, 4.120505e-07, 2.581317e-09, 5.400287e-08, 
    1.40361e-07, 7.379824e-07, 0.0002273357, -2.323578e-07, 2.857348e-07, 
    5.131379e-05, 1.013889e-06, 4.316779e-08,
  0.0001137179, 0.03232202, 0.02180147, 0.003049949, 0.0009724137, 
    0.007466129, 0.009483078, 0.01267007, 0.03936275, 0.1314448, 0.03648124, 
    0.05389371, 0.08735839, 0.05718518, 0.05376628, 0.01265134, 0.002439464, 
    0.002563406, 0.002956558, 0.0001152823, -6.534076e-05, 0.0002544913, 
    0.01235827, 0.04728849, 0.05323215, 0.02673457, 0.01124955, 0.003415498, 
    1.466779e-06,
  0.08001328, 0.1297265, 0.1100165, 0.1744668, 0.04923918, 0.01503695, 
    0.0394123, 0.01198289, 0.1235628, 0.0356989, 0.01879594, 0.06986357, 
    0.118252, 0.08186352, 0.05483827, 0.07771749, 0.0674473, 0.07489127, 
    0.07849767, 0.1070209, 0.2315357, 0.1506394, 0.1156866, 0.03100513, 
    0.03805876, 0.06769572, 0.06520365, 0.1760288, 0.1461724,
  0.02593854, 0.0002631441, 0.001041969, 0.0274202, 0.1281057, 0.1234171, 
    0.342358, 0.09827437, 0.2745677, 0.02707751, 0.1834921, 0.1282137, 
    0.06332445, 0.07389975, 0.01219728, 0.01269224, 0.0003164482, 
    0.008112929, 0.0001956919, 0.006482346, 0.02424019, 0.01923632, 
    0.007848128, 0.04336398, 0.01409362, 0.008503343, 0.01259182, 
    0.003166003, 0.02490718,
  0.07790583, 0.02329718, 0, 1.121932e-08, 0.00271541, 0.0009426934, 
    0.02734886, 0.1346678, 0.1559935, 0.04778052, 0.04515224, 0.04882387, 
    0.157247, 0.1534272, 0.09430788, 0.06133119, 0.01870316, 0.002127199, 
    0.01685391, 0.002377601, 0.07294928, 0.03948132, 0.04270916, 0.1024193, 
    0.029957, 0.009214628, 0.01152765, -8.209869e-06, 0.0295504,
  0.03522925, 0.03867953, 0.003205227, 0.001973958, 0.02486315, 0.009317487, 
    0.07625113, 0.08637077, 0.1095629, 0.1193121, 0.112074, 0.1053964, 
    0.1534906, 0.2128752, 0.1731326, 0.08006757, 0.07734209, 0.07634486, 
    0.00087008, 0.0002740089, 0.05006099, 0.02316113, 0.03904075, 0.07863102, 
    0.08919403, 0.06944406, 0.03982756, 0.01427131, 0.006386369,
  0.05826334, 0.09138659, 0.02862727, 0.08441443, 0.06475231, 0.09517168, 
    0.05627381, 0.1489804, 0.1357842, 0.1265748, 0.06461693, 0.1363725, 
    0.1390386, 0.07989889, 0.1242496, 0.1367694, 0.1182723, 0.1500775, 
    0.1357445, 0.06496751, 0.04793711, 0.0739429, 0.07815594, 0.1237706, 
    0.104198, 0.1136016, 0.1084824, 0.1186694, 0.07742453,
  0.1140429, 0.1190495, 0.09448034, 0.05971423, 0.07590321, 0.06347843, 
    0.1469503, 0.1550896, 0.09066803, 0.1022393, 0.1046883, 0.1496821, 
    0.1713057, 0.1505005, 0.1227449, 0.1944765, 0.1470544, 0.2443864, 
    0.2646902, 0.1148155, 0.1171483, 0.1028924, 0.1222451, 0.152034, 
    0.1322118, 0.1335754, 0.1067147, 0.1412734, 0.1399397,
  0.160547, 0.1677308, 0.1792074, 0.1682116, 0.1304115, 0.128991, 0.1364993, 
    0.1142531, 0.1044998, 0.1206215, 0.09039803, 0.1041902, 0.126122, 
    0.1249633, 0.1812811, 0.1763511, 0.1410575, 0.07317665, 0.1066655, 
    0.1139686, 0.1470365, 0.1328479, 0.2011062, 0.1678041, 0.1787308, 
    0.2642718, 0.2057217, 0.2011851, 0.1983401,
  0.09641407, 0.1351274, 0.2002057, 0.1163636, 0.08124293, 0.1211835, 
    0.1717721, 0.1724995, 0.1375356, 0.138544, 0.1579268, 0.1797105, 
    0.1849623, 0.1634006, 0.1271741, 0.1567363, 0.1804129, 0.1510102, 
    0.1772819, 0.1797982, 0.1534733, 0.1524899, 0.179337, 0.09351161, 
    0.2342272, 0.1815857, 0.1678036, 0.07969432, 0.08629508,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008529252, 0.06235649, 0.09070362, 
    0.09039178, 0.05788322, 0.02030272, 0.0003088322, 0.0001981691, 
    0.00232929, 0.0171681, 0.09128527, 0.08112973, 0.05764983, 0.0725171, 
    0.0123057, 0,
  0.1605815, 0.1965752, 0.2455651, 0.1891039, 0.01277403, 0.004623711, 
    0.02612289, 1.648713e-05, 0.0002329406, 0.002135935, 0.002926398, 
    0.006128022, 0.1257137, 0.2044004, 0.2305107, 0.167007, 0.157128, 
    0.1633399, 0.151611, 0.1869859, 0.232613, 0.2294222, 0.2236553, 
    0.2105159, 0.1632417, 0.08531302, 0.09309915, 0.09980202, 0.1275719,
  0.1765552, 0.1953733, 0.2866379, 0.2563235, 0.2080384, 0.1623975, 
    0.1246515, 0.130672, 0.1373328, 0.1840612, 0.276513, 0.2831365, 
    0.2934132, 0.219308, 0.2380145, 0.1637292, 0.2103679, 0.1673972, 
    0.1401455, 0.162369, 0.2198448, 0.2369523, 0.1999885, 0.2528225, 
    0.2272503, 0.2343195, 0.2391651, 0.187231, 0.1992113,
  0.2565455, 0.2794074, 0.198466, 0.194687, 0.1773669, 0.1895767, 0.1490481, 
    0.1566696, 0.2295946, 0.2382234, 0.2239544, 0.2375108, 0.2372963, 
    0.1412737, 0.1281169, 0.1690137, 0.1604992, 0.1780727, 0.1605456, 
    0.1929744, 0.2247305, 0.1998859, 0.213711, 0.2082798, 0.1458033, 
    0.1923227, 0.2270132, 0.2119115, 0.2343338,
  0.1301758, 0.06495633, 0.05177683, 0.05595439, 0.0693898, 0.1064577, 
    0.09814848, 0.109323, 0.09244122, 0.07043654, 0.08297899, 0.1075007, 
    0.06211479, 0.1004192, 0.1026864, 0.13126, 0.1404618, 0.1722372, 
    0.173645, 0.1852889, 0.2129709, 0.1642794, 0.1656009, 0.1613045, 
    0.06202871, 0.08087421, 0.09502763, 0.1409678, 0.1296774,
  0.008403518, 0.02762254, 0.01396438, 0.02734203, 0.02866278, 0.03338811, 
    0.01064594, 0.008064792, -2.154568e-05, 0.0003781789, 0.01044227, 
    0.004717728, 0.02205352, 0.01757356, 0.06131327, 0.1297704, 0.1191183, 
    0.08072625, 0.1293703, 0.05986033, 0.03747804, 0.009416194, 0.002485581, 
    0.001393247, 0.01530108, 0.05206181, 0.02921694, 0.05436573, 0.02919784,
  -3.883876e-08, -8.306188e-10, -4.735416e-05, 0.01042938, 0.01536484, 
    1.023899e-05, 0.002794925, 1.378437e-05, -9.302026e-05, 1.169671e-08, 
    7.294726e-09, 0.0001488886, 0.01680012, 0.07928629, 0.05904046, 
    0.03838304, 0.006006802, 0.007978697, 0.0008416864, -1.596878e-07, 
    -4.606579e-07, 0.0008045519, 4.284307e-08, 3.252022e-07, 0.0002930135, 
    5.063086e-05, 0.0001874086, 0.01375977, 0.001697838,
  4.038051e-08, 1.54397e-06, 3.324269e-06, 4.786467e-05, 0.00410187, 
    0.004357006, 0.01049537, 0.08287464, 0.01992748, 0.007467899, 0.01899536, 
    0.03664011, 0.1074034, 0.1101172, 0.05006593, 0.01627433, 0.007560277, 
    1.122145e-05, 4.974178e-06, 2.757676e-09, -1.340354e-11, 2.451383e-08, 
    3.61003e-07, 0.0003500572, -6.007784e-05, 9.617394e-07, 0.0001097887, 
    4.298078e-05, 1.672418e-08,
  0.0006381818, 0.02893156, 0.03115093, 0.002126324, 0.001544496, 
    0.008467222, 0.008355048, 0.009377007, 0.04306426, 0.1323413, 0.02748563, 
    0.04563517, 0.07841015, 0.0558982, 0.05256005, 0.01480503, 0.004300579, 
    0.006534307, 0.009881543, 0.001925542, -8.928958e-05, 0.0001259463, 
    0.01018774, 0.04877497, 0.06524111, 0.04916406, 0.01546419, 0.00603504, 
    -3.156379e-08,
  0.0730973, 0.1247249, 0.1073472, 0.2062287, 0.08616545, 0.01699063, 
    0.03420294, 0.0107329, 0.09382982, 0.04793585, 0.01826095, 0.06462908, 
    0.1202761, 0.0769949, 0.05282379, 0.07938338, 0.06952876, 0.09034595, 
    0.08102266, 0.1336499, 0.2383468, 0.132475, 0.1014748, 0.0318995, 
    0.03484467, 0.06266222, 0.07698481, 0.1816955, 0.1479607,
  0.04081598, 0.001990451, 0.000164449, 0.01084126, 0.100567, 0.09067037, 
    0.3572212, 0.1104701, 0.3007148, 0.023973, 0.1940107, 0.1311792, 
    0.06344845, 0.06111901, 0.01076946, 0.005579562, 9.113397e-05, 
    0.0007994988, 0.0001887406, 0.007275668, 0.02506413, 0.01845612, 
    0.006187546, 0.04803874, 0.01219879, 0.01312233, 0.0111635, 0.0107745, 
    0.02596287,
  0.05936515, 0.01752597, -5.476043e-11, 8.522089e-09, 0.0004457418, 
    0.0002525954, 0.03173804, 0.1450908, 0.1709853, 0.05371196, 0.04816563, 
    0.04708879, 0.1511622, 0.1441436, 0.08069754, 0.04322292, 0.009438039, 
    9.229407e-05, 0.01048073, 0.006533456, 0.06226332, 0.02790664, 
    0.04189223, 0.08527155, 0.02480441, 0.00787201, 0.008659098, 
    -2.208723e-06, 0.02386378,
  0.0336073, 0.03455967, 0.00248029, 0.002152759, 0.03043716, 0.009671137, 
    0.08132292, 0.06804274, 0.09276249, 0.1178714, 0.09354855, 0.09160008, 
    0.1496929, 0.2109314, 0.1457801, 0.07140651, 0.06661159, 0.06503382, 
    0.0005709328, 0.000148698, 0.08744063, 0.02475813, 0.04704247, 0.0799098, 
    0.08571489, 0.0650098, 0.04060586, 0.008930778, 0.002695287,
  0.04388157, 0.08777367, 0.02488549, 0.08135688, 0.06161904, 0.09076138, 
    0.05819868, 0.1335381, 0.1274632, 0.1255899, 0.06907724, 0.1206362, 
    0.1306363, 0.07602222, 0.1035867, 0.1325225, 0.1203428, 0.1470528, 
    0.1297487, 0.06154682, 0.04697535, 0.07146741, 0.07393462, 0.1056291, 
    0.09701311, 0.1132259, 0.1117328, 0.1264467, 0.09703761,
  0.1222384, 0.1177391, 0.09889133, 0.05254703, 0.06007931, 0.06048179, 
    0.1492257, 0.1522017, 0.09017137, 0.1035157, 0.08420844, 0.1375911, 
    0.1722792, 0.143673, 0.1180736, 0.1858046, 0.1512167, 0.24863, 0.2588844, 
    0.1131731, 0.1036864, 0.1016763, 0.1134802, 0.1528826, 0.1385664, 
    0.138137, 0.1320516, 0.166249, 0.1445069,
  0.1865558, 0.2238261, 0.1857174, 0.1668443, 0.126539, 0.1234255, 0.1284166, 
    0.1013922, 0.1021067, 0.1088883, 0.07817993, 0.1099572, 0.1186104, 
    0.1284907, 0.1746904, 0.1785632, 0.1279004, 0.06634037, 0.09213157, 
    0.09557225, 0.1575928, 0.1447032, 0.2069925, 0.1874308, 0.1935407, 
    0.2508121, 0.2189052, 0.1858294, 0.1990486,
  0.118573, 0.1580715, 0.2048942, 0.1250582, 0.08194785, 0.1122883, 
    0.1736532, 0.1709543, 0.1496985, 0.1453907, 0.1634157, 0.172125, 
    0.1935248, 0.1832755, 0.1302547, 0.1669258, 0.2003526, 0.1617721, 
    0.1827797, 0.1761394, 0.1514259, 0.1499473, 0.1916274, 0.1038737, 
    0.228054, 0.1956132, 0.1743688, 0.08974218, 0.1059471,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -2.40997e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.756987e-06, 0.06948008, 
    0.1138662, 0.1205333, 0.1179888, 0.09375037, 0.07362962, 0.0177471, 
    0.0114005, 0.005705718, 0.04107539, 0.1979206, 0.1496234, 0.1089909, 
    0.1396547, 0.05074295, 0.002552773,
  0.23333, 0.2964259, 0.3054, 0.2444976, 0.0555599, 0.02065505, 0.05669111, 
    0.006796938, 0.008280012, 0.02655772, 0.01765519, 0.03114986, 0.2079841, 
    0.2571468, 0.2716187, 0.1931723, 0.1607653, 0.1914467, 0.1721778, 
    0.2082995, 0.2392062, 0.2449895, 0.2485127, 0.2815735, 0.213992, 
    0.1489382, 0.1544851, 0.1458128, 0.2060096,
  0.1901849, 0.2148468, 0.3014463, 0.2749564, 0.2251368, 0.1819853, 
    0.1428743, 0.1741442, 0.1500285, 0.2041193, 0.2997844, 0.3029826, 
    0.2841683, 0.2387513, 0.2307111, 0.1679194, 0.2144226, 0.1595783, 
    0.1406845, 0.1661124, 0.2294405, 0.2472582, 0.221801, 0.2564074, 
    0.2172899, 0.2483499, 0.236217, 0.1974809, 0.1949051,
  0.2660362, 0.2712141, 0.1833454, 0.1921259, 0.1681855, 0.1872558, 
    0.1541546, 0.1631538, 0.2464251, 0.2589257, 0.2269678, 0.2225597, 
    0.2198699, 0.1346166, 0.1276954, 0.143632, 0.1467039, 0.1719054, 
    0.1638224, 0.1911672, 0.218406, 0.1953906, 0.2043502, 0.195024, 
    0.1389872, 0.1845332, 0.2414686, 0.2173867, 0.224908,
  0.1259812, 0.06292489, 0.05588727, 0.05506343, 0.0701485, 0.09643786, 
    0.09776723, 0.1206305, 0.09021878, 0.06791643, 0.08573245, 0.1022362, 
    0.06773561, 0.09651382, 0.1012366, 0.1299678, 0.1332078, 0.1576188, 
    0.1709599, 0.1780438, 0.194016, 0.1557809, 0.1674898, 0.1685809, 
    0.0500413, 0.07460333, 0.0953092, 0.1356365, 0.121349,
  0.01218079, 0.02685959, 0.0228107, 0.02790738, 0.03317507, 0.03007527, 
    0.01360684, 0.007093734, -3.574249e-05, 0.001343324, 0.004089763, 
    0.004615966, 0.02398365, 0.0149321, 0.05971713, 0.1026295, 0.1162348, 
    0.06975035, 0.13628, 0.06004707, 0.03350735, 0.01094689, 0.005384927, 
    0.002083398, 0.01927048, 0.05589076, 0.03206331, 0.05398563, 0.0309289,
  -5.301808e-06, 1.942084e-10, -6.37779e-05, 0.01512782, 0.01833857, 
    0.0001905874, 0.005030086, 0.001009375, -0.0002825939, 6.137433e-09, 
    3.036433e-08, 0.0009883065, 0.01997583, 0.07884488, 0.06471801, 
    0.02497299, 0.006878606, 0.01300544, 8.038773e-05, -1.518643e-06, 
    -2.571421e-06, 0.001976402, 3.674032e-08, 1.580372e-06, 0.0004288117, 
    0.0003307561, 0.0007982756, 0.01368781, 0.003667884,
  6.465918e-08, 1.123588e-06, 4.039795e-06, 5.723107e-05, 0.00595811, 
    0.009258982, 0.01380227, 0.0836353, 0.02736457, 0.008454321, 0.02917753, 
    0.02534552, 0.1091854, 0.109748, 0.05452634, 0.02168687, 0.01123869, 
    0.0003864477, 3.224178e-05, 2.52164e-08, 1.021378e-08, 7.868016e-08, 
    4.166768e-06, 0.001165355, 2.238707e-05, 3.536044e-07, 4.307165e-06, 
    1.770204e-05, 3.4185e-08,
  0.004541385, 0.03334805, 0.04587772, 0.01317254, 0.0009591164, 0.007967085, 
    0.008072313, 0.01003943, 0.0529158, 0.1344591, 0.02702929, 0.05350847, 
    0.08438893, 0.06039112, 0.05516683, 0.0164493, 0.00938811, 0.006498451, 
    0.0125529, 0.008063227, 0.0009618888, 0.0003640597, 0.009876097, 
    0.0477258, 0.07797316, 0.07108453, 0.02563488, 0.01499765, 0.003733461,
  0.06727467, 0.1141863, 0.1067248, 0.273192, 0.1047338, 0.02293442, 
    0.04292055, 0.01187303, 0.07687478, 0.06873921, 0.0278291, 0.07088409, 
    0.1248431, 0.09056055, 0.05409563, 0.09390721, 0.07414369, 0.1065917, 
    0.09035499, 0.1437631, 0.2642611, 0.1209776, 0.1097176, 0.03655181, 
    0.0362211, 0.05954925, 0.09134714, 0.1760231, 0.1550942,
  0.01247625, 0.000382884, -8.627339e-07, 0.0004801374, 0.07156949, 
    0.09387361, 0.4055862, 0.1412379, 0.3553322, 0.0322686, 0.2192836, 
    0.1413219, 0.0761776, 0.05435847, 0.01018756, 0.003326401, 0.0001776499, 
    0.0002700821, 0.009529253, 0.01378908, 0.03265736, 0.02070845, 
    0.005548627, 0.04997194, 0.01016293, 0.007178899, 0.00794854, 
    0.007313147, 0.01942103,
  0.01807385, 0.006639976, 6.353039e-08, 1.830189e-08, 0.0003369103, 
    7.738867e-05, 0.0460569, 0.1484641, 0.1849372, 0.0622341, 0.04990781, 
    0.05827723, 0.1649566, 0.1413385, 0.07186934, 0.04013902, 0.01371123, 
    0.0004888472, 0.007629007, 0.00318398, 0.05735523, 0.02751032, 
    0.05043422, 0.07680923, 0.02037355, 0.005962528, 0.005965339, 
    6.817232e-08, 0.01156304,
  0.03361938, 0.03283032, 0.003958431, 0.003046704, 0.02812652, 0.007027153, 
    0.09651844, 0.04211305, 0.07406107, 0.1245685, 0.08794537, 0.09134589, 
    0.1521965, 0.2350897, 0.134585, 0.06224634, 0.0504775, 0.05678675, 
    0.0008641644, 0.0004241197, 0.1081593, 0.03740808, 0.04784657, 
    0.08724353, 0.08758666, 0.05765109, 0.04392288, 0.008203825, 0.002114447,
  0.04526775, 0.07738274, 0.02602578, 0.07487006, 0.05949638, 0.09172992, 
    0.06652562, 0.134302, 0.1245051, 0.1278707, 0.07044377, 0.1108768, 
    0.1215461, 0.07400102, 0.1004117, 0.1307584, 0.119055, 0.1454728, 
    0.1298633, 0.05552348, 0.04589027, 0.06554497, 0.07325574, 0.1027611, 
    0.1034354, 0.09607099, 0.122384, 0.1188784, 0.09039757,
  0.0987438, 0.1129893, 0.0968587, 0.05713516, 0.0604368, 0.056984, 
    0.1316232, 0.1441949, 0.08487441, 0.1129044, 0.07842243, 0.1345612, 
    0.1775137, 0.1441871, 0.1036659, 0.1952728, 0.17806, 0.2666411, 0.271909, 
    0.1177011, 0.08027682, 0.1064739, 0.1263155, 0.1631071, 0.1635741, 
    0.1389769, 0.1284936, 0.1603931, 0.1494623,
  0.2059242, 0.1950088, 0.1880829, 0.1783135, 0.1239255, 0.1214357, 0.121895, 
    0.1240003, 0.08932364, 0.101523, 0.08729117, 0.1148643, 0.1279971, 
    0.1393185, 0.1800835, 0.1546197, 0.1174391, 0.06286895, 0.07471278, 
    0.07998108, 0.1691295, 0.1536026, 0.2072741, 0.209529, 0.2055407, 
    0.2428847, 0.230391, 0.1877061, 0.2225311,
  0.1067659, 0.1627734, 0.2061649, 0.1506784, 0.1012122, 0.1328228, 
    0.1936301, 0.2042717, 0.1793827, 0.1828871, 0.1785841, 0.1775938, 
    0.2198718, 0.2165409, 0.1773572, 0.2120808, 0.2365365, 0.2160092, 
    0.2046511, 0.1896601, 0.1932292, 0.1869949, 0.2112987, 0.1223446, 
    0.2348343, 0.1885748, 0.1871149, 0.0906347, 0.09041736,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001482421, -0.000117395, 
    -8.654799e-05, -5.570093e-05, -2.485387e-05, 5.993184e-06, 3.684024e-05, 
    0.0001033376, 7.249058e-05, 4.164353e-05, 1.079647e-05, -2.005059e-05, 
    -5.089764e-05, -8.174471e-05, 0,
  0.003624043, -9.388837e-05, -1.152685e-06, 0, -4.935778e-06, 0.0001124593, 
    0, 0, -1.352915e-08, 0, -6.931259e-07, 4.333492e-05, 0.0003577148, 
    0.1077856, 0.1122556, 0.1326034, 0.131217, 0.1407473, 0.1148979, 
    0.03399453, 0.0291867, 0.02073267, 0.0879916, 0.2439053, 0.1745735, 
    0.1388514, 0.1832169, 0.1205542, 0.02425738,
  0.3004628, 0.3324716, 0.3145302, 0.2707589, 0.09286458, 0.04793213, 
    0.07032636, 0.02713743, 0.04679818, 0.07684694, 0.07073322, 0.09673063, 
    0.2757571, 0.2726012, 0.2792889, 0.2122778, 0.1522928, 0.2027497, 
    0.1864106, 0.2356559, 0.2936829, 0.2749813, 0.2441783, 0.2989302, 
    0.2218722, 0.150556, 0.1631601, 0.1505939, 0.2578407,
  0.2065196, 0.2107854, 0.2987807, 0.2707738, 0.2281302, 0.1974006, 
    0.1580909, 0.1969909, 0.1866151, 0.2206092, 0.2879571, 0.2936513, 
    0.2653222, 0.2377739, 0.2210272, 0.1728288, 0.2127077, 0.1427544, 
    0.1450859, 0.1744292, 0.2140648, 0.2474295, 0.2026024, 0.2457781, 
    0.19315, 0.2313971, 0.2310926, 0.1979389, 0.2190623,
  0.2533253, 0.2559178, 0.1822458, 0.1900362, 0.1649896, 0.1813977, 
    0.1670037, 0.1844195, 0.2391783, 0.2477423, 0.2195246, 0.2118411, 
    0.2077709, 0.1425521, 0.1224733, 0.1446162, 0.139103, 0.1616099, 
    0.1559564, 0.1939018, 0.2123786, 0.187192, 0.1911406, 0.1750289, 
    0.1319918, 0.161849, 0.241913, 0.2282783, 0.222616,
  0.1336309, 0.07852431, 0.05837632, 0.06565691, 0.06714138, 0.0964094, 
    0.09530354, 0.1173337, 0.09452619, 0.07873084, 0.09446684, 0.09730892, 
    0.07740115, 0.1019397, 0.09390859, 0.1222556, 0.1248447, 0.1507754, 
    0.1700606, 0.1689237, 0.1873408, 0.1511768, 0.1549532, 0.1715195, 
    0.04627153, 0.06606283, 0.09650648, 0.1429023, 0.1288273,
  0.01434381, 0.02057912, 0.03656069, 0.02793623, 0.04324728, 0.02659161, 
    0.01171402, 0.0102462, 0.0002573337, 0.00309659, 0.0003813707, 
    0.01303096, 0.03573358, 0.01970804, 0.05776844, 0.08857724, 0.1153535, 
    0.064337, 0.1311736, 0.05575242, 0.03280395, 0.01472908, 0.008425495, 
    0.00333019, 0.02681288, 0.0614414, 0.03296998, 0.05666604, 0.02996191,
  -3.809653e-07, 6.128995e-09, -7.928482e-06, 0.02103801, 0.02121175, 
    0.0002278999, 0.0127674, 0.00102561, -0.0002371327, 9.649317e-08, 
    1.109345e-07, 0.0002731185, 0.02085218, 0.07932612, 0.07170223, 
    0.02228084, 0.00535951, 0.01681462, -8.694462e-06, 1.897093e-05, 
    -1.400275e-05, 0.003786725, 6.028164e-08, 5.106753e-06, 0.0006332378, 
    0.0003975254, 0.001253318, 0.01300158, 0.001012903,
  2.346473e-07, 4.660708e-06, 1.938221e-05, 0.0005257804, 0.01228878, 
    0.01061208, 0.02274432, 0.09131324, 0.03385749, 0.006573722, 0.02585299, 
    0.01731405, 0.1141523, 0.1180812, 0.06832714, 0.02706727, 0.01769269, 
    0.0005526242, 5.366555e-05, 6.933495e-08, 5.721488e-08, 2.793111e-07, 
    7.007148e-06, 0.001075015, 2.480438e-05, 1.589918e-07, -3.210161e-06, 
    5.261905e-05, 5.975213e-08,
  0.01829796, 0.05391881, 0.06013314, 0.01872153, 0.001404935, 0.009446658, 
    0.0152552, 0.01733074, 0.07505042, 0.1555183, 0.04006886, 0.07653546, 
    0.09346478, 0.06642418, 0.06115072, 0.02221144, 0.01556986, 0.004972439, 
    0.01292569, 0.003605203, 0.004898299, 0.0007080456, 0.01246554, 
    0.06167441, 0.08358212, 0.07131368, 0.02831302, 0.00267339, 0.01064548,
  0.08094769, 0.1217932, 0.1253371, 0.3351014, 0.09721321, 0.02165597, 
    0.07105862, 0.02400042, 0.07881206, 0.0988485, 0.05068254, 0.09363762, 
    0.147519, 0.1054282, 0.07002646, 0.1042519, 0.08693293, 0.1252669, 
    0.1151402, 0.1661129, 0.3013256, 0.1403348, 0.1293436, 0.04861348, 
    0.04824022, 0.07095416, 0.1063625, 0.2057187, 0.1940463,
  0.006576936, 0.001485638, 5.915855e-05, 1.381661e-05, 0.04726269, 0.101087, 
    0.4766495, 0.1886692, 0.4132676, 0.05365606, 0.2392996, 0.1664691, 
    0.1035247, 0.05305791, 0.01082803, 0.003336335, 0.0003516521, 
    0.0001184359, 0.0043996, 0.02193897, 0.05529219, 0.02930753, 0.008210157, 
    0.05312008, 0.01519182, 0.008931503, 0.005217676, 0.006483575, 0.005960529,
  0.0009617939, 0.001935343, 3.965306e-08, 4.165913e-08, 0.0003598995, 
    0.0005601795, 0.0620768, 0.1680928, 0.2229287, 0.07528026, 0.05599635, 
    0.08801353, 0.2000627, 0.1396198, 0.07147463, 0.04625504, 0.01166183, 
    0.01290965, 0.004075434, 0.002243887, 0.06763034, 0.03477554, 0.07674912, 
    0.08431034, 0.02067264, 0.00324887, 0.01173349, 1.371431e-06, 0.003299282,
  0.03695775, 0.03327243, 0.009368485, 0.004798459, 0.01267637, 0.006248905, 
    0.1105963, 0.02426089, 0.05657429, 0.1332557, 0.09585073, 0.09942316, 
    0.159965, 0.2303266, 0.1444493, 0.07326946, 0.04870527, 0.05422204, 
    0.001231835, 0.0004109344, 0.06209046, 0.03675654, 0.05123584, 0.1116815, 
    0.09873942, 0.06804861, 0.04151057, 0.01323475, 0.003015535,
  0.03583662, 0.07638266, 0.03236292, 0.07501603, 0.06031771, 0.08730045, 
    0.07366743, 0.1411431, 0.1200931, 0.1232586, 0.06551076, 0.1139278, 
    0.1175084, 0.0821582, 0.1081314, 0.1402064, 0.1220759, 0.1662159, 
    0.1241248, 0.0544741, 0.04677356, 0.07425039, 0.08379494, 0.1095683, 
    0.09758212, 0.09132496, 0.1087582, 0.1094002, 0.09147872,
  0.1116198, 0.1210703, 0.09783839, 0.06142068, 0.06397285, 0.054345, 
    0.1455414, 0.1422365, 0.08416532, 0.1294253, 0.07439055, 0.1369418, 
    0.1922671, 0.1447455, 0.1180324, 0.1826933, 0.1734923, 0.2888608, 
    0.3087839, 0.1235314, 0.06609116, 0.09149098, 0.1312914, 0.1744919, 
    0.1482518, 0.164149, 0.09140432, 0.196145, 0.1474107,
  0.2171926, 0.1989444, 0.2017544, 0.1619033, 0.1243178, 0.1172843, 
    0.1254678, 0.1093836, 0.09388164, 0.1018603, 0.08731066, 0.112758, 
    0.1207063, 0.1420469, 0.1714003, 0.1801792, 0.141999, 0.07017756, 
    0.09141152, 0.07964535, 0.1733622, 0.1814378, 0.2320247, 0.2344225, 
    0.2291954, 0.2603894, 0.2327127, 0.164181, 0.1983607,
  0.08735756, 0.1386759, 0.1775299, 0.1351916, 0.1034451, 0.1412342, 
    0.2008931, 0.1890664, 0.1591002, 0.1574737, 0.163186, 0.1936239, 
    0.2078653, 0.216248, 0.1743007, 0.2224641, 0.2405721, 0.2168447, 
    0.2412688, 0.20063, 0.1859427, 0.1866577, 0.2488444, 0.1390398, 0.232085, 
    0.1795652, 0.1784093, 0.102036, 0.08794902,
  0.0008395411, 0.0004972518, 0.0001549626, -0.0001873267, -0.000529616, 
    -0.0008719052, -0.001214195, -1.464412e-06, -9.236419e-07, -3.82872e-07, 
    1.578978e-07, 6.986677e-07, 1.239438e-06, 1.780208e-06, -0.001218705, 
    -0.0008924623, -0.0005662197, -0.0002399772, 8.626538e-05, 0.0004125079, 
    0.0007387505, -0.001243727, -0.001228221, -0.001212715, -0.001197209, 
    -0.001181703, -0.001166197, -0.001150691, 0.001113373,
  0.01985512, -0.0007198136, 0.0012222, -2.891928e-05, -1.288778e-05, 
    0.001910756, 0.0002005361, -1.904936e-05, 9.595636e-06, 0.0001668213, 
    0.0006466793, 0.0007670497, 0.001211503, 0.1113588, 0.1178139, 0.1424642, 
    0.1300147, 0.1666875, 0.1703761, 0.06799958, 0.04523987, 0.04720246, 
    0.1430673, 0.2384469, 0.167688, 0.1445559, 0.2089235, 0.1819015, 
    0.05562595,
  0.3032437, 0.3454721, 0.3360969, 0.2983675, 0.1272666, 0.06102035, 
    0.08481588, 0.0430109, 0.0986938, 0.1477798, 0.1419984, 0.2048749, 
    0.3187296, 0.2806647, 0.2801765, 0.2155134, 0.1663719, 0.2062037, 
    0.2190001, 0.2629088, 0.3090008, 0.2951112, 0.2530845, 0.3100412, 
    0.219839, 0.1461239, 0.1585653, 0.1427618, 0.2689138,
  0.2076156, 0.2092371, 0.2932253, 0.265285, 0.2305706, 0.2111304, 0.1602464, 
    0.2129824, 0.1832804, 0.2040653, 0.276655, 0.2771066, 0.2589639, 0.23534, 
    0.1893451, 0.1642384, 0.212891, 0.1564789, 0.162212, 0.2011793, 
    0.2345145, 0.2493721, 0.1948924, 0.2415741, 0.1943749, 0.225924, 
    0.2209805, 0.1766284, 0.2175556,
  0.2648045, 0.2455307, 0.1791475, 0.1877084, 0.1657099, 0.1843098, 
    0.1593998, 0.1738522, 0.23571, 0.2357166, 0.2216648, 0.2134962, 
    0.2011343, 0.1563409, 0.1223731, 0.1363353, 0.1483252, 0.152217, 
    0.1700754, 0.1894405, 0.196179, 0.1936537, 0.1945619, 0.1622296, 
    0.1178589, 0.1641269, 0.2358902, 0.2450172, 0.2414733,
  0.1298176, 0.09312527, 0.06481269, 0.07303922, 0.06840177, 0.09456026, 
    0.1022369, 0.1186739, 0.09571265, 0.09486695, 0.1097084, 0.09749332, 
    0.08442545, 0.09933324, 0.09230468, 0.1100532, 0.1185031, 0.1461746, 
    0.1559648, 0.161737, 0.1794109, 0.1526028, 0.1407939, 0.1730052, 
    0.05246743, 0.06627486, 0.09344112, 0.148937, 0.1244955,
  0.01524422, 0.02147983, 0.04542257, 0.02765956, 0.04371351, 0.02761857, 
    0.01533051, 0.01692165, 0.002396262, 0.006721085, 0.01066224, 0.02219536, 
    0.04810005, 0.02337527, 0.0621546, 0.0784274, 0.1024762, 0.06954619, 
    0.128413, 0.06476514, 0.0374582, 0.02080528, 0.01860177, 0.005649237, 
    0.02780947, 0.07086785, 0.033342, 0.0675938, 0.03415604,
  4.711731e-05, -6.105328e-06, 1.522285e-05, 0.01433001, 0.02261478, 
    0.0002596217, 0.02256552, 0.00179462, -1.845466e-05, 1.824775e-07, 
    1.499699e-07, 0.001419845, 0.01517221, 0.069221, 0.0888015, 0.02218433, 
    0.006041204, 0.02105515, 0.004642633, 0.0008519624, -1.974254e-05, 
    0.006461458, 1.065865e-07, 2.576578e-06, 0.001119469, 0.0004561042, 
    0.006864295, 0.01083971, 1.759114e-05,
  3.040292e-07, 6.89416e-06, 0.0002204941, 0.0005990088, 0.01093698, 
    0.01530215, 0.02657032, 0.09170854, 0.03681024, 0.001645931, 0.02121644, 
    0.02791787, 0.1333181, 0.1294018, 0.06832608, 0.02736744, 0.02138423, 
    0.001420112, 9.639383e-05, 6.901207e-08, 5.24011e-08, 6.39553e-07, 
    8.994312e-06, 0.001609692, 1.520259e-05, 7.550564e-07, 5.887866e-06, 
    7.607769e-05, -1.540312e-06,
  0.02504814, 0.05174163, 0.09523114, 0.01529255, 0.001002734, 0.01084544, 
    0.02324055, 0.01979535, 0.1044632, 0.173492, 0.04788901, 0.09373967, 
    0.1015179, 0.07149898, 0.05968341, 0.02355044, 0.01266187, 0.004745639, 
    0.02006863, 0.001569317, 0.002294405, 0.0004142242, 0.01296757, 
    0.08232101, 0.09694459, 0.05253223, 0.0242452, 0.002752961, 0.01089698,
  0.09192371, 0.1540945, 0.1467791, 0.3804609, 0.07144614, 0.02908066, 
    0.09731679, 0.03874893, 0.08456135, 0.1099094, 0.06668051, 0.1035067, 
    0.1684987, 0.1197592, 0.0814282, 0.1101043, 0.1008156, 0.1375521, 
    0.1369122, 0.1992053, 0.3415344, 0.1594872, 0.1622182, 0.06858031, 
    0.0565386, 0.09116457, 0.1224168, 0.2454481, 0.2278414,
  0.003494003, 0.002617121, 0.002084799, 6.467273e-06, 0.02111363, 
    0.09362827, 0.5211805, 0.2110207, 0.4695361, 0.06046429, 0.2304712, 
    0.1748354, 0.1150072, 0.06213826, 0.01147624, 0.00514308, 0.0004539902, 
    4.537833e-05, 0.009670271, 0.008990155, 0.06652705, 0.0339676, 
    0.009401056, 0.05868944, 0.01649896, 0.005575133, 0.002571019, 
    0.006107674, 0.0007503018,
  7.32593e-05, 0.0002063312, 3.564464e-08, 4.394428e-08, 3.747908e-05, 
    0.0002110584, 0.06125027, 0.2086618, 0.2457106, 0.07565457, 0.0560837, 
    0.08731017, 0.2205712, 0.1668607, 0.07384673, 0.05250602, 0.01188733, 
    0.003987883, 0.001317813, 0.0004791731, 0.08571109, 0.04319734, 
    0.09179994, 0.101644, 0.02430686, 0.002668714, 0.00306247, 2.703577e-06, 
    0.0005139915,
  0.03654432, 0.0419007, 0.009292297, 0.00763121, 0.005109017, 0.003147511, 
    0.1112741, 0.01049869, 0.04015647, 0.1375716, 0.1105913, 0.09208813, 
    0.1931449, 0.2464977, 0.1634735, 0.06355313, 0.05116822, 0.05420841, 
    0.0009731553, 0.0005559886, 0.02302042, 0.04276913, 0.06018907, 
    0.1396923, 0.1137171, 0.079546, 0.04950846, 0.008596476, 0.01267186,
  0.04709091, 0.08252452, 0.03896023, 0.09388637, 0.05362458, 0.08679219, 
    0.07933051, 0.1437661, 0.1132695, 0.1182349, 0.07480665, 0.1306109, 
    0.1199839, 0.09239322, 0.1148994, 0.1616751, 0.1494925, 0.163504, 
    0.1515786, 0.05108365, 0.05026137, 0.07421286, 0.1008179, 0.1163175, 
    0.1022034, 0.1017421, 0.1142381, 0.1154531, 0.08721361,
  0.1320728, 0.1196304, 0.1079311, 0.05487011, 0.06065188, 0.06464091, 
    0.1530881, 0.1457112, 0.08963023, 0.1282838, 0.08333796, 0.1485981, 
    0.2064221, 0.1597256, 0.1350896, 0.203424, 0.2035889, 0.2924329, 
    0.3474377, 0.1411995, 0.06294599, 0.1037056, 0.1233269, 0.1555115, 
    0.1422864, 0.1572857, 0.1123281, 0.2119907, 0.1545866,
  0.229681, 0.2173142, 0.2021413, 0.1459952, 0.1064638, 0.1218909, 0.1399694, 
    0.1249743, 0.07708359, 0.1044335, 0.09993823, 0.1156541, 0.1488355, 
    0.1340575, 0.1998343, 0.1592059, 0.1268859, 0.0717326, 0.1004839, 
    0.08096185, 0.1711735, 0.188926, 0.2317927, 0.2612351, 0.2034993, 
    0.2563075, 0.2365935, 0.1689857, 0.2072138,
  0.09759372, 0.1411532, 0.2125071, 0.1777483, 0.1653654, 0.1951587, 
    0.2029722, 0.1955519, 0.1613981, 0.1587805, 0.1925646, 0.2272929, 
    0.2489105, 0.2197576, 0.1791787, 0.2072627, 0.2595665, 0.2259119, 
    0.1790906, 0.1379564, 0.1423487, 0.1746744, 0.2501529, 0.1310918, 
    0.2226124, 0.1695552, 0.1858183, 0.1125376, 0.09752092,
  0.01197243, 0.01060774, 0.009243046, 0.007878355, 0.006513663, 0.005148972, 
    0.00378428, 0.007036214, 0.00713328, 0.007230346, 0.007327411, 
    0.007424477, 0.007521543, 0.007618609, 0.004528041, 0.005685294, 
    0.006842546, 0.007999797, 0.009157049, 0.0103143, 0.01147155, 0.0130317, 
    0.01314207, 0.01325245, 0.01336282, 0.01347319, 0.01358357, 0.01369394, 
    0.01306418,
  0.02209516, 0.0009669908, 0.005081578, 0.003535157, 0.0009405504, 
    0.00540743, 0.001574058, 7.518596e-05, 0.0008374008, 0.003498282, 
    0.001376703, 0.000725204, 0.01391206, 0.1079721, 0.1418736, 0.1719205, 
    0.1344272, 0.1757421, 0.1805501, 0.1125431, 0.1134127, 0.09089538, 
    0.2013596, 0.2271633, 0.1760281, 0.1528571, 0.2193619, 0.2012225, 
    0.1035573,
  0.3187251, 0.354613, 0.3440591, 0.3130932, 0.1517505, 0.07133466, 
    0.08828934, 0.06435654, 0.1477854, 0.2038537, 0.2000037, 0.2869061, 
    0.3311089, 0.3116233, 0.2981572, 0.2258485, 0.1691288, 0.2326697, 
    0.2448955, 0.3045903, 0.3146514, 0.2772447, 0.2643422, 0.3250493, 
    0.2278074, 0.133416, 0.1491519, 0.1314292, 0.2589212,
  0.2207565, 0.2084435, 0.2956558, 0.2725709, 0.2245713, 0.2060772, 
    0.1828285, 0.2140493, 0.1899196, 0.2012538, 0.2706113, 0.2914691, 
    0.2524208, 0.2449651, 0.1836961, 0.178953, 0.2016144, 0.1498256, 
    0.1613434, 0.2070397, 0.2266272, 0.2847866, 0.2032841, 0.238808, 
    0.1909155, 0.2467115, 0.2222958, 0.1818738, 0.2326102,
  0.259721, 0.24494, 0.1851621, 0.1865011, 0.1860442, 0.1715211, 0.1769795, 
    0.203371, 0.2552454, 0.2456844, 0.2419978, 0.2185001, 0.1981571, 
    0.1511586, 0.1318941, 0.1385368, 0.1363819, 0.1564251, 0.1715114, 
    0.1896288, 0.1967262, 0.2032071, 0.1808207, 0.1605599, 0.120037, 
    0.1593622, 0.2396554, 0.2211765, 0.231352,
  0.1391982, 0.08258277, 0.07087482, 0.06911254, 0.0729104, 0.09778152, 
    0.1112054, 0.1329495, 0.1090168, 0.1026799, 0.1095122, 0.1044332, 
    0.08950588, 0.1133239, 0.09573123, 0.1087522, 0.1176666, 0.1456531, 
    0.1431357, 0.1678704, 0.1658993, 0.1519272, 0.1378066, 0.1740975, 
    0.0552179, 0.06847999, 0.0898587, 0.1478207, 0.1322523,
  0.01738691, 0.0244735, 0.05145758, 0.02951514, 0.04928048, 0.02750725, 
    0.02588102, 0.02261106, 0.005732509, 0.009694645, 0.03570326, 0.02428671, 
    0.06120208, 0.03530242, 0.06714357, 0.07232022, 0.09763322, 0.07004, 
    0.1307389, 0.07677649, 0.04579483, 0.0338558, 0.02649248, 0.006082583, 
    0.02861591, 0.08309646, 0.03930757, 0.07315579, 0.0329491,
  1.189832e-07, -4.042222e-05, 0.000203317, 0.01897993, 0.03266922, 
    0.007066914, 0.03125308, 0.003001044, 0.0001421927, -1.802798e-06, 
    5.708776e-05, 0.000740164, 0.02728306, 0.05433907, 0.09572738, 
    0.02468633, 0.01976811, 0.02670466, 0.01182964, 0.0009592707, 
    -1.643388e-05, 0.008308239, 7.340055e-08, 1.179882e-06, 0.002555917, 
    0.0007824691, 0.01352691, 0.006838523, -0.0001452093,
  3.468716e-07, 1.979255e-05, 0.000193025, 0.0007903191, 0.02067909, 
    0.02341574, 0.02786809, 0.09143747, 0.03840341, 0.001060239, 0.01698368, 
    0.04629037, 0.1313814, 0.1182218, 0.0692925, 0.03037952, 0.02867665, 
    0.003473941, 0.0001046122, 6.966963e-08, 1.030042e-07, 7.93391e-07, 
    1.021127e-05, 0.002905905, 2.492717e-05, 1.548154e-06, 0.00110036, 
    1.602369e-05, 9.58761e-08,
  0.01547972, 0.05413838, 0.129609, 0.008715017, 0.0005206033, 0.008568848, 
    0.02349043, 0.01610112, 0.0964033, 0.1848753, 0.04058643, 0.06554839, 
    0.08118905, 0.06329747, 0.05093414, 0.02091593, 0.005803194, 0.007998, 
    0.01703973, 0.003014905, 0.0004139364, 0.0005413322, 0.01674269, 
    0.1073068, 0.1130593, 0.03779439, 0.02587671, 0.007481904, 0.01367565,
  0.0759694, 0.1696377, 0.149329, 0.4269819, 0.02994874, 0.01854701, 
    0.09415913, 0.02923797, 0.04513866, 0.07876088, 0.03210765, 0.06831833, 
    0.122049, 0.09303409, 0.072441, 0.1044915, 0.1053729, 0.1266111, 
    0.1410927, 0.2025593, 0.3255317, 0.1366472, 0.1638982, 0.07629238, 
    0.04399949, 0.09870561, 0.1059723, 0.2228295, 0.2412647,
  0.0009202826, 0.0007049699, 0.003084726, 3.235707e-06, 0.0007992476, 
    0.07334064, 0.4209527, 0.1956834, 0.4940256, 0.06050478, 0.1917354, 
    0.1430721, 0.08343714, 0.0536881, 0.01457414, 0.006158646, 0.000786202, 
    -6.424393e-06, 0.005960269, 0.001536972, 0.04162046, 0.03191712, 
    0.008493351, 0.05112408, 0.01490495, 0.003686293, 0.001415747, 
    0.004671589, 0.0002892917,
  2.495678e-05, 2.653908e-05, 1.638885e-08, 3.818273e-08, 1.487518e-05, 
    0.0002707784, 0.06753857, 0.265729, 0.2868098, 0.07398618, 0.05367191, 
    0.06889877, 0.1914337, 0.1532438, 0.07273863, 0.04949841, 0.007821437, 
    0.0006280557, 0.0006711656, 0.0001243806, 0.07146204, 0.03502401, 
    0.07056413, 0.09243178, 0.02071666, 0.002287666, 0.0005675643, 
    3.976745e-06, 0.000233859,
  0.03552385, 0.02671048, 0.01963921, 0.01074648, 0.00670248, 0.0009696411, 
    0.09476401, 0.005011234, 0.02859705, 0.1382538, 0.1092156, 0.08194749, 
    0.205152, 0.25146, 0.1877911, 0.06872357, 0.06948524, 0.05136175, 
    0.002701621, 0.0007455861, 0.009036665, 0.04199475, 0.06982372, 
    0.1482916, 0.117407, 0.07388484, 0.07962333, 0.0152996, 0.01508086,
  0.04417716, 0.08864125, 0.04270535, 0.09585692, 0.07641544, 0.09004398, 
    0.08533253, 0.1481803, 0.09852806, 0.1124175, 0.08417238, 0.1631107, 
    0.1319764, 0.1039108, 0.1349258, 0.18143, 0.1642996, 0.179635, 0.1556567, 
    0.05137958, 0.05871257, 0.07685544, 0.1198357, 0.1319928, 0.1025566, 
    0.1148363, 0.1190939, 0.1310902, 0.08291108,
  0.1269551, 0.1291656, 0.1269796, 0.07473311, 0.0782295, 0.07314364, 
    0.1578405, 0.1463052, 0.09875275, 0.1449994, 0.09537231, 0.1559707, 
    0.229974, 0.1810031, 0.1416737, 0.2465228, 0.1847102, 0.3344792, 
    0.3294988, 0.1376785, 0.06761789, 0.1171802, 0.132493, 0.176348, 
    0.1497165, 0.1493292, 0.08296818, 0.1884184, 0.1501546,
  0.237212, 0.1877133, 0.2021758, 0.1628762, 0.1217477, 0.1118423, 0.1468986, 
    0.1453518, 0.0811753, 0.09854142, 0.1012371, 0.1179462, 0.1318178, 
    0.14512, 0.2010704, 0.1733002, 0.1296732, 0.08049931, 0.07953633, 
    0.08538386, 0.1536609, 0.2130086, 0.2307472, 0.2469661, 0.2235573, 
    0.2822077, 0.2298834, 0.1676013, 0.1950062,
  0.08742815, 0.1297539, 0.192896, 0.1681977, 0.155801, 0.1606588, 0.1995293, 
    0.1820394, 0.1733443, 0.1621287, 0.2148904, 0.2606534, 0.2343236, 
    0.1907879, 0.1801759, 0.2283267, 0.1967531, 0.2140628, 0.1916612, 
    0.1106478, 0.1376172, 0.1784045, 0.2461316, 0.1272125, 0.1904334, 
    0.1903542, 0.1909029, 0.1278268, 0.07713655,
  0.02519479, 0.02431544, 0.02343608, 0.02255673, 0.02167738, 0.02079803, 
    0.01991868, 0.01984838, 0.01954909, 0.0192498, 0.01895051, 0.01865122, 
    0.01835193, 0.01805265, 0.02108839, 0.02242001, 0.02375162, 0.02508324, 
    0.02641486, 0.02774648, 0.0290781, 0.02485701, 0.02470404, 0.02455106, 
    0.02439808, 0.0242451, 0.02409213, 0.02393915, 0.02589827,
  0.05440208, 0.02059205, 0.02303825, 0.01676344, 0.01257829, 0.01941518, 
    0.01414061, 0.01574136, 0.007953998, 0.006920068, 0.006588819, 
    0.006832733, 0.03140704, 0.09704886, 0.1259976, 0.1471812, 0.1509159, 
    0.1938159, 0.1928457, 0.1516015, 0.1776972, 0.2193479, 0.2405805, 
    0.2268838, 0.1772324, 0.1616071, 0.2291335, 0.2034065, 0.1465675,
  0.3383129, 0.3712994, 0.3547804, 0.3248687, 0.1778333, 0.08272129, 
    0.09021077, 0.1160846, 0.2012419, 0.2436005, 0.2741891, 0.3343874, 
    0.3203049, 0.3303209, 0.2956414, 0.2521849, 0.1986485, 0.2544367, 
    0.2779947, 0.3387077, 0.3415267, 0.3378398, 0.2688674, 0.3809208, 
    0.2460284, 0.150613, 0.1781911, 0.1452481, 0.2892119,
  0.2531083, 0.2229791, 0.3037502, 0.2604979, 0.2218518, 0.2253819, 
    0.1749843, 0.2558889, 0.2443919, 0.2210875, 0.2825667, 0.280552, 
    0.2449595, 0.2437481, 0.1973727, 0.1791429, 0.2014182, 0.1766082, 
    0.183641, 0.2278306, 0.2530245, 0.2719839, 0.2211415, 0.2696846, 
    0.1944897, 0.2578363, 0.2204837, 0.1849314, 0.2396725,
  0.2588488, 0.2341064, 0.1904663, 0.1991715, 0.1805445, 0.1828952, 0.210085, 
    0.2294158, 0.2743786, 0.2548474, 0.26642, 0.2155897, 0.2106422, 
    0.1750499, 0.1506434, 0.1432844, 0.1368496, 0.1489721, 0.1984395, 
    0.1829138, 0.1984361, 0.2043938, 0.1803145, 0.1573571, 0.1145533, 
    0.15843, 0.2388079, 0.2171273, 0.2342816,
  0.155149, 0.0922613, 0.07424953, 0.07387773, 0.07962376, 0.116741, 
    0.1175616, 0.1318893, 0.1238124, 0.1209885, 0.1104812, 0.1200854, 
    0.1008173, 0.1102714, 0.1007634, 0.1165496, 0.1316519, 0.1534623, 
    0.1414452, 0.1600409, 0.1750802, 0.1519479, 0.1296023, 0.172029, 
    0.06033392, 0.07567777, 0.09529343, 0.160256, 0.1383308,
  0.02280967, 0.03052033, 0.06428678, 0.03085904, 0.05637475, 0.03019456, 
    0.03633972, 0.03309327, 0.007430617, 0.01174815, 0.03046889, 0.01523608, 
    0.07572104, 0.04879504, 0.07650125, 0.07151788, 0.09465992, 0.07517457, 
    0.1398556, 0.09616674, 0.05826171, 0.04228297, 0.02817415, 0.006028671, 
    0.04294973, 0.09515559, 0.04794042, 0.08278844, 0.04056495,
  8.116453e-08, 0.0007590418, 0.001773881, 0.02361943, 0.04155529, 
    0.008164095, 0.04261234, 0.005252603, 0.01391876, -1.156595e-05, 
    0.001212466, -0.0003981222, 0.02634147, 0.05040116, 0.09662011, 
    0.03152837, 0.02318397, 0.0224183, 0.02363607, 0.003764126, 0.0007903031, 
    0.008556847, 1.784059e-07, 6.889571e-07, 0.005747811, 0.003472452, 
    0.03380106, 0.009215295, 0.0007345206,
  2.526023e-07, -0.0001486136, 0.0003988828, 0.005248556, 0.02353667, 
    0.02933594, 0.02391278, 0.08048798, 0.03964917, 0.001001139, 0.01284512, 
    0.05172711, 0.1425868, 0.109538, 0.0665004, 0.03492332, 0.03248614, 
    0.006030621, 0.0002234454, 1.103245e-06, 1.654937e-07, 2.256438e-06, 
    2.479955e-05, 0.004007962, 0.001285722, 0.0005477667, 0.006054245, 
    2.17321e-05, 1.210431e-07,
  0.006613043, 0.04834189, 0.1157831, 0.01267851, 0.000513549, 0.007498223, 
    0.02190451, 0.01601424, 0.07615887, 0.1530738, 0.03915682, 0.04673529, 
    0.06787077, 0.05728288, 0.04489555, 0.02281831, 0.007733332, 0.0116313, 
    0.01444494, 0.002091519, 0.0003649761, 0.0004844033, 0.02253959, 
    0.1153039, 0.1302625, 0.02825638, 0.02216768, 0.01251375, 0.006672033,
  0.04527806, 0.1036331, 0.08426344, 0.469952, 0.01206941, 0.00972344, 
    0.09056561, 0.02629369, 0.02181557, 0.05187167, 0.01630747, 0.05075284, 
    0.09718433, 0.07562339, 0.06521432, 0.09514496, 0.1015756, 0.1239811, 
    0.1453672, 0.2061344, 0.2894263, 0.1220581, 0.1399577, 0.06833203, 
    0.03081662, 0.0829604, 0.09774849, 0.183478, 0.1916905,
  0.000150631, 0.0001112119, 0.0006279635, 1.235441e-06, 4.040334e-05, 
    0.04448915, 0.346596, 0.1997606, 0.4131761, 0.06758463, 0.1687149, 
    0.1216543, 0.06682371, 0.03572044, 0.0189636, 0.01201635, 0.0004959747, 
    0.0002059131, 0.008555464, 0.0001355733, 0.03332748, 0.0318378, 
    0.00824687, 0.03617955, 0.01562923, 0.002453191, 0.0009660602, 
    0.0009826537, 0.0001599448,
  1.095304e-05, 1.135615e-05, -4.865905e-09, 2.87566e-08, 4.536782e-06, 
    0.0001344729, 0.0622422, 0.278581, 0.3382595, 0.07684422, 0.05549885, 
    0.05454966, 0.1458586, 0.09269916, 0.06552161, 0.04205437, 0.003938975, 
    7.72106e-06, 0.00059999, 9.520007e-06, 0.03125399, 0.02126731, 
    0.06329463, 0.05048787, 0.01088773, 0.002538234, 0.0003268434, 
    2.670648e-06, 1.330155e-05,
  0.03479557, 0.01875679, 0.02485737, 0.01317856, 0.004448946, 0.002812296, 
    0.06590226, 0.0009750898, 0.01911246, 0.1063093, 0.09734862, 0.0765698, 
    0.1884734, 0.2424757, 0.1722325, 0.08577874, 0.07371712, 0.06513628, 
    0.001738006, 0.000352058, 0.003178078, 0.02816611, 0.06313934, 0.1185717, 
    0.105765, 0.0776018, 0.05384277, 0.01717945, 0.009276404,
  0.06041699, 0.1021258, 0.05028386, 0.1145544, 0.07429425, 0.08654819, 
    0.08696218, 0.177572, 0.09599635, 0.1105333, 0.0910415, 0.1622813, 
    0.1177896, 0.1219509, 0.1293517, 0.2141889, 0.1980995, 0.2178311, 
    0.175846, 0.05855974, 0.06494638, 0.0687693, 0.1204928, 0.1471044, 
    0.1031091, 0.1122792, 0.1255984, 0.1464584, 0.09577002,
  0.1631912, 0.1531613, 0.1311705, 0.09516487, 0.1143294, 0.08080551, 
    0.1704601, 0.1607114, 0.1151537, 0.1677212, 0.1276418, 0.182306, 
    0.253185, 0.1847796, 0.1505832, 0.265485, 0.1846605, 0.3581184, 0.337834, 
    0.1319474, 0.083281, 0.1407821, 0.1502267, 0.1779148, 0.1503391, 
    0.1640243, 0.1198264, 0.1916973, 0.1919588,
  0.2229498, 0.2158934, 0.2334865, 0.1758559, 0.1349458, 0.1139754, 
    0.1350941, 0.1274468, 0.09420942, 0.1067382, 0.1183482, 0.1598123, 
    0.1383467, 0.1477447, 0.1887445, 0.1324136, 0.1288847, 0.09956345, 
    0.08552088, 0.09351495, 0.1840507, 0.1969866, 0.265773, 0.2567979, 
    0.1960004, 0.3243854, 0.2743718, 0.1843556, 0.2269472,
  0.1356579, 0.1468957, 0.2402868, 0.1853112, 0.1828031, 0.1793089, 
    0.2278446, 0.2113459, 0.1835904, 0.1396302, 0.204261, 0.2314708, 
    0.2443391, 0.1954965, 0.1675218, 0.1592752, 0.2064742, 0.1978485, 
    0.1999952, 0.1365848, 0.1581923, 0.1672594, 0.2394295, 0.1399394, 
    0.1971091, 0.169297, 0.1777884, 0.1354787, 0.1251756,
  0.04534409, 0.04345874, 0.04157339, 0.03968804, 0.03780269, 0.03591734, 
    0.03403199, 0.03652577, 0.03636635, 0.03620693, 0.03604751, 0.03588809, 
    0.03572867, 0.03556925, 0.03115585, 0.03374503, 0.03633421, 0.03892339, 
    0.04151257, 0.04410176, 0.04669094, 0.03908803, 0.03854362, 0.03799921, 
    0.0374548, 0.03691039, 0.03636597, 0.03582157, 0.04685237,
  0.1037035, 0.04646025, 0.04710757, 0.03363974, 0.01939406, 0.03350266, 
    0.0252037, 0.03058842, 0.0179648, 0.02469001, 0.007517782, 0.02055088, 
    0.04843301, 0.0903734, 0.1062548, 0.1607791, 0.1729825, 0.2005058, 
    0.1904807, 0.1713867, 0.216072, 0.3145536, 0.2677806, 0.2239454, 
    0.187652, 0.1585836, 0.2495901, 0.2048783, 0.1571197,
  0.3866152, 0.4104502, 0.3561192, 0.3466551, 0.2090122, 0.07686964, 
    0.1022808, 0.1337478, 0.2460351, 0.2653879, 0.3029401, 0.3835962, 
    0.3094211, 0.3453058, 0.2901092, 0.2301022, 0.1779323, 0.2448323, 
    0.2837168, 0.3311572, 0.3457514, 0.3306856, 0.2779583, 0.3893365, 
    0.2423142, 0.1437815, 0.1759682, 0.1556767, 0.3090227,
  0.2540747, 0.2272369, 0.303331, 0.2764379, 0.2628417, 0.2501455, 0.2052671, 
    0.2766109, 0.2741711, 0.2450276, 0.3012986, 0.3078213, 0.2843589, 
    0.2711206, 0.2590408, 0.2125958, 0.2264494, 0.2042006, 0.2155848, 
    0.2568396, 0.3036112, 0.291669, 0.2144455, 0.324788, 0.1991801, 
    0.2735857, 0.2510537, 0.219641, 0.2245988,
  0.2887922, 0.2599576, 0.2186722, 0.2109117, 0.1984003, 0.1962738, 
    0.2141833, 0.2499612, 0.2772611, 0.2565618, 0.2707546, 0.2195545, 
    0.2328088, 0.1938244, 0.1471005, 0.1573281, 0.1554736, 0.1858753, 
    0.2031468, 0.1744744, 0.2083639, 0.2023743, 0.1903422, 0.1670611, 
    0.1321394, 0.1761326, 0.246678, 0.2335318, 0.2792518,
  0.1697822, 0.1087266, 0.08999779, 0.07736315, 0.08934788, 0.1347976, 
    0.1402112, 0.1465742, 0.132608, 0.1350621, 0.1255498, 0.1339062, 
    0.1163747, 0.1152044, 0.1096148, 0.1323513, 0.1471756, 0.1575501, 
    0.1558988, 0.1597855, 0.1796441, 0.171322, 0.1301289, 0.1764806, 
    0.06070203, 0.08385596, 0.1203274, 0.1781059, 0.1592895,
  0.04026543, 0.03600301, 0.0773708, 0.03237657, 0.06234017, 0.03115851, 
    0.04344392, 0.04682224, 0.01767103, 0.01544742, 0.02321664, 0.005288553, 
    0.09239417, 0.06315135, 0.09142461, 0.07433598, 0.09973057, 0.08250079, 
    0.1446583, 0.1033946, 0.07619646, 0.06534608, 0.02955061, 0.005970079, 
    0.0599584, 0.1180009, 0.06307675, 0.08975329, 0.05204868,
  -2.671141e-06, -1.535371e-05, 0.01838563, 0.03724941, 0.0578748, 
    0.02609479, 0.04605545, 0.01168715, 0.02547573, 0.02882159, 
    -4.667818e-06, 0.004465893, 0.02485007, 0.06206617, 0.08447491, 
    0.0584466, 0.04022341, 0.0174343, 0.03350374, 0.01562535, 0.003444596, 
    0.007214532, 1.448304e-06, 5.236494e-07, 0.01378238, 0.01534873, 
    0.04066177, 0.02185661, 0.005601971,
  1.586642e-07, -3.940775e-05, 0.0006846468, 0.03047432, 0.03421658, 
    0.0363614, 0.02301857, 0.07577014, 0.03880896, 0.002165058, 0.02305145, 
    0.05424191, 0.1636713, 0.1103912, 0.06902753, 0.04211541, 0.04292735, 
    0.01700846, 0.002446747, 0.0001001359, 6.826581e-07, 1.24053e-06, 
    4.597669e-06, 0.0074193, 0.04848693, 0.0186523, 0.0290074, 6.797558e-05, 
    3.615858e-07,
  0.0006112078, 0.04255466, 0.1175611, 0.02094707, 0.001081617, 0.007447607, 
    0.02057863, 0.01616227, 0.06835882, 0.1374763, 0.04172193, 0.03594901, 
    0.06142773, 0.0520282, 0.04209648, 0.03363111, 0.01603133, 0.006043512, 
    0.01380223, 0.0009247169, 0.0005380486, 0.001456816, 0.02996011, 
    0.1383936, 0.1531044, 0.03194946, 0.01553017, 0.005536393, 0.003510462,
  0.04220494, 0.06959022, 0.05172265, 0.462798, 0.007237816, 0.006440459, 
    0.08891191, 0.02720221, 0.01631197, 0.03397801, 0.01155763, 0.04139755, 
    0.08020221, 0.06360088, 0.06509651, 0.09283728, 0.09669228, 0.1279251, 
    0.1465307, 0.2059487, 0.2648637, 0.1136098, 0.1364946, 0.06256092, 
    0.02232729, 0.07700348, 0.09825055, 0.1691094, 0.1755484,
  3.45934e-05, 1.888986e-05, 6.395539e-06, 5.327715e-07, 5.270083e-07, 
    0.02629585, 0.290575, 0.2199987, 0.3998069, 0.07542863, 0.1542481, 
    0.1091963, 0.05641854, 0.03226473, 0.02301279, 0.0224738, 0.0009272288, 
    0.001694738, 0.01127371, 3.199573e-05, 0.02919568, 0.03675, 0.008709634, 
    0.02926518, 0.01803405, 0.003424709, 0.0005467217, 0.0001760404, 
    8.335795e-05,
  4.899682e-06, 5.623832e-06, 1.302337e-06, 1.310378e-08, 1.251174e-06, 
    4.334092e-05, 0.05373762, 0.2877379, 0.3596094, 0.08161961, 0.06140515, 
    0.04486796, 0.117599, 0.06570943, 0.05367707, 0.02676663, 0.00498665, 
    -2.697141e-05, 0.0001973912, 1.08187e-06, 0.009183008, 0.02317114, 
    0.06552058, 0.03194945, 0.009238206, 0.003732004, 0.001138766, 
    5.503407e-06, 6.134126e-06,
  0.02492068, 0.01847716, 0.02480895, 0.02186858, 0.001592862, 0.001662441, 
    0.03668669, 4.337698e-05, 0.0114046, 0.08382566, 0.09532727, 0.07673424, 
    0.1808817, 0.2112444, 0.1358068, 0.1010766, 0.07572775, 0.06061564, 
    0.01058795, 0.0001398981, 0.001489684, 0.01810322, 0.06574076, 0.1173074, 
    0.09508814, 0.0595854, 0.03866601, 0.01533886, 0.002366385,
  0.05969901, 0.1218847, 0.05904173, 0.1193483, 0.06492971, 0.08318692, 
    0.08209018, 0.1821088, 0.1051896, 0.09718929, 0.07308143, 0.1652364, 
    0.08881452, 0.1098674, 0.1418729, 0.230413, 0.2100079, 0.2242275, 
    0.1835259, 0.0731463, 0.07328205, 0.05776435, 0.1159936, 0.1689747, 
    0.1160208, 0.1152536, 0.1124324, 0.1412412, 0.09009706,
  0.1801012, 0.1903448, 0.1529201, 0.1317043, 0.1128423, 0.07799882, 
    0.1662076, 0.1933481, 0.1352347, 0.1837881, 0.1448446, 0.2138679, 
    0.2800452, 0.1925887, 0.1550519, 0.2911373, 0.2001879, 0.3903068, 
    0.3751693, 0.1436987, 0.1213012, 0.1825921, 0.1666525, 0.2014731, 
    0.1662037, 0.173755, 0.1242458, 0.1934772, 0.2108702,
  0.2585839, 0.233766, 0.2800903, 0.2200351, 0.173168, 0.118589, 0.1904164, 
    0.1420842, 0.1275961, 0.1232124, 0.1452796, 0.1910097, 0.1491736, 
    0.1684722, 0.2094011, 0.1467363, 0.152782, 0.09950511, 0.1011904, 
    0.1188368, 0.1802661, 0.1959095, 0.2329612, 0.2514108, 0.1862974, 
    0.3149617, 0.2747627, 0.1948234, 0.260007,
  0.1295816, 0.1826546, 0.2844512, 0.1946472, 0.1746096, 0.1587046, 
    0.2075089, 0.2221446, 0.1757355, 0.1329997, 0.1810609, 0.2240897, 
    0.2331807, 0.224327, 0.1953129, 0.195544, 0.2185483, 0.1952609, 
    0.1872726, 0.0926844, 0.1401831, 0.1724648, 0.2321156, 0.1158023, 
    0.1569012, 0.1609011, 0.174814, 0.1440143, 0.1258702,
  0.08799879, 0.08283213, 0.07766547, 0.07249881, 0.06733216, 0.0621655, 
    0.05699884, 0.06627027, 0.06789044, 0.06951062, 0.0711308, 0.07275098, 
    0.07437116, 0.07599133, 0.08310217, 0.08756315, 0.09202413, 0.09648511, 
    0.1009461, 0.1054071, 0.109868, 0.1170128, 0.1160983, 0.1151838, 
    0.1142693, 0.1133548, 0.1124403, 0.1115258, 0.09213211,
  0.1206765, 0.07544303, 0.06934929, 0.03439611, 0.0282745, 0.04526365, 
    0.03524923, 0.03831019, 0.03137563, 0.03352569, 0.02313247, 0.02691239, 
    0.05174129, 0.08120294, 0.08844616, 0.147416, 0.1729626, 0.197003, 
    0.1727092, 0.1650564, 0.2381523, 0.3451118, 0.278194, 0.2172908, 
    0.1877739, 0.1577035, 0.2649368, 0.2056656, 0.1706964,
  0.4080946, 0.4419982, 0.3713582, 0.3431622, 0.2179247, 0.07104354, 
    0.1016868, 0.1665596, 0.2716853, 0.2794996, 0.3172261, 0.4002928, 
    0.3054351, 0.3164405, 0.2550164, 0.1859214, 0.1603464, 0.2731915, 
    0.2524518, 0.2907572, 0.322331, 0.2845524, 0.2460247, 0.3450614, 
    0.2186884, 0.1313199, 0.1567606, 0.1845491, 0.3233244,
  0.2425201, 0.2230296, 0.3095685, 0.2778983, 0.2847422, 0.2638036, 
    0.1729345, 0.2559702, 0.2795216, 0.2606049, 0.2734386, 0.3207411, 
    0.2745794, 0.2623329, 0.2764705, 0.2717292, 0.2536247, 0.2198257, 
    0.2378698, 0.2857755, 0.3128208, 0.3020692, 0.2219821, 0.3288188, 
    0.2123692, 0.2595527, 0.2414472, 0.2295924, 0.2262811,
  0.2844924, 0.2800123, 0.2382806, 0.2299504, 0.2240035, 0.2330761, 
    0.2336293, 0.2877899, 0.2802695, 0.2727112, 0.2733695, 0.2264575, 
    0.2290226, 0.2033993, 0.1837116, 0.1782917, 0.1764496, 0.197083, 
    0.241449, 0.1793319, 0.2037651, 0.230297, 0.188893, 0.1796877, 0.1291387, 
    0.18289, 0.2749476, 0.2481798, 0.2872154,
  0.1807895, 0.1320447, 0.108602, 0.101816, 0.1100555, 0.1589357, 0.1663399, 
    0.1729181, 0.1651639, 0.1468514, 0.1487278, 0.1518342, 0.1163067, 
    0.1323181, 0.1222117, 0.1600524, 0.1647778, 0.1738018, 0.1794715, 
    0.1738362, 0.1914003, 0.1912398, 0.1513456, 0.1939582, 0.05731703, 
    0.1049619, 0.1466249, 0.20097, 0.185697,
  0.05896612, 0.03964099, 0.08373474, 0.03833459, 0.06048203, 0.04056244, 
    0.04844974, 0.0482518, 0.03767917, 0.02749681, 0.0256164, 0.003997027, 
    0.08949182, 0.07058388, 0.1025627, 0.08460315, 0.1126987, 0.07807803, 
    0.1472474, 0.1115163, 0.07985067, 0.08123754, 0.03331066, 0.006332465, 
    0.06034376, 0.1120718, 0.08825947, 0.09801373, 0.06813141,
  9.762296e-05, -3.780163e-06, 0.06563717, 0.04619906, 0.07739796, 
    0.04257574, 0.05361756, 0.02030947, 0.03415401, 0.02374594, 
    -6.025947e-05, 0.006257042, 0.02026632, 0.06931528, 0.08065623, 
    0.06441513, 0.03708502, 0.01847059, 0.04161828, 0.04901634, 0.01323258, 
    0.008287642, -1.8112e-05, 3.820474e-06, 0.01525016, 0.02560648, 
    0.0671454, 0.03913226, 0.007563794,
  9.87789e-08, -3.580979e-05, 0.004420651, 0.1117715, 0.04209846, 0.03925716, 
    0.02765638, 0.07452554, 0.0413225, 0.005806367, 0.04108656, 0.05488572, 
    0.1853857, 0.1149881, 0.06857806, 0.04405956, 0.04946669, 0.02591097, 
    0.01230402, 0.002825664, 0.0001199798, 1.907466e-07, 6.681857e-07, 
    0.009114181, 0.0375604, 0.01662819, 0.06919134, 0.001413076, 0.000108951,
  7.954908e-05, 0.04112974, 0.1012142, 0.03452192, 0.005581953, 0.0107241, 
    0.01810893, 0.01678869, 0.05421819, 0.1358035, 0.04390974, 0.03226011, 
    0.05438139, 0.0465242, 0.04176388, 0.04329488, 0.01806832, 0.005462116, 
    0.009833975, 0.0002418183, 0.0001471279, 0.002343617, 0.02498009, 
    0.1667064, 0.1504561, 0.02536866, 0.01774101, 0.003714388, 0.001489794,
  0.04212467, 0.0491542, 0.03673997, 0.385947, 0.005472474, 0.00720636, 
    0.08283196, 0.02943417, 0.01426671, 0.02435314, 0.01257088, 0.03613149, 
    0.06907944, 0.05540461, 0.06802602, 0.09452317, 0.09580225, 0.1381212, 
    0.1558821, 0.1955438, 0.2496304, 0.1139824, 0.1356848, 0.06644887, 
    0.02089532, 0.0774329, 0.110834, 0.1690538, 0.1620603,
  8.014408e-06, 3.302243e-07, 4.575639e-07, 1.549732e-07, 1.639631e-07, 
    0.0102622, 0.2661087, 0.2353285, 0.3788802, 0.08211672, 0.1456272, 
    0.1035185, 0.04937953, 0.02766901, 0.02303529, 0.03008866, 0.006622201, 
    0.004464117, 0.01400474, 3.85625e-05, 0.0298737, 0.04416395, 0.01077566, 
    0.02369943, 0.02447907, 0.008561159, 0.0007858832, 2.080183e-05, 
    4.519075e-05,
  2.333949e-06, 3.156422e-06, -3.856888e-07, 4.047041e-09, 5.841357e-07, 
    1.909707e-05, 0.0448553, 0.30474, 0.3532411, 0.09014053, 0.0654247, 
    0.04062191, 0.1015613, 0.04838759, 0.05030333, 0.02571188, 0.007662487, 
    0.0004700924, 1.574124e-06, 4.406195e-07, 0.002611137, 0.01583447, 
    0.06314868, 0.02370027, 0.01147933, 0.01135945, 0.001937264, 
    6.775991e-05, 4.694107e-06,
  0.01432223, 0.01469246, 0.02111023, 0.02974823, -9.886061e-05, 
    8.455729e-05, 0.01987732, 1.13002e-05, 0.006436381, 0.05857222, 
    0.1029689, 0.08416937, 0.18863, 0.2081478, 0.1235455, 0.1049165, 
    0.07296234, 0.04998044, 0.0204445, 0.0001018406, 0.0003258429, 
    0.01128229, 0.06875427, 0.1129837, 0.09047771, 0.05879845, 0.03208923, 
    0.01320846, 0.007356838,
  0.05404811, 0.1285928, 0.06160183, 0.109193, 0.03282862, 0.06951366, 
    0.09156314, 0.1938532, 0.1229218, 0.07621687, 0.0668595, 0.160039, 
    0.09215623, 0.1193838, 0.1388903, 0.2227782, 0.2549258, 0.2378762, 
    0.2046089, 0.08890979, 0.06762523, 0.05216755, 0.1105612, 0.1861419, 
    0.1375649, 0.1267492, 0.1137193, 0.1460839, 0.09067734,
  0.1869945, 0.2088919, 0.1570811, 0.1219275, 0.1247845, 0.09556184, 
    0.179954, 0.2207778, 0.128488, 0.1842479, 0.1353643, 0.2506888, 
    0.2905474, 0.1991901, 0.1398537, 0.3343588, 0.2413116, 0.419424, 
    0.3979386, 0.1583186, 0.1433916, 0.1838746, 0.1666985, 0.2434489, 
    0.1797955, 0.1911401, 0.1580986, 0.2197964, 0.2425022,
  0.2607725, 0.277209, 0.3162911, 0.2155594, 0.1644556, 0.1629199, 0.2032179, 
    0.1680653, 0.1780321, 0.1700165, 0.1551674, 0.2189602, 0.1766347, 
    0.1966071, 0.2345176, 0.1550209, 0.190501, 0.1079671, 0.1272086, 
    0.1282273, 0.1738968, 0.2117887, 0.2229754, 0.264662, 0.1912959, 
    0.305829, 0.2327801, 0.2079919, 0.2883412,
  0.1395209, 0.2104392, 0.2646813, 0.2279001, 0.1841394, 0.1801985, 
    0.2345834, 0.2565883, 0.236231, 0.2019743, 0.1883571, 0.2269476, 
    0.2668863, 0.2580527, 0.2347381, 0.2202741, 0.2373244, 0.2336987, 
    0.1906341, 0.100614, 0.1363635, 0.1953079, 0.2311392, 0.1101292, 
    0.1450158, 0.141237, 0.1440566, 0.1365709, 0.1599946,
  0.1774418, 0.1734846, 0.1695274, 0.1655701, 0.1616129, 0.1576557, 
    0.1536984, 0.1535153, 0.1542013, 0.1548873, 0.1555733, 0.1562593, 
    0.1569453, 0.1576314, 0.1538413, 0.1575649, 0.1612885, 0.1650121, 
    0.1687357, 0.1724593, 0.1761829, 0.1694759, 0.1690235, 0.1685712, 
    0.1681188, 0.1676664, 0.1672141, 0.1667617, 0.1806076,
  0.1322241, 0.1147236, 0.07926299, 0.04126721, 0.03826257, 0.04809551, 
    0.06723758, 0.06388629, 0.04746456, 0.0432979, 0.0386271, 0.02931857, 
    0.05045739, 0.0797094, 0.1068561, 0.1339823, 0.1403061, 0.1671431, 
    0.1574549, 0.1889612, 0.26086, 0.3782772, 0.3012548, 0.2255762, 
    0.1878063, 0.1655318, 0.2504834, 0.2107812, 0.1740332,
  0.4173053, 0.4384088, 0.3864378, 0.3470426, 0.2132567, 0.07417712, 
    0.1148991, 0.1918787, 0.2892382, 0.2812231, 0.3306343, 0.407066, 
    0.2986407, 0.3180883, 0.2655235, 0.1725104, 0.1632015, 0.2428997, 
    0.2437555, 0.279012, 0.3039727, 0.2695749, 0.2314582, 0.3335217, 
    0.1954302, 0.1177095, 0.1424216, 0.1942533, 0.3565082,
  0.2385785, 0.2414813, 0.3347541, 0.306112, 0.2786734, 0.2730196, 0.1843636, 
    0.2606786, 0.2640933, 0.274544, 0.2699627, 0.2975982, 0.2630004, 
    0.269563, 0.2519229, 0.2478508, 0.2681874, 0.2517248, 0.242937, 0.272761, 
    0.3168074, 0.2743319, 0.2264045, 0.2878474, 0.2011772, 0.2602438, 
    0.2047939, 0.2272629, 0.2560205,
  0.2810401, 0.2883336, 0.2684129, 0.2681332, 0.2413962, 0.2392218, 
    0.2499226, 0.3111955, 0.2904498, 0.2854399, 0.3179142, 0.2352261, 
    0.2651658, 0.2179268, 0.1982606, 0.2093266, 0.2044178, 0.2093281, 
    0.2429726, 0.1971325, 0.2255282, 0.2568066, 0.2222778, 0.1933275, 
    0.1195101, 0.1934888, 0.2776222, 0.2697371, 0.2898669,
  0.2209542, 0.151854, 0.1194984, 0.1296427, 0.1290615, 0.1767304, 0.1812236, 
    0.2050987, 0.1964413, 0.1696729, 0.13901, 0.1459013, 0.1135143, 
    0.1462392, 0.131464, 0.1751058, 0.1872537, 0.1938332, 0.2014649, 
    0.1974039, 0.2074289, 0.2042722, 0.1728482, 0.2083896, 0.06060553, 
    0.1264553, 0.1805468, 0.2286018, 0.2104347,
  0.07596153, 0.04792123, 0.06780201, 0.05425971, 0.05630739, 0.05122998, 
    0.05426713, 0.0603044, 0.071419, 0.0555601, 0.03030184, 0.01202135, 
    0.0679424, 0.07692777, 0.09325598, 0.1124413, 0.1254499, 0.07403477, 
    0.1576865, 0.128774, 0.08015072, 0.0986965, 0.04479953, 0.007548159, 
    0.05135073, 0.09934625, 0.09911947, 0.1047391, 0.08397456,
  0.002201636, 4.790566e-07, 0.03747486, 0.04800019, 0.06729531, 0.05297393, 
    0.05271097, 0.02087181, 0.04280777, 0.01518383, -3.410193e-06, 
    0.01163191, 0.02071556, 0.09180262, 0.1034353, 0.06208922, 0.02790162, 
    0.02978577, 0.05224635, 0.05838663, 0.06562859, 0.03006706, 0.002506107, 
    2.795534e-05, 0.008263484, 0.05784947, 0.08949146, 0.06726879, 0.02603124,
  8.223254e-08, -9.255044e-07, 0.01061232, 0.1817988, 0.03665683, 0.03826426, 
    0.03830231, 0.08103936, 0.04406205, 0.01402058, 0.06273168, 0.07057161, 
    0.1983397, 0.1012697, 0.0607891, 0.03914943, 0.045901, 0.02764579, 
    0.01691009, 0.008984165, 0.002271884, 9.127417e-07, 1.959684e-07, 
    0.01254059, 0.01775692, 0.001177398, 0.0678071, 0.009885323, 0.001618494,
  0.0001778037, 0.04231615, 0.06687488, 0.01921893, 0.01752127, 0.01532765, 
    0.01465629, 0.01655594, 0.05170574, 0.1393266, 0.04361843, 0.02705611, 
    0.04589138, 0.04047123, 0.03684996, 0.03895803, 0.02131992, 0.010505, 
    0.005244123, 0.0005126905, 0.0005089738, 0.0009936268, 0.01023014, 
    0.1750952, 0.1417357, 0.01739235, 0.01899591, 0.002248333, 0.0008007959,
  0.05005421, 0.04455991, 0.03082817, 0.2969128, 0.003079718, 0.008597583, 
    0.07316324, 0.02914824, 0.01272745, 0.01706847, 0.01219021, 0.03250089, 
    0.05475538, 0.04714379, 0.06182229, 0.09492882, 0.09344168, 0.1445968, 
    0.1466119, 0.1815299, 0.2240038, 0.1034739, 0.1295242, 0.07386309, 
    0.01984342, 0.07609218, 0.1222343, 0.1598519, 0.1514722,
  5.634928e-07, 7.754241e-07, 1.660333e-07, 3.732106e-08, 2.942467e-07, 
    0.0009436717, 0.2629798, 0.2352064, 0.3500805, 0.08192688, 0.1180319, 
    0.09716027, 0.04229885, 0.02408115, 0.02092927, 0.0354804, 0.02532922, 
    0.007737005, 0.01984791, 0.0009414466, 0.0270399, 0.0481187, 0.0117165, 
    0.02213276, 0.03137412, 0.02650765, 0.001031357, 1.892946e-06, 
    3.026363e-05,
  1.012458e-06, 2.023143e-06, -6.445404e-07, 9.355173e-10, 3.488765e-07, 
    3.26448e-06, 0.0367342, 0.2798128, 0.3216757, 0.1003858, 0.06860926, 
    0.04165135, 0.09644212, 0.03754985, 0.04986167, 0.04161388, 0.01685616, 
    0.006078095, 0.0001099019, 2.077311e-07, 0.001052425, 0.01302462, 
    0.06041287, 0.01878316, 0.0170505, 0.03127494, 0.006073354, 0.0009319792, 
    3.661031e-06,
  0.008581762, 0.01207769, 0.01853201, 0.03966215, -0.000154039, 
    -2.404353e-05, 0.01010391, 8.299069e-06, 0.001574757, 0.04549018, 
    0.1210399, 0.07995532, 0.1856487, 0.2105778, 0.1207568, 0.0884669, 
    0.08958033, 0.06158863, 0.01850999, 5.857098e-05, 0.0001837777, 
    0.008161369, 0.07570435, 0.1094022, 0.08714359, 0.05504199, 0.03716974, 
    0.02231167, 0.00179513,
  0.06535001, 0.145098, 0.06388059, 0.09769423, 0.02669728, 0.05359104, 
    0.09125867, 0.18704, 0.1365416, 0.05221158, 0.06490251, 0.1657424, 
    0.103764, 0.1269694, 0.1703001, 0.2080602, 0.2524812, 0.2405108, 
    0.2094112, 0.0843037, 0.05201005, 0.05392995, 0.09943971, 0.1978584, 
    0.1802811, 0.1377024, 0.1202191, 0.1447169, 0.1010654,
  0.1746654, 0.2162021, 0.1510411, 0.1028922, 0.1343566, 0.1094327, 
    0.1822844, 0.1871719, 0.1129361, 0.1753562, 0.1334649, 0.252214, 
    0.2980509, 0.2161442, 0.1361769, 0.3418524, 0.2616258, 0.4286461, 
    0.4144228, 0.1609216, 0.1576036, 0.1789792, 0.1643363, 0.2738979, 
    0.1879025, 0.1959348, 0.182648, 0.2410406, 0.2486227,
  0.2850246, 0.2786775, 0.337065, 0.1889701, 0.1492023, 0.1557429, 0.1795419, 
    0.1740877, 0.1774737, 0.2134689, 0.1615581, 0.2251007, 0.1627139, 
    0.2128453, 0.2514503, 0.1624224, 0.2104797, 0.1107594, 0.1470938, 
    0.1439882, 0.1684705, 0.244947, 0.2433004, 0.2651739, 0.1781897, 
    0.3231692, 0.2133414, 0.2135139, 0.3230153,
  0.1431168, 0.1880053, 0.2475133, 0.210549, 0.1940392, 0.193119, 0.2924473, 
    0.3209511, 0.2352571, 0.2074895, 0.1937383, 0.2414279, 0.2969501, 
    0.2497388, 0.2283069, 0.2304588, 0.2260301, 0.2522336, 0.203929, 
    0.1320567, 0.1351912, 0.2148785, 0.2108691, 0.1284156, 0.1422066, 
    0.1157489, 0.145846, 0.1595654, 0.160779,
  0.2200023, 0.2174552, 0.2149082, 0.2123611, 0.209814, 0.2072669, 0.2047199, 
    0.2206052, 0.219492, 0.2183788, 0.2172656, 0.2161524, 0.2150393, 
    0.2139261, 0.1932014, 0.1985473, 0.2038932, 0.2092392, 0.2145851, 
    0.219931, 0.2252769, 0.2229447, 0.221259, 0.2195733, 0.2178877, 0.216202, 
    0.2145163, 0.2128307, 0.22204,
  0.1361483, 0.1358824, 0.0991874, 0.06118039, 0.0518791, 0.05878922, 
    0.1017567, 0.08767674, 0.04264504, 0.05299811, 0.04509155, 0.03041872, 
    0.06188736, 0.08140144, 0.1133826, 0.1310541, 0.1240633, 0.1494489, 
    0.149521, 0.1875352, 0.282795, 0.395993, 0.319405, 0.2407586, 0.183123, 
    0.1665412, 0.2413736, 0.1983013, 0.174115,
  0.4450694, 0.4605693, 0.4291872, 0.3411198, 0.2058031, 0.07843288, 
    0.1173243, 0.2167333, 0.3014299, 0.2998927, 0.3408679, 0.4079461, 
    0.2920046, 0.3155099, 0.2638069, 0.2087741, 0.1601846, 0.233069, 
    0.2482292, 0.2838477, 0.3521986, 0.2804446, 0.2346744, 0.3382967, 
    0.1757778, 0.1229364, 0.1294496, 0.2209459, 0.335013,
  0.2480936, 0.2546054, 0.4049168, 0.3471807, 0.2773142, 0.2732204, 0.222388, 
    0.2609234, 0.2653038, 0.2901531, 0.3185495, 0.3161147, 0.2817802, 
    0.3374802, 0.3035368, 0.3129593, 0.3171412, 0.2802461, 0.2988417, 
    0.2717939, 0.3160172, 0.2951781, 0.254925, 0.3126926, 0.2101287, 
    0.2886443, 0.2177727, 0.2369501, 0.2593657,
  0.3201681, 0.3249376, 0.3260064, 0.2862928, 0.2659179, 0.2897453, 
    0.2880322, 0.3344182, 0.298537, 0.2939351, 0.308507, 0.2470779, 
    0.2818816, 0.2438441, 0.1971406, 0.2154324, 0.242218, 0.2329847, 
    0.2994041, 0.2789732, 0.2572311, 0.2662188, 0.2771623, 0.2144492, 
    0.1379129, 0.2353058, 0.3428756, 0.3381436, 0.3281738,
  0.2426528, 0.1916769, 0.1391903, 0.1511537, 0.155354, 0.2034175, 0.2009403, 
    0.2419138, 0.2072908, 0.1719946, 0.1492096, 0.1525984, 0.1173866, 
    0.1564798, 0.1507628, 0.1728904, 0.2026739, 0.2142826, 0.2101107, 
    0.2253666, 0.2394668, 0.2229364, 0.2046661, 0.2280332, 0.07589132, 
    0.1689683, 0.2045504, 0.2570219, 0.2248165,
  0.117519, 0.06497107, 0.0577166, 0.09980728, 0.0766675, 0.08084688, 
    0.07597318, 0.09740163, 0.1028003, 0.09394926, 0.01931045, 0.004180716, 
    0.06403866, 0.09527646, 0.1072745, 0.1226728, 0.137849, 0.1151838, 
    0.2043776, 0.1413074, 0.09590931, 0.1207813, 0.0936314, 0.009570894, 
    0.04316113, 0.115306, 0.145805, 0.1265836, 0.1252159,
  0.04094796, -2.861696e-05, 0.01404254, 0.06530008, 0.06367747, 0.07971612, 
    0.09006311, 0.06594113, 0.08718166, 0.03454743, -5.374884e-08, 
    0.007367549, 0.0415243, 0.106128, 0.1374959, 0.06606936, 0.04845629, 
    0.03778666, 0.05356605, 0.07383355, 0.1412593, 0.1163252, 0.03820416, 
    8.590376e-06, 0.006486698, 0.06434304, 0.09329841, 0.1837622, 0.09236676,
  5.974427e-07, 2.664685e-07, 0.003358303, 0.1723465, 0.03032792, 0.04131643, 
    0.06399574, 0.08860271, 0.04558183, 0.02733762, 0.08532497, 0.08062525, 
    0.2295974, 0.08646619, 0.05663361, 0.03496566, 0.03928812, 0.02077655, 
    0.01884919, 0.01341859, 0.006388585, 0.0001667545, 1.488743e-07, 
    0.01847003, 0.001178255, -1.795669e-06, 0.06045831, 0.02355921, 
    0.005777002,
  0.0006436871, 0.05282976, 0.04461303, 0.01658661, 0.02512563, 0.02077981, 
    0.01532305, 0.0168702, 0.04803647, 0.1343091, 0.04631166, 0.02402665, 
    0.0374408, 0.03611765, 0.03357357, 0.03096696, 0.02329895, 0.01556494, 
    0.009672575, 0.007261843, 0.001531086, 0.003794906, 0.005591261, 
    0.1627984, 0.1458402, 0.01398581, 0.02056011, 0.01258275, 0.0006810178,
  0.0526192, 0.04448458, 0.02969134, 0.243728, 0.0004601396, 0.01232923, 
    0.06046097, 0.02690968, 0.01162067, 0.01449557, 0.01393408, 0.03146045, 
    0.04268904, 0.04004864, 0.0550659, 0.08912854, 0.09615098, 0.14647, 
    0.1253883, 0.1573143, 0.1979266, 0.09393314, 0.1268055, 0.07821134, 
    0.01941134, 0.06946959, 0.1252637, 0.1528976, 0.1424675,
  -1.146562e-08, 3.257101e-07, 7.291906e-08, 1.308975e-08, 2.082374e-07, 
    0.002957597, 0.2641772, 0.2109077, 0.3197052, 0.0718088, 0.08904609, 
    0.08650474, 0.03628685, 0.02299003, 0.02225287, 0.04853585, 0.03267031, 
    0.03448134, 0.02562045, 0.00364538, 0.02433127, 0.05190875, 0.01165714, 
    0.02161087, 0.04238063, 0.04337413, 0.01000809, 3.178476e-07, 1.58858e-05,
  6.209392e-07, 1.528457e-06, 3.120545e-10, 5.246574e-10, 2.251527e-07, 
    -8.588728e-07, 0.02746721, 0.2584466, 0.3026722, 0.107021, 0.06502439, 
    0.04687399, 0.08828653, 0.03015224, 0.04388517, 0.05588782, 0.03358565, 
    0.0262547, 0.001539281, 1.231138e-07, 0.0004487558, 0.01359577, 
    0.05627881, 0.01718187, 0.01830015, 0.0428323, 0.03912527, 0.003421021, 
    3.261839e-06,
  0.005038122, 0.01104766, 0.01285312, 0.0595971, -0.0001183224, -3.1215e-06, 
    0.006607024, 5.311961e-06, -2.146802e-05, 0.04559596, 0.1619549, 
    0.07768305, 0.1964911, 0.2258766, 0.1248512, 0.1045527, 0.1249443, 
    0.1142325, 0.03087251, 5.897457e-06, 7.101724e-05, 0.006373082, 
    0.08248637, 0.1049535, 0.08338445, 0.06077177, 0.05814456, 0.03665127, 
    0.0006273148,
  0.1112742, 0.1703602, 0.09342459, 0.08625028, 0.00929754, 0.05080474, 
    0.05962829, 0.1932016, 0.1140649, 0.03721291, 0.06674001, 0.1862459, 
    0.1253488, 0.149299, 0.2086959, 0.2236061, 0.271674, 0.286922, 0.2599514, 
    0.08234902, 0.05031588, 0.07078214, 0.101321, 0.196227, 0.1726917, 
    0.12084, 0.155354, 0.1644443, 0.1461249,
  0.1918991, 0.2252394, 0.1631104, 0.126878, 0.1398931, 0.1004439, 0.2009811, 
    0.1887364, 0.1305808, 0.1762022, 0.1498655, 0.2541828, 0.3280105, 
    0.2393447, 0.1438493, 0.3223796, 0.2770315, 0.4337944, 0.4195739, 
    0.1540753, 0.1268232, 0.1879284, 0.1643708, 0.2942629, 0.1726692, 
    0.2086171, 0.2299597, 0.2771462, 0.2723507,
  0.3168791, 0.2884042, 0.329784, 0.2016705, 0.2010518, 0.1938169, 0.2028406, 
    0.1947602, 0.1785076, 0.2244393, 0.1624352, 0.2572568, 0.2217295, 
    0.2560951, 0.2711343, 0.1467631, 0.2088324, 0.1271126, 0.1601669, 
    0.1348108, 0.2081564, 0.2646042, 0.3119467, 0.2862916, 0.1700602, 
    0.3287901, 0.2327296, 0.2216547, 0.3257309,
  0.1735309, 0.2492625, 0.2830357, 0.2023301, 0.194484, 0.2288882, 0.3060858, 
    0.3245039, 0.3251057, 0.2702268, 0.2854285, 0.2996497, 0.3016313, 
    0.2283684, 0.2223077, 0.2489515, 0.2635432, 0.2837717, 0.2021448, 
    0.1773786, 0.1741433, 0.2219476, 0.2255868, 0.1427815, 0.1196929, 
    0.1561931, 0.1522163, 0.1810038, 0.1948061,
  0.2480035, 0.2453096, 0.2426156, 0.2399217, 0.2372278, 0.2345339, 0.23184, 
    0.2483516, 0.2464218, 0.2444919, 0.242562, 0.2406321, 0.2387023, 
    0.2367724, 0.2368877, 0.2429965, 0.2491054, 0.2552142, 0.2613231, 
    0.2674319, 0.2735408, 0.2622818, 0.2607968, 0.2593117, 0.2578267, 
    0.2563416, 0.2548565, 0.2533714, 0.2501586,
  0.1319932, 0.1417026, 0.1289532, 0.07698086, 0.06295826, 0.08555952, 
    0.1225173, 0.1035956, 0.04841653, 0.06650253, 0.05414107, 0.03324959, 
    0.07610444, 0.08135734, 0.1220788, 0.1198303, 0.120563, 0.1297277, 
    0.1346812, 0.1784727, 0.326004, 0.4121389, 0.3498947, 0.2322852, 
    0.2001414, 0.1803336, 0.2204499, 0.1828417, 0.1759037,
  0.4573802, 0.4366724, 0.442601, 0.3145882, 0.1908889, 0.08021621, 
    0.1126892, 0.2390303, 0.3193218, 0.3067155, 0.3616956, 0.4014786, 
    0.2801008, 0.3001378, 0.3005683, 0.2304933, 0.1903944, 0.2670886, 
    0.3045318, 0.3043165, 0.3479356, 0.2917446, 0.2450874, 0.3771789, 
    0.1625304, 0.1240551, 0.1307864, 0.2643111, 0.3485411,
  0.2806582, 0.307715, 0.4847779, 0.3623514, 0.3388978, 0.3678179, 0.2352277, 
    0.3013233, 0.3049574, 0.3184246, 0.3722305, 0.3116737, 0.3312271, 
    0.3798304, 0.3632808, 0.3681679, 0.3671173, 0.3874443, 0.3857874, 
    0.3428175, 0.3428211, 0.3029256, 0.3064808, 0.3695289, 0.3075823, 
    0.3428313, 0.259497, 0.2654782, 0.2587873,
  0.3721621, 0.3698602, 0.3484832, 0.3368813, 0.3139611, 0.2863989, 
    0.3026311, 0.3457372, 0.2777063, 0.2745222, 0.2717196, 0.2616927, 
    0.2804356, 0.2604948, 0.2396883, 0.2215758, 0.2690126, 0.2673599, 
    0.3179292, 0.3196791, 0.2890845, 0.3181155, 0.3001217, 0.2295921, 
    0.1621109, 0.2762666, 0.4099344, 0.380772, 0.3655232,
  0.2751526, 0.2223385, 0.1540222, 0.2243668, 0.2293402, 0.2430908, 
    0.2148878, 0.2356664, 0.1948004, 0.1542973, 0.1580364, 0.1459617, 
    0.1179156, 0.1454011, 0.1909739, 0.1633291, 0.2041444, 0.2320065, 
    0.2217664, 0.2286178, 0.2567473, 0.2531731, 0.2411144, 0.2637202, 
    0.1165094, 0.1846845, 0.2200544, 0.2392399, 0.2036643,
  0.1549382, 0.07995334, 0.04500671, 0.1265509, 0.1644, 0.150737, 0.1766514, 
    0.2307834, 0.2100413, 0.1444576, 0.002225414, 0.0009058882, 0.05674983, 
    0.09936617, 0.1183046, 0.1324358, 0.1269859, 0.1239602, 0.1789277, 
    0.1298121, 0.1439169, 0.1474628, 0.1788072, 0.01325541, 0.05521471, 
    0.1014623, 0.1150109, 0.1799074, 0.18885,
  0.1834824, -0.0001212308, 0.006924577, 0.1056692, 0.07262345, 0.105992, 
    0.1235308, 0.1722274, 0.2853104, 0.06198003, -2.053999e-09, 0.000791789, 
    0.1282046, 0.1798341, 0.1291955, 0.07551177, 0.07239744, 0.04222762, 
    0.05420442, 0.0958042, 0.2060112, 0.2712655, 0.1372874, 5.765608e-06, 
    0.01236443, 0.04101852, 0.08246246, 0.3024696, 0.3681349,
  0.001758546, 3.786357e-06, 0.0001740079, 0.09130018, 0.03215731, 
    0.04330386, 0.08202766, 0.08990161, 0.05104644, 0.0448469, 0.09723236, 
    0.09111333, 0.2435623, 0.0694979, 0.05169388, 0.03411512, 0.03740058, 
    0.02312164, 0.02260509, 0.02643815, 0.03101462, 0.01729257, 1.116223e-06, 
    0.01819322, 0.0001709799, -2.142166e-06, 0.071618, 0.030942, 0.03614933,
  0.009374806, 0.1118436, 0.03227926, 0.01447768, 0.03001728, 0.03096389, 
    0.02211318, 0.02088139, 0.04459481, 0.1349536, 0.04519192, 0.02304944, 
    0.03415617, 0.03308747, 0.03120793, 0.02754798, 0.01841654, 0.01573447, 
    0.01746567, 0.01916976, 0.00811062, 0.0007599076, 0.002883772, 0.1697322, 
    0.1440946, 0.0141606, 0.0261117, 0.02345211, 0.008285496,
  0.06282876, 0.04635542, 0.02501969, 0.2195579, -0.0003040804, 0.01683498, 
    0.05225125, 0.02635596, 0.01095987, 0.01598727, 0.0209746, 0.03133594, 
    0.03552834, 0.03655295, 0.05116913, 0.08111189, 0.09007207, 0.133196, 
    0.1074587, 0.1255038, 0.1665592, 0.07928817, 0.127315, 0.07508597, 
    0.02130149, 0.06346369, 0.121344, 0.1438953, 0.1353097,
  1.49029e-07, 1.893722e-07, 4.331628e-08, 7.780158e-09, 1.317578e-07, 
    0.01411346, 0.247795, 0.1816499, 0.2911935, 0.05538383, 0.0679087, 
    0.07186514, 0.03611146, 0.02640367, 0.02665997, 0.05068984, 0.08073113, 
    0.0683435, 0.03653314, 0.004935314, 0.02164622, 0.05760169, 0.01364643, 
    0.02236969, 0.05059688, 0.06119706, 0.04337643, 6.720675e-06, 5.25514e-06,
  4.632299e-07, 1.240939e-06, 2.404784e-07, 3.586123e-10, 1.630935e-07, 
    -8.58922e-07, 0.0160396, 0.2444818, 0.3054828, 0.09195215, 0.05861946, 
    0.05441047, 0.07363233, 0.02818857, 0.04489903, 0.06004554, 0.07191312, 
    0.05758093, 0.00331832, 9.40002e-08, 0.0001646569, 0.01560373, 
    0.05159745, 0.01911375, 0.02673916, 0.04731944, 0.1014803, 0.01305284, 
    4.188867e-06,
  0.001532382, 0.008061524, 0.01038835, 0.07911218, -2.709314e-05, 
    -1.257737e-06, 0.005948571, 1.672457e-06, -0.0001012302, 0.0382972, 
    0.1927395, 0.07328719, 0.2038582, 0.2356544, 0.1342149, 0.1344763, 
    0.1824868, 0.1589038, 0.07616303, 4.145872e-06, -2.734425e-05, 
    0.005466288, 0.09322046, 0.1083713, 0.0852599, 0.07893573, 0.08201934, 
    0.05278436, 0.007245413,
  0.1295117, 0.1651599, 0.08373891, 0.07881834, 0.006071336, 0.04269985, 
    0.04165691, 0.1797851, 0.09451558, 0.02767228, 0.06143462, 0.2175096, 
    0.1357346, 0.1953871, 0.2195303, 0.2566887, 0.3143288, 0.3349174, 
    0.2663375, 0.08154568, 0.03316266, 0.05709283, 0.09035466, 0.2017438, 
    0.1683476, 0.137303, 0.2224665, 0.2122285, 0.1822537,
  0.2236781, 0.223521, 0.1320778, 0.1170962, 0.1511703, 0.1114695, 0.2154061, 
    0.2097185, 0.1273748, 0.164886, 0.2077016, 0.2722505, 0.3538696, 
    0.2644596, 0.1649849, 0.3221739, 0.3075579, 0.4334857, 0.3855011, 
    0.1313246, 0.09240901, 0.173589, 0.1658695, 0.2932335, 0.1648831, 
    0.2169489, 0.2973095, 0.3704379, 0.3012195,
  0.3508092, 0.2951856, 0.3273929, 0.2135321, 0.2477088, 0.2613977, 
    0.2415803, 0.2137581, 0.202552, 0.2464868, 0.2151331, 0.2580804, 
    0.2535307, 0.2592608, 0.2409806, 0.1408588, 0.2227325, 0.1198487, 
    0.1531659, 0.1503581, 0.3139414, 0.2950206, 0.3602478, 0.3428745, 
    0.1620335, 0.3545245, 0.2378873, 0.238598, 0.3257995,
  0.2898725, 0.3549261, 0.3544366, 0.2661237, 0.2489759, 0.3081865, 0.37641, 
    0.3454144, 0.3704698, 0.290203, 0.3266203, 0.3284135, 0.3561413, 
    0.2750911, 0.2924967, 0.2940955, 0.333723, 0.3160036, 0.2131589, 
    0.2439869, 0.2243603, 0.2730358, 0.2655303, 0.1559322, 0.1272206, 
    0.1799031, 0.1688632, 0.1945408, 0.2780401,
  0.2990524, 0.29626, 0.2934675, 0.2906751, 0.2878826, 0.2850902, 0.2822978, 
    0.2814484, 0.2795157, 0.2775829, 0.2756501, 0.2737174, 0.2717847, 
    0.2698519, 0.2796295, 0.2857853, 0.2919412, 0.298097, 0.3042528, 
    0.3104086, 0.3165644, 0.3052091, 0.3037785, 0.3023479, 0.3009172, 
    0.2994866, 0.298056, 0.2966253, 0.3012864,
  0.128814, 0.1366836, 0.1460875, 0.1023117, 0.06398845, 0.09951207, 
    0.1302954, 0.1172436, 0.05695257, 0.07128917, 0.06652829, 0.03744005, 
    0.08641591, 0.07697485, 0.1234366, 0.1148938, 0.1114689, 0.1067912, 
    0.1344837, 0.1759295, 0.3642404, 0.4123657, 0.3634216, 0.2339002, 
    0.2147853, 0.1886351, 0.2206669, 0.1579697, 0.1624776,
  0.4381544, 0.4004653, 0.4456585, 0.2698456, 0.1698981, 0.09269037, 
    0.07713735, 0.2587799, 0.3355503, 0.3182198, 0.3691355, 0.3897875, 
    0.2518701, 0.2898028, 0.3150306, 0.250708, 0.2063182, 0.3024563, 
    0.3490166, 0.3604522, 0.3711888, 0.3034765, 0.2391339, 0.4176876, 
    0.1553185, 0.1307232, 0.1755782, 0.2656425, 0.3505643,
  0.3007684, 0.3814976, 0.4675092, 0.3253703, 0.3410075, 0.4239649, 
    0.2340333, 0.385433, 0.3533728, 0.3215546, 0.3795456, 0.3222513, 
    0.3633656, 0.3865162, 0.3233603, 0.3278841, 0.4071241, 0.3800329, 
    0.3508561, 0.3052142, 0.311662, 0.2783241, 0.2959276, 0.3621712, 
    0.3683035, 0.3450582, 0.2782001, 0.2847446, 0.2977111,
  0.3650855, 0.3839943, 0.3916283, 0.3932093, 0.3490472, 0.2866026, 0.305476, 
    0.2594607, 0.2464204, 0.2569778, 0.2548028, 0.2441587, 0.2882738, 
    0.2506891, 0.2788855, 0.2413616, 0.2357028, 0.2826865, 0.322978, 
    0.3244951, 0.2725137, 0.2823632, 0.2728397, 0.2609364, 0.167904, 
    0.3034722, 0.4088185, 0.3666161, 0.3575347,
  0.2657953, 0.2142392, 0.1351397, 0.2046992, 0.2458706, 0.2075807, 
    0.2037177, 0.2079448, 0.1696162, 0.1442924, 0.1390738, 0.1125748, 
    0.1118117, 0.1244869, 0.3068309, 0.1591023, 0.1912955, 0.2135738, 
    0.1925398, 0.1980147, 0.2352295, 0.2680511, 0.2221415, 0.3120869, 
    0.0900818, 0.1559357, 0.1610231, 0.1881634, 0.1760109,
  0.2025454, 0.07191452, 0.04237618, 0.1143545, 0.1445524, 0.1412946, 
    0.2509322, 0.2290304, 0.1990281, 0.0986921, 0.0004826146, 0.001059917, 
    0.0475692, 0.04532928, 0.08897625, 0.1137259, 0.1126201, 0.104807, 
    0.1613434, 0.1163647, 0.1430127, 0.1615156, 0.2134964, 0.01484301, 
    0.04623879, 0.09888674, 0.1077159, 0.1112988, 0.1590806,
  0.3356512, -0.0006733458, 0.00521534, 0.1235271, 0.08267, 0.09926496, 
    0.1313389, 0.1731391, 0.2790484, 0.02187549, 2.930266e-10, 9.23953e-05, 
    0.09789038, 0.1959748, 0.1408578, 0.09742512, 0.1209634, 0.05385378, 
    0.0709483, 0.1156159, 0.1660543, 0.345036, 0.3228491, -1.354445e-05, 
    0.01767446, 0.03458212, 0.06010893, 0.1967987, 0.3521232,
  0.02244054, 7.20058e-05, -0.0001996393, 0.05585833, 0.04638099, 0.05902695, 
    0.08081968, 0.08622503, 0.07219326, 0.08062667, 0.1289986, 0.1185379, 
    0.2328534, 0.062085, 0.05821099, 0.04216019, 0.04402879, 0.05173194, 
    0.05402102, 0.07028669, 0.1125001, 0.1190449, 2.382522e-05, 0.02291655, 
    3.2549e-05, -6.032402e-07, 0.09925277, 0.05306397, 0.1717401,
  0.05528092, 0.1587959, 0.02377117, 0.01332917, 0.0404736, 0.09047631, 
    0.06045077, 0.03741226, 0.03435454, 0.1233987, 0.04683531, 0.02535515, 
    0.03386601, 0.03798627, 0.03190625, 0.03032953, 0.02301194, 0.01564942, 
    0.01599939, 0.01824654, 0.03293806, 0.006978329, 0.002132414, 0.1992338, 
    0.1147204, 0.01821626, 0.05429486, 0.03891428, 0.04586221,
  0.06980044, 0.04497807, 0.0177072, 0.2076596, -0.0003190448, 0.01842895, 
    0.04608715, 0.03090778, 0.008846534, 0.01989419, 0.01454446, 0.03926718, 
    0.03311862, 0.03343353, 0.04946538, 0.08019844, 0.0846438, 0.1224477, 
    0.09910794, 0.1126814, 0.1416406, 0.06862541, 0.1203832, 0.06109073, 
    0.02784833, 0.06204124, 0.1126437, 0.1324388, 0.1253121,
  1.845385e-07, 1.315801e-07, 3.129545e-08, 5.613674e-09, 8.975594e-08, 
    0.02290881, 0.1909763, 0.1548566, 0.2607331, 0.03931957, 0.06196258, 
    0.06406737, 0.04220758, 0.03635706, 0.0366814, 0.05825341, 0.1271437, 
    0.1426817, 0.05585869, 0.01415012, 0.01429318, 0.0601059, 0.02045424, 
    0.02384637, 0.05428575, 0.08037392, 0.0909351, 0.0002238135, 2.164591e-07,
  3.884253e-07, 1.05413e-06, -8.381261e-08, 1.491508e-10, 1.274445e-07, 
    -4.600335e-07, 0.00753919, 0.2566019, 0.3056441, 0.07795168, 0.05650223, 
    0.07866906, 0.08192651, 0.02948622, 0.05194253, 0.07065006, 0.1194109, 
    0.1516648, 0.03847323, 1.281389e-07, 4.968177e-05, 0.01410429, 0.0459561, 
    0.02383738, 0.03243113, 0.06133877, 0.1541428, 0.05875655, -1.514122e-05,
  0.0004186877, 0.00432709, 0.008993896, 0.1117531, -8.000301e-05, 
    -5.453735e-07, 0.006020422, 1.474793e-06, -8.338953e-05, 0.03328433, 
    0.2122191, 0.07385652, 0.2101972, 0.2575714, 0.1893831, 0.2133804, 
    0.2825352, 0.2716224, 0.1816316, 2.277513e-06, -0.000154332, 0.002566915, 
    0.08519285, 0.100965, 0.09825139, 0.1418485, 0.1486787, 0.1360127, 
    0.02040746,
  0.1131836, 0.1342551, 0.06282526, 0.06686619, 0.005128035, 0.03608171, 
    0.0294539, 0.1569481, 0.08106636, 0.02022288, 0.05196245, 0.2188413, 
    0.1666633, 0.2277843, 0.2595818, 0.330388, 0.3840909, 0.450089, 
    0.3353391, 0.06575692, 0.02972075, 0.0488212, 0.08587657, 0.196261, 
    0.148762, 0.1633492, 0.3191898, 0.302247, 0.2198281,
  0.246083, 0.1809551, 0.131615, 0.09364434, 0.1173506, 0.07645237, 
    0.1973866, 0.200706, 0.1234371, 0.1377412, 0.1798997, 0.2749285, 
    0.3731932, 0.2834981, 0.1777738, 0.3510196, 0.2996557, 0.4190291, 
    0.349678, 0.08786687, 0.06664626, 0.1477881, 0.1721656, 0.2894602, 
    0.155362, 0.2094789, 0.3251648, 0.4070264, 0.3452378,
  0.4673334, 0.3459158, 0.3347064, 0.2419702, 0.2474617, 0.2651884, 
    0.2797296, 0.2588037, 0.2146674, 0.2954111, 0.2629506, 0.3499404, 
    0.2667273, 0.2639666, 0.2530478, 0.163533, 0.2473372, 0.1115454, 
    0.1342628, 0.1635102, 0.3382458, 0.3204725, 0.4068001, 0.3862343, 
    0.1601039, 0.3798568, 0.2628262, 0.248363, 0.3911759,
  0.3919265, 0.4486506, 0.4308593, 0.3569453, 0.3676963, 0.4035715, 
    0.4546183, 0.4145067, 0.4016619, 0.3456663, 0.361374, 0.4126334, 
    0.4257304, 0.3593792, 0.3581195, 0.3511496, 0.3741742, 0.3590303, 
    0.2715166, 0.2519239, 0.2858847, 0.2862189, 0.3113441, 0.2090545, 
    0.1387921, 0.2375669, 0.1631761, 0.2419702, 0.3394162,
  0.3303313, 0.328487, 0.3266427, 0.3247984, 0.3229541, 0.3211098, 0.3192654, 
    0.3159894, 0.3132561, 0.3105229, 0.3077897, 0.3050565, 0.3023232, 
    0.29959, 0.3230369, 0.3288611, 0.3346853, 0.3405095, 0.3463337, 
    0.3521579, 0.357982, 0.3317607, 0.330514, 0.3292674, 0.3280208, 
    0.3267741, 0.3255274, 0.3242808, 0.3318067,
  0.1298932, 0.1429329, 0.14397, 0.1182183, 0.07219249, 0.1078623, 0.138475, 
    0.1281251, 0.05868615, 0.07240775, 0.08651464, 0.0480414, 0.0932686, 
    0.06833944, 0.1136942, 0.1143244, 0.09659366, 0.08088047, 0.1374398, 
    0.1710274, 0.3835666, 0.4192846, 0.3686329, 0.225487, 0.2119749, 
    0.1925192, 0.2140467, 0.13853, 0.1543345,
  0.4042727, 0.3690485, 0.4476623, 0.1958687, 0.1404483, 0.1041497, 
    0.03983469, 0.2856571, 0.3565345, 0.3224506, 0.3803119, 0.357901, 
    0.2288087, 0.2756146, 0.3099086, 0.2793379, 0.2404375, 0.3539014, 
    0.3945739, 0.3561625, 0.3853871, 0.2773008, 0.2570168, 0.4313501, 
    0.1581822, 0.1911179, 0.1967503, 0.2752262, 0.3706209,
  0.3157773, 0.3792396, 0.4271565, 0.313576, 0.3234829, 0.4159324, 0.2874767, 
    0.4388279, 0.3779642, 0.2678013, 0.328085, 0.3312155, 0.3500624, 
    0.3573849, 0.3249108, 0.2878349, 0.3784876, 0.372144, 0.3335148, 
    0.2534693, 0.2556818, 0.2780762, 0.248695, 0.3452948, 0.3531769, 
    0.3627951, 0.3400635, 0.3277621, 0.3713313,
  0.3538003, 0.3839874, 0.4118967, 0.425156, 0.3759955, 0.3219606, 0.2938293, 
    0.1893474, 0.2179421, 0.2421716, 0.2511176, 0.2243796, 0.2618343, 
    0.2167456, 0.2483004, 0.1899495, 0.2042065, 0.258204, 0.2948023, 
    0.2997984, 0.2563522, 0.2759432, 0.2633618, 0.267574, 0.1948218, 
    0.2798858, 0.3658201, 0.3585834, 0.3470055,
  0.240111, 0.1955799, 0.1081264, 0.180585, 0.2018844, 0.1635518, 0.168438, 
    0.1904567, 0.1764826, 0.1344052, 0.1058897, 0.09198725, 0.05568459, 
    0.09738611, 0.3685643, 0.1331712, 0.1511796, 0.1848911, 0.1508167, 
    0.1960821, 0.1874462, 0.2735308, 0.2301986, 0.3541237, 0.05758172, 
    0.1377057, 0.1311026, 0.1633755, 0.1603708,
  0.180911, 0.04709765, 0.04397979, 0.06467257, 0.1145624, 0.102815, 
    0.1467151, 0.1408522, 0.1066625, 0.03208171, 4.785576e-05, 0.0007557899, 
    0.03466875, 0.01969474, 0.04882681, 0.07370807, 0.1009834, 0.09267581, 
    0.1258256, 0.106558, 0.09384114, 0.1210208, 0.2235365, 0.02437232, 
    0.06109559, 0.08176452, 0.09241234, 0.07274354, 0.09585278,
  0.2799423, 0.003465135, 0.003122678, 0.1075065, 0.05382061, 0.05986005, 
    0.08953983, 0.1421803, 0.1661368, 0.01619918, 2.161726e-10, 4.398618e-06, 
    0.0429407, 0.1881237, 0.153664, 0.1249175, 0.1117457, 0.0954005, 
    0.09510343, 0.06656502, 0.1303088, 0.2486028, 0.3989193, -0.0006506945, 
    0.0224626, 0.05347142, 0.03913091, 0.1103123, 0.1908982,
  0.3903741, 0.001727947, 0.000139535, 0.04430107, 0.03943755, 0.06081246, 
    0.09676085, 0.1088397, 0.06912999, 0.06543414, 0.08203006, 0.07479821, 
    0.20252, 0.07340124, 0.05563363, 0.05290673, 0.03903271, 0.04339479, 
    0.03281186, 0.05630852, 0.1372443, 0.3763618, 0.06053919, 0.01190395, 
    5.77701e-06, -9.68555e-07, 0.0465463, 0.03801014, 0.268987,
  0.2042725, 0.1768841, 0.008842833, 0.01667968, 0.04549916, 0.08037899, 
    0.1326554, 0.09596254, 0.02819687, 0.1033666, 0.07421376, 0.05442507, 
    0.08516588, 0.04390862, 0.07334856, 0.04288217, 0.03466006, 0.03286178, 
    0.043187, 0.03268744, 0.04427731, 0.04493652, 0.009553879, 0.1478869, 
    0.06803402, 0.04253536, 0.06293134, 0.07864456, 0.09433831,
  0.07550399, 0.03984339, 0.008673705, 0.2006498, -0.0001689017, 0.01891592, 
    0.04256182, 0.03555973, 0.006260123, 0.03979312, 0.009772265, 0.08611964, 
    0.04232204, 0.03805052, 0.05121926, 0.07865441, 0.0957511, 0.135687, 
    0.1233127, 0.1073272, 0.1334924, 0.07250197, 0.1090357, 0.05629463, 
    0.04267328, 0.07525944, 0.1020159, 0.1386259, 0.1015504,
  1.74074e-07, 3.99669e-08, 2.648639e-08, 3.858803e-09, 6.613442e-08, 
    0.04387481, 0.1866678, 0.1235321, 0.230692, 0.0321083, 0.05682389, 
    0.05975784, 0.04252587, 0.03905725, 0.03893607, 0.05205327, 0.09037937, 
    0.2124541, 0.1950289, 0.05414189, 0.01793888, 0.07459007, 0.05511937, 
    0.02116856, 0.05022401, 0.1076801, 0.2284359, 0.004889977, -4.002129e-07,
  3.473673e-07, 6.752291e-07, -3.499278e-06, -1.005732e-09, 1.080489e-07, 
    -2.328355e-07, 0.003549438, 0.2684144, 0.3056018, 0.05943621, 0.06625055, 
    0.0692932, 0.08980162, 0.0493562, 0.08140551, 0.07283431, 0.1472436, 
    0.2053792, 0.2136556, 1.035055e-05, 3.141613e-05, 0.009673459, 
    0.03414499, 0.03341398, 0.04817498, 0.08582067, 0.156293, 0.318518, 
    -0.000187546,
  -9.057151e-05, 0.003532479, 0.005982351, 0.147508, -8.923929e-05, 
    -2.257556e-07, 0.004834141, 1.287496e-06, -6.637353e-05, 0.03128745, 
    0.2127974, 0.0687187, 0.2518903, 0.2938572, 0.2679727, 0.3526095, 
    0.4064187, 0.3692768, 0.320895, 3.047736e-05, -0.0001218822, 0.001179832, 
    0.07896867, 0.1073402, 0.1036611, 0.1817893, 0.2027114, 0.3147454, 
    0.03909161,
  0.129237, 0.1247124, 0.05460976, 0.06411415, 0.005167633, 0.03333761, 
    0.02230939, 0.1566928, 0.07875241, 0.01772014, 0.04513996, 0.204709, 
    0.2291196, 0.3163282, 0.3553259, 0.4268543, 0.4788933, 0.4872038, 
    0.415168, 0.06430227, 0.02762663, 0.03175376, 0.07341002, 0.1649, 
    0.1443859, 0.2084183, 0.3738689, 0.4183396, 0.2790568,
  0.2437773, 0.1411031, 0.1028448, 0.07672108, 0.08414152, 0.04319092, 
    0.1476293, 0.1730874, 0.1115374, 0.1182452, 0.1425512, 0.2774352, 
    0.3743588, 0.295041, 0.2022168, 0.4374724, 0.2775891, 0.3976317, 
    0.3278239, 0.07045604, 0.06294005, 0.1257057, 0.1685701, 0.2673509, 
    0.1597993, 0.2083171, 0.3579996, 0.4546017, 0.368767,
  0.5177895, 0.3893334, 0.3376455, 0.2576051, 0.2761158, 0.2748682, 
    0.2997026, 0.2518767, 0.189318, 0.2836639, 0.2760814, 0.3711516, 
    0.2768608, 0.2910434, 0.2955977, 0.2512304, 0.314817, 0.135262, 
    0.1435095, 0.2158587, 0.3654128, 0.393455, 0.3602892, 0.3927703, 
    0.1733858, 0.3921253, 0.2790987, 0.2852077, 0.4706216,
  0.4477584, 0.4451504, 0.4630896, 0.4235719, 0.4704698, 0.5322536, 
    0.5515447, 0.5155509, 0.5217398, 0.4542019, 0.4333994, 0.5095899, 
    0.479593, 0.4458626, 0.4103152, 0.3746077, 0.3443248, 0.3631327, 
    0.3428982, 0.3805202, 0.4021837, 0.3331903, 0.3196624, 0.2692237, 
    0.1709523, 0.1940567, 0.2065699, 0.2948377, 0.4369916,
  0.3844549, 0.3842859, 0.3841168, 0.3839478, 0.3837788, 0.3836097, 
    0.3834406, 0.3774076, 0.3734662, 0.3695248, 0.3655834, 0.361642, 
    0.3577006, 0.3537592, 0.3564287, 0.3615147, 0.3666008, 0.3716869, 
    0.376773, 0.3818591, 0.3869452, 0.3577188, 0.3567432, 0.3557675, 
    0.3547919, 0.3538163, 0.3528407, 0.3518651, 0.3845902,
  0.1314287, 0.1479151, 0.1563504, 0.1359298, 0.09767906, 0.1154573, 
    0.1447812, 0.1265714, 0.05303013, 0.08163414, 0.1131244, 0.08293895, 
    0.107858, 0.05465036, 0.1236491, 0.1102961, 0.0956668, 0.07493643, 
    0.1347595, 0.1703494, 0.384513, 0.4409388, 0.3678502, 0.2196871, 
    0.1995842, 0.2118883, 0.1882909, 0.1163023, 0.1493256,
  0.3855619, 0.3423081, 0.4287825, 0.1318285, 0.1111672, 0.09967534, 
    0.02084741, 0.2937335, 0.3590184, 0.3257527, 0.3851429, 0.3416604, 
    0.2024216, 0.2506301, 0.3154421, 0.3135829, 0.287784, 0.4054781, 
    0.4459196, 0.3805624, 0.4069229, 0.2770838, 0.2784936, 0.4462643, 
    0.1587823, 0.2036138, 0.2323155, 0.2806042, 0.3933366,
  0.3607446, 0.3889992, 0.3821995, 0.3016835, 0.2798704, 0.3567311, 
    0.2807192, 0.435186, 0.3052717, 0.2077122, 0.2910679, 0.3300335, 
    0.3211934, 0.3411379, 0.3238076, 0.2887237, 0.3310826, 0.3948904, 
    0.296327, 0.2185889, 0.2446512, 0.2468244, 0.2171169, 0.3504929, 
    0.2893221, 0.3789321, 0.3742233, 0.3914893, 0.411488,
  0.3427613, 0.4086635, 0.4105162, 0.4261786, 0.4097388, 0.341754, 0.2649323, 
    0.1506198, 0.2032458, 0.2375516, 0.2655806, 0.2243408, 0.2152388, 
    0.1689695, 0.2007187, 0.1536041, 0.1573466, 0.1854326, 0.2462174, 
    0.2564612, 0.2261872, 0.2630531, 0.2668149, 0.2685728, 0.1617818, 
    0.2600661, 0.3478985, 0.3280757, 0.335224,
  0.2037465, 0.1174248, 0.07084827, 0.1435243, 0.1263901, 0.1266596, 
    0.1246304, 0.1619184, 0.1554216, 0.1045443, 0.07572746, 0.05879012, 
    0.02855275, 0.06421704, 0.3551369, 0.09702075, 0.1301893, 0.1595106, 
    0.132379, 0.1810117, 0.1766919, 0.2294488, 0.218717, 0.3790702, 
    0.04595088, 0.1146246, 0.1262785, 0.1676086, 0.1658879,
  0.1034585, 0.03228311, 0.03901932, 0.03708466, 0.05374134, 0.04467947, 
    0.06230852, 0.07199432, 0.06518468, 0.008306112, -1.245211e-05, 
    0.0001129805, 0.02404733, 0.009805739, 0.02870136, 0.05670752, 
    0.09107904, 0.07446223, 0.1207663, 0.07894548, 0.05051871, 0.08432537, 
    0.1334588, 0.02536957, 0.04768826, 0.07061005, 0.04988315, 0.04645061, 
    0.05130052,
  0.1334929, 0.01765558, 0.0008066995, 0.03451177, 0.01339034, 0.01935798, 
    0.0332323, 0.08228604, 0.06870264, 0.004508673, 5.910146e-11, 
    -2.718172e-05, 0.01860649, 0.09950249, 0.1024105, 0.09669403, 0.08916855, 
    0.1044712, 0.04111777, 0.02526059, 0.03981593, 0.09841435, 0.3046178, 
    0.00339374, 0.02079673, 0.04544188, 0.01215262, 0.051673, 0.08529771,
  0.3719439, 0.02795118, 0.0001067272, 0.03111853, 0.01495473, 0.04358573, 
    0.05160702, 0.06430754, 0.02162175, 0.02959487, 0.04743802, 0.02929073, 
    0.15206, 0.0606909, 0.03193697, 0.01816169, 0.01583469, 0.009374429, 
    0.007712436, 0.01489013, 0.04556886, 0.1923645, 0.2118362, 0.005448257, 
    9.844634e-07, -2.54198e-07, 0.002572377, 0.007726924, 0.09956174,
  0.3687949, 0.1004374, 0.003257853, 0.01995652, 0.03366698, 0.02265413, 
    0.04662263, 0.04097071, 0.02495234, 0.081836, 0.1002165, 0.07977946, 
    0.03469999, 0.02807396, 0.02454622, 0.01450707, 0.02022762, 0.01601471, 
    0.02167874, 0.02311775, 0.05751247, 0.2691202, 0.03929739, 0.06519251, 
    0.04075868, 0.02219255, 0.01809688, 0.04231627, 0.1289085,
  0.04489052, 0.0349778, 0.00559848, 0.1933002, -0.0001099513, 0.008627008, 
    0.0429854, 0.01268113, 0.0007630698, 0.01227528, 0.003805068, 0.07180306, 
    0.08309063, 0.06021395, 0.0359116, 0.05022377, 0.07495522, 0.1155217, 
    0.1041955, 0.1142274, 0.1400517, 0.09326253, 0.1369509, 0.04538086, 
    0.04300838, 0.0647573, 0.1395866, 0.1676713, 0.07056867,
  1.551213e-07, 3.555095e-08, 2.378482e-08, 2.315604e-09, 4.735797e-08, 
    0.05951853, 0.2051374, 0.08462903, 0.215722, 0.02691873, 0.06727541, 
    0.040852, 0.01755664, 0.008406108, 0.008727537, 0.01337552, 0.02291629, 
    0.09747235, 0.4405013, 0.2679122, 0.07820468, 0.08843945, 0.009255449, 
    0.005323697, 0.01968108, 0.03988183, 0.1882862, 0.1003294, -1.530868e-07,
  3.243078e-07, -1.631539e-05, -2.163224e-05, -2.804982e-08, 9.613785e-08, 
    -1.120077e-07, -0.000171127, 0.2831055, 0.3139714, 0.04425446, 0.1106149, 
    0.06644291, 0.109171, 0.04498275, 0.07943673, 0.04650248, 0.1003863, 
    0.2219022, 0.4311602, 0.005729245, 9.263699e-07, 0.009679157, 0.01741537, 
    0.04817971, 0.07862552, 0.08260384, 0.06901064, 0.3240301, -0.0008490196,
  -0.0005300931, 0.003095296, 0.005041625, 0.1785827, -6.947225e-05, 
    -5.633205e-08, 0.00406693, 1.105025e-06, -5.621139e-05, 0.03016375, 
    0.2245611, 0.06548174, 0.3871955, 0.3925686, 0.3929264, 0.4789221, 
    0.476053, 0.3866599, 0.3229005, 0.003131541, -0.0001057027, 0.004403139, 
    0.05985291, 0.1092306, 0.142965, 0.1811498, 0.1810317, 0.3777311, 
    0.08783336,
  0.1242101, 0.08940412, 0.03990248, 0.05472942, 0.004246473, 0.024701, 
    0.01912449, 0.1649157, 0.07367302, 0.01774939, 0.03524056, 0.1832208, 
    0.2897372, 0.3907409, 0.5106952, 0.5682673, 0.5855466, 0.5132779, 
    0.4892829, 0.06646441, 0.02391427, 0.02586262, 0.06624268, 0.1439417, 
    0.139253, 0.310743, 0.3726879, 0.4736965, 0.3490234,
  0.2796592, 0.1174046, 0.07346313, 0.06922181, 0.05691997, 0.02669448, 
    0.1206233, 0.1492085, 0.0807177, 0.1030985, 0.1143675, 0.2596846, 
    0.4036563, 0.3255586, 0.2260885, 0.5514532, 0.2640952, 0.3650023, 
    0.2933423, 0.06170021, 0.05482745, 0.1084719, 0.1594843, 0.2408352, 
    0.185394, 0.225604, 0.3794841, 0.4413255, 0.4304048,
  0.5601513, 0.4157969, 0.3010668, 0.2880434, 0.33922, 0.2920231, 0.2754912, 
    0.189027, 0.1327561, 0.2307029, 0.2538357, 0.3503886, 0.3144539, 
    0.3098672, 0.3434654, 0.3852281, 0.3133444, 0.1497284, 0.1595176, 
    0.2633566, 0.3703093, 0.3952205, 0.3220443, 0.3821939, 0.2432652, 
    0.3885117, 0.2875318, 0.338362, 0.6095093,
  0.5297551, 0.5396601, 0.4768395, 0.5400019, 0.6068063, 0.6242015, 
    0.6590892, 0.6110785, 0.6251673, 0.5605195, 0.5837862, 0.582101, 
    0.5943118, 0.5420534, 0.5334599, 0.5451918, 0.5186312, 0.4606344, 
    0.4817407, 0.5652398, 0.5115499, 0.4284079, 0.2866635, 0.4255223, 
    0.242185, 0.1718083, 0.2052558, 0.3532354, 0.5036977,
  0.3617402, 0.3591567, 0.3565732, 0.3539898, 0.3514063, 0.3488228, 
    0.3462393, 0.345708, 0.3447519, 0.3437957, 0.3428397, 0.3418836, 
    0.3409275, 0.3399714, 0.3495768, 0.3554351, 0.3612933, 0.3671516, 
    0.3730098, 0.3788681, 0.3847263, 0.3979757, 0.395657, 0.3933383, 
    0.3910197, 0.388701, 0.3863823, 0.3840636, 0.363807,
  0.1383659, 0.1534873, 0.1605961, 0.1469657, 0.1300232, 0.1137459, 
    0.1401971, 0.1257372, 0.04589931, 0.09652603, 0.09848002, 0.07958459, 
    0.1389201, 0.03881644, 0.117236, 0.1100603, 0.1070189, 0.09295741, 
    0.1404779, 0.1689547, 0.3751869, 0.4797868, 0.3517873, 0.2198121, 
    0.2142782, 0.2220531, 0.1679497, 0.1102215, 0.1477317,
  0.3828387, 0.2999939, 0.3773289, 0.08004151, 0.08913745, 0.09056022, 
    0.009809908, 0.2815424, 0.3536885, 0.3147259, 0.3767281, 0.3308172, 
    0.1554019, 0.2147981, 0.3268126, 0.3342724, 0.32897, 0.447677, 0.4406806, 
    0.3881612, 0.4227034, 0.3096234, 0.2832096, 0.4378684, 0.1680537, 
    0.2565883, 0.2875412, 0.3006828, 0.4195877,
  0.4042744, 0.4000178, 0.3229014, 0.2726935, 0.2362526, 0.2772164, 
    0.2750435, 0.3651496, 0.2488726, 0.1597304, 0.2661648, 0.3310784, 
    0.3129926, 0.3347636, 0.3190545, 0.268633, 0.3203453, 0.3763375, 
    0.2572581, 0.1822142, 0.2181719, 0.2107358, 0.1888788, 0.3034948, 
    0.2627471, 0.3840038, 0.4083329, 0.4318654, 0.4475037,
  0.315708, 0.4077853, 0.3929173, 0.4106795, 0.3915305, 0.3025188, 0.2244408, 
    0.1281583, 0.185932, 0.2270249, 0.2340516, 0.2098489, 0.197015, 
    0.1410171, 0.157438, 0.1172075, 0.110328, 0.1328454, 0.2069604, 
    0.2098939, 0.2006006, 0.2542223, 0.2457567, 0.2539659, 0.1465669, 
    0.2428375, 0.315977, 0.2963411, 0.3280165,
  0.1950585, 0.06830747, 0.03992307, 0.1026404, 0.08377009, 0.1005754, 
    0.0871673, 0.1180365, 0.1140787, 0.06636796, 0.04770009, 0.03325722, 
    0.01161166, 0.03860958, 0.3025144, 0.07193814, 0.1038233, 0.1419225, 
    0.1170558, 0.1539903, 0.1658431, 0.204262, 0.1837142, 0.3876232, 
    0.03456183, 0.06919283, 0.1105618, 0.1417876, 0.1507576,
  0.05302394, 0.02356108, 0.03225741, 0.02415935, 0.02433902, 0.01828594, 
    0.03573227, 0.03091195, 0.0557945, 0.003238928, -3.738528e-06, 
    -9.20628e-06, 0.0185508, 0.006061352, 0.01934474, 0.03421977, 0.07744739, 
    0.06548924, 0.1103092, 0.06601042, 0.03142923, 0.04839028, 0.06402569, 
    0.02916871, 0.03669608, 0.05183737, 0.03505667, 0.02842169, 0.02410267,
  0.06145316, 0.02113099, 6.660399e-05, 0.01171646, 0.003523028, 0.004917495, 
    0.01060546, 0.04119974, 0.02438978, 0.002109203, 5.117634e-11, 
    -2.181615e-05, 0.004724712, 0.06357975, 0.04819423, 0.04895313, 
    0.03816068, 0.03603248, 0.01222623, 0.004992512, 0.01235488, 0.03360586, 
    0.1231912, 0.0345244, 0.008402783, 0.05368793, 0.007235294, 0.01665928, 
    0.02822887,
  0.1719765, 0.141387, 7.532779e-05, 0.02245396, 0.004808895, 0.01209601, 
    0.02202059, 0.02493425, 0.005097428, 0.003810385, 0.02538052, 
    0.006251526, 0.1216998, 0.03412966, 0.01596468, 0.004365723, 0.005533124, 
    0.000784929, 0.0007559691, 0.00363296, 0.01188439, 0.06249727, 0.2334611, 
    0.001228571, 1.53931e-07, -3.289487e-08, -0.002803714, 0.0004508541, 
    0.03536141,
  0.1321645, 0.06909014, 0.00178188, 0.01201541, 0.01618256, 0.006297293, 
    0.006836374, 0.008141352, 0.04155243, 0.05713075, 0.030155, 0.01920297, 
    0.01815942, 0.008768772, 0.0114697, 0.002624568, 0.00537463, 0.003833134, 
    0.00649949, 0.01142214, 0.0313198, 0.3132552, 0.3178766, 0.03151796, 
    0.02927586, 0.002174258, 0.001869788, 0.009366098, 0.06231375,
  0.02928085, 0.03287152, 0.003285716, 0.1925773, -4.811856e-05, 0.001228077, 
    0.05311062, 0.002318725, -0.00132099, 0.00231933, 0.001163776, 
    0.01796912, 0.02835343, 0.01835684, 0.01601041, 0.03079216, 0.04339527, 
    0.06873418, 0.05607535, 0.06876431, 0.1071864, 0.09033886, 0.1902301, 
    0.03870932, 0.007605643, 0.03130411, 0.09360315, 0.1026213, 0.05713976,
  1.42297e-07, 3.298774e-08, 2.241701e-08, 8.529517e-10, 3.481723e-08, 
    0.06148892, 0.181036, 0.04548179, 0.2249862, 0.0223274, 0.0327108, 
    0.02569192, 0.004500117, 0.0006703568, 0.0009675788, 0.001546675, 
    0.004821999, 0.03198509, 0.2419678, 0.4654199, 0.1644627, 0.07310501, 
    0.001515961, 0.0003876934, 0.005142136, 0.009703196, 0.07274826, 
    0.086151, 3.796253e-08,
  3.096517e-07, -7.543254e-05, 5.491502e-05, -5.508819e-07, 8.870938e-08, 
    -3.59583e-08, -0.002437642, 0.2813126, 0.3187256, 0.03906068, 0.08899718, 
    0.05438311, 0.06879688, 0.02282155, 0.0508964, 0.0318051, 0.03722961, 
    0.1269051, 0.2655593, 0.2301213, -6.408413e-06, 0.004183036, 0.009639943, 
    0.005852835, 0.01799677, 0.01375612, 0.01231955, 0.1625428, 0.0009911794,
  -0.001032754, 0.00144152, 0.003070849, 0.1998729, -5.515407e-05, 
    7.20709e-10, 0.003366089, 9.845129e-07, -4.981189e-05, 0.02769888, 
    0.2518016, 0.08491318, 0.4515036, 0.547496, 0.4693677, 0.5400321, 
    0.4552556, 0.2877274, 0.3713159, 0.001155516, -0.0001006954, 0.004919177, 
    0.04588509, 0.1518893, 0.1778707, 0.1723999, 0.1161783, 0.2474947, 
    0.1080819,
  0.1299243, 0.06842668, 0.03323144, 0.03884167, 0.002308974, 0.01449634, 
    0.01410179, 0.1677385, 0.05963159, 0.01972824, 0.03823126, 0.1673025, 
    0.3983879, 0.5221571, 0.711403, 0.6722047, 0.686927, 0.5170817, 
    0.3777843, 0.06836052, 0.01862878, 0.01495305, 0.0651931, 0.1264058, 
    0.1442312, 0.4065016, 0.3749042, 0.4807774, 0.3197416,
  0.2781636, 0.1029476, 0.05252919, 0.05132955, 0.04963585, 0.01649274, 
    0.1085321, 0.1261207, 0.06498081, 0.09098791, 0.1007301, 0.2650275, 
    0.4452996, 0.3509616, 0.284171, 0.6689566, 0.2465055, 0.3440014, 
    0.2682356, 0.05079067, 0.0442418, 0.09814034, 0.1667188, 0.2141034, 
    0.2283643, 0.2273431, 0.3685842, 0.4010804, 0.4210087,
  0.5825889, 0.3944027, 0.2898039, 0.3064758, 0.3684457, 0.3060351, 0.258774, 
    0.1430188, 0.09242149, 0.174098, 0.2166177, 0.311589, 0.2999388, 
    0.2966421, 0.3578269, 0.4247029, 0.2850348, 0.1743268, 0.2373387, 
    0.257571, 0.3647581, 0.3634644, 0.2710839, 0.3734445, 0.2862253, 0.38043, 
    0.2640254, 0.3519894, 0.6673101,
  0.5859374, 0.5375736, 0.4756262, 0.6396128, 0.6796308, 0.679133, 0.6530554, 
    0.6210486, 0.6546491, 0.6352651, 0.6410703, 0.6388587, 0.648093, 
    0.5777162, 0.5908328, 0.6097146, 0.6091287, 0.6042949, 0.6519954, 
    0.6958514, 0.5904385, 0.4995421, 0.2508722, 0.4866375, 0.3066045, 
    0.169551, 0.2316513, 0.4531196, 0.5622666,
  0.2153607, 0.2094314, 0.203502, 0.1975727, 0.1916434, 0.1857141, 0.1797848, 
    0.1854236, 0.1914522, 0.1974807, 0.2035092, 0.2095378, 0.2155663, 
    0.2215948, 0.2556795, 0.262392, 0.2691046, 0.2758172, 0.2825298, 
    0.2892424, 0.295955, 0.324335, 0.3175232, 0.3107114, 0.3038996, 
    0.2970878, 0.2902759, 0.2834641, 0.2201041,
  0.1496406, 0.1279042, 0.1467897, 0.1357265, 0.1643043, 0.09526524, 
    0.1223057, 0.1262812, 0.03950142, 0.04667397, 0.06053007, 0.06121079, 
    0.1510386, 0.02531844, 0.127505, 0.1165333, 0.1528992, 0.1418127, 
    0.1747154, 0.1798455, 0.4012872, 0.5144444, 0.3229707, 0.1989917, 
    0.2537981, 0.2626437, 0.1932654, 0.1117268, 0.1417569,
  0.3510015, 0.2550512, 0.2944477, 0.04998814, 0.06747194, 0.08287068, 
    0.004164658, 0.2399765, 0.3420117, 0.2842283, 0.3525026, 0.3321889, 
    0.1148703, 0.1816315, 0.341752, 0.3617892, 0.361424, 0.4774465, 
    0.4095725, 0.3981017, 0.4205576, 0.3374362, 0.2994995, 0.4523402, 
    0.1743581, 0.3087287, 0.369019, 0.3964386, 0.4419927,
  0.4362466, 0.3963698, 0.2532974, 0.2389597, 0.1965167, 0.2116031, 
    0.2607381, 0.3390163, 0.2086266, 0.1367058, 0.2316199, 0.304508, 
    0.2983915, 0.3093503, 0.2897055, 0.2521197, 0.2853392, 0.3294569, 
    0.2228862, 0.1443844, 0.1776115, 0.1753041, 0.1724039, 0.2623857, 
    0.2471554, 0.3956459, 0.4266567, 0.4652029, 0.4919781,
  0.2760578, 0.3622478, 0.3470578, 0.3722609, 0.3600334, 0.2667491, 
    0.1864192, 0.1029849, 0.1536212, 0.1959121, 0.1826826, 0.1675864, 
    0.1620857, 0.1059219, 0.1237955, 0.09812151, 0.07966122, 0.09732128, 
    0.1614535, 0.1801256, 0.1776944, 0.222136, 0.2183672, 0.2214445, 
    0.1168374, 0.2034024, 0.2855388, 0.2701784, 0.30656,
  0.1591008, 0.03707909, 0.02775117, 0.0677291, 0.05305333, 0.06698193, 
    0.0604751, 0.07337813, 0.07786225, 0.04293165, 0.03333305, 0.02006985, 
    0.005706838, 0.02723796, 0.2378351, 0.04697265, 0.07566414, 0.1188366, 
    0.08535155, 0.1264612, 0.1380479, 0.1718015, 0.1410838, 0.3836365, 
    0.02451709, 0.04422718, 0.08124985, 0.1041866, 0.1112525,
  0.02154932, 0.007632617, 0.02711988, 0.00958637, 0.0106868, 0.009961965, 
    0.02452857, 0.01673171, 0.03572989, 0.001908904, -1.06982e-05, 
    -2.919973e-05, 0.01616373, 0.004515382, 0.01367578, 0.02252285, 
    0.06019066, 0.04965824, 0.07887049, 0.04788528, 0.01990738, 0.02323616, 
    0.03354578, 0.02363496, 0.0332696, 0.03996737, 0.02279988, 0.01378589, 
    0.009803339,
  0.02694639, 0.02166033, -1.562282e-05, 0.004330229, 0.0003902287, 
    0.001747658, 0.003140808, 0.02050528, 0.009271569, 0.0008116545, 
    1.021938e-10, -9.97944e-06, 0.001599214, 0.03364729, 0.02083609, 
    0.01987782, 0.01275417, 0.007373384, 0.00564039, 0.001573161, 
    0.005271267, 0.01236915, 0.04900958, 0.03389286, 0.00362245, 0.06465587, 
    0.002541802, 0.006980114, 0.01123444,
  0.08117831, 0.1134173, 0.0003685936, 0.01803388, 0.001075606, 0.004145362, 
    0.008668613, 0.009522419, 0.00146, 0.0001529478, 0.01252404, 0.001117165, 
    0.08551297, 0.01531413, 0.006085949, 0.001402285, 0.001825551, 
    0.0002978987, 0.0003142243, 0.001516628, 0.004411512, 0.02438463, 
    0.1068459, 0.0005071192, -1.286345e-07, 1.103448e-08, -0.001577422, 
    0.0001130232, 0.01509625,
  0.04890013, 0.05068066, 0.001519926, 0.0064638, 0.002238905, 0.001368201, 
    0.002350327, 0.001756766, 0.04177184, 0.04450495, 0.007547541, 
    0.003264561, 0.009339082, 0.007373221, 0.008228613, 0.0006079634, 
    0.0005747119, 0.0004048955, 0.0007012971, 0.0009760194, 0.004928382, 
    0.1301381, 0.1736126, 0.02209727, 0.02439459, 0.0003245633, 0.0001497456, 
    0.001303677, 0.01096417,
  0.01747733, 0.03297408, 0.002209374, 0.2034791, -1.056801e-05, 
    5.029687e-05, 0.05728427, 9.446037e-05, -0.001243129, 0.0005031791, 
    0.0001541314, 0.005473849, 0.008500707, 0.005434125, 0.006781379, 
    0.01821313, 0.02608719, 0.03511046, 0.03512809, 0.03176951, 0.06420612, 
    0.03184978, 0.2397768, 0.02836735, 0.0009562778, 0.01235818, 0.03260161, 
    0.04504283, 0.05743104,
  1.348378e-07, 3.119708e-08, 2.154302e-08, 3.60364e-10, 3.149603e-08, 
    0.00642888, 0.128836, 0.0184934, 0.2342247, 0.01003175, 0.01293044, 
    0.01209493, 0.0005687231, -4.925266e-06, 9.90187e-05, 0.0002380297, 
    0.001593241, 0.01275446, 0.1271608, 0.2948564, 0.04416211, 0.05823045, 
    0.0005489734, -0.0009830524, 0.001226354, 0.002407806, 0.02492243, 
    0.04876544, 1.168799e-07,
  2.999975e-07, -6.175529e-05, 0.0001379485, -9.298822e-07, 8.371359e-08, 
    -9.163772e-10, -0.002050939, 0.2631794, 0.3116757, 0.03211705, 
    0.05892168, 0.01801913, 0.03586654, 0.00932934, 0.01183329, 0.006480565, 
    0.01388793, 0.05191413, 0.1166672, 0.2649399, 6.421988e-06, 0.001139193, 
    0.004575668, 0.001143044, 0.003866266, 0.004366814, 0.003919324, 
    0.07295573, 0.003727124,
  -0.001050014, 0.0004691511, 0.0009952174, 0.2137997, -5.773698e-05, 
    1.243377e-08, 0.002356706, 9.578736e-07, -3.921401e-05, 0.0234424, 
    0.2762006, 0.1264227, 0.5495993, 0.6261411, 0.5429084, 0.4491001, 
    0.3480993, 0.1918711, 0.2446445, 0.0005022178, -0.0001143033, 
    0.004598459, 0.03755295, 0.1693006, 0.1171211, 0.1462322, 0.07094637, 
    0.1347072, 0.1065398,
  0.1295806, 0.05966073, 0.02814657, 0.02528042, 0.001013435, 0.006157552, 
    0.009172956, 0.1514595, 0.05108942, 0.02240214, 0.03394173, 0.1606087, 
    0.5652546, 0.6031076, 0.784817, 0.6591767, 0.6865959, 0.4540898, 
    0.2943805, 0.07025488, 0.013242, 0.008658934, 0.0592369, 0.1108089, 
    0.145912, 0.4403582, 0.3679233, 0.4668519, 0.291478,
  0.2351673, 0.08863444, 0.04016404, 0.03390701, 0.04091993, 0.01094654, 
    0.0949447, 0.1084297, 0.05285398, 0.08120508, 0.09408683, 0.2725951, 
    0.4549794, 0.3377624, 0.3753403, 0.7296476, 0.2350799, 0.3149626, 
    0.2441944, 0.04441449, 0.03329258, 0.09316996, 0.1878419, 0.1846164, 
    0.2625903, 0.2231503, 0.3230534, 0.3570865, 0.3827665,
  0.5950993, 0.3759687, 0.262176, 0.2515424, 0.3509574, 0.2921946, 0.2272589, 
    0.1136361, 0.07336359, 0.1388769, 0.1708824, 0.2747387, 0.2600921, 
    0.2991944, 0.3925592, 0.3861616, 0.2560893, 0.244395, 0.2809005, 
    0.2451134, 0.3289326, 0.3812246, 0.2285784, 0.3471342, 0.3612788, 
    0.3544883, 0.2284672, 0.3445371, 0.6559324,
  0.5653106, 0.4290563, 0.5258231, 0.6317275, 0.6352857, 0.6756567, 
    0.6450062, 0.6284469, 0.6453456, 0.6174866, 0.6283579, 0.6553645, 
    0.6753824, 0.5876059, 0.6139921, 0.6141595, 0.6534009, 0.655934, 
    0.6456422, 0.6245809, 0.6126712, 0.4595977, 0.1872443, 0.4239225, 
    0.2984222, 0.1878597, 0.2420944, 0.5176029, 0.5640803,
  0.1088469, 0.1050996, 0.1013524, 0.09760512, 0.09385785, 0.09011059, 
    0.08636332, 0.07237325, 0.078968, 0.08556275, 0.09215751, 0.09875226, 
    0.105347, 0.1119418, 0.1171891, 0.1215309, 0.1258726, 0.1302143, 
    0.1345561, 0.1388978, 0.1432396, 0.1577201, 0.1505309, 0.1433417, 
    0.1361524, 0.1289632, 0.121774, 0.1145848, 0.1118447,
  0.1408638, 0.1114772, 0.09382199, 0.1195962, 0.1282496, 0.08315786, 
    0.100616, 0.1235511, 0.02093117, 0.0211061, 0.04482591, 0.07985314, 
    0.1365293, 0.013219, 0.1625617, 0.1719732, 0.2023368, 0.180907, 
    0.1817555, 0.2046867, 0.4149312, 0.5490335, 0.2713513, 0.1764455, 
    0.250313, 0.3346728, 0.1862669, 0.1037849, 0.1347601,
  0.3074715, 0.2041989, 0.2244881, 0.0342613, 0.04410474, 0.07816404, 
    0.001678207, 0.18673, 0.3399846, 0.2585168, 0.3037617, 0.3279039, 
    0.08618055, 0.153201, 0.3416246, 0.3530822, 0.3726217, 0.4530495, 
    0.3683291, 0.4105369, 0.3803118, 0.3536494, 0.3112559, 0.4517628, 
    0.1630246, 0.3462551, 0.4109849, 0.4786026, 0.4335979,
  0.4108361, 0.3653119, 0.1982093, 0.1903906, 0.1529025, 0.1555476, 
    0.2584056, 0.2876276, 0.173194, 0.1093865, 0.1947506, 0.2589885, 
    0.2531779, 0.2764333, 0.2509883, 0.2224055, 0.2376872, 0.2736477, 
    0.1896363, 0.1056093, 0.1423583, 0.1313001, 0.1449766, 0.218039, 
    0.2248882, 0.3842322, 0.4233702, 0.4745043, 0.4716766,
  0.2358217, 0.2960607, 0.296387, 0.3329685, 0.3139971, 0.2144843, 0.1491563, 
    0.0772476, 0.1193976, 0.1501148, 0.1306084, 0.1172448, 0.1105231, 
    0.07302839, 0.08750726, 0.07895969, 0.05272282, 0.06689775, 0.1172088, 
    0.1351048, 0.1478944, 0.1939433, 0.1797503, 0.1872451, 0.07872213, 
    0.1532979, 0.2394861, 0.2203399, 0.2757739,
  0.1122509, 0.02029041, 0.01844172, 0.04041772, 0.03184171, 0.04043463, 
    0.03296853, 0.041876, 0.04684506, 0.02886868, 0.02546592, 0.01068711, 
    0.002746205, 0.01885046, 0.1847744, 0.03103455, 0.05445635, 0.0945183, 
    0.0619718, 0.09529877, 0.1057155, 0.1297394, 0.08983599, 0.3637067, 
    0.02016386, 0.03021626, 0.05608507, 0.06714062, 0.07726371,
  0.01154485, 0.002589346, 0.02303739, 0.005225331, 0.003900005, 0.006518988, 
    0.0152109, 0.009750731, 0.02250042, 0.001327314, -1.345335e-05, 
    -1.687875e-05, 0.0130878, 0.002697718, 0.008905591, 0.01526304, 
    0.04212357, 0.03629292, 0.05327713, 0.02700627, 0.01280023, 0.00954862, 
    0.01831563, 0.01489482, 0.02664918, 0.02058241, 0.009907354, 0.006086303, 
    0.005221087,
  0.01583698, 0.01642274, -2.467979e-05, 0.002299515, -0.00112163, 
    0.0006836837, 0.001246204, 0.01079871, 0.004262296, 0.00042694, 
    1.109676e-10, -3.181038e-06, 0.0009181913, 0.01451548, 0.009539291, 
    0.008272198, 0.005351767, 0.002864925, 0.002818497, 0.0008397329, 
    0.002303918, 0.00590903, 0.02629965, 0.02859288, 0.002331675, 0.06610505, 
    0.000955001, 0.003184542, 0.005984305,
  0.04562482, 0.06937375, 0.0005029056, 0.01312369, 0.0001268096, 
    0.001014211, 0.003507388, 0.002951805, 0.000591986, -0.0001230447, 
    0.007573788, 0.0004509073, 0.04456481, 0.005704758, 0.002163347, 
    0.0004749004, 0.0006510309, 0.0001713188, 0.0001751443, 0.0008035242, 
    0.002237803, 0.01276198, 0.05994137, 0.0004207208, -2.979514e-06, 
    1.179921e-08, -0.001015904, 4.946563e-05, 0.008363839,
  0.02435477, 0.04534165, 0.001193444, 0.002928435, 0.0001709112, 
    0.0006239614, 0.001284303, 0.0007862588, 0.03455542, 0.04950992, 
    0.002531183, 0.001357632, 0.005410143, 0.004749769, 0.004682046, 
    0.0002798444, 0.0002174762, 0.0001144326, 0.0003292613, 0.0002017595, 
    0.001490849, 0.05225784, 0.09114993, 0.02425772, 0.03091716, 
    0.0001636997, 6.728306e-05, 0.0006219246, 0.004117484,
  0.0107492, 0.0272899, 0.001052971, 0.2023634, -3.561929e-06, 1.010109e-05, 
    0.0449274, 1.522026e-05, -0.0004682817, 0.0002378279, 1.982439e-05, 
    0.002308715, 0.003663553, 0.001644279, 0.002811571, 0.01117071, 
    0.0125691, 0.02034562, 0.02273512, 0.01281502, 0.03088885, 0.01163725, 
    0.2117409, 0.0222767, 0.0003141583, 0.006593566, 0.01454023, 0.02118941, 
    0.0442579,
  1.274703e-07, 3.007161e-08, 2.092556e-08, 2.090328e-11, 3.100791e-08, 
    0.001087322, 0.06356609, 0.005166671, 0.2116558, 0.0017473, 0.005930555, 
    0.00483369, 0.0001653916, -1.20538e-06, 4.859638e-05, 0.0001036299, 
    0.000749933, 0.006511558, 0.07253543, 0.1607074, 0.0214478, 0.04784984, 
    0.0003087987, -0.001088104, 0.0003826348, 0.0009791538, 0.01072136, 
    0.03018329, 1.21685e-07,
  2.9327e-07, -2.825881e-06, 0.0009663907, -1.710053e-06, 8.045879e-08, 
    2.377639e-09, -0.00279382, 0.2333161, 0.2940192, 0.02020111, 0.06675421, 
    0.009873299, 0.01523155, 0.002572687, 0.003528549, 0.001352679, 
    0.006672028, 0.02501271, 0.05761937, 0.175895, 1.1129e-06, 0.000413746, 
    0.002358578, 0.0004093401, 0.001772858, 0.002360577, 0.002054587, 
    0.03495244, 0.0040187,
  -0.0008345894, 7.203439e-05, 0.0002154953, 0.20327, -5.061991e-05, 
    1.185105e-08, 0.00138305, 9.642476e-07, -2.692913e-05, 0.01808785, 
    0.2770875, 0.2114978, 0.5752453, 0.586791, 0.4846178, 0.3689589, 
    0.2563036, 0.1648124, 0.1657561, 0.00182103, -0.0001036768, 0.003116465, 
    0.0317191, 0.1511638, 0.07032223, 0.08154552, 0.02918228, 0.0667002, 
    0.09784327,
  0.1042797, 0.04702177, 0.01919581, 0.01400956, 0.0003816853, 0.002209329, 
    0.004893612, 0.1346037, 0.04531101, 0.02445631, 0.03585041, 0.1455887, 
    0.6377694, 0.61185, 0.7159677, 0.5931665, 0.5925037, 0.3740901, 
    0.2413753, 0.06373294, 0.008676843, 0.004400709, 0.04909897, 0.09662271, 
    0.1478103, 0.4539511, 0.3575107, 0.4160733, 0.26594,
  0.1667838, 0.07529371, 0.02990561, 0.02154865, 0.03455736, 0.00922397, 
    0.08418041, 0.09712481, 0.04761497, 0.07519288, 0.09200812, 0.2536575, 
    0.4480277, 0.3135251, 0.4526026, 0.722241, 0.2132528, 0.280421, 0.195542, 
    0.04294002, 0.02433098, 0.08955936, 0.2372559, 0.1494372, 0.2785271, 
    0.2167065, 0.2775139, 0.310595, 0.3221135,
  0.566789, 0.353642, 0.2285468, 0.2298957, 0.3399266, 0.3179046, 0.1856091, 
    0.09063239, 0.06104139, 0.1146981, 0.1386803, 0.2317434, 0.2255185, 
    0.3090822, 0.3806322, 0.3712137, 0.2287846, 0.3045749, 0.2826506, 
    0.2308423, 0.2583206, 0.3730511, 0.1916692, 0.3296003, 0.4169371, 
    0.3065461, 0.1905841, 0.328123, 0.6081567,
  0.5776352, 0.3945624, 0.4972169, 0.6017081, 0.56172, 0.6385328, 0.691795, 
    0.6303123, 0.6376181, 0.6345653, 0.6180805, 0.6647699, 0.6704503, 
    0.6147646, 0.6136701, 0.6103399, 0.6479477, 0.6541075, 0.5922518, 
    0.5686816, 0.5720673, 0.389039, 0.1518653, 0.3526908, 0.2663208, 
    0.1788727, 0.2425303, 0.5018646, 0.555146,
  0.06157084, 0.05859252, 0.05561421, 0.05263589, 0.04965757, 0.04667926, 
    0.04370094, 0.03555692, 0.03746512, 0.03937331, 0.04128151, 0.0431897, 
    0.04509789, 0.04700609, 0.04893584, 0.05282786, 0.05671988, 0.0606119, 
    0.06450393, 0.06839595, 0.07228798, 0.06948602, 0.06666412, 0.06384222, 
    0.06102033, 0.05819843, 0.05537653, 0.05255463, 0.06395349,
  0.1128692, 0.09530069, 0.0555566, 0.07591258, 0.07245249, 0.06545538, 
    0.07852213, 0.08890609, 0.03124996, 0.01705839, 0.0196008, 0.08155773, 
    0.1117494, 0.008269981, 0.1887605, 0.2522455, 0.2413242, 0.2017786, 
    0.1657746, 0.1956088, 0.4586862, 0.5684311, 0.2238982, 0.1312849, 
    0.2706109, 0.408549, 0.1913636, 0.08555074, 0.1273826,
  0.2484381, 0.1638754, 0.1643388, 0.02609182, 0.03081217, 0.07412963, 
    0.001495546, 0.1358923, 0.3150848, 0.236571, 0.2856219, 0.296632, 
    0.06585309, 0.1233488, 0.3342778, 0.3256878, 0.3285304, 0.3709375, 
    0.3164943, 0.4080731, 0.3309833, 0.3504006, 0.3193659, 0.4417105, 
    0.16745, 0.3519391, 0.3896955, 0.4835603, 0.3725024,
  0.3559808, 0.3077239, 0.1499659, 0.1394458, 0.1083, 0.117111, 0.2317594, 
    0.2445704, 0.1401142, 0.0829829, 0.1513133, 0.2120365, 0.192439, 
    0.2248928, 0.197301, 0.1824028, 0.1823843, 0.2139724, 0.145807, 
    0.07831676, 0.1089837, 0.09401403, 0.1081286, 0.1701032, 0.1914977, 
    0.3522665, 0.3780089, 0.4379774, 0.4182739,
  0.2016278, 0.229506, 0.2541234, 0.2804847, 0.2564195, 0.1625428, 0.1147649, 
    0.05541033, 0.08924549, 0.1100197, 0.08896028, 0.07156633, 0.06433308, 
    0.04288861, 0.05268171, 0.05395519, 0.0326217, 0.0438201, 0.07955539, 
    0.08929189, 0.1110335, 0.1402744, 0.1309175, 0.1601623, 0.04759292, 
    0.1152977, 0.1871526, 0.1718217, 0.2458878,
  0.07835416, 0.0114615, 0.01339865, 0.02235684, 0.01853943, 0.02277285, 
    0.01874797, 0.02509183, 0.02581104, 0.01710067, 0.01528151, 0.005492264, 
    0.001559843, 0.011347, 0.1449911, 0.01883454, 0.03578078, 0.06865524, 
    0.04215515, 0.06660762, 0.0725921, 0.08710149, 0.05295413, 0.3395848, 
    0.01468124, 0.0179758, 0.03630028, 0.03776814, 0.04709496,
  0.007494041, 0.001508192, 0.01765551, 0.003377308, 0.001866039, 
    0.004122145, 0.009706102, 0.006409109, 0.01121082, 0.00100645, 
    -6.779464e-05, -1.78896e-05, 0.00972207, 0.001412002, 0.004368738, 
    0.008476635, 0.02567414, 0.02233294, 0.03190465, 0.01254412, 0.004867348, 
    0.004366259, 0.0116726, 0.009556354, 0.02063414, 0.008446349, 0.00404838, 
    0.002778234, 0.003264465,
  0.01076836, 0.01158926, -2.218035e-05, 0.001560966, -0.001483894, 
    0.0003558448, 0.0007136385, 0.00454043, 0.002481887, 0.0002909077, 
    1.31168e-10, -1.351836e-06, 0.0006442349, 0.006403429, 0.004319127, 
    0.003477424, 0.002396374, 0.001720723, 0.001276425, 0.0005542761, 
    0.001332234, 0.003565188, 0.01731813, 0.02333538, 0.002570064, 
    0.05837523, 0.0004588608, 0.001804317, 0.003865886,
  0.03037186, 0.0406929, 0.0003750026, 0.008456844, 2.863064e-05, 
    0.000427028, 0.001300158, 0.001250051, 0.0003036559, -7.433681e-05, 
    0.004517019, 0.0002545904, 0.01869437, 0.001867994, 0.0006942404, 
    0.0001997423, 0.000263259, 0.0001153062, 0.0001153549, 0.0005137667, 
    0.00140262, 0.008183644, 0.03934407, 0.00141487, -1.436421e-06, 
    1.132981e-08, -0.0005525744, 2.868894e-05, 0.005529733,
  0.01539978, 0.04092987, 0.001120499, 0.001288157, 6.444068e-05, 
    0.0003990336, 0.0008386222, 0.0004971005, 0.02223494, 0.04949411, 
    0.001353451, 0.0007920751, 0.002583476, 0.002429535, 0.002135317, 
    0.0002091495, 0.0001374867, 7.049609e-05, 0.0002010758, 0.0001079907, 
    0.0007971117, 0.02781389, 0.05937847, 0.02494685, 0.03511036, 
    0.0001083027, 4.06603e-05, 0.0003828211, 0.00241169,
  0.006292129, 0.01663794, 0.0003305849, 0.1796839, -1.601088e-06, 
    4.545815e-06, 0.0267585, 7.232746e-06, -0.0001681626, 0.0001410801, 
    1.194527e-05, 0.001267576, 0.001722247, 0.0006755709, 0.0009690937, 
    0.005236076, 0.005646079, 0.01098255, 0.01182975, 0.005059161, 
    0.01306322, 0.004440405, 0.1750303, 0.02501579, 0.0001798056, 
    0.003177028, 0.006734813, 0.01000076, 0.03064593,
  1.230926e-07, 2.934387e-08, 2.047558e-08, -2.441969e-10, 3.076351e-08, 
    0.0004679343, 0.01837347, 0.001433457, 0.152208, 0.0004373221, 
    0.002567296, 0.001107128, 7.668243e-05, 6.310236e-07, 2.917901e-05, 
    6.100072e-05, 0.0004551802, 0.003168105, 0.04163817, 0.08750445, 
    0.0105621, 0.03703971, 0.0002045087, -0.001042904, 0.0001348458, 
    0.0005576649, 0.006077277, 0.01621304, 1.193677e-07,
  2.891443e-07, 3.408415e-06, 0.001480995, -2.22888e-06, 7.844528e-08, 
    2.251171e-09, -0.003427361, 0.2040001, 0.260843, 0.01174609, 0.05059787, 
    0.006904236, 0.004989022, 0.001324978, 0.001810168, 0.0007195332, 
    0.003982949, 0.0150198, 0.03429606, 0.1220467, -9.466784e-07, 
    0.0007428179, 0.001465685, 0.0002472433, 0.00109912, 0.001571803, 
    0.001349204, 0.02072131, 0.003930038,
  -0.0006149236, -6.966142e-05, -4.478632e-05, 0.1878634, -4.19986e-05, 
    1.153309e-08, 0.0007454009, 9.436783e-07, -1.851553e-05, 0.0117091, 
    0.2562256, 0.2719858, 0.5301136, 0.5259427, 0.402316, 0.3016191, 
    0.1719161, 0.1292378, 0.1137628, 0.001543675, -6.392763e-05, 0.001758043, 
    0.02180712, 0.1313705, 0.03903867, 0.03656306, 0.01107479, 0.03686926, 
    0.0809689,
  0.07631549, 0.03234093, 0.01524565, 0.006789085, 0.0001727391, 0.001067413, 
    0.002474682, 0.125931, 0.03845872, 0.02168944, 0.03478416, 0.1258995, 
    0.6090064, 0.5701859, 0.6273124, 0.4852394, 0.4320893, 0.2658047, 
    0.1762196, 0.05557942, 0.006356097, 0.002255861, 0.03829414, 0.07718748, 
    0.1520506, 0.40416, 0.2870888, 0.3149147, 0.2062817,
  0.1191234, 0.05979616, 0.01942722, 0.01366664, 0.02946022, 0.01187397, 
    0.068197, 0.08335462, 0.04633552, 0.06648213, 0.08725297, 0.2219939, 
    0.4245436, 0.2719944, 0.492465, 0.6148791, 0.1827408, 0.2474984, 
    0.1317776, 0.03731563, 0.01877482, 0.08106932, 0.2768424, 0.1210337, 
    0.2982509, 0.2007534, 0.2118252, 0.2400704, 0.2326454,
  0.4690737, 0.2954933, 0.1925459, 0.2130139, 0.340663, 0.4069498, 0.1485365, 
    0.06820745, 0.04984186, 0.09419389, 0.1104906, 0.1952139, 0.1990744, 
    0.2996388, 0.3559285, 0.3382278, 0.1873901, 0.3033371, 0.2934454, 
    0.2423032, 0.1959862, 0.354702, 0.1545736, 0.3032347, 0.3871447, 
    0.263199, 0.1677129, 0.3055037, 0.5348902,
  0.5545886, 0.3494624, 0.419138, 0.5487894, 0.4878587, 0.5676509, 0.6692324, 
    0.6140918, 0.6124959, 0.6197401, 0.5748131, 0.6074207, 0.608235, 
    0.5535924, 0.5363376, 0.5609047, 0.5647518, 0.5706628, 0.4995225, 
    0.4782394, 0.4976035, 0.325407, 0.1264843, 0.2914785, 0.239935, 
    0.1655939, 0.2292967, 0.4520253, 0.5310248,
  0.03505328, 0.03292828, 0.03080329, 0.02867829, 0.0265533, 0.0244283, 
    0.02230331, 0.007307196, 0.008067641, 0.008828087, 0.009588532, 
    0.01034898, 0.01110942, 0.01186987, 0.0179125, 0.02050726, 0.02310202, 
    0.02569677, 0.02829153, 0.03088628, 0.03348104, 0.04002209, 0.03879188, 
    0.03756168, 0.03633147, 0.03510127, 0.03387106, 0.03264086, 0.03675328,
  0.1021594, 0.07812624, 0.02261529, 0.04158026, 0.05145697, 0.05094141, 
    0.0628814, 0.03268674, 0.02208889, 0.0157183, 0.01507861, 0.06874411, 
    0.0903502, 0.004626061, 0.2440147, 0.2513964, 0.2271319, 0.2236593, 
    0.1500857, 0.2396312, 0.5058821, 0.5725491, 0.201923, 0.1050233, 
    0.3206761, 0.4485282, 0.1933128, 0.06343085, 0.09277356,
  0.2020329, 0.1311905, 0.1285879, 0.02157205, 0.0198475, 0.06896826, 
    0.001393334, 0.1142682, 0.2784537, 0.2211834, 0.2663349, 0.2807753, 
    0.05409815, 0.1024194, 0.311652, 0.3065823, 0.2751406, 0.3051821, 
    0.2636572, 0.3633128, 0.2965129, 0.3214675, 0.3017925, 0.4247591, 
    0.1561743, 0.342483, 0.3370048, 0.3967181, 0.2998423,
  0.3012634, 0.2556286, 0.1207744, 0.1111899, 0.08358298, 0.09514232, 
    0.2113059, 0.2139276, 0.1122216, 0.06868408, 0.1220814, 0.1799509, 
    0.1520518, 0.1854418, 0.1503491, 0.142612, 0.1441677, 0.1738389, 
    0.1183084, 0.06156812, 0.08720604, 0.07517039, 0.08437937, 0.1341156, 
    0.1625165, 0.3220254, 0.3354351, 0.3880773, 0.3592029,
  0.1758533, 0.1890089, 0.2166386, 0.2385491, 0.2120568, 0.1337268, 
    0.09425074, 0.04164558, 0.07098381, 0.08346511, 0.06435175, 0.04811487, 
    0.04094295, 0.02757751, 0.03623496, 0.03649019, 0.02255988, 0.02706608, 
    0.05460985, 0.06377139, 0.08172469, 0.1028144, 0.09341498, 0.1546591, 
    0.03162127, 0.0885654, 0.1490611, 0.1403241, 0.2135597,
  0.0534455, 0.007452558, 0.01054878, 0.01279017, 0.01214249, 0.01380968, 
    0.01100496, 0.01624609, 0.01646176, 0.01101339, 0.009215429, 0.003482437, 
    0.001199647, 0.007107377, 0.1208571, 0.01126842, 0.02027033, 0.04765211, 
    0.02708363, 0.04621951, 0.04664091, 0.0614211, 0.03291192, 0.3149194, 
    0.009231516, 0.01111494, 0.02385701, 0.02271204, 0.0282963,
  0.005665439, 0.001091402, 0.01464304, 0.002225091, 0.001315145, 
    0.002213762, 0.006366022, 0.004885712, 0.005688957, 0.0008128181, 
    0.0001374842, -1.416031e-05, 0.009137728, 0.0006996676, 0.002125856, 
    0.00484154, 0.01549008, 0.01245789, 0.0187133, 0.006320253, 0.002668498, 
    0.002735332, 0.008532412, 0.007218906, 0.01713477, 0.004328744, 
    0.002179361, 0.001784429, 0.002386825,
  0.008198988, 0.008776663, -1.943854e-05, 0.001195031, -0.001251494, 
    0.0002490545, 0.0005061373, 0.002552907, 0.001719881, 0.000224744, 
    1.460598e-10, -6.747048e-07, 0.0004998056, 0.003431173, 0.002354604, 
    0.001974114, 0.00149526, 0.001237649, 0.000836101, 0.0004141068, 
    0.000945156, 0.002525402, 0.01291728, 0.02000389, 0.002389678, 
    0.05151621, 0.0002715074, 0.001238615, 0.002846756,
  0.02279903, 0.02575296, 0.0002032373, 0.005129271, 1.770749e-05, 
    0.0002771413, 0.0006836465, 0.0006909849, 0.0002022921, -6.19737e-06, 
    0.00267476, 0.0001885095, 0.009119974, 0.0007390496, 0.0003062297, 
    0.000127742, 0.0001514285, 8.721706e-05, 8.629406e-05, 0.0003764472, 
    0.001016029, 0.006004929, 0.02935433, 0.004811014, -5.132563e-07, 
    1.150843e-08, -0.000295562, 1.972187e-05, 0.004148074,
  0.01121853, 0.04304994, 0.0006941147, 0.0005774936, 3.781565e-05, 
    0.0002961236, 0.000619438, 0.0003647826, 0.01785162, 0.05847623, 
    0.000891596, 0.0004733432, 0.001350875, 0.001176591, 0.0009727489, 
    0.0001341229, 0.0001005406, 5.077914e-05, 0.0001431702, 7.229962e-05, 
    0.0005278625, 0.01862947, 0.04375745, 0.02440174, 0.0315897, 
    8.147423e-05, 2.925069e-05, 0.0002763608, 0.00169272,
  0.006987884, 0.01037741, 0.000106712, 0.1520645, -8.801387e-07, 
    2.844648e-06, 0.01707571, 4.878036e-06, -0.0001085437, 9.98721e-05, 
    9.762567e-06, 0.0008399441, 0.001009662, 0.000377818, 0.0004087881, 
    0.002519094, 0.002853266, 0.005471938, 0.005736262, 0.002294073, 
    0.005436418, 0.00190411, 0.1518647, 0.0296074, 0.0001252788, 0.001548897, 
    0.003076229, 0.005097186, 0.01942076,
  1.184021e-07, 2.872377e-08, 2.014095e-08, -3.237745e-10, 3.004999e-08, 
    0.0002661387, 0.006915106, 0.000468345, 0.09374934, 0.0001490197, 
    0.001190376, 0.0004772766, 5.064646e-05, 1.108814e-06, 2.086399e-05, 
    4.248319e-05, 0.0003274947, 0.001924813, 0.02688631, 0.05611035, 
    0.006848668, 0.02930532, 0.0001522511, -0.001039213, 7.859947e-05, 
    0.0003802178, 0.004117753, 0.01028379, 1.180466e-07,
  2.862151e-07, -1.201229e-06, 0.0008537637, -1.536576e-06, 7.745622e-08, 
    2.16887e-09, -0.003317599, 0.1830167, 0.2336379, 0.007479284, 0.03229794, 
    0.004470568, 0.002437199, 0.0009089152, 0.001264507, 0.0004960424, 
    0.002788835, 0.01069654, 0.02398504, 0.09520131, -5.490599e-07, 
    0.005392363, 0.004286674, 0.0001743783, 0.0007950867, 0.001183081, 
    0.0009668246, 0.01459756, 0.003445781,
  -0.0003605343, -0.0001214066, -0.0001187548, 0.1702048, -3.559018e-05, 
    1.185427e-08, 0.0004378276, 9.307768e-07, -1.351116e-05, 0.007797398, 
    0.2286177, 0.250878, 0.4412635, 0.4553729, 0.318183, 0.2339541, 
    0.1124435, 0.0829374, 0.07665169, 0.001353564, -4.405111e-05, 
    0.0009321441, 0.0127015, 0.08823719, 0.01958272, 0.01742356, 0.005019893, 
    0.02451807, 0.06392123,
  0.05928189, 0.0235438, 0.01323572, 0.003903629, 0.0001012408, 0.0006132502, 
    0.001424014, 0.1179137, 0.03285502, 0.0185148, 0.03848313, 0.1095983, 
    0.5415937, 0.4925522, 0.5254434, 0.3453323, 0.3139049, 0.1789141, 
    0.1133097, 0.04916872, 0.005043216, 0.001394616, 0.03199289, 0.06148452, 
    0.1563694, 0.35647, 0.2161039, 0.2327407, 0.1421288,
  0.08505931, 0.04903989, 0.0134148, 0.009145653, 0.02801359, 0.01747282, 
    0.0584996, 0.07184506, 0.05052247, 0.06294629, 0.08313367, 0.1961373, 
    0.3882692, 0.2272353, 0.4541849, 0.4534497, 0.158511, 0.2209217, 
    0.09234186, 0.03253162, 0.01594151, 0.07620218, 0.28244, 0.09921295, 
    0.2754927, 0.1745079, 0.1656098, 0.1739686, 0.1584934,
  0.3568857, 0.2274225, 0.1702814, 0.2037468, 0.3244137, 0.4700761, 
    0.1192644, 0.05257645, 0.04119784, 0.07791516, 0.08930013, 0.1678712, 
    0.1735625, 0.3022981, 0.3412845, 0.2943307, 0.1578169, 0.3012725, 
    0.2822816, 0.3147643, 0.1504245, 0.3342206, 0.1237125, 0.2720335, 
    0.3287781, 0.2310552, 0.1523927, 0.2696913, 0.4201473,
  0.494372, 0.3325116, 0.3733929, 0.4736796, 0.4063359, 0.488213, 0.5734901, 
    0.5389142, 0.5584798, 0.5270516, 0.4889741, 0.5153818, 0.4992881, 
    0.4725831, 0.4423166, 0.4649698, 0.467852, 0.4559934, 0.4081459, 
    0.3993465, 0.4209278, 0.2836224, 0.1100766, 0.2550731, 0.2118922, 
    0.1552393, 0.2105795, 0.4164398, 0.4818656,
  0.01659864, 0.01489006, 0.01318148, 0.01147291, 0.009764326, 0.008055747, 
    0.006347168, 0.004423565, 0.005405005, 0.006386446, 0.007367886, 
    0.008349326, 0.009330766, 0.01031221, 0.0133326, 0.0151613, 0.01698999, 
    0.01881869, 0.02064738, 0.02247607, 0.02430477, 0.02402119, 0.02291964, 
    0.02181808, 0.02071653, 0.01961497, 0.01851341, 0.01741186, 0.0179655,
  0.05469336, 0.04078356, 0.01370184, 0.01676823, 0.0123397, 0.08193307, 
    0.0649535, 0.02398636, 0.01273317, 0.01487323, 0.01215826, 0.05555873, 
    0.08411688, 0.003732261, 0.3211586, 0.205086, 0.1839748, 0.2425941, 
    0.1636467, 0.2789591, 0.4940423, 0.5506493, 0.1814796, 0.1069568, 
    0.2841282, 0.4790941, 0.2103533, 0.06718975, 0.07141609,
  0.1839368, 0.1193964, 0.1148402, 0.01932714, 0.02526634, 0.06993914, 
    0.001379131, 0.1074349, 0.2599667, 0.2113623, 0.2601813, 0.2740537, 
    0.05076759, 0.09499212, 0.2929518, 0.2846334, 0.2599905, 0.2796078, 
    0.2274302, 0.3329414, 0.2764637, 0.3141552, 0.2830509, 0.4085752, 
    0.1480495, 0.3267215, 0.3105437, 0.354802, 0.2748878,
  0.271198, 0.2288879, 0.1053295, 0.09697204, 0.07202376, 0.08391006, 
    0.2076671, 0.199755, 0.09905928, 0.05905479, 0.1038161, 0.1566655, 
    0.1311229, 0.1583447, 0.1220649, 0.120092, 0.1227546, 0.1483734, 
    0.1033975, 0.05208494, 0.07361884, 0.06430992, 0.06973557, 0.1136915, 
    0.1484236, 0.3033347, 0.3126843, 0.3549272, 0.3209326,
  0.149278, 0.1622777, 0.1829612, 0.1997313, 0.1774472, 0.1153597, 
    0.08173953, 0.03568043, 0.06139238, 0.07190636, 0.05342432, 0.03814073, 
    0.03066974, 0.02037735, 0.02662032, 0.02719957, 0.01732874, 0.01910167, 
    0.04151675, 0.04995996, 0.06370189, 0.08024794, 0.07372201, 0.1952118, 
    0.02526719, 0.07068818, 0.1245624, 0.1201706, 0.1852129,
  0.03964472, 0.005931291, 0.008216738, 0.009060761, 0.0095772, 0.009714055, 
    0.00790999, 0.01203992, 0.0124898, 0.008211993, 0.006778158, 0.002760396, 
    0.001020634, 0.005135804, 0.119043, 0.008043671, 0.01285193, 0.0352763, 
    0.02007811, 0.03543597, 0.03348102, 0.04526167, 0.02404605, 0.310608, 
    0.005678041, 0.008299306, 0.01785095, 0.01598143, 0.02059308,
  0.004774612, 0.0009075704, 0.01697667, 0.001695566, 0.001103011, 
    0.00173565, 0.004783501, 0.004183452, 0.003831108, 0.0006568088, 
    0.0004045634, -9.578327e-06, 0.01684624, 0.0004739782, 0.001307298, 
    0.003289574, 0.009488982, 0.008167841, 0.01249674, 0.003997426, 
    0.002028474, 0.002150855, 0.00706296, 0.0060499, 0.02078218, 0.003104137, 
    0.001506742, 0.001429864, 0.00199078,
  0.006926459, 0.00792309, -2.197618e-05, 0.001008071, -0.001251754, 
    0.0001979077, 0.0004205591, 0.001900955, 0.001395124, 0.0001924837, 
    1.594836e-10, -3.430364e-07, 0.0004292195, 0.002397749, 0.001542279, 
    0.001483201, 0.001147203, 0.001002175, 0.0006671135, 0.000345497, 
    0.0007715816, 0.002054009, 0.01075496, 0.01788968, 0.004777731, 
    0.05327289, 0.0002032679, 0.0009858636, 0.002365189,
  0.01901726, 0.02078145, 0.0001450907, 0.006287499, 1.473659e-05, 
    0.0002187828, 0.000482655, 0.0005129082, 0.0001614103, -3.144845e-05, 
    0.001981742, 0.0001608071, 0.006106955, 0.000492747, 0.0002099434, 
    9.893728e-05, 0.000115255, 7.381714e-05, 7.334734e-05, 0.0003130047, 
    0.0008411643, 0.004982592, 0.02434153, 0.01101717, -2.428388e-07, 
    1.399993e-08, -0.0002331599, 1.592434e-05, 0.003473952,
  0.009157529, 0.0739775, 0.004140604, 0.0004085147, 2.910341e-05, 
    0.0002465835, 0.0005076379, 0.0002998412, 0.02533481, 0.07641672, 
    0.0006850214, 0.0003572483, 0.0009339903, 0.0007574511, 0.0005838319, 
    0.0001130627, 8.350621e-05, 4.229066e-05, 0.0001179251, 5.812748e-05, 
    0.0004059592, 0.01446026, 0.03544978, 0.05394949, 0.04311571, 
    6.826791e-05, 2.469305e-05, 0.0002270293, 0.001358224,
  0.08132263, 0.009105268, 0.0001908783, 0.1488662, -5.702668e-07, 
    2.175028e-06, 0.02617265, 4.025824e-06, -0.0022327, 8.373428e-05, 
    8.531562e-06, 0.0006608101, 0.0007347374, 0.0002792896, 0.0002637888, 
    0.001526943, 0.001677964, 0.003266672, 0.003484163, 0.001479145, 
    0.003284874, 0.001186367, 0.2023132, 0.04178039, 9.776656e-05, 
    0.000970309, 0.001816878, 0.003304271, 0.04713063,
  1.196629e-07, 2.848706e-08, 1.987702e-08, -3.309145e-10, 3.006095e-08, 
    0.0002027328, 0.003389566, 0.0002298087, 0.1247355, -0.0006573694, 
    0.0007521514, 0.0003078234, 4.101986e-05, 1.187447e-06, 1.743532e-05, 
    3.738721e-05, 0.0002662112, 0.001508557, 0.0191632, 0.04178672, 
    0.005222408, 0.02595001, 0.0001253683, -0.001740486, 5.92092e-05, 
    0.0003075759, 0.003281664, 0.008055734, 1.177452e-07,
  2.844593e-07, -3.473028e-06, 0.0004831856, -1.052105e-06, 7.737454e-08, 
    2.091037e-09, -0.00250877, 0.1754651, 0.2425628, 0.005392119, 0.02385581, 
    0.002429309, 0.001595352, 0.0007251297, 0.0009441144, 0.0003948293, 
    0.002234485, 0.008628018, 0.01920103, 0.08069547, -2.307227e-07, 
    0.03540466, 0.05052494, 0.0001399821, 0.0006497835, 0.0009824383, 
    0.0007814871, 0.01177826, 0.003100573,
  -0.0003328502, -0.0001994079, -0.0003677467, 0.1729158, -3.301576e-05, 
    1.21487e-08, 0.0003111988, 9.161557e-07, -1.101156e-05, 0.005787853, 
    0.2248781, 0.2033057, 0.3389779, 0.3370912, 0.2236053, 0.1842539, 
    0.08036208, 0.05871839, 0.05265179, 0.0008405675, -5.712821e-05, 
    0.0009689445, 0.02021828, 0.06203251, 0.01189011, 0.01047134, 
    0.003245627, 0.0169652, 0.05666757,
  0.05000852, 0.02363943, 0.0170846, 0.002839347, 7.005924e-05, 0.0004426503, 
    0.001056907, 0.1232305, 0.04619617, 0.02368286, 0.09536354, 0.1324212, 
    0.4512988, 0.4112386, 0.4217646, 0.25157, 0.2341279, 0.1308212, 
    0.07857611, 0.04814633, 0.006772056, 0.001050727, 0.04134656, 0.08668251, 
    0.1571084, 0.3098969, 0.1628344, 0.1790009, 0.1015304,
  0.06413408, 0.05147226, 0.01475326, 0.01139261, 0.05328047, 0.05173115, 
    0.08059154, 0.09824641, 0.09226233, 0.09076963, 0.104442, 0.2093709, 
    0.3760817, 0.2034588, 0.3816906, 0.3370676, 0.1639703, 0.2056016, 
    0.09269153, 0.04095707, 0.0254156, 0.08279784, 0.245588, 0.1007312, 
    0.2289591, 0.154285, 0.1325059, 0.1341698, 0.119178,
  0.2819078, 0.1801, 0.1768436, 0.1819965, 0.2956652, 0.5296214, 0.1106133, 
    0.05058873, 0.03948003, 0.07594947, 0.08503001, 0.1610087, 0.1677374, 
    0.3092085, 0.3455245, 0.2599709, 0.1486718, 0.3195153, 0.2668172, 
    0.3280223, 0.1238611, 0.3231358, 0.1014581, 0.2493805, 0.2790931, 
    0.2124365, 0.146931, 0.2330919, 0.3347872,
  0.4325749, 0.3112368, 0.3346589, 0.4158682, 0.349699, 0.4287481, 0.5042844, 
    0.4725358, 0.4894852, 0.4437249, 0.4069052, 0.4336484, 0.419528, 
    0.4011412, 0.372764, 0.3950136, 0.3986776, 0.3922375, 0.3562623, 
    0.345318, 0.3666757, 0.2594659, 0.09981476, 0.2322471, 0.1960595, 
    0.1506246, 0.1966322, 0.3921521, 0.4121178 ;

 average_DT = 730 ;

 average_T1 = 197.5 ;

 average_T2 = 927.5 ;

 climatology_bounds =
  197.5, 927.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
