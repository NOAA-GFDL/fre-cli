netcdf atmos_month.198101-198112.aliq {
dimensions:
	time = UNLIMITED ; // (12 currently)
	pfull = 65 ;
	lat = 2 ;
	lon = 2 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:cell_methods = "time: mean" ;
		aliq:interp_method = "conserve_order2" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19810101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 11 19:59:00 2025" ;
		:hostname = "pp030" ;
		:history = "Tue Sep 23 14:27:36 2025: ncks -d lon,0,1 atmos_month.198101-198112.aliq.nc_lat01 atmos_month.198101-198112.aliq.nc_lat01_lon01\n",
			"Tue Sep 23 14:26:18 2025: ncks -d lat,0,1 atmos_month.198101-198112.aliq.nc atmos_month.198101-198112.aliq.nc_lat01\n",
			"Mon Aug 11 16:17:05 2025: ncks -d lat,,,10 -d lon,,,10 atmos_month.198101-198112.aliq.nc reduced/atmos_month.198101-198112.aliq.nc\n",
			"Mon Aug 11 20:01:59 2025: cdo --history splitname 19810101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/split/regrid-xy/180_288.conserve_order2/19810101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --input_file 19810101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f9d8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run1/share/cycle/19810101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19810101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:NCO = "netCDF Operators version 5.3.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -4.491342e-05, 0,
  0.02296697, 0.02169413,
  0.0009700851, -9.700741e-06,
  0.03809136, 0.03797016,
  0.06700874, -0.002116767,
  0.07488589, 0.07580532,
  0.1655094, 0.03911929,
  0.06676793, 0.06918348,
  0.1666038, 0.09632391,
  0.04636255, 0.05091704,
  0.1564192, 0.1190029,
  0.03815215, 0.04370495,
  0.1479255, 0.1209658,
  0.04313901, 0.04795041,
  0.1471429, 0.1154234,
  0.02838382, 0.03280894,
  0.156526, 0.1384603,
  0.01250187, 0.01664344,
  0.1523077, 0.1374102,
  0.001425399, 0.005074626,
  0.1776326, 0.1497964,
  0.05075943, 0.05286239,
  0.2353781, 0.1482287,
  0.1081508, 0.108836,
  0.3321565, 0.2291835,
  0.1397576, 0.1457741,
  0.3102934, 0.2428513,
  0.2326029, 0.2407883,
  0.2703567, 0.2392209,
  0.2384491, 0.2508228,
  0.2067465, 0.1889161,
  0.2435669, 0.2561018,
  0.1352055, 0.1311978,
  0.1939361, 0.2054376,
  0.09318246, 0.08330628,
  0.1153693, 0.1234577,
  0.07297079, 0.06063513,
  0.07150491, 0.07684118,
  0.07309344, 0.05491544,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.004711038, -0.0001543938,
  0.00256033, 0.001952785,
  0.09316878, 0.003576081,
  0.01556732, 0.01544515,
  0.1029392, 0.0490526,
  0.1294536, 0.1206586,
  0.1116929, 0.1003812,
  0.2422447, 0.2411297,
  0.1337328, 0.1191146,
  0.256148, 0.2574337,
  0.1633203, 0.1435377,
  0.2635781, 0.2676706,
  0.1995254, 0.1901483,
  0.2649513, 0.270602,
  0.2281703, 0.2253346,
  0.2521323, 0.2565313,
  0.2523987, 0.2356615,
  0.2345039, 0.2399323,
  0.275351, 0.2403952,
  0.230301, 0.235682,
  0.3093794, 0.2580776,
  0.254095, 0.2581178,
  0.4140086, 0.3246003,
  0.2995879, 0.3040421,
  0.4318767, 0.4084997,
  0.358198, 0.3646259,
  0.4401007, 0.4582294,
  0.4173191, 0.4248479,
  0.4079661, 0.5115343,
  0.4153857, 0.4225698,
  0.3494994, 0.4846241,
  0.3278913, 0.3377218,
  0.2879099, 0.3980478,
  0.2220206, 0.2291644,
  0.2400485, 0.3074589,
  0.1362991, 0.1385082,
  0.2256765, 0.2887464,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -4.678266e-06, 0,
  0.01948665, 0.01714497,
  -0.001379295, -1.435289e-05,
  0.07102598, 0.06937036,
  0.014405, -0.0001785445,
  0.08739972, 0.08723405,
  0.01928135, 0.007921161,
  0.1346407, 0.1336931,
  0.05033576, 0.02380863,
  0.1739201, 0.1771531,
  0.05990031, 0.06550848,
  0.1799833, 0.1854659,
  0.0734354, 0.1228403,
  0.1714773, 0.1784899,
  0.08743396, 0.1434198,
  0.1606044, 0.1686554,
  0.1164846, 0.1950328,
  0.1634839, 0.1715128,
  0.1344189, 0.2055568,
  0.1690997, 0.1775773,
  0.1294883, 0.2164367,
  0.1861326, 0.1933555,
  0.1323456, 0.2038834,
  0.2259647, 0.2321153,
  0.1449854, 0.2216627,
  0.2810682, 0.2852596,
  0.1853099, 0.2378492,
  0.2707836, 0.2743719,
  0.2587493, 0.2474534,
  0.3068349, 0.3060478,
  0.2940012, 0.2136553,
  0.164152, 0.1618822,
  0.2767366, 0.214793,
  0.08443969, 0.08230194,
  0.2978669, 0.2364064,
  0.08015239, 0.07858247,
  0.2703884, 0.2191936,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -9.199804e-05, 0,
  0, 0,
  0.001440697, 0,
  0, 0,
  0.091052, -0.003702047,
  0.006848796, 0.006259379,
  0.2699322, 0.02864366,
  0.04017341, 0.03704654,
  0.40229, 0.186595,
  0.1169933, 0.1078761,
  0.5538808, 0.3293002,
  0.2205237, 0.2104179,
  0.6179182, 0.4483205,
  0.2861318, 0.281342,
  0.6023822, 0.5506296,
  0.3371134, 0.3364006,
  0.5823221, 0.5602188,
  0.3471834, 0.348908,
  0.5693925, 0.5608546,
  0.3724307, 0.3750005,
  0.5662165, 0.5662276,
  0.400697, 0.4055333,
  0.5854999, 0.590511,
  0.3868661, 0.3872755,
  0.5967954, 0.6180573,
  0.1366692, 0.1245681,
  0.5546175, 0.570996,
  0.04669929, 0.04464187,
  0.4912306, 0.4536555,
  0.04971619, 0.04916412,
  0.4878913, 0.3927369,
  0.04410319, 0.04345647,
  0.4162822, 0.281952,
  0.0358117, 0.03473014,
  0.3148237, 0.2041708,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0001745938, 0,
  0, 0,
  -0.002553057, -6.159259e-05,
  0, 0,
  0.01601959, -0.0001822365,
  8.814842e-05, 5.609445e-05,
  0.04672474, 0.0002231111,
  0.005642292, 0.003587275,
  0.06294678, 0.02191081,
  0.06900441, 0.06432658,
  0.08861378, 0.04432161,
  0.1122268, 0.1080231,
  0.1294441, 0.07652675,
  0.155934, 0.1508025,
  0.1624188, 0.09191135,
  0.1991826, 0.194491,
  0.1594303, 0.1140424,
  0.2526399, 0.2478842,
  0.1593583, 0.1334233,
  0.278973, 0.2743315,
  0.1681137, 0.1527701,
  0.3066899, 0.3023382,
  0.1790444, 0.1725224,
  0.3144235, 0.3095978,
  0.1805746, 0.1941278,
  0.3212804, 0.3160094,
  0.2010247, 0.2315549,
  0.3120373, 0.3075071,
  0.2171474, 0.2365611,
  0.282757, 0.2802002,
  0.2394395, 0.2503728,
  0.2543121, 0.248078,
  0.2536327, 0.2485329,
  0.1638406, 0.1553347,
  0.2580993, 0.2101724,
  0.1325901, 0.124773,
  0.2852113, 0.1308956,
  0.1097378, 0.1046833,
  0.3703603, 0.09421147,
  0.1035665, 0.09938545,
  0.30685, 0.0655206,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0.0001204821, -3.668194e-05,
  0, 0,
  0.0004958096, 0.0005761356,
  0, 0,
  0.02516185, 0.007534817,
  0.001202133, 0.0006541673,
  0.0335715, 0.01821303,
  0.02846045, 0.02513455,
  0.07290995, 0.02468314,
  0.07693093, 0.07670315,
  0.08872149, 0.05468274,
  0.1006265, 0.1005999,
  0.1012162, 0.07676516,
  0.1411746, 0.1400149,
  0.1092212, 0.09070639,
  0.1754344, 0.1767438,
  0.1202212, 0.1171027,
  0.1895771, 0.1931944,
  0.1233328, 0.1466324,
  0.2042726, 0.2089887,
  0.1450891, 0.1761244,
  0.2365253, 0.2409665,
  0.1425191, 0.216225,
  0.2447793, 0.2482699,
  0.121621, 0.2582647,
  0.1370479, 0.1357534,
  0.1399632, 0.2589181,
  0.06687903, 0.06453998,
  0.150223, 0.233447,
  0.01312607, 0.01031134,
  0.1709878, 0.138003,
  0.004821852, 0.004244498,
  0.1662404, 0.07912147,
  0.003101829, 0.003021918,
  0.1139426, 0.06065706,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -4.819941e-05, 0,
  0, 0,
  0.007347177, -0.0001837689,
  0.001665664, 0.0009907245,
  0.04188894, -0.001239319,
  0.02388384, 0.02115944,
  0.04975493, 0.00279889,
  0.0499032, 0.04821989,
  0.07182139, 0.03350017,
  0.08085403, 0.07733684,
  0.1194001, 0.07778943,
  0.1517885, 0.1415054,
  0.1371081, 0.1055079,
  0.3133529, 0.3057201,
  0.1468954, 0.1349598,
  0.3800527, 0.377435,
  0.1548824, 0.1613692,
  0.4115606, 0.4109752,
  0.1654784, 0.1634051,
  0.4590726, 0.4590345,
  0.1793326, 0.1650474,
  0.4964442, 0.497359,
  0.1812605, 0.1707458,
  0.5531421, 0.5556651,
  0.1793602, 0.1831701,
  0.5002319, 0.4986661,
  0.1927524, 0.2122944,
  0.3106402, 0.3028205,
  0.215673, 0.1980826,
  0.1824317, 0.1766734,
  0.21429, 0.1708363,
  0.1078733, 0.1031233,
  0.1589639, 0.122722,
  0.06280475, 0.0592671,
  0.152738, 0.1112433,
  0.02716677, 0.02403313,
  0.09622999, 0.06526627,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -4.035057e-05, 0,
  0, 0,
  -0.0002515528, 0,
  0, 0,
  0.002864336, -5.411986e-05,
  0, 0,
  0.008581975, 0.004736247,
  0.0002160266, 2.046304e-05,
  0.009659011, 0.02200538,
  0.007446679, 0.006876235,
  0.02753555, 0.03381344,
  0.0214645, 0.01854335,
  0.03801402, 0.03988358,
  0.06314979, 0.05838,
  0.05340203, 0.05676458,
  0.1342186, 0.1304251,
  0.0712808, 0.07508865,
  0.1592852, 0.1587761,
  0.07618497, 0.07596207,
  0.1759438, 0.1774538,
  0.08203961, 0.06799297,
  0.1763586, 0.1788832,
  0.08330896, 0.06205471,
  0.1922017, 0.1938577,
  0.09728622, 0.06295542,
  0.1948528, 0.1955874,
  0.151472, 0.05482477,
  0.1568702, 0.156603,
  0.1758619, 0.06834692,
  0.1284978, 0.1314706,
  0.1845847, 0.06501874,
  0.0700592, 0.07063691,
  0.1635979, 0.05191122,
  0.03026015, 0.02723086,
  0.137531, 0.02514263,
  0.01819965, 0.01728851,
  0.06960107, 0.03516091,
  0.0121508, 0.01135126,
  0.05753171, 0.04256249,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0001932691, 0,
  0, 0,
  0.005609978, -0.0002503169,
  0, 0,
  0.0198053, -0.0006658328,
  0, 0,
  0.04101567, 0.007911535,
  0, 0,
  0.0587402, 0.02080031,
  0.001833516, 0.001156008,
  0.07647536, 0.03489848,
  0.005529186, 0.003127942,
  0.1005232, 0.04536717,
  0.03075307, 0.02672863,
  0.1389418, 0.06027723,
  0.07431089, 0.06730748,
  0.1732562, 0.08541671,
  0.13739, 0.1291475,
  0.2023837, 0.1321262,
  0.1638758, 0.155448,
  0.2326793, 0.1633229,
  0.1769939, 0.1683514,
  0.2709692, 0.2048606,
  0.1627824, 0.1533676,
  0.3283429, 0.2398203,
  0.1071833, 0.09966077,
  0.376786, 0.2500581,
  0.03902563, 0.03444779,
  0.3743533, 0.2554266,
  0.0139429, 0.01239912,
  0.3576486, 0.1941382,
  0.003736889, 0.002856296,
  0.3155184, 0.1105515,
  0.003819135, 0.003142179,
  0.1553686, 0.08050427,
  0.003320626, 0.002881413,
  0.1088076, 0.06422083,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.0002600058, 0,
  0, 0,
  -0.00105901, 0,
  0, 0,
  0.02500182, -6.618957e-06,
  0.000794057, 0.0004321011,
  0.02761946, 0.04008167,
  0.02086262, 0.01861147,
  0.06077183, 0.0501748,
  0.05324561, 0.05175487,
  0.09489982, 0.05906706,
  0.06050764, 0.05912954,
  0.1610091, 0.06941463,
  0.1016514, 0.09597941,
  0.2190153, 0.1294457,
  0.1688053, 0.1615343,
  0.3086219, 0.1982387,
  0.2082218, 0.2005184,
  0.3383916, 0.255904,
  0.2529767, 0.2434386,
  0.3649154, 0.3365712,
  0.3260913, 0.3162608,
  0.3782505, 0.393324,
  0.3594762, 0.3494927,
  0.4146209, 0.4263366,
  0.3837712, 0.3730008,
  0.4284412, 0.454033,
  0.4011571, 0.3904168,
  0.4379379, 0.4876425,
  0.3687391, 0.3569036,
  0.4419533, 0.502968,
  0.3176644, 0.307829,
  0.422233, 0.4866165,
  0.2415785, 0.2322704,
  0.3670374, 0.4349916,
  0.1916758, 0.183056,
  0.3217882, 0.3519646,
  0.1450771, 0.1399068,
  0.2666386, 0.2702276,
  0.1148572, 0.1120314,
  0.2275236, 0.1835084,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -1.71803e-05, 0,
  0, 0,
  0.0005680366, 0.0003388887,
  0.005770106, 0.005239251,
  0.001159403, 0.003063783,
  0.01464422, 0.01385491,
  -9.875018e-05, 0.01295865,
  0.02625817, 0.02518668,
  0.008766535, 0.02011747,
  0.06238401, 0.06150869,
  0.02986054, 0.03213101,
  0.1222565, 0.1170061,
  0.02774042, 0.07342289,
  0.1194098, 0.1170025,
  0.02739816, 0.08381601,
  0.1272156, 0.125129,
  0.03114708, 0.08020636,
  0.1474065, 0.1454343,
  0.04245842, 0.07979512,
  0.1521569, 0.1505543,
  0.05448104, 0.07823371,
  0.162397, 0.1620773,
  0.05930302, 0.07474802,
  0.190781, 0.1941935,
  0.04880956, 0.07337786,
  0.2558433, 0.2643838,
  0.0318316, 0.06975681,
  0.4036934, 0.4097953,
  0.02305798, 0.05787795,
  0.5170724, 0.5234949,
  0.01807222, 0.05745756,
  0.5832077, 0.5919046,
  0.01817741, 0.07435265,
  0.5544297, 0.5636647,
  0.02246189, 0.07595833,
  0.404533, 0.4135377,
  0.03188274, 0.06713018,
  0.2443429, 0.2501571,
  0.0532366, 0.06128776,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  0, 0,
  -0.00100424, -1.481948e-08,
  0, 0,
  0.04740304, -0.002822329,
  0.01928804, 0.01793282,
  0.06665791, 0.01341033,
  0.0173764, 0.01779843,
  0.08174979, 0.01748203,
  0.01373157, 0.01418531,
  0.07081497, 0.05544846,
  0.01948795, 0.01999178,
  0.06006323, 0.04815568,
  0.02719259, 0.02769588,
  0.0475177, 0.04383528,
  0.04373394, 0.04407591,
  0.0341759, 0.03787872,
  0.05982209, 0.06071055,
  0.03490298, 0.03459252,
  0.06886089, 0.07022113,
  0.05226711, 0.04197386,
  0.1022699, 0.1038334,
  0.08949219, 0.05606827,
  0.1907186, 0.1937128,
  0.1125208, 0.07677264,
  0.2481331, 0.2487615,
  0.1134536, 0.1115486,
  0.2357024, 0.2390266,
  0.1648434, 0.1219504,
  0.1903012, 0.1965569,
  0.1320664, 0.0900026,
  0.2090821, 0.2139375,
  0.09585206, 0.06167449,
  0.1642161, 0.1686779,
  0.06492731, 0.03827018,
  0.1151061, 0.1179393,
  0.05076362, 0.02477964,
  0.08991197, 0.09149998,
  0.04553084, 0.01698917,
  0.0681904, 0.06946099,
  0.04449594, 0.01249589 ;

 lat = -89.5, -79.5 ;

 lat_bnds =
  -90, -89,
  -80, -79 ;

 lon = 0.625, 13.125 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 746.5, 776, 805.5, 836, 866.5, 897, 927.5, 958.5, 989, 1019.5, 1050, 
    1080.5 ;

 time_bnds =
  731, 762,
  762, 790,
  790, 821,
  821, 851,
  851, 882,
  882, 912,
  912, 943,
  943, 974,
  974, 1004,
  1004, 1035,
  1035, 1065,
  1065, 1096 ;
}
