netcdf atmos.1980-1981.aliq.09 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:22 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.09.nc reduced/atmos.1980-1981.aliq.09.nc\n",
			"Mon Aug 25 14:40:51 2025: cdo -O -s -select,month=9 merged_output.nc monthly_nc_files/all_years.9.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.890948e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -4.942857e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.200513e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.442674e-06, 0, -2.395512e-06, 0, 7.199851e-07, 
    -9.670194e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 7.630036e-05, 0, 0, 0, 9.5472e-06, 0, 0, 0, 0, 0, 0, -4.177581e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.300543e-06, 6.26679e-05, -2.941278e-05, 
    0, 0, 0, 0, 0, 0, -3.65719e-06, 0.0004054295, 0, 1.24653e-05, 0, 0, 
    -4.500419e-06, 0, 0,
  0, 0, 0, 0, 0, 0, -1.991695e-05, 0, -1.479316e-05, 0, 0.000119363, 
    0.0004514212, 0, 0, 0, 0, 0, 0, 0, 0, -7.435316e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.764067e-05, 0, 0, 0, 0, 0, 0, -7.078443e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000198472, 0, 0, 0, 0.001651188, 0, 0, 0, 0, 0, 0, -4.525451e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -4.045842e-06, 0, 0, 0, 0, 0, 0, 0, -3.341342e-06, 0, 0.0001633562, 
    0.0003047668, -6.805423e-05, 0, 0.00164807, -1.658086e-05, 0.0003932315, 
    0, -2.192379e-05, -1.383152e-05, 0.0025475, -4.025054e-05, 1.038925e-05, 
    0.0001207451, 0, -5.624367e-05, 0.0001425201, 0,
  0, 0, 0, 0, 0, 0, 0.001094071, 0, -3.178011e-05, 0, 0.002134509, 
    0.00125673, -1.476104e-05, 0, 0, 0, 0, 0, 0, 0, -8.841633e-05, 
    -4.342038e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.208927e-05, 0, 0, 0, -1.311439e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.131009e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002168997, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.000581336, 0, 0, 0, 0, -7.153341e-07, 0, -3.001078e-07, 
    -2.39399e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0003529919, -1.12767e-05, 0, 0, 0.002887616, -1.076987e-05, 
    0.0009806736, -6.939963e-06, 7.00979e-05, 0, -4.154277e-06, 
    -3.374125e-05, 1.636134e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -3.305467e-05, 5.523111e-05, 1.588287e-05, 0, 0, 0, 0, 0, 0, -2.057306e-05, 
    0, 0.001149393, 0.001355443, 0.0001614362, 0.0007067209, 0.001823427, 
    0.0003386862, 0.0006699085, -1.896761e-05, 0.001278676, 0.001132247, 
    0.005407074, 0.0003245804, 9.875497e-05, 0.0006243605, 0, 0.00146881, 
    0.001241537, 0.0003048564,
  0, 0, 0, 0, 0, 0, 0.003265449, -1.12349e-05, -3.775236e-05, -6.655159e-06, 
    0.005663434, 0.003016175, 0.0003092884, 0, 0, 0, 0, 0, 0, -8.706059e-07, 
    0.0001958079, -0.000257074, 0, 0, 0.000117686, -2.528906e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 6.432066e-05, 0.0008257954, -4.001927e-05, 0, 
    4.394981e-05, -8.289239e-06, 0, -8.907203e-06, 0, 0, 0, 0, 0, 
    -5.51035e-05, 0, 0, 0.0003725305, 0, -3.603805e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007716138, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.209982e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001254156, 0, 0, 0, 0, -1.213253e-05, 0.003674189, 
    0.000671039, 0.0004145988, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0007967941, 0.0001132876, 0, 0, 0.007937665, -3.756663e-05, 
    0.001943952, -4.710382e-05, 0.001181427, 1.726026e-05, -1.909708e-05, 
    -0.0001174802, 3.565564e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.585945e-06, 0, 
    0, 0, 0, 0,
  -4.576025e-05, 0.0003249689, 2.38243e-05, 0, 0, 0, 0, 0, 0.001402969, 
    0.0004031322, 0, 0.004235953, 0.005381284, 0.002664287, 0.002488594, 
    0.006532396, 0.0004521189, 0.001632436, 0.000231619, 0.008419986, 
    0.003250509, 0.01175858, 0.001968866, 0.0001468686, 0.001075797, 
    1.732296e-07, 0.004387385, 0.00354331, 0.0006499298,
  0, 0, 0, 0, 0, 0, 0.008561241, 0.0003816446, 0.001439779, 0.000781487, 
    0.01101498, 0.006729014, 0.002151066, -1.08219e-05, -5.113286e-07, 0, 0, 
    0, 0, -2.119191e-06, 0.0007459613, -0.000413486, -4.399777e-06, 0, 
    0.0006185261, -0.0001290277, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0006368664, 0.001652776, 2.260493e-05, 4.988779e-05, 
    0.0001355347, -4.539149e-05, 1.130682e-05, -3.775871e-05, -8.428137e-06, 
    0, 0, 0, 0, 0.0001207478, 0, 0, 0.001820459, 0, -1.969612e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001387704, 0, 0.005786975, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.505764e-06, 0, -4.3596e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.000137095, -9.636965e-06, -4.114074e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.120534e-05, 0.0002016767, -3.502818e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.456228e-06, 5.90218e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.004218065, 1.716349e-05, 0, 0, -5.819902e-11, 
    0.0001035926, 0.005916753, 0.003076197, 0.001257158, -6.933219e-05, 0, 0, 
    0, 0, 0, 0, 0, 2.277994e-05, 0, 0, 0, 0, 0,
  0, 0.003207975, 0.002596363, 0, 0, 0.01470231, -1.635908e-05, 0.007027639, 
    -0.0001341993, 0.005010516, 0.001734924, -1.254962e-05, -8.896491e-05, 
    4.100033e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005683515, 0, 0, 0, 0, 0,
  -3.21742e-05, 0.0004764144, 6.984735e-05, -2.062521e-06, 0, 0, 0, 
    -1.457836e-05, 0.002116674, 0.001902025, 0, 0.006525875, 0.01162416, 
    0.0066834, 0.003961013, 0.01191254, 0.002182791, 0.00417174, 0.001391533, 
    0.0171184, 0.01077732, 0.0224872, 0.007309983, 0.0002994104, 0.002070919, 
    -9.946823e-06, 0.008739177, 0.005530623, 0.001546079,
  0, 0, 0, 0, 0, 0, 0.01378287, 0.0006371329, 0.002102905, 0.002258431, 
    0.01703449, 0.01243297, 0.006292663, -2.628341e-05, -1.223911e-06, 
    -6.792192e-06, 0, 0, 0, -9.597615e-06, 0.003473328, 0.001693866, 
    -0.0001007395, -1.012966e-05, 0.001840965, -9.88742e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001925956, 0.002409209, 0.0007619994, 0.001213035, 
    0.0004237362, 0.0001751644, 2.104288e-05, -0.0001185004, -4.370063e-05, 
    0, 0, 0, 0, 0.0004207177, 0, -4.379416e-05, 0.00299854, -1.642262e-05, 
    -4.317325e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.205786e-05, -2.637188e-08, 0, 0.003544142, 
    -2.844115e-05, 0.00900941, 0.0002680694, -7.841772e-06, -2.625841e-06, 0, 
    0, 0, 0, -1.394954e-05, 0.0002646688, -1.386154e-05, 0.0001197231, 
    -4.696636e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.609816e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, -1.462074e-05, 3.142185e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -9.624287e-07, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -1.009919e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002933218, 
    0, 0, 0, 0, 0, 0, 0, 0.001546509, 0.001030601, 0.0008475709, 0, 0,
  0, 0, -1.128695e-05, 1.881353e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.019585e-07, 0.001138846, 0, 0, 0, 0, 0, 0, 0, 0, 2.153618e-06, 
    0.0009663118, -0.0001074439, 0.0005889887, 0,
  0, 0, 0, 0, 0, 0, -2.030435e-05, 0, 0, 0, 0, 0, 0, 0, 0, -1.814575e-05, 
    0.001535439, 0, 0, 0, 0, 0, 0, -4.643726e-08, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -9.967535e-06, 0, 0.008872089, 9.267254e-05, -9.309976e-06, 0, 
    -3.271758e-07, 0.0003558941, 0.009427761, 0.008972259, 0.00436852, 
    0.0005419637, 0, 0, 0, 0, 0, 0, 0, 0.0007493261, 2.492209e-05, 0, 0, 0, 0,
  0, 0.01115875, 0.004440827, 0, 0, 0.02067092, -7.154229e-05, 0.01410659, 
    -0.0002574653, 0.01233416, 0.004411678, 0.001189543, 0.0005308524, 
    7.46219e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007621704, 0, 0, 0, 0, 0,
  -7.603e-05, 0.002272513, 0.0004088454, 0.0001948045, 0, 0, 0, 0.0001243061, 
    0.004405111, 0.005593121, -1.086121e-05, 0.009200322, 0.02496331, 
    0.01300529, 0.009667031, 0.02205934, 0.005846417, 0.009344937, 
    0.005036582, 0.02537658, 0.0270225, 0.03828961, 0.01405908, 0.0009743958, 
    0.002480329, 0.0002822427, 0.01161262, 0.01344706, 0.003456126,
  0, 0, 0, 0, 0, -1.788318e-05, 0.01928738, 0.00345634, 0.003303006, 
    0.007917896, 0.02869478, 0.02407573, 0.01376691, -4.419625e-05, 
    -2.344163e-06, 0.0003661429, 0, 0, 0, -4.397242e-05, 0.006835322, 
    0.005830103, -7.799087e-05, -6.464953e-05, 0.003713211, 0.001611072, 
    0.0001648426, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.003361629, 0.002813375, 0.006113529, 0.004118009, 
    0.001720327, 0.004270113, -2.909041e-05, -0.0002621766, 0.000859473, 
    -5.738821e-06, 0, 0, 0, 0.00153321, 4.49115e-05, 0.000170414, 
    0.004342506, 3.408208e-05, 6.587173e-05, 0, 0, 0,
  0, -2.365189e-06, 0, 0, 0, 0, 0, 0, -1.738255e-05, -1.114778e-05, 
    0.0007999849, 0.009812274, 0.002312362, 0.01521851, 0.003077089, 
    0.0003887371, 0.0001873718, 0, 0, 0, 0, 0.0002431315, 0.0006623068, 
    -5.941413e-05, 0.0006164307, 0.0001316329, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003248714, 4.927295e-05, 0.0006835769, 
    -5.872433e-06, 0.001140963, -1.684449e-06, 2.111657e-06, 0, 0, 0, 0, 
    0.0002848544, 0.006799348, 0.0006926818, 0.0008592589, 0.0001342688, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009198954, -5.111194e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0006159814, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0001581275, 0, 0, 0,
  0, 0, 0, 0.001768288, -2.040096e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -4.465261e-07, 0, 0.0007982599, 0, -1.848302e-05, 0.0007611474, 
    -1.081906e-05, 0, 0, 0, 0.001868112, 0.003341355, 0.002823781, 0, 0,
  0, -2.245335e-05, 4.602398e-05, 0.0006054785, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001338734, 7.934551e-05, 0.008478917, 0, 0, 0.0004205397, 0, 0, 0, 0, 
    0, 0.0005873342, 0.008425767, 0.002646676, 0.001891159, 0,
  0, 0, 0, 0, -1.214914e-05, -1.670057e-05, -0.0001369438, 0, 0, 0, 0, 0, 0, 
    0, 2.327165e-06, 0.005372484, 0.004577283, 0.001336929, 0, 0, 0, 0, 
    -4.12362e-06, -9.287453e-08, 0, -2.834468e-05, 0, 0, 0,
  0, -8.32376e-06, -1.070686e-06, 0, -1.93784e-05, 0, 0.01369471, 
    0.002038882, 0.001742469, 0, -3.962718e-05, 0.001623282, 0.0132656, 
    0.02130237, 0.01000574, 0.001342112, -9.662081e-05, 0, 0, 0, 0, 0, 0, 
    0.001433113, 6.619575e-05, 0, 0, 0, 0,
  0, 0.0217995, 0.006351945, 0, 0, 0.02892383, 0.0025352, 0.0291185, 
    0.0006823139, 0.02225261, 0.006651757, 0.01281332, 0.00547921, 
    0.002665264, -2.285879e-06, 0, 0, 0, 0, -8.211713e-10, 0, -1.487604e-06, 
    -1.713855e-05, 0.001594631, -4.156341e-06, 0, 0, -3.703644e-06, 
    -1.222183e-05,
  0.001108801, 0.005368973, 0.0008192896, 0.0008718347, 0, 1.825793e-08, 0, 
    0.000173135, 0.007515171, 0.01523523, 0.0002932252, 0.01624596, 
    0.04461482, 0.0292635, 0.02536419, 0.037671, 0.01369348, 0.01588837, 
    0.007327657, 0.04539867, 0.06036917, 0.0802377, 0.02183079, 0.002162467, 
    0.005172146, 0.002371438, 0.01609587, 0.031271, 0.005580007,
  0, 0, 0, 0, -3.937858e-07, -6.453497e-05, 0.02596847, 0.008144604, 
    0.007352162, 0.01270157, 0.04126269, 0.04440503, 0.02825567, 
    6.984419e-05, 0.0001880158, 0.0009666664, 0, 0, 0, -8.023914e-05, 
    0.01471666, 0.01469075, 0.001040342, 0.0003988144, 0.006734042, 
    0.00533999, 0.0008152519, 0, 0,
  0, 0, 0, 0, 0, 0, -7.150439e-12, 0.006186493, 0.005069556, 0.01240065, 
    0.01177282, 0.007329386, 0.01043162, 0.003547668, -0.0002409978, 
    0.003704099, 0.0001780052, 0, 0, 0, 0.002196583, 0.003146436, 
    0.002293618, 0.007391956, 7.826614e-05, 0.0008914717, 0.0001227673, 0, 0,
  -2.411498e-05, 0.000277357, 0, 0, 0, 0, -2.219067e-06, 0, -1.736534e-05, 
    0.0003925178, 0.003559012, 0.02411587, 0.009498915, 0.02285479, 
    0.006316751, 0.00330251, 0.0003908321, 3.997358e-07, 0, 0, 0, 
    0.002378383, 0.007940529, 0.002276784, 0.002949468, 0.01396121, 
    0.000538107, 0, 0,
  0, -2.391212e-06, 0, -4.805449e-05, 0, 0, 0, 0, 0, 0, 0.0009025702, 
    0.00195332, 0.003845128, 0.002941801, 0.003124913, 0.004389107, 
    0.0005712763, 0.0009741351, 0, 0, 4.657147e-05, 0.0009590364, 
    0.002532032, 0.01425502, 0.003831849, 0.003092474, 0.002319116, 
    -1.584067e-05, 0,
  -5.076517e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.200081e-06, 
    0.001606952, 0, 0, 0, 0, 0, 0, 0.002017934, 2.426327e-05, 0.001213379, 
    -3.737661e-05, 0, 0, 6.015331e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, -8.97581e-06, 0, -1.061751e-05, 0.002166917, 0.0005532616, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001435771, 0, 0, 0, 0, 0, 0.0006585616, 0, 
    0, 0,
  0, 0, 0, 0.003874587, 0.000451011, 0, -9.95518e-07, 0, 0, 0, 0, 0, 0, 0, 
    0.001617217, 0, 0.003595042, 6.41039e-06, 0.001700204, 0.002260302, 
    0.001580753, 0, 0, 0, 0.002391716, 0.008774817, 0.009136036, 
    8.612038e-05, -1.909914e-05,
  0, -5.460265e-05, 0.0003747614, 0.002199988, 0, -9.454212e-07, 0, 0, 0, 0, 
    0, 1.194307e-07, 0, 0.002284358, 0.00885186, 0.02236322, 0.0009401366, 
    3.108504e-05, 0.004469174, 0.002511116, 6.821091e-05, -1.014207e-06, 0, 
    0, 0.001967807, 0.02123229, 0.01083475, 0.002812545, 8.585925e-06,
  0, -1.109702e-10, 3.062098e-05, 2.978952e-09, 2.961232e-05, 5.338198e-05, 
    -9.882458e-05, 1.999973e-08, 0, 0, 0, 0, 0.0003472559, -1.5276e-09, 
    0.007534576, 0.01909912, 0.009400794, 0.003550747, -7.475509e-05, 0, 
    -6.793532e-09, 0, -6.036836e-07, -1.043826e-06, 0.0001534855, 
    0.000248378, -5.133587e-07, 0, 0,
  0, -1.033389e-05, 2.135306e-05, -3.286738e-07, -2.648131e-05, 0, 
    0.02392091, 0.006747292, 0.003603998, 0, 0.0007488584, 0.008949857, 
    0.02083653, 0.04433241, 0.02636291, 0.004133576, -0.0001077714, 0, 0, 0, 
    0, 0, -3.301235e-10, 0.004735761, 0.0007287182, 0, 0, 0, 0,
  1.508587e-06, 0.04108162, 0.01218089, 1.361442e-08, -9.443388e-07, 
    0.04259498, 0.01474165, 0.05815049, 0.008367551, 0.03997804, 0.01064865, 
    0.03353941, 0.02151142, 0.01144545, 5.505063e-06, 0.0002255841, 0, 0, 0, 
    -5.006563e-06, 9.69792e-07, 0.0005041242, 0.0009517123, 0.01161666, 
    -1.348111e-05, -7.974765e-06, 0, -1.140051e-05, -1.803274e-05,
  0.009873477, 0.01163421, 0.004960547, 0.001344895, 0, 3.730099e-05, 
    0.000754517, 0.008316975, 0.01976266, 0.03855341, 0.002079746, 
    0.03216207, 0.08152413, 0.06209296, 0.04557923, 0.05945538, 0.02209977, 
    0.02202459, 0.01081256, 0.06970298, 0.1053471, 0.1444385, 0.04668429, 
    0.01286311, 0.01216066, 0.007577863, 0.03112428, 0.04628551, 0.01296923,
  0, 0, 0.0001876917, 0, -4.082655e-05, 0.0007893622, 0.03813424, 0.02800473, 
    0.02340839, 0.0239446, 0.05617009, 0.06513496, 0.05459892, 0.002033497, 
    0.002069448, 0.001415671, 0.001307558, -1.868567e-08, 0, 0.0002064141, 
    0.03274233, 0.04857852, 0.004267905, 0.002795144, 0.007146718, 
    0.01428226, 0.001603433, 0, 0,
  0, 0, 0, 0, 0, 0, -8.092076e-06, 0.01282414, 0.009345516, 0.01620899, 
    0.02321533, 0.01651718, 0.01930121, 0.01385587, 0.0009119636, 
    0.008270074, 0.000764099, -4.596731e-08, 0, 0, 0.007008221, 0.01059102, 
    0.01557227, 0.0113768, 0.005531813, 0.006227378, 0.00174114, 0, 
    -2.879863e-06,
  3.127315e-06, 0.001477898, -1.738543e-05, -1.701393e-11, 6.01638e-13, 0, 
    -3.527728e-05, -1.484806e-08, 2.498048e-05, 0.00340783, 0.01040805, 
    0.04702411, 0.02229274, 0.03543206, 0.01259153, 0.01236271, 0.0040106, 
    -9.933357e-06, 0, 0, 7.901056e-05, 0.003639051, 0.0154471, 0.006458249, 
    0.008896182, 0.0346618, 0.0009869426, -2.419284e-05, -3.28137e-06,
  -6.052896e-06, 0.0006043371, 0, 0.0005593611, -8.309371e-08, -3.562315e-05, 
    0, 0, 0, 0.0004392108, 0.006898359, 0.004427579, 0.008991363, 0.01057302, 
    0.005658254, 0.008014087, 0.003454466, 0.004681389, -8.410365e-11, 0, 
    0.0004281729, 0.001491864, 0.007887877, 0.02361027, 0.01634093, 
    0.007006047, 0.01124977, 0.002578838, -7.75579e-05,
  4.762156e-05, -5.821549e-07, -9.124633e-06, -9.871915e-06, 0.002113841, 
    0.0006296516, 0, 0, 0, 0, -3.930118e-05, 0, 0, 3.26384e-05, 0.003114721, 
    0.003330511, 0.0007211685, 0, 0.0004869913, -4.308236e-11, -6.177888e-10, 
    -9.884006e-11, 0.002060788, 0.003073859, 0.004811421, 0.001076743, 
    -2.519043e-05, -1.290625e-05, 0.0007022558,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009695442, -3.800468e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.065963e-09, 
    0, 0, 0, 0, 0, 0, 0, 0,
  -2.572303e-05, 0.0004362886, -1.701548e-05, -2.073045e-05, 0.0005823618, 
    0.004464213, 0.002104528, 0.0002668727, 0, 0, 0, 0, 0, -1.813419e-06, 
    -3.48035e-06, 0, 0, -2.235084e-06, -7.819501e-06, 0.001704837, 
    0.0001439164, 0.0002975532, 1.183421e-07, 0, 0, 0.00192107, 0, 
    6.627991e-05, -6.16228e-07,
  -4.517406e-06, -0.000106122, 2.012114e-06, 0.00638152, 0.001603174, 
    0.004437178, 0.001756414, -3.311404e-06, 0, 0, 0, 0.0008950271, 
    0.0003183396, -2.814946e-05, 0.002601183, 0, 0.006805505, 0.003543174, 
    0.006138313, 0.01254911, 0.007183665, 0.0001915175, 0.0002618099, 
    0.000227483, 0.004744397, 0.01415681, 0.02312423, 0.002793102, 0.005254095,
  3.428947e-05, 0.0005606847, 0.0007140075, 0.004476387, 0, 1.62121e-05, 0, 
    2.620322e-09, 2.79652e-08, -1.925895e-08, -1.275509e-10, 0.0002390479, 0, 
    0.003712632, 0.01931235, 0.04186612, 0.006419219, 0.006399672, 
    0.03013668, 0.00367869, 0.0004158457, 0.001265661, 1.590657e-05, 
    -4.272238e-08, 0.005529297, 0.03718016, 0.02103684, 0.004623499, 
    1.693316e-05,
  0, 6.298968e-06, 0.004731199, 2.738798e-07, 0.0006885469, 0.002019764, 
    0.0003494494, 0.0001642091, 1.008576e-06, 1.364713e-06, 3.324194e-07, 
    1.507119e-07, 0.00603752, 1.525892e-05, 0.01550084, 0.05054583, 
    0.02862025, 0.01677933, 0.0015878, -4.239075e-06, 5.573242e-06, 
    2.313051e-07, 2.971562e-06, 0.0003118939, 0.000634774, 0.002656522, 
    5.995405e-05, 1.394784e-07, -2.112104e-07,
  -1.09209e-08, -1.449568e-05, 0.0001449308, 0.0001007782, 9.851811e-06, 
    8.571333e-07, 0.0328031, 0.04433942, 0.007464611, -1.102894e-05, 
    0.01029174, 0.05710056, 0.07645257, 0.1513529, 0.1135114, 0.03000866, 
    0.0007002041, -8.80626e-07, 1.41451e-07, 7.953906e-06, 9.654703e-05, 
    2.733113e-05, 6.931133e-05, 0.01675876, 0.01202877, 3.704137e-05, 
    -1.339647e-05, -7.685646e-09, 0,
  0.004453319, 0.09160927, 0.03861441, 0.0001313759, -8.505329e-06, 
    0.06235743, 0.03336569, 0.1664807, 0.07077584, 0.08065508, 0.05577544, 
    0.1129976, 0.09332235, 0.06287925, 0.002983977, 0.0002390232, 
    0.000189174, 8.182915e-08, -5.101762e-07, 3.98485e-05, 0.007709589, 
    0.00322731, 0.01453854, 0.08372481, 0.001885725, 2.891942e-05, 
    -8.947833e-08, 0.003001111, 4.963172e-05,
  0.04982138, 0.03548205, 0.02307862, 0.001615467, -1.154428e-06, 
    0.002171023, 0.02924514, 0.3596317, 0.418376, 0.3897806, 0.2530107, 
    0.2858467, 0.2713496, 0.2187322, 0.1561057, 0.1286132, 0.04575422, 
    0.02412446, 0.01664578, 0.1186038, 0.2982286, 0.3561081, 0.08526489, 
    0.06521927, 0.0323801, 0.01598238, 0.06334908, 0.07722548, 0.02996064,
  7.918973e-05, -5.404649e-05, 0.0008242139, 0.0002221104, 0.003941667, 
    0.05607595, 0.2786134, 0.1441351, 0.1950109, 0.08421706, 0.1355553, 
    0.1998219, 0.1789856, 0.03904531, 0.00821011, 0.004395347, 0.005730255, 
    0.001099876, 2.505498e-06, 0.02481995, 0.1505807, 0.1600378, 0.05908523, 
    0.06290947, 0.01006503, 0.02239452, 0.01091221, 0.002093685, 0.001428216,
  -4.232181e-06, -1.533275e-09, 0, 5.396137e-10, 3.478066e-08, -8.163291e-07, 
    7.255236e-05, 0.01916813, 0.01539935, 0.07239117, 0.08620033, 0.07061912, 
    0.09169368, 0.1046423, 0.02666874, 0.01964514, 0.01291779, -1.477242e-05, 
    4.370815e-10, -5.605702e-08, 0.0254594, 0.0661118, 0.06321127, 
    0.02441999, 0.01320865, 0.02422599, 0.004043276, 9.865355e-06, 
    0.0002584409,
  0.000472493, 0.0045586, 0.0004032286, -6.40696e-10, -1.3156e-06, 
    8.965784e-06, -3.036975e-05, 0.0006828935, 0.002387304, 0.009189141, 
    0.03038035, 0.08760544, 0.06913434, 0.07980603, 0.04165563, 0.03598223, 
    0.01331298, 0.0005017563, 0.0002549562, 0, 0.0006260502, 0.005330867, 
    0.02745959, 0.01513978, 0.01529982, 0.04451859, 0.002588695, 
    -3.309475e-05, 0.0003124301,
  3.720825e-05, 0.00390201, 0.0009336676, 0.002300692, -4.605463e-05, 
    -1.303926e-05, 0, 0, -7.109527e-05, 0.003762956, 0.01391062, 0.01181077, 
    0.02743703, 0.02538268, 0.01517816, 0.01430907, 0.01903615, 0.01008797, 
    0.0002096475, 0, 0.001697345, 0.004411076, 0.01700957, 0.0304339, 
    0.02994545, 0.01974029, 0.04036088, 0.01214835, 0.00270002,
  0.003321539, -5.470845e-05, 0.003699178, 0.0002944916, 0.004488586, 
    0.001180692, 0, 0, 0, 0, -0.0001133223, -7.174458e-06, 0, 0.002249302, 
    0.006962833, 0.006204387, 0.004873302, 9.083585e-05, 0.002477174, 
    0.0002402755, -2.140125e-10, -6.950869e-05, 0.002348467, 0.004113985, 
    0.01621325, 0.008992009, 0.000819894, 0.0006690708, 0.005177666,
  0, 2.363701e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.562505e-05, 
    6.146011e-06, 0, 0, 0, 0, 0, 0, 0, -8.999094e-06, 0.003308674, 
    -1.651533e-05, 0, 0.0001779001, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.286617e-06, 0, 0, -1.075817e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.736596e-06, 0, 0, 0, 0.001399997, 0, 0, 0, 0,
  0.000692127, 0.002176247, 6.440295e-06, -0.0001838397, 0.004640635, 
    0.008365745, 0.004319167, 0.0006383971, 0, 0, 0, 0, 0, 0.0007438203, 
    0.0001772134, 2.410374e-05, 0, -3.484606e-06, -0.000117513, 0.004119703, 
    0.0012678, 0.002624018, 0.004122166, 0.0003277751, 5.427812e-05, 
    0.005150575, -4.459916e-07, 0.001210956, 3.678952e-05,
  0.0002683816, 0.001314957, 0.001933835, 0.009839475, 0.009205398, 
    0.01048181, 0.004684286, -2.184722e-05, 3.760872e-08, -1.075884e-08, 
    -2.083013e-07, 0.002906721, 0.004447996, 0.003500924, 0.004727295, 
    0.0007161088, 0.008937062, 0.01147069, 0.01417218, 0.02849005, 
    0.01921787, 0.003736325, 0.003018772, 0.001945499, 0.008130534, 
    0.02276714, 0.03588716, 0.01217857, 0.01999038,
  0.0003905048, 0.001531109, 0.001999132, 0.009881185, 0.0001841655, 
    0.00123595, 2.834363e-08, 3.418001e-07, 0.0002475031, -1.16492e-05, 
    5.894481e-08, 0.0008766324, -3.298836e-06, 0.005101994, 0.03787221, 
    0.06442177, 0.03375065, 0.02933997, 0.07272174, 0.02059578, 0.006130055, 
    0.008420336, 0.004213098, 0.001035463, 0.01583634, 0.08396518, 0.0558025, 
    0.02619347, 0.001429849,
  2.194243e-06, 0.0001533416, 0.009112344, 0.0001014616, 0.006175471, 
    0.007934654, 0.003570031, 0.001885612, 6.394551e-06, 1.423052e-06, 
    3.72001e-07, 5.558749e-07, 0.01622756, 0.00134056, 0.03734666, 0.1038161, 
    0.0893594, 0.06424949, 0.0123972, 0.001298701, 5.086985e-06, 
    7.299658e-06, 1.483394e-05, 0.03229476, 0.1157205, 0.01903526, 
    0.002773936, 0.0001507844, 0.004720461,
  5.861423e-06, -0.0004310943, 0.01796374, 0.003956061, 0.0001333691, 
    0.009079427, 0.06358478, 0.09670699, 0.01486465, 8.880467e-05, 
    0.01568265, 0.04929257, 0.06929433, 0.1544722, 0.1493729, 0.09344795, 
    0.01476653, -1.80888e-06, 2.49127e-06, 6.824981e-05, 0.007036715, 
    0.0002865909, 0.000547834, 0.1412219, 0.1978158, 0.002052451, 
    0.000109968, 4.685893e-05, 1.723331e-05,
  0.08221238, 0.4420458, 0.4185854, 0.006401857, 0.0002950415, 0.1336188, 
    0.1651622, 0.3304788, 0.3179869, 0.2498091, 0.07856417, 0.1105061, 
    0.08582318, 0.06058647, 0.002035816, 0.001539045, 0.0002045276, 
    1.690205e-05, 3.034389e-05, 0.02193896, 0.05952459, 0.08190501, 
    0.08528274, 0.2550744, 0.04365836, 0.00147861, 0.001301604, 0.02982118, 
    0.01716107,
  0.2231912, 0.174384, 0.175843, 0.003318752, 0.001871987, 0.005433955, 
    0.08293208, 0.3076586, 0.3539612, 0.2742016, 0.1500449, 0.2354721, 
    0.2457371, 0.2064234, 0.1643228, 0.1721873, 0.09863613, 0.02959871, 
    0.01786901, 0.1522344, 0.3540224, 0.3939888, 0.2261969, 0.1884006, 
    0.08176054, 0.05315562, 0.1222848, 0.1777081, 0.1897784,
  0.01402703, 0.01549249, 0.01519739, 6.348114e-05, 0.002087247, 0.04046558, 
    0.2677094, 0.09167865, 0.1708968, 0.06580669, 0.1129248, 0.1461324, 
    0.1538034, 0.0782207, 0.09678829, 0.08030218, 0.05643497, 0.008909679, 
    5.961101e-06, 0.01494883, 0.1083257, 0.1686892, 0.08142343, 0.1328888, 
    0.09071814, 0.07976773, 0.05370439, 0.07314494, 0.07381409,
  0.0003635712, 0.003663002, 0.0001008507, 0.0005301854, -1.009277e-08, 
    -1.777477e-07, 0.0004433529, 0.02755022, 0.02871227, 0.06825001, 
    0.07109444, 0.06270292, 0.1020548, 0.1214778, 0.08597702, 0.07946663, 
    0.07644136, 0.05064287, 3.233798e-05, 5.017583e-06, 0.1045391, 0.1425683, 
    0.1849887, 0.1296316, 0.1063064, 0.1053794, 0.03723283, 0.03604241, 
    0.002233235,
  0.001097755, 0.0104239, 0.001331561, -1.524086e-06, 0.0003827666, 
    0.001016691, 0.0004024027, 0.01083857, 0.01921166, 0.04853494, 0.1002168, 
    0.1964317, 0.1835305, 0.2095793, 0.1639192, 0.1767578, 0.04072536, 
    0.0368404, 0.01687399, 0.0004104497, 0.001495216, 0.04175297, 0.1013984, 
    0.06282891, 0.1006301, 0.1091256, 0.04372123, 0.007793638, 0.009049784,
  0.00189325, 0.01619142, 0.002178099, 0.006387671, 0.001956362, 0.00388199, 
    -1.082876e-06, 0.0005123903, 4.611436e-05, 0.005865905, 0.02377338, 
    0.0218134, 0.0604732, 0.08292977, 0.04563885, 0.03794529, 0.07051495, 
    0.02838972, 0.01349731, 0.0002125748, 0.00432342, 0.00923224, 0.02630876, 
    0.04295028, 0.05756754, 0.05722316, 0.1002941, 0.03201256, 0.005130492,
  0.01458458, 0.001491625, 0.008253303, 0.002541049, 0.006404892, 
    0.001197739, -6.731482e-05, -2.638197e-06, 0.0003122162, -1.039032e-05, 
    0.0009852281, 0.0005965616, -5.233475e-05, 0.004562809, 0.01320141, 
    0.02431479, 0.01087207, 0.004580798, 0.005746569, 0.001702887, 
    0.0004481284, 0.0004770586, 0.00244167, 0.00661731, 0.03327664, 
    0.02980196, 0.01014275, 0.006786376, 0.01214173,
  -2.407863e-05, 0.001568744, 7.012323e-05, 0.0008113873, 0, 0, 
    -1.032797e-05, 0, 0, 0, 0, 0, 0, 0, -7.699627e-05, 0.0003884753, 
    0.001312449, 0.0002704604, -1.154822e-05, -4.409435e-07, 0, 0, 0, 
    -1.567588e-05, 0.006554468, 4.770537e-05, 7.748682e-06, 0.002842247, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.484175e-06, 
    3.119195e-05, 0, 0, 0, 0, -1.129514e-05, -3.454579e-08, 0, 0, 
    -6.933297e-14, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00062775, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0003380186, -7.033306e-06, 5.641097e-05, -1.115837e-06, 0, 0, 
    -3.919375e-06, -5.178449e-05, -2.944129e-05, 0.0004639687, -2.196272e-05, 
    -6.837006e-08, -1.092506e-05, 0, 0, 0, 0.0007235869, 0, 1.045488e-05, 0, 
    0.002032917, -3.461899e-05, 0, 0, 0,
  0.003941321, 0.007414282, 0.0002093284, 0.003500848, 0.01125752, 
    0.01669279, 0.008427877, 0.00198069, 0.0001535967, 0.0007680577, 
    0.0009330139, 9.107891e-05, 1.484897e-07, 0.00462669, 0.004649783, 
    0.001344194, -6.226192e-06, 0.0003653975, 0.00240863, 0.01272514, 
    0.01108637, 0.008875009, 0.008446151, 0.003441487, 0.002550686, 
    0.005467977, -2.921078e-05, 0.007855125, 0.00476354,
  0.02834737, 0.02386586, 0.01609094, 0.02710455, 0.02477537, 0.03862889, 
    0.01476704, 0.0001054832, 2.195983e-05, -1.590245e-05, 0.0001943722, 
    0.007424492, 0.00798545, 0.01208435, 0.01237007, 0.002239035, 0.01452186, 
    0.02369606, 0.03103996, 0.04206904, 0.05377949, 0.0299224, 0.01288796, 
    0.008346652, 0.01346692, 0.04270434, 0.0900572, 0.04907859, 0.05346262,
  0.0345564, 0.02750031, 0.005969771, 0.05337053, 0.02160338, 0.006507008, 
    0.002228573, -2.288556e-05, 0.01099869, 0.004073096, 0.005326081, 
    0.00917554, 0.006589704, 0.007691731, 0.04796933, 0.103985, 0.102847, 
    0.1047125, 0.175771, 0.1027038, 0.02491785, 0.01492118, 0.01762531, 
    0.01178455, 0.03523385, 0.1274407, 0.1144566, 0.09020159, 0.03833282,
  5.474719e-07, 0.002504649, 0.05660294, 0.0109836, 0.01336163, 0.007812624, 
    0.001616197, 0.00271159, 4.968551e-06, 8.77458e-07, 2.017191e-07, 
    5.38687e-08, 0.01213581, 0.0001654027, 0.04050533, 0.1019476, 0.08661698, 
    0.07542592, 0.007728597, 0.0007497623, 2.097989e-06, 2.274629e-06, 
    2.974856e-06, 0.03299641, 0.0972409, 0.08204639, 0.0001436935, 
    0.001503608, 0.0004402277,
  2.309607e-06, -0.0001259751, 0.01429074, 0.0005505349, 0.0007176696, 
    0.005425254, 0.03946623, 0.07315753, 0.01140226, 0.0001093941, 
    0.01260396, 0.03301184, 0.05842841, 0.1266149, 0.1097355, 0.0663554, 
    0.01042124, 2.658729e-06, 8.217265e-08, 2.481196e-06, 6.249318e-05, 
    1.769883e-05, 8.085009e-06, 0.1094807, 0.1394639, 4.041742e-05, 
    1.171257e-05, 3.228691e-06, 5.359978e-07,
  0.02830475, 0.4037915, 0.315528, 0.001897844, 3.517133e-06, 0.1104039, 
    0.110342, 0.2660657, 0.2482888, 0.1970868, 0.05560782, 0.09425892, 
    0.05713639, 0.04646517, 0.001026735, 0.0003159754, 2.436767e-05, 
    3.02729e-06, 9.403e-06, 0.005521677, 0.01701265, 0.02825779, 0.06665082, 
    0.1969332, 0.01623894, 0.001217365, 0.0001315397, 0.009395925, 0.003826078,
  0.1848066, 0.1412087, 0.1218017, 0.03073549, 0.0006654801, 0.002584956, 
    0.04772633, 0.2099333, 0.2648616, 0.171959, 0.08959877, 0.1747572, 
    0.1984193, 0.177983, 0.1370729, 0.1459343, 0.07345114, 0.0243086, 
    0.01613928, 0.1132097, 0.2754105, 0.3657511, 0.2005909, 0.1350192, 
    0.05612336, 0.03352504, 0.08650903, 0.1510188, 0.1402037,
  0.009100021, 0.01122434, 0.007886615, 8.999238e-05, 0.004761101, 
    0.03303385, 0.2434317, 0.08299557, 0.1244366, 0.061191, 0.1038209, 
    0.1248579, 0.1284021, 0.04385491, 0.05388984, 0.06736505, 0.04459167, 
    0.005162699, 1.705509e-06, 0.01541845, 0.08090271, 0.1326718, 0.05820045, 
    0.1091212, 0.06475902, 0.06019751, 0.04470792, 0.07782821, 0.0923593,
  0.07924399, 0.03536113, 5.76881e-05, 0.0001323192, -1.60556e-07, 
    -2.728441e-08, 0.0004159935, 0.0357337, 0.06654844, 0.07036609, 
    0.0618313, 0.05404379, 0.09641925, 0.08804053, 0.05729778, 0.06804985, 
    0.07721224, 0.05764378, 0.01108981, 2.268486e-06, 0.1020298, 0.1084744, 
    0.1485932, 0.09959914, 0.09418944, 0.07754779, 0.06449575, 0.05289105, 
    0.04125429,
  0.06255765, 0.06275021, 0.01233345, 0.0002509301, 0.004485843, 0.01372982, 
    0.002626213, 0.02995879, 0.05945976, 0.07488218, 0.1594819, 0.1977375, 
    0.1984531, 0.1837344, 0.1591622, 0.2320928, 0.1199187, 0.1371463, 
    0.06093162, 0.009773762, 0.02589722, 0.1000174, 0.1236418, 0.09852426, 
    0.1253168, 0.1477752, 0.09400325, 0.06285444, 0.07360178,
  0.03924175, 0.03083539, 0.0306426, 0.0182489, 0.01725762, 0.008270673, 
    0.001701717, 0.001514046, 0.001050442, 0.01518475, 0.04407778, 
    0.03875344, 0.07245541, 0.1402444, 0.07745461, 0.09354413, 0.1441721, 
    0.1291864, 0.1005396, 0.01594732, 0.01746015, 0.05469716, 0.04783292, 
    0.07731087, 0.1198574, 0.1451886, 0.1864088, 0.1156853, 0.06403343,
  0.04506896, 0.01155874, 0.01240889, 0.008492383, 0.009532674, 0.003425913, 
    0.00095457, 0.0005543588, 0.002752585, 0.0006819479, 0.007653522, 
    0.001856824, 0.0001632517, 0.04128325, 0.0219115, 0.02086024, 0.03065157, 
    0.02085734, 0.01369713, 0.01109536, 0.008693877, 0.01167784, 0.003172928, 
    0.01957108, 0.050317, 0.04711196, 0.05316892, 0.01493928, 0.03688025,
  0.001704775, 0.006543613, 0.0002168734, 0.002507197, 0.0001323354, 
    -1.741072e-07, 0.002672473, 0, 0, -3.818434e-06, 2.970869e-05, 
    -1.993629e-05, 0, 0, 0.0007788358, 0.00588805, 0.01158104, 0.01536862, 
    0.009943199, 0.01312167, 0.004647734, 2.867659e-05, 9.935944e-07, 
    -0.0001283525, 0.01390963, 0.0004252963, 0.001428448, 0.01555833, 
    0.009253046,
  0, 0, -5.465908e-08, 0, -1.279808e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.743708e-05, -4.383576e-05, -2.23684e-05, 0.0004982221, 1.424199e-07, 
    1.729498e-06, 7.628089e-05, -1.545367e-07, -1.842116e-05, -0.0001147612, 
    1.000034e-05, -1.58397e-10, -2.516723e-05, 1.454719e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003492455, 0, 0, 0, 0,
  0, -9.119271e-06, -4.061323e-06, 0, 0.001041075, 4.663298e-05, 
    -8.927095e-05, -1.277286e-05, 0.0001947757, 0, -1.219264e-05, 
    -0.00015313, 0.0006760309, 0.001145128, 0.0003130976, 0.0001516447, 
    4.806752e-05, 0, 0.0003324146, 0.001545974, 0.003916014, 0.001553762, 
    0.001043864, 7.200222e-06, 0.002462114, 0.001490619, -6.286884e-06, 
    0.0005255134, 0,
  0.01526213, 0.035595, 0.01063785, 0.03460615, 0.05932593, 0.0554723, 
    0.03622633, 0.01821184, 0.005257154, 0.003928144, 0.00271347, 
    0.0005988176, 0.002624143, 0.0135819, 0.0112817, 0.005096164, 
    0.001015534, 0.004979125, 0.009145747, 0.02470387, 0.03085918, 
    0.02401944, 0.02760924, 0.01799719, 0.02784652, 0.01354033, 0.003298396, 
    0.01779342, 0.02358685,
  0.0953467, 0.07098947, 0.1075502, 0.1313155, 0.1770668, 0.1158404, 
    0.06647612, 0.03542699, 0.02119149, 0.01109558, 0.007158981, 0.02018914, 
    0.02843045, 0.05164206, 0.03210387, 0.04103858, 0.04100688, 0.04763193, 
    0.05465887, 0.07325047, 0.1259932, 0.08602323, 0.0715568, 0.02663798, 
    0.06808761, 0.08120624, 0.1335973, 0.08845171, 0.1234912,
  0.04583514, 0.02216552, 0.0539795, 0.07652301, 0.02305882, 0.008055667, 
    0.0001872726, -0.0001232111, 0.01150155, 0.00502244, 0.00583264, 
    0.0103489, 0.006398342, 0.01603451, 0.06028786, 0.1177705, 0.1080003, 
    0.1359442, 0.2285103, 0.1276065, 0.0280376, 0.03483994, 0.03562856, 
    0.02530881, 0.05084881, 0.1179416, 0.1018192, 0.07634009, 0.05220214,
  3.973359e-07, 0.004125102, 0.07533513, 0.007653493, 0.01465307, 
    0.007751067, 0.0001903521, 0.008347655, 1.627373e-06, 4.821773e-07, 
    1.616454e-07, -3.33594e-07, 0.005780566, 0.002993798, 0.04771814, 
    0.09620225, 0.07329594, 0.06239852, 0.003332827, 9.465079e-06, 
    2.404901e-07, 6.67442e-07, 3.073863e-07, 0.03379693, 0.08663794, 
    0.06806453, -0.0002587454, 0.0005391932, 3.037994e-06,
  1.05494e-06, -6.697844e-05, 0.009409389, 0.001106095, 0.0007819495, 
    0.001476745, 0.0331424, 0.06621757, 0.01139732, 0.0003098912, 0.01496478, 
    0.02441315, 0.05638639, 0.1184037, 0.09688996, 0.05323455, 0.007631939, 
    3.368206e-06, 1.559169e-07, 1.297706e-06, 7.266401e-06, 1.373079e-06, 
    6.026583e-06, 0.09583334, 0.0934635, 1.693169e-06, 1.73409e-06, 
    1.174207e-06, 2.217649e-07,
  0.005200746, 0.3701589, 0.2245832, 7.054731e-05, 0.0002891786, 0.09497947, 
    0.09402759, 0.2222418, 0.2062322, 0.1697304, 0.04690225, 0.08684819, 
    0.0524819, 0.04478535, 0.002169047, 2.65361e-05, 3.67149e-05, 
    3.855623e-06, 2.438717e-06, 0.000338336, 0.0003644426, 0.009566014, 
    0.04944995, 0.1776194, 0.008123728, 0.00119234, 9.037952e-05, 
    0.001026726, 4.95279e-05,
  0.166543, 0.134052, 0.09890001, 0.01808647, 0.0005464569, 0.00182738, 
    0.03583365, 0.1249658, 0.2096751, 0.1218816, 0.0575313, 0.1433392, 
    0.1765324, 0.1583021, 0.1373999, 0.1417208, 0.06531227, 0.02442825, 
    0.01663642, 0.09604388, 0.2208393, 0.3295276, 0.1780058, 0.110296, 
    0.05259434, 0.02789118, 0.06943895, 0.1440807, 0.1365592,
  0.01072509, 0.005620804, 0.002140753, 3.312591e-05, 0.0003816476, 
    0.02633714, 0.2284776, 0.07220685, 0.1097414, 0.05321782, 0.08917272, 
    0.1089761, 0.121171, 0.0389495, 0.04529326, 0.05157007, 0.03939841, 
    0.0001810823, 5.70935e-07, 0.01100138, 0.06284891, 0.1253329, 0.05579701, 
    0.09600732, 0.05262156, 0.05199916, 0.04491112, 0.06506572, 0.08454467,
  0.0760935, 0.01601411, 1.088656e-05, 1.46522e-05, -2.059431e-09, 
    6.682542e-08, 0.0006163482, 0.0918766, 0.1374673, 0.09597524, 0.05348199, 
    0.0493196, 0.08197589, 0.07253136, 0.04832872, 0.05263843, 0.05267692, 
    0.03875773, 0.00580347, -3.067973e-06, 0.08123891, 0.09402537, 0.1372331, 
    0.09155881, 0.0840396, 0.05068535, 0.05216708, 0.03431509, 0.05018264,
  0.1275724, 0.09964047, 0.02055779, 0.004170343, 0.01318255, 0.02298484, 
    0.006711189, 0.1161446, 0.1438561, 0.1442002, 0.1991195, 0.2040113, 
    0.1908797, 0.1650562, 0.1428836, 0.2401862, 0.1180128, 0.1212982, 
    0.05974545, 0.04833418, 0.1082582, 0.08327693, 0.09834162, 0.09965107, 
    0.1116075, 0.1267466, 0.08895326, 0.05901636, 0.09500259,
  0.0855248, 0.1431223, 0.141894, 0.126337, 0.1050222, 0.1026315, 0.02606463, 
    0.003508483, 0.005901521, 0.02432422, 0.06628312, 0.09569788, 0.1078789, 
    0.1728294, 0.1272183, 0.1094415, 0.1811367, 0.1846421, 0.1575481, 
    0.04581665, 0.05219689, 0.1223134, 0.1045369, 0.1042058, 0.1247785, 
    0.151824, 0.1968993, 0.1630235, 0.1355331,
  0.1259813, 0.06576274, 0.05166562, 0.05834337, 0.04092716, 0.02060405, 
    0.0453311, 0.01699864, 0.008351998, 0.01905978, 0.02878107, 0.02897823, 
    0.05143956, 0.06563311, 0.03497338, 0.06052169, 0.04906413, 0.08151589, 
    0.04648504, 0.06057434, 0.05726595, 0.07886803, 0.02307354, 0.05114175, 
    0.1012004, 0.1148556, 0.1390072, 0.05884877, 0.1118007,
  0.01156603, 0.02088801, 0.01105589, 0.0344875, 0.01160695, 0.005756257, 
    0.004218264, -0.0002332655, 0, 0.0006733335, 0.002226841, -0.0001971528, 
    0.01804731, 0.02295905, 0.03224026, 0.02880818, 0.02281412, 0.0250274, 
    0.04131855, 0.04764983, 0.03396314, 0.02138852, 0.01802543, 0.003983051, 
    0.04270078, 0.002847867, 0.005112309, 0.03717317, 0.01783592,
  0.0007511006, -1.926415e-05, 9.088102e-05, 0.000281333, 0.0003331595, 
    0.0004324738, 2.210203e-05, -1.362152e-05, 0.0009599487, -1.871918e-05, 
    0, 0, 0, -1.427544e-05, -1.526391e-05, 0.0001312652, 0.000681737, 
    0.007860795, 0.01747324, 0.01393012, 0.001057001, 0.0001335236, 
    -1.653958e-05, 0.0001437955, 0.001824308, 0.0001700768, -0.000370576, 
    0.002721934, 0.002266382,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 5.526361e-05, -3.929999e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003241539, 0.003146578, 0.0003177033, 0, 0, 0, 3.68042e-05, 
    -0.0001249226, 0.0002813287, 0.003331475, 0.01075998, 0.000194623, 
    -2.176948e-06, 0, 0,
  0.002153286, -3.614142e-05, 1.301678e-05, -2.14396e-05, 0.003999887, 
    0.002891596, 0.01049621, 0.009386914, 0.007887278, 0.002787023, 
    -5.360223e-05, 0.002913267, 0.002410092, 0.006937004, 0.00716194, 
    0.01180332, 0.007653472, 0.001247055, 0.004401793, 0.00781248, 
    0.01228958, 0.01532962, 0.008863374, 0.007486863, 0.01470659, 
    0.007948684, 0.00148016, 0.002500752, 0.002074753,
  0.07487527, 0.08190738, 0.0826539, 0.09935696, 0.1297061, 0.1302279, 
    0.1053276, 0.08835877, 0.05652831, 0.03199342, 0.04624666, 0.07305576, 
    0.079999, 0.08639333, 0.07749511, 0.04961868, 0.05137542, 0.05335718, 
    0.03854099, 0.07292865, 0.07287668, 0.06468399, 0.06658338, 0.03732157, 
    0.05692189, 0.05939817, 0.0430328, 0.08160913, 0.07892305,
  0.1681898, 0.1045977, 0.1251509, 0.168435, 0.1834641, 0.1150328, 0.1040052, 
    0.07549627, 0.0612676, 0.04392808, 0.04005411, 0.07214469, 0.07013464, 
    0.1084165, 0.06473089, 0.08220927, 0.1044949, 0.1013947, 0.1400533, 
    0.1044887, 0.157183, 0.1218379, 0.1100138, 0.05986895, 0.1339494, 
    0.1158877, 0.1763233, 0.1293979, 0.1851993,
  0.05236163, 0.0128764, 0.05117329, 0.06130595, 0.02838387, 0.01373724, 
    0.0005837815, -0.0001507934, 0.00186272, 0.002107081, 0.001927709, 
    0.01134682, 0.009667562, 0.01931541, 0.07416528, 0.11749, 0.09521037, 
    0.1181905, 0.2069603, 0.1148191, 0.03077017, 0.03720532, 0.03112263, 
    0.02184777, 0.05402513, 0.1091081, 0.08716574, 0.05298751, 0.04744155,
  5.461999e-07, 0.005328562, 0.06773327, 0.004722583, 0.01279374, 
    0.009782062, -0.0001442091, 0.01251488, 4.057724e-06, 1.016386e-08, 
    -1.54435e-07, -8.583368e-08, 0.001393755, 0.01496483, 0.05105766, 
    0.08892431, 0.06876832, 0.05122978, 0.001851692, 2.765958e-07, 
    4.860109e-09, 4.428348e-08, 5.213708e-08, 0.04067788, 0.06929035, 
    0.05921768, -1.894593e-06, 0.003558549, 1.48701e-06,
  3.659831e-07, -4.443825e-05, 0.008029686, 0.0005565663, 0.001799837, 
    0.000400183, 0.02700334, 0.06214213, 0.01305656, 0.0005160071, 
    0.01241176, 0.02009209, 0.05774133, 0.1179532, 0.08126867, 0.03601265, 
    0.006425541, -1.15466e-06, 2.058745e-07, 3.89834e-06, 1.650717e-06, 
    1.207394e-06, 9.660356e-06, 0.07054541, 0.06872158, 9.814463e-07, 
    5.972414e-07, 1.511739e-07, 3.973074e-07,
  0.0002851545, 0.3250106, 0.1486107, 0.002204038, 0.0007860261, 0.08123574, 
    0.07133742, 0.1690295, 0.1598462, 0.153223, 0.03884658, 0.07967994, 
    0.04314713, 0.04128944, 0.003780437, 1.246543e-05, 1.696287e-05, 
    6.944095e-07, 2.504539e-06, 4.026265e-06, 3.340334e-05, 0.003292705, 
    0.03118196, 0.1456107, 0.005567144, 4.502796e-06, 2.875726e-05, 
    8.339885e-05, -1.357811e-05,
  0.1368878, 0.1198605, 0.08215228, 0.01349948, 0.0003528027, 0.003261972, 
    0.02187494, 0.07642338, 0.1682159, 0.09049761, 0.03997959, 0.1048965, 
    0.1463034, 0.136468, 0.1204484, 0.1369211, 0.05808891, 0.02592907, 
    0.02033699, 0.09948958, 0.1864162, 0.3077461, 0.1455474, 0.07661127, 
    0.04628494, 0.02582568, 0.05900625, 0.1261254, 0.1239635,
  0.01233058, 0.001438834, 0.000975986, 4.139109e-05, 0.0002151033, 
    0.01482132, 0.2035601, 0.06004274, 0.08996929, 0.04744252, 0.07590662, 
    0.09276015, 0.1057827, 0.03146774, 0.0341701, 0.03787455, 0.02863808, 
    1.095125e-06, 2.68243e-07, 0.03021883, 0.05434955, 0.1157382, 0.04246271, 
    0.07304128, 0.04143578, 0.04269872, 0.04717951, 0.05812034, 0.05113046,
  0.06351229, 0.002974032, 6.121471e-06, 8.348779e-07, -3.940045e-08, 
    5.617304e-09, 0.0007442042, 0.1003114, 0.1456212, 0.1205897, 0.04804949, 
    0.04262727, 0.06163727, 0.06386046, 0.04112649, 0.04735966, 0.03484552, 
    0.02148888, 0.003550191, 4.528256e-05, 0.05970809, 0.08517633, 0.1218741, 
    0.079124, 0.07328543, 0.03617469, 0.03419773, 0.01969319, 0.04445228,
  0.1102456, 0.08678946, 0.01288139, 0.007161299, 0.01159406, 0.01730404, 
    0.01241927, 0.1618724, 0.1581833, 0.1747745, 0.1841293, 0.2073636, 
    0.1851398, 0.1615437, 0.1354708, 0.2473588, 0.1134817, 0.1386475, 
    0.05801293, 0.0367594, 0.1065293, 0.0707401, 0.08809396, 0.08888073, 
    0.09783935, 0.1197247, 0.08361389, 0.05094523, 0.0814346,
  0.09595677, 0.1840113, 0.1437941, 0.1446652, 0.1419067, 0.1591331, 
    0.09637282, 0.01678029, 0.02835599, 0.09056971, 0.1220791, 0.1171831, 
    0.1379518, 0.2027244, 0.1429733, 0.1129842, 0.2018906, 0.1889707, 
    0.1595258, 0.08537778, 0.08646949, 0.1147606, 0.1399389, 0.1377954, 
    0.1293172, 0.1629545, 0.1936381, 0.1534389, 0.1386456,
  0.1788305, 0.134872, 0.1161027, 0.09216075, 0.1015111, 0.1092056, 
    0.1260755, 0.1247959, 0.1001861, 0.1212661, 0.06013207, 0.07836089, 
    0.08941545, 0.1269944, 0.06793862, 0.1070821, 0.1144769, 0.1651574, 
    0.1357522, 0.119812, 0.1036032, 0.1799104, 0.1116791, 0.1165175, 
    0.1881698, 0.1973732, 0.1773903, 0.1197185, 0.170446,
  0.08686709, 0.1015473, 0.1000979, 0.1047516, 0.1544672, 0.1426771, 
    0.1209415, 0.1104403, 0.03138326, 0.01708369, 0.01707165, 0.03319837, 
    0.04584585, 0.05154015, 0.06734733, 0.07837291, 0.07732439, 0.1323238, 
    0.08824427, 0.1239867, 0.07492201, 0.04795307, 0.04733472, 0.04426087, 
    0.1034588, 0.01662819, 0.01351202, 0.1241057, 0.09219049,
  0.05742595, 0.06831773, 0.06867951, 0.07040943, 0.06348024, 0.03933807, 
    0.02881903, 0.02982516, 0.0148454, 0.01048348, 0.007866488, 0.01371767, 
    0.01762603, 0.02125534, 0.01771979, 0.01801152, 0.03161687, 0.02998902, 
    0.04225304, 0.03995681, 0.01301641, 0.009495252, 0.002636638, 
    -4.881842e-05, 0.002558418, 0.004205242, 0.003848481, 0.007827082, 
    0.06487799,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001287971, -7.606003e-05, 0,
  4.122146e-05, 0.0008327399, 0.003978805, 5.552812e-05, 0, 0, 0, 0, 0, 0, 0, 
    -6.810701e-06, -1.87331e-05, -0.0001654801, 0.006073967, 0.006617492, 
    0.007203278, 0.003020267, -7.339196e-06, -0.0001172573, 0.001016654, 
    0.007500705, 0.008050353, 0.01785943, 0.01828754, 0.001499568, 
    0.00645658, 0.002896523, 0.00181792,
  0.009928527, 0.01420034, 0.01157101, 0.01006804, 0.02317179, 0.01928685, 
    0.02778693, 0.02679947, 0.02031418, 0.01536578, 0.0176398, 0.03036746, 
    0.0616752, 0.08219982, 0.07010522, 0.08358379, 0.05905047, 0.04897546, 
    0.05112363, 0.03473722, 0.03966644, 0.03972438, 0.05554828, 0.05647323, 
    0.05962396, 0.03939361, 0.03169036, 0.01633097, 0.009370743,
  0.1585878, 0.1777366, 0.1538041, 0.1752622, 0.2053042, 0.191425, 0.1575463, 
    0.151803, 0.1380432, 0.130852, 0.1663441, 0.1774176, 0.1614316, 
    0.1531144, 0.1275666, 0.1309436, 0.1440924, 0.1554067, 0.1205658, 
    0.1691146, 0.1328491, 0.1282537, 0.1336641, 0.08256417, 0.121587, 
    0.1104303, 0.1100139, 0.1589309, 0.1436506,
  0.1672581, 0.08928992, 0.1211232, 0.1591019, 0.1519915, 0.09102233, 
    0.1070398, 0.07993504, 0.06199744, 0.05438204, 0.04660016, 0.08568281, 
    0.09179679, 0.1405602, 0.07863813, 0.09828736, 0.1067771, 0.1269125, 
    0.1239117, 0.1119975, 0.1598229, 0.1413001, 0.1342275, 0.08520482, 
    0.112104, 0.1198468, 0.171184, 0.1233256, 0.1840676,
  0.04670987, 0.005938546, 0.0358762, 0.05252842, 0.02922379, 0.01171106, 
    0.001945229, -0.0001632835, 0.00300109, 0.003025294, 0.0006804581, 
    0.0159655, 0.01528853, 0.02438586, 0.07745223, 0.1205539, 0.07256443, 
    0.09121045, 0.1964014, 0.09360614, 0.0231581, 0.02357607, 0.01876518, 
    0.01535641, 0.05262065, 0.09603912, 0.0669046, 0.04551079, 0.04650953,
  7.205722e-08, 0.005712418, 0.0583904, 0.004160208, 0.01098904, 0.02301906, 
    0.0005754823, 0.009644652, 1.136961e-06, 4.480432e-07, -3.044755e-06, 
    -1.042039e-08, 0.0001990783, 0.01920195, 0.05338975, 0.1003811, 
    0.04784504, 0.04515935, 0.001085726, -9.198083e-07, 4.157247e-09, 
    5.258539e-09, 5.14648e-09, 0.04442933, 0.05317022, 0.05260064, 
    -0.0003169177, 0.002790798, -5.760057e-07,
  4.167694e-07, 0.0006255354, 0.005891565, 6.934509e-05, 0.003280619, 
    0.0003520053, 0.02869955, 0.0619449, 0.01429662, 0.0005156894, 
    0.02094051, 0.02546398, 0.06006617, 0.1169313, 0.0668878, 0.0249311, 
    0.006808446, -6.870047e-07, 1.784422e-07, 4.878215e-07, 4.454491e-07, 
    5.477225e-07, 3.555724e-06, 0.05887948, 0.04922742, 5.945882e-07, 
    1.261335e-07, 1.86016e-08, 7.327156e-08,
  0.0006817334, 0.289989, 0.1094873, 0.002345412, 0.001353148, 0.06844917, 
    0.05739423, 0.1257469, 0.1147099, 0.1536954, 0.03913476, 0.06954806, 
    0.0350489, 0.02948395, 0.005756819, 0.0001241509, 6.014008e-06, 
    -3.578781e-05, 1.008651e-06, -1.965131e-05, 1.312704e-05, 0.003233706, 
    0.02621273, 0.09938192, 0.006282201, -7.68469e-05, 3.245686e-06, 
    1.533744e-05, 5.219218e-05,
  0.1172451, 0.1050971, 0.07445288, 0.02003067, 0.001117303, 0.003093179, 
    0.0159634, 0.03848044, 0.1141977, 0.0664243, 0.02346858, 0.07201648, 
    0.1136068, 0.1185503, 0.09513678, 0.126331, 0.05282527, 0.02610629, 
    0.03214623, 0.1180597, 0.1409997, 0.2715399, 0.1219755, 0.05109165, 
    0.04045399, 0.02118786, 0.05404838, 0.1159522, 0.1103698,
  0.01077048, 0.0005388345, 0.0003680886, 9.187386e-05, 0.0001732068, 
    0.0142115, 0.1787851, 0.05153802, 0.0674153, 0.04522753, 0.06975093, 
    0.07416017, 0.09740974, 0.02220566, 0.02409466, 0.0364203, 0.01364518, 
    -7.220301e-06, 2.321075e-07, 0.01751084, 0.05162707, 0.1088496, 
    0.02707966, 0.04834393, 0.03292898, 0.04011709, 0.06417869, 0.06071606, 
    0.02436161,
  0.06171252, 0.001914233, 1.311297e-06, 7.292435e-07, -3.00659e-06, 
    1.815161e-08, 0.0007693107, 0.09995667, 0.1569141, 0.113874, 0.04406853, 
    0.03071973, 0.04101977, 0.05320711, 0.03817194, 0.03939433, 0.03221158, 
    0.008329035, 0.0001582177, 0.00724184, 0.03690715, 0.07078871, 0.0973382, 
    0.06045194, 0.06337775, 0.02820833, 0.02707478, 0.009248562, 0.04674184,
  0.1060669, 0.08245353, 0.01114043, 0.006621741, 0.0107544, 0.01625273, 
    0.03053722, 0.1497339, 0.15452, 0.1557191, 0.1627946, 0.2006004, 
    0.1751127, 0.1566236, 0.1311066, 0.2345311, 0.1015863, 0.09934831, 
    0.04550987, 0.0304135, 0.07423308, 0.05538959, 0.09338523, 0.08297717, 
    0.08119442, 0.1139911, 0.08040798, 0.04245231, 0.07034269,
  0.08125752, 0.1849255, 0.1232991, 0.1359311, 0.1320142, 0.1428416, 
    0.107726, 0.0772509, 0.08060797, 0.134629, 0.1524769, 0.1266322, 
    0.1738232, 0.2154395, 0.154615, 0.1189457, 0.2256134, 0.185891, 
    0.1395129, 0.1117969, 0.08954988, 0.102134, 0.1403868, 0.1558411, 
    0.1271778, 0.165787, 0.1776675, 0.1517397, 0.1196551,
  0.2039131, 0.1742427, 0.1157946, 0.1484763, 0.1640129, 0.1170686, 
    0.1251849, 0.1782172, 0.1457728, 0.2038732, 0.1199204, 0.1383931, 
    0.1358982, 0.1617635, 0.1266242, 0.1471114, 0.1727865, 0.2220066, 
    0.2266232, 0.1498289, 0.1387076, 0.2131701, 0.1690735, 0.1701176, 
    0.2373686, 0.2041368, 0.194652, 0.1478261, 0.1760062,
  0.1978033, 0.1666226, 0.1603618, 0.1204207, 0.1869843, 0.2066938, 0.159034, 
    0.1452682, 0.09551622, 0.1262422, 0.1347104, 0.08647072, 0.1442626, 
    0.1313373, 0.1190739, 0.1302372, 0.154998, 0.1858361, 0.1292192, 
    0.1820687, 0.1182117, 0.1340026, 0.1297005, 0.1056837, 0.2209235, 
    0.02613135, 0.01682158, 0.2150661, 0.1759284,
  0.1662969, 0.1575533, 0.1230663, 0.1581227, 0.1897723, 0.167728, 0.1562424, 
    0.1268394, 0.1034592, 0.09063857, 0.08518183, 0.06760073, 0.05292009, 
    0.05251251, 0.05806673, 0.0887122, 0.1154723, 0.1253511, 0.1570449, 
    0.1189608, 0.0679348, 0.076947, 0.02737379, -0.005509798, 0.01801281, 
    0.004429696, 0.0008158188, 0.03061601, 0.166796,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.369178e-07, 0.0001577853, -3.648839e-05, 0, 0.0003569836, 
    -0.0001989028, 0,
  0.001959333, 0.007700481, 0.007866877, 0.002758801, -9.23535e-06, 
    -5.652511e-07, -1.694524e-05, 0, 0, 0, 0, -4.325582e-05, -0.0001979919, 
    0.01862042, 0.02718727, 0.01803755, 0.01593863, 0.02677911, 0.01743886, 
    0.005338683, 0.01954276, 0.02794685, 0.02313133, 0.03433292, 0.0467451, 
    0.03350352, 0.02917348, 0.01207314, 0.009972153,
  0.0441568, 0.04767249, 0.04461224, 0.04910167, 0.07897454, 0.08402409, 
    0.07351375, 0.06332771, 0.04832274, 0.02644514, 0.07481956, 0.1204554, 
    0.1769302, 0.1841997, 0.1801077, 0.1942642, 0.2012831, 0.1789224, 
    0.1070476, 0.1260808, 0.107323, 0.1319776, 0.1303999, 0.125005, 
    0.1363843, 0.1100559, 0.09629014, 0.0791308, 0.05697239,
  0.1918462, 0.2100758, 0.1965543, 0.2214145, 0.2098883, 0.2140613, 
    0.1896047, 0.1898137, 0.1636024, 0.1948799, 0.2132222, 0.2147357, 
    0.1805116, 0.1711134, 0.1750534, 0.1645857, 0.1935883, 0.1979782, 
    0.1761592, 0.2344911, 0.1879496, 0.1757673, 0.1907924, 0.1460084, 
    0.1726927, 0.158533, 0.1687769, 0.2135775, 0.1867513,
  0.1591383, 0.08358049, 0.1093842, 0.1395165, 0.1162153, 0.07923067, 
    0.1015557, 0.07191855, 0.05626255, 0.04825713, 0.04327526, 0.0912384, 
    0.08318627, 0.1318404, 0.08939861, 0.1130901, 0.1078311, 0.1290461, 
    0.1229426, 0.1216241, 0.1639625, 0.1420724, 0.1327102, 0.1046417, 
    0.08298485, 0.1145405, 0.1543798, 0.1244399, 0.1796179,
  0.034052, 0.004583641, 0.03033211, 0.04791763, 0.02788012, 0.01094504, 
    0.0002330993, -4.011133e-06, 0.0002035617, 0.00261666, 0.01108244, 
    0.03884596, 0.02492893, 0.0313981, 0.06148532, 0.1082097, 0.06843183, 
    0.0767297, 0.175164, 0.073867, 0.02392431, 0.01516859, 0.01339209, 
    0.01029202, 0.04941612, 0.08328498, 0.05972529, 0.04160835, 0.04523851,
  -7.01319e-10, 0.004183413, 0.05116417, 0.002228281, 0.007175968, 
    0.01920344, 0.0008156076, 0.01025582, -1.355506e-07, 3.393571e-07, 
    7.658104e-05, 1.651591e-07, 0.0001557284, 0.015134, 0.04985488, 
    0.1050555, 0.04273598, 0.03517624, 0.0006657851, -3.023446e-07, 
    4.258365e-09, 3.627295e-08, 1.253555e-08, 0.04538321, 0.03701295, 
    0.04454323, 0.002557539, 7.733917e-05, 9.911504e-08,
  4.817597e-07, 0.009215194, 0.00347847, 4.558824e-05, 0.004011115, 
    0.0008469002, 0.03442767, 0.0670145, 0.01505264, 0.0006985128, 
    0.02202305, 0.04487772, 0.09489559, 0.1263729, 0.0469253, 0.02067677, 
    0.006025247, 7.980809e-07, 5.698143e-08, 3.351081e-08, 3.184138e-07, 
    8.34478e-08, 3.995844e-05, 0.0528724, 0.03186355, 4.310291e-06, 
    2.062639e-08, 2.979268e-08, 7.887794e-08,
  0.007375727, 0.2626242, 0.08544597, 0.000782076, 0.002034611, 0.06677847, 
    0.05218237, 0.1013666, 0.06926066, 0.1613334, 0.04482597, 0.06161166, 
    0.0299762, 0.02295587, 0.006979582, 0.0007200368, 3.604981e-07, 
    -0.0001802484, -1.867118e-05, -7.740736e-05, 7.63016e-06, 0.003487429, 
    0.02138422, 0.06156179, 0.007151179, 5.581174e-05, -9.592782e-06, 
    -5.501756e-05, 0.0004451931,
  0.101109, 0.08980689, 0.07257638, 0.01919694, 0.0008423245, 0.002694279, 
    0.01782127, 0.022863, 0.0866495, 0.06538558, 0.01572956, 0.05285069, 
    0.09039318, 0.1097353, 0.08141971, 0.1233136, 0.04961998, 0.02885385, 
    0.04748974, 0.1522856, 0.1263623, 0.2405934, 0.115398, 0.03862036, 
    0.04059095, 0.01928467, 0.0570428, 0.1105001, 0.1002281,
  0.009300476, 0.0001803048, 0.0004187891, 0.0002910731, -5.959238e-05, 
    0.01645542, 0.1369584, 0.04852425, 0.06578165, 0.04442259, 0.06696311, 
    0.0650808, 0.09124924, 0.01836427, 0.01599553, 0.03443287, 0.003129122, 
    -1.777257e-05, 1.782224e-07, 0.01991504, 0.0526637, 0.1101409, 
    0.01854359, 0.03456868, 0.02647831, 0.03760836, 0.06124318, 0.05047755, 
    0.01405581,
  0.04522781, 0.0008423949, 4.722329e-07, 1.062158e-05, -4.145095e-05, 
    4.061985e-05, 0.001523112, 0.1018619, 0.1710544, 0.1210905, 0.03652733, 
    0.02827634, 0.02681716, 0.05421816, 0.03923332, 0.02989464, 0.0106283, 
    0.003527681, 3.685719e-05, 0.009217773, 0.02496801, 0.05543838, 
    0.07784113, 0.04672304, 0.05066973, 0.02048886, 0.02005346, 0.002753342, 
    0.05031813,
  0.0905631, 0.08937261, 0.01029059, 0.007188727, 0.01415098, 0.02019124, 
    0.05449586, 0.1232198, 0.134107, 0.1296299, 0.1403337, 0.2000329, 
    0.1537027, 0.1467004, 0.1306348, 0.2281242, 0.1035791, 0.08634706, 
    0.04233487, 0.02900819, 0.05457185, 0.0478923, 0.082535, 0.0818852, 
    0.07245076, 0.1080975, 0.08155259, 0.03547059, 0.05693643,
  0.08921851, 0.1680712, 0.1170779, 0.1217476, 0.1223551, 0.1263849, 
    0.09662928, 0.1453909, 0.1229811, 0.1775846, 0.1562395, 0.1318938, 
    0.1672067, 0.2036395, 0.1517733, 0.1275655, 0.2261769, 0.1937693, 
    0.1170655, 0.1074279, 0.07867411, 0.09443201, 0.1438406, 0.1579279, 
    0.1222331, 0.1552583, 0.1808403, 0.1527065, 0.113602,
  0.1918052, 0.203957, 0.1058573, 0.1577612, 0.1761301, 0.1200005, 0.1362143, 
    0.190739, 0.1626581, 0.2291217, 0.1366465, 0.1660076, 0.1771286, 
    0.1900013, 0.1712617, 0.2146948, 0.2200935, 0.2927543, 0.2683738, 
    0.1804218, 0.1434696, 0.2238695, 0.1678274, 0.2025835, 0.280683, 
    0.2151057, 0.1931604, 0.1375077, 0.1826826,
  0.2229306, 0.1757236, 0.18946, 0.1738949, 0.2107439, 0.2030658, 0.1782134, 
    0.2000746, 0.1254636, 0.1894547, 0.186996, 0.2371693, 0.190664, 
    0.1720305, 0.1382303, 0.1433593, 0.1823241, 0.2056254, 0.1735895, 
    0.2049113, 0.1601861, 0.1409351, 0.1406479, 0.1825004, 0.2315405, 
    0.07796622, 0.02191773, 0.2117448, 0.2386733,
  0.2108484, 0.1962178, 0.1534809, 0.2100744, 0.2172834, 0.1665718, 
    0.1738373, 0.1717326, 0.1652272, 0.2136088, 0.1788484, 0.1238199, 
    0.1151327, 0.1258445, 0.1694687, 0.2006046, 0.2019063, 0.2491759, 
    0.2656363, 0.2377457, 0.1674902, 0.1426132, 0.1117463, 0.06111781, 
    0.072172, 0.02286233, 0.03086204, 0.08364662, 0.2107399,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004779946, 0.004955797, 
    0.0116395, 0.009657743, -0.0002412439, 0, 0, -5.148037e-06, 
    -1.187745e-05, 0.002924164, 0.01915498, 0.01835811, -0.002069158, 
    0.001943837, 0.0002078158, 0,
  0.02583488, 0.02187859, 0.01978535, 0.006603842, -0.0001431403, 
    -1.738656e-05, 0.005781434, 0, 0, 0, -3.965897e-06, -6.606725e-05, 
    0.00451916, 0.07074612, 0.082941, 0.09975579, 0.1113814, 0.109599, 
    0.1024735, 0.08225259, 0.1372004, 0.1340436, 0.1460345, 0.1510524, 
    0.1808172, 0.1135506, 0.09341513, 0.05900367, 0.04122525,
  0.09830767, 0.1013571, 0.1127168, 0.1441536, 0.1271763, 0.1365809, 
    0.1300398, 0.1140821, 0.1125757, 0.1111726, 0.1512958, 0.1984883, 
    0.2581064, 0.2615045, 0.2194613, 0.2354033, 0.2374613, 0.2414834, 
    0.1546658, 0.1666596, 0.1730827, 0.1921162, 0.2210605, 0.2096368, 
    0.2019526, 0.1679665, 0.1639787, 0.1355998, 0.1478039,
  0.2143296, 0.2447284, 0.2113384, 0.2263388, 0.1925757, 0.2077225, 
    0.1933813, 0.2006978, 0.1746023, 0.226288, 0.2307534, 0.209386, 0.179707, 
    0.1685469, 0.16889, 0.1510266, 0.1798523, 0.1852616, 0.1686773, 
    0.2521978, 0.2214023, 0.2074266, 0.2184289, 0.1768654, 0.1815836, 
    0.1650692, 0.1769752, 0.2272772, 0.2148098,
  0.1448564, 0.06808812, 0.09667134, 0.1237695, 0.09495264, 0.08200964, 
    0.09379869, 0.07258317, 0.05507357, 0.03863564, 0.04109036, 0.09020105, 
    0.07245138, 0.1225183, 0.08872847, 0.1197991, 0.1156077, 0.1199489, 
    0.1221974, 0.1261001, 0.1681919, 0.1463651, 0.1282141, 0.1066, 
    0.06141788, 0.1047315, 0.1490043, 0.1213047, 0.1746702,
  0.02077482, 0.008143356, 0.03617333, 0.04831691, 0.02254117, 0.002862044, 
    1.023071e-05, -0.0001339195, 0.001837801, 0.001231154, 0.01944241, 
    0.04782233, 0.03393302, 0.04018834, 0.06541553, 0.09940673, 0.08235876, 
    0.07228859, 0.1712196, 0.06634317, 0.01744294, 0.005865691, 0.004260607, 
    0.01056435, 0.04725075, 0.08242124, 0.05905671, 0.0449505, 0.04067545,
  -6.841176e-10, 0.005212944, 0.04686072, 0.0008769194, 0.004922908, 
    0.01372142, 0.003121826, 0.01702655, 0.0007795463, 6.647032e-07, 
    2.327214e-05, 5.046062e-07, 0.0005284716, 0.01675034, 0.05235998, 
    0.1016959, 0.0360989, 0.0370442, 0.001277502, -9.533626e-09, 0, 
    3.835234e-08, -5.791033e-08, 0.03183956, 0.02934237, 0.03587928, 
    0.005535075, -1.732683e-05, 5.068082e-08,
  3.724152e-07, 0.00121587, 0.003068857, 2.096051e-05, 0.003190004, 
    0.001875111, 0.05083996, 0.05705712, 0.01255007, 0.0009268071, 
    0.02773374, 0.0634883, 0.09780413, 0.1253407, 0.04880945, 0.02247057, 
    0.005537844, 6.833468e-06, 1.634312e-08, 4.373702e-08, 1.386053e-07, 
    2.126116e-08, 0.001371448, 0.05066948, 0.02119853, 6.126846e-06, 
    9.943204e-09, 1.06016e-07, 1.517908e-07,
  0.008972704, 0.2358898, 0.08615745, 0.0004641643, 0.008322564, 0.07509716, 
    0.04863606, 0.08895987, 0.04817438, 0.1669243, 0.04068362, 0.0575968, 
    0.03064832, 0.02126398, 0.008562785, 0.002645353, 5.218066e-05, 
    0.0006320719, -2.148041e-05, -0.0001342652, 2.952789e-06, 0.00563001, 
    0.02682319, 0.04903057, 0.01223333, 0.0003802605, 0.0003295217, 
    7.632971e-05, 0.01346585,
  0.08965738, 0.07821323, 0.07525099, 0.02079372, 0.0009314298, 0.003019517, 
    0.01727473, 0.017222, 0.08841562, 0.06299922, 0.01210318, 0.04436061, 
    0.07498564, 0.1011762, 0.08018188, 0.1269252, 0.04734574, 0.03031785, 
    0.0592576, 0.1802801, 0.1239155, 0.220582, 0.1091, 0.03042057, 
    0.03903184, 0.02218432, 0.07297352, 0.1122073, 0.08738692,
  0.01107444, 6.2748e-05, 0.001042127, 0.002515629, 0.0004837926, 0.02690186, 
    0.1117096, 0.04474781, 0.0673669, 0.05778228, 0.07037763, 0.06695419, 
    0.08649289, 0.01675913, 0.0137174, 0.0269889, 0.001155509, -5.931025e-07, 
    6.86987e-08, 0.02180981, 0.05559465, 0.111304, 0.01876791, 0.02800061, 
    0.02011669, 0.03833713, 0.05640155, 0.03095458, 0.008353079,
  0.03764774, 0.001694051, 1.566618e-05, 0.0001825263, -2.964778e-05, 
    0.002544207, 0.002132245, 0.1119874, 0.1874321, 0.1436474, 0.03833467, 
    0.03135366, 0.02305202, 0.04928845, 0.04347505, 0.02659384, 0.008094575, 
    0.001172159, 0.0002748272, 0.001304105, 0.02125732, 0.04445338, 
    0.07269873, 0.04205755, 0.03862565, 0.01652167, 0.01873479, 0.00159303, 
    0.05199011,
  0.07339334, 0.09640758, 0.007218845, 0.006712496, 0.02562998, 0.02270211, 
    0.07128829, 0.08833551, 0.1120386, 0.1057821, 0.1189106, 0.1823286, 
    0.1396723, 0.1372362, 0.1171719, 0.2093363, 0.1030106, 0.05791328, 
    0.03444609, 0.03488173, 0.04330286, 0.04303345, 0.07429646, 0.07682028, 
    0.05542406, 0.1018201, 0.06694648, 0.02345276, 0.05392873,
  0.09592428, 0.1483975, 0.1162206, 0.1130063, 0.1109653, 0.1149924, 
    0.08208725, 0.1523477, 0.1644378, 0.1708771, 0.1508457, 0.1252488, 
    0.1587302, 0.1958838, 0.1433169, 0.1284169, 0.1998459, 0.1791866, 
    0.09996985, 0.09636259, 0.07252125, 0.0910989, 0.1443252, 0.1606487, 
    0.1192839, 0.146969, 0.1739839, 0.1443926, 0.1080349,
  0.1957745, 0.2017166, 0.1016334, 0.1498778, 0.1755047, 0.1226225, 0.134238, 
    0.1814228, 0.175633, 0.2048334, 0.1298157, 0.167411, 0.1768741, 
    0.1911136, 0.2008895, 0.2158353, 0.2131448, 0.3197674, 0.2944181, 
    0.1712664, 0.1326115, 0.2147992, 0.1703453, 0.2043765, 0.2800069, 
    0.2325643, 0.2091178, 0.142654, 0.1721386,
  0.2236229, 0.1777001, 0.1933713, 0.1785441, 0.2368755, 0.2186718, 
    0.1873945, 0.2117052, 0.1454598, 0.2029783, 0.2011807, 0.2455421, 
    0.1976204, 0.1896515, 0.1526884, 0.1352325, 0.1895562, 0.2007391, 
    0.162788, 0.1901256, 0.188139, 0.1561104, 0.1689817, 0.2175727, 
    0.2237561, 0.1164829, 0.05666674, 0.1934728, 0.2325683,
  0.2307594, 0.2160852, 0.1640778, 0.195122, 0.2143631, 0.1906929, 0.1889413, 
    0.1946472, 0.2014857, 0.2602201, 0.2451057, 0.2147983, 0.1932741, 
    0.1728429, 0.2090557, 0.2456149, 0.2477945, 0.273591, 0.2649589, 
    0.2774596, 0.2206335, 0.193553, 0.1487519, 0.1291554, 0.1333064, 
    0.07099395, 0.08008353, 0.104917, 0.2276064,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01485593, 0.04817046, 0.05447889, 
    0.04770369, 0.01719767, 0.0005480276, 1.317845e-05, -0.0001381089, 
    3.701916e-05, 0.008664897, 0.08562338, 0.1018529, 0.04150483, 0.07192023, 
    0.0005998794, 0,
  0.06155948, 0.06014332, 0.09893552, 0.03574114, -0.0006225406, 
    0.0005251642, 0.02756365, -8.563136e-05, -7.040913e-09, -0.0001422993, 
    -0.0001671895, -0.0003844316, 0.0330237, 0.136154, 0.1612683, 0.1758648, 
    0.1778575, 0.2040627, 0.219767, 0.1885239, 0.2297099, 0.2423025, 
    0.2390195, 0.2799577, 0.2830207, 0.235004, 0.2372516, 0.1534414, 0.108678,
  0.1392827, 0.1674454, 0.1790974, 0.1962149, 0.1973055, 0.1784629, 
    0.1773826, 0.1683312, 0.1514898, 0.1541738, 0.2019677, 0.2643349, 
    0.2955058, 0.3105733, 0.2526061, 0.2381407, 0.2404852, 0.2751302, 
    0.1893739, 0.1964416, 0.206632, 0.2203056, 0.2564289, 0.2233139, 
    0.2185221, 0.1974236, 0.1971035, 0.1879349, 0.2119039,
  0.2041441, 0.2403037, 0.2182281, 0.2025279, 0.1737686, 0.207658, 0.1963664, 
    0.2035751, 0.1808528, 0.2330172, 0.2317159, 0.2055649, 0.1879297, 
    0.160775, 0.1638434, 0.1444254, 0.1571943, 0.1675443, 0.1751646, 
    0.2498519, 0.218607, 0.2061451, 0.2162729, 0.1878586, 0.1672295, 
    0.1455413, 0.1740498, 0.2163276, 0.2024879,
  0.1333588, 0.06840448, 0.08862171, 0.1205302, 0.09057741, 0.08781621, 
    0.09032431, 0.06949469, 0.05381974, 0.03480154, 0.0403853, 0.08618202, 
    0.06681293, 0.1161861, 0.0946992, 0.113501, 0.1042713, 0.1130723, 
    0.1102849, 0.1111542, 0.1505981, 0.1426488, 0.1274949, 0.1074393, 
    0.0516789, 0.09731966, 0.1353544, 0.1270279, 0.1752757,
  0.01151698, 0.02906129, 0.05175245, 0.04509763, 0.02194662, 0.000493263, 
    -2.391178e-05, -8.327731e-05, 0.004460746, 0.000122068, 0.03132769, 
    0.05430347, 0.04346941, 0.04723438, 0.07214667, 0.09047608, 0.07592208, 
    0.06934754, 0.1551071, 0.05406979, 0.005390947, 0.00217665, 0.002140911, 
    0.01274373, 0.04556345, 0.08606354, 0.0623848, 0.04414883, 0.0288185,
  -2.402452e-07, 0.01945842, 0.04998313, 0.003560224, 0.006917284, 
    0.008068987, 0.01177678, 0.02122515, 0.006207697, 0.0003032268, 
    0.002950174, 0.0001847784, -9.074506e-05, 0.01330637, 0.04854873, 
    0.09584402, 0.02069151, 0.04709017, 0.0005217257, -2.300786e-10, 
    -3.388753e-10, 4.739775e-10, -5.86801e-07, 0.01601772, 0.0250911, 
    0.02809266, 0.007588627, -5.337841e-06, 4.742733e-08,
  7.029467e-07, 0.0003258349, 0.003419869, 0.0003995528, 0.003280088, 
    0.001932097, 0.05625825, 0.05442384, 0.008538559, 0.001504626, 
    0.02623777, 0.05463324, 0.1093747, 0.105539, 0.04736712, 0.02661514, 
    0.008985233, 3.844803e-06, -1.023266e-10, 5.592067e-08, 4.162904e-08, 
    1.947303e-08, 0.000146964, 0.03757697, 0.01454338, 1.665912e-05, 
    1.789111e-09, 7.917921e-08, 1.782012e-07,
  0.01827687, 0.2100999, 0.09840162, 0.003872849, 0.02212724, 0.07934952, 
    0.05023968, 0.08735929, 0.04229166, 0.1669442, 0.03680202, 0.0515312, 
    0.02651433, 0.01575032, 0.008601809, 0.002749944, 0.002249443, 
    -3.334301e-05, 0.002406734, -8.323452e-06, 4.345542e-06, 0.003444453, 
    0.03337574, 0.04463653, 0.008137476, 0.002123135, 0.0009606547, 
    0.005481166, 0.02576132,
  0.08650054, 0.06771607, 0.08891311, 0.0253098, 0.002814936, 0.005140054, 
    0.01796166, 0.0137537, 0.08349133, 0.06260838, 0.01195414, 0.03587444, 
    0.07347937, 0.09411979, 0.06971166, 0.1096211, 0.05057548, 0.0356052, 
    0.07342661, 0.2159881, 0.1376458, 0.1920934, 0.1083137, 0.02527614, 
    0.03653784, 0.02633063, 0.07799746, 0.1201742, 0.07881431,
  0.00179949, 0.0001191325, 0.001535265, 0.006853619, 0.0002494456, 
    0.02362485, 0.09219494, 0.0555362, 0.07690366, 0.04978353, 0.07650848, 
    0.0734998, 0.08746588, 0.02111479, 0.0123064, 0.02188736, 0.000928961, 
    1.573926e-06, -3.605622e-05, 0.0208184, 0.05376672, 0.1168269, 
    0.01453209, 0.02382411, 0.01627508, 0.03857795, 0.05213024, 0.02182205, 
    0.00379426,
  0.02903178, 0.0005197569, 5.301598e-06, 0.0006424562, 1.809701e-05, 
    0.003948244, 0.003204924, 0.1200089, 0.2194092, 0.1558593, 0.04438466, 
    0.035944, 0.02196471, 0.04675652, 0.04265678, 0.02064288, 0.006467719, 
    0.000130534, 0.0003456311, 0.0001394375, 0.02276856, 0.03932239, 
    0.06409533, 0.03793842, 0.03396943, 0.01608099, 0.0164155, 0.001615759, 
    0.0463714,
  0.06542149, 0.1035478, 0.007760641, 0.006982159, 0.04173703, 0.01729383, 
    0.08633316, 0.06247225, 0.08940515, 0.0834652, 0.09942965, 0.1616313, 
    0.1217672, 0.1287149, 0.103026, 0.1894177, 0.1161042, 0.05218251, 
    0.0371458, 0.03454105, 0.0438676, 0.06020328, 0.07244199, 0.08022976, 
    0.05312946, 0.09634723, 0.06033399, 0.02362316, 0.04976324,
  0.07886411, 0.137794, 0.1083178, 0.1119993, 0.09283589, 0.1104427, 
    0.07777151, 0.149558, 0.1651877, 0.1582845, 0.1469311, 0.1195895, 
    0.1554344, 0.2015304, 0.1363391, 0.1200204, 0.1813919, 0.1772166, 
    0.09404531, 0.09220283, 0.07988921, 0.07825851, 0.1423755, 0.1630902, 
    0.1246054, 0.1417071, 0.1617185, 0.1374865, 0.110053,
  0.1965162, 0.1927755, 0.1011562, 0.1546259, 0.1733575, 0.1192378, 
    0.1180148, 0.1664711, 0.1688639, 0.1875763, 0.114241, 0.1725183, 
    0.184229, 0.1868201, 0.1988471, 0.2111421, 0.2055957, 0.3389433, 
    0.2861342, 0.1633395, 0.1345461, 0.2169372, 0.1697098, 0.2050472, 
    0.2771889, 0.2406206, 0.2110598, 0.1383384, 0.1715303,
  0.2196001, 0.1632975, 0.1970949, 0.1837589, 0.2272721, 0.2207773, 0.189965, 
    0.2425455, 0.1772316, 0.2111881, 0.2051385, 0.2459284, 0.1914493, 
    0.1890644, 0.1582406, 0.1447307, 0.2088899, 0.2005243, 0.1564244, 
    0.1781108, 0.1884778, 0.1544298, 0.1580719, 0.2487112, 0.2249233, 
    0.1782502, 0.0964159, 0.1764841, 0.219339,
  0.2282251, 0.2329289, 0.1757008, 0.1836524, 0.217242, 0.2013323, 0.2102471, 
    0.216659, 0.2117251, 0.270711, 0.2487571, 0.2242985, 0.2058155, 
    0.1826554, 0.2077027, 0.2897451, 0.2798254, 0.2779989, 0.2504251, 
    0.2732227, 0.2197488, 0.1836106, 0.1749527, 0.1456603, 0.1500739, 
    0.1150236, 0.1428636, 0.09574911, 0.2331337,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -9.663455e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.943128e-05, 0.05473837, 
    0.06584632, 0.126816, 0.1612839, 0.09139181, 0.01257625, -8.699507e-05, 
    0.0002298236, 0.0008268371, 0.03382694, 0.1792278, 0.2162021, 0.1849014, 
    0.1640618, 0.02878859, 0.0009228116,
  0.1152341, 0.124045, 0.1384567, 0.1151714, -0.000449763, -0.001853888, 
    0.0558965, -0.001577515, -0.0005236699, -0.0003760352, -0.0002243341, 
    -0.0008599329, 0.08527213, 0.2384328, 0.2496838, 0.2175259, 0.2127262, 
    0.2332026, 0.2799594, 0.2602257, 0.2647365, 0.286696, 0.2739946, 
    0.3330673, 0.3493202, 0.2770327, 0.2867156, 0.1826587, 0.1715481,
  0.1740741, 0.2110482, 0.2093743, 0.2010044, 0.2335484, 0.2394841, 
    0.2463736, 0.2137401, 0.2493564, 0.2464115, 0.2855278, 0.314375, 
    0.3039077, 0.3155584, 0.2508509, 0.2283767, 0.2362729, 0.2696253, 
    0.1829272, 0.2075889, 0.216028, 0.2227455, 0.2650903, 0.2323831, 
    0.2270192, 0.1887238, 0.1806664, 0.1850711, 0.2084841,
  0.200655, 0.2373574, 0.2097457, 0.1895466, 0.1592196, 0.2099303, 0.1993957, 
    0.2206855, 0.1987333, 0.2392395, 0.2369912, 0.2081726, 0.1829747, 
    0.154309, 0.1575778, 0.1359093, 0.1284155, 0.1598441, 0.1608015, 
    0.2273206, 0.2081003, 0.2033197, 0.2020898, 0.1797635, 0.150533, 
    0.1532885, 0.170057, 0.2015474, 0.1936381,
  0.1233494, 0.0755187, 0.07465582, 0.1139661, 0.08565747, 0.08065279, 
    0.08078483, 0.0671966, 0.04909704, 0.03483112, 0.04175149, 0.08188927, 
    0.06384613, 0.1177196, 0.0974151, 0.1039838, 0.10269, 0.09752855, 
    0.1113372, 0.09410863, 0.1357633, 0.1276262, 0.1337942, 0.1092385, 
    0.04752751, 0.08988601, 0.1258017, 0.1218505, 0.1697497,
  0.01346716, 0.05631879, 0.07477645, 0.04965209, 0.01581847, 0.0001054028, 
    3.494603e-05, -1.904072e-05, 0.005809089, -0.0001816112, 0.05592389, 
    0.06273592, 0.04924753, 0.0467174, 0.07445031, 0.07973858, 0.07798146, 
    0.06196775, 0.1426114, 0.05284123, 0.001299074, 0.005503687, 0.00348434, 
    0.01586858, 0.05141827, 0.1033785, 0.06250122, 0.04596177, 0.02920893,
  -9.797699e-06, 0.02467594, 0.0528511, 0.001342011, 0.005731971, 0.02012139, 
    0.02630705, 0.02802862, 0.00391254, 2.373155e-06, 0.006915026, 
    0.004375826, -8.040019e-06, 0.01284056, 0.04366205, 0.08310291, 
    0.01361001, 0.0509792, 0.0002904252, 3.091148e-09, 5.352967e-11, 
    3.870105e-09, -1.555308e-06, 0.01152673, 0.02664816, 0.02044611, 
    0.009311857, 3.371791e-05, 7.119506e-08,
  5.021175e-07, 0.001853443, 0.003544405, 0.0005161975, 0.004448966, 
    0.002348281, 0.06623542, 0.06018075, 0.008001979, 0.002531317, 
    0.02209699, 0.04692788, 0.1161461, 0.09683095, 0.04223959, 0.02591737, 
    0.0095868, 7.836699e-05, 8.53499e-08, 1.411988e-07, 2.285238e-07, 
    6.768279e-08, 0.003732443, 0.03165305, 0.01412715, 0.0002170165, 
    6.280294e-07, 8.624651e-08, 3.914055e-08,
  0.01693424, 0.1973648, 0.1162215, 0.004015811, 0.02110573, 0.07883071, 
    0.05143993, 0.09792559, 0.0564631, 0.1673223, 0.03739174, 0.04873804, 
    0.03136459, 0.017158, 0.009204077, 0.002922342, 0.0002522117, 
    0.003538694, 0.009109182, 0.0007467417, 0.001139699, 0.0002702416, 
    0.03189681, 0.04955227, 0.0127545, 0.00919223, 0.00518163, 0.01990575, 
    0.0156002,
  0.09956916, 0.06392813, 0.08865757, 0.03734691, 0.01317006, 0.006724756, 
    0.02037154, 0.02064065, 0.1004595, 0.07861037, 0.01196104, 0.0321881, 
    0.08000946, 0.09508368, 0.06771722, 0.1114804, 0.06771504, 0.06783047, 
    0.09238318, 0.2416854, 0.1531957, 0.1787406, 0.1166633, 0.02734126, 
    0.0342177, 0.02867292, 0.09315121, 0.1289101, 0.08708175,
  0.003793489, 0.0001028915, 0.002218679, 0.005030434, 0.0001439413, 
    0.02704897, 0.1033014, 0.07063535, 0.08272326, 0.05034367, 0.08839351, 
    0.08063375, 0.09453115, 0.0232209, 0.01173619, 0.01617419, 0.001039092, 
    2.736563e-06, -4.043685e-07, 0.02025158, 0.05676074, 0.119898, 
    0.01425399, 0.02726997, 0.01761264, 0.04347819, 0.0488123, 0.01103138, 
    0.004897011,
  0.02463286, 0.0006570501, 2.901269e-06, 0.001778889, 0.002349466, 
    0.00114214, 0.002382442, 0.1221094, 0.2362449, 0.1701992, 0.05416856, 
    0.05050331, 0.02402254, 0.05005257, 0.04588021, 0.02129877, 0.006112205, 
    0.0001190575, 0.0002890835, -1.112286e-05, 0.0224, 0.03180796, 
    0.06153968, 0.03912635, 0.03452245, 0.01603471, 0.01629311, 0.001562114, 
    0.03467102,
  0.05475279, 0.1181278, 0.009521948, 0.007484973, 0.0459629, 0.0112744, 
    0.1049334, 0.04610939, 0.06261088, 0.06651741, 0.08412948, 0.1379696, 
    0.09442762, 0.1179835, 0.09113705, 0.1852846, 0.1159742, 0.05333105, 
    0.03104202, 0.03804135, 0.06047448, 0.0730481, 0.08408834, 0.07393958, 
    0.04613054, 0.09435998, 0.05390657, 0.02545035, 0.05506809,
  0.07284311, 0.1262476, 0.09999305, 0.1251602, 0.09033532, 0.1090576, 
    0.07144217, 0.1481705, 0.1613849, 0.1476257, 0.142258, 0.1065806, 
    0.1543768, 0.1778963, 0.1376076, 0.1224668, 0.1737691, 0.1742506, 
    0.09884599, 0.08490955, 0.07777996, 0.06174902, 0.1462298, 0.1856399, 
    0.1299907, 0.143816, 0.1399987, 0.138919, 0.1158811,
  0.1735301, 0.1990469, 0.1075291, 0.1480679, 0.1743897, 0.1230556, 
    0.1152682, 0.1511428, 0.1722173, 0.1823936, 0.09336273, 0.1686293, 
    0.1835682, 0.1903868, 0.1847747, 0.1985087, 0.1957136, 0.3527402, 
    0.2823105, 0.1608195, 0.1266444, 0.2083085, 0.1572752, 0.2388215, 
    0.2694943, 0.269355, 0.2128226, 0.1398772, 0.1646439,
  0.2426533, 0.1634837, 0.2252645, 0.2022309, 0.1976691, 0.2178996, 
    0.1899118, 0.2422024, 0.1974146, 0.2047855, 0.198691, 0.2515736, 
    0.1893531, 0.1801672, 0.1692903, 0.1501247, 0.2145123, 0.2062974, 
    0.1628937, 0.1918273, 0.2024609, 0.1485435, 0.1689844, 0.269919, 
    0.2437893, 0.215704, 0.1476598, 0.1609921, 0.2063996,
  0.237659, 0.2590778, 0.1754699, 0.1909032, 0.2219686, 0.2042369, 0.2141665, 
    0.2334039, 0.2299536, 0.2781639, 0.2600011, 0.2337137, 0.2021021, 
    0.1741637, 0.2048109, 0.3046924, 0.3043568, 0.2824842, 0.2412365, 
    0.2671279, 0.233075, 0.1943682, 0.1835439, 0.1575319, 0.1556405, 
    0.136531, 0.1621225, 0.09453128, 0.2404062,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.002804989, -0.0001251584, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002351855, 
    0.08352937, 0.169513, 0.2101979, 0.2112742, 0.1899384, 0.0656561, 
    0.004153368, 0.0007726399, 0.004165943, 0.07681195, 0.2963034, 0.2635133, 
    0.2324509, 0.208997, 0.09658788, 0.01002638,
  0.127846, 0.1844692, 0.1995898, 0.196435, 0.007483675, 0.01362814, 
    0.09293235, 3.296265e-05, 0.003013361, -0.001507973, 0.004642332, 
    0.01118385, 0.1728036, 0.2772609, 0.2708402, 0.2394427, 0.2313108, 
    0.2507542, 0.3000412, 0.2783239, 0.2603954, 0.2803578, 0.2967055, 
    0.3692427, 0.3678586, 0.2754331, 0.2769777, 0.1604382, 0.1773435,
  0.1903567, 0.2301267, 0.2252837, 0.2116803, 0.2628014, 0.2956609, 
    0.2721399, 0.2281256, 0.2780651, 0.2807301, 0.3038253, 0.3170935, 
    0.2887941, 0.3051301, 0.2395311, 0.227567, 0.230059, 0.2620533, 
    0.1969727, 0.2040039, 0.2149968, 0.2097578, 0.261047, 0.2194016, 
    0.2209639, 0.1821803, 0.179683, 0.1890094, 0.2175796,
  0.1989818, 0.2272488, 0.210271, 0.1878294, 0.146471, 0.2109512, 0.2151046, 
    0.2202101, 0.2055551, 0.2239946, 0.236905, 0.1939349, 0.1733158, 
    0.1554765, 0.1545675, 0.1384883, 0.1160359, 0.1720209, 0.1680735, 
    0.233062, 0.2087722, 0.1935517, 0.1949005, 0.1582229, 0.1379983, 
    0.1356696, 0.1597317, 0.1962766, 0.1907704,
  0.1143462, 0.06851315, 0.07654407, 0.102462, 0.08221403, 0.08081493, 
    0.08722275, 0.0695144, 0.05571154, 0.03204667, 0.04481648, 0.08294103, 
    0.06119639, 0.1141233, 0.09774446, 0.104394, 0.09518883, 0.08615926, 
    0.1027789, 0.08424998, 0.1357898, 0.1231227, 0.1382945, 0.110333, 
    0.04766271, 0.08866283, 0.1176266, 0.1200214, 0.1693541,
  0.007634751, 0.03284304, 0.0925112, 0.0502805, 0.01631159, 0.001291048, 
    4.063049e-05, 0.0001192707, 0.006382557, 0.0004168724, 0.06198725, 
    0.06581502, 0.05251983, 0.04240881, 0.07289396, 0.0773495, 0.09188356, 
    0.05923843, 0.1294584, 0.04363273, 0.00264524, 0.009155842, 0.003251332, 
    0.01980884, 0.07697126, 0.1084736, 0.06404226, 0.05803264, 0.02808641,
  0.00332822, 0.03131365, 0.0570271, 0.0005195054, 0.007428344, 0.02993665, 
    0.0349429, 0.03882788, 0.00526031, -1.000215e-05, 0.007217048, 
    0.01666553, 0.00115857, 0.009042728, 0.04985296, 0.05693741, 0.01414078, 
    0.06080827, 0.0002230024, 2.062835e-08, 1.462007e-09, 1.991518e-08, 
    -2.245903e-09, 0.005368189, 0.03330097, 0.03194686, 0.008404699, 
    1.715155e-05, 2.154607e-09,
  6.536528e-05, 0.01372063, 0.02244235, 0.001358128, 0.005809451, 
    0.004081558, 0.07360414, 0.08150645, 0.004578973, 0.001711018, 
    0.02316143, 0.04433776, 0.1298189, 0.1101929, 0.06065603, 0.03260629, 
    0.01320602, 0.0003461731, 2.121267e-06, 5.881075e-07, 1.050625e-06, 
    2.846243e-07, 0.008752208, 0.0380955, 0.01981981, 0.005590243, 
    -5.475245e-06, 9.32959e-07, -9.821788e-07,
  0.01566817, 0.2089858, 0.1607961, 0.004385365, 0.01768057, 0.07377686, 
    0.05984112, 0.1122674, 0.08949345, 0.1719741, 0.04905518, 0.05302463, 
    0.04016026, 0.01906108, 0.009745684, 0.003675856, 0.0008175762, 
    0.006067217, 0.012659, 0.005773011, 0.0002433263, 0.0008558091, 
    0.03693746, 0.07486687, 0.0137833, 0.01701219, 0.01289633, 0.03037151, 
    0.02933578,
  0.1208397, 0.07901267, 0.1000206, 0.05050182, 0.02196156, 0.00787139, 
    0.02830825, 0.03704362, 0.1514828, 0.1121618, 0.02411683, 0.03859245, 
    0.09978209, 0.1124392, 0.08226658, 0.1327306, 0.07733577, 0.08747683, 
    0.1151436, 0.2743033, 0.1917987, 0.1944453, 0.1413488, 0.0370333, 
    0.03831284, 0.04884544, 0.11526, 0.1410261, 0.1215471,
  0.00990075, 0.001563983, 0.003450442, 0.003633082, -2.190628e-05, 
    0.02096078, 0.1493547, 0.09897687, 0.1100849, 0.05484189, 0.09839569, 
    0.09604587, 0.1128853, 0.03000376, 0.01333836, 0.01652887, 0.001330973, 
    1.079758e-06, 4.475823e-05, 0.02597694, 0.07479793, 0.1336875, 
    0.01879426, 0.04585271, 0.02414212, 0.05145098, 0.05119723, 0.01172661, 
    0.008482466,
  0.01994094, 0.008364289, 2.334628e-06, 0.0004880789, 0.0004552743, 
    6.184493e-05, 0.004020694, 0.1295823, 0.2726772, 0.1722284, 0.06283537, 
    0.06405, 0.03647892, 0.05882024, 0.05114258, 0.02476521, 0.008631201, 
    0.0003543995, 0.003376246, 2.311398e-05, 0.03069777, 0.03401297, 
    0.06410819, 0.04565881, 0.03766435, 0.01990435, 0.020651, 0.002259636, 
    0.02725939,
  0.03914251, 0.09973545, 0.008340321, 0.01233351, 0.02879105, 0.007539607, 
    0.1212976, 0.03599365, 0.0411105, 0.05529919, 0.07476307, 0.121904, 
    0.0821788, 0.1221756, 0.09622028, 0.1839456, 0.1200858, 0.04893527, 
    0.03061727, 0.03636544, 0.0592266, 0.07440878, 0.08065987, 0.06799431, 
    0.04120703, 0.09494804, 0.05739774, 0.03432176, 0.05249414,
  0.08406184, 0.1285111, 0.1033761, 0.1303865, 0.08133423, 0.1021345, 
    0.06742309, 0.1465642, 0.1574965, 0.1438695, 0.1451168, 0.1140253, 
    0.1759358, 0.1750463, 0.1366988, 0.1345517, 0.1602154, 0.1667952, 
    0.1079428, 0.08377682, 0.07996227, 0.06099203, 0.1491681, 0.1894025, 
    0.1394092, 0.1377118, 0.1250471, 0.1440279, 0.1124061,
  0.17741, 0.1907024, 0.1232158, 0.1555537, 0.193004, 0.1292043, 0.1254356, 
    0.1482363, 0.1737087, 0.1756389, 0.08849276, 0.1741964, 0.1694029, 
    0.1982387, 0.180812, 0.193426, 0.2136205, 0.36009, 0.2788225, 0.1515805, 
    0.1284194, 0.1955589, 0.1500207, 0.2487686, 0.2968711, 0.2775773, 
    0.1917018, 0.139386, 0.170344,
  0.2499409, 0.1967962, 0.2783855, 0.2220724, 0.1919761, 0.2235444, 0.200986, 
    0.2498475, 0.2135749, 0.1865809, 0.2106743, 0.260393, 0.1974901, 
    0.1598485, 0.1766413, 0.1579826, 0.2279556, 0.1997503, 0.1787391, 
    0.2153048, 0.2188767, 0.1679687, 0.1775699, 0.2922515, 0.2600981, 
    0.220032, 0.1835361, 0.1434076, 0.2023814,
  0.2391687, 0.2494704, 0.1795939, 0.162153, 0.2027955, 0.1962512, 0.2106436, 
    0.2768526, 0.2598063, 0.2939274, 0.2527878, 0.2556698, 0.2304303, 
    0.170177, 0.2015115, 0.3318893, 0.3299339, 0.3087475, 0.2797178, 
    0.2929874, 0.2517509, 0.1925272, 0.1975168, 0.1681143, 0.1720557, 
    0.1336994, 0.1688771, 0.1037925, 0.2299957,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.009624109, -0.0003329164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008847316, 
    0.1332055, 0.1912823, 0.2103679, 0.241684, 0.2652742, 0.1566752, 
    0.08249711, 0.02234884, 0.01361641, 0.166717, 0.3090961, 0.2577283, 
    0.2311835, 0.2294139, 0.1374096, 0.03363602,
  0.1520853, 0.2340963, 0.2159724, 0.2532582, 0.02699933, 0.04987812, 
    0.1092372, 0.01077295, 0.01006302, 0.003979418, 0.02705508, 0.04670997, 
    0.2345296, 0.2729662, 0.2733484, 0.2428688, 0.24415, 0.257085, 0.3142532, 
    0.3003575, 0.2596096, 0.2651525, 0.2955266, 0.3696513, 0.3767931, 
    0.2867244, 0.2663105, 0.1558328, 0.1719329,
  0.1856982, 0.2284755, 0.2248127, 0.2035242, 0.2586911, 0.2879656, 
    0.2822117, 0.22634, 0.2842585, 0.277056, 0.2998624, 0.3200411, 0.2765306, 
    0.2939969, 0.2368458, 0.2255293, 0.2283148, 0.2502354, 0.201706, 
    0.2123013, 0.2272497, 0.2124037, 0.2488732, 0.2199344, 0.2154798, 
    0.1708575, 0.1813325, 0.1789424, 0.2219472,
  0.2005166, 0.2241189, 0.2061454, 0.1847448, 0.1465272, 0.2205486, 0.214529, 
    0.2200475, 0.2057082, 0.2182821, 0.2325306, 0.1996373, 0.1840578, 
    0.1480116, 0.1547358, 0.1527622, 0.111192, 0.177654, 0.1476135, 
    0.2222986, 0.1916593, 0.1808157, 0.1987972, 0.1556735, 0.1330362, 
    0.1276996, 0.146995, 0.1830175, 0.1805263,
  0.1271988, 0.07707974, 0.08352327, 0.0938586, 0.101347, 0.08055675, 
    0.08857542, 0.08164617, 0.06960429, 0.04785238, 0.04581918, 0.07941675, 
    0.05644424, 0.1071273, 0.09676643, 0.09589742, 0.09302045, 0.07674119, 
    0.1012599, 0.08062001, 0.1260994, 0.1211562, 0.1395597, 0.1159316, 
    0.04509296, 0.08775876, 0.1003605, 0.1178727, 0.1670075,
  0.008225973, 0.02118088, 0.08990812, 0.05108567, 0.02435478, 0.005146133, 
    4.004327e-05, 0.0004291667, 0.006815604, 0.002081256, 0.03942682, 
    0.04084117, 0.04985345, 0.04693675, 0.07008005, 0.0844302, 0.08504639, 
    0.05583959, 0.1251805, 0.04259131, 0.008173596, 0.01400123, 0.008752052, 
    0.02348317, 0.1007104, 0.1020868, 0.06402443, 0.05098718, 0.02515927,
  0.0002854977, 0.02629771, 0.07053663, 0.005482825, 0.008265449, 0.03374515, 
    0.03758473, 0.03168363, 0.003759608, 0.000876957, 0.01662862, 
    0.008640866, 0.0003752533, 0.01589872, 0.05505165, 0.04690154, 
    0.01925809, 0.06678425, 0.002522229, 4.698526e-08, -7.8133e-08, 
    5.111112e-08, 5.024761e-08, 0.003074826, 0.05494104, 0.06537274, 
    0.01301594, 0.0001010992, -3.533057e-05,
  0.002444966, 0.02641441, 0.09413371, 0.0006394865, 0.007414867, 
    0.006854698, 0.07730776, 0.09206745, 0.005640864, 0.002969639, 
    0.02664049, 0.05684188, 0.1433944, 0.1330392, 0.0822991, 0.03654081, 
    0.01192411, 0.001148788, 4.803696e-05, 4.39054e-07, 7.524673e-07, 
    6.62556e-07, 0.0129105, 0.04658648, 0.04749648, 0.04314767, 7.405508e-06, 
    1.212653e-06, 2.631361e-06,
  0.01937453, 0.2491387, 0.2194102, 0.00568051, 0.01196695, 0.06919138, 
    0.07440224, 0.1365733, 0.1185792, 0.2055258, 0.05403301, 0.06010441, 
    0.05070788, 0.02042583, 0.00669536, 0.00270705, 0.0007119452, 
    0.002050076, 0.008136578, 0.001152216, 0.0003074356, 0.004889703, 
    0.04967985, 0.1134846, 0.01500155, 0.008236559, 0.01163528, 0.02687458, 
    0.03688532,
  0.1485467, 0.09972759, 0.1244791, 0.09520835, 0.01811804, 0.006282208, 
    0.0344338, 0.04656661, 0.1872998, 0.1188901, 0.03990779, 0.04758569, 
    0.1111402, 0.1140933, 0.1020212, 0.1408085, 0.08274175, 0.113837, 
    0.1372814, 0.3082618, 0.2358491, 0.2155176, 0.1730462, 0.04978345, 
    0.03834508, 0.05994295, 0.1306477, 0.1716366, 0.16752,
  0.02045116, 0.006474494, 0.01350565, 0.0003598159, 0.002193255, 0.01215066, 
    0.2120606, 0.1100855, 0.1690931, 0.06165197, 0.09908839, 0.1024916, 
    0.116485, 0.03597508, 0.01626463, 0.01854714, 0.001865246, 4.506921e-07, 
    0.001128611, 0.03480775, 0.08641367, 0.1541751, 0.02018267, 0.063269, 
    0.02573478, 0.05557378, 0.05964377, 0.01008931, 0.009525074,
  0.004841643, 0.002487515, 1.063839e-05, 0.0001231354, 0.0009479934, 
    -1.099497e-05, 0.008678659, 0.1542422, 0.2884434, 0.1759253, 0.07810415, 
    0.07417894, 0.04147812, 0.05614788, 0.05700291, 0.03152831, 0.01382976, 
    0.001482064, 0.0001007289, 0.0001229377, 0.04354205, 0.04190405, 
    0.06850549, 0.05198411, 0.03707944, 0.02549874, 0.02399719, 0.002621099, 
    0.01255651,
  0.0295431, 0.07266346, 0.006699917, 0.01800651, 0.0251581, 0.006125575, 
    0.1340541, 0.03262054, 0.0270129, 0.0573041, 0.06197971, 0.1160953, 
    0.07827346, 0.1379927, 0.1059453, 0.2005292, 0.1178449, 0.04867189, 
    0.03113537, 0.03000922, 0.05079592, 0.08629642, 0.07783278, 0.07169995, 
    0.04745255, 0.09893927, 0.06862973, 0.0448285, 0.05042183,
  0.0768605, 0.1276992, 0.09970762, 0.1399866, 0.09010028, 0.09489607, 
    0.07201409, 0.1476794, 0.1499347, 0.1447489, 0.1492298, 0.1160705, 
    0.1564545, 0.1686028, 0.1431431, 0.1374402, 0.1632332, 0.1701997, 
    0.1109873, 0.08470026, 0.0802159, 0.05868461, 0.1596485, 0.1928801, 
    0.1428509, 0.1394948, 0.1308893, 0.1429586, 0.1235821,
  0.1617943, 0.1865348, 0.1309289, 0.1727579, 0.1834216, 0.1466254, 
    0.1372205, 0.1638868, 0.2007523, 0.1798512, 0.09597373, 0.1680517, 
    0.1614795, 0.187672, 0.1727869, 0.2061589, 0.2102473, 0.365714, 
    0.2687201, 0.1523239, 0.12538, 0.1994735, 0.1539255, 0.2796549, 
    0.3034987, 0.2939731, 0.2031265, 0.1431422, 0.1712125,
  0.2698921, 0.1990992, 0.2331713, 0.1954845, 0.1883671, 0.2123851, 
    0.2090057, 0.2805823, 0.2213598, 0.1916503, 0.2413815, 0.2736373, 
    0.2116972, 0.1509933, 0.2034362, 0.1861058, 0.2584356, 0.2029929, 
    0.1932942, 0.2433328, 0.2488654, 0.1465003, 0.189085, 0.3439594, 
    0.2528016, 0.2230437, 0.1898296, 0.1526338, 0.1984798,
  0.2375392, 0.2665178, 0.1789733, 0.1741454, 0.2346915, 0.2345441, 
    0.2123916, 0.2715541, 0.2514491, 0.2822925, 0.2304918, 0.2541724, 
    0.226525, 0.2021065, 0.2204291, 0.356393, 0.368032, 0.3847283, 0.3101217, 
    0.3454267, 0.2645283, 0.2175426, 0.2226923, 0.197917, 0.1829353, 
    0.1397093, 0.1668993, 0.1076412, 0.2297553,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.02194746, 0.003793808, -1.667902e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    -3.812882e-05, 0.01067143, 0.1622583, 0.1594512, 0.182184, 0.2331237, 
    0.3120196, 0.2093992, 0.1506223, 0.07948527, 0.08844966, 0.2032453, 
    0.3087524, 0.260134, 0.2255779, 0.2279863, 0.1707747, 0.06949261,
  0.1765525, 0.240117, 0.2174758, 0.2460482, 0.06685093, 0.07850636, 
    0.1137418, 0.02701082, 0.01733972, 0.04488172, 0.06732306, 0.1084043, 
    0.2839054, 0.285203, 0.2843232, 0.2586438, 0.2587981, 0.2337922, 
    0.3122653, 0.30804, 0.2524412, 0.2703878, 0.2999921, 0.3779509, 
    0.3756724, 0.2835336, 0.2727925, 0.1654265, 0.1871362,
  0.1907599, 0.2413038, 0.2271184, 0.2045261, 0.2603253, 0.2803306, 
    0.2926878, 0.2353421, 0.2818629, 0.2737369, 0.2862298, 0.3163189, 
    0.269345, 0.2814039, 0.2431761, 0.2459849, 0.2360329, 0.2556399, 
    0.2093849, 0.209885, 0.223106, 0.2262089, 0.2597685, 0.2121913, 
    0.2126367, 0.1830911, 0.1967461, 0.1970661, 0.2288769,
  0.2004718, 0.2128005, 0.2082874, 0.1832342, 0.1470763, 0.2097951, 
    0.2131901, 0.236182, 0.2119399, 0.2265893, 0.2400992, 0.2116766, 
    0.1842665, 0.1339782, 0.1409389, 0.1390067, 0.1168613, 0.1838269, 
    0.1544499, 0.2244369, 0.1975394, 0.1757534, 0.2002533, 0.1571119, 
    0.1236698, 0.1215569, 0.1542377, 0.2066513, 0.1872166,
  0.1228283, 0.08187303, 0.08766436, 0.07707488, 0.1043677, 0.09277232, 
    0.08814728, 0.07700762, 0.07101161, 0.04920848, 0.04163384, 0.06557922, 
    0.05454499, 0.1125008, 0.1015932, 0.09443986, 0.07420829, 0.07354792, 
    0.1037211, 0.09195956, 0.1225197, 0.1207166, 0.1397164, 0.1286972, 
    0.04316367, 0.09377049, 0.09602089, 0.1195559, 0.1629,
  0.009804332, 0.00638116, 0.07125892, 0.04675854, 0.03880028, 0.01119668, 
    0.0003588261, 0.003484802, 0.009328221, 0.005062848, 0.01396271, 
    0.02546834, 0.0493845, 0.05788581, 0.07076681, 0.08968166, 0.08994298, 
    0.06583917, 0.1212268, 0.05113368, 0.01821207, 0.02286138, 0.01073718, 
    0.01713265, 0.1014365, 0.09881181, 0.06783177, 0.04495315, 0.04047546,
  5.254355e-06, 0.01200355, 0.0762729, 0.01033717, 0.01291886, 0.03353059, 
    0.04532381, 0.03314879, 0.001797851, 0.003101929, 0.03873942, 0.03912945, 
    0.00194839, 0.02051054, 0.05544745, 0.04581919, 0.0326313, 0.0715396, 
    0.00939195, 4.80166e-07, 7.225226e-06, 4.951105e-08, 4.107497e-08, 
    8.611842e-05, 0.03622982, 0.09326853, 0.006522289, 1.860846e-05, 
    0.0001278664,
  0.0001694533, 0.01906755, 0.1599339, 0.008862035, 0.01052399, 0.01213576, 
    0.07749789, 0.08046259, 0.004446686, 0.002929797, 0.03219132, 0.03245148, 
    0.142671, 0.1032356, 0.08155534, 0.03895092, 0.01357477, 0.002931949, 
    1.798283e-05, 4.618456e-07, 2.976045e-07, -4.431198e-06, 0.007914877, 
    0.05307086, 0.05638129, 0.1567495, 7.366542e-05, -2.874516e-06, 
    0.0004255794,
  0.02782124, 0.2810246, 0.2404787, 0.002870817, 0.00855105, 0.06486867, 
    0.08089866, 0.1172221, 0.1223591, 0.2163649, 0.05026576, 0.03868581, 
    0.04042023, 0.0181159, 0.005124647, 0.002083245, 0.003547896, 
    0.003526077, 0.007863075, 0.001839484, 0.002402669, 0.01376369, 0.055213, 
    0.1243415, 0.01894411, 0.003482548, 0.0155924, 0.01829303, 0.01906986,
  0.1346652, 0.1146287, 0.1219822, 0.1433261, 0.01598223, 0.005445519, 
    0.0386815, 0.03806127, 0.1083838, 0.0996725, 0.02501104, 0.03264831, 
    0.08017153, 0.08351047, 0.08425839, 0.1313583, 0.08468561, 0.1276277, 
    0.1426564, 0.3115648, 0.227323, 0.192613, 0.1908694, 0.04960573, 
    0.03470764, 0.0613631, 0.117046, 0.1453449, 0.1922235,
  0.006020289, 0.005183662, 0.01055932, -8.086779e-06, 4.510081e-05, 
    0.0004708652, 0.1898082, 0.08968706, 0.1962977, 0.05669787, 0.08546747, 
    0.0778345, 0.08146003, 0.03106073, 0.0150682, 0.01871074, 0.001263705, 
    3.72703e-07, 0.001706252, 0.05208083, 0.06425375, 0.1462614, 0.01644149, 
    0.05620012, 0.02692618, 0.05291141, 0.05049472, 0.00361589, 0.005706262,
  0.0004715948, 0.007963839, 2.091424e-05, 2.921287e-06, 6.697084e-05, 
    -1.051477e-06, 0.005744047, 0.1801832, 0.3185577, 0.1756442, 0.07135427, 
    0.06634179, 0.03621036, 0.04051222, 0.06030161, 0.0373295, 0.01853286, 
    0.005271276, -2.668982e-06, 0.0001298211, 0.0643469, 0.03978726, 
    0.07198068, 0.05120129, 0.03447821, 0.0278564, 0.02821451, 0.003035956, 
    0.01062986,
  0.02747053, 0.04203236, 0.006125196, 0.02243398, 0.02301354, 0.008305209, 
    0.1263974, 0.03083563, 0.02187592, 0.05646453, 0.0622778, 0.11135, 
    0.07794847, 0.1453351, 0.1237087, 0.2202212, 0.1291458, 0.05615231, 
    0.02555258, 0.02279113, 0.04772608, 0.08142147, 0.08656988, 0.07244888, 
    0.06433667, 0.1029785, 0.07178394, 0.05949846, 0.05383949,
  0.08229928, 0.1302555, 0.104202, 0.1523248, 0.06998709, 0.07882852, 
    0.08903071, 0.1675355, 0.1466116, 0.1487486, 0.1493728, 0.130052, 
    0.1720599, 0.1654859, 0.1461707, 0.15078, 0.1554777, 0.162782, 0.1095228, 
    0.08266304, 0.07984544, 0.04786918, 0.1631895, 0.1964188, 0.1539796, 
    0.1347687, 0.1410336, 0.1529602, 0.1185203,
  0.1529784, 0.1935447, 0.145097, 0.185789, 0.1986099, 0.1533656, 0.1351963, 
    0.1814712, 0.2330638, 0.1806915, 0.104914, 0.1614901, 0.1819512, 
    0.2047202, 0.1816571, 0.198968, 0.2056377, 0.3877822, 0.2644104, 
    0.152264, 0.124935, 0.2201142, 0.1797547, 0.2921407, 0.2906669, 
    0.2840699, 0.2051685, 0.1441338, 0.1899454,
  0.2882379, 0.2153921, 0.2428, 0.2615846, 0.1941506, 0.2017323, 0.2308192, 
    0.2888961, 0.2346148, 0.1910826, 0.2628819, 0.2602377, 0.2379372, 
    0.1530802, 0.2374292, 0.1770444, 0.274377, 0.2321165, 0.1851987, 
    0.2528875, 0.2344759, 0.1548863, 0.2096708, 0.3614374, 0.289837, 
    0.2331915, 0.1922065, 0.1594895, 0.1925561,
  0.2002656, 0.2399133, 0.1714368, 0.1588054, 0.2260175, 0.2031688, 
    0.2250478, 0.304006, 0.2998686, 0.3014959, 0.256741, 0.255301, 0.2505347, 
    0.1911924, 0.2237498, 0.346882, 0.3615286, 0.3668728, 0.2925438, 
    0.3197186, 0.2542928, 0.2209184, 0.2559877, 0.2230214, 0.2092365, 
    0.1521074, 0.1777569, 0.1291526, 0.2200513,
  0, 0, 0, 0, 0, 0, 0, -3.572356e-07, -2.361388e-07, -1.15042e-07, 
    6.05484e-09, 1.271517e-07, 2.482485e-07, 3.693453e-07, -0.0001041714, 
    -8.105735e-05, -5.794332e-05, -3.482928e-05, -1.171525e-05, 1.139879e-05, 
    3.451282e-05, -0.0002308829, -0.000254118, -0.0002773532, -0.0003005883, 
    -0.0003238234, -0.0003470586, -0.0003702937, 0,
  0.03563856, 0.01123731, 0.003990224, -3.852637e-05, 0, 0, 0, 0, 0, 0, 0, 
    -2.584748e-05, 0.02436654, 0.1553961, 0.1388894, 0.175653, 0.2219451, 
    0.3297989, 0.2414134, 0.1918734, 0.1520897, 0.1825484, 0.2427357, 
    0.3141524, 0.2580209, 0.212554, 0.2329712, 0.1864506, 0.1230872,
  0.1822962, 0.2530506, 0.2257268, 0.2484309, 0.1262239, 0.08961345, 
    0.1256472, 0.06299917, 0.02343558, 0.1373934, 0.1167029, 0.1728072, 
    0.2894153, 0.3093781, 0.3011045, 0.3128322, 0.2797208, 0.3029, 0.3554741, 
    0.3275495, 0.2887209, 0.3314649, 0.3330384, 0.3908418, 0.3717337, 
    0.2727942, 0.3046204, 0.1806522, 0.2054948,
  0.2061434, 0.2429442, 0.2293467, 0.2164723, 0.2748675, 0.2761948, 
    0.2890453, 0.2460789, 0.2889969, 0.2936573, 0.2928298, 0.3249703, 
    0.2661575, 0.2731171, 0.2628109, 0.2434846, 0.2455521, 0.2575926, 
    0.2508537, 0.2235209, 0.2245752, 0.2326045, 0.2813739, 0.1945234, 
    0.2108333, 0.1994168, 0.207371, 0.2022602, 0.221091,
  0.2092751, 0.1981454, 0.199628, 0.1771058, 0.1565009, 0.2209963, 0.2325439, 
    0.2490819, 0.2229516, 0.2490273, 0.25025, 0.2078657, 0.1714628, 
    0.1361458, 0.1382312, 0.146708, 0.1383864, 0.1884505, 0.1612398, 
    0.2179008, 0.192209, 0.1663528, 0.1853895, 0.1682599, 0.1165867, 
    0.130749, 0.1566588, 0.1875792, 0.1919124,
  0.130817, 0.09322953, 0.1006157, 0.08312371, 0.1107522, 0.1055336, 
    0.09191251, 0.09151666, 0.07797456, 0.05614759, 0.04326595, 0.0693969, 
    0.04953384, 0.1249548, 0.09913746, 0.09816473, 0.07670892, 0.07366474, 
    0.107684, 0.085739, 0.1153962, 0.1211814, 0.1387994, 0.1431858, 
    0.03853121, 0.09456794, 0.09857289, 0.1306278, 0.1747723,
  0.01293756, 0.003274258, 0.04877726, 0.04082248, 0.03786992, 0.01779946, 
    0.003458255, 0.01574789, 0.01289141, 0.007283039, 0.003135481, 
    0.02317791, 0.0590107, 0.06484964, 0.07054408, 0.09529357, 0.09164165, 
    0.05776578, 0.1165449, 0.05555873, 0.03441694, 0.03634035, 0.01247234, 
    0.008279295, 0.0922618, 0.09529731, 0.07431425, 0.05323058, 0.0451006,
  3.489061e-07, 0.001708571, 0.07072932, 0.01084353, 0.02100992, 0.03623083, 
    0.05591844, 0.02190741, 0.001042876, 0.003036333, 0.02935066, 0.02462156, 
    0.002930935, 0.04370839, 0.05702652, 0.04870409, 0.03948939, 0.07860532, 
    0.02294736, 3.489566e-05, 0.0005397545, 2.207789e-08, -1.011845e-07, 
    4.889891e-06, 0.02743865, 0.09461988, 0.0030223, 1.385627e-05, 
    0.0002820972,
  -8.439661e-07, 0.005969724, 0.1221171, 0.03586733, 0.01463676, 0.01224698, 
    0.07046531, 0.07152795, 0.003116216, 0.001719594, 0.03479172, 0.02344485, 
    0.1396565, 0.08298944, 0.08161154, 0.04082976, 0.01865048, 0.004652241, 
    0.0002087899, 1.489814e-06, 2.270225e-07, -1.337473e-07, 0.002925798, 
    0.0361034, 0.04174046, 0.09212957, 0.0001878991, 1.189862e-06, 
    2.791092e-05,
  0.007285421, 0.2364485, 0.1629415, 0.00243762, 0.007687267, 0.04939299, 
    0.07063204, 0.08580595, 0.09493662, 0.1831813, 0.04633665, 0.02535215, 
    0.03495961, 0.0195571, 0.00675933, 0.002638664, 0.0006080136, 
    0.002702593, 0.005592122, 0.001746362, 0.0006782591, 0.01471282, 
    0.06373386, 0.08070125, 0.05041086, 0.002577594, 0.003239172, 0.01393101, 
    0.008862369,
  0.09083977, 0.07219489, 0.06213118, 0.1974085, 0.02823218, 0.005397674, 
    0.0548687, 0.03725504, 0.07144336, 0.08586095, 0.01719737, 0.02610535, 
    0.06102235, 0.06339891, 0.07319906, 0.1151466, 0.08555822, 0.1309857, 
    0.1443014, 0.3015375, 0.2257707, 0.174024, 0.1740166, 0.04043878, 
    0.02979108, 0.05485189, 0.1062225, 0.1004714, 0.1505721,
  0.0004609932, 0.0008778119, 0.01212509, -1.270031e-05, 4.088208e-06, 
    -0.0001266301, 0.1557958, 0.08288603, 0.1741226, 0.05802713, 0.08068754, 
    0.06287318, 0.06456968, 0.02820159, 0.01485184, 0.02216699, 0.001659433, 
    -2.281332e-05, 0.001052656, 0.05137265, 0.05031291, 0.1428845, 
    0.01572727, 0.04415883, 0.0267686, 0.04722912, 0.03690098, 0.0002475508, 
    0.001295477,
  5.310255e-05, 0.006724284, 4.67584e-05, 5.31176e-07, 6.96507e-06, 
    5.548655e-07, 0.005004559, 0.2427503, 0.3710336, 0.1771258, 0.06030938, 
    0.07423589, 0.0331273, 0.03210939, 0.04966702, 0.0364951, 0.01895529, 
    0.01200105, -4.592532e-08, 0.0001008176, 0.07571646, 0.03710124, 
    0.05992508, 0.04464118, 0.0271481, 0.02796812, 0.02000167, 0.003654898, 
    0.006916346,
  0.02742912, 0.02904835, 0.008795138, 0.02779123, 0.01833935, 0.004597155, 
    0.110495, 0.01692146, 0.02032861, 0.07519288, 0.06018797, 0.1131534, 
    0.07900582, 0.1477958, 0.1167846, 0.2197052, 0.1379822, 0.07458831, 
    0.02693022, 0.01642969, 0.05173416, 0.08317158, 0.08435708, 0.06317024, 
    0.0628557, 0.0965706, 0.07445354, 0.06749007, 0.06318576,
  0.08605784, 0.1401101, 0.1296538, 0.1757283, 0.07826942, 0.06779727, 
    0.1145426, 0.1941404, 0.1483597, 0.1521952, 0.1617346, 0.163403, 
    0.1823962, 0.1762857, 0.157028, 0.1533304, 0.1554438, 0.1678318, 
    0.113305, 0.08279338, 0.09535523, 0.04178656, 0.1802512, 0.2114082, 
    0.1497954, 0.1299327, 0.1554846, 0.1734982, 0.120799,
  0.1591745, 0.1941426, 0.1377882, 0.1847906, 0.2225422, 0.1508803, 
    0.1581436, 0.1993033, 0.2169504, 0.2062103, 0.1189961, 0.188741, 
    0.2101541, 0.2217321, 0.1878748, 0.1995481, 0.205594, 0.4106222, 
    0.2765845, 0.1392532, 0.1196337, 0.236326, 0.1607581, 0.2901156, 
    0.3321701, 0.2891545, 0.2295007, 0.1534294, 0.1841101,
  0.2634615, 0.1884094, 0.2754271, 0.2348477, 0.2214242, 0.2323062, 
    0.2221579, 0.2730104, 0.2310135, 0.2076871, 0.2770037, 0.2693018, 
    0.2377112, 0.1906162, 0.2808139, 0.2246691, 0.2634747, 0.2191048, 
    0.207177, 0.248669, 0.2193793, 0.1257925, 0.2422445, 0.3677977, 
    0.2812917, 0.2534493, 0.2010567, 0.1541633, 0.1846134,
  0.2172959, 0.2250656, 0.181371, 0.123762, 0.183523, 0.199247, 0.2212053, 
    0.2871294, 0.2910866, 0.3254135, 0.2950467, 0.3031387, 0.2651393, 
    0.2387603, 0.2790129, 0.4086791, 0.3734909, 0.3351331, 0.3354441, 
    0.29981, 0.248556, 0.22812, 0.2896617, 0.2778525, 0.2446454, 0.1819944, 
    0.207784, 0.1470039, 0.2223031,
  0.0009261662, 0.0005840055, 0.0002418447, -0.0001003161, -0.0004424768, 
    -0.0007846376, -0.001126798, 6.510878e-05, 6.539975e-05, 6.569072e-05, 
    6.598169e-05, 6.627267e-05, 6.656363e-05, 6.685461e-05, -0.001592777, 
    -0.001163497, -0.0007342161, -0.0003049354, 0.0001243453, 0.000553626, 
    0.0009829067, 0.0008662564, 0.0007788455, 0.0006914346, 0.0006040237, 
    0.0005166128, 0.000429202, 0.0003417911, 0.001199895,
  0.07053213, 0.02067724, 0.01231779, 0.0007895799, 0, -4.66224e-07, 0, 0, 0, 
    0, 0, 0.001015556, 0.04264818, 0.1321044, 0.1371365, 0.1676212, 
    0.2343255, 0.3224269, 0.2622012, 0.2114625, 0.199059, 0.2655875, 
    0.2523085, 0.3259247, 0.2618999, 0.2021465, 0.2288687, 0.1989189, 
    0.1584441,
  0.1751445, 0.2568839, 0.2389455, 0.242033, 0.1785496, 0.09455516, 
    0.1289227, 0.1231228, 0.09485202, 0.2155415, 0.2218405, 0.2305718, 
    0.2707044, 0.3219022, 0.3145698, 0.3272596, 0.2888626, 0.2701962, 
    0.3845508, 0.3657356, 0.3060566, 0.3083004, 0.3257445, 0.4292985, 
    0.3611889, 0.2732037, 0.3065584, 0.2143723, 0.20979,
  0.2373168, 0.2682312, 0.2433439, 0.2182987, 0.296389, 0.2500109, 0.2993559, 
    0.2735295, 0.305202, 0.3075108, 0.2914982, 0.3155926, 0.2619209, 
    0.280776, 0.2590643, 0.2622175, 0.257147, 0.2788801, 0.2601846, 
    0.2575511, 0.2463889, 0.2503296, 0.2908127, 0.2202853, 0.2123243, 
    0.2076733, 0.1877458, 0.218869, 0.2635674,
  0.2392704, 0.2185539, 0.21578, 0.1826201, 0.1801481, 0.2215719, 0.235459, 
    0.2551594, 0.2281919, 0.2683184, 0.2564189, 0.2048443, 0.1682747, 
    0.1501009, 0.1419321, 0.1470952, 0.1448373, 0.2312839, 0.1986997, 
    0.2295529, 0.2098955, 0.1963941, 0.2159652, 0.1731927, 0.1380641, 
    0.1363141, 0.1709194, 0.2229377, 0.2009772,
  0.1472225, 0.1239089, 0.1091695, 0.07951859, 0.1229802, 0.1216637, 
    0.1126528, 0.1172807, 0.08592449, 0.07746855, 0.04949547, 0.07096595, 
    0.05462178, 0.132301, 0.1017374, 0.1120136, 0.09069074, 0.075371, 
    0.1253924, 0.08963025, 0.1140006, 0.1370777, 0.1625145, 0.1606322, 
    0.04552501, 0.1005067, 0.1059762, 0.1515831, 0.1867872,
  0.01463036, 0.001056538, 0.04208257, 0.04333793, 0.03522103, 0.02058639, 
    0.01533064, 0.02452384, 0.01718711, 0.008799658, 0.002581637, 0.01828416, 
    0.07701258, 0.07660577, 0.09092079, 0.1121203, 0.09789361, 0.06782691, 
    0.125448, 0.08150826, 0.05805369, 0.05194421, 0.01504551, 0.00135135, 
    0.06373198, 0.09328471, 0.07893161, 0.06083306, 0.05833345,
  3.750977e-08, 0.0002875326, 0.07781917, 0.01076896, 0.04367834, 0.04359193, 
    0.05737744, 0.008914403, 0.004627614, 0.0006448552, 0.004847449, 
    0.00685059, 0.005447062, 0.05262152, 0.06389858, 0.04301195, 0.04362581, 
    0.08287912, 0.0500293, 0.006847689, 0.0008009452, 8.041054e-05, 
    3.276233e-08, 3.959926e-05, 0.02375443, 0.05936035, 0.002855042, 
    0.0001161203, 0.001433376,
  6.02639e-07, 0.002719047, 0.06989861, 0.1136832, 0.01821878, 0.01237355, 
    0.06605269, 0.07022545, 0.003928022, 0.001879138, 0.03541985, 0.02324453, 
    0.1516145, 0.07533652, 0.08290795, 0.04530941, 0.03160897, 0.009160042, 
    0.003789824, 1.338102e-05, 4.289398e-07, -1.075978e-07, 0.001262419, 
    0.03559056, 0.02143053, 0.02694173, 0.003666596, 3.227184e-06, 7.22719e-07,
  0.001316248, 0.2000039, 0.08568753, 0.006080138, 0.007070825, 0.03746386, 
    0.06176095, 0.07263616, 0.08619489, 0.1759259, 0.03768288, 0.02139074, 
    0.03354066, 0.02086697, 0.01224227, 0.004442816, 0.0009399223, 
    0.0003113642, 0.001606928, 0.0002492912, 0.0008444472, 0.01296983, 
    0.07707424, 0.06802242, 0.08764577, 0.001767375, 0.003638498, 
    0.004255163, 0.001212099,
  0.07059366, 0.05278471, 0.04001066, 0.2499295, 0.04597667, 0.008722829, 
    0.07138248, 0.03676353, 0.05207545, 0.07899322, 0.0154677, 0.02521708, 
    0.05080393, 0.05488982, 0.06785947, 0.1044489, 0.1030552, 0.1542033, 
    0.1569075, 0.28901, 0.2097595, 0.1631635, 0.1682559, 0.03741549, 
    0.02542748, 0.04545863, 0.09547284, 0.08446956, 0.1202755,
  7.673221e-05, 4.296908e-05, 0.01462782, -8.686687e-06, 2.126617e-07, 
    -1.912914e-05, 0.1362799, 0.08495042, 0.1932978, 0.06674464, 0.09016247, 
    0.05794664, 0.05679305, 0.02876925, 0.01980973, 0.03141077, 0.005517376, 
    0.007898608, 0.0005296412, 0.06867921, 0.04869629, 0.1530583, 0.01733806, 
    0.03729647, 0.0268204, 0.04504991, 0.03036962, 6.632171e-05, 0.0005053746,
  1.41123e-05, 0.001261279, 0.00271405, 2.025546e-07, 2.776181e-06, 
    3.054534e-07, 0.008803095, 0.3104926, 0.3773448, 0.1793032, 0.0604437, 
    0.08257459, 0.03744268, 0.03095822, 0.0454849, 0.03614708, 0.02484648, 
    0.02199741, 4.979387e-07, -1.217522e-05, 0.07129419, 0.05231675, 
    0.06325854, 0.04974789, 0.02351565, 0.03209518, 0.018899, 0.004882633, 
    0.004704251,
  0.02981915, 0.01887551, 0.007747712, 0.0348231, 0.01170938, 0.006109488, 
    0.1045508, 0.007004883, 0.02197117, 0.09274344, 0.06600922, 0.107339, 
    0.0813536, 0.1514278, 0.1250752, 0.2129367, 0.1542422, 0.07586461, 
    0.03197113, 0.006840153, 0.04048376, 0.07890876, 0.0817679, 0.05822675, 
    0.06065861, 0.09171352, 0.06463188, 0.08264399, 0.06549909,
  0.09788552, 0.1525592, 0.1477801, 0.2005485, 0.08119789, 0.07875174, 
    0.1449382, 0.2131899, 0.1498182, 0.1535951, 0.1749165, 0.182769, 
    0.2167926, 0.1997967, 0.1580626, 0.1669952, 0.1655847, 0.174692, 
    0.1433445, 0.08470321, 0.1049337, 0.0488593, 0.2350536, 0.2334449, 
    0.2065682, 0.1473385, 0.1694733, 0.1932677, 0.1396737,
  0.1746032, 0.2012568, 0.1797356, 0.1866535, 0.2288971, 0.1942155, 
    0.1610803, 0.2090711, 0.2343148, 0.2275366, 0.1792311, 0.1987702, 
    0.2322547, 0.232378, 0.1818537, 0.2439069, 0.2182393, 0.4361308, 
    0.2838562, 0.1464265, 0.1361473, 0.2513435, 0.1811398, 0.3149451, 
    0.3428115, 0.2899394, 0.2226772, 0.1746689, 0.2175215,
  0.3129886, 0.2228683, 0.3019511, 0.282691, 0.2788437, 0.2647687, 0.2466758, 
    0.2904619, 0.2394893, 0.2272471, 0.2928209, 0.327761, 0.2324388, 
    0.1997678, 0.3754412, 0.2246851, 0.2679956, 0.2482629, 0.1883392, 
    0.2280234, 0.2132785, 0.148097, 0.2128917, 0.3706177, 0.256055, 
    0.3080208, 0.208013, 0.1345438, 0.232704,
  0.22518, 0.2104521, 0.1708455, 0.1801379, 0.1949755, 0.2278146, 0.2771189, 
    0.2968743, 0.3028378, 0.3077325, 0.3182146, 0.3520962, 0.3355657, 
    0.2669483, 0.2631475, 0.3956856, 0.3730019, 0.3299981, 0.3267498, 
    0.3431441, 0.289735, 0.2694151, 0.3080603, 0.3040997, 0.2979459, 
    0.2619396, 0.2202826, 0.1588534, 0.2649069,
  0.004401739, 0.002623893, 0.0008460466, -0.0009317995, -0.002709646, 
    -0.004487492, -0.006265338, 0.0003786708, 0.0004416573, 0.0005046438, 
    0.0005676302, 0.0006306167, 0.0006936032, 0.0007565896, -0.006945321, 
    -0.004726696, -0.002508071, -0.0002894451, 0.00192918, 0.004147806, 
    0.006366431, 0.007205737, 0.006701972, 0.006198206, 0.005694441, 
    0.005190674, 0.004686909, 0.004183143, 0.005824015,
  0.0965343, 0.03723691, 0.02267187, 0.01029129, 0.001088939, 7.841366e-05, 
    1.120343e-05, 0, 0, 0, 0.0001807813, 0.01034521, 0.06677813, 0.1270462, 
    0.1153727, 0.1547068, 0.2285951, 0.324154, 0.2751013, 0.2352626, 
    0.2255888, 0.2923073, 0.2696922, 0.3293661, 0.2554217, 0.1953174, 
    0.2387203, 0.2176369, 0.1899604,
  0.1655038, 0.2339451, 0.2400238, 0.2421901, 0.2085947, 0.09466959, 
    0.1349989, 0.1747558, 0.2130831, 0.2577484, 0.2637981, 0.2740916, 
    0.2746601, 0.3117579, 0.3184642, 0.2954114, 0.2741709, 0.2475792, 
    0.3508556, 0.3055331, 0.2696507, 0.2719652, 0.3146818, 0.4411638, 
    0.3451611, 0.2794592, 0.2721571, 0.1945353, 0.2229038,
  0.2202868, 0.266057, 0.2471934, 0.2439672, 0.3113344, 0.2613739, 0.3055986, 
    0.2672265, 0.3046577, 0.3018965, 0.2923722, 0.3169588, 0.2583876, 
    0.287125, 0.2843164, 0.2931679, 0.2691566, 0.2873178, 0.2639608, 
    0.2650373, 0.2617732, 0.2700067, 0.3021841, 0.2499684, 0.2131929, 
    0.1956135, 0.221984, 0.2297381, 0.2628531,
  0.238412, 0.2353284, 0.2213778, 0.1831878, 0.1970273, 0.2245091, 0.2513155, 
    0.2699082, 0.230638, 0.2875236, 0.2654837, 0.2013594, 0.1693219, 
    0.1667248, 0.1545822, 0.1781421, 0.1740114, 0.2583966, 0.2400685, 
    0.2343073, 0.2140368, 0.2240748, 0.2188518, 0.1766626, 0.1212206, 
    0.1507419, 0.1812044, 0.2452032, 0.2027397,
  0.1764089, 0.1490572, 0.1261, 0.0878247, 0.1263317, 0.1556606, 0.1451755, 
    0.1259923, 0.105393, 0.1014155, 0.06599063, 0.07636814, 0.06890165, 
    0.127796, 0.1074594, 0.1118658, 0.10353, 0.0913697, 0.1517229, 0.116768, 
    0.1380531, 0.1480131, 0.1920691, 0.1801375, 0.03712182, 0.119165, 
    0.1250773, 0.1740809, 0.2014361,
  0.02148343, 0.001273177, 0.0330206, 0.0374691, 0.04018262, 0.02480739, 
    0.01923792, 0.02521645, 0.02363184, 0.009613793, 0.003160001, 0.01357771, 
    0.09044898, 0.08105282, 0.1063048, 0.1235022, 0.1017219, 0.07830882, 
    0.1382943, 0.1014893, 0.07637842, 0.08054236, 0.02197372, 0.0003821831, 
    0.04230709, 0.08580993, 0.08127832, 0.06771494, 0.06819241,
  2.095705e-08, 0.0002358944, 0.0512097, 0.006495514, 0.05478007, 0.04947461, 
    0.05693822, 0.006278918, 0.005739423, 0.0001291254, 0.0001000278, 
    0.007075067, 0.01151088, 0.06936941, 0.06807971, 0.04287225, 0.04432262, 
    0.09300441, 0.07102565, 0.03813249, 0.008744188, 0.002028076, 
    8.720214e-08, 1.264313e-05, 0.01266656, 0.02554267, 0.01752142, 
    0.000747134, 0.001994293,
  1.534232e-07, 0.0002562006, 0.0222793, 0.1488534, 0.02568595, 0.01362182, 
    0.06043803, 0.07926568, 0.007800998, 0.003939388, 0.03056277, 0.0249512, 
    0.1661563, 0.07273264, 0.07436118, 0.04360607, 0.03628521, 0.0168863, 
    0.006062986, 0.0006667653, 1.45899e-06, -1.029006e-07, 0.001239274, 
    0.02981735, 0.01180764, 0.003402752, 0.01191803, 0.0003248884, 
    4.524099e-07,
  9.062581e-05, 0.1867194, 0.05937026, 0.01899047, 0.009856851, 0.03250619, 
    0.0546882, 0.06407771, 0.08222303, 0.1741012, 0.03217422, 0.02086551, 
    0.03229543, 0.02120087, 0.01362755, 0.007723778, 0.002749109, 
    0.0006062376, 8.694087e-05, 2.450416e-05, 0.000229738, 0.006291241, 
    0.06347387, 0.05700698, 0.08973879, 0.001399173, 0.005533355, 
    6.155699e-05, 0.0001361129,
  0.05137887, 0.04392551, 0.03024796, 0.2071013, 0.02301032, 0.01024016, 
    0.07748267, 0.03573997, 0.04100494, 0.07041425, 0.01758343, 0.0250904, 
    0.04858591, 0.04585005, 0.05847152, 0.09155621, 0.1125246, 0.1520199, 
    0.1688741, 0.2774399, 0.1991654, 0.1591281, 0.1726112, 0.03818154, 
    0.02433253, 0.03805718, 0.07941931, 0.063439, 0.1038588,
  1.128851e-05, 3.506237e-06, 0.008755147, -6.708402e-06, -1.989948e-07, 
    -6.197961e-07, 0.1196965, 0.08551839, 0.2011468, 0.07533132, 0.0955383, 
    0.05845786, 0.0504709, 0.03171281, 0.02306385, 0.0409492, 0.01792145, 
    0.008062034, 0.001810266, 0.08100677, 0.04712075, 0.1662362, 0.01750726, 
    0.02973363, 0.02596982, 0.04902476, 0.02611804, 3.194085e-05, 0.0001910251,
  5.363264e-06, 0.0001799789, 0.00052148, 1.142438e-07, 1.033604e-06, 
    1.557459e-07, 0.003046889, 0.3094688, 0.3598052, 0.1805414, 0.06473124, 
    0.08837982, 0.042086, 0.03184215, 0.04617926, 0.03623625, 0.03383167, 
    0.02731615, 0.000218745, 0.0001786819, 0.05572722, 0.05513026, 
    0.05897211, 0.05004234, 0.02244649, 0.03499964, 0.0258153, 0.009422284, 
    0.001822979,
  0.02770865, 0.01098993, 0.01002396, 0.04221956, 0.006828585, 0.004023006, 
    0.08338657, 0.006463748, 0.01572086, 0.08552321, 0.07134537, 0.1056227, 
    0.08330166, 0.1627526, 0.1202438, 0.2190404, 0.1561041, 0.08263806, 
    0.04186737, 0.002276356, 0.02694498, 0.07518701, 0.07805744, 0.06114403, 
    0.06522327, 0.08554627, 0.0722613, 0.07872625, 0.0603562,
  0.1060088, 0.1804494, 0.156125, 0.1972959, 0.0862506, 0.1014241, 0.126372, 
    0.2039872, 0.1547368, 0.1577386, 0.1808574, 0.236526, 0.2405561, 
    0.2172633, 0.1753359, 0.2121172, 0.1965921, 0.1896676, 0.147742, 
    0.115212, 0.1126914, 0.05465925, 0.2342252, 0.2533319, 0.2143364, 
    0.1499058, 0.1762717, 0.2060752, 0.13501,
  0.194353, 0.2122712, 0.2014786, 0.2260874, 0.2624344, 0.1814884, 0.1963572, 
    0.259496, 0.2483301, 0.216236, 0.1998666, 0.2084173, 0.2354436, 
    0.2409669, 0.2069287, 0.2494849, 0.2534773, 0.4323323, 0.2720378, 
    0.1735481, 0.1462665, 0.2801979, 0.1759941, 0.3537757, 0.3546706, 
    0.2965113, 0.2313349, 0.1963299, 0.2309112,
  0.3388517, 0.2401393, 0.3193125, 0.2785808, 0.2754557, 0.242196, 0.2310406, 
    0.2847554, 0.2380979, 0.2594136, 0.3589527, 0.3593022, 0.2329447, 
    0.2505902, 0.3536493, 0.2642438, 0.3372416, 0.2671182, 0.188013, 
    0.2363316, 0.1821418, 0.1445324, 0.2301332, 0.3383991, 0.2623593, 
    0.3555645, 0.2042359, 0.1355148, 0.2484,
  0.2209311, 0.2193173, 0.1898413, 0.1907889, 0.2517821, 0.2617549, 
    0.2208866, 0.2659387, 0.3087118, 0.3235507, 0.3028685, 0.2843891, 
    0.2561416, 0.2143693, 0.2500076, 0.3904978, 0.3612173, 0.2837852, 
    0.331526, 0.3696049, 0.2788651, 0.2828245, 0.3225878, 0.2983404, 
    0.2603402, 0.2740878, 0.2150081, 0.1530307, 0.2600569,
  0.03917853, 0.03258736, 0.0259962, 0.01940504, 0.01281387, 0.006222705, 
    -0.0003684596, 0.01254012, 0.01288152, 0.01322292, 0.01356432, 
    0.01390573, 0.01424713, 0.01458853, -0.003237842, 0.004150103, 
    0.01153805, 0.01892599, 0.02631394, 0.03370188, 0.04108983, 0.06418753, 
    0.06304934, 0.06191116, 0.06077297, 0.05963479, 0.05849661, 0.05735843, 
    0.04445146,
  0.1434845, 0.06105592, 0.03414427, 0.01568282, 0.003915498, 0.0002732708, 
    4.893649e-06, -9.557181e-07, 0, 9.04249e-05, 0.005225695, 0.03631523, 
    0.1042475, 0.1350215, 0.1078324, 0.1339934, 0.2420543, 0.3165401, 
    0.2811877, 0.2483685, 0.2662652, 0.3157215, 0.2881704, 0.3248044, 
    0.2612175, 0.1813799, 0.2593555, 0.225798, 0.207602,
  0.1807716, 0.2241158, 0.2334034, 0.2432243, 0.2163528, 0.09195219, 
    0.1437454, 0.206879, 0.2669397, 0.2774721, 0.2675229, 0.2938297, 
    0.2770253, 0.3127552, 0.2990394, 0.2938421, 0.2630826, 0.2452624, 
    0.334224, 0.3104205, 0.2499372, 0.2824069, 0.3139511, 0.4263249, 
    0.3458217, 0.2845304, 0.2622484, 0.1936137, 0.2237918,
  0.2499135, 0.2470314, 0.2703664, 0.2835243, 0.3404617, 0.2887094, 
    0.3462591, 0.2897763, 0.3186381, 0.3375586, 0.306678, 0.3311748, 
    0.2748446, 0.3085665, 0.3039788, 0.315362, 0.2957276, 0.2867739, 
    0.2919475, 0.2568711, 0.2679192, 0.2688321, 0.3301108, 0.2301033, 
    0.2364281, 0.2040731, 0.2197168, 0.2614061, 0.2739246,
  0.2511505, 0.2496738, 0.2278961, 0.1950975, 0.2023827, 0.2401927, 
    0.2815413, 0.2990935, 0.2515187, 0.2904702, 0.2946224, 0.2170911, 
    0.1781321, 0.1879108, 0.1938496, 0.2019965, 0.1991631, 0.2387491, 
    0.2480773, 0.2665076, 0.2279681, 0.2298929, 0.2282681, 0.1803603, 
    0.1211006, 0.1614033, 0.1652318, 0.2207473, 0.2274506,
  0.1975468, 0.1667234, 0.1424921, 0.1097332, 0.1322138, 0.1721028, 
    0.1523508, 0.1567527, 0.1439784, 0.1340927, 0.0981565, 0.09575307, 
    0.0703872, 0.1427647, 0.1234712, 0.1225888, 0.1316162, 0.1117713, 
    0.1703259, 0.1493163, 0.1707164, 0.1781775, 0.1997906, 0.1977651, 
    0.03388933, 0.1284453, 0.1432344, 0.1939019, 0.2226745,
  0.02688327, 0.001209687, 0.02238772, 0.04105997, 0.03654592, 0.04295654, 
    0.02579424, 0.03294734, 0.02728045, 0.03125148, 0.004159758, 0.012503, 
    0.06701404, 0.1001133, 0.1024825, 0.125207, 0.1137901, 0.1127042, 
    0.1403504, 0.1056031, 0.09329977, 0.1182182, 0.04715946, 0.0006628102, 
    0.03357411, 0.08336645, 0.0909962, 0.07241992, 0.07844968,
  -2.276786e-07, 0.0003686135, 0.02487663, 0.002900567, 0.04840557, 
    0.06478371, 0.06989495, 0.0113116, 0.0087906, 2.715042e-05, 2.757143e-06, 
    0.0008154749, 0.01299033, 0.08187678, 0.075355, 0.04302717, 0.04113281, 
    0.09526673, 0.06109729, 0.04944691, 0.02707483, 0.005752457, 
    1.379907e-05, 1.03449e-05, 0.006897748, 0.01087555, 0.03847365, 
    0.01060077, 0.005033723,
  8.223178e-08, 0.0002583411, 0.004147482, 0.1075414, 0.02935041, 0.0218325, 
    0.05959506, 0.09368937, 0.01182891, 0.008118331, 0.02769028, 0.02785591, 
    0.1688681, 0.0715948, 0.06121755, 0.03733598, 0.03239478, 0.02031539, 
    0.01111856, 0.01240439, 0.0001243979, 5.475641e-07, 0.0004273515, 
    0.02552951, 0.01002866, 0.000170905, 0.02540594, 0.0004617308, 
    6.057082e-07,
  0.0002363443, 0.1823908, 0.04880023, 0.02050367, 0.01468231, 0.03012096, 
    0.04732396, 0.05699975, 0.07723759, 0.181225, 0.03189675, 0.02006595, 
    0.02645384, 0.0207248, 0.01330637, 0.01221368, 0.01257347, 0.005286783, 
    0.001606378, 8.685076e-05, 0.0008282363, 0.005107966, 0.04184482, 
    0.05202245, 0.04443257, 0.00148821, 0.009674292, 0.0004798013, 
    5.375992e-05,
  0.0381708, 0.04181547, 0.02588412, 0.149581, 0.005364419, 0.008825793, 
    0.07745355, 0.03301758, 0.03157971, 0.05660449, 0.02579761, 0.02785846, 
    0.04224192, 0.03883436, 0.04938186, 0.08004697, 0.1121151, 0.1445851, 
    0.1797925, 0.2716955, 0.1985273, 0.1484337, 0.1745438, 0.04312588, 
    0.02269974, 0.03158151, 0.06718151, 0.05580821, 0.09174601,
  -1.834084e-07, 1.280424e-06, 0.00241661, -7.666984e-06, -2.337028e-07, 
    4.098099e-06, 0.09663554, 0.08052421, 0.2085568, 0.07638594, 0.09310091, 
    0.05590302, 0.04391824, 0.02944315, 0.02212042, 0.03566016, 0.0462578, 
    0.01625623, 0.00650426, 0.09639144, 0.04501904, 0.1678182, 0.01699246, 
    0.02260408, 0.02549528, 0.05205262, 0.01844187, 2.031654e-05, 6.686839e-05,
  2.360159e-06, 4.500719e-05, 0.0004139489, 7.592053e-08, 5.577425e-07, 
    6.830494e-08, 0.001222594, 0.2517336, 0.3477178, 0.1774782, 0.06137509, 
    0.09169275, 0.04510149, 0.03992166, 0.05022689, 0.03245988, 0.04731338, 
    0.04697675, 0.003741814, 0.0004985869, 0.03935156, 0.04859878, 0.050574, 
    0.0486988, 0.02549597, 0.03733857, 0.0376464, 0.01383964, 0.0004394013,
  0.01835801, 0.009452856, 0.009950077, 0.05254716, 0.002666154, 0.001586839, 
    0.07268041, 0.002629553, 0.01094927, 0.08935802, 0.08328071, 0.1079407, 
    0.08884956, 0.1720199, 0.1398661, 0.2364879, 0.1657391, 0.1015907, 
    0.03455558, 0.001244651, 0.01656824, 0.0414753, 0.08394028, 0.06282253, 
    0.0729617, 0.08364034, 0.0790152, 0.08581744, 0.04886505,
  0.1014165, 0.1940203, 0.1421786, 0.1774841, 0.07605751, 0.0981771, 
    0.1188767, 0.1991866, 0.1408631, 0.1620538, 0.1983576, 0.2604592, 
    0.2177931, 0.2335342, 0.1850608, 0.2371016, 0.2324107, 0.1851717, 
    0.1394245, 0.1289342, 0.1116145, 0.08184826, 0.2121757, 0.3094811, 
    0.1853112, 0.1614416, 0.1894066, 0.2267547, 0.1380159,
  0.2097883, 0.2129238, 0.2103345, 0.2340632, 0.248522, 0.1861085, 0.2225133, 
    0.220854, 0.2360568, 0.2547424, 0.1895702, 0.1945183, 0.2463266, 
    0.254231, 0.2118743, 0.2620727, 0.2880515, 0.4429691, 0.3016355, 
    0.1725062, 0.1443521, 0.2575426, 0.1854225, 0.3524384, 0.358513, 
    0.2661198, 0.2443007, 0.2108409, 0.2539454,
  0.3214436, 0.2994163, 0.3084016, 0.2369354, 0.2389063, 0.2563937, 
    0.2370385, 0.3084783, 0.237931, 0.2490277, 0.3556826, 0.3390427, 
    0.2205555, 0.2742147, 0.2370223, 0.2486744, 0.270143, 0.2710176, 
    0.1817719, 0.2325979, 0.1900229, 0.1707768, 0.2612616, 0.3356391, 
    0.2411221, 0.3457078, 0.1835084, 0.1419792, 0.2113508,
  0.1959645, 0.2129967, 0.1550671, 0.1566483, 0.2464324, 0.2048692, 
    0.2043802, 0.246276, 0.2782914, 0.3224862, 0.2428981, 0.2141231, 
    0.2412916, 0.2407945, 0.2296076, 0.3639591, 0.3234137, 0.2874656, 
    0.312085, 0.3100352, 0.2631603, 0.26663, 0.2909261, 0.3048402, 0.2587951, 
    0.3167688, 0.2045751, 0.156625, 0.2121501,
  0.1213749, 0.1112122, 0.1010495, 0.09088679, 0.08072407, 0.07056135, 
    0.06039863, 0.06443267, 0.06584486, 0.06725706, 0.06866926, 0.07008146, 
    0.07149366, 0.07290586, 0.05443146, 0.06620253, 0.07797359, 0.08974466, 
    0.1015157, 0.1132868, 0.1250578, 0.1718337, 0.1688131, 0.1657926, 
    0.162772, 0.1597515, 0.1567309, 0.1537104, 0.1295051,
  0.1711613, 0.07861319, 0.05565824, 0.03169759, 0.004173213, -0.0001722278, 
    0.001931222, -3.063577e-05, -3.555952e-06, 0.00011523, 0.006737018, 
    0.06557356, 0.1643698, 0.134728, 0.111766, 0.129141, 0.2712778, 
    0.3118476, 0.2803142, 0.2375126, 0.3169533, 0.3423423, 0.2957038, 
    0.3251994, 0.2593186, 0.1822161, 0.2664967, 0.2261235, 0.2216873,
  0.1943351, 0.2319981, 0.243529, 0.2322613, 0.216023, 0.08557612, 0.1390087, 
    0.2429397, 0.286669, 0.2892935, 0.2678346, 0.2742844, 0.2765391, 
    0.3183796, 0.3141679, 0.2740669, 0.2594205, 0.2490997, 0.3436419, 
    0.3331302, 0.2555071, 0.2890776, 0.3189363, 0.4276751, 0.335249, 
    0.2886636, 0.2992084, 0.2391797, 0.2176188,
  0.2834424, 0.2397308, 0.2767537, 0.3294933, 0.3723969, 0.3219675, 
    0.3730319, 0.3371754, 0.3593558, 0.4043587, 0.3504781, 0.3422979, 
    0.2925765, 0.3487498, 0.3189792, 0.3267622, 0.3477434, 0.3323385, 
    0.3152398, 0.3005427, 0.2857537, 0.3035613, 0.3626554, 0.259408, 
    0.2592302, 0.2292148, 0.262398, 0.2755246, 0.2969169,
  0.2954124, 0.2818518, 0.2625131, 0.2408321, 0.2324604, 0.2754604, 
    0.2875211, 0.3137327, 0.2769536, 0.3085797, 0.2918063, 0.2438096, 
    0.2119997, 0.2503401, 0.2324451, 0.2549095, 0.2802882, 0.3209884, 
    0.3022966, 0.3232645, 0.265492, 0.2418597, 0.2815997, 0.2059298, 
    0.1285513, 0.1482243, 0.1868042, 0.2499354, 0.2509675,
  0.2200726, 0.2030305, 0.1651228, 0.1625322, 0.1701067, 0.1927339, 
    0.1674818, 0.2057676, 0.1926389, 0.1988701, 0.1121935, 0.115742, 
    0.06011878, 0.1818116, 0.1396607, 0.1554922, 0.16461, 0.1579629, 
    0.2070244, 0.200792, 0.2046356, 0.2010248, 0.2178355, 0.2198513, 
    0.04330821, 0.1559771, 0.186651, 0.2270993, 0.2696856,
  0.05362944, 0.02024782, 0.01794415, 0.05769318, 0.05613438, 0.06065995, 
    0.04810726, 0.0634369, 0.05777471, 0.05453314, 0.003064163, 0.008910296, 
    0.04211136, 0.1139271, 0.1216277, 0.1302574, 0.1454846, 0.1450363, 
    0.1556233, 0.1263835, 0.1466813, 0.1497824, 0.084817, 0.0003952879, 
    0.02842952, 0.09165221, 0.1099981, 0.09409182, 0.1020579,
  -7.13699e-06, 0.0002850941, 0.01405672, 0.002362917, 0.04062877, 
    0.07139257, 0.09317359, 0.02727941, 0.03304695, 0.0001021173, 
    1.442802e-07, 8.247443e-05, 0.04089818, 0.08943015, 0.09287471, 
    0.04763888, 0.05241133, 0.1033262, 0.0494458, 0.04632249, 0.08102369, 
    0.02977525, 0.0005010284, 6.840318e-06, 0.002264081, 0.00488578, 
    0.05330472, 0.05148074, 0.009380138,
  1.304441e-06, -5.205979e-05, 0.0007508501, 0.07216623, 0.02873353, 
    0.02769804, 0.06558787, 0.08894812, 0.01397161, 0.01068802, 0.02814066, 
    0.03886136, 0.1783985, 0.07689247, 0.04720419, 0.0326732, 0.02851735, 
    0.02266208, 0.01316996, 0.02882811, 0.009821842, 7.147318e-05, 
    9.059038e-07, 0.02591308, 0.009774219, 3.60931e-05, 0.04481709, 
    0.005783976, 1.766586e-06,
  0.001392511, 0.1829635, 0.0415085, 0.02345224, 0.02014749, 0.02841859, 
    0.03951059, 0.0480005, 0.07308646, 0.1929757, 0.0311559, 0.01794456, 
    0.02327652, 0.01934612, 0.01487596, 0.01260644, 0.01967699, 0.01220405, 
    0.01002934, 0.003237945, 0.001440121, 0.00191782, 0.02014439, 0.05098187, 
    0.02468032, 0.002188187, 0.01632368, 0.004136217, 0.0001055299,
  0.03300584, 0.04116868, 0.02142633, 0.1112301, 0.001225046, 0.009152762, 
    0.07055634, 0.02890322, 0.02344903, 0.04234416, 0.03634865, 0.02833142, 
    0.0345805, 0.03123169, 0.04088988, 0.06650187, 0.1073957, 0.141059, 
    0.1774806, 0.2571244, 0.1863351, 0.1348289, 0.1729679, 0.05075905, 
    0.02200127, 0.02984731, 0.05871293, 0.05195423, 0.08202457,
  -3.265168e-07, 5.293942e-07, 0.0009515632, 7.946381e-05, -2.207351e-07, 
    -6.747581e-06, 0.08018993, 0.07248555, 0.2259743, 0.0743596, 0.08288072, 
    0.04770708, 0.03711621, 0.02883806, 0.02234755, 0.02967753, 0.05193251, 
    0.06983868, 0.007221739, 0.1151062, 0.04978491, 0.169773, 0.01734122, 
    0.01755484, 0.02536173, 0.04938675, 0.01778152, 1.207975e-05, 3.413058e-05,
  1.375597e-06, 4.340124e-06, 2.442136e-05, 5.505883e-08, 3.627917e-07, 
    2.834668e-08, 0.0002657179, 0.2037305, 0.3650646, 0.1630189, 0.05995058, 
    0.08591662, 0.04679428, 0.03719923, 0.05162911, 0.04308248, 0.05201516, 
    0.07620095, 0.008818541, 0.001225265, 0.0337024, 0.03558331, 0.05282617, 
    0.04813436, 0.03844875, 0.03694094, 0.05173561, 0.02343963, 1.218531e-05,
  0.01403314, 0.01021314, 0.008332351, 0.0671199, 0.001998648, 0.0001347038, 
    0.06423524, 0.0008056122, 0.006496941, 0.07890958, 0.08156617, 0.1042113, 
    0.09773585, 0.1737682, 0.1765817, 0.2523285, 0.2061256, 0.134723, 
    0.04427933, 0.0006108679, 0.01341107, 0.02557938, 0.08763305, 0.09831899, 
    0.09471924, 0.1113436, 0.104238, 0.09514657, 0.04936461,
  0.1129075, 0.1662057, 0.1545108, 0.1999121, 0.0733217, 0.09254464, 
    0.0947689, 0.2142622, 0.1396169, 0.155241, 0.1995538, 0.2409361, 
    0.2154091, 0.2695964, 0.2130002, 0.2511778, 0.2535258, 0.2051024, 
    0.1676109, 0.1275494, 0.110612, 0.07971793, 0.2115137, 0.3532327, 
    0.1952421, 0.1832736, 0.2124797, 0.241679, 0.1442063,
  0.222369, 0.2052092, 0.1912346, 0.2385741, 0.2198533, 0.1869799, 0.1871581, 
    0.1999452, 0.2233631, 0.2823237, 0.2050976, 0.2465897, 0.2647218, 
    0.2419368, 0.2282701, 0.2998477, 0.3110411, 0.4581761, 0.3166702, 
    0.1740916, 0.1646053, 0.2984564, 0.2399817, 0.4080939, 0.3904541, 
    0.2329416, 0.3099839, 0.260761, 0.2662242,
  0.3657474, 0.3150508, 0.3207929, 0.2605292, 0.2824204, 0.2051135, 
    0.2542297, 0.3155577, 0.2539337, 0.2677712, 0.3767031, 0.3910815, 
    0.2211482, 0.329535, 0.2407846, 0.2519287, 0.2807307, 0.2772719, 
    0.1939518, 0.2619765, 0.206302, 0.2381797, 0.2836311, 0.3518597, 
    0.2265582, 0.3246672, 0.2099499, 0.1270105, 0.2669324,
  0.1850989, 0.1977324, 0.1568952, 0.1671267, 0.2435889, 0.2000478, 
    0.2287923, 0.2603845, 0.2724745, 0.2675831, 0.2849878, 0.2429832, 
    0.2993946, 0.3219927, 0.2697972, 0.3352343, 0.3031558, 0.3063172, 
    0.3578641, 0.330669, 0.2378041, 0.2744085, 0.2827675, 0.3058191, 
    0.2902368, 0.3085239, 0.2273048, 0.1590723, 0.1909989,
  0.1951121, 0.186414, 0.177716, 0.1690179, 0.1603199, 0.1516218, 0.1429238, 
    0.1468352, 0.1507186, 0.154602, 0.1584854, 0.1623688, 0.1662522, 
    0.1701356, 0.1521343, 0.1609326, 0.1697309, 0.1785292, 0.1873275, 
    0.1961258, 0.2049241, 0.227042, 0.2230583, 0.2190746, 0.215091, 
    0.2111073, 0.2071236, 0.2031399, 0.2020705,
  0.1928088, 0.1081057, 0.07449674, 0.03673007, 0.007604667, -0.0007183034, 
    0.003142192, 0.0003480726, 0.001599986, 0.006356436, 0.01077659, 
    0.1202895, 0.1921048, 0.1248837, 0.1207103, 0.1342229, 0.263792, 
    0.3207531, 0.3002343, 0.22957, 0.3254432, 0.3507724, 0.3018674, 
    0.3123254, 0.2537887, 0.1898249, 0.2605059, 0.2250832, 0.2341958,
  0.2029628, 0.2259854, 0.2382673, 0.2131683, 0.2026676, 0.08270422, 
    0.1238143, 0.2617976, 0.290284, 0.2983815, 0.2602801, 0.2555873, 
    0.2745197, 0.2957896, 0.3279999, 0.2727129, 0.244501, 0.2524188, 
    0.3381099, 0.3694456, 0.2521485, 0.3219217, 0.338107, 0.4505152, 
    0.3218257, 0.2967444, 0.3349277, 0.2443751, 0.2455249,
  0.2902384, 0.2532194, 0.3235277, 0.4320933, 0.4438227, 0.351596, 0.3634565, 
    0.3576929, 0.4255157, 0.4209102, 0.3631885, 0.3355519, 0.3057683, 
    0.3510033, 0.3331837, 0.3558346, 0.3639414, 0.4131459, 0.3856409, 
    0.3187914, 0.3492557, 0.3319311, 0.4033612, 0.337895, 0.3042938, 
    0.2624426, 0.3020321, 0.2844867, 0.3096309,
  0.3453451, 0.3163232, 0.3445675, 0.2761694, 0.274236, 0.293642, 0.3041803, 
    0.3088138, 0.2874694, 0.2976111, 0.2669414, 0.2540013, 0.2534138, 
    0.2943102, 0.2665669, 0.3041853, 0.2708078, 0.3711772, 0.3582078, 
    0.341833, 0.2984967, 0.2652726, 0.3244986, 0.2239128, 0.132109, 
    0.2096487, 0.2953542, 0.349201, 0.3041142,
  0.2990969, 0.2211816, 0.1924278, 0.2110656, 0.2333041, 0.2168324, 
    0.2134143, 0.2329129, 0.2395576, 0.2003046, 0.1477344, 0.1189649, 
    0.07905076, 0.2386982, 0.180979, 0.2230161, 0.1616459, 0.2462429, 
    0.3070898, 0.2364725, 0.2388538, 0.2140847, 0.2416384, 0.2516824, 
    0.06166175, 0.161902, 0.2305275, 0.2998321, 0.3254929,
  0.08440562, 0.03009957, 0.01684112, 0.083903, 0.07367601, 0.09579787, 
    0.08789795, 0.1137198, 0.1482329, 0.07963549, 0.003030055, 0.006186679, 
    0.03459505, 0.1351424, 0.1635207, 0.170468, 0.1755822, 0.1534944, 
    0.1894653, 0.2218383, 0.213436, 0.180532, 0.1612449, 0.001224778, 
    0.04112896, 0.1619603, 0.1840085, 0.1422906, 0.1562412,
  0.0003307527, 0.0002064724, 0.008652373, 0.006454844, 0.04435415, 
    0.07207746, 0.1377921, 0.1024135, 0.111762, 0.0002058695, 1.057186e-07, 
    5.359612e-06, 0.07067911, 0.1041574, 0.1021748, 0.0541411, 0.06880394, 
    0.1116697, 0.04898981, 0.05510728, 0.2283289, 0.2703941, 0.07516576, 
    1.219315e-06, 0.001019507, 0.005206138, 0.06891157, 0.1098592, 0.06766315,
  1.55322e-05, 3.482002e-05, 0.0001555744, 0.04295718, 0.03269098, 
    0.03259284, 0.07176047, 0.07947484, 0.02485796, 0.02279548, 0.02847262, 
    0.04798572, 0.1735439, 0.07752395, 0.03926822, 0.03328153, 0.02898895, 
    0.02661493, 0.0165809, 0.02980915, 0.07892438, 0.0101116, 1.139233e-05, 
    0.02865293, 0.009404369, 1.005002e-05, 0.06098954, 0.05953179, 
    0.0007693357,
  0.01861475, 0.1843108, 0.0367558, 0.0217742, 0.02457296, 0.03043886, 
    0.03511133, 0.04195919, 0.07241805, 0.2093523, 0.03263082, 0.01814565, 
    0.0238963, 0.0223544, 0.01881086, 0.01454867, 0.02043363, 0.01564794, 
    0.02217021, 0.02675485, 0.003417391, 0.001040722, 0.008884856, 
    0.04909574, 0.01770534, 0.006452534, 0.02149427, 0.01949357, 0.00221401,
  0.02925317, 0.03649272, 0.01468317, 0.07917653, 0.0002084224, 0.01243495, 
    0.0623, 0.02871086, 0.02051315, 0.03319435, 0.03924906, 0.03000943, 
    0.03148644, 0.02741358, 0.03620481, 0.05783867, 0.0908011, 0.120055, 
    0.1610847, 0.2311288, 0.1649604, 0.1086492, 0.1814299, 0.0493796, 
    0.02438208, 0.03001664, 0.05698496, 0.04804906, 0.07559304,
  -2.071372e-07, 2.445325e-07, 3.216115e-05, 0.000281928, -1.874252e-07, 
    -2.001128e-05, 0.06408598, 0.06234059, 0.2233168, 0.0877096, 0.08332784, 
    0.04537282, 0.03485614, 0.03064026, 0.02630108, 0.03053829, 0.05303921, 
    0.1160484, 0.03370254, 0.1274561, 0.05439394, 0.171641, 0.02187766, 
    0.0199405, 0.02988333, 0.04883241, 0.02407608, -2.695877e-06, 1.547816e-05,
  9.498954e-07, 5.2448e-06, 0.0004924507, 4.265219e-08, 2.542701e-07, 
    1.346111e-08, -2.205377e-06, 0.1803184, 0.3783165, 0.1617491, 0.07623191, 
    0.09462297, 0.05323193, 0.05274513, 0.06183246, 0.08075085, 0.06739653, 
    0.1170437, 0.05707426, 0.001256062, 0.02892759, 0.0302806, 0.0684597, 
    0.04754166, 0.03856446, 0.04317411, 0.0521419, 0.07310413, 0.0007029054,
  0.01218476, 0.009608208, 0.006969751, 0.08933677, 0.0008308199, 
    -3.864531e-05, 0.05442274, -1.00533e-05, 0.00237791, 0.06522848, 
    0.08661585, 0.1016976, 0.1175129, 0.2104005, 0.2453827, 0.3132465, 
    0.2601112, 0.1866077, 0.1053685, -0.0001310054, 0.008175581, 0.02575504, 
    0.1014856, 0.1216971, 0.1308148, 0.1273452, 0.1552294, 0.1706683, 
    0.05303266,
  0.1307201, 0.1856063, 0.1539606, 0.1878822, 0.05379036, 0.0526706, 
    0.0794278, 0.2131673, 0.1498444, 0.1333922, 0.1521877, 0.2288204, 
    0.240739, 0.2861157, 0.2856231, 0.3008058, 0.2782522, 0.2229739, 
    0.1795973, 0.1245417, 0.09921568, 0.05799156, 0.2044868, 0.3412333, 
    0.1917326, 0.2010417, 0.2634582, 0.2741455, 0.1612442,
  0.2632113, 0.2217319, 0.2287448, 0.2472343, 0.2394829, 0.2182793, 
    0.1751772, 0.2258541, 0.2197179, 0.2952103, 0.2530857, 0.3381962, 
    0.2933675, 0.3146251, 0.2683048, 0.3757805, 0.3400657, 0.4749259, 
    0.3241241, 0.1769027, 0.1973871, 0.3094897, 0.3191063, 0.4907129, 
    0.4280574, 0.2205655, 0.3515864, 0.3088295, 0.2678243,
  0.425976, 0.3453422, 0.3759169, 0.3193132, 0.341225, 0.2606203, 0.3373109, 
    0.336159, 0.2684451, 0.3516088, 0.4237585, 0.4288676, 0.2988651, 
    0.3505588, 0.3443798, 0.2683164, 0.3596459, 0.3060631, 0.2540456, 
    0.3198486, 0.3061628, 0.3336404, 0.335536, 0.3474858, 0.2547495, 
    0.3208982, 0.2281159, 0.1382548, 0.4081695,
  0.1969433, 0.2491952, 0.215323, 0.2083118, 0.2815795, 0.2275431, 0.2580539, 
    0.2798437, 0.4011386, 0.3347519, 0.3520424, 0.3578363, 0.3748994, 
    0.3446078, 0.382571, 0.3738519, 0.4088122, 0.3698559, 0.409224, 
    0.3923014, 0.2993541, 0.3033663, 0.3043856, 0.315381, 0.2499625, 
    0.3040589, 0.2304032, 0.1893927, 0.2189193,
  0.2252364, 0.2185184, 0.2118005, 0.2050825, 0.1983646, 0.1916466, 
    0.1849287, 0.1908921, 0.196694, 0.2024958, 0.2082976, 0.2140994, 
    0.2199013, 0.2257031, 0.23205, 0.2372765, 0.2425031, 0.2477297, 
    0.2529563, 0.2581829, 0.2634094, 0.246283, 0.2419725, 0.2376621, 
    0.2333516, 0.2290412, 0.2247307, 0.2204203, 0.2306107,
  0.2156706, 0.1283169, 0.08776911, 0.04318815, 0.01557702, -0.001220985, 
    0.001490046, 0.002673762, 0.002139498, 0.006945495, 0.03223624, 
    0.1503941, 0.2096138, 0.1182278, 0.1326202, 0.1543233, 0.2667013, 
    0.3258752, 0.303102, 0.2389508, 0.3507884, 0.3476583, 0.2943254, 
    0.2876507, 0.2518879, 0.1934766, 0.2506382, 0.2125817, 0.2449509,
  0.207159, 0.2257005, 0.2274632, 0.1945985, 0.182249, 0.08151168, 0.1094109, 
    0.2749383, 0.2943265, 0.302501, 0.2581106, 0.2176412, 0.2533187, 
    0.2593141, 0.3199009, 0.3047283, 0.2709653, 0.2592151, 0.3373895, 
    0.3667083, 0.2993736, 0.3588562, 0.3420358, 0.4791186, 0.318812, 
    0.3053173, 0.3180178, 0.2763007, 0.2483976,
  0.3095613, 0.3431898, 0.4504934, 0.4594601, 0.4599719, 0.3760066, 
    0.3547311, 0.3785115, 0.4563568, 0.3710277, 0.2961919, 0.3373762, 
    0.386424, 0.343956, 0.2987196, 0.3557753, 0.3806489, 0.4615834, 
    0.3812202, 0.3271312, 0.3676793, 0.3000318, 0.3894811, 0.3295092, 
    0.3582082, 0.2960998, 0.3221902, 0.3294802, 0.3196156,
  0.3466106, 0.3318236, 0.3517769, 0.2857034, 0.3322475, 0.3100288, 
    0.2984744, 0.2776874, 0.2733706, 0.2825197, 0.2735593, 0.2620989, 
    0.2108142, 0.2498263, 0.2435166, 0.2695885, 0.2788491, 0.3509945, 
    0.3410628, 0.3791575, 0.3229263, 0.2817288, 0.327799, 0.2406228, 
    0.1517549, 0.2774818, 0.3760578, 0.4233619, 0.3890072,
  0.2802989, 0.2282418, 0.1907922, 0.2461782, 0.2792359, 0.2571294, 
    0.2164864, 0.2507268, 0.2495266, 0.2102046, 0.1235731, 0.1094849, 
    0.05130167, 0.2263187, 0.228608, 0.2344282, 0.1938725, 0.2348442, 
    0.2601909, 0.2074136, 0.2026922, 0.1745617, 0.2137895, 0.2977574, 
    0.07333137, 0.1581081, 0.2320142, 0.3238795, 0.3188945,
  0.1904577, 0.05173267, 0.01557406, 0.09237481, 0.08208233, 0.191782, 
    0.1640503, 0.1935725, 0.2270369, 0.06866534, 0.006099591, 0.003535225, 
    0.03267758, 0.1669493, 0.1916881, 0.2345925, 0.1509899, 0.1728352, 
    0.2242274, 0.1952965, 0.1890361, 0.2550409, 0.1997481, 0.003292635, 
    0.05199513, 0.1624548, 0.2543598, 0.2110884, 0.1814136,
  0.09679393, 7.267092e-05, 0.008446915, 0.01507314, 0.06059728, 0.07400852, 
    0.1465632, 0.173552, 0.1799336, 0.004035003, 2.610619e-08, 1.50874e-06, 
    0.09470034, 0.1286984, 0.1100213, 0.06594308, 0.08486679, 0.129009, 
    0.05880889, 0.08507749, 0.3185311, 0.5306457, 0.3966503, -4.54378e-06, 
    0.008204036, 0.01588451, 0.07816723, 0.186287, 0.2974034,
  0.003378009, 0.003093734, 5.980134e-05, 0.02427898, 0.04758491, 0.0629163, 
    0.0832465, 0.07797753, 0.05199336, 0.0460484, 0.03044062, 0.06145983, 
    0.1561615, 0.07940999, 0.03879464, 0.04364296, 0.03790614, 0.04791129, 
    0.03844101, 0.05320299, 0.1723934, 0.1295149, 0.0009836366, 0.02216029, 
    0.00654162, 4.019044e-06, 0.08524568, 0.1602927, 0.04290976,
  0.0995717, 0.1817962, 0.03020905, 0.02746077, 0.03335737, 0.03977329, 
    0.03828437, 0.04184037, 0.06537395, 0.198865, 0.03851957, 0.02618184, 
    0.02985467, 0.04198803, 0.04949498, 0.04157797, 0.02794317, 0.01380419, 
    0.02542236, 0.04638042, 0.03865995, 0.003508843, 0.001672552, 0.0364299, 
    0.008054622, 0.01887848, 0.04865347, 0.03814989, 0.02870297,
  0.02299401, 0.03086407, 0.009711243, 0.05760173, 4.407721e-05, 0.02126359, 
    0.05676261, 0.03686299, 0.0168704, 0.03156483, 0.02859889, 0.03405871, 
    0.04039473, 0.03042597, 0.03765516, 0.05549302, 0.08764349, 0.1072679, 
    0.1535364, 0.1945663, 0.134646, 0.09945095, 0.1640693, 0.04281408, 
    0.04988185, 0.04059173, 0.06154175, 0.04696681, 0.06232847,
  -2.695212e-08, 1.451403e-07, -9.210002e-06, 0.0001958951, -1.346614e-07, 
    0.0004614919, 0.04475014, 0.05622826, 0.2159357, 0.08185823, 0.09475829, 
    0.04442449, 0.03777214, 0.03838852, 0.03698161, 0.03948536, 0.06939279, 
    0.1267827, 0.1960685, 0.1475942, 0.05540829, 0.1734885, 0.0338562, 
    0.02275233, 0.04835784, 0.06827376, 0.04864104, 0.0001195774, 1.131581e-05,
  7.060974e-07, -4.728311e-05, 0.001273132, 3.485924e-08, 1.928045e-07, 
    8.24773e-09, -9.383347e-05, 0.1834635, 0.3932168, 0.1473637, 0.1201566, 
    0.07694508, 0.06053343, 0.04675535, 0.08539238, 0.08514662, 0.1031843, 
    0.1401495, 0.2081096, 0.0009842073, 0.01797869, 0.02883036, 0.06788132, 
    0.05275595, 0.04276923, 0.05434045, 0.06390188, 0.1332713, 0.001000783,
  0.01000041, 0.01090255, 0.002046587, 0.1073782, 0.001011774, -2.999293e-05, 
    0.04951748, -0.0001266839, 0.003485364, 0.04565807, 0.08841363, 
    0.09679464, 0.1470704, 0.2520592, 0.2658859, 0.3088145, 0.2643894, 
    0.2277077, 0.1978344, -6.471357e-05, 0.005712067, 0.02277187, 0.1253921, 
    0.1179166, 0.139311, 0.15968, 0.2052267, 0.2438226, 0.06863617,
  0.1237649, 0.2098336, 0.1987044, 0.1881867, 0.05350204, 0.03080274, 
    0.06907298, 0.2115863, 0.1292536, 0.133365, 0.1396316, 0.2084896, 
    0.293072, 0.288088, 0.3264594, 0.3191527, 0.2723791, 0.2706367, 
    0.2466675, 0.1229888, 0.07360441, 0.03946798, 0.1787419, 0.312078, 
    0.1906917, 0.2141342, 0.3042057, 0.2856802, 0.1798633,
  0.2635817, 0.2361807, 0.2423695, 0.2453453, 0.2528414, 0.1918868, 
    0.1697322, 0.1733906, 0.2251574, 0.2756784, 0.2299224, 0.341119, 
    0.2714936, 0.3438844, 0.3085551, 0.4392048, 0.3875198, 0.4642935, 
    0.303013, 0.1609571, 0.2414852, 0.3232375, 0.3891634, 0.5720423, 
    0.4032747, 0.224056, 0.3674642, 0.34577, 0.2884052,
  0.5347744, 0.354484, 0.3964396, 0.3835983, 0.4200199, 0.3080596, 0.3639268, 
    0.3945873, 0.2912726, 0.3447883, 0.4551296, 0.3891775, 0.4089782, 
    0.4199914, 0.4060994, 0.3651935, 0.4188094, 0.3878252, 0.3662704, 
    0.3958443, 0.3380153, 0.3922388, 0.3497646, 0.3634599, 0.3150179, 
    0.3404754, 0.2270781, 0.1619002, 0.4599569,
  0.2679272, 0.3256769, 0.3266959, 0.3249779, 0.3485104, 0.3435943, 
    0.3502916, 0.3687497, 0.4545061, 0.4196598, 0.3998592, 0.3748301, 
    0.3893088, 0.4273799, 0.4374208, 0.492457, 0.4415141, 0.4010563, 
    0.4439419, 0.4233954, 0.3204893, 0.3131693, 0.3291671, 0.3251218, 
    0.2513669, 0.3415896, 0.2414801, 0.2188413, 0.2720211,
  0.2395736, 0.2340011, 0.2284286, 0.2228561, 0.2172837, 0.2117112, 
    0.2061387, 0.2040376, 0.2111001, 0.2181625, 0.225225, 0.2322875, 
    0.2393499, 0.2464124, 0.2754536, 0.2785833, 0.2817129, 0.2848425, 
    0.2879722, 0.2911018, 0.2942314, 0.2636922, 0.2590726, 0.254453, 
    0.2498334, 0.2452138, 0.2405942, 0.2359746, 0.2440316,
  0.2400474, 0.1554688, 0.1062718, 0.05176242, 0.0162116, -0.001532695, 
    0.0004041645, 0.004266083, 0.001880359, 0.005526513, 0.05770263, 
    0.1758853, 0.2009387, 0.09511228, 0.1285448, 0.1640708, 0.2451456, 
    0.340981, 0.2960405, 0.2276626, 0.3690258, 0.3448224, 0.2851574, 
    0.2670419, 0.2542538, 0.212183, 0.2185785, 0.1979376, 0.2541658,
  0.2203993, 0.1984069, 0.2207164, 0.1633335, 0.1603984, 0.07204795, 
    0.08781681, 0.2844357, 0.2947707, 0.3130295, 0.2698859, 0.1855672, 
    0.2261825, 0.2346239, 0.317428, 0.358138, 0.2935418, 0.3060902, 
    0.3619449, 0.3744955, 0.3403287, 0.3801473, 0.3551257, 0.5043327, 
    0.3279133, 0.3097202, 0.3378046, 0.3057862, 0.2702256,
  0.3535663, 0.3792453, 0.5186436, 0.3772174, 0.4181711, 0.4139863, 
    0.3434146, 0.4350273, 0.4191697, 0.2769238, 0.2371584, 0.3436315, 
    0.3652987, 0.3493869, 0.2824728, 0.359986, 0.3924962, 0.4682066, 
    0.4022358, 0.2946231, 0.3000529, 0.2723382, 0.3339444, 0.3083694, 
    0.3580299, 0.3629075, 0.3641843, 0.374313, 0.3391917,
  0.3386403, 0.3355647, 0.3166193, 0.3190978, 0.3453578, 0.3150455, 
    0.3085905, 0.2530683, 0.2555383, 0.2737579, 0.2757458, 0.2791601, 
    0.2327331, 0.2172099, 0.2229798, 0.2403982, 0.2675931, 0.3234379, 
    0.3254557, 0.370483, 0.3303932, 0.3249099, 0.3127105, 0.2401464, 
    0.1574286, 0.2463825, 0.3903161, 0.4637512, 0.3839413,
  0.2592426, 0.2065403, 0.1492887, 0.2277877, 0.2696479, 0.2612501, 
    0.2390466, 0.2460648, 0.2535433, 0.1884207, 0.1628974, 0.08727415, 
    0.03213163, 0.176416, 0.2327745, 0.2127571, 0.1787252, 0.1909344, 
    0.183372, 0.1497323, 0.1393123, 0.1230961, 0.1670104, 0.3343055, 
    0.04403096, 0.1400898, 0.226027, 0.2615349, 0.3161769,
  0.2463034, 0.1011316, 0.01110562, 0.1156443, 0.134733, 0.2319153, 
    0.2383916, 0.1829551, 0.2119611, 0.06822837, 0.00902236, 0.0009869217, 
    0.03054243, 0.1387147, 0.18134, 0.1581681, 0.1218963, 0.1622237, 
    0.1573878, 0.1557097, 0.1436072, 0.202265, 0.2694557, 0.007721143, 
    0.04895336, 0.1694569, 0.202058, 0.2159307, 0.2145529,
  0.3886753, -6.590714e-05, 0.006286164, 0.05229766, 0.05466304, 0.04542024, 
    0.08081874, 0.08975054, 0.1559514, 0.001420924, 1.538003e-08, 
    9.809685e-07, 0.06855298, 0.1414155, 0.1447008, 0.08697703, 0.08290964, 
    0.1202728, 0.06849263, 0.06444341, 0.1668179, 0.3166459, 0.5106356, 
    -0.0002269994, 0.01234485, 0.02002149, 0.1102697, 0.1508903, 0.3469635,
  0.103631, 0.03082881, 2.840784e-05, 0.01934237, 0.05401529, 0.05483839, 
    0.08736831, 0.06532285, 0.07073641, 0.05355344, 0.0316276, 0.04479747, 
    0.1654492, 0.09255987, 0.04569718, 0.04068948, 0.04765934, 0.03608484, 
    0.03218894, 0.02841573, 0.1323794, 0.4530831, 0.04561565, 0.009198743, 
    0.002462036, 4.541014e-07, 0.104512, 0.2161563, 0.4829162,
  0.1650167, 0.1594304, 0.02742848, 0.03875858, 0.06498664, 0.07651364, 
    0.05685329, 0.04532517, 0.0422373, 0.1569959, 0.06361432, 0.07574987, 
    0.06546366, 0.07010308, 0.08186442, 0.05053903, 0.04249504, 0.03315729, 
    0.04523259, 0.05368543, 0.1086265, 0.03086582, 0.007272136, 0.01611386, 
    0.002784276, 0.08807278, 0.09813521, 0.09363797, 0.1159889,
  0.014423, 0.02519039, 0.006419653, 0.04551905, -1.322314e-05, 0.04948336, 
    0.0561659, 0.04449367, 0.01490799, 0.03804513, 0.01523749, 0.1482354, 
    0.06093097, 0.06454384, 0.04257312, 0.09245357, 0.1081291, 0.1576793, 
    0.1645529, 0.1645965, 0.1283518, 0.1125494, 0.1470858, 0.03878014, 
    0.06806345, 0.1064825, 0.083674, 0.06000329, 0.04454742,
  2.232155e-08, 1.051523e-07, -2.84954e-06, 0.0005363838, -6.60076e-08, 
    0.0160306, 0.02838805, 0.05322696, 0.1639587, 0.08970445, 0.0975365, 
    0.04798596, 0.05184948, 0.06259605, 0.06896718, 0.04178172, 0.04302391, 
    0.1150361, 0.2866512, 0.2346784, 0.08898278, 0.1799054, 0.0818215, 
    0.01956107, 0.07117908, 0.1132863, 0.1443511, 0.03640039, 7.234424e-06,
  5.538007e-07, 0.0004876002, 0.000507665, 2.927974e-08, 1.581276e-07, 
    5.788086e-09, -0.0001328894, 0.1951264, 0.4093938, 0.152952, 0.1364289, 
    0.06484738, 0.07514767, 0.06846597, 0.101355, 0.1193224, 0.1263742, 
    0.1316743, 0.2456998, 0.0003284371, 0.01426721, 0.04047472, 0.05828947, 
    0.0805696, 0.0632868, 0.0976714, 0.127432, 0.1541791, 0.003288209,
  0.008600293, 0.007952698, 0.0005541645, 0.1297771, 0.0004040916, 
    -2.098596e-05, 0.04917159, -3.825548e-05, 0.001786825, 0.03358639, 
    0.08867235, 0.09954125, 0.2065356, 0.2776291, 0.2736768, 0.2986108, 
    0.2244054, 0.258154, 0.2818385, -0.0001083333, 0.00148671, 0.01654791, 
    0.114283, 0.1054332, 0.125381, 0.131169, 0.1924241, 0.1746944, 0.06877548,
  0.1086741, 0.2255057, 0.1843108, 0.1993335, 0.0371009, 0.02238486, 
    0.05449325, 0.204796, 0.1121969, 0.1319596, 0.1127021, 0.1871188, 
    0.3241743, 0.3235698, 0.3158139, 0.3022556, 0.2833435, 0.2768818, 
    0.2792404, 0.1146447, 0.06880967, 0.03068965, 0.1554935, 0.2960354, 
    0.1896783, 0.3041353, 0.3627356, 0.2789647, 0.1597579,
  0.2325525, 0.2311222, 0.2190237, 0.2078965, 0.2387683, 0.1643577, 
    0.1411845, 0.1393023, 0.2220179, 0.2518913, 0.2006011, 0.3507173, 
    0.2853428, 0.3343498, 0.3322807, 0.3751827, 0.3858016, 0.4528495, 
    0.303418, 0.152785, 0.1818252, 0.3053313, 0.4109611, 0.5179665, 
    0.4072148, 0.2274745, 0.3659414, 0.2772282, 0.2885474,
  0.5700276, 0.3218551, 0.3815709, 0.436201, 0.4299708, 0.2849755, 0.3430048, 
    0.373086, 0.2942241, 0.2553714, 0.453625, 0.3911729, 0.4144407, 
    0.4807237, 0.4266027, 0.4769713, 0.4636304, 0.4043025, 0.4298682, 
    0.3986807, 0.40168, 0.4101719, 0.3816347, 0.4071346, 0.4048485, 
    0.3598689, 0.2209353, 0.1918508, 0.5053412,
  0.412816, 0.5376177, 0.4390885, 0.4352348, 0.4407827, 0.4172868, 0.4586699, 
    0.4732398, 0.4271543, 0.4574525, 0.3940642, 0.3722445, 0.4007604, 
    0.4251493, 0.4493251, 0.4980696, 0.4625223, 0.5632046, 0.5343688, 
    0.4756297, 0.4860911, 0.319008, 0.3346866, 0.3791524, 0.2778798, 
    0.3476476, 0.2201634, 0.2307157, 0.3430249,
  0.2175003, 0.2119045, 0.2063085, 0.2007127, 0.1951168, 0.1895209, 0.183925, 
    0.1868439, 0.195198, 0.2035521, 0.2119062, 0.2202603, 0.2286144, 
    0.2369685, 0.2709782, 0.2737545, 0.2765307, 0.279307, 0.2820833, 
    0.2848596, 0.2876359, 0.2771186, 0.2715841, 0.2660496, 0.2605151, 
    0.2549806, 0.2494462, 0.2439117, 0.2219771,
  0.2783583, 0.1802773, 0.1162474, 0.060112, 0.01630667, -0.001395482, 
    -0.0002046527, 0.004358501, 0.001479713, 0.003347794, 0.05158898, 
    0.1825486, 0.2155878, 0.07173327, 0.1241134, 0.1835702, 0.2577255, 
    0.317641, 0.2602449, 0.2269797, 0.3722082, 0.351782, 0.2751155, 
    0.2471628, 0.2458496, 0.227472, 0.171098, 0.1804021, 0.2749103,
  0.2185187, 0.1671016, 0.2130125, 0.1019697, 0.1395055, 0.05597309, 
    0.05817714, 0.2947642, 0.2837543, 0.3151703, 0.2829841, 0.1651198, 
    0.1929186, 0.2101596, 0.3381988, 0.3837433, 0.3330528, 0.3701892, 
    0.4069566, 0.4304295, 0.3594004, 0.4005995, 0.387795, 0.5369902, 
    0.3118021, 0.3452646, 0.3746758, 0.3556703, 0.2950397,
  0.4138884, 0.3803319, 0.4832564, 0.2897852, 0.3324779, 0.3741231, 
    0.3378914, 0.4585074, 0.352572, 0.1969331, 0.1849717, 0.304588, 
    0.3134509, 0.3419307, 0.2891285, 0.3579868, 0.3820378, 0.430311, 
    0.3539162, 0.25518, 0.2583615, 0.2498516, 0.3362779, 0.2628039, 
    0.3306943, 0.3990863, 0.4109485, 0.4243774, 0.3663609,
  0.3100432, 0.2944967, 0.3048167, 0.3118501, 0.3299177, 0.3170606, 
    0.3253641, 0.2311675, 0.2378009, 0.2563688, 0.2586362, 0.2644473, 
    0.209138, 0.2118575, 0.1749163, 0.2259584, 0.231253, 0.2935976, 
    0.3033537, 0.3274996, 0.295266, 0.3258078, 0.289735, 0.2191656, 0.134064, 
    0.2692992, 0.3864523, 0.413464, 0.3642905,
  0.2202491, 0.149751, 0.1243173, 0.2228902, 0.2688572, 0.2502086, 0.2382512, 
    0.2205184, 0.2174278, 0.1203141, 0.1270684, 0.05047294, 0.01949758, 
    0.1322657, 0.2124812, 0.1731798, 0.1445387, 0.1429324, 0.1545159, 
    0.1132387, 0.1045771, 0.1146341, 0.1277723, 0.3526389, 0.02831369, 
    0.1002883, 0.187959, 0.1958174, 0.2538636,
  0.1337495, 0.0838071, 0.008823113, 0.106153, 0.1198273, 0.1654768, 
    0.09317039, 0.1015211, 0.1104996, 0.02795513, 0.01224175, 0.0003311452, 
    0.03091315, 0.09200995, 0.1317015, 0.1195699, 0.1128861, 0.1418768, 
    0.1299703, 0.1306577, 0.1051182, 0.0972458, 0.1699836, 0.00874659, 
    0.04653554, 0.1671828, 0.1446519, 0.135013, 0.100414,
  0.3386116, -0.0003604239, 0.006063188, 0.07609227, 0.005148379, 0.02199621, 
    0.03488808, 0.03952342, 0.09009855, 0.0004176478, 1.398264e-08, 
    -1.040574e-06, 0.03457148, 0.1220702, 0.1401996, 0.1019003, 0.06374205, 
    0.07722598, 0.02472005, 0.02148052, 0.04972458, 0.09695457, 0.2448013, 
    0.009787343, 0.003673953, 0.02710491, 0.03446441, 0.05384465, 0.1789524,
  0.634236, 0.1257122, -2.967688e-06, 0.02610999, 0.02637232, 0.02628165, 
    0.04907491, 0.04308196, 0.01632309, 0.02688178, 0.02703515, 0.02026346, 
    0.1390282, 0.0735643, 0.03120134, 0.01546087, 0.01463317, 0.008102444, 
    0.008009435, 0.004998842, 0.04002155, 0.2576224, 0.3201898, 0.003803473, 
    0.0006901201, 1.439043e-07, 0.02879066, 0.06979722, 0.3314675,
  0.1747132, 0.1208207, 0.01774453, 0.05403296, 0.07804032, 0.04269854, 
    0.03892268, 0.04402574, 0.04496701, 0.1142129, 0.07238338, 0.06588567, 
    0.02569572, 0.01555572, 0.01116929, 0.013101, 0.0261375, 0.02052912, 
    0.03149598, 0.04403574, 0.1545624, 0.2724883, 0.05656823, 0.00644567, 
    0.001022336, 0.04279033, 0.02970411, 0.08758648, 0.3069291,
  0.01231938, 0.02250182, 0.004320612, 0.03643258, -8.108808e-05, 0.02483127, 
    0.06167163, 0.02282635, 0.006973164, 0.0261936, 0.006168792, 0.09036021, 
    0.02927469, 0.03902717, 0.04826434, 0.05740826, 0.06899393, 0.1190257, 
    0.1318006, 0.1538486, 0.08958225, 0.1111949, 0.154514, 0.02651874, 
    0.01681513, 0.04683174, 0.06860991, 0.1324271, 0.03143943,
  3.416097e-08, 8.62734e-08, -1.231951e-06, 0.0003815558, -4.086008e-08, 
    0.09705719, 0.01548649, 0.04267349, 0.1136176, 0.07085202, 0.09665762, 
    0.03547765, 0.01666636, 0.02027817, 0.01580072, 0.01451179, 0.01575975, 
    0.06199588, 0.2095201, 0.2537523, 0.0901657, 0.1782611, 0.01188082, 
    0.004389918, 0.04288698, 0.08247896, 0.2153084, 0.1082468, 3.440666e-06,
  4.688338e-07, 0.002787599, 0.0004559392, -6.964432e-09, 1.352226e-07, 
    5.167663e-09, -0.0001110913, 0.2114022, 0.3942137, 0.1414627, 0.1202742, 
    0.07655258, 0.104154, 0.08492453, 0.1176166, 0.07406255, 0.06489697, 
    0.09016801, 0.2334026, 0.05357355, 0.01661368, 0.03514583, 0.04093098, 
    0.06714411, 0.0478643, 0.0440364, 0.09051215, 0.1262583, 0.006175794,
  0.005893644, 0.007731486, 0.0006184092, 0.1512624, 0.0002206587, 
    -1.246941e-05, 0.0526196, -1.825955e-05, -3.647307e-05, 0.02715823, 
    0.0918588, 0.1052473, 0.2009922, 0.2807402, 0.2926633, 0.2922831, 
    0.2259659, 0.3177362, 0.3127607, 0.0002204052, 0.0003051626, 0.01931216, 
    0.1035049, 0.09905062, 0.1097039, 0.1089371, 0.1407943, 0.1068604, 
    0.07920726,
  0.0927614, 0.2418229, 0.166885, 0.1962443, 0.03186165, 0.01937624, 
    0.04194052, 0.198809, 0.09629081, 0.1195177, 0.09920168, 0.1636844, 
    0.3333993, 0.3500822, 0.2554213, 0.3119635, 0.3455126, 0.292461, 
    0.2397914, 0.1119095, 0.06980333, 0.02660705, 0.1315241, 0.2994614, 
    0.2039659, 0.3270988, 0.3371266, 0.2746337, 0.1856934,
  0.2154544, 0.2427255, 0.169727, 0.1792382, 0.2149942, 0.1577508, 0.1277343, 
    0.1309904, 0.2054285, 0.2317924, 0.2295047, 0.3593999, 0.2998248, 
    0.290415, 0.3216661, 0.3165444, 0.3826392, 0.4196082, 0.3095686, 
    0.1325765, 0.1317041, 0.2663589, 0.420001, 0.4567596, 0.3664483, 
    0.212263, 0.3360831, 0.227228, 0.2258841,
  0.5049893, 0.309576, 0.3859973, 0.3614475, 0.3943682, 0.3529729, 0.3630015, 
    0.3554841, 0.2850235, 0.2295271, 0.4488031, 0.3588002, 0.3948055, 
    0.3889221, 0.4267176, 0.4684021, 0.4722255, 0.3446546, 0.3344565, 
    0.3496285, 0.4165515, 0.4779038, 0.4416514, 0.4580062, 0.3643933, 
    0.3482598, 0.2161186, 0.1547261, 0.4609103,
  0.5429076, 0.4807582, 0.4952365, 0.5325277, 0.6590031, 0.5635175, 
    0.5278287, 0.5261879, 0.4579364, 0.4530974, 0.4360262, 0.3913153, 
    0.3860343, 0.3786293, 0.4050117, 0.4752868, 0.5332646, 0.6312798, 
    0.6092086, 0.5734485, 0.4962335, 0.3448243, 0.3362615, 0.4491107, 
    0.3003839, 0.3264813, 0.2216529, 0.2465069, 0.4003975,
  0.1701497, 0.1656838, 0.1612179, 0.156752, 0.1522861, 0.1478202, 0.1433543, 
    0.125723, 0.1337861, 0.1418493, 0.1499125, 0.1579756, 0.1660388, 
    0.174102, 0.2031372, 0.2062439, 0.2093506, 0.2124573, 0.215564, 
    0.2186707, 0.2217773, 0.2381786, 0.2314746, 0.2247707, 0.2180667, 
    0.2113628, 0.2046588, 0.1979549, 0.1737224,
  0.2971594, 0.1920792, 0.114117, 0.0655183, 0.01744704, -0.001074829, 
    -0.0004721635, 0.003386967, 0.0008388155, 0.003160056, 0.02049858, 
    0.1318347, 0.2558601, 0.04577217, 0.1376514, 0.2056413, 0.2900065, 
    0.3004135, 0.221242, 0.2255727, 0.3713909, 0.3515099, 0.2407506, 
    0.2336111, 0.214007, 0.2149927, 0.1578802, 0.1690565, 0.2977414,
  0.2065277, 0.1432674, 0.2010062, 0.06004888, 0.1157907, 0.04575486, 
    0.04006269, 0.2974037, 0.2707042, 0.2979814, 0.2710364, 0.1631531, 
    0.1674786, 0.1860923, 0.3523506, 0.4241579, 0.3869197, 0.4065892, 
    0.4202935, 0.4515051, 0.3649368, 0.4021229, 0.4023888, 0.5620699, 
    0.2718676, 0.3867953, 0.4344539, 0.4037154, 0.309435,
  0.4575455, 0.416659, 0.4105227, 0.2267853, 0.2586693, 0.3347939, 0.3379273, 
    0.4011508, 0.3223519, 0.1490808, 0.1512045, 0.250698, 0.2804205, 
    0.3181038, 0.277027, 0.3421996, 0.3619058, 0.3728538, 0.3060391, 
    0.2229259, 0.2352293, 0.219777, 0.3299696, 0.2213399, 0.3227853, 
    0.4186658, 0.4272016, 0.4575431, 0.4161536,
  0.2912691, 0.2946765, 0.2788876, 0.273205, 0.3051, 0.3052609, 0.3058538, 
    0.2056947, 0.2089285, 0.2289646, 0.2066711, 0.2294817, 0.1559368, 
    0.1828511, 0.1326199, 0.1999518, 0.2024267, 0.2611506, 0.2650392, 
    0.2767669, 0.2302153, 0.2766242, 0.2428806, 0.1920506, 0.1002567, 
    0.2638951, 0.3771704, 0.3863732, 0.3383392,
  0.1596072, 0.08978999, 0.1042289, 0.2035531, 0.2834147, 0.2207262, 
    0.1906027, 0.1696355, 0.1554635, 0.07184045, 0.06896085, 0.02908527, 
    0.008603917, 0.117494, 0.1924333, 0.128885, 0.1048442, 0.09868847, 
    0.1352741, 0.09865619, 0.09258548, 0.1034869, 0.1049179, 0.3531644, 
    0.02166347, 0.09209459, 0.1447302, 0.1708073, 0.2074865,
  0.04676183, 0.05025037, 0.009568989, 0.07563698, 0.06623099, 0.055586, 
    0.03273454, 0.03926232, 0.04195385, 0.01140639, 0.01009192, 0.0003394008, 
    0.02588105, 0.06258054, 0.1002448, 0.1066576, 0.1204315, 0.1041889, 
    0.11766, 0.1060188, 0.07002987, 0.05472261, 0.06512438, 0.006037064, 
    0.03384756, 0.1541815, 0.1028282, 0.07500012, 0.04793116,
  0.1459396, 0.000732156, 0.00606467, 0.02570526, -0.00312283, 0.01464429, 
    0.01714284, 0.008155859, 0.02748096, 0.01930949, 9.703624e-09, 
    -3.738028e-07, 0.009773189, 0.08927515, 0.1067258, 0.04774154, 
    0.02117254, 0.033167, 0.01094701, 0.004529264, 0.01392686, 0.03029906, 
    0.09386291, 0.02220114, 0.001050409, 0.03572024, 0.01110525, 0.01537191, 
    0.06304972,
  0.3632317, 0.2631751, -1.147735e-05, 0.05101311, 0.01000638, 0.007816956, 
    0.02341985, 0.02321405, 0.002002235, 0.003862225, 0.02171494, 
    0.007911863, 0.111861, 0.03818862, 0.009473201, 0.003152907, 0.001743137, 
    0.0003734692, 0.0002313938, 0.0003197358, 0.01059021, 0.08815686, 
    0.3038557, 0.001120337, 0.0002681695, 1.629925e-07, 0.001853543, 
    0.01833657, 0.1264694,
  0.1169108, 0.1028886, 0.01310337, 0.04392088, 0.02712252, 0.009380437, 
    0.01237597, 0.02492212, 0.04284766, 0.0775425, 0.02853279, 0.01311976, 
    0.004440646, 0.003422957, 0.002031166, 0.001689633, 0.006343174, 
    0.005724269, 0.01466731, 0.01878385, 0.06591097, 0.4405597, 0.2951544, 
    0.00421428, 0.000401938, 0.008544302, 0.005562871, 0.01543092, 0.1921003,
  0.006165201, 0.02031611, 0.004946264, 0.0345208, -1.759281e-05, 
    0.006055089, 0.07346046, 0.003141764, 0.0006790479, 0.01328407, 
    0.002314238, 0.02085974, 0.008223576, 0.01367006, 0.01398933, 0.03091761, 
    0.0324451, 0.0511102, 0.07071908, 0.1192818, 0.04538772, 0.05956919, 
    0.1744168, 0.01741166, 0.003747495, 0.009121815, 0.01977289, 0.08402843, 
    0.02347559,
  4.351245e-08, 7.387884e-08, -4.455799e-07, -9.490113e-06, -1.450657e-08, 
    0.2006969, 0.02024966, 0.02674928, 0.08093502, 0.04033971, 0.03404699, 
    0.01188409, 0.00439179, 0.005386471, 0.003769812, 0.001923746, 
    0.002417478, 0.01847689, 0.09788069, 0.2001319, 0.09828949, 0.1492973, 
    0.001772764, -0.001036968, 0.008292914, 0.02315784, 0.1010811, 0.1033071, 
    1.773543e-06,
  4.18409e-07, 0.005184643, 0.0005533636, -7.690873e-08, 1.201686e-07, 
    4.865122e-09, -7.780117e-05, 0.2281697, 0.3603827, 0.1214325, 0.106406, 
    0.04449507, 0.04526564, 0.03582254, 0.05942903, 0.02507439, 0.03082155, 
    0.04765284, 0.1528675, 0.1475054, 0.01765074, 0.02488909, 0.024892, 
    0.01528531, 0.01298569, 0.007418736, 0.02314811, 0.04352634, 0.009013576,
  0.004793922, 0.01410196, 0.0004909478, 0.1672707, -0.0003408044, 
    -1.516808e-05, 0.04697334, -8.451265e-06, -5.021751e-05, 0.02808786, 
    0.0991226, 0.08450697, 0.2066752, 0.2359341, 0.2930702, 0.2672647, 
    0.2743596, 0.2563041, 0.2523539, 0.0002084674, 5.70595e-05, 0.02855684, 
    0.08690129, 0.1394013, 0.09001304, 0.08200229, 0.09338513, 0.06008351, 
    0.09748691,
  0.06870224, 0.2284279, 0.162112, 0.1767766, 0.0261756, 0.02150546, 
    0.03758973, 0.1928097, 0.08082254, 0.1155119, 0.08647253, 0.1593271, 
    0.3380235, 0.3205759, 0.2251909, 0.2978879, 0.2979674, 0.2601981, 
    0.2178085, 0.1096579, 0.06474593, 0.02078475, 0.1144775, 0.2901702, 
    0.1994763, 0.2959841, 0.2714354, 0.2522196, 0.1887978,
  0.1848283, 0.2402498, 0.1387195, 0.1694304, 0.2145857, 0.1480408, 
    0.1115127, 0.123016, 0.2001756, 0.2223856, 0.2234216, 0.3925237, 
    0.3168225, 0.2568498, 0.2570699, 0.2665805, 0.3900846, 0.3903675, 
    0.3199793, 0.1194797, 0.09971906, 0.2273365, 0.3237233, 0.4219509, 
    0.3738253, 0.1778103, 0.3115392, 0.2236429, 0.1901411,
  0.414206, 0.2278935, 0.4006046, 0.3073168, 0.3898213, 0.3372683, 0.3594623, 
    0.3218771, 0.26055, 0.2193554, 0.4572676, 0.3264952, 0.3254877, 
    0.3497207, 0.3894425, 0.3867567, 0.4150034, 0.2705697, 0.2496531, 
    0.2842372, 0.3913799, 0.4602062, 0.4669501, 0.5122231, 0.3273657, 
    0.3347009, 0.2123106, 0.1141961, 0.4075949,
  0.5069418, 0.3886043, 0.4337086, 0.5345371, 0.5981673, 0.5361886, 
    0.4962772, 0.5140857, 0.4606839, 0.4547338, 0.4822758, 0.4162745, 
    0.3733894, 0.3719513, 0.3695988, 0.480632, 0.5765515, 0.6180604, 
    0.6154264, 0.5559211, 0.4475475, 0.2885213, 0.3655686, 0.5197038, 
    0.3051027, 0.3023787, 0.2138086, 0.280832, 0.3646699,
  0.07365185, 0.07002918, 0.0664065, 0.06278384, 0.05916116, 0.05553849, 
    0.05191582, 0.03673611, 0.04481424, 0.05289238, 0.06097051, 0.06904864, 
    0.07712676, 0.0852049, 0.0982684, 0.1002923, 0.1023163, 0.1043403, 
    0.1063642, 0.1083882, 0.1104121, 0.129479, 0.1229996, 0.1165202, 
    0.1100408, 0.1035614, 0.09708195, 0.09060254, 0.07654998,
  0.2948656, 0.1838551, 0.08708198, 0.06065741, 0.02055692, -0.0008092605, 
    -0.0002014484, 0.001387496, 0, 2.161349e-08, 0.009298888, 0.06692966, 
    0.2376788, 0.0268416, 0.1548609, 0.2271246, 0.3097567, 0.2717972, 
    0.1955988, 0.2267171, 0.3748837, 0.35313, 0.2085514, 0.2081199, 
    0.1901496, 0.2338191, 0.1502164, 0.1463305, 0.3064364,
  0.197607, 0.1092328, 0.1845827, 0.03780575, 0.07902084, 0.03860783, 
    0.02516349, 0.2781068, 0.2367606, 0.2722762, 0.2611706, 0.1638136, 
    0.1479933, 0.1605164, 0.3547617, 0.4207038, 0.4030818, 0.4283158, 
    0.4259156, 0.4620897, 0.3707197, 0.3897406, 0.4054064, 0.5650203, 
    0.2391495, 0.4526308, 0.4766018, 0.4266214, 0.304406,
  0.4596169, 0.4221462, 0.3360587, 0.166464, 0.2052333, 0.2739741, 0.3235108, 
    0.3442317, 0.2868958, 0.1138737, 0.1199357, 0.1989004, 0.2547718, 
    0.2812774, 0.2432258, 0.3080369, 0.3257743, 0.3430952, 0.250658, 
    0.1870573, 0.1935645, 0.1810592, 0.2815212, 0.1921967, 0.2965046, 
    0.401283, 0.4040264, 0.45367, 0.4210372,
  0.2545547, 0.2739779, 0.2439707, 0.2324411, 0.2894306, 0.276798, 0.2658766, 
    0.171822, 0.1751475, 0.1866858, 0.1496548, 0.1698814, 0.1047254, 
    0.1484185, 0.09710826, 0.15376, 0.1528496, 0.2135234, 0.2181728, 
    0.223564, 0.1786517, 0.216723, 0.182448, 0.1566363, 0.07503069, 
    0.2377559, 0.3284967, 0.3641624, 0.296436,
  0.1160145, 0.0529923, 0.07540019, 0.1733544, 0.2590671, 0.1803193, 
    0.1334553, 0.1183107, 0.09747462, 0.04304454, 0.04749676, 0.01424618, 
    0.004838378, 0.1035649, 0.1555748, 0.09295428, 0.07446324, 0.07352551, 
    0.1129397, 0.08633627, 0.08295934, 0.08308873, 0.08283633, 0.3301689, 
    0.01809554, 0.08179104, 0.1084654, 0.139781, 0.1797387,
  0.02004582, 0.02350111, 0.008444505, 0.0401656, 0.03754363, 0.02377901, 
    0.01360238, 0.01622812, 0.01961978, 0.006101665, 0.006387373, 
    0.0001781972, 0.01981403, 0.04262714, 0.07871635, 0.08279733, 0.09173286, 
    0.07592408, 0.09934294, 0.07828856, 0.03668838, 0.03495076, 0.02747853, 
    0.003530668, 0.02243681, 0.1299721, 0.06007284, 0.04538802, 0.02463593,
  0.0683159, 0.004531578, 0.003624054, 0.006960474, -0.003403286, 
    0.008456178, 0.00725337, 0.002693314, 0.01168469, 0.01685091, 
    7.364769e-09, 5.066829e-08, 0.003146651, 0.04947303, 0.06801908, 
    0.01627755, 0.005466027, 0.01027257, 0.003471137, 0.001387696, 
    0.00558744, 0.01236225, 0.04205802, 0.01862244, 0.0004493681, 0.04355686, 
    0.001745575, 0.004399906, 0.02430713,
  0.1621465, 0.1773962, -4.856804e-06, 0.08092777, 0.00281264, 0.001281876, 
    0.006409046, 0.008569619, 0.0007346662, -0.001171673, 0.01418689, 
    0.002852591, 0.06799442, 0.007415767, 0.001034274, 0.0007127048, 
    0.0003751034, 6.110925e-05, 6.503306e-05, 0.0001325437, 0.003946496, 
    0.03456335, 0.1400613, 0.0004084492, 0.0002043158, 8.811676e-08, 
    0.0004725137, 0.007483009, 0.04912522,
  0.02503854, 0.1026144, 0.01061788, 0.03052501, 0.005889304, 0.002642527, 
    0.004778859, 0.01089738, 0.0471979, 0.0630746, 0.004969304, 0.002353994, 
    0.0003538904, 0.0006972899, 0.0007726195, 0.0005471141, 0.000626238, 
    0.0006225383, 0.001540736, 0.002266562, 0.01416039, 0.1943876, 0.1476553, 
    0.002797041, 0.000190131, 0.003058954, 0.001355349, 0.003888984, 
    0.05880943,
  0.00501445, 0.01868585, 0.002647264, 0.03641082, 5.441926e-05, 
    0.0009160301, 0.07351863, 0.0002060693, -0.0008788376, 0.003453422, 
    0.0002962815, 0.008025607, 0.003164258, 0.00387424, 0.005546118, 
    0.01263269, 0.01107966, 0.03046092, 0.04323058, 0.06527974, 0.01825744, 
    0.02619887, 0.1785285, 0.0158567, 0.001149328, 0.002925338, 0.004769133, 
    0.02233571, 0.02254891,
  4.747962e-08, 6.453077e-08, -1.359109e-07, -1.622418e-05, -6.963068e-10, 
    0.1596394, 0.017457, 0.009401361, 0.0647405, 0.01431113, 0.01711102, 
    0.002750882, 0.0006044729, 0.002099704, 0.0007847436, 0.0003675467, 
    0.0009196657, 0.006643929, 0.04147745, 0.1337554, 0.0205247, 0.1115672, 
    0.0005470818, -0.001324981, 0.002265009, 0.007958075, 0.03680041, 
    0.03630281, 6.784326e-07,
  3.850029e-07, 0.004310717, 0.0004109627, 2.594481e-06, 1.099642e-07, 
    4.79778e-09, -4.096074e-05, 0.2306634, 0.3286141, 0.09570121, 0.06513146, 
    0.01278946, 0.01273081, 0.01234409, 0.01682383, 0.006934867, 0.006857442, 
    0.02720346, 0.05843538, 0.2981738, 0.01562279, 0.02002831, 0.01737746, 
    0.005807113, 0.002657394, 0.001927869, 0.007333633, 0.02044796, 0.0144135,
  0.00483295, 0.005149534, 0.00157136, 0.1784635, -0.0004862183, 
    -1.198506e-05, 0.04454616, -4.315908e-06, -0.000108778, 0.02591855, 
    0.09900783, 0.06646955, 0.1764181, 0.1852826, 0.2514716, 0.2260052, 
    0.2287678, 0.154288, 0.1792406, 0.0001937509, -0.0001337237, 0.03474851, 
    0.069093, 0.1419531, 0.06155197, 0.07720549, 0.05904529, 0.03448045, 
    0.07173759,
  0.06018337, 0.2124285, 0.1531486, 0.1565722, 0.02001759, 0.01640979, 
    0.02741722, 0.1811334, 0.07206379, 0.1092164, 0.07726332, 0.1533309, 
    0.3356216, 0.292501, 0.1954461, 0.2658952, 0.2191435, 0.2077955, 
    0.1993596, 0.1036631, 0.05359168, 0.01573022, 0.09978552, 0.2741869, 
    0.1864561, 0.263094, 0.2357052, 0.1973634, 0.1391318,
  0.1408251, 0.2233958, 0.1220047, 0.1538037, 0.2175043, 0.1285937, 
    0.09349705, 0.1099202, 0.1951757, 0.2154371, 0.1974933, 0.4252678, 
    0.3179562, 0.2246034, 0.1952511, 0.2385598, 0.379404, 0.3591202, 
    0.3043355, 0.1136521, 0.08207648, 0.213768, 0.2744896, 0.4059684, 
    0.3460527, 0.1636708, 0.2791256, 0.1798764, 0.1668085,
  0.3496708, 0.1592428, 0.3743796, 0.2703945, 0.3645288, 0.2981898, 
    0.3358246, 0.2947485, 0.2365661, 0.2273042, 0.454425, 0.3199482, 
    0.2782314, 0.2954502, 0.3354656, 0.3242244, 0.3581926, 0.2140784, 
    0.2043543, 0.228445, 0.3903778, 0.411029, 0.4273463, 0.5397006, 
    0.2755679, 0.2946779, 0.2048155, 0.09727945, 0.3552438,
  0.4330071, 0.2906175, 0.3664359, 0.4912907, 0.5007913, 0.4663919, 
    0.4635757, 0.4861827, 0.4687148, 0.4755304, 0.4428943, 0.3732213, 
    0.3639584, 0.3888425, 0.3657696, 0.4531916, 0.5555384, 0.5507431, 
    0.5803194, 0.4962723, 0.378009, 0.2502054, 0.3469117, 0.5336725, 
    0.2805723, 0.2673048, 0.1954232, 0.2771929, 0.3149886,
  0.00980832, 0.008894199, 0.007980078, 0.007065956, 0.006151835, 
    0.005237714, 0.004323594, -0.006020077, -0.002871081, 0.0002779146, 
    0.00342691, 0.006575905, 0.009724901, 0.0128739, 0.01094162, 0.01140001, 
    0.0118584, 0.01231678, 0.01277517, 0.01323356, 0.01369195, 0.02410211, 
    0.02140884, 0.01871558, 0.01602232, 0.01332906, 0.0106358, 0.007942535, 
    0.01053962,
  0.2988582, 0.1383386, 0.06833239, 0.045164, 0.01356459, -0.0003234005, 
    0.0001872448, -5.916665e-06, 0, 0, -0.0002183428, 0.03156929, 0.1676084, 
    0.01785026, 0.1891961, 0.2867711, 0.3829582, 0.2570856, 0.1582277, 
    0.2664829, 0.3951151, 0.3449228, 0.1625803, 0.1497994, 0.1926753, 
    0.2895325, 0.1915673, 0.1184471, 0.2924014,
  0.2107595, 0.09483878, 0.1629201, 0.02265855, 0.05012039, 0.02666391, 
    0.01696078, 0.2266569, 0.1836768, 0.2029155, 0.2325689, 0.143315, 
    0.1325624, 0.1355549, 0.3639204, 0.4148858, 0.3713494, 0.3842729, 
    0.3881734, 0.4226032, 0.3644035, 0.3523638, 0.3757908, 0.5318422, 
    0.2349081, 0.4917661, 0.4788727, 0.4323131, 0.3103553,
  0.4049028, 0.3880407, 0.2701667, 0.1212298, 0.1498997, 0.2098338, 
    0.2827878, 0.2744154, 0.2218079, 0.08247627, 0.08814852, 0.1511238, 
    0.207136, 0.2303482, 0.1921851, 0.2603508, 0.2791956, 0.2867603, 
    0.1920067, 0.148129, 0.1547599, 0.1398696, 0.2124682, 0.1519147, 
    0.2510371, 0.3445125, 0.3717562, 0.4125816, 0.3899398,
  0.211639, 0.2259119, 0.1968516, 0.1878996, 0.2443772, 0.2270321, 0.219529, 
    0.131752, 0.1358203, 0.1400342, 0.1013798, 0.1167191, 0.06646208, 
    0.1047231, 0.07353311, 0.1035082, 0.09904689, 0.1643804, 0.1483139, 
    0.1532151, 0.1343407, 0.1477058, 0.1243779, 0.122734, 0.05945228, 
    0.1866212, 0.2439933, 0.3076053, 0.2407297,
  0.08916818, 0.02976594, 0.04844699, 0.1345486, 0.1956919, 0.123906, 
    0.08806528, 0.07096268, 0.05333433, 0.02681387, 0.02468111, 0.007332355, 
    0.002343411, 0.07625741, 0.1233207, 0.06457753, 0.04457375, 0.05342049, 
    0.08390453, 0.06395413, 0.06617048, 0.06090314, 0.05719781, 0.2958562, 
    0.01533847, 0.07265694, 0.08268933, 0.1021373, 0.1445929,
  0.01087351, 0.01377521, 0.007093037, 0.01807355, 0.01973979, 0.01616811, 
    0.007779481, 0.009644603, 0.01166646, 0.003717542, 0.003959297, 
    7.275233e-05, 0.01379528, 0.03320935, 0.05560397, 0.06110533, 0.04805475, 
    0.05763367, 0.06854942, 0.04575306, 0.01970838, 0.02094196, 0.01600819, 
    0.002527389, 0.02025527, 0.08713864, 0.0376176, 0.02533554, 0.01397005,
  0.03927196, 0.007663419, 0.001343252, 0.003142182, -0.003008681, 
    0.003993605, 0.003004797, 0.001450236, 0.00647985, 0.007327797, 
    6.076137e-09, 6.641289e-08, 0.001670281, 0.02573149, 0.04032007, 
    0.005150573, 0.001751017, 0.002725295, 0.0009715504, 0.0006086613, 
    0.002978395, 0.006722358, 0.02351175, 0.01650787, 0.0002009739, 
    0.0486404, 0.0007921893, 0.002176784, 0.01237329,
  0.08255801, 0.08143108, -1.298408e-06, 0.07616416, 0.0007374111, 
    0.0002574647, 0.0016139, 0.002571041, 0.0004013671, -0.001910791, 
    0.008777949, 0.001036062, 0.03415002, 0.00149278, 0.0001333226, 
    0.0002368634, 0.0001376996, 3.067985e-05, 2.896959e-05, 7.281723e-05, 
    0.002030691, 0.0179569, 0.07629935, 0.0002758979, 0.0001485195, 
    8.17647e-08, 0.0004588525, 0.004114958, 0.02487987,
  0.0106013, 0.1081898, 0.008370994, 0.01970175, 0.001224239, 0.0008889914, 
    0.002030728, 0.005141631, 0.04076486, 0.06389458, 0.001267092, 
    0.0008029847, 6.172612e-05, 0.0002942846, 0.0004263937, 0.0002761889, 
    0.0002731222, 0.0002736165, 0.0004702825, 0.000739112, 0.005372317, 
    0.08175952, 0.07988334, 0.001576184, 8.065946e-05, 0.001624012, 
    0.0007060264, 0.001869895, 0.0256004,
  0.005340301, 0.01466143, 0.001678268, 0.03515205, 2.56754e-05, 0.000363179, 
    0.04691941, 5.628737e-05, -0.0009567988, 0.001064813, 5.20323e-05, 
    0.004723202, 0.001031666, 0.001273855, 0.003217089, 0.005920738, 
    0.006021374, 0.0205157, 0.02754956, 0.03075096, 0.006941699, 0.01122693, 
    0.1572069, 0.01619865, 0.000486567, 0.00139493, 0.002066971, 0.007293589, 
    0.02225436,
  4.47212e-08, 5.880788e-08, 7.02689e-09, -1.087264e-05, 2.814975e-09, 
    0.08949606, 0.01146299, 0.002734977, 0.05610227, 0.005540949, 
    0.008416375, 0.0008845042, 9.78818e-05, 0.0006564855, 0.0003069693, 
    9.010825e-05, 0.0005085961, 0.0033157, 0.01731199, 0.09064846, 
    0.006409692, 0.0889293, 0.0002965639, -0.001197428, 0.0008935879, 
    0.003447458, 0.01699683, 0.01479561, 3.35846e-07,
  3.622228e-07, 0.00395327, 0.001195503, 1.766187e-06, 1.026348e-07, 
    4.793947e-09, -2.925057e-05, 0.2174227, 0.2959171, 0.06241737, 
    0.02591436, 0.004437874, 0.004715761, 0.00488247, 0.007466945, 
    0.003048881, 0.002632914, 0.007621925, 0.02985042, 0.2726017, 0.01225971, 
    0.01322848, 0.01104557, 0.003045885, 0.001229372, 0.0009915468, 
    0.003424039, 0.01241252, 0.01382636,
  0.004499676, 0.001906416, 0.002082808, 0.1773043, -0.0004639578, 
    -3.475914e-06, 0.04174653, -3.148831e-06, -0.0001669863, 0.0193347, 
    0.09462553, 0.0586887, 0.1434614, 0.1372169, 0.20514, 0.19846, 0.148769, 
    0.09000632, 0.133585, 1.189639e-05, 0.000383727, 0.03849517, 0.05027332, 
    0.1072235, 0.03709617, 0.04972217, 0.03829128, 0.0195935, 0.05458511,
  0.04354844, 0.1938827, 0.1364602, 0.1233552, 0.01273227, 0.009888474, 
    0.01918878, 0.1604373, 0.06343532, 0.0978348, 0.07023077, 0.1468971, 
    0.3151495, 0.2572003, 0.1637994, 0.2126002, 0.1787405, 0.1646708, 
    0.1835018, 0.09557273, 0.04219434, 0.01199893, 0.07856034, 0.244334, 
    0.1648587, 0.2426083, 0.1960675, 0.1573988, 0.07915291,
  0.09279644, 0.1997663, 0.1016306, 0.130065, 0.1975663, 0.1132643, 
    0.07725541, 0.09661338, 0.1778082, 0.1910006, 0.1706778, 0.3951636, 
    0.3005376, 0.181802, 0.1477591, 0.1967494, 0.3575015, 0.3213106, 
    0.2631091, 0.1074979, 0.06877691, 0.193732, 0.2089593, 0.3744649, 
    0.2962903, 0.1381109, 0.2486798, 0.1426515, 0.1423475,
  0.2850103, 0.113011, 0.3318022, 0.2247386, 0.3085566, 0.2805671, 0.3033749, 
    0.2675427, 0.2010412, 0.2102105, 0.4262122, 0.2953333, 0.2528228, 
    0.2338988, 0.294112, 0.279677, 0.3058926, 0.1675165, 0.1733267, 
    0.1816697, 0.3492021, 0.364044, 0.3721021, 0.5517449, 0.2277931, 
    0.2531992, 0.2076295, 0.08167446, 0.2931336,
  0.3906845, 0.2275443, 0.3185859, 0.4299718, 0.4241523, 0.41494, 0.43317, 
    0.439761, 0.3928406, 0.4517646, 0.3956183, 0.3171236, 0.344022, 
    0.3767863, 0.3338538, 0.4047678, 0.4748385, 0.4683235, 0.4764604, 
    0.4393076, 0.3308302, 0.224325, 0.3257116, 0.5160327, 0.2547778, 
    0.2473545, 0.1654406, 0.2606813, 0.2875293,
  0.003417513, 0.003094498, 0.002771482, 0.002448467, 0.002125452, 
    0.001802436, 0.001479421, 0.003928916, 0.005239491, 0.006550066, 
    0.00786064, 0.009171216, 0.01048179, 0.01179237, 0.009125848, 
    0.008355989, 0.00758613, 0.006816271, 0.006046412, 0.005276552, 
    0.004506694, 0.004603487, 0.004385787, 0.004168087, 0.003950386, 
    0.003732685, 0.003514985, 0.003297285, 0.003675925,
  0.2740516, 0.09424415, 0.05737121, 0.0206297, -0.001198352, -6.544229e-05, 
    -4.574569e-05, -2.599942e-06, 0, 0, 0.000299844, 0.008123701, 0.09197147, 
    0.009642414, 0.2249262, 0.338808, 0.3770384, 0.2261725, 0.1340213, 
    0.2800514, 0.4186938, 0.3759786, 0.1207509, 0.1030278, 0.1918025, 
    0.3644189, 0.1840231, 0.1031269, 0.3030601,
  0.1963727, 0.07799517, 0.1434179, 0.01476667, 0.03893095, 0.01593057, 
    0.01017745, 0.1168132, 0.08699615, 0.1409165, 0.1867821, 0.1067282, 
    0.1189409, 0.1099619, 0.346481, 0.3752227, 0.3270426, 0.3017992, 
    0.3305807, 0.3581219, 0.3162827, 0.3118177, 0.3292125, 0.4773097, 
    0.2214907, 0.4561383, 0.4396273, 0.3937865, 0.2794225,
  0.3392662, 0.313752, 0.2215842, 0.09497114, 0.1156845, 0.1639057, 0.23975, 
    0.2243594, 0.1780007, 0.05874592, 0.06674244, 0.1166708, 0.1597517, 
    0.1818719, 0.1418985, 0.1999583, 0.2187211, 0.2275286, 0.147633, 
    0.1134328, 0.1190504, 0.09998385, 0.1576319, 0.1071922, 0.1974714, 
    0.2846303, 0.3303897, 0.3472645, 0.3279799,
  0.1675631, 0.1811796, 0.1549392, 0.1499802, 0.2081136, 0.1864132, 
    0.1761801, 0.09995186, 0.104845, 0.09845741, 0.06630497, 0.07069745, 
    0.03902531, 0.06701784, 0.04982632, 0.06688043, 0.06253006, 0.1120005, 
    0.09683405, 0.1016477, 0.09038793, 0.09678476, 0.07729658, 0.09694201, 
    0.04660776, 0.1347563, 0.1762281, 0.236631, 0.1900813,
  0.05819861, 0.01651817, 0.03304226, 0.0926976, 0.1303476, 0.07580318, 
    0.05341195, 0.0405634, 0.02805919, 0.01305626, 0.01362064, 0.00400861, 
    0.001269856, 0.04799145, 0.09481905, 0.04271912, 0.02474873, 0.03435077, 
    0.05796303, 0.03821838, 0.04113419, 0.03700672, 0.03305742, 0.2632295, 
    0.01265874, 0.0578973, 0.05675809, 0.06666837, 0.09567813,
  0.007209056, 0.00841438, 0.005397661, 0.00861102, 0.01078025, 0.01048883, 
    0.005539527, 0.006906436, 0.008196888, 0.00252517, 0.002340765, 
    4.442206e-05, 0.009011059, 0.02217181, 0.03538015, 0.04325113, 
    0.02108063, 0.03978266, 0.03815601, 0.02508349, 0.01030182, 0.01221506, 
    0.01128059, 0.001698488, 0.01936926, 0.05113565, 0.0209389, 0.01212031, 
    0.008144506,
  0.02653511, 0.009644415, 0.0005979617, 0.002002733, -0.002305503, 
    0.001801896, 0.001428488, 0.00094783, 0.004268437, 0.003764907, 
    5.334589e-09, 5.431397e-08, 0.001103784, 0.01377872, 0.01664891, 
    0.002375765, 0.0009897941, 0.0009258842, 0.0004050999, 0.0003381039, 
    0.001893671, 0.004316805, 0.01559454, 0.01321043, 0.0001001641, 
    0.04565823, 0.0006634677, 0.001362848, 0.007795132,
  0.05133304, 0.0389597, -1.158779e-08, 0.05393265, 0.0002682749, 
    0.0001232901, 0.0006697869, 0.0007835904, 0.0002635988, -0.001191105, 
    0.006026003, 0.0004557848, 0.0154206, 0.0004993783, 6.428788e-05, 
    9.360925e-05, 7.19132e-05, 2.031836e-05, 1.662657e-05, 4.815626e-05, 
    0.001277589, 0.01141146, 0.04890135, 0.0001952712, 0.0001083695, 
    5.719564e-08, 0.0005045137, 0.00269384, 0.01564692,
  0.006190693, 0.08956794, 0.00731815, 0.01266064, 0.0006090624, 
    0.0003856527, 0.0007995427, 0.002388198, 0.03313753, 0.06335085, 
    0.0005891883, 0.0004332773, 3.258501e-05, 0.000199321, 0.0002786594, 
    0.0001714546, 0.0001592809, 0.0001675816, 0.0002771927, 0.0004258193, 
    0.003026936, 0.04451871, 0.05204863, 0.002221575, 8.546618e-05, 
    0.00103934, 0.0004358287, 0.001145236, 0.01523592,
  0.00488134, 0.00985314, 0.0007728518, 0.03025318, 1.49697e-06, 
    0.0002088435, 0.02436705, 2.970212e-05, -0.000626579, 0.0003278184, 
    2.831255e-05, 0.00276376, 0.0003576196, 0.0005631367, 0.001548649, 
    0.002761438, 0.003733966, 0.01100139, 0.0133005, 0.01274936, 0.002727694, 
    0.004793966, 0.124357, 0.01525958, 0.0002520084, 0.0008046365, 
    0.001062018, 0.00314882, 0.01983164,
  4.332605e-08, 5.594983e-08, 1.010115e-07, -4.875749e-06, 2.907696e-09, 
    0.04788462, 0.005605544, 0.0009548337, 0.04745258, 0.002105033, 
    0.00256675, 0.0004131743, 3.749117e-05, 0.0002805625, 0.0001948627, 
    3.945166e-05, 0.0003347545, 0.002073483, 0.01009548, 0.05599212, 
    0.003378348, 0.07128306, 0.0001957496, -0.001020737, 0.0005141629, 
    0.002020611, 0.009941597, 0.008865904, 3.29699e-07,
  3.443938e-07, 0.003083155, 0.0009036204, -1.838775e-06, 9.685556e-08, 
    4.928664e-09, -2.223727e-05, 0.2013748, 0.2610281, 0.03173558, 
    0.01137135, 0.001972022, 0.002142182, 0.001548935, 0.003801342, 
    0.001788521, 0.001615018, 0.002545612, 0.01860378, 0.2299119, 
    0.009262824, 0.009148744, 0.007753875, 0.001513015, 0.000771616, 
    0.0006529237, 0.002060196, 0.005941896, 0.01144129,
  0.002853013, 0.000729888, 0.002285581, 0.1649996, -0.0003925508, 
    -1.75741e-06, 0.03997265, -3.501706e-06, -0.0001766058, 0.01309032, 
    0.08338366, 0.04075347, 0.1092362, 0.09168971, 0.1595018, 0.1516438, 
    0.1045955, 0.04975083, 0.110572, -9.891496e-05, 0.0004437595, 0.03449037, 
    0.03418253, 0.07250101, 0.02171728, 0.02666478, 0.02010594, 0.007851336, 
    0.03941946,
  0.03335718, 0.1733502, 0.1176833, 0.08856852, 0.008570374, 0.006681235, 
    0.01280065, 0.1401086, 0.05445203, 0.08790135, 0.06115451, 0.1285293, 
    0.2646235, 0.2106906, 0.121389, 0.1611842, 0.1298908, 0.1193577, 
    0.1412945, 0.08671262, 0.0325145, 0.009372913, 0.05618439, 0.2104872, 
    0.1408057, 0.2219894, 0.1510383, 0.1159695, 0.04732099,
  0.0568509, 0.1707891, 0.08356194, 0.1031384, 0.1745027, 0.09571263, 
    0.06870803, 0.08906882, 0.1579616, 0.1648154, 0.1448106, 0.3550479, 
    0.2736332, 0.1455474, 0.1033507, 0.1435867, 0.3237019, 0.2777017, 
    0.2107798, 0.1014791, 0.05388995, 0.168326, 0.1599925, 0.3309403, 
    0.2254232, 0.1031821, 0.1981874, 0.09436998, 0.1035051,
  0.2091701, 0.07162326, 0.2778214, 0.1766406, 0.2734072, 0.2543312, 
    0.2571486, 0.2211849, 0.1720293, 0.1907378, 0.380513, 0.2592379, 
    0.2210194, 0.1853777, 0.2569845, 0.2332359, 0.2589317, 0.1377109, 
    0.1552781, 0.1407112, 0.3050805, 0.3276749, 0.3074723, 0.5087547, 
    0.1959607, 0.2085449, 0.244592, 0.07189749, 0.2245674,
  0.3330445, 0.1979678, 0.2711374, 0.3686793, 0.3515797, 0.3634382, 
    0.3822607, 0.3589551, 0.3151352, 0.3632222, 0.3198253, 0.2552766, 
    0.2933069, 0.3345177, 0.2820622, 0.3439654, 0.3724516, 0.371581, 
    0.3637574, 0.3645405, 0.2898034, 0.2001247, 0.3002318, 0.5015839, 
    0.2285869, 0.2082347, 0.1420781, 0.2474498, 0.2674426,
  0.002934038, 0.002616038, 0.002298038, 0.001980038, 0.001662038, 
    0.001344039, 0.001026039, 0.000568916, 0.001316641, 0.002064367, 
    0.002812092, 0.003559818, 0.004307543, 0.005055268, 0.005859287, 
    0.005486066, 0.005112846, 0.004739625, 0.004366405, 0.003993184, 
    0.003619964, 0.001500383, 0.001443877, 0.001387372, 0.001330868, 
    0.001274363, 0.001217858, 0.001161352, 0.003188438,
  0.1610906, 0.07620952, 0.03845834, 0.001322674, 8.337238e-05, 
    -4.550656e-05, -1.125374e-05, -3.730526e-06, 0, 0, 1.957395e-05, 
    0.005247859, 0.05964634, 0.007274087, 0.2270814, 0.2560956, 0.3133415, 
    0.2268437, 0.1152902, 0.3265097, 0.4335591, 0.4063494, 0.1062279, 
    0.07684942, 0.1769819, 0.3971704, 0.1823589, 0.09620941, 0.2696639,
  0.1745262, 0.06610703, 0.1118199, 0.01035917, 0.02168396, 0.005432013, 
    0.006012891, 0.07584591, 0.04164222, 0.0983033, 0.1537073, 0.09923603, 
    0.1090519, 0.09789057, 0.32894, 0.3286604, 0.2880421, 0.2612449, 
    0.2844464, 0.3076084, 0.2776436, 0.270472, 0.2927868, 0.4372506, 
    0.2142882, 0.3898957, 0.3726239, 0.3385864, 0.2521476,
  0.2909156, 0.2624708, 0.1912764, 0.07986518, 0.09689683, 0.1432575, 
    0.2131673, 0.1936805, 0.151542, 0.04496626, 0.05400513, 0.09430884, 
    0.1313659, 0.1504055, 0.110367, 0.1591973, 0.177893, 0.1887854, 0.121801, 
    0.09241351, 0.09767804, 0.075045, 0.1256904, 0.08226683, 0.1609577, 
    0.2454517, 0.2979373, 0.3023174, 0.2782535,
  0.1407389, 0.1500728, 0.1284692, 0.1290395, 0.1816592, 0.1593767, 0.149058, 
    0.08029734, 0.08455859, 0.07245457, 0.04616229, 0.0469196, 0.02675968, 
    0.04592022, 0.03502808, 0.0444894, 0.04376648, 0.07670953, 0.06864758, 
    0.07210138, 0.05860963, 0.06806807, 0.05470268, 0.08361216, 0.03382117, 
    0.1024369, 0.1333208, 0.1869131, 0.1553347,
  0.03796095, 0.009752802, 0.02227255, 0.06606084, 0.08938206, 0.04758881, 
    0.03451511, 0.02495558, 0.01731869, 0.007333602, 0.008967839, 
    0.002627549, 0.0009030087, 0.03060499, 0.07211168, 0.02888685, 
    0.01553376, 0.02302185, 0.04144243, 0.0234215, 0.02626295, 0.02284096, 
    0.02053413, 0.2337895, 0.01094898, 0.04405656, 0.03724134, 0.04542052, 
    0.06315763,
  0.005546215, 0.005141171, 0.003759464, 0.004977455, 0.006742258, 
    0.006894987, 0.004381824, 0.005499555, 0.0064251, 0.001920165, 
    0.001620613, 3.609073e-05, 0.007153162, 0.01161411, 0.02108305, 
    0.02551643, 0.01069088, 0.02806537, 0.02052191, 0.01525222, 0.005910451, 
    0.007381698, 0.008867893, 0.001299178, 0.01912165, 0.03256156, 
    0.01115046, 0.006800933, 0.005132324,
  0.02011066, 0.007455015, 0.0003306762, 0.001460589, -0.001656366, 
    0.0008396452, 0.0008685576, 0.0007078919, 0.003187083, 0.002548521, 
    4.740253e-09, 4.572251e-08, 0.0008279663, 0.007822372, 0.009632415, 
    0.001539036, 0.0006962101, 0.0005522785, 0.0002512451, 0.0002236926, 
    0.001375116, 0.003166898, 0.01172112, 0.0108808, 6.228512e-05, 
    0.04114569, 0.0005421178, 0.0009937861, 0.005673834,
  0.03675558, 0.02466962, 7.570022e-07, 0.03815999, 0.0001658432, 
    8.138167e-05, 0.0004201063, 0.0003621692, 0.0001967875, -0.0006152733, 
    0.004551655, 0.0002221302, 0.007776052, 0.0002925229, 4.1556e-05, 
    5.805582e-05, 4.84073e-05, 1.54851e-05, 1.178291e-05, 3.617703e-05, 
    0.0009279498, 0.00832459, 0.0358227, 0.001527103, 3.175895e-05, 
    3.759047e-08, 0.0004252217, 0.00200071, 0.01132534,
  0.004341895, 0.0700105, 0.0037448, 0.008776409, 0.0004192572, 0.0002505872, 
    0.0004037254, 0.001079604, 0.02572145, 0.06117655, 0.0003751382, 
    0.0003055913, 3.387456e-05, 0.0001298166, 0.0002050209, 0.0001230224, 
    0.00011101, 0.0001199621, 0.0001979377, 0.0002970523, 0.002065734, 
    0.03037567, 0.03856228, 0.002393407, 0.0004740382, 0.0007603246, 
    0.0003137865, 0.0008167813, 0.01076322,
  0.003537709, 0.006352606, 0.0003293918, 0.02289487, 1.598791e-07, 
    0.0001443818, 0.01028472, 2.05501e-05, -0.0004696161, 0.0001565234, 
    2.290668e-05, 0.001546408, 0.0002090061, 0.0003636322, 0.0008358087, 
    0.001404505, 0.001696312, 0.005388524, 0.006020721, 0.005488359, 
    0.001241645, 0.002184204, 0.1079542, 0.02454773, 0.0001748036, 
    0.0005244416, 0.0006196667, 0.001779136, 0.01790052,
  4.243586e-08, 5.446264e-08, 1.956454e-07, -2.626721e-06, 6.570245e-10, 
    0.03183872, 0.003766056, 0.0004033704, 0.04355975, 0.0007463339, 
    0.001154959, 0.0002578813, 2.931562e-05, 0.0001427732, 0.0001436243, 
    2.607424e-05, 0.0002496527, 0.001486518, 0.006983588, 0.0355493, 
    0.002251001, 0.06084874, 0.0001438312, -0.000983546, 0.0003643364, 
    0.00141075, 0.006836777, 0.00623538, 3.263019e-07,
  3.267956e-07, 0.001895179, 0.000457767, -1.293206e-06, 9.254346e-08, 
    5.050695e-09, -4.56399e-06, 0.1924581, 0.2398407, 0.01578331, 
    0.005147229, 0.001132533, 0.0013359, 0.0009384258, 0.002255548, 
    0.001327169, 0.001173973, 0.001402057, 0.01350925, 0.1945065, 
    0.007412976, 0.01109179, 0.00774226, 0.0008897761, 0.000562837, 
    0.0004915987, 0.001451281, 0.004223487, 0.008842548,
  0.002614192, 0.0003043483, 0.001853154, 0.1488165, -0.0003376071, 
    -1.071801e-06, 0.03518821, -2.845005e-06, -0.0001556591, 0.009184758, 
    0.07587083, 0.02575232, 0.07876668, 0.05984714, 0.110599, 0.1158809, 
    0.06787832, 0.03083304, 0.08591861, -0.0001220948, 0.0004150078, 
    0.02951699, 0.02440476, 0.05143975, 0.01263633, 0.01199457, 0.01201205, 
    0.004569023, 0.03065492,
  0.02790728, 0.1566552, 0.09830368, 0.06796356, 0.006490131, 0.00485292, 
    0.00953912, 0.1255952, 0.0496757, 0.08041157, 0.05218592, 0.1178397, 
    0.2018516, 0.1537718, 0.08496454, 0.1183697, 0.09485683, 0.08907713, 
    0.1024803, 0.08062987, 0.02643653, 0.007465923, 0.04187705, 0.18267, 
    0.1228269, 0.1872596, 0.110197, 0.07877641, 0.02601431,
  0.03429984, 0.1475082, 0.07075257, 0.08863072, 0.1561674, 0.08531775, 
    0.06684655, 0.08338848, 0.1464469, 0.1454587, 0.1287462, 0.320939, 
    0.2452045, 0.1152316, 0.07252645, 0.1073135, 0.292263, 0.2452453, 
    0.1796197, 0.09703776, 0.04608571, 0.1512847, 0.1106747, 0.2864664, 
    0.1680677, 0.07988054, 0.1453425, 0.06137721, 0.07176155,
  0.1510207, 0.04563023, 0.2381247, 0.1377694, 0.2185523, 0.2347154, 
    0.2265369, 0.1850081, 0.149851, 0.1646812, 0.3413446, 0.2247205, 
    0.1932679, 0.1558535, 0.2278719, 0.1966155, 0.227241, 0.1156964, 
    0.1422846, 0.1108634, 0.268788, 0.2979459, 0.2592376, 0.4667439, 
    0.1656125, 0.1737592, 0.301477, 0.0633624, 0.164262,
  0.2881562, 0.1715532, 0.2476558, 0.3029453, 0.2948164, 0.3238411, 
    0.3270094, 0.2967885, 0.2563834, 0.2903196, 0.2611259, 0.2097282, 
    0.2558788, 0.2799698, 0.2328264, 0.2733348, 0.3014063, 0.3031743, 
    0.2841941, 0.3025358, 0.2414221, 0.1759632, 0.2628367, 0.4826691, 
    0.2116829, 0.1707979, 0.1298408, 0.232293, 0.2456003,
  0.002596252, 0.002384338, 0.002172425, 0.001960511, 0.001748597, 
    0.001536683, 0.001324769, 0.001301845, 0.001628738, 0.00195563, 
    0.002282522, 0.002609415, 0.002936307, 0.003263199, 0.00191772, 
    0.001845153, 0.001772586, 0.001700018, 0.001627451, 0.001554884, 
    0.001482317, 0.001644555, 0.001602144, 0.001559733, 0.001517321, 
    0.00147491, 0.001432499, 0.001390088, 0.002765783,
  0.105376, 0.05251485, 0.01796146, 0.0009102614, 9.786032e-05, -3.38977e-05, 
    -3.889091e-06, 0, 0, 0, 4.679741e-05, 0.004841651, 0.03327391, 
    0.007469258, 0.2242991, 0.1978484, 0.2646521, 0.2446704, 0.127692, 
    0.3472591, 0.4403311, 0.4395891, 0.1057115, 0.07264496, 0.1562695, 
    0.3493662, 0.1802782, 0.1019857, 0.2014898,
  0.1705736, 0.06754848, 0.10597, 0.009916702, 0.01693694, 0.004533617, 
    0.006160171, 0.07027902, 0.03151315, 0.08817104, 0.1280811, 0.08247763, 
    0.104995, 0.0909303, 0.3181164, 0.3080032, 0.2676597, 0.2379128, 
    0.2561362, 0.2845519, 0.251624, 0.2538763, 0.2719931, 0.4139014, 
    0.2056098, 0.3438004, 0.338978, 0.3001933, 0.2259779,
  0.2622477, 0.2419705, 0.1789266, 0.0730243, 0.08862568, 0.136178, 0.202177, 
    0.1790645, 0.1411539, 0.03854301, 0.04731515, 0.08337301, 0.1188204, 
    0.1312993, 0.09428418, 0.1384589, 0.1587543, 0.1644556, 0.1075069, 
    0.08099861, 0.08459133, 0.06167216, 0.1056713, 0.06894693, 0.146191, 
    0.2260659, 0.282896, 0.2834307, 0.2491984,
  0.1212981, 0.1264899, 0.108865, 0.1090489, 0.1600232, 0.1347767, 0.1297469, 
    0.07006801, 0.07428576, 0.05999606, 0.03667053, 0.03662544, 0.02182811, 
    0.03557894, 0.02727506, 0.0338745, 0.03469768, 0.05917478, 0.05498125, 
    0.05832642, 0.04438882, 0.05230299, 0.04403342, 0.09554572, 0.0270475, 
    0.08501393, 0.1102379, 0.1573237, 0.1343066,
  0.02943381, 0.006954442, 0.01665318, 0.05184363, 0.06675214, 0.03315328, 
    0.02509625, 0.0178733, 0.01255197, 0.005144784, 0.006998838, 0.002054356, 
    0.0007197885, 0.02255787, 0.05950315, 0.02145133, 0.01166864, 0.01768163, 
    0.0317447, 0.01738587, 0.01894512, 0.01636118, 0.01399425, 0.2285744, 
    0.01004229, 0.03567439, 0.02669187, 0.0348778, 0.04412705,
  0.004728835, 0.004022381, 0.006328119, 0.003558868, 0.004879807, 
    0.005477035, 0.003773651, 0.004751866, 0.005499078, 0.001609863, 
    0.001261982, 3.013071e-05, 0.0092515, 0.006714164, 0.01401616, 0.0157163, 
    0.006629543, 0.01944884, 0.01341159, 0.009249841, 0.004148794, 
    0.005376383, 0.007592066, 0.001151842, 0.02282304, 0.02251158, 
    0.006829512, 0.0047889, 0.003766412,
  0.01692857, 0.006275828, 0.0002156316, 0.001202514, -0.001529826, 
    0.0005345027, 0.0006647854, 0.0006041426, 0.002678112, 0.002005032, 
    4.976628e-09, 4.631089e-08, 0.0006938627, 0.004796874, 0.00555486, 
    0.001196996, 0.0005629401, 0.0004327414, 0.0001932998, 0.0001739435, 
    0.001136017, 0.00263598, 0.009890867, 0.009514339, 3.983778e-05, 
    0.05409951, 0.0004675632, 0.000822085, 0.00466543,
  0.02974863, 0.01877844, 2.711934e-05, 0.03043302, 0.0001292992, 
    6.607663e-05, 0.0003303746, 0.0002525204, 0.0001667711, -0.0005025648, 
    0.003663765, 0.0001370681, 0.005149849, 0.0002230871, 3.448178e-05, 
    4.518047e-05, 3.868475e-05, 1.319864e-05, 9.899512e-06, 3.077178e-05, 
    0.000774201, 0.006896401, 0.02934891, 0.02320418, -0.0001368881, 
    7.829954e-08, 0.0003629212, 0.001671224, 0.009298288,
  0.003472346, 0.1113394, 0.005876204, 0.008096944, 0.0003292596, 
    0.0001966326, 0.0002788221, 0.0006849193, 0.03279375, 0.07682419, 
    0.0002956763, 0.0002450988, 3.194434e-05, 9.436214e-05, 0.0001684023, 
    0.0001005893, 9.051516e-05, 9.875485e-05, 0.0001656619, 0.0002412552, 
    0.001611887, 0.02390128, 0.03174774, 0.00743626, 0.008896923, 
    0.0006263375, 0.0002540614, 0.0006633712, 0.008613924,
  0.01389731, 0.005875775, 0.0002398184, 0.01879934, -1.764389e-07, 
    0.0001183763, 0.0081633, 2.205116e-05, -0.00251492, 0.0001061548, 
    2.041561e-05, 0.001103582, 0.000149309, 0.0002871861, 0.0005781076, 
    0.0009324611, 0.0009995253, 0.003298092, 0.003601329, 0.00322804, 
    0.0008065756, 0.001351951, 0.1681031, 0.03381877, 0.0001397772, 
    0.0004146313, 0.0004533317, 0.001343592, 0.04114576,
  4.193323e-08, 5.361244e-08, 1.915632e-07, -1.742812e-06, -2.349951e-09, 
    0.02400865, 0.006387298, 0.0002397128, 0.08792168, -0.0002570375, 
    0.0007617762, 0.0001891159, 2.440769e-05, 9.790799e-05, 0.0001185554, 
    2.088529e-05, 0.0002076192, 0.001204906, 0.005551052, 0.02399292, 
    0.00178149, 0.05720038, 0.0001181728, -0.001723776, 0.0002945828, 
    0.001136619, 0.005406935, 0.005008041, 3.279649e-07,
  3.20697e-07, 0.00116417, 0.000168014, -7.681957e-07, 8.953988e-08, 
    5.131276e-09, 0.0004821274, 0.2118967, 0.2437821, 0.01220261, 
    0.003509409, 0.0008241027, 0.001002937, 0.0007800626, 0.001697367, 
    0.001101317, 0.0009696586, 0.001053858, 0.01104706, 0.1723732, 
    0.007305696, 0.04192092, 0.02725017, 0.0006615417, 0.0004611012, 
    0.0004098393, 0.001116756, 0.003500655, 0.006860832,
  0.003283849, -7.324597e-05, 0.001660037, 0.1409272, -0.0003159053, 
    -7.18279e-07, 0.03127336, -2.811606e-06, -0.0001417714, 0.007006565, 
    0.08880006, 0.01402484, 0.06174459, 0.03931408, 0.07944445, 0.08410771, 
    0.04478681, 0.01950002, 0.06224018, -0.0001952107, 0.0003902782, 
    0.02821468, 0.02840114, 0.03673097, 0.008324106, 0.00782819, 0.008035191, 
    0.003407311, 0.02625275,
  0.02417996, 0.1609573, 0.09605683, 0.06621003, 0.005458427, 0.003872102, 
    0.008080946, 0.1247521, 0.0550339, 0.08713989, 0.06998407, 0.1343911, 
    0.1608768, 0.1121073, 0.06002498, 0.08866131, 0.07049435, 0.06840295, 
    0.0704333, 0.08256869, 0.02467717, 0.007411915, 0.04779936, 0.199867, 
    0.1169112, 0.1487569, 0.08221481, 0.05554338, 0.01736699,
  0.02347351, 0.1554027, 0.07042623, 0.08608415, 0.1765047, 0.103264, 
    0.09286677, 0.1144578, 0.1774188, 0.1691082, 0.1389377, 0.3217874, 
    0.2431914, 0.1186292, 0.05856074, 0.08430865, 0.3018844, 0.2408487, 
    0.1901197, 0.102784, 0.04901949, 0.1664815, 0.07966308, 0.279991, 
    0.1318077, 0.06786311, 0.1177798, 0.04522204, 0.05232713,
  0.110281, 0.03223731, 0.2342202, 0.101621, 0.1717434, 0.2125323, 0.2336094, 
    0.1820748, 0.1498761, 0.1667361, 0.351512, 0.2325107, 0.1900254, 
    0.1335622, 0.2033661, 0.1736731, 0.2125544, 0.1082006, 0.1308237, 
    0.09142415, 0.2408467, 0.2712071, 0.2450939, 0.4347994, 0.135121, 
    0.1527294, 0.3680051, 0.0550643, 0.1287003,
  0.2689984, 0.1515133, 0.2270271, 0.2592645, 0.2609915, 0.2962985, 
    0.2892244, 0.2610482, 0.2196645, 0.2544477, 0.2196346, 0.180237, 
    0.2187798, 0.2365726, 0.1977849, 0.2247463, 0.2604181, 0.2629024, 
    0.243546, 0.2619882, 0.2042587, 0.1664079, 0.246944, 0.455097, 0.1946045, 
    0.1519052, 0.1306085, 0.2219917, 0.2254549 ;

 average_DT = 730 ;

 average_T1 = 259 ;

 average_T2 = 989 ;

 climatology_bounds =
  259, 989 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
