netcdf atmos.1980-1981.alb_sfc {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:bounds = "time_bnds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double time_bnds(time, bnds) ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 11:53:26 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.nc reduced/atmos.1980-1981.alb_sfc.nc\n",
			"Mon Aug 25 14:39:16 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  37.45993, 37.45993, 37.45993, 37.45993, 37.45993, 37.45993, 37.45993, 
    37.45878, 37.45878, 37.45878, 37.45878, 37.45878, 37.45878, 37.45878, 
    37.44279, 37.44279, 37.44279, 37.44279, 37.44279, 37.44279, 37.44279, 
    37.45418, 37.45418, 37.45418, 37.45418, 37.45418, 37.45418, 37.45418, 
    37.45993,
  38.03535, 37.95234, 37.91778, 37.87039, 37.86663, 37.86129, 37.85198, 
    37.84583, 37.85187, 37.87751, 37.90581, 37.9373, 37.99785, 37.73974, 
    37.60143, 37.11834, 37.33641, 36.96517, 36.8639, 37.77762, 38.04186, 
    38.14217, 38.0373, 36.40692, 37.00923, 36.1885, 36.81783, 36.80325, 
    38.07371,
  30.33605, 28.33545, 29.43709, 36.53866, 38.61345, 38.64645, 35.0915, 
    38.64052, 38.59653, 38.62041, 38.59209, 38.57387, 37.98376, 31.91109, 
    24.97525, 23.30625, 22.75709, 24.0446, 22.65203, 26.55817, 27.58533, 
    25.56068, 34.9426, 35.59814, 37.40865, 31.40498, 24.89729, 22.5753, 
    25.76643,
  19.26042, 20.85573, 10.1349, 5.2674, 4.797372, 6.081092, 14.62923, 
    8.422602, 7.176382, 4.097719, 4.114795, 3.977645, 3.761458, 3.870051, 
    4.036924, 3.925717, 3.800187, 3.799801, 3.98992, 4.127749, 4.204319, 
    4.199813, 4.13286, 4.054861, 6.229377, 13.05438, 19.62386, 17.92866, 
    19.35307,
  3.774479, 3.838792, 3.8345, 3.87201, 3.855156, 3.858616, 3.884374, 3.96393, 
    3.984507, 3.976398, 3.965414, 3.944838, 3.946605, 3.931716, 3.915069, 
    3.916279, 3.878623, 3.847686, 3.908394, 3.931341, 3.960512, 3.984962, 
    3.935166, 8.041118, 4.38075, 3.979097, 3.761329, 3.785665, 3.761953,
  3.777115, 3.893794, 4.024122, 3.887876, 3.820014, 3.869495, 3.854475, 
    3.81674, 3.788136, 3.916249, 3.900683, 4.005403, 4.1674, 3.969128, 
    10.48656, 3.886335, 3.874708, 3.812052, 3.787953, 3.779731, 3.754786, 
    3.787159, 3.868348, 9.646874, 4.305488, 3.938987, 3.833462, 3.805404, 
    3.776341,
  3.824853, 4.034652, 12.08973, 3.862848, 3.851677, 3.818546, 3.832149, 
    3.84521, 3.817913, 4.103725, 9.49978, 14.2443, 10.35399, 3.956338, 
    3.860187, 3.799219, 3.771741, 3.67976, 3.578305, 3.678083, 3.81165, 
    3.91877, 3.792727, 4.46473, 8.968763, 3.73048, 3.744849, 3.843025, 
    3.859042,
  3.479322, 9.758091, 10.61068, 3.762444, 3.682558, 3.727141, 3.75803, 
    3.737916, 3.636152, 3.86576, 11.94082, 11.60274, 3.767761, 3.649697, 
    3.587939, 3.60775, 3.590988, 3.599503, 3.723098, 3.841023, 3.83588, 
    3.681329, 3.397042, 3.581701, 8.992791, 9.038381, 3.760325, 3.780236, 
    3.671401,
  3.292887, 6.306999, 8.915585, 9.098597, 3.478494, 3.449342, 3.416554, 
    3.407036, 3.401942, 3.434816, 4.683577, 3.417869, 4.289854, 3.361482, 
    3.399756, 3.489893, 3.55491, 3.709733, 3.699762, 3.798621, 3.698399, 
    3.557586, 3.336347, 8.671864, 8.58602, 9.422429, 3.730154, 3.629855, 
    3.527236,
  3.180231, 8.521408, 8.35378, 9.900547, 3.456246, 3.366768, 3.304661, 
    3.270167, 8.574446, 8.299625, 3.310154, 3.325699, 3.322168, 3.417664, 
    3.443453, 3.564374, 3.598329, 3.748667, 3.628184, 3.715953, 3.558012, 
    3.38276, 3.299225, 8.42738, 8.488513, 3.383074, 3.39954, 3.384226, 
    3.238375,
  9.847279, 10.18859, 10.28258, 9.513283, 14.71262, 3.366705, 5.187101, 
    3.337696, 3.501173, 3.311682, 4.186483, 3.312178, 3.286719, 3.342498, 
    3.364689, 3.36715, 3.434729, 3.437693, 3.423315, 3.371299, 3.323021, 
    3.340537, 8.718559, 7.439555, 3.428066, 3.358228, 3.190545, 3.260875, 
    8.828611,
  17.63745, 20.10217, 22.0703, 3.527292, 22.25309, 3.549904, 10.52603, 
    3.553025, 9.142807, 3.361149, 3.445198, 3.52735, 3.605648, 3.695551, 
    3.739467, 3.761205, 3.754842, 3.753906, 3.550002, 3.494633, 3.673942, 
    6.306129, 3.618136, 4.300377, 3.645838, 3.657512, 3.528582, 3.457198, 
    22.85155,
  22.90774, 19.02185, 19.85403, 18.55453, 12.37888, 14.15996, 12.1651, 
    16.85423, 9.138701, 10.30511, 3.500245, 3.629782, 3.695691, 3.703731, 
    3.711864, 3.706154, 3.771835, 3.77705, 3.658345, 3.915842, 11.019, 
    11.59688, 9.381607, 3.62171, 3.684407, 3.755291, 3.811707, 3.79545, 
    10.74925,
  6.862579, 4.136683, 6.067963, 12.79179, 1.946488, 14.24467, 14.70746, 
    14.73052, 12.52858, 13.45459, 8.335635, 3.785952, 3.759634, 3.747746, 
    3.740135, 3.688364, 3.593117, 3.593329, 3.696813, 11.94578, 14.73228, 
    14.42592, 13.59047, 4.557602, 3.680932, 3.695635, 3.749509, 3.837311, 
    5.125711,
  5.63048, 12.25049, 13.79066, 16.13728, 16.06226, 17.23173, 9.679915, 
    21.90686, 10.53441, 7.279898, 7.830172, 12.54683, 6.740848, 3.930022, 
    3.892049, 3.857399, 3.802904, 3.819779, 3.934446, 13.97994, 12.56317, 
    15.15049, 12.95065, 16.43394, 7.620394, 3.792377, 3.87215, 3.944572, 
    4.027317,
  4.240577, 11.10437, 10.9065, 12.15293, 12.39044, 12.3108, 14.09149, 
    15.70507, 13.61311, 13.60658, 12.02155, 23.38995, 24.87297, 17.58506, 
    4.606345, 13.32736, 17.63372, 13.94056, 21.50202, 11.44591, 12.20459, 
    22.96399, 24.61838, 23.8048, 3.84124, 8.560878, 4.162157, 4.112668, 
    4.143772,
  3.818251, 4.147723, 12.67614, 3.950956, 13.39264, 27.10033, 23.90227, 
    23.81619, 23.6854, 24.00868, 15.72201, 13.24643, 22.39485, 29.01567, 
    32.92902, 24.35602, 24.32892, 23.49706, 24.72709, 23.5178, 25.31774, 
    28.98533, 25.82146, 30.33984, 21.66751, 37.66063, 38.99792, 24.06214, 
    3.857056,
  33.20492, 26.20865, 29.51533, 30.61344, 27.12186, 31.48092, 35.97458, 
    32.51833, 35.11747, 37.20291, 37.23371, 37.21825, 37.22918, 37.11561, 
    37.14951, 37.11675, 36.90792, 36.77555, 36.84005, 36.83963, 36.87662, 
    33.82414, 32.9637, 35.65375, 37.11012, 37.24373, 38.22337, 35.10448, 
    33.50555 ;

 average_DT = 720 ;

 average_T1 = 350.5 ;

 average_T2 = 1080.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 715.5 ;

 time_bnds =
  350.5, 1080.5 ;
}
