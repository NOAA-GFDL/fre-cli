netcdf atmos_cmip.ua_unmsk {
dimensions:
	bnds = 2 ;
	lat = 10 ;
	lon = 10 ;
	plev19 = 19 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double bnds(bnds) ;
		bnds:long_name = "vertex number" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
		lat_bnds:long_name = "latitude bounds" ;
		lat_bnds:units = "degrees_N" ;
		lat_bnds:axis = "Y" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
		lon_bnds:long_name = "longitude bounds" ;
		lon_bnds:units = "degrees_E" ;
		lon_bnds:axis = "X" ;
	double plev19(plev19) ;
		plev19:units = "Pa" ;
		plev19:long_name = "pressure" ;
		plev19:axis = "Z" ;
		plev19:positive = "down" ;
	double time(time) ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, bnds) ;
		time_bnds:units = "days since 1979-01-01 00:00:00" ;
		time_bnds:long_name = "time axis boundaries" ;
	float ua_unmsk(time, plev19, lat, lon) ;
		ua_unmsk:_FillValue = 1.e+20f ;
		ua_unmsk:missing_value = 1.e+20f ;
		ua_unmsk:units = "m s-1" ;
		ua_unmsk:long_name = "Eastward Wind" ;
		ua_unmsk:cell_methods = "time: mean" ;
		ua_unmsk:cell_measures = "area: area" ;
		ua_unmsk:standard_name = "eastward_wind" ;
		ua_unmsk:interp_method = "conserve_order2" ;
        ua_unmsk:pressure_mask = ".false." ;

// global attributes:
		:title = "c96L65_am5f9d7r0_amip" ;
		:associated_files = "area: 20050101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Thu Jun 26 22:27:29 2025" ;
		:hostname = "pp208" ;
		:history = "Tue Jul  1 23:47:57 2025: ncks -d lat,10,19 -d lon,10,19 -d time,0,0 atmos_cmip.200501-200512.ua_unmsk.nc atmos_cmip.ua_unmsk.nc\n",
			"fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_file 20050101.atmos_month_cmip --interp_method conserve_order2 --remap_file .fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field tas,ts,psl,ps,uas,height10m,vas,sfcWind,hurs,height2m,huss,pr,prsn,prc,evspsbl,tauu,tauv,hfls,hfss,rlds,rlus,rsds,rsus,rsdscs,rsuscs,rldscs,rsdt,rsut,rlut,rlutcs,rsutcs,prw,clt,clwvi,clivi,rtmt,ccb,cct,ci,sci,ta_unmsk,ua_unmsk,va_unmsk,hus_unmsk,hur_unmsk,wap_unmsk,zg_unmsk,ap,b,ap_bnds,b_bnds,lev_bnds,utendnogw,utendogw,time_bnds --output_file out.nc" ;
		:external_variables = "area" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 bnds = 1, 2 ;

 lat = -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5 ;

 lat_bnds =
  -80, -79,
  -79, -78,
  -78, -77,
  -77, -76,
  -76, -75,
  -75, -74,
  -74, -73,
  -73, -72,
  -72, -71,
  -71, -70 ;

 lon = 13.125, 14.375, 15.625, 16.875, 18.125, 19.375, 20.625, 21.875, 
    23.125, 24.375 ;

 lon_bnds =
  12.5, 13.75,
  13.75, 15,
  15, 16.25,
  16.25, 17.5,
  17.5, 18.75,
  18.75, 20,
  20, 21.25,
  21.25, 22.5,
  22.5, 23.75,
  23.75, 25 ;

 plev19 = 100000, 92500, 85000, 70000, 60000, 50000, 40000, 30000, 25000, 
    20000, 15000, 10000, 7000, 5000, 3000, 2000, 1000, 500, 100 ;

 time = 9512.5 ;

 time_bnds =
  9497, 9528 ;

 ua_unmsk =
  -0.3975942, -0.2708012, -0.1832284, -0.09187625, 0.001559797, 0.07204625, 
    0.0783459, 0.09246785, 0.1097215, 0.1203732,
  -0.5745555, -0.5160208, -0.4475087, -0.3612338, -0.3011235, -0.2559909, 
    -0.2050162, -0.1434478, -0.08277573, -0.06627619,
  -0.6454812, -0.6330528, -0.6397436, -0.6381702, -0.6238125, -0.5942059, 
    -0.5442353, -0.5295258, -0.5248909, -0.527373,
  -0.8545123, -0.8994937, -0.9365253, -1.021321, -1.10686, -1.154233, 
    -1.184383, -1.207665, -1.235654, -1.261622,
  -1.426775, -1.437999, -1.512454, -1.57849, -1.644708, -1.758953, -1.863996, 
    -1.918497, -1.973612, -2.010429,
  -2.151411, -2.133208, -2.145542, -2.198483, -2.335929, -2.401734, 
    -2.460874, -2.553266, -2.576532, -2.571083,
  -2.586592, -2.56783, -2.469594, -2.440526, -2.463234, -2.546937, -2.664745, 
    -2.762299, -2.825696, -2.793565,
  -2.590438, -2.542438, -2.476797, -2.352731, -2.229772, -2.188571, 
    -2.246655, -2.410638, -2.534509, -2.572949,
  -1.956838, -1.938947, -1.808724, -1.627707, -1.515042, -1.380297, 
    -1.431068, -1.480767, -1.527824, -1.59102,
  -0.5315368, -0.5231183, -0.4564048, -0.3944708, -0.1738839, -0.07352839, 
    0.01055507, 0.1166717, 0.1312627, 0.2858787,
  -0.3975942, -0.2708012, -0.1832284, -0.09187625, 0.001559797, 0.07204625, 
    0.0783459, 0.09246785, 0.1097215, 0.1203732,
  -0.5745555, -0.5160208, -0.4475087, -0.3612338, -0.3011235, -0.2559909, 
    -0.2050162, -0.1434478, -0.08277573, -0.06627619,
  -0.6454812, -0.6330528, -0.6397436, -0.6381702, -0.6238125, -0.5942059, 
    -0.5442353, -0.5295258, -0.5248909, -0.527373,
  -0.8545123, -0.8994937, -0.9365253, -1.021321, -1.10686, -1.154233, 
    -1.184383, -1.207665, -1.235654, -1.261622,
  -1.426775, -1.437999, -1.512454, -1.57849, -1.644708, -1.758953, -1.863996, 
    -1.918497, -1.973612, -2.010429,
  -2.151411, -2.133208, -2.145542, -2.198483, -2.335929, -2.401734, 
    -2.460874, -2.553266, -2.576532, -2.571083,
  -2.586592, -2.56783, -2.469594, -2.440526, -2.463234, -2.546937, -2.664745, 
    -2.76217, -2.823994, -2.793565,
  -2.56729, -2.51979, -2.476788, -2.342977, -2.180678, -2.173315, -2.202794, 
    -2.382988, -2.51635, -2.56469,
  -2.164203, -2.002625, -1.769979, -1.522183, -1.529329, -1.788184, 
    -1.570996, -1.601109, -2.148522, -2.238381,
  -1.765279, -1.833698, -1.684174, -1.374214, -1.259788, -1.473578, 
    -1.366698, -1.105641, -1.151468, -1.052101,
  -0.3975942, -0.2708012, -0.1832284, -0.09187625, 0.001559797, 0.07204625, 
    0.0783459, 0.09246785, 0.1097215, 0.1203732,
  -0.5745555, -0.5160208, -0.4475087, -0.3612338, -0.3011235, -0.2559909, 
    -0.2050162, -0.1434478, -0.08277573, -0.06627619,
  -0.6454812, -0.6330528, -0.6397436, -0.6381702, -0.6238125, -0.5942059, 
    -0.5442353, -0.5295258, -0.5248909, -0.527373,
  -0.8545123, -0.8994937, -0.9365253, -1.021321, -1.10686, -1.154233, 
    -1.184383, -1.207665, -1.235654, -1.261622,
  -1.426775, -1.437999, -1.512454, -1.57849, -1.644708, -1.758953, -1.863996, 
    -1.918497, -1.973612, -2.010429,
  -2.151411, -2.133208, -2.145542, -2.198483, -2.335929, -2.401734, 
    -2.460874, -2.553266, -2.576532, -2.571083,
  -2.586592, -2.559288, -2.461631, -2.440526, -2.46086, -2.4672, -2.609189, 
    -2.751828, -2.816938, -2.793565,
  -2.410764, -2.404498, -2.467111, -2.314096, -1.887833, -2.113094, 
    -2.547507, -2.529567, -2.430087, -2.455852,
  -2.803633, -2.214195, -2.758755, -3.378312, -3.186033, -3.65111, -4.398364, 
    -4.396877, -4.207345, -3.572534,
  -5.248218, -4.912538, -4.553966, -4.296717, -4.063207, -4.280607, 
    -4.150732, -3.721014, -3.682456, -3.493971,
  -0.4638011, -0.2794998, -0.1847423, -0.1013127, -0.01874243, 0.05095983, 
    0.07407396, 0.09246785, 0.1097215, 0.1203732,
  -0.5747783, -0.5167099, -0.4489113, -0.3624935, -0.3011871, -0.2559909, 
    -0.2050162, -0.1434478, -0.08277573, -0.06627619,
  -0.6454812, -0.6330528, -0.6397436, -0.6381702, -0.6238125, -0.5942059, 
    -0.5442353, -0.5295258, -0.5248909, -0.527373,
  -0.8545123, -0.8994937, -0.9365253, -1.021321, -1.10686, -1.154233, 
    -1.184383, -1.207665, -1.235654, -1.261622,
  -1.426775, -1.437999, -1.512454, -1.57849, -1.644708, -1.758953, -1.863996, 
    -1.918497, -1.973612, -2.010429,
  -2.046627, -2.075339, -2.133872, -2.192768, -2.29642, -2.385374, -2.421421, 
    -2.375845, -2.522865, -2.570514,
  -2.329157, -2.661558, -2.550557, -2.222389, -2.452235, -2.64684, -2.825807, 
    -3.021084, -2.930932, -2.340356,
  -4.449573, -5.811647, -6.238008, -5.904782, -5.536724, -5.204103, 
    -5.139505, -6.584569, -7.315174, -6.587632,
  -7.759037, -7.923704, -7.657747, -7.342247, -7.189469, -6.957999, 
    -6.869977, -6.911683, -6.890206, -6.571945,
  -5.766199, -5.629292, -5.500316, -5.457587, -5.137841, -4.946566, 
    -4.747363, -4.453594, -4.333026, -4.211693,
  1.063227, 1.156564, 1.210127, 1.265683, 1.325263, 1.37135, 1.379399, 
    1.395321, 1.408047, 1.413615,
  0.8057297, 0.823011, 0.8517545, 0.8839636, 0.8734952, 0.8716547, 0.8792083, 
    0.8959213, 0.933274, 0.9308779,
  0.3776965, 0.3511574, 0.3064211, 0.2771505, 0.2723292, 0.26952, 0.2818037, 
    0.2319987, 0.165376, 0.1122594,
  -0.2686788, -0.3904975, -0.4879307, -0.5713966, -0.6487127, -0.7579689, 
    -0.879656, -1.019151, -1.160378, -1.290107,
  -1.44353, -1.544772, -1.67499, -1.812897, -1.98716, -2.274205, -2.556359, 
    -2.771371, -2.97445, -3.201544,
  -3.11445, -3.268162, -3.425929, -3.644483, -3.970347, -4.194717, -4.426955, 
    -4.785159, -4.986393, -5.121875,
  -4.842557, -4.942987, -5.010421, -5.153152, -5.254729, -5.326348, 
    -5.648958, -6.018217, -6.451276, -6.772595,
  -6.110239, -6.028393, -5.95482, -5.914704, -5.883089, -5.694447, -5.721324, 
    -5.85588, -6.038979, -6.222065,
  -6.000411, -6.046391, -5.883338, -5.710005, -5.577016, -5.360312, 
    -5.450391, -5.419651, -5.09429, -4.927251,
  -4.122381, -4.0073, -3.920688, -3.890532, -3.619308, -3.348911, -3.164834, 
    -3.032901, -2.999816, -2.981941,
  1.021295, 1.058732, 1.055263, 1.055828, 1.06735, 1.085502, 1.072789, 
    1.066372, 1.055719, 1.03737,
  0.5644462, 0.5258871, 0.505933, 0.5047766, 0.4665931, 0.4326979, 0.4054725, 
    0.3554713, 0.3202047, 0.2826239,
  -0.09909091, -0.1695052, -0.2423104, -0.308107, -0.3618009, -0.4362217, 
    -0.5038798, -0.5690737, -0.6322247, -0.6912587,
  -0.8452172, -0.9907208, -1.12432, -1.275977, -1.407145, -1.514558, 
    -1.611202, -1.70489, -1.787341, -1.840466,
  -1.660944, -1.836267, -2.043581, -2.208486, -2.365314, -2.544751, 
    -2.701359, -2.791034, -2.877407, -2.950873,
  -2.49663, -2.691726, -2.876794, -3.089699, -3.315934, -3.422023, -3.487426, 
    -3.497974, -3.590583, -3.699841,
  -3.409052, -3.454748, -3.579855, -3.723231, -3.777681, -3.849489, 
    -3.761075, -3.758978, -3.830392, -3.977781,
  -4.332948, -4.30478, -4.268668, -4.142052, -4.038466, -3.906201, -3.853595, 
    -3.97838, -4.061214, -3.96847,
  -4.037989, -3.923016, -3.725387, -3.504999, -3.335768, -3.048127, 
    -2.881483, -2.777315, -2.57696, -2.525698,
  -2.675588, -2.521989, -2.357147, -2.217182, -1.92482, -1.59737, -1.311503, 
    -1.052147, -0.8554193, -0.7043628,
  0.868393, 0.8096983, 0.7342755, 0.6706711, 0.6231919, 0.5861326, 0.5235301, 
    0.4832453, 0.4458269, 0.403123,
  0.3249699, 0.203376, 0.09710471, 0.005840228, -0.09959703, -0.186581, 
    -0.2659973, -0.3638777, -0.4377598, -0.5044919,
  -0.4682975, -0.6448929, -0.7865676, -0.9014125, -1.010695, -1.141248, 
    -1.26495, -1.354475, -1.432743, -1.508723,
  -1.302762, -1.487646, -1.667504, -1.870815, -2.038251, -2.165048, 
    -2.268736, -2.35599, -2.422225, -2.462221,
  -1.897165, -2.089815, -2.293899, -2.467101, -2.626223, -2.795213, 
    -2.938092, -3.009527, -3.077491, -3.088423,
  -2.338803, -2.44815, -2.576407, -2.714023, -2.881914, -2.990129, -3.088588, 
    -3.162073, -3.200975, -3.280721,
  -2.629382, -2.617197, -2.644625, -2.714817, -2.728057, -2.764721, 
    -2.755495, -2.804715, -2.900975, -3.060241,
  -2.806314, -2.699975, -2.604603, -2.467385, -2.316504, -2.181494, 
    -2.104434, -2.068235, -2.089983, -2.092961,
  -2.350076, -2.191863, -2.015235, -1.808842, -1.591449, -1.298141, 
    -1.055869, -0.8611979, -0.6329716, -0.4672858,
  -1.417739, -1.253469, -1.085745, -0.9032833, -0.6274295, -0.3408952, 
    -0.04521877, 0.2827266, 0.5437686, 0.7892594,
  0.08603396, -0.01244956, -0.1302382, -0.230692, -0.3224648, -0.4244072, 
    -0.5279509, -0.5862728, -0.6336403, -0.6853408,
  -0.5083337, -0.6752201, -0.8401579, -1.021567, -1.198536, -1.330774, 
    -1.454516, -1.586487, -1.691136, -1.77504,
  -1.209975, -1.465892, -1.672402, -1.836556, -2.003343, -2.175733, 
    -2.340954, -2.462788, -2.570125, -2.671328,
  -1.835453, -2.040931, -2.250755, -2.488194, -2.693811, -2.848905, 
    -2.973454, -3.076011, -3.155657, -3.221975,
  -2.087997, -2.262499, -2.42809, -2.583258, -2.728339, -2.874663, -3.012026, 
    -3.105144, -3.219588, -3.292633,
  -2.219754, -2.239856, -2.291842, -2.338402, -2.416109, -2.477032, 
    -2.551712, -2.625169, -2.696625, -2.812562,
  -2.214184, -2.120897, -2.02604, -1.978979, -1.914884, -1.861667, -1.797479, 
    -1.808812, -1.854385, -1.959785,
  -2.145867, -1.937978, -1.761547, -1.585332, -1.406883, -1.215052, 
    -1.064301, -0.9400889, -0.883372, -0.8476374,
  -1.6123, -1.449645, -1.277987, -1.08922, -0.8639328, -0.5785105, 
    -0.3019016, -0.06757384, 0.1769251, 0.3469639,
  -0.4829444, -0.3573219, -0.2495783, -0.1331687, 0.03723535, 0.2394148, 
    0.4937723, 0.8273596, 1.081453, 1.332125,
  -0.8436456, -0.9486177, -1.059377, -1.153291, -1.241334, -1.344937, 
    -1.442711, -1.494026, -1.531425, -1.569082,
  -1.363601, -1.517111, -1.673566, -1.853703, -2.024385, -2.153884, 
    -2.277348, -2.399244, -2.49864, -2.581057,
  -1.900008, -2.121459, -2.298829, -2.446108, -2.600936, -2.75574, -2.91209, 
    -3.041326, -3.159974, -3.291958,
  -2.332246, -2.485257, -2.649413, -2.831298, -2.996419, -3.138222, 
    -3.260611, -3.390049, -3.512205, -3.606771,
  -2.484051, -2.582164, -2.656566, -2.747351, -2.843552, -2.953647, 
    -3.080211, -3.176885, -3.30392, -3.404524,
  -2.524805, -2.482363, -2.478343, -2.466771, -2.482541, -2.493074, 
    -2.524661, -2.568022, -2.622594, -2.706606,
  -2.361249, -2.253306, -2.134065, -2.054415, -1.964403, -1.889408, 
    -1.791761, -1.750293, -1.718029, -1.732389,
  -2.014955, -1.839144, -1.68769, -1.535044, -1.384408, -1.211162, -1.050033, 
    -0.8907735, -0.7928692, -0.7119153,
  -1.236629, -1.093662, -0.9508283, -0.8085872, -0.6442373, -0.4315634, 
    -0.1945382, -0.002699569, 0.1975364, 0.3391424,
  -0.113028, 0.03701114, 0.1509672, 0.244096, 0.3440107, 0.4850455, 0.659207, 
    0.8812482, 1.058411, 1.222257,
  -1.854996, -1.890166, -1.915619, -1.932104, -1.946811, -1.971547, 
    -1.988159, -1.97958, -1.964028, -1.948233,
  -2.224256, -2.271724, -2.324106, -2.393641, -2.449779, -2.481474, 
    -2.509733, -2.527462, -2.532758, -2.527077,
  -2.520393, -2.60658, -2.663467, -2.701849, -2.744738, -2.780796, -2.817967, 
    -2.841355, -2.859165, -2.87995,
  -2.696981, -2.736231, -2.781672, -2.833747, -2.878667, -2.9107, -2.931204, 
    -2.952544, -2.963497, -2.964039,
  -2.669573, -2.676523, -2.663651, -2.663748, -2.672803, -2.703568, -2.73891, 
    -2.744817, -2.765156, -2.767472,
  -2.476536, -2.429364, -2.405869, -2.377028, -2.36033, -2.332005, -2.306961, 
    -2.277795, -2.2701, -2.287573,
  -2.063781, -1.986485, -1.90999, -1.85632, -1.792651, -1.720523, -1.636689, 
    -1.607912, -1.594598, -1.61015,
  -1.519658, -1.429246, -1.343379, -1.238522, -1.116604, -1.015946, 
    -0.9358807, -0.8798366, -0.8500427, -0.8273263,
  -0.7674065, -0.6452081, -0.5515807, -0.4693587, -0.3846785, -0.3116637, 
    -0.2242767, -0.1593899, -0.1116388, -0.06896764,
  -0.01183324, 0.1091698, 0.2188423, 0.312474, 0.3854575, 0.4438081, 
    0.5140151, 0.5824342, 0.6187019, 0.6379458,
  -2.684902, -2.610719, -2.535948, -2.460751, -2.387049, -2.321111, 
    -2.254766, -2.182338, -2.107151, -2.031494,
  -2.820069, -2.740268, -2.659949, -2.584899, -2.516798, -2.444206, 
    -2.371544, -2.295798, -2.221301, -2.142587,
  -2.920424, -2.834318, -2.745224, -2.660668, -2.577662, -2.494831, -2.4213, 
    -2.345643, -2.268257, -2.192751,
  -2.919983, -2.838565, -2.757891, -2.677184, -2.599998, -2.519447, 
    -2.432564, -2.343707, -2.255901, -2.170567,
  -2.795936, -2.718457, -2.634572, -2.554108, -2.473378, -2.391261, 
    -2.312509, -2.233216, -2.158018, -2.077407,
  -2.562569, -2.481418, -2.403707, -2.320077, -2.236581, -2.159199, 
    -2.083839, -2.011575, -1.949767, -1.892647,
  -2.250703, -2.162687, -2.078802, -2.00374, -1.924842, -1.843397, -1.762613, 
    -1.697863, -1.633513, -1.583002,
  -1.825546, -1.773501, -1.720045, -1.646263, -1.569409, -1.491826, 
    -1.415384, -1.344221, -1.289576, -1.235646,
  -1.16891, -1.113447, -1.082653, -1.06613, -1.038724, -1.014261, -0.971841, 
    -0.9325086, -0.8841423, -0.8362257,
  -0.4466377, -0.3950162, -0.3640113, -0.3467484, -0.3497896, -0.3435763, 
    -0.3285452, -0.3093777, -0.3015329, -0.2992152,
  -3.47265, -3.349887, -3.225127, -3.099491, -2.975098, -2.858005, -2.742823, 
    -2.620348, -2.497191, -2.375009,
  -3.669024, -3.520918, -3.372771, -3.233594, -3.098513, -2.952549, 
    -2.805939, -2.665119, -2.521485, -2.376583,
  -3.875113, -3.713779, -3.561024, -3.408706, -3.2558, -3.100774, -2.95319, 
    -2.807744, -2.659667, -2.510706,
  -3.950386, -3.795719, -3.641412, -3.475792, -3.323338, -3.181724, 
    -3.039761, -2.904638, -2.775108, -2.650002,
  -3.947389, -3.783504, -3.606038, -3.452417, -3.30665, -3.171729, -3.049297, 
    -2.93359, -2.822966, -2.726708,
  -3.906445, -3.746139, -3.594896, -3.442577, -3.297046, -3.1648, -3.036906, 
    -2.916452, -2.812173, -2.712864,
  -3.83857, -3.71836, -3.602963, -3.481781, -3.346611, -3.205612, -3.061509, 
    -2.923938, -2.794568, -2.691266,
  -3.559861, -3.530004, -3.478284, -3.396861, -3.302307, -3.188716, 
    -3.069149, -2.94336, -2.817003, -2.663864,
  -2.915129, -2.919575, -2.929287, -2.93514, -2.908199, -2.866826, -2.797559, 
    -2.709057, -2.578434, -2.428774,
  -2.010599, -2.042224, -2.077676, -2.104624, -2.122853, -2.120454, 
    -2.097497, -2.047853, -1.992431, -1.92157,
  -4.22112, -4.07559, -3.922843, -3.768222, -3.614719, -3.473573, -3.340809, 
    -3.200793, -3.061464, -2.926893,
  -4.502892, -4.344226, -4.183433, -4.026276, -3.878217, -3.729609, -3.58069, 
    -3.431968, -3.287462, -3.145941,
  -4.631217, -4.473382, -4.315218, -4.164486, -4.013389, -3.85793, -3.710944, 
    -3.570176, -3.429156, -3.28708,
  -4.626989, -4.476557, -4.326241, -4.174338, -4.032887, -3.895635, 
    -3.756263, -3.619544, -3.485802, -3.356973,
  -4.556738, -4.395508, -4.235921, -4.096162, -3.958964, -3.832275, 
    -3.715655, -3.600988, -3.489401, -3.387974,
  -4.468916, -4.302645, -4.15163, -4.001896, -3.865624, -3.743882, -3.626797, 
    -3.521506, -3.429111, -3.338457,
  -4.44977, -4.292527, -4.144361, -4.001679, -3.853956, -3.707088, -3.567008, 
    -3.438192, -3.317925, -3.220261,
  -4.439157, -4.329401, -4.202333, -4.056956, -3.905393, -3.736642, 
    -3.568599, -3.403389, -3.260043, -3.114572,
  -4.203069, -4.12499, -4.031964, -3.926179, -3.793952, -3.63649, -3.470912, 
    -3.312045, -3.139288, -2.968029,
  -3.549062, -3.518938, -3.466148, -3.407319, -3.308811, -3.204609, 
    -3.090285, -2.963688, -2.832902, -2.702063,
  -4.634931, -4.510322, -4.387384, -4.262967, -4.13814, -4.019274, -3.907151, 
    -3.793168, -3.677498, -3.562162,
  -4.812496, -4.685526, -4.557202, -4.432652, -4.315062, -4.196854, 
    -4.077685, -3.961596, -3.849445, -3.737238,
  -4.926235, -4.801914, -4.682349, -4.564368, -4.445381, -4.328474, 
    -4.217326, -4.105275, -3.991226, -3.87654,
  -4.974308, -4.86126, -4.746056, -4.629657, -4.521437, -4.412365, -4.300677, 
    -4.186651, -4.075935, -3.968378,
  -4.938999, -4.831478, -4.722439, -4.619403, -4.516479, -4.414182, 
    -4.313823, -4.215149, -4.114635, -4.01406,
  -4.802555, -4.709178, -4.621257, -4.533046, -4.446228, -4.362994, 
    -4.278905, -4.198927, -4.114691, -4.029364,
  -4.646967, -4.549815, -4.467683, -4.393793, -4.318109, -4.249639, 
    -4.184724, -4.118573, -4.056467, -3.996501,
  -4.553621, -4.461698, -4.370646, -4.279413, -4.197869, -4.108099, 
    -4.025449, -3.951957, -3.882595, -3.806807,
  -4.450593, -4.350024, -4.254059, -4.160119, -4.047391, -3.930037, 
    -3.814608, -3.705483, -3.598191, -3.498837,
  -4.176404, -4.088185, -3.99167, -3.888712, -3.763858, -3.636919, -3.503574, 
    -3.371032, -3.253147, -3.15005,
  -5.305916, -5.228198, -5.149081, -5.066242, -4.979733, -4.891483, 
    -4.805131, -4.715399, -4.625538, -4.536609,
  -5.409827, -5.338651, -5.264568, -5.190886, -5.118539, -5.040178, 
    -4.958767, -4.879787, -4.798156, -4.714354,
  -5.436405, -5.377537, -5.321352, -5.260819, -5.19785, -5.135309, -5.069129, 
    -4.99902, -4.925947, -4.848398,
  -5.425586, -5.371675, -5.315626, -5.258965, -5.205391, -5.147702, 
    -5.090356, -5.029489, -4.966897, -4.903516,
  -5.421552, -5.364684, -5.306411, -5.247279, -5.189979, -5.13738, -5.082496, 
    -5.023454, -4.961823, -4.898187,
  -5.399646, -5.353481, -5.305019, -5.255711, -5.203397, -5.146911, 
    -5.086962, -5.023842, -4.958927, -4.891607,
  -5.324206, -5.285987, -5.253324, -5.216431, -5.17214, -5.119621, -5.066675, 
    -5.011673, -4.952978, -4.889044,
  -5.201594, -5.185238, -5.161349, -5.129875, -5.091774, -5.047886, 
    -5.002157, -4.954802, -4.903096, -4.845263,
  -5.027672, -5.009829, -4.996872, -4.982873, -4.957479, -4.928816, 
    -4.894786, -4.855186, -4.809749, -4.755376,
  -4.800905, -4.790343, -4.778637, -4.76788, -4.754467, -4.730603, -4.70276, 
    -4.672376, -4.637187, -4.600635,
  -5.877733, -5.806942, -5.737911, -5.665781, -5.589697, -5.508978, 
    -5.428902, -5.346344, -5.262498, -5.177478,
  -5.999748, -5.93775, -5.871769, -5.80268, -5.736236, -5.664495, -5.589656, 
    -5.515277, -5.436458, -5.355067,
  -6.105768, -6.050148, -5.99489, -5.934047, -5.869964, -5.807178, -5.740132, 
    -5.669778, -5.59723, -5.518231,
  -6.204219, -6.156556, -6.104576, -6.049919, -5.996562, -5.93629, -5.873829, 
    -5.805651, -5.734739, -5.662208,
  -6.283307, -6.238613, -6.188774, -6.136417, -6.083857, -6.031115, 
    -5.974864, -5.914575, -5.849953, -5.782243,
  -6.327734, -6.29085, -6.250577, -6.207967, -6.160203, -6.109562, -6.055408, 
    -5.996362, -5.935081, -5.871264,
  -6.328987, -6.301887, -6.276907, -6.244695, -6.205217, -6.156336, 
    -6.106204, -6.054013, -5.999475, -5.941885,
  -6.286625, -6.282731, -6.267518, -6.242774, -6.20835, -6.168219, -6.125497, 
    -6.080946, -6.031807, -5.975547,
  -6.193247, -6.187342, -6.183197, -6.175198, -6.155711, -6.131026, -6.09807, 
    -6.059319, -6.013174, -5.959172,
  -6.058994, -6.055746, -6.05086, -6.046446, -6.038727, -6.018096, -5.98981, 
    -5.954857, -5.918507, -5.881165,
  -6.561323, -6.499266, -6.438377, -6.375708, -6.310773, -6.244139, 
    -6.180099, -6.115896, -6.051152, -5.986147,
  -6.845045, -6.786884, -6.725439, -6.661109, -6.601454, -6.540991, 
    -6.479097, -6.417562, -6.355603, -6.293946,
  -7.102453, -7.045627, -6.989235, -6.932842, -6.874574, -6.816972, 
    -6.758873, -6.701811, -6.644189, -6.583754,
  -7.351357, -7.301179, -7.248499, -7.19398, -7.142448, -7.089523, -7.035904, 
    -6.981055, -6.926404, -6.871471,
  -7.598204, -7.549111, -7.497645, -7.447221, -7.397934, -7.350796, 
    -7.304009, -7.256029, -7.20568, -7.155462,
  -7.82113, -7.78062, -7.739799, -7.69751, -7.652907, -7.609156, -7.56383, 
    -7.517503, -7.472572, -7.428266,
  -8.020307, -7.985536, -7.955499, -7.923059, -7.885509, -7.841635, 
    -7.801394, -7.76416, -7.727195, -7.691062,
  -8.203031, -8.185472, -8.161825, -8.130711, -8.093474, -8.056222, 
    -8.020072, -7.988377, -7.958443, -7.925798,
  -8.343966, -8.324842, -8.308795, -8.291328, -8.267859, -8.240988, -8.21365, 
    -8.186219, -8.156057, -8.126547,
  -8.44836, -8.431485, -8.415438, -8.404657, -8.391961, -8.373449, -8.350844, 
    -8.326425, -8.308137, -8.293455,
  -7.418903, -7.380289, -7.343199, -7.30528, -7.266068, -7.225653, -7.186882, 
    -7.148771, -7.1104, -7.071782,
  -7.886793, -7.851552, -7.814201, -7.774897, -7.739104, -7.703277, 
    -7.666594, -7.630272, -7.594023, -7.558314,
  -8.341415, -8.308264, -8.274553, -8.240778, -8.205718, -8.171395, 
    -8.137189, -8.103981, -8.07057, -8.035443,
  -8.796901, -8.767877, -8.73701, -8.704835, -8.674766, -8.644069, -8.61279, 
    -8.580782, -8.54905, -8.517601,
  -9.253543, -9.225341, -9.195226, -9.165483, -9.137247, -9.111868, 
    -9.086359, -9.059315, -9.030994, -9.003092,
  -9.699064, -9.677286, -9.654745, -9.63162, -9.607246, -9.582701, -9.557117, 
    -9.531214, -9.505648, -9.481256,
  -10.12736, -10.10717, -10.09253, -10.07685, -10.05586, -10.03019, 
    -10.00788, -9.988334, -9.96856, -9.949014,
  -10.53594, -10.52901, -10.51833, -10.50091, -10.47864, -10.45729, 
    -10.43758, -10.42123, -10.40631, -10.38915,
  -10.90329, -10.89263, -10.88709, -10.88161, -10.87157, -10.86071, 
    -10.84752, -10.83391, -10.81815, -10.80181,
  -11.248, -11.23781, -11.23062, -11.22926, -11.23034, -11.22393, -11.21365, 
    -11.20186, -11.19413, -11.18977,
  -13.83239, -13.82074, -13.808, -13.79507, -13.78222, -13.76985, -13.75674, 
    -13.74387, -13.73124, -13.71895,
  -14.99369, -14.98229, -14.97097, -14.96008, -14.94822, -14.9366, -14.92516, 
    -14.9145, -14.90532, -14.89437,
  -16.12242, -16.11533, -16.10389, -16.09248, -16.08173, -16.06978, 
    -16.06084, -16.05067, -16.03975, -16.03102,
  -17.2117, -17.20174, -17.1923, -17.18274, -17.17234, -17.16337, -17.15279, 
    -17.14514, -17.13551, -17.12395,
  -18.23167, -18.22563, -18.21396, -18.20369, -18.19536, -18.19025, -18.1865, 
    -18.17599, -18.1694, -18.16037,
  -19.16084, -19.15458, -19.15068, -19.14543, -19.14352, -19.13608, 
    -19.12984, -19.12499, -19.11406, -19.10741,
  -19.96635, -19.96284, -19.96158, -19.96541, -19.9607, -19.95777, -19.95134, 
    -19.94964, -19.94552, -19.9427,
  -20.64782, -20.64862, -20.65172, -20.64795, -20.64328, -20.63709, -20.6386, 
    -20.63893, -20.64199, -20.63851,
  -21.1739, -21.17439, -21.17778, -21.18302, -21.18665, -21.19431, -21.1958, 
    -21.1981, -21.19873, -21.19386,
  -21.59861, -21.59514, -21.59659, -21.60578, -21.61945, -21.62407, 
    -21.62483, -21.62446, -21.6267, -21.63452 ;
}
