netcdf \00010101.ocean_static {
dimensions:
	yq = 10 ;
	xq = 15 ;
	yh = 10 ;
	xh = 15 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float Coriolis(yq, xq) ;
		Coriolis:_FillValue = 1.e+20f ;
		Coriolis:missing_value = 1.e+20f ;
		Coriolis:units = "s-1" ;
		Coriolis:long_name = "Coriolis parameter at corner (Bu) points" ;
		Coriolis:cell_methods = "time: point" ;
		Coriolis:interp_method = "none" ;
	float areacello(yh, xh) ;
		areacello:_FillValue = 1.e+20f ;
		areacello:missing_value = 1.e+20f ;
		areacello:units = "m2" ;
		areacello:long_name = "Ocean Grid-Cell Area" ;
		areacello:cell_methods = "area:sum yh:sum xh:sum time: point" ;
		areacello:standard_name = "cell_area" ;
	float areacello_bu(yq, xq) ;
		areacello_bu:_FillValue = 1.e+20f ;
		areacello_bu:missing_value = 1.e+20f ;
		areacello_bu:units = "m2" ;
		areacello_bu:long_name = "Ocean Grid-Cell Area" ;
		areacello_bu:cell_methods = "area:sum yq:sum xq:sum time: point" ;
		areacello_bu:standard_name = "cell_area" ;
	float areacello_cu(yh, xq) ;
		areacello_cu:_FillValue = 1.e+20f ;
		areacello_cu:missing_value = 1.e+20f ;
		areacello_cu:units = "m2" ;
		areacello_cu:long_name = "Ocean Grid-Cell Area" ;
		areacello_cu:cell_methods = "area:sum yh:sum xq:sum time: point" ;
		areacello_cu:standard_name = "cell_area" ;
	float areacello_cv(yq, xh) ;
		areacello_cv:_FillValue = 1.e+20f ;
		areacello_cv:missing_value = 1.e+20f ;
		areacello_cv:units = "m2" ;
		areacello_cv:long_name = "Ocean Grid-Cell Area" ;
		areacello_cv:cell_methods = "area:sum yq:sum xh:sum time: point" ;
		areacello_cv:standard_name = "cell_area" ;
	float deptho(yh, xh) ;
		deptho:_FillValue = 1.e+20f ;
		deptho:missing_value = 1.e+20f ;
		deptho:units = "m" ;
		deptho:long_name = "Sea Floor Depth" ;
		deptho:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		deptho:cell_measures = "area: areacello" ;
		deptho:standard_name = "sea_floor_depth_below_geoid" ;
	float dxCu(yh, xq) ;
		dxCu:_FillValue = 1.e+20f ;
		dxCu:missing_value = 1.e+20f ;
		dxCu:units = "m" ;
		dxCu:long_name = "Delta(x) at u points (meter)" ;
		dxCu:cell_methods = "time: point" ;
		dxCu:interp_method = "none" ;
	float dxCv(yq, xh) ;
		dxCv:_FillValue = 1.e+20f ;
		dxCv:missing_value = 1.e+20f ;
		dxCv:units = "m" ;
		dxCv:long_name = "Delta(x) at v points (meter)" ;
		dxCv:cell_methods = "time: point" ;
		dxCv:interp_method = "none" ;
	float dxt(yh, xh) ;
		dxt:_FillValue = 1.e+20f ;
		dxt:missing_value = 1.e+20f ;
		dxt:units = "m" ;
		dxt:long_name = "Delta(x) at thickness/tracer points (meter)" ;
		dxt:cell_methods = "time: point" ;
		dxt:interp_method = "none" ;
	float dyCu(yh, xq) ;
		dyCu:_FillValue = 1.e+20f ;
		dyCu:missing_value = 1.e+20f ;
		dyCu:units = "m" ;
		dyCu:long_name = "Delta(y) at u points (meter)" ;
		dyCu:cell_methods = "time: point" ;
		dyCu:interp_method = "none" ;
	float dyCv(yq, xh) ;
		dyCv:_FillValue = 1.e+20f ;
		dyCv:missing_value = 1.e+20f ;
		dyCv:units = "m" ;
		dyCv:long_name = "Delta(y) at v points (meter)" ;
		dyCv:cell_methods = "time: point" ;
		dyCv:interp_method = "none" ;
	float dyt(yh, xh) ;
		dyt:_FillValue = 1.e+20f ;
		dyt:missing_value = 1.e+20f ;
		dyt:units = "m" ;
		dyt:long_name = "Delta(y) at thickness/tracer points (meter)" ;
		dyt:cell_methods = "time: point" ;
		dyt:interp_method = "none" ;
	float geolat(yh, xh) ;
		geolat:_FillValue = 1.e+20f ;
		geolat:missing_value = 1.e+20f ;
		geolat:units = "degrees_north" ;
		geolat:long_name = "Latitude of tracer (T) points" ;
		geolat:cell_methods = "time: point" ;
	float geolat_c(yq, xq) ;
		geolat_c:_FillValue = 1.e+20f ;
		geolat_c:missing_value = 1.e+20f ;
		geolat_c:units = "degrees_north" ;
		geolat_c:long_name = "Latitude of corner (Bu) points" ;
		geolat_c:cell_methods = "time: point" ;
		geolat_c:interp_method = "none" ;
	float geolat_u(yh, xq) ;
		geolat_u:_FillValue = 1.e+20f ;
		geolat_u:missing_value = 1.e+20f ;
		geolat_u:units = "degrees_north" ;
		geolat_u:long_name = "Latitude of zonal velocity (Cu) points" ;
		geolat_u:cell_methods = "time: point" ;
		geolat_u:interp_method = "none" ;
	float geolat_v(yq, xh) ;
		geolat_v:_FillValue = 1.e+20f ;
		geolat_v:missing_value = 1.e+20f ;
		geolat_v:units = "degrees_north" ;
		geolat_v:long_name = "Latitude of meridional velocity (Cv) points" ;
		geolat_v:cell_methods = "time: point" ;
		geolat_v:interp_method = "none" ;
	float geolon(yh, xh) ;
		geolon:_FillValue = 1.e+20f ;
		geolon:missing_value = 1.e+20f ;
		geolon:units = "degrees_east" ;
		geolon:long_name = "Longitude of tracer (T) points" ;
		geolon:cell_methods = "time: point" ;
	float geolon_c(yq, xq) ;
		geolon_c:_FillValue = 1.e+20f ;
		geolon_c:missing_value = 1.e+20f ;
		geolon_c:units = "degrees_east" ;
		geolon_c:long_name = "Longitude of corner (Bu) points" ;
		geolon_c:cell_methods = "time: point" ;
		geolon_c:interp_method = "none" ;
	float geolon_u(yh, xq) ;
		geolon_u:_FillValue = 1.e+20f ;
		geolon_u:missing_value = 1.e+20f ;
		geolon_u:units = "degrees_east" ;
		geolon_u:long_name = "Longitude of zonal velocity (Cu) points" ;
		geolon_u:cell_methods = "time: point" ;
		geolon_u:interp_method = "none" ;
	float geolon_v(yq, xh) ;
		geolon_v:_FillValue = 1.e+20f ;
		geolon_v:missing_value = 1.e+20f ;
		geolon_v:units = "degrees_east" ;
		geolon_v:long_name = "Longitude of meridional velocity (Cv) points" ;
		geolon_v:cell_methods = "time: point" ;
		geolon_v:interp_method = "none" ;
	float hfgeou(yh, xh) ;
		hfgeou:_FillValue = 1.e+20f ;
		hfgeou:missing_value = 1.e+20f ;
		hfgeou:units = "W m-2" ;
		hfgeou:long_name = "Upward geothermal heat flux at sea floor" ;
		hfgeou:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		hfgeou:standard_name = "upward_geothermal_heat_flux_at_sea_floor" ;
	float sftof(yh, xh) ;
		sftof:_FillValue = 1.e+20f ;
		sftof:missing_value = 1.e+20f ;
		sftof:units = "%" ;
		sftof:long_name = "Sea Area Fraction" ;
		sftof:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		sftof:standard_name = "SeaAreaFraction" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
	float wet(yh, xh) ;
		wet:_FillValue = 1.e+20f ;
		wet:missing_value = 1.e+20f ;
		wet:long_name = "0 if land, 1 if ocean at tracer points" ;
		wet:cell_methods = "time: point" ;
		wet:cell_measures = "area: areacello" ;
	float wet_c(yq, xq) ;
		wet_c:_FillValue = 1.e+20f ;
		wet_c:missing_value = 1.e+20f ;
		wet_c:long_name = "0 if land, 1 if ocean at corner (Bu) points" ;
		wet_c:cell_methods = "time: point" ;
		wet_c:interp_method = "none" ;
	float wet_u(yh, xq) ;
		wet_u:_FillValue = 1.e+20f ;
		wet_u:missing_value = 1.e+20f ;
		wet_u:long_name = "0 if land, 1 if ocean at zonal velocity (Cu) points" ;
		wet_u:cell_methods = "time: point" ;
		wet_u:interp_method = "none" ;
	float wet_v(yq, xh) ;
		wet_v:_FillValue = 1.e+20f ;
		wet_v:missing_value = 1.e+20f ;
		wet_v:long_name = "0 if land, 1 if ocean at meridional velocity (Cv) points" ;
		wet_v:cell_methods = "time: point" ;
		wet_v:interp_method = "none" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Jun 13 14:06:58 2025: ncks -d xh,532,546 -d yh,526,535 -d xq,532,546 -d yq,526,535 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.ocean_static.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.ocean_static.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 Coriolis =
  -3.643884e-05, -3.643884e-05, -3.643884e-05, -3.643884e-05, -3.643884e-05, 
    -3.643884e-05, -3.643884e-05, -3.643884e-05, -3.643884e-05, 
    -3.643884e-05, -3.643884e-05, -3.643884e-05, -3.643884e-05, 
    -3.643884e-05, -3.643884e-05,
  -3.584156e-05, -3.584156e-05, -3.584156e-05, -3.584156e-05, -3.584156e-05, 
    -3.584156e-05, -3.584156e-05, -3.584156e-05, -3.584156e-05, 
    -3.584156e-05, -3.584156e-05, -3.584156e-05, -3.584156e-05, 
    -3.584156e-05, -3.584156e-05,
  -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05, 
    -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05, 
    -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05, -3.5243e-05,
  -3.464318e-05, -3.464318e-05, -3.464318e-05, -3.464318e-05, -3.464318e-05, 
    -3.464318e-05, -3.464318e-05, -3.464318e-05, -3.464318e-05, 
    -3.464318e-05, -3.464318e-05, -3.464318e-05, -3.464318e-05, 
    -3.464318e-05, -3.464318e-05,
  -3.404211e-05, -3.404211e-05, -3.404211e-05, -3.404211e-05, -3.404211e-05, 
    -3.404211e-05, -3.404211e-05, -3.404211e-05, -3.404211e-05, 
    -3.404211e-05, -3.404211e-05, -3.404211e-05, -3.404211e-05, 
    -3.404211e-05, -3.404211e-05,
  -3.343981e-05, -3.343981e-05, -3.343981e-05, -3.343981e-05, -3.343981e-05, 
    -3.343981e-05, -3.343981e-05, -3.343981e-05, -3.343981e-05, 
    -3.343981e-05, -3.343981e-05, -3.343981e-05, -3.343981e-05, 
    -3.343981e-05, -3.343981e-05,
  -3.283631e-05, -3.283631e-05, -3.283631e-05, -3.283631e-05, -3.283631e-05, 
    -3.283631e-05, -3.283631e-05, -3.283631e-05, -3.283631e-05, 
    -3.283631e-05, -3.283631e-05, -3.283631e-05, -3.283631e-05, 
    -3.283631e-05, -3.283631e-05,
  -3.223163e-05, -3.223163e-05, -3.223163e-05, -3.223163e-05, -3.223163e-05, 
    -3.223163e-05, -3.223163e-05, -3.223163e-05, -3.223163e-05, 
    -3.223163e-05, -3.223163e-05, -3.223163e-05, -3.223163e-05, 
    -3.223163e-05, -3.223163e-05,
  -3.162577e-05, -3.162577e-05, -3.162577e-05, -3.162577e-05, -3.162577e-05, 
    -3.162577e-05, -3.162577e-05, -3.162577e-05, -3.162577e-05, 
    -3.162577e-05, -3.162577e-05, -3.162577e-05, -3.162577e-05, 
    -3.162577e-05, -3.162577e-05,
  -3.101877e-05, -3.101877e-05, -3.101877e-05, -3.101877e-05, -3.101877e-05, 
    -3.101877e-05, -3.101877e-05, -3.101877e-05, -3.101877e-05, 
    -3.101877e-05, -3.101877e-05, -3.101877e-05, -3.101877e-05, 
    -3.101877e-05, -3.101877e-05 ;

 areacello =
  7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08, 
    7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08, 
    7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08, 7.253149e+08,
  7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08, 
    7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08, 
    7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08, 7.268721e+08,
  7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08, 
    7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08, 
    7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08, 7.284065e+08,
  7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08, 
    7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08, 
    7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08, 7.29918e+08,
  7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08, 
    7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08, 
    7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08, 7.314063e+08,
  7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08, 
    7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08, 
    7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08, 7.328712e+08,
  7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08, 
    7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08, 
    7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08, 7.343126e+08,
  7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08, 
    7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08, 
    7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08, 7.357302e+08,
  7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08, 
    7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08, 
    7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08, 7.371238e+08,
  7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08, 
    7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08, 
    7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08, 7.384932e+08 ;

 areacello_bu =
  7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08, 
    7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08, 
    7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08, 7.245278e+08,
  7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08, 
    7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08, 
    7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08, 7.260963e+08,
  7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08, 
    7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08, 
    7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08, 7.276422e+08,
  7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08, 
    7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08, 
    7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08, 7.291651e+08,
  7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08, 
    7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08, 
    7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08, 7.306651e+08,
  7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08, 
    7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08, 
    7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08, 7.321417e+08,
  7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08, 
    7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08, 
    7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08, 7.335949e+08,
  7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08, 
    7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08, 
    7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08, 7.350244e+08,
  7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 
    7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 7.3643e+08, 
    7.3643e+08, 7.3643e+08, 7.3643e+08,
  7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08, 
    7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08, 
    7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08, 7.378115e+08 ;

 areacello_cu =
  7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08, 
    7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08, 
    7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08, 7.253153e+08,
  7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08, 
    7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08, 
    7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08, 7.268725e+08,
  7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08, 
    7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08, 
    7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08, 7.28407e+08,
  7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08, 
    7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08, 
    7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08, 7.299185e+08,
  7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08, 
    7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08, 
    7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08, 7.314068e+08,
  7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08, 
    7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08, 
    7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08, 7.328717e+08,
  7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08, 
    7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08, 
    7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08, 7.343131e+08,
  7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08, 
    7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08, 
    7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08, 7.357306e+08,
  7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08, 
    7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08, 
    7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08, 7.371242e+08,
  7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08, 
    7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08, 
    7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08, 7.384936e+08 ;

 areacello_cv =
  7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08, 
    7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08, 
    7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08, 7.245283e+08,
  7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08, 
    7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08, 
    7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08, 7.260968e+08,
  7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08, 
    7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08, 
    7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08, 7.276426e+08,
  7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08, 
    7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08, 
    7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08, 7.291656e+08,
  7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08, 
    7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08, 
    7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08, 7.306655e+08,
  7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08, 
    7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08, 
    7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08, 7.321421e+08,
  7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08, 
    7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08, 
    7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08, 7.335953e+08,
  7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08, 
    7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08, 
    7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08, 7.350248e+08,
  7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08, 
    7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08, 
    7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08, 7.364305e+08,
  7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08, 
    7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08, 
    7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08, 7.37812e+08 ;

 deptho =
  5459.581, 5518.351, 5471.555, 5464.517, 5493.351, 5443.992, 5481.438, 
    5399.232, 5437.585, 5564.116, 5508.024, 5278.302, 5339.634, 5338.516, 
    5362.45,
  5444.997, 5526.517, 5558.977, 5506.794, 5539.163, 5464.714, 5371.029, 
    5283.403, 5344.632, 5276.831, 5453.903, 5460.983, 5401.993, 5373.839, 
    5222.505,
  5469.43, 5485.55, 5484.331, 5534.783, 5515.036, 5381.512, 5379.43, 
    5436.272, 5353.861, 5308.952, 5356.044, 5565.796, 5455.912, 5291.331, 
    5030.697,
  5377.339, 5432.107, 5414.18, 5474.686, 5430.449, 5403.279, 5411.458, 
    5495.017, 5410.293, 5379.038, 5393.203, 5604.945, 5393.119, 4742.138, 
    4438.138,
  5412.795, 5426.14, 5400.57, 5435.193, 5439.468, 5473.852, 5430.786, 
    5391.758, 5547.167, 5492.971, 5509.514, 5286.06, 4352.004, 4455.662, 
    3532.009,
  5441.89, 5533.067, 5532.043, 5451.808, 5465.8, 5563.95, 5503.784, 5289.503, 
    5447.585, 5495.046, 5438.338, 5136.738, 4889.081, 4330.568, 3322.158,
  5367.564, 5623.584, 5646.252, 5546.898, 5537.195, 5522.411, 4901.873, 
    5396.403, 5512.202, 5424.177, 5183.489, 5008.471, 5015.458, 3874.39, 
    3237.326,
  5536.536, 5390.403, 5186.029, 5572.206, 5660.611, 5683.173, 5679.197, 
    5480.841, 5338.633, 5219.022, 5189.761, 4972.972, 4596.265, 3853.92, 3078,
  5527.949, 5094.13, 4281.74, 5565.208, 5684.5, 5743.412, 5613.496, 5286.793, 
    5167.222, 5019.19, 4948.869, 4768.419, 4239.951, 3896.296, 3292.449,
  5542.585, 5490.353, 5468.412, 5531.694, 5649.889, 5580.06, 5496.899, 
    4881.083, 4591.047, 4642.272, 4266.763, 3973.73, 3807.69, 3853.071, 
    3504.758 ;

 dxCu =
  26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 
    26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 
    26931.69,
  26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 
    26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 
    26960.58,
  26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 
    26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 
    26989.03,
  27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 
    27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 
    27017.01,
  27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 
    27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 
    27044.54,
  27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 
    27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 
    27071.61,
  27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 
    27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 
    27098.22,
  27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 
    27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 
    27124.37,
  27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 
    27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 
    27150.04,
  27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 
    27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 
    27175.25 ;

 dxCv =
  26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 
    26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 26917.07, 
    26917.07,
  26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 
    26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 26946.19, 
    26946.19,
  26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 
    26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 26974.86, 
    26974.86,
  27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 
    27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 27003.08, 
    27003.08,
  27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 
    27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 27030.83, 
    27030.83,
  27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 
    27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 27058.13, 
    27058.13,
  27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 
    27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 27084.97, 
    27084.97,
  27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 
    27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 27111.35, 
    27111.35,
  27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 
    27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 27137.26, 
    27137.26,
  27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 
    27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 27162.71, 
    27162.71 ;

 dxt =
  26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 
    26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 26931.69, 
    26931.69,
  26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 
    26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 26960.58, 
    26960.58,
  26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 
    26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 26989.03, 
    26989.03,
  27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 
    27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 27017.01, 
    27017.01,
  27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 
    27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 27044.54, 
    27044.54,
  27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 
    27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 27071.61, 
    27071.61,
  27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 
    27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 27098.22, 
    27098.22,
  27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 
    27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 27124.37, 
    27124.37,
  27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 
    27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 27150.04, 
    27150.04,
  27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 
    27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 27175.25, 
    27175.25 ;

 dyCu =
  26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 
    26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 
    26931.67,
  26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 
    26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 
    26960.56,
  26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 
    26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 
    26989.01,
  27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 
    27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 
    27016.99,
  27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 
    27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 
    27044.52,
  27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 
    27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 
    27071.59,
  27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 
    27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2,
  27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 
    27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 
    27124.35,
  27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 
    27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 
    27150.02,
  27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 
    27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 
    27175.23 ;

 dyCv =
  26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 
    26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 26917.05, 
    26917.05,
  26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 
    26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 26946.17, 
    26946.17,
  26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 
    26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 26974.84, 
    26974.84,
  27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 
    27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 27003.06, 
    27003.06,
  27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 
    27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 27030.82, 
    27030.82,
  27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 
    27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 27058.12, 
    27058.12,
  27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 
    27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 27084.96, 
    27084.96,
  27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 
    27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 27111.33, 
    27111.33,
  27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 
    27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 27137.24, 
    27137.24,
  27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 
    27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 27162.69, 
    27162.69 ;

 dyt =
  26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 
    26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 26931.67, 
    26931.67,
  26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 
    26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 26960.56, 
    26960.56,
  26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 
    26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 26989.01, 
    26989.01,
  27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 
    27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 27016.99, 
    27016.99,
  27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 
    27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 27044.52, 
    27044.52,
  27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 
    27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 27071.59, 
    27071.59,
  27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 
    27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2, 27098.2,
  27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 
    27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 27124.35, 
    27124.35,
  27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 
    27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 27150.02, 
    27150.02,
  27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 
    27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 27175.23, 
    27175.23 ;

 geolat =
  -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, 
    -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, 
    -14.34766, -14.34766, -14.34766,
  -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, 
    -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, 
    -14.10532, -14.10532, -14.10532,
  -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, 
    -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, 
    -13.86273, -13.86273, -13.86273,
  -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, 
    -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, 
    -13.61989, -13.61989, -13.61989,
  -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, 
    -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, 
    -13.37679, -13.37679, -13.37679,
  -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, 
    -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, 
    -13.13345, -13.13345, -13.13345,
  -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, 
    -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, 
    -12.88987, -12.88987, -12.88987,
  -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, 
    -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, 
    -12.64606, -12.64606, -12.64606,
  -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, 
    -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402,
  -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, 
    -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, 
    -12.15772, -12.15772, -12.15772 ;

 geolat_c =
  -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, 
    -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, 
    -14.46872, -14.46872, -14.46872,
  -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, 
    -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, 
    -14.22652, -14.22652, -14.22652,
  -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, 
    -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, 
    -13.98406, -13.98406, -13.98406,
  -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, 
    -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, 
    -13.74134, -13.74134, -13.74134,
  -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, 
    -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, 
    -13.49837, -13.49837, -13.49837,
  -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, 
    -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, 
    -13.25515, -13.25515, -13.25515,
  -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, 
    -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, 
    -13.01169, -13.01169, -13.01169,
  -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, 
    -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, 
    -12.76799, -12.76799, -12.76799,
  -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, 
    -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, 
    -12.52406, -12.52406, -12.52406,
  -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, 
    -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, 
    -12.27989, -12.27989, -12.27989 ;

 geolat_u =
  -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, 
    -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, -14.34766, 
    -14.34766, -14.34766, -14.34766,
  -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, 
    -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, -14.10532, 
    -14.10532, -14.10532, -14.10532,
  -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, 
    -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, -13.86273, 
    -13.86273, -13.86273, -13.86273,
  -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, 
    -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, -13.61989, 
    -13.61989, -13.61989, -13.61989,
  -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, 
    -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, -13.37679, 
    -13.37679, -13.37679, -13.37679,
  -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, 
    -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, -13.13345, 
    -13.13345, -13.13345, -13.13345,
  -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, 
    -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, -12.88987, 
    -12.88987, -12.88987, -12.88987,
  -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, 
    -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, -12.64606, 
    -12.64606, -12.64606, -12.64606,
  -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, 
    -12.402, -12.402, -12.402, -12.402, -12.402, -12.402, -12.402,
  -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, 
    -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, -12.15772, 
    -12.15772, -12.15772, -12.15772 ;

 geolat_v =
  -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, 
    -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, -14.46872, 
    -14.46872, -14.46872, -14.46872,
  -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, 
    -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, -14.22652, 
    -14.22652, -14.22652, -14.22652,
  -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, 
    -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, -13.98406, 
    -13.98406, -13.98406, -13.98406,
  -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, 
    -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, -13.74134, 
    -13.74134, -13.74134, -13.74134,
  -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, 
    -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, -13.49837, 
    -13.49837, -13.49837, -13.49837,
  -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, 
    -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, -13.25515, 
    -13.25515, -13.25515, -13.25515,
  -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, 
    -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, -13.01169, 
    -13.01169, -13.01169, -13.01169,
  -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, 
    -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, -12.76799, 
    -12.76799, -12.76799, -12.76799,
  -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, 
    -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, -12.52406, 
    -12.52406, -12.52406, -12.52406,
  -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, 
    -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, -12.27989, 
    -12.27989, -12.27989, -12.27989 ;

 geolon =
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 geolon_c =
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 geolon_u =
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5,
  -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 geolon_v =
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375,
  -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 hfgeou =
  0.07096534, 0.07089603, 0.07082672, 0.0707574, 0.07068809, 0.07061878, 
    0.07054947, 0.07048015, 0.07044549, 0.07044549, 0.07044549, 0.07044549, 
    0.07044549, 0.07044549, 0.07044549,
  0.07095248, 0.07085741, 0.07076235, 0.07066729, 0.07057223, 0.07047717, 
    0.0703821, 0.07028704, 0.07023951, 0.07023951, 0.07023951, 0.07023951, 
    0.07023951, 0.07023951, 0.07023951,
  0.07093959, 0.07081874, 0.07069791, 0.07057708, 0.07045624, 0.0703354, 
    0.07021457, 0.07009373, 0.07003331, 0.07003331, 0.07003331, 0.07003331, 
    0.07003331, 0.07003331, 0.07003331,
  0.07092668, 0.07078005, 0.0706334, 0.07048677, 0.07034013, 0.07019349, 
    0.07004685, 0.06990021, 0.06982689, 0.06982689, 0.06982689, 0.06982689, 
    0.06982689, 0.06982689, 0.06982689,
  0.07091377, 0.0707413, 0.07056884, 0.07039636, 0.0702239, 0.07005143, 
    0.06987897, 0.0697065, 0.06962027, 0.06962027, 0.06962027, 0.06962027, 
    0.06962027, 0.06962027, 0.06962027,
  0.07090084, 0.07070252, 0.0705042, 0.07030588, 0.07010756, 0.06990923, 
    0.06971091, 0.06951259, 0.06941342, 0.06941342, 0.06941342, 0.06941342, 
    0.06941342, 0.06941342, 0.06941342,
  0.07061216, 0.07041199, 0.07021181, 0.07001164, 0.06981146, 0.06961128, 
    0.06941111, 0.06921093, 0.06912883, 0.0691648, 0.06920077, 0.06923673, 
    0.0692727, 0.06930867, 0.06934464,
  0.07001173, 0.06983684, 0.06966195, 0.06948706, 0.06931216, 0.06913728, 
    0.06896238, 0.06878749, 0.06875634, 0.06886895, 0.06898155, 0.06909415, 
    0.06920676, 0.06931936, 0.06943196,
  0.06940359, 0.06925463, 0.06910566, 0.0689567, 0.06880774, 0.06865878, 
    0.06850982, 0.06836086, 0.0683815, 0.06857174, 0.06876198, 0.06895223, 
    0.06914247, 0.0693327, 0.06952295,
  0.06879488, 0.06867187, 0.06854886, 0.06842586, 0.06830285, 0.06817984, 
    0.06805684, 0.06793383, 0.0680063, 0.06827425, 0.0685422, 0.06881016, 
    0.06907811, 0.06934606, 0.06961402 ;

 sftof =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100 ;

 time = 0 ;

 wet =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wet_c =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wet_u =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 wet_v =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 xh = -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 xq = -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 yh = -14.3476556382336, -14.1053228834302, -13.862732304759, 
    -13.6198879813569, -13.3767940148509, -13.1334545290505, 
    -12.889873669635, -12.6460556038367, -12.4020045201193, -12.1577246278516 ;

 yq = -14.4687240631789, -14.2265217428746, -13.9840595676627, 
    -13.7413416053212, -13.4983719462701, -13.2551547032665, 
    -13.011694011094, -12.7679940262485, -12.5240589266184, -12.279892911161 ;
}
