netcdf \00010101.tas.atmos_daily.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	grid_xt = 15 ;
	grid_yt = 10 ;
	scalar_axis = 1 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:_FillValue = NaN ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	float tas(time, grid_yt, grid_xt) ;
		tas:_FillValue = 1.e+20f ;
		tas:missing_value = 1.e+20f ;
		tas:units = "K" ;
		tas:long_name = "Near-Surface Air Temperature" ;
		tas:cell_methods = "time: mean" ;
		tas:cell_measures = "area: area" ;
		tas:coordinates = "height2m" ;
		tas:time_avg_info = "average_T1,average_T2,average_DT" ;
		tas:standard_name = "air_temperature" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Wed Apr 30 14:48:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.atmos_daily.tile3.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.atmos_daily.tile3.nc\nFri Apr 25 14:15:06 2025: ncks -x -v sphum,psl 00010101.atmos_daily.tile3.nc -o reduce/00010101.atmos_daily.tile3.nc\nFri Apr 25 13:47:12 2025: ncks -d grid_xt,35,55 -d grid_yt,30,45 00010101.atmos_daily.tile3.nc var_select/00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 grid_xt = 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50 ;

 grid_yt = 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 height10m = 10 ;

 height2m = 2 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 scalar_axis = 0 ;

 tas =
  257.3323, 260.88, 257.5914, 259.1828, 258.3731, 255.5161, 256.0681, 
    256.0787, 254.784, 245.458, 247.9986, 247.0397, 242.3113, 243.4877, 
    238.1712,
  261.7868, 261.0693, 259.9989, 260.6577, 257.3373, 254.8879, 256.6866, 
    255.6404, 255.6418, 252.3849, 248.9996, 251.1672, 249.5659, 242.117, 
    238.2685,
  261.2714, 260.4882, 260.0078, 259.9549, 256.8253, 247.2238, 254.6864, 
    254.5843, 254.7667, 253.9407, 252.5523, 252.8993, 252.4525, 250.1712, 
    245.3846,
  262.394, 260.1046, 259.1379, 258.8006, 257.9276, 254.2534, 241.7579, 
    250.6201, 254.1058, 253.2135, 252.5095, 253.0166, 253.0879, 252.2941, 
    248.6708,
  264.9443, 261.4029, 259.3835, 258.444, 257.8813, 256.7296, 253.1776, 
    239.6601, 239.8034, 245.3244, 251.4951, 252.5442, 253.1486, 253.2319, 
    251.9598,
  265.8576, 263.0153, 260.1853, 258.9289, 258.0598, 257.1744, 255.4048, 
    253.9191, 249.6825, 246.9975, 247.8435, 252.8719, 253.466, 254.0337, 
    253.442,
  265.8682, 263.2753, 260.8395, 259.4356, 258.5786, 257.6841, 256.6308, 
    255.1561, 253.8207, 253.3743, 253.2192, 253.4531, 253.9817, 254.3997, 
    254.1335,
  264.7134, 262.8682, 261.0251, 259.8904, 258.8793, 258.1032, 257.1086, 
    256.0076, 255.1823, 254.9045, 254.5466, 254.4372, 254.9967, 255.3217, 
    255.2251,
  264.0444, 262.2692, 260.952, 259.9066, 259.0594, 258.1192, 257.2582, 
    256.5033, 255.9284, 255.4713, 255.2423, 255.1285, 255.3839, 255.2261, 
    254.2033,
  263.4248, 262.0819, 261.0137, 260.0119, 259.1375, 258.1608, 257.1331, 
    255.9644, 254.3446, 251.7746, 253.3735, 254.8599, 254.9076, 254.7921, 
    254.2934,
  258.4195, 263.5067, 257.9645, 261.2277, 258.3206, 256.5709, 256.9903, 
    255.5727, 253.5879, 250.0532, 251.866, 252.4058, 250.5711, 249.7602, 
    246.6446,
  265.9001, 264.9107, 263.3162, 261.9574, 257.01, 255.5386, 257.9186, 
    256.5347, 255.1877, 253.2882, 252.6958, 254.0507, 252.3513, 246.4025, 
    244.6697,
  265.9961, 265.311, 264.2448, 262.6939, 258.1933, 246.9427, 257.6172, 
    257.5423, 256.6671, 255.294, 255.1433, 254.9729, 253.8484, 252.1565, 
    247.8858,
  265.7617, 264.8673, 264.0826, 262.6717, 260.953, 257.4916, 245.9679, 
    256.7961, 257.4683, 256.1368, 255.9548, 255.5407, 254.4773, 252.6647, 
    249.0741,
  265.794, 264.7625, 263.8561, 262.7377, 261.4766, 260.1553, 257.4985, 
    246.6585, 247.5201, 253.6317, 256.0474, 255.7959, 255.1737, 253.8013, 
    252.096,
  265.9899, 265.0357, 264.1097, 263.1571, 262.0897, 261.0681, 260.0819, 
    258.9783, 256.0976, 254.7907, 253.9639, 256.3376, 255.8681, 255.2225, 
    253.9363,
  266.321, 265.3523, 264.4941, 263.6087, 262.7368, 261.795, 260.968, 
    260.1318, 259.3445, 258.7122, 257.3122, 256.7181, 256.4186, 255.9225, 
    254.7222,
  266.5473, 265.7186, 264.8308, 264.1199, 263.3368, 262.6262, 261.8524, 
    261.0756, 260.3412, 259.5369, 258.0516, 257.0339, 256.8534, 256.5387, 
    255.6746,
  266.6315, 265.8673, 265.058, 264.3089, 263.6638, 263.0876, 262.5147, 
    261.9573, 261.2803, 260.2654, 258.9274, 257.6666, 257.4537, 256.9272, 
    255.7152,
  266.4758, 265.7392, 265.1261, 264.3718, 263.6382, 262.9539, 262.3299, 
    261.4855, 260.2487, 257.9246, 258.24, 258.1395, 257.8662, 257.3954, 
    256.1844,
  264.8817, 266.1729, 261.5373, 264.5287, 262.3291, 259.007, 259.615, 
    259.4613, 258.6757, 251.8968, 252.1595, 250.7152, 249.4279, 250.7593, 
    248.4598,
  267.0686, 266.3005, 265.59, 264.7638, 259.4618, 257.2405, 260.2491, 
    259.6976, 259.0996, 255.5653, 252.9476, 253.2618, 253.5601, 249.1061, 
    247.1831,
  267.0357, 266.2807, 265.7342, 265.3151, 262.6158, 250.0694, 259.1555, 
    259.5745, 259.4631, 256.877, 255.4082, 255.2333, 255.3061, 255.176, 
    251.4025,
  267.2388, 266.3228, 265.816, 265.4993, 265.3268, 262.2662, 247.7221, 
    258.1014, 259.5406, 257.5139, 256.6819, 256.5837, 256.5259, 255.7676, 
    253.0708,
  267.3807, 266.4816, 265.8221, 265.4841, 265.3559, 264.9973, 261.8337, 
    249.009, 251.1543, 256.7899, 257.9844, 257.7597, 257.3172, 256.5182, 
    255.2087,
  267.6126, 266.6355, 265.8995, 265.423, 265.2278, 265.0688, 264.3217, 
    262.0578, 259.6971, 258.9327, 258.1954, 258.3993, 257.8901, 257.4043, 
    256.267,
  267.7957, 266.8461, 265.9867, 265.3514, 264.9988, 264.8388, 264.5434, 
    263.5232, 262.6237, 261.9224, 259.7923, 258.9445, 258.3191, 258.0836, 
    257.421,
  267.8984, 266.9873, 266.0725, 265.3731, 264.8644, 264.5803, 264.4041, 
    263.9573, 263.426, 262.7862, 260.4153, 259.2509, 258.9382, 259.2151, 
    257.565,
  267.8848, 267.0353, 266.1555, 265.3666, 264.7422, 264.3532, 264.1173, 
    264.025, 263.7627, 262.9115, 260.6421, 259.4606, 259.4912, 258.6704, 
    256.0655,
  267.6209, 266.9453, 266.1505, 265.377, 264.6075, 264.1338, 263.8115, 
    263.4282, 262.5659, 260.7712, 260.062, 259.6225, 259.5226, 257.9076, 
    256.8581,
  265.3307, 267.6815, 265.287, 267.8759, 265.5076, 262.0374, 260.0273, 
    257.0714, 254.9016, 247.5133, 248.7244, 245.7773, 243.3002, 244.8995, 
    239.732,
  268.028, 268.6091, 268.3418, 268.0414, 259.3233, 258.0249, 262.9699, 
    260.1566, 257.6875, 252.7958, 249.4796, 249.2399, 249.4608, 242.7653, 
    239.8356,
  268.4381, 268.4102, 268.0788, 267.9126, 263.3148, 251.0186, 262.8719, 
    261.701, 259.5234, 255.1543, 252.4168, 250.9049, 250.8231, 251.2972, 
    247.365,
  268.7743, 268.3102, 267.9783, 267.7755, 267.7915, 264.0586, 252.6809, 
    260.3331, 259.163, 255.3308, 252.7828, 251.7216, 251.828, 252.2741, 
    249.7016,
  268.7004, 268.1188, 267.8112, 267.6877, 267.6169, 267.3391, 262.8741, 
    251.5352, 251.3353, 252.9356, 253.0122, 252.493, 253.1935, 253.8443, 
    252.6036,
  268.5504, 267.9759, 267.6951, 267.5922, 267.491, 267.5509, 264.7845, 
    262.036, 257.3742, 254.9909, 253.2083, 253.6988, 254.4558, 254.9148, 
    252.493,
  268.2882, 267.7722, 267.6339, 267.5068, 267.4101, 267.6233, 265.4738, 
    262.8179, 260.6687, 258.7798, 255.6227, 255.1654, 255.8626, 254.9632, 
    254.0325,
  267.9258, 267.5067, 267.5434, 267.58, 267.5914, 267.6478, 265.5717, 
    263.3784, 261.6208, 259.8746, 257.0966, 256.6601, 256.2859, 255.5382, 
    255.3462,
  267.3932, 267.054, 267.3965, 267.7781, 267.9869, 267.5893, 265.5294, 
    264.0406, 262.9866, 261.807, 258.539, 257.4994, 256.7362, 256.3883, 
    255.4601,
  266.7253, 266.4741, 267.3094, 267.9643, 268.0405, 267.1465, 265.7646, 
    264.8501, 263.4009, 260.1739, 258.4481, 258.1371, 257.4215, 256.8218, 
    256.9749,
  263.7388, 266.0892, 265.4207, 266.9755, 265.2805, 262.3929, 259.4987, 
    253.5452, 250.2994, 245.2825, 243.9145, 243.9747, 241.4598, 242.739, 
    235.3501,
  265.9181, 267.6089, 268.7134, 269.0177, 262.9244, 260.5416, 257.6, 
    253.9688, 251.7829, 248.5843, 245.8003, 249.1544, 250.5551, 239.6949, 
    234.32,
  266.5021, 268.1301, 269.2892, 269.4607, 264.3605, 254.7613, 257.9884, 
    255.2591, 252.874, 251.1072, 251.0354, 251.4341, 252.3463, 252.3648, 
    244.0658,
  267.2164, 268.7383, 269.6263, 269.7397, 267.1771, 261.2646, 252.4242, 
    255.4957, 254.4852, 253.5311, 252.3909, 252.3478, 253.1502, 252.9475, 
    247.9922,
  268.5041, 269.4616, 269.9313, 269.8966, 268.2724, 265.3022, 260.1832, 
    248.791, 247.1405, 251.7392, 252.8014, 253.1189, 254.1465, 254.6502, 
    254.6848,
  269.3052, 269.9691, 270.0798, 269.9434, 268.9583, 267.1946, 263.7658, 
    260.6551, 255.8736, 254.2922, 252.9526, 254.0236, 254.8953, 255.5856, 
    255.2288,
  270.028, 270.3344, 270.2048, 269.9011, 269.3083, 268.4337, 265.7514, 
    262.9851, 260.5612, 258.9066, 255.5496, 254.7047, 255.5749, 256.1443, 
    256.1703,
  270.6265, 270.5545, 270.1304, 269.8701, 269.5591, 269.0082, 266.5813, 
    264.2596, 262.1822, 260.2392, 255.8436, 255.3813, 256.3909, 256.7803, 
    256.7982,
  270.814, 270.4677, 270.0374, 269.8725, 269.7862, 269.2297, 266.8498, 
    264.8079, 263.4128, 261.1481, 256.7253, 256.0993, 257.0399, 257.2335, 
    257.0342,
  270.6309, 270.0197, 269.8553, 269.9848, 269.8315, 268.8926, 266.6781, 
    265.0884, 263.1579, 258.8529, 256.6241, 256.9835, 257.5314, 257.8186, 
    258.7262,
  258.3063, 261.551, 260.2991, 262.2397, 259.9857, 259.3553, 258.6271, 
    254.4759, 250.7405, 243.0442, 240.9002, 246.4113, 245.3392, 245.946, 
    238.3521,
  263.3137, 264.3396, 264.6923, 265.2455, 261.2976, 260.6928, 258.859, 
    254.5084, 251.6618, 247.9678, 243.3592, 251.8633, 254.8414, 243.1928, 
    238.2208,
  265.3065, 266.0053, 266.6342, 267.2016, 263.7721, 257.0653, 258.2126, 
    254.6103, 252.3125, 251.6917, 251.4116, 253.8957, 255.9269, 255.8112, 
    244.9305,
  266.1934, 267.2254, 267.8137, 268.5279, 266.7154, 261.7221, 252.1434, 
    253.5658, 252.9459, 253.1155, 252.6291, 254.2436, 256.045, 255.97, 
    249.6488,
  266.9051, 268.2055, 268.7317, 269.4453, 268.362, 265.1328, 258.9236, 
    246.5046, 244.0697, 249.687, 252.7664, 254.4636, 256.8286, 257.5292, 
    257.0929,
  267.4735, 268.9209, 269.3939, 270.0673, 269.5184, 267.262, 263.5881, 
    259.794, 255.7822, 253.6775, 251.9246, 255.5171, 257.1812, 257.8877, 
    258.0675,
  268.3259, 269.4926, 269.9936, 270.5302, 270.0976, 268.4454, 266.0225, 
    263.1385, 260.7491, 259.2345, 256.5536, 256.5992, 257.6497, 258.2121, 
    258.5763,
  269.2356, 270.1424, 270.5977, 270.8854, 270.3857, 268.9815, 267.0448, 
    264.7777, 262.7721, 260.8242, 257.3461, 257.1121, 258.0515, 258.5029, 
    258.8497,
  269.868, 270.6047, 271.0951, 271.1353, 270.4793, 269.2056, 267.456, 
    265.4526, 263.8731, 262.805, 258.3032, 257.598, 258.194, 258.7524, 
    259.2857,
  270.432, 271.0936, 271.3484, 271.1643, 270.4685, 269.2498, 267.5949, 
    265.9238, 264.1153, 261.0602, 257.914, 257.8605, 258.3088, 259.7871, 
    261.2979,
  255.3701, 260.928, 258.5592, 260.9637, 255.0942, 253.6112, 255.0205, 
    254.1837, 253.5668, 248.7037, 249.9864, 252.9385, 246.9239, 245.2027, 
    241.4923,
  262.3604, 264.0266, 263.6255, 263.4198, 255.7087, 255.3233, 256.5335, 
    254.4964, 254.3558, 254.4374, 252.6316, 257.0331, 254.7976, 242.6002, 
    240.3795,
  265.3595, 265.868, 265.651, 265.0709, 258.4506, 253.2494, 257.0582, 
    254.9836, 254.7559, 255.5965, 256.4105, 257.7479, 257.4135, 253.9538, 
    247.2568,
  266.9849, 267.091, 266.9767, 266.3509, 263.0956, 259.6412, 252.7452, 
    252.1804, 254.6701, 254.9503, 255.7989, 257.6583, 258.0068, 255.5361, 
    249.9919,
  267.9501, 268.2303, 267.9731, 267.5301, 265.3629, 263.5778, 259.3444, 
    245.8192, 241.6189, 249.5746, 255.2323, 257.7849, 258.593, 258.5909, 
    256.616,
  268.392, 269.0404, 268.868, 268.3834, 266.8857, 265.3727, 263.2414, 
    261.0809, 256.6454, 253.7554, 252.1223, 258.1288, 258.8893, 258.9619, 
    258.3636,
  268.7065, 269.5462, 269.5273, 269.2124, 268.0806, 266.9845, 265.5435, 
    263.9173, 262.3361, 261.3988, 258.6118, 258.3318, 259.3222, 259.322, 
    258.5659,
  269.2516, 270.0721, 270.108, 269.757, 268.9299, 268.2076, 267.2894, 
    266.2817, 264.5863, 262.7567, 258.6912, 258.3693, 259.5806, 260.3229, 
    259.6628,
  269.923, 270.3307, 270.4813, 270.3736, 269.6035, 269.0188, 268.49, 
    267.9973, 266.0159, 264.999, 259.2526, 258.3116, 259.2861, 260.7971, 
    260.6741,
  270.4945, 270.7377, 270.7202, 270.5041, 270.0132, 269.626, 269.3617, 
    269.0343, 267.1696, 262.9804, 258.5841, 258.5986, 258.9982, 260.8708, 
    261.4591,
  256.4575, 259.9048, 256.4776, 259.5357, 255.0092, 251.5162, 256.6388, 
    256.0074, 254.4076, 247.4821, 245.6482, 245.321, 242.5082, 243.5111, 
    239.5751,
  263.2191, 263.9157, 262.8735, 262.8359, 253.9149, 249.998, 256.9035, 
    256.8688, 256.2853, 253.7083, 248.7869, 251.4239, 250.5897, 241.1054, 
    239.1102,
  265.7437, 266.0631, 265.2372, 264.6524, 257.3415, 249.0667, 255.2661, 
    257.1474, 257.5252, 256.5814, 255.0711, 254.8181, 253.7286, 251.9109, 
    247.5736,
  267.1178, 267.3866, 266.7699, 266.229, 262.6827, 258.7065, 244.651, 
    254.0385, 258.0002, 257.3736, 256.69, 255.9005, 254.7933, 253.8242, 
    250.8465,
  267.9803, 268.3077, 267.7059, 267.3175, 264.9569, 263.5102, 259.8525, 
    244.5168, 245.8031, 253.3241, 257.5503, 257.0543, 256.0875, 255.2596, 
    254.4334,
  269.1581, 269.2145, 268.5342, 268.0807, 266.4607, 265.6214, 263.3329, 
    262.3401, 257.959, 256.6778, 255.1406, 257.9311, 257.1925, 256.8945, 
    256.2876,
  269.8601, 269.8972, 269.2123, 268.8992, 267.6745, 266.706, 265.2883, 
    264.2144, 263.3942, 261.83, 259.5067, 258.7238, 258.0258, 257.5331, 
    257.0362,
  270.7344, 270.5959, 270.0337, 269.5263, 268.6087, 267.8835, 266.2408, 
    265.7575, 264.8265, 262.7571, 259.5919, 259.3922, 259.0826, 258.1584, 
    256.9856,
  270.9873, 271.0766, 270.6587, 270.3081, 269.4305, 268.7176, 267.2906, 
    266.1491, 265.7184, 263.1708, 259.5326, 259.556, 259.5015, 258.5802, 
    257.0432,
  271.6677, 271.5526, 271.2346, 270.6179, 269.9028, 269.3555, 268.1402, 
    267.0258, 265.8508, 261.3515, 258.9904, 259.6124, 259.8883, 259.6475, 
    259.3957,
  259.1815, 259.3047, 254.4991, 256.6562, 254.4741, 252.5574, 252.2175, 
    250.7111, 249.1012, 242.3536, 242.8511, 244.7068, 242.4206, 243.7421, 
    238.8272,
  264.1339, 263.3508, 260.9655, 260.6194, 253.7837, 252.3157, 253.9767, 
    252.3288, 251.2334, 249.4319, 244.0919, 251.0351, 251.8144, 239.4827, 
    238.3457,
  266.3381, 265.8158, 264.0619, 262.9222, 256.6343, 248.1566, 255.2931, 
    254.2214, 253.0384, 252.1161, 252.2245, 253.3104, 253.8183, 252.9664, 
    247.2123,
  267.4371, 267.4362, 265.9833, 264.7889, 261.1805, 257.7495, 248.2008, 
    253.5465, 253.6865, 253.0365, 252.4984, 253.3332, 254.3906, 254.0646, 
    251.6165,
  268.6385, 268.6681, 267.2677, 266.2262, 263.507, 262.2214, 258.65, 
    247.3203, 245.3662, 250.1917, 253.1784, 253.9184, 255.0528, 255.3199, 
    255.6216,
  269.664, 269.5162, 268.2135, 267.135, 265.2359, 264.68, 262.6611, 260.6188, 
    256.9706, 254.7033, 252.7623, 254.6399, 255.4936, 255.9221, 256.3023,
  270.4502, 270.2771, 268.9267, 268.0286, 266.4771, 266.0728, 265.0828, 
    263.8836, 262.2934, 259.844, 256.6294, 255.8884, 255.8844, 256.2808, 
    256.9631,
  271.149, 270.6967, 269.4602, 268.5069, 267.3358, 267.1356, 266.4841, 
    266.2786, 265.0051, 262.8345, 258.0592, 256.9977, 256.3794, 256.8242, 
    256.9965,
  271.6605, 270.9505, 269.9962, 269.3027, 268.2464, 267.8611, 267.2777, 
    267.1649, 266.745, 264.7853, 258.8828, 257.9467, 257.0554, 257.1374, 
    256.2411,
  271.7729, 271.1689, 270.3295, 269.5067, 268.7239, 268.6031, 267.9097, 
    267.6945, 266.6959, 262.1588, 259.3223, 258.8812, 257.7623, 257.6142, 
    256.9861,
  254.0506, 256.4793, 252.272, 254.7029, 252.1729, 250.9539, 253.2732, 
    253.3156, 253.6395, 248.759, 248.3612, 251.5975, 248.1538, 246.5371, 
    241.212,
  260.6561, 261.0045, 259.2006, 258.3174, 250.6835, 249.3638, 253.586, 
    253.6698, 253.7142, 253.4234, 249.7865, 254.9774, 255.7064, 247.0429, 
    245.3867,
  263.9216, 263.5658, 262.1027, 260.7979, 253.8179, 245.3074, 252.2366, 
    253.675, 253.7082, 253.7276, 254.0407, 255.1429, 256.5381, 257.1322, 
    252.6691,
  266.2963, 265.5283, 264.357, 263.2907, 260.0318, 255.5875, 245.5522, 
    250.082, 253.1901, 252.7981, 253.1886, 254.5677, 256.2807, 257.4915, 
    256.7227,
  268.0628, 267.1038, 265.8939, 265.2008, 262.9655, 261.4009, 257.5215, 
    242.1269, 241.3891, 247.4654, 252.5798, 254.5748, 256.4317, 258.0105, 
    259.4053,
  269.2281, 268.4021, 267.2635, 266.6292, 265.2382, 263.9161, 262.1067, 
    260.6917, 255.0324, 251.4244, 249.7093, 254.8932, 256.4221, 258.1982, 
    259.5412,
  270.4202, 269.6149, 268.4474, 267.8961, 266.8626, 266.2625, 264.4746, 
    263.7126, 261.8652, 259.3484, 256.3375, 255.4884, 256.7355, 258.3315, 
    259.7367,
  271.238, 270.5978, 269.4223, 268.9442, 267.8956, 267.5809, 266.7641, 
    265.7844, 264.672, 261.7613, 256.8034, 256.1253, 256.8166, 258.1479, 
    259.1524,
  272.1782, 271.4579, 270.2673, 269.7816, 269.0089, 268.5497, 268.0008, 
    267.4334, 266.0517, 263.92, 257.4783, 256.5437, 256.6637, 258.075, 
    258.3637,
  272.5002, 272.0954, 271.0434, 270.4287, 269.3546, 269.1471, 268.6277, 
    268.2167, 266.9148, 261.5544, 258.0495, 257.3105, 256.4568, 257.6357, 
    258.6771,
  251.3518, 256.2884, 251.4619, 256.9149, 253.4772, 250.5583, 254.6365, 
    254.9102, 256.0606, 253.1933, 252.6712, 254.5661, 249.8551, 248.4561, 
    243.4991,
  259.598, 261.1288, 260.5751, 259.9828, 248.5528, 248.3379, 254.2906, 
    254.9738, 255.7016, 256.7656, 255.2564, 258.4642, 257.4947, 246.4094, 
    246.3481,
  263.03, 263.4658, 263.1879, 262.4984, 254.8296, 244.8416, 251.85, 254.7777, 
    256.1688, 257.0882, 258.6998, 259.9112, 260.2076, 259.5191, 256.0626,
  265.4008, 265.3688, 264.952, 264.0642, 263.0612, 258.5235, 244.5497, 
    251.6597, 255.6372, 256.6847, 258.8714, 260.2693, 261.035, 260.8629, 
    259.7185,
  267.0507, 266.7151, 266.2579, 265.8519, 264.6588, 264.6275, 261.4017, 
    244.717, 248.2613, 254.5169, 258.9848, 260.5207, 261.2843, 261.2169, 
    261.6492,
  268.5258, 268.0256, 267.4233, 267.07, 266.4538, 265.7045, 265.459, 
    262.7587, 255.312, 255.1304, 257.9082, 260.6659, 261.1242, 261.1045, 
    261.5522,
  270.3939, 269.8238, 269.0287, 268.5173, 268.0542, 267.4944, 266.3038, 
    265.203, 262.1508, 260.3956, 260.005, 261.2099, 261.8083, 261.1433, 
    261.2982,
  271.8787, 271.4192, 270.585, 269.9702, 269.3982, 268.7705, 268.0168, 
    267.0116, 264.659, 261.1327, 259.3006, 260.9161, 261.7086, 261.369, 
    261.3121,
  273.5677, 272.7421, 271.8651, 270.8911, 270.3731, 269.8552, 269.1769, 
    268.2859, 266.0712, 261.8447, 258.4483, 260.3934, 261.3514, 261.6814, 
    261.2168,
  274.4818, 273.4496, 272.6642, 271.7126, 270.6299, 270.0741, 269.4341, 
    268.746, 266.658, 261.0377, 257.1858, 259.7336, 260.4872, 261.3504, 
    261.5387,
  251.1298, 258.1656, 255.5475, 260.3839, 255.4176, 250.9586, 257.0022, 
    258.4987, 259.6558, 255.2812, 255.0891, 257.7087, 255.3968, 254.5242, 
    251.3313,
  260.3768, 262.8015, 264.9719, 264.9512, 252.4708, 249.3505, 256.5626, 
    258.2149, 259.023, 258.9817, 256.84, 260.058, 260.4131, 253.2544, 253.5606,
  263.9255, 264.9151, 265.9559, 266.2476, 259.7042, 249.1599, 252.9063, 
    258.3165, 259.1786, 259.0241, 258.9068, 259.585, 260.128, 260.2863, 
    259.0736,
  266.3262, 266.5, 266.8105, 267.1654, 267.4748, 261.5528, 244.6734, 
    253.1207, 258.3088, 258.3365, 258.3602, 258.6823, 259.3047, 259.5177, 
    259.6159,
  267.532, 267.9963, 268.153, 268.3928, 267.9773, 267.5358, 260.8789, 
    244.9849, 250.5103, 253.3208, 257.5185, 258.0836, 258.5456, 258.7548, 
    259.4143,
  268.3642, 269.0548, 269.322, 269.3376, 268.9871, 268.1062, 265.5541, 
    262.0913, 255.7416, 255.9015, 257.1538, 257.8635, 258.0925, 258.2563, 
    258.5999,
  269.3878, 269.7446, 270.0349, 270.1533, 270.1119, 269.3662, 267.5756, 
    264.1504, 262.1534, 261.6409, 258.8441, 258.3434, 258.1793, 258.1318, 
    258.1965,
  272.4273, 271.6618, 271.1078, 270.6648, 270.4993, 270.0649, 269.1066, 
    266.8956, 264.5838, 262.2139, 258.444, 258.401, 258.3921, 258.3224, 
    258.1372,
  273.9364, 273.3746, 273.1069, 272.5089, 271.6328, 270.855, 270.122, 
    268.916, 267.2025, 263.3419, 258.6857, 258.1458, 258.1569, 258.6447, 
    258.4234,
  272.9722, 272.5993, 272.6881, 272.6526, 272.2683, 271.4107, 270.5769, 
    269.6532, 267.9703, 261.5422, 258.8666, 259.1099, 257.8772, 258.508, 
    258.8515,
  251.4748, 257.5754, 257.2615, 261.0736, 258.5512, 252.1471, 257.5969, 
    257.6201, 257.6039, 253.7898, 253.2618, 256.1915, 255.8161, 255.619, 
    252.4745,
  260.0081, 262.8299, 265.7643, 266.9464, 255.953, 250.3214, 255.5097, 
    257.6269, 256.8755, 256.5717, 255.3365, 257.215, 258.1912, 254.1223, 
    253.4846,
  263.6912, 264.7297, 266.079, 267.9213, 263.1982, 251.4658, 253.3917, 
    256.1476, 256.4131, 256.3041, 256.1578, 257.2644, 258.0121, 258.7026, 
    258.1937,
  265.8808, 266.2977, 266.8733, 267.8567, 269.0905, 264.144, 250.2079, 
    251.8205, 255.4237, 255.6549, 255.6418, 256.9537, 257.4998, 258.2439, 
    258.8829,
  266.75, 267.2828, 267.7473, 268.4853, 269.4026, 269.257, 263.5428, 
    245.1172, 245.5228, 253.0838, 255.9471, 256.9338, 256.9729, 257.4362, 
    259.0293,
  267.4753, 268.1281, 268.5903, 269.1103, 269.7966, 269.9477, 267.8034, 
    263.5957, 256.3686, 254.8085, 255.7297, 257.5543, 257.0799, 257.0828, 
    258.0797,
  268.1358, 268.8087, 269.3417, 269.5492, 269.9612, 270.1977, 269.3914, 
    267.2127, 263.9999, 262.1199, 259.8435, 258.9919, 257.8955, 256.9095, 
    257.6931,
  269.8609, 269.6261, 269.8396, 269.8454, 270.0608, 270.2669, 270.2097, 
    269.1236, 267.7457, 265.4017, 261.7457, 260.3145, 259.0547, 257.4308, 
    257.6157,
  272.0969, 271.6987, 271.3592, 271.0307, 270.8008, 270.7146, 270.641, 
    270.2245, 269.5156, 268.0262, 264.5821, 262.106, 260.1104, 258.2088, 
    258.4668,
  272.5998, 272.2103, 272.3004, 272.0987, 271.8099, 271.4663, 271.2104, 
    270.7668, 269.5345, 268.0632, 266.6506, 264.089, 261.4739, 259.3144, 
    258.1603,
  254.2537, 256.6355, 255.215, 256.0981, 256.0715, 254.9958, 256.4727, 
    256.1218, 255.3531, 252.0851, 252.8211, 254.6061, 254.5131, 255.122, 
    251.2309,
  260.7879, 262.1843, 261.8053, 260.9195, 254.8061, 252.9814, 255.7133, 
    256.8172, 255.7622, 254.2496, 253.0187, 257.3255, 258.6928, 253.271, 
    252.875,
  264.1798, 265.1383, 265.0622, 264.5359, 260.5747, 248.7373, 257.4516, 
    256.4265, 255.5803, 254.8189, 255.5682, 259.0695, 259.7122, 259.4858, 
    258.2783,
  266.0857, 266.679, 266.6833, 266.6926, 266.0689, 263.5092, 254.3378, 
    254.0643, 256.9022, 255.6139, 256.0433, 259.742, 260.0753, 259.9286, 
    259.0698,
  267.3743, 267.6232, 267.6528, 267.8461, 268.0077, 268.1451, 266.5733, 
    256.9766, 254.0376, 256.8496, 256.933, 260.8406, 261.0727, 260.6074, 
    259.7874,
  268.347, 268.4664, 268.466, 268.6172, 268.8451, 269.1697, 269.3747, 
    268.3267, 263.8708, 260.3939, 259.2392, 262.2594, 262.8353, 261.8409, 
    260.9899,
  268.9131, 269.0905, 269.0804, 269.1468, 269.3216, 269.5037, 269.7141, 
    269.7245, 268.4256, 266.8198, 264.5587, 264.487, 264.7357, 263.6543, 
    262.1187,
  269.288, 269.4678, 269.5529, 269.6391, 269.7632, 269.9025, 269.9716, 
    270.1122, 269.912, 268.6442, 267.4773, 266.7428, 266.2063, 264.8476, 
    263.8139,
  269.6566, 269.8512, 270.0358, 270.0811, 270.1688, 270.2596, 270.2822, 
    270.2683, 270.2663, 268.6268, 267.5895, 266.9169, 266.8442, 265.7008, 
    264.9578,
  270.4185, 270.4069, 270.6117, 270.7422, 270.7599, 270.7462, 270.7188, 
    270.6073, 269.8381, 267.9555, 269.0469, 268.7271, 267.9242, 266.8677, 
    265.9135,
  256.2137, 257.3112, 256.4611, 256.6671, 254.5339, 252.9526, 254.4218, 
    254.8028, 254.3801, 250.8562, 250.7362, 254.1186, 254.8167, 257.0892, 
    251.5103,
  260.0779, 261.5323, 261.0429, 258.7359, 253.8519, 252.9793, 255.7135, 
    255.5629, 255.8301, 255.5578, 253.7564, 257.1118, 260.6888, 259.3639, 
    252.1589,
  263.2432, 264.1591, 263.8033, 261.7774, 256.4984, 249.2654, 255.5865, 
    257.1783, 258.1305, 258.7439, 258.9772, 261.5886, 262.9193, 263.3693, 
    256.0394,
  265.2905, 265.831, 265.3568, 264.0045, 262.1704, 258.6005, 249.4777, 
    253.4638, 260.9959, 263.316, 262.2112, 264.0138, 264.7979, 264.1145, 
    258.0883,
  266.7109, 266.9538, 266.4325, 265.5354, 264.4614, 263.6372, 261.7689, 
    253.4247, 257.2867, 263.4835, 264.5669, 265.4135, 265.6237, 265.2708, 
    260.6685,
  267.847, 267.8317, 267.332, 266.7224, 266.2701, 265.8301, 265.4892, 
    265.6698, 263.7954, 265.5586, 265.3403, 266.2545, 266.291, 265.8899, 
    263.1181,
  268.7971, 268.687, 268.0964, 267.7002, 267.5462, 267.3982, 267.1606, 
    267.6716, 267.4936, 268.0496, 267.4427, 266.9215, 266.7505, 266.2032, 
    264.2181,
  269.7565, 269.4162, 268.9122, 268.5903, 268.4969, 268.4546, 268.4716, 
    268.7126, 269.1453, 267.2132, 266.0023, 266.6056, 267.1425, 266.99, 
    265.4037,
  270.2204, 269.9352, 269.465, 269.1904, 269.1461, 269.1446, 269.2343, 
    269.3748, 269.6686, 267.9492, 266.8137, 267.7103, 267.8554, 267.6166, 
    266.9872,
  270.5508, 270.1873, 269.9648, 269.754, 269.6401, 269.6602, 269.7353, 
    269.8294, 269.1209, 266.7704, 268.1525, 268.6438, 268.414, 268.3237, 
    268.1249,
  254.1298, 255.5388, 254.5988, 255.6738, 253.5808, 251.3834, 253.1429, 
    254.1715, 256.3159, 257.9981, 256.9775, 256.8521, 251.3451, 247.0907, 
    240.5879,
  260.0175, 260.9012, 260.1412, 257.258, 252.6201, 250.7279, 254.7021, 
    255.0525, 257.628, 260.9386, 260.963, 261.355, 259.1384, 250.2626, 
    246.2203,
  263.8754, 264.1461, 263.776, 261.4308, 255.8932, 247.1763, 254.0671, 
    255.8237, 259.2769, 263.309, 264.8919, 265.4019, 263.3325, 261.0386, 
    253.957,
  266.1323, 266.1333, 265.7102, 264.2238, 262.1826, 258.119, 248.0931, 
    253.502, 260.8589, 264.7313, 265.3195, 265.9071, 265.6678, 264.2436, 
    259.0954,
  267.6771, 267.5475, 267.1957, 266.1473, 264.8078, 263.6344, 260.4076, 
    248.6175, 255.1071, 262.4748, 265.4934, 266.1083, 265.9584, 265.6263, 
    262.4261,
  268.6801, 268.6203, 268.3064, 267.5637, 266.5449, 265.6842, 264.3877, 
    263.1108, 259.9316, 263.5818, 264.7414, 266.2664, 266.2771, 264.3532, 
    265.0981,
  269.5336, 269.5723, 269.3247, 268.7288, 267.8742, 267.2273, 266.271, 
    265.7421, 265.3509, 265.4273, 266.1663, 266.2698, 266.4872, 265.3557, 
    266.5482,
  270.201, 270.3211, 270.1051, 269.6121, 268.7678, 268.1039, 267.3481, 
    267.1068, 266.6769, 265.092, 265.3545, 266.1168, 266.6178, 266.7683, 
    267.2131,
  270.6389, 270.7616, 270.6375, 270.2094, 269.5559, 268.9904, 268.306, 
    267.7634, 267.6354, 266.3441, 264.1261, 263.5951, 265.8702, 266.3677, 
    267.2739,
  271.1161, 270.9012, 270.6461, 270.2625, 269.7005, 269.1601, 268.766, 
    268.3674, 267.7031, 263.6053, 265.0871, 265.1579, 265.0616, 266.5992, 
    267.409,
  251.7237, 253.8636, 252.609, 255.3042, 252.996, 249.8794, 256.3229, 
    258.7831, 261.4239, 261.2432, 261.0261, 262.7396, 261.4745, 259.2573, 
    251.3283,
  258.4475, 259.2883, 259.081, 256.4693, 249.2268, 247.1966, 254.6468, 
    257.5096, 260.3648, 262.6546, 262.3673, 263.9315, 264.2355, 259.8533, 
    252.4997,
  262.2755, 262.8363, 263.0106, 261.3116, 255.52, 242.1468, 252.7805, 
    255.4937, 259.3125, 262.0901, 263.4311, 264.211, 264.5453, 262.1547, 
    255.4236,
  264.5323, 264.9497, 265.0546, 264.5194, 262.9933, 259.7906, 247.401, 
    253.5792, 258.0662, 261.3265, 262.8623, 263.8898, 264.5527, 262.5461, 
    256.749,
  266.1783, 266.5874, 266.7079, 266.5326, 265.8266, 265.3184, 262.9197, 
    249.3638, 247.635, 257.4023, 262.0176, 262.9948, 264.3946, 263.4464, 
    259.5081,
  267.4649, 267.7794, 267.7647, 267.6729, 267.5071, 267.3572, 266.8393, 
    265.0044, 261.1906, 258.9012, 258.7775, 262.5439, 264.0942, 263.7837, 
    260.7712,
  268.4588, 268.8421, 268.7882, 268.7321, 268.656, 268.5356, 268.3555, 
    267.8655, 266.4265, 263.7966, 262.1871, 262.1856, 263.9459, 264.1615, 
    262.2215,
  269.5579, 269.7522, 269.7327, 269.6562, 269.5591, 269.4687, 269.1848, 
    268.9517, 268.2514, 265.4143, 262.4869, 262.06, 262.8097, 263.4444, 
    263.5883,
  270.8296, 270.7701, 270.7469, 270.5829, 270.3504, 270.1627, 269.9298, 
    269.3371, 268.9962, 267.1087, 263.5089, 262.1199, 261.5534, 261.5568, 
    264.5491,
  271.6739, 271.5235, 271.4148, 271.2572, 271.0411, 270.7413, 270.4317, 
    270.0614, 268.9737, 265.9923, 265.2143, 263.4498, 261.1575, 260.8115, 
    264.4354,
  253.7856, 257.5047, 256.6837, 257.4397, 253.7209, 251.006, 255.7431, 
    256.3353, 256.8138, 251.4669, 251.2189, 250.0179, 242.4027, 238.5717, 
    233.8269,
  261.4966, 262.0888, 262.0203, 258.639, 248.0699, 248.7615, 255.9968, 
    257.4632, 257.9191, 255.2384, 252.3415, 253.2758, 247.0114, 236.0046, 
    233.379,
  264.2643, 264.1443, 263.9852, 263.0138, 258.0779, 246.4182, 255.7867, 
    258.6252, 259.4067, 257.8009, 256.284, 254.2632, 249.3259, 244.8745, 
    238.9988,
  265.6555, 265.35, 265.2653, 265.3431, 266.0331, 264.5169, 255.2161, 
    259.6151, 261.0479, 258.8628, 256.9828, 255.6261, 250.66, 246.4339, 
    242.7386,
  266.8566, 266.8657, 266.9783, 267.3582, 267.7369, 268.4116, 267.7143, 
    257.1516, 257.9552, 258.5409, 257.6161, 256.1548, 252.6582, 248.7307, 
    247.5664,
  268.4935, 268.1674, 268.1861, 268.4235, 268.9429, 269.2134, 269.4856, 
    268.6324, 264.9613, 261.564, 257.036, 257.0927, 254.7279, 250.7239, 
    249.4696,
  268.7256, 269.4347, 269.5846, 269.8102, 270.0112, 270.1443, 270.0646, 
    269.7838, 268.3782, 265.1837, 261.0966, 258.5589, 257.4573, 252.9461, 
    251.0309,
  268.8826, 269.7399, 270.2597, 270.4238, 270.619, 270.5218, 270.3092, 
    270.0799, 269.2502, 266.1258, 262.3786, 260.012, 260.0596, 255.4888, 
    253.0093,
  269.1195, 269.9045, 270.4773, 270.7093, 270.7286, 270.5913, 270.4294, 
    270.082, 269.7229, 267.3597, 263.2688, 261.3626, 259.7808, 259.5333, 
    254.8144,
  270.2254, 270.6527, 270.9997, 271.1496, 270.9953, 270.7122, 270.1931, 
    269.8551, 268.8622, 265.9586, 265.0269, 262.5645, 260.4671, 259.1024, 
    259.8987,
  257.8344, 259.7687, 254.79, 258.9764, 256.9288, 255.4048, 258.4957, 
    256.9781, 251.3993, 240.9667, 239.272, 240.1165, 238.5169, 240.8279, 
    239.3152,
  263.1894, 263.4779, 263.7202, 262.2582, 257.0233, 256.3729, 260.8437, 
    260.6736, 255.3237, 248.4787, 242.7727, 246.0395, 246.8322, 239.0157, 
    239.9033,
  265.0423, 265.474, 266.0788, 266.42, 263.1072, 255.5142, 262.0499, 
    262.9249, 259.5766, 253.8702, 250.1864, 249.1053, 248.2043, 248.2803, 
    246.6315,
  266.8898, 266.5982, 266.7494, 267.6369, 269.4573, 268.5824, 260.9962, 
    263.5713, 260.7029, 256.3194, 252.1355, 250.1828, 249.1695, 248.9374, 
    248.7763,
  267.6216, 267.5119, 267.7652, 268.9803, 269.9666, 270.7905, 269.7197, 
    261.7962, 259.5465, 257.4852, 254.3103, 251.8103, 249.9066, 249.8912, 
    250.8224,
  269.0637, 269.0292, 269.283, 270.0934, 270.7227, 271.0383, 270.7975, 
    268.8441, 262.7065, 258.7459, 254.3557, 253.0943, 251.2292, 250.4276, 
    251.2654,
  269.5643, 270.2242, 270.5268, 270.7543, 270.9443, 271.0456, 270.7656, 
    270.0775, 267.053, 262.5625, 258.5246, 255.0458, 252.6822, 251.539, 
    251.9698,
  269.4225, 270.1541, 270.6562, 270.7984, 270.9957, 270.9279, 270.5227, 
    270.1148, 268.7034, 264.0434, 259.7708, 256.7861, 254.9198, 252.7532, 
    252.7088,
  269.5384, 270.185, 270.6951, 270.7838, 270.8942, 270.6533, 270.2433, 
    269.5279, 269.1212, 267.3609, 263.5305, 260.7921, 258.0723, 255.2641, 
    252.902,
  269.8277, 270.2248, 270.3401, 270.5643, 270.4968, 270.0232, 269.3397, 
    268.8289, 266.9342, 264.1447, 264.6771, 262.6597, 260.3912, 257.401, 
    254.0941,
  254.271, 257.6601, 255.49, 259.5291, 259.6518, 260.0761, 262.4342, 
    261.9334, 257.9815, 254.3659, 251.7252, 250.6417, 245.698, 246.419, 
    244.7365,
  260.9462, 262.5102, 264.3029, 263.9657, 259.8729, 260.2091, 263.3759, 
    262.4229, 260.1621, 259.443, 255.228, 254.8116, 251.6022, 245.166, 
    245.2663,
  264.2034, 265.1469, 266.3984, 267.4143, 265.2741, 259.5515, 263.74, 
    263.1988, 261.7181, 259.9156, 259.2646, 256.8235, 252.4866, 252.2813, 
    251.1718,
  265.9799, 266.4868, 267.3884, 268.1222, 269.3961, 268.7299, 259.4549, 
    263.0106, 263.0056, 261.2347, 259.6438, 257.3289, 253.2549, 252.8575, 
    252.4457,
  267.5647, 267.9013, 268.3119, 268.9786, 269.8465, 270.5596, 269.5997, 
    263.5286, 262.3862, 260.9483, 259.6681, 257.4217, 254.3604, 253.4064, 
    254.1855,
  267.7407, 268.7747, 269.2903, 269.8101, 270.4078, 270.6476, 270.6185, 
    269.1063, 264.9124, 264.1298, 261.0513, 259.0657, 255.4013, 253.7199, 
    254.3574,
  267.4933, 268.7953, 269.5848, 270.0937, 270.4296, 270.5516, 270.5421, 
    270.235, 268.7501, 266.1606, 264.0876, 260.3978, 257.285, 253.854, 
    254.2986,
  267.8911, 268.872, 269.611, 270.0942, 270.3641, 270.4494, 270.3687, 
    270.0744, 268.9959, 266.6592, 264.0078, 261.3468, 258.7222, 255.0726, 
    254.1864,
  268.783, 269.3548, 269.9934, 270.2041, 270.3257, 270.3144, 270.1609, 
    269.4116, 269.0736, 266.6812, 263.7678, 262.2555, 259.9921, 257.1347, 
    253.3985,
  269.9877, 270.1105, 270.2962, 270.271, 270.2601, 269.9309, 269.2354, 
    269.1106, 268.1334, 263.3872, 263.4807, 263.3427, 261.0455, 260.1496, 
    253.8775,
  255.4069, 256.9309, 256.0608, 257.0029, 256.6743, 256.7037, 258.241, 
    259.3499, 259.6894, 259.0974, 258.3986, 258.0316, 256.2029, 251.7117, 
    245.1268,
  260.0361, 260.7087, 262.1197, 261.2943, 256.9012, 257.0031, 259.9251, 
    260.6518, 261.2182, 260.9911, 259.7808, 260.2472, 259.1828, 250.4243, 
    243.017,
  263.6713, 264.1853, 264.8343, 265.6076, 264.0156, 256.3794, 261.535, 
    262.0851, 262.3372, 262.1799, 262.112, 261.7324, 260.057, 256.0956, 
    245.9969,
  265.0417, 265.8643, 266.6034, 267.077, 267.9865, 266.9644, 257.7343, 
    261.9766, 263.3617, 263.543, 263.1222, 262.5661, 260.9306, 256.8888, 
    247.1881,
  266.2933, 267.2607, 267.8829, 268.5442, 269.0599, 269.4815, 268.8994, 
    260.8501, 262.3922, 263.6018, 263.6846, 262.719, 260.8986, 257.1858, 
    250.1077,
  266.9616, 268.2073, 269.0388, 269.4793, 269.9507, 270.1185, 270.1895, 
    269.2418, 266.2339, 264.0376, 263.317, 263.2898, 261.4755, 257.7567, 
    252.0161,
  268.3389, 269.3392, 269.9666, 270.3301, 270.5866, 270.6443, 270.5847, 
    270.3639, 269.5152, 267.4001, 265.7501, 264.541, 262.0485, 257.5496, 
    252.8913,
  270.7804, 271.265, 271.5578, 271.5699, 271.4505, 271.229, 270.9357, 
    270.557, 269.6799, 267.7984, 266.0793, 264.6606, 262.5312, 257.7641, 
    252.5165,
  272.9351, 272.8693, 272.7895, 272.3145, 271.7802, 271.3979, 270.8096, 
    269.5717, 269.1667, 267.8662, 266.5225, 265.6629, 262.8972, 257.6485, 
    251.7264,
  273.7505, 273.2648, 272.744, 272.1843, 271.6802, 270.8782, 269.1656, 
    268.6997, 268.4132, 267.3793, 267.6388, 266.5082, 263.2381, 257.8376, 
    251.115,
  254.6025, 256.6662, 256.32, 257.0552, 256.2419, 255.9602, 256.7661, 
    256.4427, 256.2146, 254.8094, 254.8647, 254.7841, 254.904, 255.3461, 
    251.1108,
  259.5368, 259.9802, 261.4609, 260.3441, 255.723, 255.5828, 257.9084, 
    257.6319, 257.5477, 257.1013, 258.2742, 259.4896, 259.6608, 256.527, 
    249.6689,
  264.0153, 264.5183, 264.9369, 265.3447, 262.55, 257.5446, 260.2477, 
    260.2872, 260.1925, 260.6375, 261.7357, 262.7443, 262.3443, 260.6801, 
    250.4634,
  265.4158, 266.2932, 266.8226, 267.0667, 267.7005, 266.1432, 257.3379, 
    261.6977, 263.949, 264.6225, 265.8311, 265.4355, 264.5834, 261.9901, 
    249.1572,
  266.5512, 267.3652, 267.8382, 268.2959, 268.6169, 269.0224, 268.4316, 
    262.8643, 263.132, 267.5884, 268.2818, 266.069, 265.3011, 262.1951, 
    249.5864,
  268.4015, 268.4976, 268.5403, 268.9719, 269.3764, 269.7245, 270.0496, 
    269.8838, 269.0453, 268.9806, 267.4838, 264.9507, 264.992, 261.9881, 
    249.2243,
  270.7576, 270.3713, 269.9791, 269.9019, 270.2342, 270.4829, 270.7439, 
    270.8663, 270.5903, 268.9401, 265.5971, 264.664, 265.0036, 259.8151, 
    248.3624,
  272.7094, 272.1364, 271.5446, 271.1421, 271.0473, 271.1291, 271.0146, 
    270.8792, 269.692, 266.9723, 263.5905, 265.3908, 264.8295, 257.6038, 
    247.4078,
  273.8392, 273.2565, 272.7864, 272.015, 271.3741, 271.2135, 271.0898, 
    270.334, 269.2184, 266.9017, 263.7219, 265.8914, 262.9471, 253.8571, 
    244.2384,
  274.2626, 273.6176, 272.9914, 272.3781, 271.7513, 271.0574, 270.3246, 
    269.2733, 267.9839, 264.0583, 266.4434, 266.4375, 260.183, 250.6655, 
    244.6742,
  251.4518, 252.6309, 251.6436, 251.8808, 251.2999, 251.2402, 252.6035, 
    252.5155, 252.2221, 250.4683, 250.8584, 252.4182, 252.5967, 254.7872, 
    257.4705,
  257.3138, 257.0725, 257.2541, 255.7015, 250.9328, 252.5265, 254.5112, 
    253.7322, 253.6288, 253.0277, 252.3004, 254.7079, 256.4677, 258.2939, 
    258.6741,
  265.04, 263.544, 263.1587, 262.522, 256.4473, 250.3372, 256.0941, 255.9711, 
    255.2193, 254.8817, 255.4615, 256.9464, 259.4075, 261.5337, 254.8186,
  268.744, 267.8903, 266.7715, 266.113, 264.9064, 259.6106, 252.8219, 
    256.5002, 257.4211, 257.0174, 257.4586, 259.3693, 261.132, 261.5757, 
    250.5222,
  271.7055, 271.0109, 270.0084, 268.9932, 268.1934, 266.5665, 262.6368, 
    253.9166, 254.299, 259.3082, 260.7131, 261.623, 262.3359, 261.3553, 
    251.2902,
  273.1543, 273.0106, 272.4008, 271.4443, 270.5364, 269.6591, 267.9141, 
    264.9682, 260.5959, 260.1493, 260.9815, 262.5561, 263.2163, 259.2898, 
    250.0233,
  273.7628, 273.7663, 273.5549, 273.002, 272.226, 271.5085, 270.4946, 
    269.0688, 266.5399, 262.9309, 262.3425, 263.2092, 262.461, 256.0575, 
    249.2123,
  274.5389, 274.1824, 273.87, 273.5213, 272.9269, 272.3814, 271.5643, 
    270.7833, 269.3595, 265.3036, 263.5764, 263.7194, 261.7719, 253.6242, 
    248.0725,
  273.6856, 273.1642, 272.8891, 272.5515, 272.307, 272.0742, 271.6982, 
    271.0827, 270.2232, 267.4928, 264.7062, 264.281, 260.3667, 251.1544, 
    245.0355,
  272.4845, 271.7585, 271.3555, 271.3227, 271.4752, 271.4279, 271.1706, 
    270.8909, 270.3623, 268.3745, 266.0652, 264.5957, 258.5688, 248.9919, 
    245.6174,
  253.8294, 253.7306, 250.5761, 251.527, 250.3228, 249.7378, 252.2662, 
    250.8877, 249.6094, 244.7276, 245.0758, 246.7842, 244.6623, 245.5289, 
    243.3905,
  257.5174, 257.5992, 255.641, 253.2682, 249.5562, 251.5857, 253.0532, 
    251.5852, 250.9596, 248.8249, 246.5643, 249.1901, 249.6812, 245.9623, 
    241.456,
  263.9174, 262.5746, 261.7383, 259.423, 251.7274, 248.2406, 255.1562, 
    253.3063, 252.0019, 250.3203, 250.2546, 250.5388, 250.6511, 251.1246, 
    247.0174,
  269.1427, 265.8322, 264.8964, 263.8657, 259.464, 254.7554, 250.4061, 
    254.7505, 254.4092, 252.6575, 251.3674, 251.3532, 251.6656, 252.7154, 
    249.1906,
  272.7073, 269.0832, 266.9424, 266.2973, 263.559, 261.4281, 258.7791, 
    250.2728, 250.6438, 255.094, 254.9889, 253.9179, 252.7715, 254.0808, 
    252.1056,
  272.4389, 270.9568, 268.7537, 268.1843, 266.4459, 265.133, 263.8551, 
    261.8457, 257.5115, 256.3677, 255.5808, 255.7772, 254.6835, 254.9926, 
    253.0106,
  272.8619, 271.4088, 269.5767, 269.102, 268.0033, 267.1311, 266.3147, 
    265.7324, 264.566, 260.7626, 258.2795, 256.9275, 255.8395, 255.8706, 
    252.5907,
  273.059, 272.4354, 271.1997, 270.5976, 269.7689, 269.3698, 268.5338, 
    267.6062, 267.0265, 263.8188, 260.8142, 258.7465, 256.9585, 255.8303, 
    252.0087,
  270.5561, 271.1409, 271.1126, 270.5932, 270.0966, 269.9601, 270.3142, 
    270.0979, 269.3068, 266.6734, 263.1512, 260.3868, 257.6914, 255.9008, 
    248.922,
  268.4809, 267.7795, 267.4077, 267.5069, 267.4533, 267.0973, 267.3674, 
    268.9953, 269.9175, 268.8475, 265.3886, 262.1211, 258.6325, 255.4803, 
    249.2142,
  254.9344, 255.4674, 254.2969, 255.5628, 253.6789, 253.4601, 255.4815, 
    251.429, 249.8419, 244.9745, 244.3768, 244.2875, 239.485, 239.4465, 
    235.0734,
  257.4767, 258.2437, 256.8203, 255.8839, 252.4035, 255.1025, 255.5468, 
    251.8493, 251.1106, 248.9291, 246.3724, 248.903, 247.4267, 237.882, 
    233.8557,
  262.2518, 261.9927, 260.9042, 258.5446, 254.5374, 251.2881, 256.148, 
    252.7515, 251.8245, 250.7208, 251.1598, 249.892, 248.1163, 245.7767, 
    238.585,
  265.0984, 264.7672, 263.8337, 262.3599, 259.8007, 257.2198, 250.8872, 
    253.4176, 253.0147, 251.4319, 251.301, 250.4667, 249.1244, 247.8438, 
    242.459,
  267.2321, 266.6828, 265.7492, 264.6064, 262.9363, 262.2989, 259.2452, 
    248.973, 248.5843, 252.4363, 252.7126, 252.2426, 250.5325, 250.536, 
    248.2404,
  268.946, 267.9343, 267.0714, 266.3399, 264.8366, 264.5852, 263.7196, 
    260.8985, 256.461, 254.075, 253.8697, 254.1859, 252.1376, 251.5852, 
    249.5818,
  270.2735, 269.6514, 268.502, 267.7086, 266.5656, 266.2188, 265.7389, 
    264.887, 263.1118, 258.4178, 256.331, 255.3684, 253.4958, 252.5137, 
    250.7727,
  271.174, 270.1313, 269.2571, 268.647, 267.6208, 267.3024, 266.8573, 
    266.4341, 265.5904, 260.8087, 257.2965, 255.839, 254.5372, 252.7431, 
    250.6457,
  271.3635, 271.0718, 270.4024, 269.4578, 268.4909, 268.0689, 267.7899, 
    267.3475, 266.6758, 262.635, 258.4158, 257.0247, 255.2808, 252.9227, 
    249.4806,
  269.1846, 269.3809, 269.754, 269.5374, 268.945, 268.5482, 267.9033, 
    267.4524, 266.4843, 262.421, 260.3568, 258.337, 256.2558, 253.6362, 
    250.1978,
  254.7403, 256.09, 255.5772, 255.7057, 252.4061, 251.9036, 253.115, 
    248.4167, 247.4482, 241.5884, 240.4483, 241.6776, 239.4111, 239.6681, 
    237.0863,
  258.1314, 259.1637, 258.3538, 255.2431, 251.9299, 253.1212, 251.9077, 
    249.437, 248.9967, 246.9587, 244.2095, 247.5394, 246.2874, 236.9948, 
    235.4777,
  262.5245, 262.2864, 261.1275, 257.248, 254.3362, 248.1296, 251.695, 
    250.4918, 250.3695, 249.8784, 250.104, 247.5501, 246.5494, 245.3616, 
    239.4452,
  265.2258, 264.9855, 264.0801, 262.1003, 260.1199, 255.2475, 246.7024, 
    250.744, 250.8323, 249.8261, 249.3103, 247.6398, 246.9012, 246.2508, 
    244.5141,
  266.899, 266.5443, 265.7835, 264.6136, 263.4546, 260.8606, 257.2317, 
    246.5622, 245.0766, 247.7517, 250.4103, 249.4973, 248.3804, 248.611, 
    248.5164,
  268.4202, 267.91, 267.1288, 266.2944, 265.42, 264.0065, 262.6815, 260.3487, 
    256.1042, 252.6789, 250.892, 252.2068, 249.9002, 249.3161, 248.1465,
  269.4828, 269.0039, 268.1921, 267.4134, 266.8228, 265.7867, 265.0719, 
    264.053, 262.1282, 258.5424, 256.2073, 253.9738, 251.6148, 250.4508, 
    248.7678,
  270.6628, 270.0765, 269.1769, 268.4723, 267.7883, 267.1627, 266.3921, 
    265.7415, 264.1909, 259.8369, 256.3274, 254.0934, 252.5564, 250.6302, 
    248.6828,
  271.1619, 270.6148, 269.8683, 269.1507, 268.5896, 267.9727, 267.3014, 
    266.858, 265.6673, 260.3665, 256.588, 255.0572, 253.5659, 251.2, 248.721,
  271.8706, 271.2625, 270.4525, 269.6755, 269.0349, 268.4794, 267.909, 
    267.3435, 264.4676, 259.0315, 258.296, 256.4433, 254.4872, 252.5456, 
    250.4972,
  254.1245, 254.6193, 253.5227, 252.9894, 249.8337, 249.0968, 250.4192, 
    248.6225, 249.493, 244.8709, 244.2537, 246.1366, 242.9227, 241.3076, 
    238.1742,
  257.8153, 257.602, 256.1628, 252.0901, 248.9701, 248.645, 249.6064, 
    249.1868, 249.7213, 250.0027, 246.9811, 249.3849, 248.9714, 240.4497, 
    238.6157,
  261.569, 260.212, 258.473, 253.5618, 251.6279, 244.3641, 249.5987, 
    250.3243, 250.4349, 250.1739, 250.3155, 249.3473, 249.4753, 248.6732, 
    243.1879,
  264.1302, 263.0695, 261.4289, 258.7092, 257.3309, 252.5994, 244.9445, 
    249.8006, 250.3266, 249.4082, 249.3573, 249.2446, 249.5824, 249.9085, 
    248.59,
  265.611, 264.5825, 263.4147, 262.2108, 261.0655, 258.7325, 256.7459, 
    244.6779, 242.611, 246.7544, 250.583, 250.8709, 250.2733, 250.8632, 
    251.7422,
  266.6496, 265.8312, 264.8943, 264.1785, 263.2554, 261.918, 261.2184, 
    259.6088, 254.6148, 252.0993, 250.4324, 252.3071, 251.0279, 250.8435, 
    251.2571,
  267.4627, 267.0146, 266.1665, 265.5194, 264.8748, 264.1985, 263.6572, 
    262.4313, 260.4793, 257.3338, 254.6197, 252.995, 252.0955, 251.2728, 
    251.006,
  268.5669, 268.0163, 267.0552, 266.6213, 266.06, 265.7644, 265.1773, 
    263.6754, 261.3614, 257.1083, 254.3146, 253.2361, 252.9159, 251.2585, 
    251.4207,
  269.1378, 268.5876, 267.9807, 267.4522, 266.9922, 266.5119, 265.7486, 
    264.5628, 262.2381, 256.42, 254.8884, 254.7053, 254.2031, 252.4397, 
    251.8086,
  269.9203, 269.3222, 268.704, 268.1318, 267.5829, 267.0384, 266.1143, 
    264.6069, 259.317, 252.7294, 255.1218, 256.0401, 255.2269, 253.9685, 
    252.9035,
  253.4429, 254.4542, 252.8337, 253.3812, 250.4828, 249.5889, 251.334, 
    250.0262, 250.1194, 244.1068, 242.3596, 243.2862, 241.8342, 241.9851, 
    239.2046,
  258.4196, 257.7101, 256.5602, 252.8265, 248.7693, 248.3273, 251.0332, 
    251.0813, 251.2445, 251.3772, 248.2155, 250.5647, 250.4594, 243.7441, 
    242.5945,
  262.0973, 260.1934, 259.041, 254.9648, 253.5465, 243.8292, 250.7801, 
    252.1271, 252.5719, 252.5678, 252.7514, 252.7178, 253.2208, 253.0051, 
    248.8503,
  264.6978, 263.4819, 262.6506, 260.6115, 260.2642, 255.4448, 244.1148, 
    252.2472, 253.2645, 253.069, 253.1514, 253.6952, 254.2885, 254.9311, 
    253.737,
  266.1619, 265.3094, 264.7766, 264.121, 263.7684, 262.3981, 260.6048, 
    246.1054, 247.3247, 253.0687, 254.219, 255.0503, 255.0486, 256.077, 
    256.6451,
  267.4742, 266.7286, 266.2148, 265.792, 265.6368, 264.6534, 263.8437, 
    261.4801, 257.3014, 255.7974, 254.0365, 255.548, 256.0728, 256.5729, 
    257.8781,
  268.3125, 267.7153, 267.2033, 266.9404, 266.6558, 266.2046, 265.3845, 
    263.6989, 261.4302, 257.9686, 256.1897, 255.5868, 255.9387, 256.55, 
    257.7249,
  269.2293, 268.6713, 268.0364, 267.5834, 267.2339, 266.5397, 265.6033, 
    264.2739, 261.1514, 257.7209, 256.3498, 255.5093, 255.3744, 255.7063, 
    257.0988,
  269.5367, 269.1429, 268.6187, 268.1179, 267.4401, 266.8471, 265.7998, 
    264.5761, 262.4322, 258.3467, 257.8693, 256.3998, 255.0111, 255.2461, 
    255.8835,
  270.1047, 269.6962, 269.057, 268.3976, 267.6778, 266.7005, 265.2241, 
    263.862, 259.543, 256.6582, 259.0646, 256.998, 254.9604, 254.434, 255.4191,
  253.0482, 255.2662, 252.1839, 252.942, 249.9681, 248.251, 249.1833, 
    248.3802, 247.9729, 241.6935, 241.2899, 243.6366, 242.9558, 244.1236, 
    241.8619,
  258.7006, 257.426, 255.4464, 252.8099, 248.7758, 247.9607, 251.0197, 
    250.3673, 249.9715, 248.6348, 245.2622, 249.1803, 249.8341, 242.1981, 
    240.1861,
  262.6014, 260.0507, 259.1484, 255.0994, 253.3533, 243.1097, 252.0102, 
    253.4194, 253.2091, 252.6755, 251.6771, 251.6931, 251.5986, 250.5896, 
    245.1759,
  265.3433, 264.1152, 263.561, 261.0372, 260.5608, 256.4655, 247.1589, 
    253.9081, 255.1055, 254.2005, 252.9647, 252.607, 252.5278, 252.4861, 
    249.2013,
  266.8533, 266.8441, 266.9091, 266.403, 265.3268, 263.1397, 260.678, 
    249.9527, 249.9547, 253.0877, 254.4801, 253.8027, 253.8856, 254.5889, 
    252.5216,
  268.3339, 268.4125, 268.4491, 268.4327, 267.7057, 266.4685, 264.6215, 
    261.8528, 259.2495, 256.9516, 254.7615, 256.2589, 255.7073, 254.9045, 
    253.8125,
  269.3713, 269.511, 269.2607, 268.856, 268.3183, 267.6891, 266.2446, 
    264.3118, 261.7804, 260.1038, 258.9518, 257.4735, 256.6402, 255.3241, 
    254.6093,
  270.2344, 269.9422, 269.3459, 268.8485, 268.0868, 267.3398, 265.9603, 
    264.1264, 261.0452, 259.9779, 259.418, 259.1617, 258.7077, 259.0002, 
    259.5789,
  270.6172, 270.2419, 269.5312, 268.7218, 267.8791, 267.0808, 265.7959, 
    263.9706, 261.3953, 259.8116, 259.4912, 259.3142, 258.6062, 257.7733, 
    256.7182,
  270.8839, 270.1913, 269.2031, 268.2498, 267.2755, 266.2671, 265.0345, 
    263.4804, 260.526, 258.9443, 258.612, 257.202, 256.8262, 256.3876, 
    256.4753,
  251.0935, 252.4892, 250.4183, 251.8904, 249.4217, 249.0215, 252.0478, 
    252.7473, 253.5793, 251.2714, 250.7846, 250.5393, 247.6704, 246.928, 
    243.3438,
  256.6962, 255.6113, 253.7245, 252.1179, 247.9935, 247.8488, 252.0989, 
    252.9522, 253.7437, 254.3497, 252.4441, 253.5788, 252.2697, 245.7241, 
    243.6249,
  261.1811, 258.9503, 257.4614, 253.5274, 251.3763, 243.5003, 251.3697, 
    253.087, 253.9165, 254.4773, 254.4906, 253.9734, 253.6972, 251.0991, 
    247.3427,
  264.5677, 262.4405, 261.4731, 258.2936, 257.7713, 253.913, 245.099, 
    251.4995, 253.2869, 253.3873, 253.557, 253.4732, 253.3115, 251.7705, 
    249.6481,
  266.7997, 265.6086, 264.6387, 262.6565, 262.2184, 260.2084, 258.4059, 
    246.2201, 244.9203, 251.2249, 254.1654, 254.4901, 254.487, 253.9958, 
    252.888,
  268.6561, 267.6961, 267.077, 265.8823, 265.4427, 263.3938, 262.1805, 
    259.9344, 257.3104, 255.1075, 253.9393, 255.8009, 255.4221, 254.625, 
    254.1677,
  270.1436, 269.9218, 268.9554, 267.8259, 267.3945, 266.2346, 265.0676, 
    263.1734, 260.8587, 257.7953, 257.077, 256.022, 255.3651, 254.1293, 
    254.0837,
  271.4292, 270.8195, 270.0245, 269.1058, 268.4963, 267.4186, 266.4632, 
    264.6848, 260.5805, 258.3085, 257.466, 256.7656, 256.7768, 255.9604, 
    254.9748,
  271.742, 271.1148, 270.5552, 269.6984, 269.0514, 268.0428, 267.1401, 
    264.7419, 260.9783, 259.3988, 258.9554, 258.738, 257.1929, 254.7893, 
    252.934,
  271.5043, 270.6198, 269.9792, 269.2568, 268.734, 267.6567, 266.4417, 
    264.3575, 260.8306, 259.6736, 259.9026, 258.4732, 255.2982, 253.8892, 
    253.6462,
  248.7666, 252.1441, 249.1589, 252.8328, 249.4505, 250.8002, 255.2465, 
    254.585, 253.0387, 248.6657, 248.6528, 247.2599, 243.8844, 242.1261, 
    239.1706,
  254.3926, 255.3076, 254.926, 253.6489, 247.2904, 249.7479, 255.7767, 
    255.3511, 254.3897, 252.8007, 248.28, 249.5623, 247.403, 241.3979, 
    241.6279,
  260.1533, 259.2884, 259.0645, 256.576, 255.1331, 249.4233, 255.5211, 
    256.2871, 255.5168, 253.7734, 251.9441, 250.9094, 249.809, 248.2706, 
    245.1266,
  263.6346, 263.1014, 262.9057, 261.2315, 259.9736, 257.0423, 250.1331, 
    254.2728, 253.3745, 252.7642, 251.4056, 250.3537, 249.7231, 249.1974, 
    248.8335,
  265.8798, 265.4927, 265.2992, 265.0987, 264.192, 261.397, 259.1819, 
    248.1339, 246.8125, 250.2838, 251.3067, 250.4062, 250.4376, 250.8833, 
    251.1537,
  267.3501, 266.6562, 266.6279, 266.7164, 266.2637, 264.1418, 262.6386, 
    259.7623, 257.0219, 254.0663, 251.4473, 251.4547, 251.28, 251.5351, 
    251.8776,
  268.6952, 268.0078, 267.792, 267.7439, 267.4499, 266.1938, 264.6582, 
    262.4021, 259.7284, 255.6936, 253.6077, 252.3732, 251.9551, 251.6558, 
    252.0491,
  270.0186, 269.061, 268.316, 268.1641, 267.8401, 266.9155, 265.9635, 
    264.2564, 259.5103, 256.262, 254.0733, 253.0837, 252.4279, 251.9311, 
    252.1834,
  270.9118, 270.0594, 269.2278, 268.6221, 268.0793, 267.434, 266.4455, 
    263.7827, 259.1767, 256.3512, 254.6617, 253.6852, 252.4753, 251.8957, 
    251.8991,
  271.7854, 270.9714, 269.9166, 269.0598, 268.4617, 267.4078, 266.0602, 
    263.1773, 258.2383, 256.6402, 255.4324, 254.2293, 252.8123, 252.4672, 
    252.5443,
  247.7522, 252.6288, 249.3089, 253.8739, 252.6243, 252.8434, 254.7493, 
    253.0042, 251.6352, 246.8546, 245.5932, 245.1327, 243.2722, 241.9044, 
    238.8201,
  254.6161, 255.7615, 256.0773, 254.7797, 248.7077, 250.7053, 253.7364, 
    252.3443, 251.394, 249.5687, 247.5774, 248.3365, 247.7011, 240.7431, 
    239.642,
  260.8919, 260.2257, 260.3538, 258.7361, 253.3071, 244.8758, 251.937, 
    252.3296, 252.0711, 251.8296, 251.177, 249.9775, 249.6373, 247.9999, 
    243.7921,
  264.1709, 264.1699, 264.2807, 263.6304, 261.9274, 256.4068, 245.2068, 
    249.9616, 251.4307, 251.6515, 250.7878, 249.0834, 249.0586, 248.196, 
    247.3888,
  265.8847, 266.3324, 266.5786, 266.7083, 266.0818, 262.7855, 258.2549, 
    243.871, 242.8467, 248.2458, 249.9115, 248.967, 249.2077, 249.7059, 
    250.5128,
  266.8521, 267.7565, 268.0204, 268.0861, 267.8755, 266.0082, 262.7077, 
    258.3098, 254.2723, 251.7088, 249.4872, 249.5425, 249.6523, 250.2703, 
    250.9584,
  267.7892, 268.7429, 269.1784, 269.0957, 268.8632, 267.874, 265.5093, 
    261.5191, 256.9249, 253.0281, 251.4347, 250.3775, 250.2348, 250.4322, 
    251.1641,
  268.8499, 269.6081, 269.7186, 269.701, 269.4053, 268.6261, 266.8578, 
    264.2294, 258.0613, 253.4086, 251.6816, 250.921, 250.7029, 250.4111, 
    251.0148,
  269.6824, 270.1542, 270.4039, 270.0943, 269.774, 268.9867, 267.8395, 
    265.6327, 258.4047, 253.0019, 251.5632, 251.3284, 250.8876, 250.4705, 
    250.9488,
  270.6019, 270.5483, 270.1774, 269.6782, 269.4431, 268.5459, 267.7056, 
    265.8274, 257.7309, 252.9315, 252.5228, 252.0021, 251.455, 251.2631, 
    251.6939,
  249.5589, 253.0275, 250.87, 255.6792, 253.3538, 251.9492, 252.1326, 
    249.4244, 245.9809, 240.0936, 240.2738, 243.5079, 243.2372, 240.6642, 
    236.9258,
  254.2885, 255.0474, 256.4373, 256.8326, 250.411, 248.6176, 251.5943, 
    250.5772, 248.0564, 245.9588, 242.4038, 246.9072, 248.7713, 239.1631, 
    236.5905,
  260.4038, 260.1696, 260.7216, 259.7815, 256.3128, 245.1972, 249.1736, 
    250.7993, 249.386, 248.5661, 247.2188, 248.9117, 250.6378, 247.9492, 
    242.4419,
  264.1982, 264.0781, 264.45, 264.4139, 263.9019, 258.2065, 243.5099, 
    249.2152, 250.887, 250.0584, 248.1687, 248.1076, 249.5461, 249.2599, 
    245.6069,
  265.9767, 266.0494, 266.3659, 266.6915, 267.6678, 266.5732, 258.4681, 
    243.6673, 243.3442, 249.4624, 248.4733, 247.8976, 248.8995, 249.4675, 
    248.8259,
  266.7506, 267.1673, 267.5213, 267.7704, 268.3687, 268.838, 265.4965, 
    257.9388, 254.2538, 253.4061, 250.0195, 248.6169, 248.6625, 248.9428, 
    248.9585,
  267.4393, 267.9624, 268.2475, 268.45, 268.8743, 269.3095, 268.9406, 
    264.115, 259.1467, 255.8515, 252.7509, 249.4457, 248.9096, 248.7142, 
    249.0221,
  268.194, 268.6089, 268.877, 269.0787, 269.3059, 269.5285, 269.4123, 
    267.4668, 261.7386, 256.3394, 253.0589, 250.2036, 249.131, 248.5925, 
    248.8305,
  268.6022, 268.864, 269.2724, 269.4917, 269.6496, 269.7258, 269.7005, 
    268.1786, 261.4572, 255.411, 252.9572, 251.0186, 249.5121, 248.6308, 
    248.9701,
  269.1863, 269.3643, 269.6765, 269.7433, 269.8038, 269.291, 269.0117, 
    267.7009, 260.5249, 255.5973, 254.0868, 251.7621, 250.2227, 249.5518, 
    249.3616,
  253.3038, 252.8749, 251.3058, 253.1404, 252.5593, 248.9452, 246.7713, 
    247.3382, 245.3347, 238.6775, 239.2395, 241.7776, 240.0576, 238.5325, 
    234.9197,
  255.7251, 255.1571, 254.3794, 254.6564, 251.4566, 247.4901, 247.7245, 
    247.4369, 245.8929, 244.2708, 241.9967, 247.3556, 247.4468, 237.02, 
    234.5432,
  260.4554, 259.0342, 257.3635, 256.159, 252.9043, 243.5659, 247.2493, 
    247.5746, 246.6809, 247.3325, 247.3446, 249.7501, 250.7338, 246.8859, 
    241.3292,
  265.2589, 263.3406, 262.0751, 260.0443, 257.2137, 251.5026, 242.551, 
    246.201, 246.8557, 247.1744, 247.2, 249.0443, 251.6058, 249.0213, 244.6355,
  267.5256, 266.0771, 264.6008, 263.4127, 262.1027, 259.1297, 254.7203, 
    242.2355, 240.8953, 245.8985, 247.1074, 247.9634, 250.9881, 251.5793, 
    247.7372,
  268.5226, 267.8467, 266.5658, 265.2754, 264.5308, 263.3882, 261.2917, 
    256.763, 253.4693, 252.3499, 249.2209, 248.5616, 249.2282, 250.4991, 
    249.0576,
  269.2393, 269.0182, 267.8823, 266.6476, 266.0925, 265.4129, 264.9167, 
    262.7869, 260.1039, 256.6119, 252.7437, 249.4846, 249.1381, 249.6609, 
    249.1102,
  269.9039, 269.8633, 269.0954, 267.808, 267.1943, 266.7863, 266.5753, 
    266.1575, 264.067, 260.3564, 254.7683, 250.3946, 249.2236, 248.8291, 
    248.4567,
  270.2861, 270.2515, 269.6826, 268.6949, 267.992, 267.4976, 267.3686, 
    267.136, 264.1254, 261.5165, 258.4165, 253.7622, 250.1417, 248.4814, 
    248.0072,
  270.6791, 270.7314, 270.3304, 269.2112, 268.4643, 267.6906, 267.3094, 
    266.5975, 263.081, 260.8634, 260.6632, 257.7524, 253.9977, 250.6404, 
    248.5979,
  262.8506, 260.7293, 255.2831, 251.2219, 248.5856, 246.429, 246.3678, 
    247.6643, 246.3354, 239.0907, 238.7567, 238.905, 236.8127, 237.3087, 
    233.5581,
  265.1185, 262.3278, 257.9655, 252.5137, 248.0857, 245.7247, 246.8578, 
    247.4984, 247.0571, 244.2973, 241.3474, 244.2233, 243.6461, 235.6686, 
    233.5406,
  268.7076, 265.6897, 259.8381, 253.8433, 249.6451, 242.6891, 246.3418, 
    247.339, 247.2149, 247.2912, 246.8532, 247.3079, 246.7662, 244.4435, 
    240.2677,
  270.9497, 269.2826, 264.3149, 257.5515, 253.3627, 249.6044, 242.0874, 
    245.406, 246.6623, 247.2984, 247.4218, 248.0654, 248.1626, 246.4025, 
    243.1051,
  271.9689, 271.0374, 267.3251, 262.2997, 258.8472, 255.7892, 252.7451, 
    241.732, 240.7302, 245.3395, 247.3204, 248.3491, 248.8299, 248.3486, 
    246.1557,
  272.3784, 271.822, 269.3277, 265.0997, 262.2574, 260.3826, 258.0993, 
    254.973, 252.0629, 250.8953, 248.4393, 249.1571, 248.9574, 248.8275, 
    247.1789,
  272.7544, 272.252, 270.6891, 267.0162, 264.5328, 262.775, 261.6405, 
    258.9583, 256.376, 254.6493, 251.856, 249.6997, 249.3443, 248.9105, 
    247.8364,
  272.7711, 272.397, 271.4491, 268.497, 266.0243, 264.7951, 263.6979, 
    262.3078, 259.3281, 255.629, 252.5704, 250.0974, 249.5615, 248.668, 
    247.8902,
  272.3517, 272.1354, 271.9764, 269.5377, 267.4437, 265.821, 264.8022, 
    263.8055, 259.795, 255.822, 253.5046, 250.9439, 249.7071, 248.4601, 
    247.3718,
  271.7225, 271.7291, 271.8998, 270.2086, 268.046, 266.5836, 265.3748, 
    263.6705, 258.6762, 256.0919, 256.0753, 253.8184, 251.4563, 249.3598, 
    247.9033,
  264.0908, 266.0256, 265.5446, 260.6745, 254.0777, 249.0366, 248.6367, 
    248.1364, 244.3559, 237.2431, 237.1096, 236.7274, 234.9033, 235.4747, 
    233.1305,
  267.194, 268.2869, 267.076, 259.4436, 250.2189, 247.9662, 247.9467, 
    247.4494, 244.8632, 241.853, 239.3235, 241.3936, 240.3664, 233.8186, 
    232.241,
  269.9052, 269.934, 267.6149, 259.0541, 251.0231, 243.5362, 246.8871, 
    247.1824, 245.8928, 244.6366, 243.5319, 243.3756, 242.9451, 240.9717, 
    237.7097,
  271.3913, 272.0094, 270.1413, 261.4544, 254.7928, 250.4687, 242.11, 
    245.2688, 245.6936, 245.4894, 244.6221, 244.3771, 243.866, 242.5895, 
    240.796,
  271.8747, 272.2094, 271.4749, 265.7189, 259.3149, 255.7658, 252.1641, 
    240.5631, 238.9321, 243.6122, 244.676, 244.9338, 244.854, 244.2449, 
    243.7457,
  272.3105, 272.5349, 272.2054, 268.2236, 263.4376, 260.5667, 257.1634, 
    253.3607, 250.335, 248.9644, 246.1911, 246.1543, 245.6829, 245.3167, 
    244.6875,
  273.0097, 272.8757, 272.5512, 269.7962, 265.8564, 262.9125, 260.6111, 
    256.6427, 253.5599, 251.93, 249.1574, 247.2543, 246.608, 245.9211, 
    245.4841,
  272.8454, 272.3759, 272.3437, 270.6349, 267.0033, 264.8642, 262.8369, 
    259.7956, 256.1306, 252.7605, 250.0253, 247.9375, 247.3421, 246.5696, 
    246.1283,
  272.0919, 271.9382, 272.2977, 271.197, 267.9807, 265.4604, 263.8752, 
    262.3001, 256.5533, 252.2042, 250.1159, 248.7482, 248.0546, 246.8721, 
    245.9734,
  271.3104, 271.2877, 272.0851, 271.0394, 268.0495, 266.2811, 264.5119, 
    261.6613, 254.5181, 251.8149, 251.3182, 249.5982, 248.9935, 247.8557, 
    246.3559,
  262.6943, 263.219, 263.269, 263.6774, 261.7937, 257.809, 255.0205, 
    251.7626, 245.5509, 238.5603, 238.2284, 237.553, 235.2973, 235.5883, 
    233.2229,
  264.3852, 264.029, 263.9565, 263.9624, 260.0817, 255.0389, 252.9187, 
    249.8412, 245.757, 242.5975, 240.0458, 241.8068, 241.0598, 233.0741, 
    231.148,
  267.9749, 267.4307, 266.1333, 264.7356, 260.1091, 249.9319, 249.6497, 
    248.8352, 245.9158, 244.8136, 243.6986, 243.9942, 243.3327, 241.0636, 
    237.0025,
  269.7502, 269.7085, 269.3058, 267.3139, 262.3618, 255.0402, 244.9186, 
    245.2025, 245.3096, 244.8907, 244.8699, 244.1803, 243.2949, 241.8459, 
    239.6696,
  271.1783, 270.9205, 270.6189, 269.8372, 265.0799, 259.1804, 254.5368, 
    241.5834, 239.2346, 243.0664, 244.5132, 244.2572, 243.5501, 242.7469, 
    242.0813,
  271.5493, 271.4496, 271.2005, 270.8562, 267.8687, 263.5054, 259.5598, 
    255.1103, 250.4961, 247.7468, 245.3516, 244.9105, 244.0473, 242.8981, 
    242.4616,
  272.0428, 271.817, 271.5953, 271.2714, 269.1326, 265.6458, 263.0309, 
    257.6094, 253.0777, 251.0774, 248.4146, 245.5898, 244.4886, 243.1666, 
    242.7457,
  272.4411, 271.9314, 271.7233, 271.3942, 269.2945, 266.7482, 263.9439, 
    259.4122, 254.4364, 250.6548, 248.0518, 245.7675, 244.7203, 243.3678, 
    243.115,
  272.1861, 272.0602, 271.908, 271.3399, 269.2112, 266.7495, 264.3022, 
    260.5367, 253.3694, 249.2602, 247.1347, 245.7195, 244.8493, 243.6804, 
    243.1679,
  271.7621, 271.6933, 271.6472, 270.8184, 268.6271, 266.4592, 263.4646, 
    257.7635, 249.9064, 248.2134, 247.6281, 246.0576, 245.5406, 244.5406, 
    244.0675,
  263.9433, 263.9797, 263.4465, 262.872, 262.0839, 261.087, 261.1264, 
    259.0579, 255.1249, 247.2821, 243.3532, 241.0384, 236.5639, 236.1323, 
    236.0284,
  266.5383, 265.4626, 264.4411, 263.6589, 262.1114, 260.9287, 260.1535, 
    257.7693, 254.0765, 248.8649, 244.6369, 244.442, 242.765, 234.1708, 
    233.6745,
  269.6002, 268.7456, 266.9421, 264.2925, 262.357, 257.0748, 257.4047, 
    255.9693, 252.2849, 249.379, 246.9353, 246.9132, 245.6122, 243.0478, 
    238.6829,
  271.2154, 270.9353, 270.1024, 267.1462, 264.3262, 261.0269, 250.2625, 
    249.642, 249.2413, 248.5394, 247.4376, 246.3742, 245.5495, 243.6108, 
    241.1098,
  272.5965, 272.0525, 271.2972, 269.5035, 265.9091, 262.9956, 257.8077, 
    244.7673, 242.6931, 245.8563, 246.502, 245.9575, 245.3058, 244.5157, 
    243.9864,
  273.2101, 272.7924, 271.9736, 270.2732, 267.6766, 265.0334, 262.0503, 
    257.6155, 253.724, 249.6355, 247.4733, 246.6304, 245.4088, 244.0847, 
    243.2529,
  273.2088, 272.8108, 272.2313, 270.5924, 268.2931, 266.3731, 263.9543, 
    260.4995, 257.5767, 253.6283, 250.5345, 246.8029, 245.3902, 243.3642, 
    242.8346,
  273.1067, 272.4241, 271.9639, 270.3419, 268.7574, 267.2696, 265.2564, 
    262.2634, 257.1655, 252.356, 249.6232, 246.5509, 245.1401, 242.8985, 
    242.353,
  273.1272, 272.5693, 271.7251, 270.2223, 268.8835, 267.4633, 265.8453, 
    262.2762, 254.0511, 249.8001, 247.4679, 245.9617, 244.2845, 242.6801, 
    241.938,
  271.612, 271.4201, 270.8608, 269.6561, 268.6541, 267.0518, 263.7503, 
    255.349, 249.1012, 248.0319, 247.8472, 245.8316, 244.5699, 243.4969, 
    243.2263,
  262.0768, 262.3657, 261.7885, 261.3797, 260.4338, 259.0156, 259.3637, 
    259.0531, 258.7426, 254.1198, 252.6363, 251.6151, 247.6525, 245.904, 
    244.2554,
  266.6063, 264.5942, 263.2912, 262.1343, 260.6281, 259.7449, 259.7573, 
    258.925, 258.4021, 257.6325, 254.6977, 254.3565, 250.8188, 242.853, 
    240.9643,
  270.9912, 269.8725, 267.9634, 265.0829, 262.4236, 257.8489, 259.1364, 
    258.527, 257.0845, 256.8485, 256.0024, 254.3657, 251.0688, 246.7144, 
    242.8006,
  272.634, 272.3821, 271.8617, 270.1521, 266.4357, 262.9402, 254.5467, 
    254.7783, 254.2933, 254.6861, 254.4503, 252.8819, 250.03, 246.216, 
    242.6128,
  273.037, 272.7084, 272.415, 272.2636, 269.8649, 266.9171, 262.4595, 
    252.857, 250.7311, 250.9811, 252.2121, 251.3832, 248.6583, 246.2213, 
    243.8356,
  272.8491, 272.6157, 272.4357, 272.2721, 271.3037, 268.6798, 265.0471, 
    261.5623, 257.974, 255.1628, 252.3789, 250.3786, 247.8277, 245.3663, 
    243.6246,
  272.3712, 272.1456, 272.0665, 271.69, 270.4877, 268.0754, 264.9841, 261.19, 
    258.7518, 256.8864, 253.877, 249.6925, 246.9461, 244.5755, 243.1186,
  271.6371, 270.895, 270.2167, 269.6552, 268.1902, 266.6759, 264.3876, 
    261.5752, 257.3368, 254.8596, 252.2554, 248.2216, 246.4926, 243.5347, 
    242.7614,
  271.2688, 270.4009, 269.6069, 268.5495, 267.6044, 266.0104, 264.1707, 
    260.8277, 253.8954, 250.9166, 248.9621, 247.2774, 245.0467, 243.2713, 
    242.8738,
  270.0797, 269.8926, 269.1741, 268.3717, 267.176, 265.5191, 262.3956, 
    255.4685, 249.6524, 248.3647, 248.6135, 246.3965, 245.4091, 244.0467, 
    244.7596,
  263.1688, 263.8552, 262.6599, 261.2572, 259.4884, 255.7898, 255.8235, 
    254.8477, 253.6488, 246.9433, 246.9718, 248.7368, 246.9221, 246.8111, 
    245.5369,
  270.049, 268.9383, 267.3722, 265.0991, 261.5718, 258.8812, 257.5257, 
    255.2363, 254.0636, 252.026, 249.877, 251.9254, 251.5361, 246.0267, 
    244.7982,
  271.9753, 271.3306, 270.3013, 268.6072, 264.6819, 258.6422, 259.2517, 
    257.7192, 255.5658, 254.1712, 253.504, 253.8794, 253.6952, 251.8714, 
    247.7131,
  271.917, 271.7359, 271.6392, 271.2179, 268.5466, 263.5566, 257.0865, 
    256.4355, 255.5629, 255.37, 254.6697, 254.4375, 253.9999, 252.5814, 
    248.3469,
  271.6361, 271.1617, 271.0895, 271.2979, 270.7111, 267.8721, 262.9848, 
    254.2943, 251.8688, 255.1587, 254.8647, 254.6672, 254.0693, 252.6416, 
    249.7301,
  271.3321, 270.7871, 270.5542, 270.4985, 270.6104, 269.2771, 265.9247, 
    264.2054, 262.0387, 259.5934, 256.5626, 255.6221, 254.351, 251.4271, 
    248.5783,
  270.9744, 270.2658, 269.5756, 269.0033, 268.6492, 268.1222, 265.8779, 
    263.8411, 262.2361, 261.8429, 258.6653, 255.9306, 253.341, 249.6524, 
    247.3386,
  270.7769, 269.796, 268.8402, 267.9633, 267.0182, 265.9464, 264.4284, 
    262.2042, 259.2235, 258.8704, 256.753, 254.2254, 251.6826, 248.0985, 
    246.2101,
  270.5775, 269.3307, 268.2115, 267.0828, 265.9168, 264.3157, 262.4613, 
    259.286, 253.994, 253.8556, 253.3893, 252.0091, 248.8331, 245.8068, 
    243.496,
  269.8627, 268.1393, 266.5544, 265.2901, 263.9178, 262.1487, 259.6654, 
    254.5294, 250.4778, 249.6868, 251.2534, 249.2957, 247.3788, 245.3781, 
    243.9167,
  267.7863, 268.6148, 266.6905, 267.318, 265.8895, 263.1842, 262.2788, 
    260.5118, 257.5328, 249.154, 248.7162, 250.5875, 248.6412, 248.3924, 
    247.6231,
  267.9656, 266.8387, 265.7867, 267.0241, 265.6293, 264.5129, 263.163, 
    261.1185, 259.4403, 253.818, 251.2179, 252.3497, 251.064, 245.6664, 
    245.5027,
  270.7511, 269.8711, 267.699, 265.7058, 265.6493, 262.199, 262.6397, 
    261.5227, 260.239, 257.9617, 255.2996, 254.1671, 252.1956, 249.6303, 
    246.918,
  270.8911, 270.1711, 269.6771, 268.5713, 266.1687, 264.4556, 258.3242, 
    257.7973, 257.641, 257.1425, 255.3484, 253.3954, 252.5537, 250.823, 
    247.7772,
  271.0041, 270.015, 269.4663, 268.9843, 267.9474, 266.8616, 263.6259, 
    250.5947, 253.9746, 256.4804, 256.1917, 254.5409, 252.8965, 251.7233, 
    249.5858,
  271.1481, 270.1139, 269.5749, 268.958, 268.2763, 267.0576, 264.8261, 
    262.1749, 260.1076, 260.6525, 257.6543, 255.7665, 253.7376, 252.1065, 
    250.007,
  271.4608, 270.4962, 269.826, 269.0526, 268.2444, 266.9683, 264.944, 
    261.5182, 259.4787, 261.2557, 259.474, 255.8206, 253.9167, 252.0356, 
    249.8531,
  271.6227, 270.7175, 270.2774, 269.4042, 268.1926, 266.7885, 264.8339, 
    261.3386, 256.9551, 257.3804, 257.6481, 255.4708, 253.9159, 251.4696, 
    249.0414,
  271.7539, 271.2639, 270.7467, 269.3451, 267.7935, 266.0371, 264.4139, 
    260.3301, 254.6712, 254.3477, 256.0283, 254.7685, 253.0839, 249.5363, 
    245.5176,
  272.3646, 271.8401, 270.8658, 268.8056, 267.0063, 265.2363, 263.1993, 
    259.3886, 252.2476, 248.4972, 253.7421, 253.959, 251.8065, 247.923, 
    245.774,
  263.169, 264.5944, 258.6185, 263.0885, 261.6458, 260.9203, 262.488, 
    262.0604, 261.5646, 256.98, 255.566, 255.4101, 252.8149, 251.8595, 
    250.3383,
  264.0971, 262.4641, 261.6211, 262.3641, 260.2362, 261.2544, 262.3335, 
    261.7151, 261.5206, 259.5127, 257.239, 257.5412, 257.0135, 251.4337, 
    249.5768,
  269.268, 269.239, 267.5538, 265.5025, 262.7046, 259.5861, 262.4204, 
    262.0031, 261.4075, 259.3283, 258.2659, 258.1288, 256.6204, 254.8363, 
    251.4972,
  270.7683, 270.9543, 271.1736, 270.8842, 269.1964, 267.4284, 262.8054, 
    261.0829, 260.3354, 258.6367, 255.7572, 254.7498, 254.6185, 253.8257, 
    251.8284,
  271.7383, 271.6194, 271.6187, 271.7597, 271.5165, 271.069, 269.3174, 
    260.8564, 256.7919, 255.8666, 254.9935, 254.791, 253.8355, 254.2057, 
    252.33,
  271.826, 272.0589, 272.2297, 272.1854, 272.007, 271.4455, 269.8683, 
    267.1856, 262.1695, 258.901, 254.8387, 255.1017, 254.1907, 253.2474, 
    251.5158,
  272.2154, 272.8236, 272.8709, 272.0062, 271.7413, 270.6972, 269.26, 
    266.1579, 262.6311, 260.2815, 255.6454, 252.9385, 253.5236, 253.1454, 
    250.9677,
  273.2097, 273.5606, 272.9954, 271.548, 271.0468, 269.5872, 267.9679, 
    266.3353, 261.5033, 257.2874, 253.0029, 251.086, 253.1514, 251.9592, 
    250.1361,
  274.2391, 273.9297, 272.856, 270.8637, 270.2109, 268.1727, 266.4182, 
    264.82, 259.572, 254.7667, 251.1674, 251.3002, 251.9006, 250.2284, 247.739,
  274.311, 273.3345, 272.0373, 269.513, 268.7564, 266.7596, 264.2067, 
    262.1466, 256.6273, 250.114, 248.2784, 251.4378, 251.4658, 249.3186, 
    247.5066,
  258.6635, 261.1371, 258.2024, 261.1918, 260.9119, 260.8918, 261.8811, 
    261.7139, 261.6069, 260.4472, 260.8883, 261.617, 260.4763, 259, 254.8627,
  261.8028, 263.5138, 262.9565, 262.839, 261.9552, 262.5255, 262.541, 
    261.9367, 261.0012, 260.4373, 261.2064, 262.4939, 261.6104, 256.3985, 
    253.4859,
  269.1162, 269.8835, 269.2061, 267.3868, 264.1616, 259.7909, 262.607, 
    262.5788, 261.0064, 259.3848, 260.6182, 260.7984, 259.2096, 256.9158, 
    253.6237,
  272.0401, 272.1914, 271.8552, 270.6639, 267.6512, 262.6422, 257.5469, 
    259.6842, 259.661, 257.1188, 257.336, 257.8438, 257.4774, 256.6657, 
    254.6561,
  273.1839, 272.5248, 271.9429, 270.7081, 269.6986, 267.7358, 262.4229, 
    255.1963, 254.9776, 254.6807, 254.5922, 254.9846, 255.7494, 257.1158, 
    256.1364,
  273.9048, 273.2353, 272.2158, 270.739, 269.7886, 267.9887, 265.3049, 
    262.2473, 258.3923, 256.0755, 252.9431, 254.7074, 256.2245, 256.9616, 
    254.1185,
  274.5775, 273.8227, 272.561, 271.0849, 269.9857, 268.1706, 266.2282, 
    262.2341, 258.7585, 256.4319, 253.1278, 252.4771, 255.029, 253.9821, 
    251.414,
  274.5937, 273.8951, 272.853, 271.4782, 270.2738, 268.4314, 266.2536, 
    263.5356, 257.9089, 255.0555, 251.4453, 251.1033, 250.752, 249.8048, 
    249.2263,
  274.453, 273.8481, 273.1104, 271.7352, 270.4537, 268.2712, 266.2789, 
    263.6389, 257.7419, 253.19, 250.51, 249.3409, 248.8304, 248.2025, 247.7762,
  274.1073, 273.1954, 272.5917, 271.4049, 270.1366, 268.4052, 265.9328, 
    262.8889, 257.5339, 251.5628, 248.3076, 249.2648, 248.6117, 248.1436, 
    247.4132,
  259.2279, 261.0458, 257.6045, 258.9395, 256.8625, 257.1918, 259.3607, 
    258.0882, 255.9027, 251.3605, 253.6622, 255.9443, 253.6259, 252.4285, 
    249.7113,
  264.0531, 262.5532, 259.4736, 259.3662, 256.5844, 259.3896, 260.6067, 
    259.6576, 257.3364, 253.6494, 253.4829, 255.9784, 254.3649, 248.6358, 
    246.9582,
  268.4846, 267.2875, 266.3527, 264.8488, 261.2386, 257.5072, 263.087, 
    261.8771, 259.8969, 254.5051, 254.838, 255.8496, 254.5131, 252.0629, 
    248.4249,
  270.3838, 270.8715, 271.3845, 270.7095, 268.1674, 265.1416, 262.1192, 
    261.8771, 261.5681, 256.3747, 254.0759, 256.2333, 255.4796, 252.2247, 
    249.8582,
  271.6515, 271.928, 272.2332, 272.0981, 271.7956, 271.1044, 268.716, 
    261.8825, 260.31, 259.3718, 254.1754, 255.6068, 255.2384, 254.0168, 
    254.4482,
  272.963, 272.8867, 272.8131, 272.4956, 272.2561, 271.8759, 270.9706, 
    269.0348, 267.0274, 263.6659, 254.3812, 255.5952, 254.1544, 252.054, 
    249.8734,
  273.6179, 273.3776, 272.8464, 272.4615, 272.2842, 272.0738, 271.6223, 
    270.274, 268.6829, 266.1559, 258.4167, 253.6909, 254.4591, 249.5151, 
    247.8057,
  274.0197, 273.6103, 272.9734, 272.573, 272.3913, 272.1237, 271.4951, 
    270.8281, 269.554, 267.5014, 262.0617, 254.9142, 253.3186, 250.6224, 
    246.4803,
  274.0799, 273.4398, 272.8362, 272.4221, 272.2516, 271.2825, 271.4826, 
    270.722, 270.0869, 268.3237, 263.8764, 257.4038, 253.4553, 249.2082, 
    246.4996,
  273.6839, 273.0387, 272.2125, 271.6125, 271.08, 270.3759, 270.5194, 
    270.4666, 270.4387, 268.8354, 265.1953, 259.7311, 254.8096, 250.4771, 
    247.8623,
  260.0614, 261.8847, 263.0836, 267.2129, 266.7986, 266.9416, 267.6535, 
    264.7412, 257.2058, 246.4539, 249.5696, 251.9783, 247.6819, 244.842, 
    243.595,
  262.5533, 264.4663, 266.9095, 268.0559, 266.8942, 267.5154, 267.8645, 
    265.5784, 262.241, 252.6593, 248.2447, 253.0999, 250.866, 242.136, 
    241.0401,
  267.6944, 268.3831, 269.8945, 269.1579, 267.5816, 264.9914, 268.1428, 
    267.0281, 266.8817, 260.0077, 254.5544, 252.9232, 251.8643, 251.1447, 
    247.7076,
  269.7811, 270.8647, 271.0291, 270.5288, 269.5054, 268.2753, 265.1374, 
    264.1214, 268.1351, 265.4573, 259.2185, 254.9314, 251.271, 250.6312, 
    251.0093,
  271.137, 271.259, 271.0687, 270.8314, 270.7222, 270.6854, 269.2571, 
    264.4454, 264.8584, 267.4768, 263.0941, 259.7236, 253.5252, 251.0871, 
    252.5185,
  271.8848, 271.614, 271.3183, 271.0889, 270.9875, 270.9937, 270.6313, 
    269.4264, 268.2801, 268.5046, 265.9068, 263.3052, 258.7989, 253.4025, 
    250.8071,
  272.902, 272.4072, 271.5804, 271.5874, 271.3822, 271.4276, 271.1814, 
    270.0526, 269.3413, 268.511, 267.883, 264.7619, 261.7825, 256.3799, 
    251.639,
  273.4579, 273.2601, 272.4931, 271.8533, 271.9018, 271.7842, 271.2404, 
    270.5801, 269.6386, 268.3701, 268.1678, 265.9777, 263.6407, 259.2256, 
    253.8908,
  273.9552, 273.8623, 273.5475, 272.6309, 272.1854, 271.3867, 271.0806, 
    270.3991, 269.7718, 269.0927, 268.7469, 266.6042, 264.8795, 261.5191, 
    256.2153,
  274.2715, 273.8742, 273.2573, 272.5346, 271.9591, 271.1178, 270.0865, 
    268.6121, 269.325, 268.3856, 268.5924, 267.3635, 265.1217, 262.4358, 
    258.6502,
  265.3177, 265.9339, 265.4383, 265.568, 265.1721, 264.6693, 264.8794, 
    263.314, 260.9942, 252.1173, 247.7316, 249.0532, 242.6261, 243.2028, 
    242.539,
  266.8461, 266.914, 266.5734, 265.4836, 264.3116, 264.9651, 263.9286, 
    265.1325, 264.3637, 261.9961, 254.2427, 253.3399, 251.9021, 246.3038, 
    243.7477,
  268.7466, 268.2538, 268.246, 267.4678, 266.0223, 261.3643, 266.2375, 
    265.427, 265.2031, 264.3812, 261.8047, 259.3466, 256.6964, 254.8578, 
    250.6589,
  269.8652, 269.7325, 269.7879, 269.4975, 268.3337, 266.4284, 263.6829, 
    262.8399, 263.4169, 263.4955, 263.4392, 262.4708, 260.7839, 258.6125, 
    256.7463,
  270.683, 270.4331, 270.2536, 270.2679, 270.2077, 270.1014, 268.9068, 
    263.7361, 263.7973, 265.3405, 265.7706, 265.4061, 264.142, 261.6703, 
    259.4034,
  271.4201, 271.0062, 271.0031, 270.9836, 271.0775, 271.0338, 270.7215, 
    269.5373, 269.0359, 268.0943, 267.7149, 266.2705, 265.971, 264.6667, 
    262.2038,
  272.3861, 272.2396, 272.138, 271.9463, 271.9364, 271.8117, 271.7072, 
    270.8912, 270.1316, 269.1808, 268.4367, 267.0734, 266.519, 265.8201, 
    264.6048,
  273.4067, 273.3718, 273.2454, 272.8258, 272.644, 272.5082, 272.0342, 
    271.5992, 270.9762, 270.2194, 269.8187, 268.282, 267.4513, 266.7802, 
    265.4939,
  273.8502, 273.9094, 273.9005, 273.4257, 273.0339, 272.5143, 272.2783, 
    271.9539, 271.498, 270.9088, 270.4562, 269.5117, 268.7364, 267.1139, 
    265.7809,
  274.3715, 274.0842, 273.7704, 273.1477, 272.7553, 272.3351, 272.2442, 
    271.6078, 271.8951, 271.2683, 271.0115, 270.3958, 269.6441, 267.9907, 
    265.5884,
  264.8485, 261.8226, 258.6352, 257.6251, 255.3609, 255.5244, 257.393, 
    258.2917, 259.5434, 258.7411, 259.711, 260.4534, 259.6194, 258.6164, 
    259.5721,
  264.939, 263.0526, 260.3246, 258.4973, 254.8922, 255.9321, 259.9143, 
    260.6246, 261.2311, 260.9344, 260.7349, 262.501, 263.4799, 262.049, 
    261.492,
  266.2, 264.54, 262.9667, 260.3157, 256.848, 252.86, 259.7895, 260.9037, 
    262.6068, 263.3028, 264.2262, 265.6049, 266.4745, 266.4392, 265.5472,
  268.5297, 267.8394, 267.5831, 266.612, 264.0532, 259.9436, 259.2373, 
    262.5152, 266.3743, 267.8515, 268.6158, 268.9484, 268.1826, 267.2114, 
    266.3065,
  270.2729, 269.4604, 269.2813, 269.3356, 269.2596, 269.1568, 268.6426, 
    265.1255, 266.2174, 269.6277, 270.5103, 269.7284, 268.3326, 267.2939, 
    266.5962,
  271.3229, 270.7757, 270.5661, 270.5894, 270.8535, 271.0863, 271.0916, 
    270.3247, 270.6325, 270.8199, 270.549, 268.6082, 267.5322, 266.8448, 
    265.9256,
  272.0076, 271.8544, 271.6376, 271.4204, 271.6872, 271.7862, 271.9788, 
    271.9507, 271.9904, 271.2619, 268.7916, 267.3141, 266.5057, 265.6406, 
    264.9945,
  272.6185, 272.4817, 272.4352, 272.3002, 272.3837, 272.5126, 272.4305, 
    272.2393, 271.9162, 268.6684, 266.9358, 265.8091, 265.1102, 264.1141, 
    263.9026,
  272.875, 272.9942, 273.0544, 272.9423, 272.7875, 272.5612, 272.5253, 
    272.2034, 269.2076, 266.2335, 265.4373, 264.2348, 263.1352, 262.4741, 
    262.4961,
  272.931, 272.9554, 273.0541, 272.8298, 272.6575, 272.381, 272.0609, 
    268.4085, 265.4445, 262.8032, 263.3811, 262.2981, 261.5197, 261.0798, 
    260.9415,
  265.5403, 263.6495, 260.6133, 259.0172, 256.2054, 254.0725, 255.1621, 
    253.4954, 252.5941, 251.0489, 252.5064, 255.7144, 258.0702, 260.4646, 
    258.7979,
  266.6209, 266.0385, 262.7542, 260.0208, 256.0629, 254.4143, 256.0239, 
    254.3988, 254.0996, 253.5834, 254.6351, 258.7436, 261.6854, 259.2861, 
    256.787,
  268.0536, 267.4197, 265.9497, 262.8373, 257.362, 253.8849, 257.9664, 
    257.9171, 257.3526, 256.7491, 258.1457, 261.0197, 261.5963, 259.546, 
    256.5813,
  268.9415, 269.286, 269.0554, 268.0204, 263.7998, 258.2495, 255.8471, 
    257.4802, 259.4228, 259.7006, 261.6896, 262.9056, 261.2722, 259.748, 
    257.38,
  269.7518, 270.0609, 269.9567, 269.7798, 269.0753, 266.8888, 263.4088, 
    258.8187, 258.1178, 263.8979, 266.1998, 264.5225, 262.4261, 261.0362, 
    259.496,
  269.8826, 270.5561, 270.6652, 270.5509, 270.4174, 270.0964, 269.1163, 
    267.1282, 265.8627, 266.8729, 267.0042, 264.9345, 263.476, 261.743, 
    259.2586,
  270.2211, 271.0021, 271.3236, 271.1268, 271.0575, 270.8814, 270.7457, 
    270.2508, 269.1502, 268.7309, 267.5009, 265.4391, 263.7412, 261.5622, 
    258.7955,
  270.9122, 271.5308, 271.7738, 271.6427, 271.4578, 271.4291, 271.2041, 
    270.9188, 269.903, 268.893, 267.4731, 265.1534, 263.4657, 260.7397, 
    258.2483,
  271.7098, 272.0356, 272.2161, 272.0922, 271.8315, 271.4651, 271.2294, 
    270.7267, 269.9523, 269.0116, 267.7866, 265.2607, 262.8379, 259.7573, 
    257.7498,
  272.6574, 272.3954, 272.3125, 271.8692, 271.2566, 270.8552, 270.5324, 
    269.7841, 269.464, 267.5574, 266.7633, 264.2271, 261.5103, 258.7262, 
    256.5848,
  267.3575, 266.9081, 266.6282, 266.5485, 265.469, 263.8641, 263.3209, 
    260.4984, 257.6758, 251.243, 249.6114, 250.4836, 248.6773, 247.6875, 
    247.0486,
  267.4657, 267.4993, 267.4184, 267.0396, 265.6382, 263.7386, 263.869, 
    261.2101, 258.3578, 256.0573, 253.5131, 253.8221, 253.1025, 249.3301, 
    249.5855,
  269.6455, 269.4814, 269.2007, 268.4765, 267.0401, 262.445, 264.4413, 
    263.2775, 259.5389, 258.4264, 257.8071, 257.5917, 257.0345, 257.5107, 
    257.0558,
  270.1795, 270.8748, 271.5123, 271.3553, 269.9694, 266.1339, 262.2182, 
    262.4231, 261.7585, 261.3696, 261.0946, 260.7076, 261.2744, 260.2775, 
    257.7611,
  270.9989, 271.5085, 271.791, 271.8543, 271.6082, 270.6885, 267.8422, 
    261.3446, 261.1185, 264.3135, 265.212, 264.3931, 262.8683, 259.2249, 
    257.7284,
  272.2804, 272.661, 272.6176, 272.3181, 272.032, 271.6338, 270.8952, 
    269.634, 267.6513, 266.6804, 267.2761, 265.7482, 261.3607, 258.2755, 
    257.0865,
  273.8977, 273.8228, 273.3608, 272.5939, 272.1495, 271.7275, 271.3522, 
    270.8399, 267.8189, 267.9675, 266.2703, 261.844, 258.2894, 256.6212, 
    255.5872,
  274.7892, 274.2829, 273.5883, 272.7967, 272.2466, 271.7763, 271.3283, 
    270.8642, 269.1584, 266.8531, 261.6937, 257.8683, 256.0136, 254.7434, 
    253.8795,
  275.3344, 274.6486, 273.8036, 272.7817, 272.0796, 271.3981, 270.8852, 
    270.3618, 268.3464, 264.8964, 261.3063, 256.356, 254.3837, 252.8896, 
    252.5486,
  275.1146, 274.0818, 273.2229, 272.0893, 271.0113, 270.3938, 269.8427, 
    267.8777, 265.0213, 260.2686, 259.3781, 255.8064, 253.0573, 251.5296, 
    250.7068,
  263.0947, 264.4114, 264.273, 266.5201, 266.5958, 267.5556, 268.6792, 
    268.8694, 268.0929, 265.1974, 261.9846, 260.4694, 256.389, 253.5354, 
    249.9489,
  266.1737, 266.4007, 267.7921, 269.3639, 268.9775, 269.8933, 270.8493, 
    269.9776, 268.376, 265.0948, 263.2322, 262.1044, 260.027, 254.4835, 
    251.9726,
  270.2901, 270.5654, 271.0823, 271.7177, 271.6249, 269.8162, 271.1732, 
    270.605, 268.606, 265.6819, 264.6625, 263.4937, 262.1636, 260.7929, 
    257.7831,
  271.7909, 273.1651, 273.5901, 273.1176, 272.8971, 272.0681, 269.9541, 
    270.3673, 268.7551, 267.1021, 265.5376, 264.2716, 264.0773, 262.9802, 
    261.3563,
  273.8167, 274.0745, 273.8706, 273.5955, 273.1483, 272.7563, 271.8872, 
    268.0272, 266.968, 267.807, 267.8332, 267.2339, 266.2543, 264.5327, 
    262.6671,
  275.0386, 275.1586, 274.6175, 273.8611, 273.4276, 272.934, 272.4229, 
    271.4908, 270.3918, 269.5043, 268.3937, 267.8011, 266.7861, 264.9158, 
    261.738,
  275.9571, 275.8017, 274.9576, 273.8707, 273.4206, 273.1108, 272.5638, 
    271.9609, 269.5184, 268.1507, 267.1776, 267.3395, 265.8302, 262.8465, 
    258.161,
  276.1331, 275.6703, 274.8687, 274.0609, 273.5352, 273.1333, 272.4353, 
    271.8048, 270.1402, 269.2122, 268.6177, 266.95, 264.1366, 258.5068, 
    254.1736,
  276.4084, 275.8928, 275.2474, 274.0858, 273.4352, 272.5723, 272.1399, 
    271.2573, 270.3276, 269.5412, 268.8912, 264.4546, 258.1282, 253.4822, 
    251.9091,
  276.0071, 275.0815, 274.4444, 273.4997, 272.7832, 272.121, 271.2561, 
    270.2334, 270.1922, 268.4736, 265.369, 258.2039, 253.0696, 250.1324, 
    248.6276,
  259.3624, 261.4762, 261.6631, 263.4342, 264.0183, 265.6605, 267.2164, 
    267.6118, 267.0166, 265.7116, 265.4065, 265.9933, 264.7307, 264.9822, 
    264.2793,
  264.5115, 264.5706, 264.3839, 264.4126, 264.6867, 267.5938, 268.284, 
    267.6667, 267.0644, 266.0706, 265.6584, 265.9405, 266.483, 265.9027, 
    265.6907,
  268.5271, 268.5727, 268.1205, 267.0983, 267.9855, 266.6612, 269.5164, 
    268.3981, 267.4268, 266.7759, 267.2242, 267.9608, 269.1502, 268.8445, 
    267.9128,
  269.1639, 270.3744, 271.3803, 271.4299, 270.4538, 270.1019, 268.3503, 
    269.3216, 269.1724, 269.0254, 269.4775, 270.157, 270.0469, 269.4313, 
    266.6648,
  270.283, 271.0813, 271.7307, 271.9655, 271.9151, 271.3869, 270.726, 
    267.6033, 267.6989, 271.1296, 271.4535, 270.8934, 270.248, 269.315, 
    265.5179,
  271.0208, 271.8442, 272.3998, 272.3536, 272.0451, 271.8564, 271.7572, 
    271.3281, 270.9268, 271.336, 270.9568, 270.3364, 270.1184, 268.723, 
    262.7292,
  272.1153, 272.9245, 273.2115, 272.7509, 272.2892, 272.0999, 272.0335, 
    271.9087, 271.3495, 270.539, 269.9566, 269.997, 269.975, 266.1209, 
    258.6475,
  273.2315, 273.8623, 273.7813, 273.2559, 272.7805, 272.737, 272.2997, 
    271.9778, 271.2527, 270.5348, 270.0558, 270.4289, 268.7307, 260.5231, 
    253.4387,
  274.5909, 274.7023, 274.4686, 273.6895, 273.2391, 272.6398, 272.3389, 
    271.6986, 271.0112, 270.6447, 270.9023, 270.3268, 264.0445, 254.0008, 
    249.8935,
  275.2657, 274.7519, 274.2804, 273.4292, 272.7243, 272.3388, 271.6585, 
    270.5888, 270.4495, 270.141, 270.8017, 267.6187, 256.2754, 250.2784, 
    247.326,
  257.8682, 259.5708, 259.2859, 259.8305, 258.4313, 257.8258, 260.2449, 
    260.9185, 262.4491, 263.2286, 263.9341, 264.9049, 264.7842, 265.03, 
    265.4256,
  263.2325, 262.998, 261.5425, 260.3114, 258.7835, 261.5176, 264.0681, 
    264.199, 265.2673, 265.7779, 265.9154, 266.2169, 265.5007, 264.8946, 
    266.236,
  267.7505, 268.2319, 267.6952, 266.3755, 266.9188, 264.8181, 267.5521, 
    267.8035, 267.3995, 266.7791, 265.995, 265.9982, 266.8009, 268.4207, 
    269.3419,
  268.1485, 269.3958, 269.8564, 270.424, 269.8422, 268.907, 266.6004, 
    269.2094, 268.6047, 266.4489, 266.7748, 267.8141, 269.1793, 269.9204, 
    269.686,
  268.9169, 269.6117, 270.1954, 270.5443, 270.7586, 270.7969, 270.2353, 
    266.1879, 266.2992, 269.6832, 270.35, 270.0219, 270.2699, 270.1921, 
    269.5981,
  269.4378, 270.1848, 270.782, 270.9825, 271.231, 271.3811, 271.3305, 
    270.8661, 270.2703, 270.6105, 270.7205, 270.5642, 270.4455, 270.2578, 
    268.6846,
  270.4115, 271.1595, 271.63, 271.6684, 271.8439, 271.897, 271.8841, 
    271.6833, 271.3225, 271.0349, 270.9319, 270.7695, 270.5466, 270.1268, 
    266.2776,
  272.076, 272.657, 272.8225, 272.723, 272.5344, 272.5811, 272.2365, 
    271.9829, 271.7236, 271.3618, 271.0889, 270.9075, 270.7157, 269.1418, 
    263.9988,
  273.6617, 273.8341, 273.835, 273.2968, 272.9111, 272.3804, 272.3092, 
    272.087, 271.8428, 271.644, 271.5849, 271.1895, 270.6163, 267.4682, 
    261.6223,
  274.6987, 274.3608, 274.0688, 273.3465, 272.8084, 272.4658, 272.2238, 
    271.9539, 271.9542, 272.1474, 271.9623, 271.4267, 269.6972, 265.3763, 
    259.2643,
  256.8493, 258.9137, 258.6238, 259.7126, 258.8105, 258.0927, 258.7505, 
    257.8284, 258.0055, 258.2924, 259.7855, 260.6229, 261.2462, 262.4113, 
    263.1736,
  261.7213, 260.7687, 259.1979, 258.7398, 257.1306, 259.6302, 262.1279, 
    261.694, 261.4322, 261.8712, 262.407, 263.4191, 264.0541, 263.6643, 
    264.834,
  267.5515, 267.7336, 266.3335, 263.9576, 260.8201, 260.0146, 265.3737, 
    265.4568, 264.7851, 264.475, 264.4403, 265.0034, 265.6437, 266.206, 
    266.6403,
  267.9786, 269.2007, 269.674, 269.9977, 268.762, 265.06, 263.4809, 267.4039, 
    267.5684, 266.8687, 266.343, 265.6663, 266.2333, 266.8741, 267.2255,
  268.6444, 269.3383, 269.9446, 270.2164, 270.5403, 270.1754, 268.8782, 
    264.6807, 264.9342, 267.9044, 268.8698, 267.2382, 266.9881, 267.7279, 
    267.3901,
  269.3558, 269.9133, 270.236, 270.4522, 270.6342, 270.8443, 270.7448, 
    269.9867, 268.8574, 269.119, 268.949, 267.9306, 267.6292, 268.0237, 
    268.3936,
  270.6895, 271.058, 271.1782, 271.1189, 271.1929, 271.2156, 271.2136, 
    271.1263, 270.4355, 269.0664, 268.6523, 268.2352, 268.5215, 268.6787, 
    268.9609,
  271.1405, 271.1455, 271.2592, 271.43, 271.5284, 271.6467, 271.4476, 
    271.3189, 270.8854, 269.7386, 268.9716, 268.5667, 268.5114, 268.4895, 
    268.978,
  270.892, 270.4137, 270.4556, 270.8594, 271.2714, 271.3776, 271.5348, 
    271.4427, 270.8758, 270.2891, 270.3409, 269.3478, 269.2075, 269.1888, 
    269.1517,
  269.1743, 268.0608, 267.8809, 268.5642, 269.0726, 269.5894, 270.0638, 
    270.4805, 270.7936, 270.9609, 271.2675, 270.9454, 270.4378, 269.9927, 
    269.6765,
  255.8503, 257.5167, 257.5086, 258.6912, 256.8679, 255.8806, 256.6182, 
    255.2778, 253.5481, 253.265, 253.8766, 254.4177, 253.5024, 253.2239, 
    252.6853,
  259.8263, 258.3006, 257.4296, 257.0131, 255.5756, 257.5812, 259.5323, 
    257.5812, 255.2237, 254.3563, 254.4975, 255.4081, 255.3611, 253.5198, 
    254.4896,
  265.7859, 265.1779, 263.3063, 260.7703, 255.6649, 253.5741, 262.1373, 
    261.3721, 259.1032, 256.0064, 256.5193, 256.8929, 256.4135, 256.3578, 
    256.8908,
  268.4403, 268.5872, 268.0628, 267.8289, 265.2447, 258.4762, 256.8315, 
    263.407, 263.3001, 261.5055, 259.8199, 259.7155, 259.9979, 260.5411, 
    260.7705,
  270.8928, 270.5329, 270.1813, 269.8887, 269.6806, 267.6935, 263.4295, 
    259.7749, 260.7627, 264.4222, 265.4767, 264.8249, 264.5487, 264.5466, 
    264.4024,
  271.1862, 271.0484, 270.8838, 270.6646, 270.5812, 270.4662, 269.4578, 
    267.9977, 265.4199, 265.7588, 265.7306, 266.1811, 266.2205, 266.1724, 
    266.0433,
  269.959, 269.3881, 269.0178, 268.8051, 268.8563, 269.0866, 269.5031, 
    269.7585, 269.3753, 267.5952, 267.6264, 267.5479, 267.3996, 267.178, 
    266.9016,
  268.7261, 267.9503, 267.3855, 267.012, 267.0724, 267.6283, 268.0348, 
    268.3358, 268.4369, 266.1867, 266.7257, 266.8719, 267.2261, 267.2537, 
    267.0433,
  267.2368, 266.1775, 265.3784, 264.7603, 264.5547, 264.8162, 265.1833, 
    265.7398, 265.9726, 265.9678, 267.4965, 267.2953, 267.2589, 266.9695, 
    266.8216,
  265.9286, 264.4647, 263.6256, 263.038, 261.8318, 260.7729, 259.0909, 
    258.4657, 262.1078, 264.1967, 266.6842, 267.566, 266.3856, 266.5431, 
    266.8129,
  258.2806, 259.208, 259.2132, 259.9489, 259.0641, 258.3542, 258.962, 
    257.4665, 256.1637, 254.2435, 253.4662, 254.0699, 252.3887, 251.8591, 
    250.1291,
  261.7192, 260.0826, 259.0724, 258.6781, 257.3004, 258.9473, 260.0568, 
    258.9023, 256.6451, 255.5452, 255.114, 255.64, 254.4766, 251.3158, 
    250.2378,
  268.6279, 267.6459, 265.3756, 262.0088, 258.069, 255.5063, 261.1068, 
    260.6042, 258.966, 256.0526, 256.6022, 256.0454, 255.0323, 253.3615, 
    251.725,
  270.6183, 270.7796, 270.4751, 269.7201, 266.3409, 259.1387, 256.5433, 
    261.5446, 261.6965, 259.8147, 257.913, 257.4832, 256.1951, 255.5166, 
    253.8376,
  270.1686, 269.8361, 269.8859, 270.0005, 270.0059, 267.4293, 262.0248, 
    257.0414, 256.609, 261.683, 262.305, 260.5566, 258.3811, 256.4889, 
    254.7444,
  269.4949, 269.0154, 268.6774, 268.7291, 268.9562, 269.0956, 267.8463, 
    265.3768, 262.5332, 260.8917, 261.8284, 262.4015, 262.3908, 261.9073, 
    261.0554,
  269.162, 268.5274, 267.6753, 267.1015, 267.0242, 267.3453, 267.6766, 
    267.6513, 267.2298, 265.778, 264.7718, 264.8461, 264.5049, 264.2105, 
    264.1913,
  268.7305, 267.9916, 266.9782, 266.1841, 265.6374, 265.3069, 264.4906, 
    264.4176, 263.7897, 258.7258, 257.4785, 256.5891, 256.3236, 256.9306, 
    257.5249,
  268.509, 267.4057, 266.1234, 265.0316, 263.7841, 262.8721, 261.7977, 
    260.6737, 259.2197, 258.0067, 259.7229, 256.4367, 255.3977, 254.6799, 
    255.4227,
  268.1432, 266.743, 265.1683, 264.3249, 262.6115, 260.3572, 256.2273, 
    253.336, 253.3184, 252.6122, 255.3591, 254.6203, 254.4555, 254.7815, 
    255.573,
  258.2304, 259.5573, 259.3303, 260.1291, 259.1146, 258.9696, 259.5122, 
    258.9996, 257.8643, 255.6636, 255.39, 255.8432, 255.4655, 254.899, 254.482,
  263.526, 262.5023, 260.5592, 259.847, 257.7102, 259.6003, 260.8481, 
    259.9616, 258.7305, 257.5278, 257.0488, 256.9957, 256.3514, 254.2678, 
    254.2251,
  269.5044, 268.9904, 267.2719, 264.3009, 259.1603, 256.8311, 261.8976, 
    261.6319, 260.571, 258.8101, 258.5776, 258.0593, 257.1048, 256.3936, 
    255.3579,
  270.5539, 270.5271, 270.2363, 269.8046, 266.7958, 260.4024, 257.7167, 
    262.4615, 262.5589, 260.8507, 259.9726, 259.2396, 258.1275, 257.3085, 
    256.2359,
  271.0057, 270.3913, 269.7939, 269.268, 269.1585, 267.3846, 263.6034, 
    258.7626, 258.9117, 262.2118, 262.9216, 261.4752, 260.3725, 258.7647, 
    257.7252,
  270.763, 270.1643, 269.4188, 268.8133, 268.0532, 267.8364, 267.7683, 
    266.6237, 264.0682, 260.9309, 260.5773, 260.7088, 260.1596, 259.9282, 
    259.5031,
  270.0787, 269.4432, 268.5655, 267.4905, 266.9211, 266.3417, 265.9256, 
    265.9537, 265.4214, 263.5662, 261.8905, 261.511, 261.6174, 260.9754, 
    259.2881,
  269.1478, 268.2094, 266.931, 265.6994, 264.3509, 263.7261, 262.5805, 
    261.593, 260.0035, 256.7271, 256.5318, 255.9436, 255.5623, 255.876, 
    254.9148,
  267.5387, 266.4879, 264.9886, 263.0361, 260.8343, 259.0997, 257.79, 
    256.7774, 255.4758, 254.5878, 256.6902, 252.5045, 253.1409, 251.8668, 
    251.0908,
  265.3193, 264.1526, 262.5792, 260.2933, 257.2401, 254.7634, 251.8561, 
    250.5691, 250.1908, 248.4616, 250.6518, 249.2617, 249.2608, 248.4975, 
    250.217,
  259.5765, 260.3142, 259.9316, 259.996, 258.7019, 257.1671, 258.2904, 
    257.5752, 256.7611, 253.2079, 254.0952, 254.3368, 252.9014, 251.5793, 
    250.673,
  264.7212, 263.2678, 261.4464, 259.9783, 258.8015, 259.6718, 260.0662, 
    258.3376, 256.6794, 254.7453, 255.2578, 256.1824, 255.3902, 252.0262, 
    252.2162,
  269.696, 269.2352, 267.8322, 264.299, 259.6219, 256.8372, 261.7048, 
    260.8216, 258.6968, 255.0511, 256.3751, 256.7003, 255.9293, 255.0012, 
    253.6202,
  270.1526, 270.2483, 270.2084, 269.7584, 266.339, 260.3199, 257.8156, 
    262.0714, 261.3394, 258.0151, 257.2246, 256.9819, 256.1886, 256.116, 
    255.2486,
  269.4493, 268.735, 268.5261, 268.8205, 269.0553, 266.2853, 262.1081, 
    257.953, 257.6644, 260.6484, 260.3659, 258.9103, 257.4579, 256.6655, 
    255.9288,
  269.1696, 267.8738, 266.8421, 266.4544, 267.0945, 267.2213, 265.9675, 
    264.7986, 262.5349, 261.1851, 260.6603, 260.0343, 258.9456, 257.887, 
    256.7629,
  268.6405, 266.7607, 265.3185, 264.4139, 263.8358, 263.9912, 264.3458, 
    264.0586, 262.2545, 261.0371, 260.4705, 259.8442, 259.6586, 258.9742, 
    258.2451,
  267.9431, 265.9431, 263.9236, 262.5793, 261.3265, 260.0359, 258.5466, 
    257.65, 255.6314, 254.707, 256.428, 256.8822, 257.3791, 257.5423, 257.5015,
  267.493, 265.471, 263.3966, 261.6335, 259.7771, 257.9201, 256.2343, 
    254.8426, 253.5123, 252.2588, 253.2061, 251.0104, 251.8296, 252.3166, 
    253.2559,
  267.2025, 264.6978, 261.9988, 259.8304, 257.8416, 254.3114, 251.3504, 
    249.3238, 248.1792, 245.9162, 247.4318, 246.3468, 245.9716, 246.8663, 
    248.2567,
  262.519, 262.1592, 260.9081, 261.037, 259.0621, 257.4977, 258.0021, 
    256.8572, 256.2811, 252.9934, 252.8911, 252.9163, 249.5578, 248.3189, 
    246.4758,
  265.1408, 264.1084, 262.2445, 261.4221, 259.079, 260.1812, 260.4561, 
    258.2373, 256.4998, 255.3257, 254.4316, 255.1806, 253.4978, 248.6598, 
    247.3654,
  268.67, 267.7108, 266.4572, 263.6375, 260.6833, 258.057, 262.2372, 261.261, 
    258.6005, 255.6259, 256.7066, 256.8607, 255.1329, 253.1202, 250.0469,
  270.1092, 269.6364, 268.7363, 267.7716, 266.0578, 262.0961, 258.6283, 
    262.0018, 261.3663, 257.9258, 256.8596, 257.0083, 256.2312, 254.9252, 
    252.5094,
  270.7804, 269.5921, 267.9908, 267.0809, 267.3621, 266.0792, 263.3871, 
    258.1598, 255.6961, 259.6073, 259.946, 258.0358, 257.2911, 256.1572, 
    254.0561,
  271.1431, 269.5194, 267.4882, 266.2968, 266.2279, 266.5073, 265.2539, 
    263.0181, 257.9952, 256.6224, 257.8137, 258.8496, 257.6965, 256.8841, 
    254.8739,
  271.21, 269.3677, 267.0395, 265.3314, 264.3618, 264.1625, 263.3239, 
    260.8801, 257.4973, 255.8823, 256.4927, 257.2144, 257.3887, 256.7846, 
    255.8023,
  270.6951, 268.7843, 266.4247, 265.4009, 264.5265, 263.2781, 261.0489, 
    258.5249, 254.4439, 252.1544, 252.1454, 254.0443, 257.0293, 256.7541, 
    256.0692,
  268.5573, 266.2968, 264.3085, 262.8271, 262.2754, 260.6915, 258.5765, 
    255.9376, 253.2142, 250.509, 250.5535, 249.839, 253.7069, 256.4217, 
    256.0323,
  263.8773, 262.1024, 260.0594, 258.0189, 255.5393, 253.0343, 251.5419, 
    250.0156, 246.9678, 243.1668, 245.1929, 246.2654, 250.1486, 255.276, 
    255.8916,
  265.7296, 265.9221, 264.8035, 263.7965, 261.2394, 259.1031, 260.0065, 
    257.8787, 257.9314, 254.8714, 255.3755, 254.9765, 251.3626, 248.9453, 
    246.274,
  266.3174, 265.7651, 264.6776, 263.4742, 260.7194, 260.8499, 260.9579, 
    258.7911, 258.1895, 257.9209, 256.7571, 257.0025, 254.9601, 249.8288, 
    247.4076,
  268.599, 267.6929, 265.9992, 263.5721, 260.8211, 257.8207, 261.9285, 
    260.7358, 258.7666, 257.0639, 258.958, 258.9943, 256.912, 254.0613, 
    250.619,
  269.5299, 269.5062, 268.1469, 265.9574, 262.3697, 260.0174, 257.0594, 
    261.1732, 260.446, 257.8027, 257.8254, 257.997, 257.5853, 256.1739, 
    253.2655,
  270.8765, 269.8094, 268.5551, 267.1246, 265.3295, 262.768, 260.7346, 
    256.9649, 256.7739, 259.0754, 259.2433, 257.8517, 257.131, 257.0187, 
    255.7498,
  271.0287, 269.782, 268.8055, 267.7647, 266.9299, 266.288, 265.0495, 
    262.5808, 259.1078, 257.6788, 257.3604, 258.2994, 257.4521, 256.5569, 
    255.7219,
  271.0442, 269.9397, 268.7471, 267.2491, 266.2018, 265.7957, 266.1642, 
    265.2466, 261.1222, 257.8339, 254.9673, 253.7502, 254.6792, 255.0965, 
    255.1504,
  270.2902, 268.419, 265.8513, 263.5885, 262.0587, 261.8935, 263.544, 
    264.7274, 260.3332, 255.6183, 251.8418, 250.4309, 249.4586, 249.5005, 
    251.1094,
  266.1916, 264.0845, 261.3191, 259.0779, 257.3664, 257.532, 261.5709, 
    262.8397, 259.3735, 255.207, 251.1419, 248.271, 246.6143, 245.9008, 
    246.7469,
  261.8166, 259.6794, 257.3674, 254.1465, 252.1602, 250.7876, 252.6101, 
    255.5708, 253.8783, 249.97, 247.0669, 245.3542, 244.0988, 244.6384, 
    246.3533,
  260.1137, 264.4708, 264.451, 265.6428, 264.9502, 264.1336, 264.0491, 
    261.486, 259.0717, 255.6937, 253.8002, 251.6237, 247.9421, 247.7948, 
    248.2999,
  262.8621, 263.3867, 264.0115, 264.2947, 263.101, 264.6518, 264.8719, 
    261.8455, 259.4596, 256.7419, 255.282, 255.1322, 252.4654, 246.2941, 
    247.5082,
  266.646, 266.6809, 265.4124, 263.9413, 263.3382, 261.9774, 264.8224, 
    262.4066, 259.9672, 257.7833, 258.0743, 257.0597, 253.1557, 251.2511, 
    249.1424,
  268.0626, 268.2538, 267.9571, 266.7161, 264.7049, 263.119, 260.765, 
    261.661, 259.9545, 257.7208, 257.7203, 257.7876, 254.7279, 252.3661, 
    250.8445,
  269.9186, 269.1553, 268.5104, 267.5331, 266.286, 264.299, 261.9523, 256.3, 
    255.191, 257.3157, 257.3785, 257.2142, 255.9085, 254.4288, 251.7493,
  270.1235, 269.3401, 268.5209, 267.7331, 266.8968, 265.7173, 264.4611, 
    261.8102, 259.4704, 257.5637, 256.7379, 257.192, 257.2705, 256.7483, 
    253.2874,
  269.4857, 268.4139, 267.5032, 266.4738, 265.8264, 265.0855, 264.367, 
    263.7572, 261.9448, 259.6951, 257.2626, 256.5491, 256.8992, 257.5317, 
    255.9789,
  266.7759, 264.9875, 263.4538, 261.568, 260.2572, 259.1936, 258.3834, 
    258.6205, 258.5764, 258.1844, 258.2538, 256.9541, 256.6722, 256.846, 
    256.6342,
  264.2048, 262.5214, 260.5893, 258.3626, 255.8397, 254.4026, 253.9166, 
    253.4482, 252.8414, 254.3448, 259.0063, 257.8785, 256.508, 255.7217, 
    254.8214,
  261.5355, 259.6007, 257.1347, 253.8145, 251.5995, 249.7448, 248.9353, 
    249.5137, 249.8664, 251.8266, 256.8755, 257.2367, 255.5982, 254.6436, 
    254.2259,
  258.9515, 261.7861, 260.2559, 262.7343, 262.6916, 262.2028, 262.3142, 
    260.8023, 257.8969, 257.0753, 256.8641, 256.7953, 256.7757, 256.4402, 
    255.4928,
  262.8762, 262.6437, 261.6558, 261.1584, 261.6647, 262.6978, 263.0255, 
    262.0791, 259.3283, 258.739, 258.4235, 259.0119, 258.2946, 254.7165, 
    254.3462,
  267.9726, 266.6229, 264.4937, 261.7786, 260.2181, 258.6007, 263.5027, 
    263.3984, 262.0354, 260.0244, 260.6469, 259.9033, 258.4273, 256.7143, 
    254.0131,
  269.2778, 268.6816, 268.3456, 266.6597, 262.7507, 261.858, 259.9557, 
    263.4502, 262.8788, 260.762, 260.3755, 260.092, 258.2784, 256.5479, 
    253.9696,
  269.2502, 268.8187, 268.6051, 267.8567, 266.8408, 264.497, 263.5087, 
    259.9793, 259.3461, 260.4725, 260.5223, 259.4872, 257.3534, 255.6873, 
    253.1993,
  267.745, 267.4123, 267.5164, 267.7109, 267.5835, 266.821, 266.0487, 
    264.8187, 263.0082, 261.4704, 260.6462, 259.6751, 257.1773, 254.8302, 
    252.4746,
  266.3126, 265.276, 264.7988, 264.6681, 265.3491, 265.5324, 265.588, 
    265.3077, 263.9749, 262.4993, 261.0302, 258.8835, 256.2444, 253.8124, 
    251.0933,
  264.8168, 263.5313, 262.0832, 260.721, 259.8764, 259.6368, 259.8839, 
    261.3268, 261.2073, 261.3552, 259.9937, 258.101, 255.5562, 252.9709, 
    250.8201,
  264.2637, 262.3512, 260.537, 258.069, 255.5051, 254.3804, 253.4011, 
    253.5042, 256.1054, 258.4733, 258.9552, 257.2526, 254.053, 252.1856, 
    250.4113,
  263.5679, 260.313, 257.4388, 253.5232, 250.6752, 249.0834, 248.9118, 
    249.9523, 249.8245, 251.7583, 256.2933, 255.2076, 253.4559, 251.9927, 
    251.5037,
  259.3647, 261.1281, 257.6736, 261.4642, 260.4628, 259.3979, 259.2791, 
    257.6154, 256.5186, 255.1845, 256.3615, 258.0822, 258.4315, 258.3835, 
    257.1985,
  262.7127, 260.5942, 258.1318, 259.827, 259.9902, 259.9719, 259.4239, 
    257.679, 256.4288, 257.2317, 257.4703, 259.2896, 259.3737, 256.1886, 
    255.8067,
  267.6808, 266.5638, 261.7386, 258.6731, 259.295, 254.6455, 259.7766, 
    258.6017, 257.6889, 258.2065, 259.2343, 259.0093, 258.2181, 257.5839, 
    256.3385,
  268.3203, 268.4325, 267.0402, 263.9083, 260.3575, 258.602, 255.9849, 
    258.878, 258.776, 258.7666, 259.0222, 258.7038, 257.3813, 257.0477, 
    256.9563,
  266.8659, 267.5876, 268.0358, 267.0499, 264.3426, 261.6275, 260.0832, 
    253.4382, 254.25, 258.0576, 258.8567, 258.2426, 257.36, 257.1375, 257.2946,
  265.9573, 265.6636, 266.7537, 267.3863, 266.6514, 265.2334, 263.2896, 
    261.0786, 259.8253, 259.0999, 259.4756, 258.9443, 257.727, 256.6853, 
    256.3159,
  265.0841, 264.3748, 263.8925, 265.4633, 266.6917, 266.4443, 265.5981, 
    264.0904, 261.855, 260.9465, 260.011, 258.6042, 257.3086, 256.5957, 
    256.5806,
  264.4642, 263.0626, 261.5211, 260.8034, 262.5921, 264.3416, 264.5669, 
    264.2077, 261.7162, 260.295, 258.7784, 258.7396, 257.6906, 256.7689, 
    256.8138,
  263.1194, 261.8072, 259.7455, 257.4241, 255.1464, 256.5617, 258.4937, 
    260.3317, 260.4142, 259.946, 258.6271, 259.0291, 258.007, 256.9186, 
    255.4392,
  260.5927, 258.795, 256.5107, 253.0553, 250.4969, 249.7306, 252.1907, 
    256.6321, 256.8598, 257.5459, 258.9302, 259.3798, 258.2708, 257.2096, 
    254.6716,
  262.5491, 264.2681, 260.9857, 262.6975, 261.69, 260.3424, 260.5331, 
    260.1221, 259.3933, 255.4837, 255.9528, 256.6461, 254.8307, 254.5248, 
    253.5761,
  266.7186, 264.7673, 263.0605, 262.5315, 260.6611, 259.1898, 260.044, 
    259.1767, 257.6461, 257.3087, 256.4319, 258.45, 258.3035, 253.1466, 
    252.7337,
  268.6942, 268.2741, 265.5894, 263.2716, 259.7481, 254.4153, 258.4943, 
    257.7011, 256.9889, 257.5829, 258.3227, 258.1978, 258.1505, 257.5843, 
    254.372,
  268.1731, 268.953, 268.5168, 265.7288, 260.6806, 257.1396, 251.2706, 
    256.3083, 257.0477, 257.4733, 257.6559, 257.8509, 257.53, 257.4424, 
    256.4164,
  267.8203, 268.0166, 268.2791, 267.1393, 263.6847, 259.3195, 257.5828, 
    251.0237, 252.091, 255.7845, 257.095, 257.6774, 257.517, 257.6652, 
    257.2274,
  267.0742, 267.5505, 267.9668, 267.7, 265.8532, 263.4252, 260.6225, 259.556, 
    258.7724, 259.159, 258.7552, 258.2989, 257.4672, 256.1897, 255.3148,
  266.0034, 266.1209, 266.7069, 267.1967, 267.0973, 265.3281, 263.9731, 
    262.1664, 261.3322, 261.2005, 259.7767, 258.1454, 256.7071, 254.7737, 
    252.2021,
  265.0225, 264.6651, 264.4318, 265.1044, 266.0088, 265.8589, 264.225, 
    263.0288, 260.7294, 260.0538, 258.2347, 257.1195, 254.838, 251.3865, 
    249.6933,
  263.2936, 262.756, 261.9857, 261.0374, 261.3395, 262.6452, 262.5064, 
    260.9498, 259.5047, 257.9142, 256.2209, 254.7819, 252.2962, 251.1539, 
    250.4302,
  260.4746, 259.4309, 257.9364, 255.6375, 256.204, 258.5423, 259.7288, 
    259.4344, 256.8571, 255.7941, 254.7109, 253.4585, 252.5274, 251.7395, 
    251.854,
  262.8008, 265.5046, 264.2134, 262.9893, 261.0971, 261.8185, 260.251, 
    258.4093, 257.2448, 255.2774, 256.7703, 257.0499, 255.6754, 254.0527, 
    252.4962,
  267.4897, 265.128, 261.972, 258.153, 256.0536, 260.3367, 260.9488, 
    258.7765, 257.3415, 257.0778, 256.8732, 258.3445, 257.7018, 252.2411, 
    250.8405,
  268.6677, 266.6702, 262.3041, 257.7321, 256.1638, 256.6758, 260.3617, 
    258.6697, 257.8424, 257.6944, 257.7835, 258.1364, 257.3242, 255.3496, 
    252.164,
  268.7987, 267.7111, 265.5858, 262.0323, 259.066, 258.9456, 254.9093, 
    257.615, 257.7805, 257.4851, 257.2905, 257.0805, 256.2536, 256.9085, 
    255.1356,
  268.9128, 267.7718, 266.4286, 264.1713, 261.8866, 259.9359, 259.0498, 
    252.2242, 252.5081, 254.0979, 255.8879, 255.835, 255.8709, 256.7921, 
    257.0762,
  268.9334, 268.282, 267.1697, 265.5428, 264.1026, 262.3861, 259.7806, 
    258.8087, 257.7039, 256.8735, 255.4381, 255.8028, 255.8846, 256.4763, 
    256.4601,
  268.7224, 268.2008, 267.6755, 266.6083, 265.3511, 264.2231, 262.6752, 
    260.8864, 259.5746, 259.4274, 257.6776, 255.7511, 255.5908, 255.2082, 
    254.5137,
  267.8798, 267.6974, 267.3541, 267.0071, 266.2329, 264.9384, 263.6749, 
    261.581, 258.341, 257.361, 255.9715, 255.1099, 253.8744, 252.9095, 251.205,
  265.9893, 265.9068, 265.6517, 264.7605, 264.0768, 263.4591, 261.7858, 
    259.2862, 256.5165, 253.9953, 253.0697, 253.9533, 252.1865, 250.5223, 
    249.0369,
  262.7968, 262.0086, 261.2825, 259.4465, 258.527, 258.1184, 257.9107, 
    257.4862, 253.9854, 251.6408, 250.9177, 251.7802, 250.3561, 248.9652, 
    248.7043,
  260.1582, 260.5937, 257.5218, 259.3511, 256.5665, 255.6309, 257.4353, 
    257.7431, 256.4259, 249.8255, 250.8193, 256.9603, 256.5003, 255.8158, 
    259.262,
  263.0614, 259.7917, 258.5364, 257.61, 256.7174, 258.3456, 259.0949, 
    257.5255, 254.2365, 256.6063, 254.8395, 259.3376, 258.7904, 255.0002, 
    255.6796,
  266.7009, 263.9693, 261.1272, 259.6118, 259.53, 255.6739, 257.1904, 
    256.0883, 255.7719, 256.5471, 257.7572, 258.256, 258.8859, 257.957, 
    256.1837,
  267.7941, 266.2822, 264.5872, 261.7119, 259.5012, 258.1497, 252.0787, 
    253.5284, 255.2595, 255.5293, 255.8687, 256.6576, 257.7457, 258.1452, 
    257.0709,
  268.1383, 266.6704, 265.5092, 263.6796, 260.8338, 259.4535, 258.0981, 
    247.3064, 251.0675, 255.1502, 255.8579, 256.1041, 256.8285, 258.4649, 
    257.8303,
  268.7042, 267.5868, 266.2706, 265.0709, 263.4953, 261.2373, 259.2246, 
    258.666, 255.9721, 257.1442, 256.1632, 256.3618, 257.1744, 257.3633, 
    256.5391,
  269.1887, 268.2482, 267.0765, 265.9666, 264.9578, 263.6075, 261.6677, 
    259.1955, 258.3399, 257.4933, 256.2592, 255.8588, 256.1735, 255.9995, 
    255.0491,
  269.4417, 268.5548, 267.7073, 266.7417, 265.7743, 264.2832, 262.5178, 
    259.5918, 256.838, 255.821, 254.5765, 254.4962, 253.4864, 253.0546, 
    251.6514,
  268.5591, 267.6459, 266.3099, 264.748, 263.1602, 262.5417, 260.4155, 
    257.3625, 254.2086, 251.4961, 250.4802, 251.1407, 250.6754, 250.6327, 
    250.7236,
  265.0728, 264.2779, 262.0401, 258.5061, 257.1894, 255.9195, 255.9106, 
    255.2943, 251.6093, 248.6673, 249.457, 251.1379, 251.1704, 250.5969, 
    251.3561,
  257.9644, 258.0091, 255.6467, 255.8412, 252.9235, 252.999, 255.1488, 
    256.0185, 256.3629, 255.3064, 255.8495, 259.6469, 259.0942, 258.2689, 
    257.4859,
  260.5505, 258.9678, 256.6179, 255.0483, 253.1602, 253.0346, 255.1703, 
    254.8212, 254.789, 256.7829, 256.1165, 259.3869, 259.8803, 256.5662, 
    255.8643,
  264.0381, 261.3195, 258.7736, 256.9182, 255.4938, 248.8047, 254.1784, 
    254.6776, 254.9256, 253.8706, 256.0666, 257.2714, 258.6552, 258.5058, 
    257.3299,
  266.8465, 265.303, 263.4409, 260.4852, 257.9162, 255.7293, 247.5808, 
    250.001, 252.3343, 252.4616, 252.8667, 255.8846, 256.2092, 257.4569, 
    257.7965,
  267.3848, 265.8771, 264.7803, 262.7169, 259.9536, 259.1902, 257.9879, 
    249.4279, 250.9509, 252.2629, 252.3411, 253.2151, 254.3418, 256.8184, 
    258.0437,
  268.2387, 267.0825, 265.9339, 264.7117, 263.2306, 260.8304, 258.6119, 
    258.2117, 255.0852, 255.286, 251.9159, 254.8976, 254.5607, 256.5997, 
    256.9116,
  269.1262, 268.099, 266.9952, 265.9009, 264.8884, 263.2811, 260.6697, 
    257.2203, 255.06, 253.1945, 252.0741, 254.4123, 255.5329, 257.1703, 
    256.2548,
  269.8292, 268.8161, 267.7433, 266.7978, 265.6845, 263.7257, 261.2489, 
    257.258, 252.6069, 250.7507, 250.1187, 253.5325, 256.4871, 256.761, 
    254.6348,
  269.7912, 268.3937, 266.8028, 265.0577, 263.3669, 261.6619, 259.1346, 
    255.0638, 251.2154, 249.6709, 248.7415, 249.9481, 253.6655, 254.8763, 
    253.7361,
  268.5211, 266.154, 263.2618, 257.9738, 256.7384, 253.2819, 253.3299, 
    252.9447, 249.2121, 247.7163, 246.5856, 248.8676, 249.3638, 252.4926, 
    252.6355,
  256.4721, 257.5781, 255.621, 256.9161, 256.0211, 254.8228, 255.8035, 
    255.1345, 256.0108, 256.7404, 257.4541, 257.7039, 255.0597, 254.7662, 
    256.2505,
  259.8851, 258.127, 257.4997, 256.7454, 256.0506, 253.1707, 256.0845, 
    254.9425, 255.5624, 257.3906, 258.2926, 259.3844, 257.2887, 253.447, 
    253.5788,
  264.569, 261.8409, 259.5902, 257.5487, 256.0846, 251.7613, 256.2069, 
    254.8638, 255.4803, 256.7134, 258.875, 259.8923, 258.0545, 256.4498, 
    255.0079,
  266.8842, 265.8691, 264.5504, 261.7615, 259.0237, 258.812, 253.8055, 
    253.1197, 255.1046, 255.9028, 257.8905, 258.9549, 257.6884, 256.6732, 
    256.6505,
  267.9582, 266.6742, 265.7675, 264.6625, 261.0193, 260.2082, 258.3888, 
    250.56, 250.7349, 255.2787, 256.56, 257.1966, 256.9368, 256.822, 257.5318,
  269.6251, 268.6273, 267.4679, 266.1002, 264.7416, 262.265, 258.5814, 
    256.6274, 254.7124, 255.4906, 255.5805, 256.1548, 255.7933, 255.8612, 
    256.612,
  270.8566, 270.3976, 269.4339, 268.1096, 266.51, 264.3634, 261.2987, 
    256.6786, 254.4491, 253.8769, 255.1931, 255.6109, 255.07, 255.0488, 
    255.2842,
  271.5371, 271.0473, 270.1776, 268.8645, 267.7426, 265.28, 261.2697, 
    256.776, 252.7271, 252.6949, 252.9075, 254.8871, 254.7777, 254.099, 
    253.6758,
  271.9225, 271.1337, 270.139, 268.2844, 266.2176, 263.3201, 259.4117, 
    254.1694, 251.5908, 250.9631, 250.1951, 251.4462, 253.8402, 253.4712, 
    253.8113,
  272.3265, 270.8173, 269.2588, 264.2263, 260.8695, 258.3783, 256.649, 
    253.7998, 249.6589, 249.3002, 246.757, 248.7086, 249.162, 252.0854, 
    253.4763,
  255.3948, 257.3109, 257.8781, 258.8806, 258.7012, 257.4215, 257.7094, 
    257.0739, 257.0902, 254.8787, 252.4065, 251.5688, 252.3782, 254.8404, 
    255.754,
  259.5216, 258.3977, 258.4005, 257.972, 258.1831, 256.2743, 258.1434, 
    257.5681, 256.7863, 256.7904, 254.5416, 254.8147, 255.6751, 254.1184, 
    254.537,
  265.3436, 263.8683, 262.2882, 260.7336, 260.7462, 257.0123, 259.8248, 
    257.5578, 256.6073, 257.0542, 256.2798, 255.5361, 255.8719, 257.6377, 
    256.5939,
  267.2279, 267.3952, 267.6779, 266.8819, 264.4803, 263.3724, 254.4501, 
    255.7629, 256.5479, 257.1497, 257.2856, 256.2344, 255.6092, 257.0347, 
    257.643,
  268.4406, 268.4764, 268.5846, 268.1969, 264.7822, 260.9399, 257.8286, 
    249.7699, 250.3181, 256.3066, 256.7588, 255.5468, 255.5473, 257.1457, 
    258.5019,
  269.5281, 269.3827, 268.935, 267.715, 265.6223, 261.4318, 258.3323, 
    257.1279, 256.3342, 256.9212, 255.5778, 254.8762, 255.3038, 257.8293, 
    257.9351,
  270.3022, 269.5055, 268.5154, 266.9298, 265.1103, 262.5214, 260.2624, 
    257.8064, 256.9536, 256.1147, 255.1301, 254.515, 255.3376, 257.4582, 
    257.144,
  270.4604, 269.223, 267.6744, 265.6277, 263.7799, 261.4872, 259.3673, 
    256.6844, 255.3249, 254.634, 253.8669, 253.7752, 255.8722, 256.473, 
    254.6808,
  270.1495, 268.6578, 266.2406, 263.0292, 259.6804, 257.7516, 255.9151, 
    254.389, 253.7932, 253.1405, 253.0492, 253.6203, 254.7221, 254.8627, 
    253.2182,
  269.178, 266.6733, 263.1808, 257.4813, 255.3477, 253.5261, 252.9972, 
    252.8817, 250.8657, 249.9269, 250.1884, 252.1461, 252.6351, 252.031, 
    251.6833,
  258.1159, 258.0019, 256.9135, 256.0568, 255.1978, 254.5105, 255.2814, 
    254.6886, 254.6572, 253.4547, 253.2172, 254.3491, 254.3583, 254.3321, 
    252.6348,
  260.6983, 258.9394, 258.0656, 256.9722, 255.6802, 255.596, 256.6505, 
    256.3278, 256.0279, 256.9195, 255.8878, 256.6416, 258.1593, 253.4421, 
    250.7647,
  263.1993, 260.2472, 259.1696, 257.7864, 256.8615, 253.4834, 257.3403, 
    257.8212, 257.4596, 258.6369, 257.542, 255.9469, 257.9187, 257.9741, 
    253.4127,
  265.657, 263.7017, 263.3908, 262.207, 259.9038, 259.4326, 254.0213, 
    256.3853, 257.7206, 256.8319, 255.0568, 253.3591, 256.4509, 255.8403, 
    253.8074,
  268.1214, 267.1533, 266.2969, 265.0422, 260.8422, 259.6048, 260.3523, 
    252.0682, 251.1162, 250.8697, 251.1602, 254.2961, 255.9211, 255.2305, 
    254.2304,
  268.3538, 267.4265, 266.4547, 265.6134, 263.437, 261.3891, 260.0529, 
    258.6929, 255.8614, 254.3798, 252.3544, 255.6105, 255.4263, 254.5918, 
    253.2174,
  267.9075, 267.2919, 266.5291, 265.4812, 264.352, 262.9178, 260.5021, 
    257.5981, 256.0724, 255.2233, 254.8559, 253.997, 253.1128, 251.327, 
    250.4268,
  267.3879, 266.6723, 265.8954, 265.1609, 264.3798, 262.8622, 260.703, 
    256.9752, 254.7249, 253.9542, 253.4862, 252.8308, 251.6149, 250.0122, 
    248.5515,
  266.2979, 265.4027, 264.5079, 263.0174, 261.5652, 260.0173, 257.8925, 
    255.6128, 253.9617, 253.4452, 253.2407, 252.9701, 251.9832, 250.981, 
    250.5781,
  263.4525, 262.1016, 259.8285, 256.5739, 256.1638, 255.1827, 255.0073, 
    255.1714, 253.3384, 252.5773, 252.4239, 252.7886, 252.5892, 251.0793, 
    251.3906,
  259.6594, 259.6959, 258.1198, 258.0266, 256.0356, 253.9415, 254.9071, 
    253.1229, 251.2142, 245.6282, 246.1011, 247.7277, 245.9202, 246.4142, 
    246.5402,
  261.832, 261.4528, 259.9399, 258.6236, 256.3426, 255.7336, 255.717, 
    253.6452, 252.5464, 250.9685, 249.6693, 251.9886, 252.878, 249.3361, 
    248.8318,
  265.1669, 262.4283, 260.5244, 259.0469, 257.0696, 253.2839, 255.646, 
    254.2268, 252.5174, 252.9063, 253.4852, 254.3932, 255.6874, 257.2113, 
    256.4086,
  265.2683, 264.628, 263.2094, 260.7904, 258.0748, 257.462, 251.5555, 
    252.3004, 252.0209, 252.4069, 254.0186, 254.8592, 256.5003, 257.3758, 
    257.6135,
  266.0085, 264.9321, 264.0466, 262.2733, 258.8578, 258.2462, 257.6523, 
    247.7184, 246.3637, 248.8479, 249.347, 252.819, 254.6036, 254.6872, 
    255.0399,
  266.6751, 265.5574, 264.3076, 262.9364, 261.155, 259.9201, 258.4742, 
    258.5613, 254.6217, 253.913, 249.264, 251.9627, 251.8257, 251.2547, 
    251.9254,
  267.7079, 266.5639, 265.4038, 264.5212, 264.2095, 263.4015, 260.2778, 
    257.6334, 254.2996, 252.6492, 251.0964, 250.4809, 249.7196, 248.7232, 
    249.2599,
  268.6736, 267.7421, 266.8856, 266.0229, 265.2056, 263.4338, 260.7358, 
    255.4098, 252.2218, 249.771, 248.6612, 248.4994, 247.7053, 246.8563, 
    247.1276,
  268.7979, 267.8493, 266.7884, 265.1939, 263.3028, 260.6954, 257.1738, 
    252.8428, 250.241, 247.7646, 247.0839, 247.1858, 246.8276, 247.0256, 
    246.4516,
  266.1679, 264.4897, 261.7177, 257.7212, 256.6281, 254.9033, 253.4504, 
    252.864, 248.5993, 244.5812, 244.1757, 246.8428, 246.9509, 247.0382, 
    247.0666,
  258.5774, 260.6189, 260.2931, 260.2328, 257.3164, 255.4136, 256.1617, 
    253.6047, 249.9416, 245.0064, 244.9604, 245.9501, 243.3434, 244.1499, 
    243.2958,
  260.4047, 260.5326, 260.4219, 259.1315, 255.6835, 255.6696, 255.7246, 
    252.7113, 249.7059, 248.3403, 246.5258, 250.0797, 250.988, 246.8193, 
    246.591,
  266.0965, 262.0516, 259.9335, 258.1371, 256.3777, 252.0197, 254.1913, 
    251.5973, 249.414, 250.0994, 250.8402, 251.7469, 252.9874, 254.6717, 
    254.1205,
  267.1063, 264.3196, 262.2508, 259.5925, 257.7479, 256.232, 247.9765, 
    249.4947, 248.1381, 248.6578, 250.6091, 252.0432, 253.7582, 255.4126, 
    255.5776,
  267.2736, 265.0971, 263.9026, 262.061, 258.4732, 257.9911, 256.6007, 
    245.9048, 242.6245, 248.0638, 248.0199, 250.2049, 253.1985, 253.5503, 
    253.6897,
  267.5551, 266.1518, 265.0611, 263.5836, 261.2599, 259.4914, 257.7028, 
    258.369, 252.9639, 250.6239, 246.0374, 249.9731, 250.8133, 250.3887, 
    250.9305,
  268.0159, 266.8268, 265.7053, 264.607, 263.9703, 263.1259, 259.6385, 
    256.4885, 252.6686, 250.1809, 249.2863, 248.7474, 248.7206, 247.7333, 
    248.9965,
  268.4824, 267.5332, 266.6922, 266.1322, 265.5109, 264.2926, 261.5811, 
    256.7534, 250.8323, 248.7858, 248.097, 247.9361, 247.8722, 247.5554, 
    248.6399,
  268.97, 268.0811, 267.3339, 266.1606, 265.0433, 263.0916, 259.2831, 
    252.8412, 249.2458, 246.8169, 246.2315, 246.8588, 247.1963, 247.9853, 
    247.8836,
  266.6983, 265.4028, 263.253, 259.3777, 258.1079, 255.3893, 254.7502, 
    251.659, 247.559, 242.6547, 241.7149, 245.5303, 246.0513, 246.6784, 
    246.8521,
  258.0059, 258.8195, 258.5302, 257.8868, 256.6859, 253.5025, 257.5994, 
    256.4013, 254.3907, 251.451, 250.5824, 249.6832, 246.4888, 245.4361, 
    242.9893,
  259.5219, 257.4793, 258.5789, 257.8935, 252.911, 254.4139, 255.623, 
    254.7021, 253.4869, 252.5461, 250.5965, 250.9819, 249.437, 243.0071, 
    243.2703,
  265.6495, 261.9388, 259.0667, 257.161, 254.9939, 250.0034, 253.0238, 
    252.7666, 252.481, 252.321, 251.1425, 250.2771, 250.0998, 250.2841, 
    250.6487,
  266.9125, 264.9817, 262.7342, 258.9626, 256.268, 254.6963, 246.9224, 
    249.7817, 249.7729, 248.1743, 249.6371, 249.9652, 250.9657, 252.5072, 
    253.5663,
  266.9763, 265.2303, 263.8553, 261.1294, 256.5816, 256.96, 255.6432, 
    244.8055, 241.5123, 244.0162, 246.4627, 248.9542, 250.9506, 251.7242, 
    253.8277,
  267.4496, 265.9491, 264.5937, 262.5787, 259.8923, 257.7766, 257.4117, 
    258.2398, 252.2645, 248.6028, 246.302, 248.6378, 249.7678, 250.672, 
    252.8029,
  268.1994, 266.7817, 265.5354, 264.1758, 263.3491, 261.8943, 258.3188, 
    254.9035, 251.309, 249.8726, 248.5455, 247.8868, 247.7928, 248.9589, 
    250.9866,
  268.8254, 267.5342, 266.4628, 265.74, 265.1662, 263.3675, 259.9871, 
    253.7122, 250.1109, 248.5167, 247.5579, 247.3777, 247.1825, 248.275, 
    249.1139,
  269.553, 268.6124, 267.8318, 266.633, 265.0303, 262.2306, 257.5836, 
    251.7797, 249.5715, 247.6569, 247.362, 247.8406, 248.0916, 248.4775, 
    248.2801,
  268.7804, 267.6051, 265.9899, 262.2742, 259.0039, 256.6665, 254.893, 
    250.5663, 248.0371, 244.5039, 245.2915, 247.5106, 247.7732, 247.5647, 
    247.999,
  259.0284, 259.8473, 258.0078, 254.7704, 252.0541, 251.1824, 254.2499, 
    254.7914, 255.2475, 251.2113, 249.8004, 250.6264, 248.9603, 245.782, 
    243.0556,
  259.9423, 257.7087, 255.7597, 253.5094, 250.2335, 250.5144, 252.0702, 
    252.7414, 253.5447, 253.6026, 251.1177, 251.5519, 250.1759, 241.3667, 
    238.5403,
  262.9949, 259.3202, 255.9584, 254.2023, 252.5719, 245.3555, 249.6425, 
    250.7464, 251.7484, 253.143, 253.1496, 252.3768, 252.2323, 250.0451, 
    246.4305,
  265.9828, 264.0309, 261.5624, 258.0708, 254.6804, 254.8826, 242.6286, 
    248.5753, 250.1164, 250.2434, 252.5932, 252.9911, 253.2057, 252.3953, 
    249.7578,
  267.2928, 265.5014, 263.6001, 260.8304, 255.2016, 257.19, 257.1932, 
    242.9928, 242.9809, 248.1917, 249.9506, 251.4641, 251.9682, 251.4976, 
    250.6571,
  267.9243, 266.0272, 264.5043, 262.1361, 259.7361, 256.8954, 256.3801, 
    256.1794, 250.2441, 249.9967, 248.6546, 250.4011, 250.9138, 250.5373, 
    250.4019,
  268.5893, 267.0604, 265.4266, 264.1982, 263.5098, 260.4021, 254.8714, 
    252.0904, 250.6156, 249.2694, 248.6583, 248.5815, 248.9998, 248.9175, 
    249.7604,
  269.0281, 267.6465, 266.4735, 265.5531, 263.959, 261.3344, 257.1103, 
    251.5949, 249.6135, 248.1003, 247.8559, 247.7771, 247.9761, 248.6548, 
    249.1576,
  269.356, 268.2973, 267.1055, 264.9839, 262.0266, 258.0993, 253.2444, 
    250.7823, 248.6716, 247.3019, 247.2639, 247.4846, 247.7111, 247.9413, 
    248.2922,
  269.6069, 267.8799, 263.6764, 257.2151, 254.1857, 252.3663, 251.5543, 
    250.3849, 247.5301, 245.2651, 245.3819, 247.2824, 246.9727, 246.884, 
    247.3805,
  257.876, 257.0536, 254.2812, 253.5517, 250.1691, 248.6535, 250.8203, 
    250.7206, 251.7251, 246.5428, 245.4075, 247.9005, 246.9226, 243.8067, 
    241.6829,
  257.71, 255.7431, 254.4021, 251.6137, 247.5431, 245.9989, 248.3129, 
    248.8654, 249.7561, 250.6095, 247.1209, 249.9343, 249.8888, 240.4554, 
    237.8413,
  260.3861, 257.2267, 255.0307, 253.1865, 250.9202, 241.6804, 245.7986, 
    247.677, 247.6981, 248.7203, 249.9335, 249.9665, 249.894, 247.9689, 
    241.7384,
  263.5769, 262.6713, 261.1942, 258.5932, 255.2706, 254.5045, 239.9321, 
    245.9468, 248.2638, 247.3346, 248.4372, 249.2489, 249.5513, 247.9859, 
    244.1102,
  265.8023, 264.7993, 263.9865, 261.3872, 255.3505, 257.1505, 255.599, 
    239.9338, 241.8472, 246.6889, 247.5758, 248.1644, 249.4386, 249.1907, 
    248.5938,
  267.2552, 265.7821, 264.6235, 262.451, 259.176, 255.9548, 255.517, 
    254.4709, 249.5677, 249.4999, 247.1919, 247.948, 248.7904, 249.3092, 
    249.604,
  268.3365, 266.8053, 265.7267, 264.5714, 262.873, 259.4453, 254.596, 
    252.0619, 250.8789, 249.7486, 248.777, 247.5258, 247.0005, 247.1273, 
    248.4106,
  268.7824, 267.8351, 266.8495, 265.5885, 264.079, 261.2432, 256.9369, 
    251.5045, 250.0666, 248.7102, 247.7932, 247.058, 246.1901, 246.3162, 
    247.3087,
  269.2777, 268.4276, 266.7452, 264.2142, 261.2216, 257.3724, 253.6097, 
    251.218, 249.3324, 246.7232, 246.0439, 245.8245, 245.6946, 245.6895, 
    245.1427,
  269.1054, 266.7966, 261.8371, 255.5249, 252.6957, 251.6857, 251.6552, 
    251.0093, 247.1475, 243.0779, 241.7871, 244.7034, 243.8594, 243.7276, 
    244.1755,
  256.6599, 256.5467, 254.8409, 254.6406, 252.9212, 252.2557, 252.4648, 
    251.7065, 251.2259, 246.696, 245.2852, 245.5665, 242.6854, 241.5082, 
    238.638,
  256.7458, 255.4921, 254.2405, 252.3535, 250.1277, 247.5259, 249.7661, 
    249.9189, 250.1143, 249.3074, 244.9404, 247.4422, 247.856, 240.2423, 
    239.0351,
  259.7303, 256.0284, 254.4834, 252.7243, 250.6799, 242.9125, 246.1318, 
    247.786, 247.852, 248.1072, 247.694, 247.7227, 248.468, 248.5647, 243.9123,
  264.0709, 262.3303, 259.6281, 255.9552, 254.2945, 252.2228, 240.8928, 
    245.1656, 246.5321, 245.6478, 245.9555, 247.3484, 248.3038, 247.7635, 
    245.079,
  266.2387, 264.8563, 263.1977, 260.1337, 254.2564, 255.8058, 253.9489, 
    240.1434, 238.1977, 242.3841, 245.1443, 247.0604, 248.2383, 248.0652, 
    247.3827,
  267.0397, 265.6577, 263.9299, 261.3298, 258.3053, 255.4616, 256.2739, 
    255.1662, 249.5353, 245.8868, 243.5443, 246.3338, 248.2595, 248.2523, 
    247.7071,
  268.1464, 266.9281, 265.5539, 264.0707, 262.671, 259.5289, 255.2141, 
    252.7764, 249.2472, 247.3237, 245.55, 245.008, 245.0215, 245.686, 245.8244,
  269.0644, 268.3521, 267.3498, 266.0388, 264.8964, 262.0558, 257.0996, 
    251.6295, 248.5406, 245.6402, 244.4374, 243.9791, 243.3494, 243.9897, 
    245.4905,
  269.329, 268.5735, 267.2836, 265.1455, 263.206, 260.3545, 255.4121, 
    250.7063, 247.3772, 244.0895, 243.6806, 243.6074, 243.5201, 244.5879, 
    246.0986,
  268.4879, 266.2004, 262.9817, 258.1853, 256.5522, 255.072, 252.8244, 
    250.3794, 245.9437, 240.8761, 240.6544, 243.9499, 244.3354, 245.4191, 
    247.2434,
  257.6534, 257.1696, 256.0907, 256.0968, 256.1346, 255.6765, 256.2966, 
    256.2422, 256.3652, 253.7203, 253.0426, 252.7678, 250.9005, 249.8198, 
    246.8205,
  258.6379, 257.2559, 256.6555, 255.7425, 254.3215, 252.5266, 253.8782, 
    254.2753, 254.5867, 253.8321, 251.7958, 252.3161, 251.0191, 244.9118, 
    242.8307,
  261.5189, 258.3492, 257.2446, 256.2082, 254.3726, 247.6956, 249.7632, 
    251.0965, 251.3792, 251.9871, 251.3622, 250.7609, 250.4125, 248.9603, 
    244.751,
  265.0075, 263.1511, 260.0472, 256.7011, 255.4361, 253.3163, 244.8342, 
    247.7593, 247.9833, 247.6109, 248.7502, 248.898, 249.2532, 248.9196, 
    246.5193,
  265.9355, 264.0772, 262.2758, 258.8134, 254.7124, 254.9444, 254.2378, 
    241.2036, 238.9444, 242.9063, 245.8715, 247.9547, 248.2251, 248.1255, 
    248.5173,
  266.5632, 265.0357, 263.1125, 260.5689, 257.4915, 255.0435, 256.0384, 
    255.5443, 248.9308, 244.7469, 242.6082, 245.1721, 246.0486, 246.3783, 
    246.4744,
  268.0515, 266.3745, 264.7047, 263.0196, 261.6094, 258.8288, 254.6888, 
    251.3848, 247.3441, 246.1, 244.5679, 244.1575, 244.3878, 244.6586, 
    244.6558,
  270.2744, 268.5372, 266.9242, 265.6774, 264.5819, 261.5216, 256.4971, 
    250.9706, 248.0181, 246.5921, 245.5253, 245.0445, 244.1939, 243.9906, 
    245.3907,
  271.3337, 270.2887, 269.3305, 267.5347, 264.682, 260.3914, 255.2283, 
    251.5913, 249.6163, 248.596, 248.0809, 247.8637, 247.0867, 247.2299, 
    247.2598,
  270.8653, 269.9562, 268.1028, 262.7797, 257.9006, 254.7256, 252.8739, 
    252.4314, 251.5233, 249.8307, 250.2469, 250.8237, 249.9356, 249.3598, 
    249.0487,
  260.0637, 260.317, 258.8404, 258.3915, 257.5928, 257.3151, 260.4439, 
    261.7486, 262.6024, 260.7192, 261.2584, 262.7766, 261.4214, 260.1268, 
    257.759,
  260.6817, 260.7257, 259.9838, 259.9689, 257.3117, 255.1311, 255.954, 
    259.2961, 260.9457, 261.5568, 260.3261, 261.877, 260.8979, 256.3554, 
    254.2461,
  264.7346, 262.4854, 260.7064, 260.48, 259.0038, 252.5278, 253.7742, 
    254.1523, 256.6237, 258.8573, 259.6022, 259.7994, 259.3892, 257.7575, 
    254.0407,
  267.3033, 266.4411, 263.5952, 260.18, 259.7365, 258.4846, 250.1878, 
    251.7533, 251.16, 253.1218, 255.6697, 256.0696, 256.0179, 254.5565, 
    252.3663,
  267.7947, 266.9154, 266.0499, 262.4676, 258.749, 259.0016, 258.3595, 
    245.101, 242.8686, 248.2848, 251.176, 253.0632, 253.7927, 253.0495, 
    252.0669,
  268.9783, 268.1241, 266.5815, 264.9035, 259.7155, 257.214, 257.5908, 
    256.7145, 248.8318, 246.6227, 246.0754, 249.0799, 251.0614, 251.3829, 
    250.893,
  270.7299, 269.8989, 268.1954, 267.5406, 266.1744, 263.0154, 256.8508, 
    253.5522, 249.7066, 247.5318, 245.476, 246.2766, 247.4314, 248.2367, 
    248.9575,
  271.768, 271.0946, 269.5869, 267.7655, 266.1647, 264.7244, 261.4221, 
    256.0359, 254.797, 251.0467, 247.9198, 246.4197, 245.2865, 245.0201, 
    248.1645,
  271.21, 270.357, 268.4422, 265.3167, 263.2051, 260.738, 258.0819, 256.3715, 
    255.0648, 254.2804, 252.2738, 249.2388, 247.1624, 246.5938, 246.8565,
  268.703, 266.8038, 263.5915, 260.3408, 259.0716, 258.0712, 256.9851, 
    255.4743, 252.586, 250.319, 253.4517, 253.4742, 250.3395, 248.8098, 
    248.1336,
  261.1028, 264.3786, 261.0157, 260.9495, 260.6249, 257.4952, 258.5872, 
    261.2825, 262.0763, 258.925, 259.0091, 263.4232, 260.9319, 261.3927, 
    258.949,
  262.5479, 264.4611, 262.4197, 261.8893, 260.7649, 256.5119, 256.4279, 
    258.7471, 262.7434, 263.0523, 260.4877, 264.2518, 263.7233, 260.4979, 
    258.5842,
  267.0847, 266.8354, 264.1225, 262.2155, 261.8356, 255.2746, 255.5515, 
    255.6326, 256.5225, 260.0204, 262.7573, 263.2587, 263.6512, 263.0572, 
    259.8454,
  269.3189, 270.5638, 269.6831, 262.4533, 262.5017, 261.7285, 251.1071, 
    254.1203, 253.6411, 253.2225, 257.4241, 260.5916, 261.747, 261.4439, 
    259.9188,
  269.7968, 270.5943, 270.8484, 266.8501, 261.391, 262.3037, 260.5976, 
    245.667, 246.0316, 249.8499, 251.1335, 255.8334, 258.1954, 259.6416, 
    259.5418,
  270.4972, 271.4072, 270.8634, 267.8438, 264.9358, 263.5155, 260.4861, 
    258.7508, 250.8205, 248.5162, 247.2448, 249.8435, 253.4752, 256.3217, 
    257.4745,
  271.0858, 271.5854, 270.8914, 268.9676, 267.8754, 266.0789, 260.295, 
    256.353, 254.4741, 250.6452, 247.5655, 246.6173, 248.0246, 250.8229, 
    254.0832,
  271.3492, 271.6323, 270.3814, 267.6031, 266.2973, 264.3627, 259.7764, 
    254.9478, 255.394, 254.2371, 251.4736, 246.0122, 245.2981, 246.6249, 
    249.4339,
  270.7331, 270.946, 269.3089, 266.1959, 263.1867, 259.0613, 255.2632, 
    252.7742, 251.0909, 250.0568, 249.1961, 249.0681, 247.0579, 245.5893, 
    245.4096,
  269.8059, 269.4997, 266.5637, 261.4491, 257.5835, 253.6455, 252.4355, 
    252.0262, 249.2615, 246.7694, 249.4261, 249.4059, 247.0037, 245.2497, 
    245.0282,
  260.8829, 261.9394, 261.1346, 258.5712, 257.4577, 251.0935, 253.0556, 
    256.223, 260.2246, 258.897, 256.1236, 259.6638, 259.9738, 257.1188, 
    256.2936,
  261.9608, 261.804, 261.1706, 261.8146, 259.0328, 249.2265, 251.6654, 
    252.9536, 256.6494, 258.8356, 259.7083, 263.4425, 263.7397, 258.3134, 
    256.315,
  265.4524, 263.1298, 262.4997, 263.0119, 262.1482, 252.135, 250.0246, 
    251.0629, 252.3555, 253.5127, 256.9505, 259.738, 261.7581, 262.6728, 
    260.9633,
  268.4407, 267.9208, 267.3, 264.5869, 264.1224, 262.5852, 249.7851, 
    250.3957, 251.8368, 250.4225, 251.412, 255.6365, 257.6915, 258.8285, 
    258.3204,
  269.6594, 269.1191, 269.1233, 267.6697, 264.0604, 264.3884, 262.4544, 
    246.0444, 243.9348, 247.7994, 248.4974, 250.4386, 253.7933, 255.8815, 
    257.6169,
  270.4543, 270.1154, 269.6102, 268.6727, 266.093, 263.7835, 262.9648, 
    261.7061, 253.9722, 248.8724, 245.5997, 247.7858, 249.1303, 251.5937, 
    254.2268,
  270.8652, 270.8497, 270.52, 269.8833, 269.2615, 267.2118, 261.4087, 
    258.408, 255.5772, 253.4957, 248.5114, 246.2481, 246.4833, 247.5666, 
    250.2276,
  271.2932, 271.3318, 270.9859, 270.0933, 269.4631, 268.0984, 261.4778, 
    257.0187, 254.8069, 254.274, 251.1797, 245.9965, 244.6948, 245.6359, 
    247.4842,
  271.481, 271.661, 271.4068, 270.1234, 268.2069, 265.0509, 259.2281, 
    255.1774, 253.3228, 251.425, 250.0747, 246.9956, 244.5953, 244.7572, 
    245.9229,
  271.7939, 271.7543, 270.7791, 266.621, 262.4282, 259.6477, 256.9182, 
    255.2092, 251.8687, 250.1677, 251.597, 247.492, 244.0579, 243.7696, 
    244.781,
  260.6008, 260.3606, 259.9613, 260.2395, 259.0491, 252.9159, 251.4477, 
    252.6375, 257.7824, 260.132, 260.2067, 261.5946, 260.2161, 253.9372, 
    253.4044,
  264.4338, 261.0062, 260.8837, 261.1497, 259.0976, 251.8181, 250.9502, 
    250.9923, 253.196, 256.8785, 259.9229, 262.7326, 261.9814, 259.0647, 
    255.5632,
  267.576, 263.058, 261.5318, 262.3688, 260.7592, 253.9361, 250.4972, 
    249.6007, 250.5345, 251.969, 253.9505, 256.5417, 257.6434, 258.0143, 
    256.0576,
  270.3281, 268.4039, 265.3904, 263.5663, 263.0084, 260.9738, 253.5386, 
    249.9283, 250.4224, 249.3041, 251.5182, 252.518, 252.8056, 252.7045, 
    252.406,
  271.227, 270.3535, 268.5625, 266.048, 263.8501, 263.6195, 262.212, 
    255.2642, 253.777, 248.6871, 248.6259, 249.9695, 250.8402, 250.975, 
    251.3713,
  271.8091, 271.3784, 270.0891, 267.8949, 265.1209, 263.9411, 263.8776, 
    263.3947, 257.708, 252.06, 247.1785, 247.8608, 247.9474, 248.8828, 
    250.1562,
  272.1795, 272.0506, 271.4099, 269.5378, 267.8481, 266.3207, 263.8125, 
    261.1723, 257.0714, 252.5327, 248.9272, 247.3535, 246.1143, 246.6575, 
    249.157,
  272.4298, 272.387, 271.9955, 270.6154, 269.1089, 268.3754, 264.9655, 
    259.6112, 254.4989, 252.2401, 249.3826, 247.6537, 244.4574, 245.8636, 
    248.7314,
  272.4262, 272.5506, 272.2674, 271.0751, 269.7483, 267.873, 263.7225, 
    257.8506, 253.3802, 251.8234, 248.9926, 247.8916, 243.7197, 245.4383, 
    248.178,
  272.3618, 272.3305, 271.6823, 269.2392, 267.5069, 265.8585, 261.493, 
    255.6307, 251.9318, 250.3427, 249.3547, 246.5162, 243.202, 244.3683, 
    247.105,
  266.7954, 264.8641, 261.2032, 260.1254, 256.5337, 255.6778, 257.3259, 
    259.2567, 260.8551, 259.9248, 259.7749, 259.7748, 258.81, 255.3881, 
    253.1534,
  267.5334, 265.2255, 261.2124, 259.3311, 254.4268, 253.4218, 256.2536, 
    258.2867, 260.0592, 261.2058, 261.0555, 261.8406, 260.4839, 251.53, 
    252.5892,
  269.3399, 266.668, 262.6329, 260.882, 256.8801, 250.4463, 253.7244, 
    255.6661, 257.8669, 258.6987, 259.4218, 259.4116, 257.3853, 255.6662, 
    248.762,
  270.8094, 269.4923, 265.1404, 261.766, 259.5809, 257.7723, 250.7223, 
    253.4878, 254.6753, 255.454, 256.249, 254.9161, 253.8412, 252.1647, 
    249.2646,
  271.7874, 270.6711, 267.425, 264.464, 260.4601, 260.2717, 258.3009, 
    249.9441, 250.0451, 251.6951, 253.1485, 253.1571, 252.3929, 250.8875, 
    249.8934,
  272.1921, 271.4194, 268.4739, 266.0086, 262.0763, 260.8713, 260.6358, 
    260.7253, 258.3102, 253.6713, 250.7855, 250.7553, 249.6125, 248.5384, 
    249.1073,
  272.6105, 272.2195, 269.8142, 267.6233, 265.4202, 263.9022, 261.5412, 
    261.1909, 257.9514, 253.9897, 251.383, 249.1882, 247.2914, 247.0613, 
    248.9023,
  272.8763, 272.5352, 270.6331, 268.7399, 267.1568, 266.2077, 263.3004, 
    259.4962, 255.7039, 252.6179, 250.1147, 247.6718, 244.7015, 246.6852, 
    249.1173,
  273.1739, 272.9634, 271.4288, 269.5934, 268.4226, 266.5982, 262.8102, 
    258.5883, 253.9947, 251.1695, 248.5868, 245.9017, 243.7928, 246.0191, 
    248.4309,
  273.1314, 272.8669, 271.4553, 268.1433, 265.3489, 265.0621, 261.9369, 
    256.1927, 251.4903, 249.2096, 247.2871, 245.0699, 243.2149, 245.11, 
    247.9552,
  268.0684, 267.3236, 266.2241, 264.2011, 257.6318, 251.5071, 255.0965, 
    257.4162, 258.8625, 256.2567, 256.0692, 255.6537, 254.6039, 253.1459, 
    250.3564,
  268.201, 267.5345, 266.5482, 262.4604, 255.0045, 249.7355, 253.1128, 
    256.6039, 259.0661, 259.2827, 258.1435, 258.2502, 256.8552, 251.2782, 
    250.5759,
  269.2666, 267.8542, 266.0331, 262.11, 257.129, 248.2511, 251.6671, 
    255.5246, 258.8327, 260.393, 260.3261, 259.3636, 258.1381, 256.5537, 
    252.783,
  270.5854, 270.0132, 267.4551, 262.0438, 259.7654, 258.6317, 249.7322, 
    254.856, 257.3658, 258.757, 258.9697, 257.7708, 256.8396, 254.991, 
    251.6607,
  271.0164, 270.5996, 268.6869, 263.5178, 258.0506, 259.9889, 259.8188, 
    249.6078, 249.9033, 255.0181, 255.9946, 255.4467, 255.0093, 253.7527, 
    252.2014,
  271.7444, 270.8727, 268.3725, 264.4334, 259.1734, 257.6871, 260.5975, 
    260.1467, 257.2342, 255.0995, 253.5127, 253.3602, 253.0253, 252.3941, 
    251.2242,
  272.2029, 271.1333, 268.4575, 265.8225, 264.4048, 262.7538, 260.3662, 
    258.9084, 256.2635, 254.6629, 252.8003, 251.6533, 250.7379, 250.5664, 
    250.0114,
  272.4822, 271.1324, 268.6963, 267.3414, 266.6529, 264.1864, 259.0387, 
    256.8868, 254.3798, 253.0125, 250.8612, 249.6407, 247.6063, 248.8622, 
    249.3098,
  272.471, 271.1118, 269.2062, 268.292, 266.5302, 262.4503, 257.384, 255.489, 
    252.2037, 250.2068, 248.5372, 247.2088, 245.4076, 247.7276, 248.0648,
  272.3849, 270.9058, 268.772, 264.8286, 260.2728, 259.0836, 255.7056, 
    253.504, 250.2086, 247.7431, 246.4589, 246.0067, 244.3046, 246.3254, 
    247.3923,
  269.6004, 269.142, 268.5959, 268.0669, 267.2488, 265.1859, 262.7436, 
    260.9488, 259.0965, 255.6682, 255.1961, 255.3326, 254.2891, 254.108, 
    252.3644,
  269.7783, 269.3154, 268.5876, 267.5515, 265.2092, 259.2639, 258.0577, 
    256.8094, 256.7891, 256.4044, 256.0789, 257.2599, 256.8693, 252.4637, 
    251.0113,
  270.3182, 269.2735, 267.5585, 265.8639, 262.314, 254.9964, 256.3411, 
    257.1928, 256.2166, 256.6801, 257.2454, 257.856, 258.0792, 257.3734, 
    254.2838,
  270.8723, 269.7661, 267.3135, 264.2696, 261.7995, 258.3276, 251.8291, 
    254.5012, 254.1536, 255.1264, 256.0966, 257.3326, 258.2644, 257.7371, 
    254.7972,
  270.2425, 268.749, 267.2075, 263.9149, 261.3718, 260.9544, 259.4833, 
    249.2739, 245.9563, 253.3617, 255.6794, 257.1024, 258.0936, 257.4458, 
    255.4237,
  269.9822, 268.3296, 266.5009, 264.2281, 261.7514, 260.0423, 260.4567, 
    259.248, 256.5026, 254.9287, 255.1195, 256.6739, 257.1214, 256.5045, 
    255.2702,
  269.8946, 268.5143, 266.9819, 265.2266, 263.6756, 261.162, 258.5153, 
    257.8963, 256.3833, 256.0569, 255.8008, 255.9288, 255.7281, 255.2304, 
    254.5512,
  269.9018, 268.6573, 267.1882, 265.6965, 263.9609, 261.169, 257.0237, 
    256.0326, 255.0755, 254.9141, 254.7238, 254.5823, 254.1345, 254.1442, 
    253.481,
  269.6904, 268.209, 266.4523, 264.1335, 261.801, 258.3135, 255.1885, 
    254.1011, 253.0759, 252.8749, 252.8521, 252.6915, 252.0486, 251.7924, 
    249.617,
  269.0289, 266.8565, 263.5863, 258.2561, 255.8964, 255.6517, 253.8161, 
    252.579, 251.0765, 250.1797, 250.1692, 250.5565, 249.2942, 248.7699, 
    247.8147,
  265.4997, 263.6583, 261.6736, 261.3554, 261.5286, 258.2263, 256.3366, 
    256.5118, 257.5844, 257.493, 257.3208, 257.9751, 258.3494, 259.1495, 
    258.6077,
  265.481, 263.7651, 261.7453, 261.1088, 259.9757, 257.215, 255.3384, 
    253.4409, 254.9182, 256.2061, 255.7042, 257.2585, 256.572, 252.2933, 
    255.5111,
  268.5437, 264.3391, 262.0826, 261.1472, 260.376, 254.3178, 254.9925, 
    253.866, 254.5771, 255.7491, 256.8998, 257.4868, 257.2721, 257.4859, 
    256.6911,
  270.3712, 268.8553, 266.3455, 262.3069, 260.8351, 259.2595, 251.4593, 
    252.4354, 254.073, 255.4193, 256.6281, 257.8134, 257.5404, 257.6867, 
    256.3897,
  270.6061, 268.8571, 267.1792, 263.7752, 260.3475, 259.2908, 258.5996, 
    246.8006, 247.9316, 254.5833, 256.3479, 257.1236, 258.2039, 257.998, 
    256.8336,
  270.7648, 268.9734, 266.7991, 264.3627, 261.1275, 258.2655, 257.4066, 
    257.0528, 255.9131, 256.6956, 256.1032, 257.3052, 258.0309, 257.4934, 
    256.43,
  270.8494, 269.0946, 266.8255, 264.5434, 262.8469, 259.0115, 255.9612, 
    255.5643, 255.9863, 257.2596, 257.5019, 257.5804, 257.4677, 256.8121, 
    256.1771,
  270.7877, 268.9775, 266.3166, 263.6406, 261.7796, 259.1285, 255.0981, 
    254.4692, 254.2908, 255.4678, 256.6198, 256.9608, 256.5858, 256.0437, 
    255.4768,
  270.7019, 268.7552, 265.7413, 262.2308, 259.2494, 255.9234, 254.2968, 
    253.6871, 253.2197, 253.1316, 254.1394, 254.4551, 253.9922, 253.4067, 
    251.2995,
  270.4047, 268.0675, 264.1531, 257.4339, 253.7102, 253.2267, 253.2097, 
    252.9708, 251.8914, 251.1344, 251.2495, 252.0951, 251.6897, 251.2161, 
    250.0843,
  267.3148, 264.0945, 260.5145, 258.6043, 257.9495, 254.086, 253.6156, 
    253.0169, 254.6548, 254.4919, 255.3802, 256.9027, 256.7657, 255.902, 
    256.0283,
  268.7187, 264.6782, 262.2138, 258.7942, 257.1547, 252.6349, 253.6649, 
    252.7318, 254.2753, 256.2349, 256.2526, 258.3516, 258.5232, 252.9321, 
    255.3599,
  270.3004, 265.8877, 263.4634, 259.4316, 258.7805, 250.4047, 253.2193, 
    254.3057, 255.7507, 257.1288, 258.2225, 259.0155, 258.8682, 258.4095, 
    259.3749,
  271.844, 270.362, 267.7935, 261.1361, 260.2521, 257.0864, 249.4837, 
    252.5665, 255.4727, 257.2701, 258.5659, 258.9848, 258.923, 258.5425, 
    257.6621,
  272.6513, 270.7925, 268.9156, 264.3446, 258.6709, 257.3973, 256.6653, 
    245.9881, 249.8818, 256.4369, 257.8448, 258.3895, 258.5911, 257.9807, 
    257.5894,
  273.4034, 271.9113, 269.3595, 265.951, 261.1537, 256.8413, 255.753, 
    255.0049, 254.9531, 256.8237, 256.3205, 257.6236, 257.9473, 257.4868, 
    256.8775,
  273.9173, 272.7036, 270.6903, 267.1986, 264.2336, 259.1548, 254.5935, 
    253.3178, 253.6246, 255.1006, 255.2874, 256.03, 256.3316, 256.1486, 
    255.8095,
  274.347, 273.3325, 271.4576, 268.0238, 264.6183, 260.1163, 253.7461, 
    252.4168, 251.7589, 252.5846, 253.304, 253.7927, 253.7665, 253.9407, 
    253.5026,
  274.5925, 273.6701, 272.283, 269.0248, 264.9224, 257.5329, 253.5311, 
    251.8047, 250.5404, 249.877, 250.6917, 251.1137, 251.445, 251.3886, 
    250.4163,
  274.4341, 273.4126, 272.1496, 268.7931, 262.2628, 254.8345, 252.682, 
    251.8191, 249.1947, 247.0312, 247.6441, 249.6714, 249.7101, 250.1694, 
    250.5863,
  272.6105, 270.2405, 265.0441, 259.1518, 253.7956, 249.9952, 249.4255, 
    250.7493, 255.5508, 255.2104, 256.0825, 256.8036, 254.5312, 253.3158, 
    250.4442,
  272.5873, 269.7185, 264.2938, 257.5938, 252.2655, 249.1004, 250.1599, 
    251.1345, 254.8138, 256.4559, 256.1455, 258.7286, 258.0419, 251.57, 
    247.7076,
  272.3963, 269.356, 263.8915, 258.5716, 255.3537, 247.6354, 250.1719, 
    252.7014, 255.7138, 257.1852, 257.8807, 258.0112, 257.1393, 255.7388, 
    253.7176,
  273.0765, 270.6021, 265.9456, 260.344, 258.984, 255.2781, 246.6548, 
    252.1047, 254.6974, 256.3559, 257.7632, 257.5809, 257.0649, 256.5201, 
    256.4238,
  273.6658, 271.0897, 268.1408, 262.6125, 258.8972, 258.2281, 256.5176, 
    246.3942, 250.1321, 254.2498, 256.3485, 257.3075, 257.8797, 257.4579, 
    256.9706,
  273.9759, 271.636, 268.4533, 263.7936, 259.4553, 257.49, 257.0168, 
    255.2696, 252.9272, 254.8535, 254.3011, 256.1914, 256.7373, 256.535, 
    256.4321,
  273.9793, 272.0229, 269.1105, 265.079, 261.9019, 257.9943, 255.0377, 
    252.8041, 252.1232, 252.683, 252.9138, 254.5011, 255.0123, 255.4888, 
    255.6418,
  273.7067, 271.8667, 269.5683, 266.1689, 263.6786, 259.8467, 254.1556, 
    252.3784, 250.6851, 250.3177, 250.7938, 251.8692, 252.5606, 253.7428, 
    253.8062,
  273.1565, 271.744, 269.8755, 266.8398, 264.05, 258.2624, 253.5531, 
    251.8285, 250.0232, 249.2187, 249.7525, 250.7105, 251.4075, 252.5653, 
    252.9431,
  272.5478, 271.2395, 269.1297, 265.233, 260.5634, 255.7888, 253.601, 
    252.3272, 250.1458, 248.2337, 248.8574, 251.2019, 251.8091, 252.8015, 
    253.2278,
  260.4928, 257.0429, 254.8857, 254.102, 253.1862, 252.6977, 253.7801, 
    250.2335, 251.8498, 249.3235, 250.9195, 252.9305, 251.6905, 249.9854, 
    248.6843,
  260.3258, 257.6094, 256.5923, 255.0678, 253.7612, 252.5028, 254.0056, 
    252.0898, 252.5378, 251.7066, 251.4509, 254.0907, 253.6183, 247.0001, 
    246.2013,
  262.5733, 259.1353, 258.1833, 257.8946, 256.7807, 249.4965, 253.2675, 
    254.1357, 255.5548, 254.5593, 254.432, 254.6806, 253.8349, 252.2401, 
    249.9038,
  265.6536, 264.0303, 261.5507, 259.3354, 259.6651, 257.7146, 251.022, 
    254.0033, 255.4636, 256.3404, 257.0803, 256.4823, 255.1488, 254.197, 
    252.0966,
  267.0149, 265.8542, 264.1914, 260.9657, 259.6871, 259.3008, 258.0548, 
    248.175, 250.4137, 255.21, 256.4853, 257.7396, 257.8399, 256.895, 255.3672,
  267.5959, 266.358, 264.6427, 262.1827, 259.6617, 257.957, 257.6263, 
    256.4494, 255.286, 256.1224, 255.4207, 256.4841, 257.3096, 257.4784, 
    256.7832,
  268.2599, 267.2505, 266.0003, 264.1964, 262.4747, 258.3703, 256.5636, 
    255.6758, 255.278, 255.6352, 256.4518, 256.4521, 256.6992, 257.1162, 
    257.2582,
  268.732, 267.8212, 266.3664, 264.9851, 263.2563, 259.6299, 256.5356, 
    255.6972, 254.9321, 255.015, 256.0063, 257.1942, 256.8902, 257.2568, 
    257.3638,
  268.6311, 267.4252, 265.5807, 263.8882, 261.6197, 258.5783, 256.9807, 
    256.1588, 255.2975, 254.9476, 254.9538, 256.8583, 257.7205, 257.9196, 
    257.9947,
  267.7841, 265.7376, 263.171, 260.4626, 258.5331, 258.0233, 257.1341, 
    257.169, 255.326, 254.2072, 254.1255, 255.2068, 257.155, 258.324, 258.4791,
  260.2317, 259.2618, 259.1632, 259.0428, 255.383, 252.1691, 251.9708, 
    251.1579, 251.4645, 247.2258, 246.7727, 250.546, 251.239, 251.3111, 
    252.352,
  261.0541, 259.3742, 259.6942, 258.9018, 256.5041, 252.6372, 253.3419, 
    251.996, 252.965, 250.6103, 247.1888, 251.2306, 253.6097, 247.819, 
    249.0595,
  265.5073, 262.3291, 260.4585, 259.7549, 258.8957, 250.8978, 253.381, 
    253.6601, 254.443, 253.719, 251.9293, 251.5573, 253.1019, 253.7202, 
    252.181,
  268.0821, 266.8173, 264.1206, 260.2559, 259.6622, 257.8626, 250.9774, 
    252.728, 254.676, 253.9127, 254.701, 252.7367, 252.4388, 253.5168, 
    252.3873,
  268.5608, 267.344, 265.671, 261.8581, 259.19, 257.8902, 257.1445, 247.1492, 
    249.1362, 253.3212, 253.4452, 254.0848, 252.8575, 253.0676, 253.2935,
  268.6194, 267.4917, 265.6865, 263.0172, 260.5025, 257.1999, 256.1515, 
    254.9999, 254.4398, 255.7369, 251.4342, 254.1438, 254.5739, 253.0678, 
    252.7811,
  268.5, 267.0482, 265.7853, 263.6333, 261.8162, 257.7519, 255.7011, 
    253.8335, 253.8724, 255.9527, 254.843, 254.2915, 253.9422, 253.1311, 
    252.6355,
  267.7762, 266.13, 264.0195, 262.4899, 260.5859, 257.9325, 255.5735, 
    253.4086, 252.1864, 253.538, 256.2678, 255.3748, 253.7567, 254.1608, 
    252.9329,
  266.8823, 264.8945, 262.7061, 259.9534, 257.3691, 255.3783, 255.5378, 
    253.9195, 252.0081, 252.0946, 253.2535, 256.8018, 256.0643, 254.9733, 
    254.3022,
  264.9372, 262.7198, 259.3931, 255.1453, 253.3392, 253.541, 253.4312, 
    254.6595, 251.4506, 250.2411, 251.093, 254.0375, 257.1607, 257.2508, 
    256.113,
  259.9323, 258.0286, 257.9573, 257.5659, 252.8399, 249.8221, 249.4607, 
    250.3635, 251.2419, 249.7533, 249.4332, 249.6688, 248.3231, 248.4315, 
    248.6284,
  259.7163, 258.3471, 259.1657, 258.3513, 255.6008, 248.431, 249.201, 
    249.5708, 250.8479, 251.6515, 250.0076, 251.2419, 252.7856, 248.1417, 
    247.6555,
  264.7288, 259.5027, 257.8497, 258.1735, 257.6359, 248.9049, 250.1537, 
    250.4523, 251.1623, 251.5043, 252.028, 252.0883, 252.6983, 253.9364, 
    252.431,
  267.2568, 265.2956, 262.1996, 257.7621, 257.9976, 255.6531, 247.7099, 
    250.208, 251.6056, 253.6937, 253.6251, 253.1484, 252.93, 254.127, 253.4311,
  267.4121, 265.7039, 263.5561, 259.5856, 257.1547, 256.0654, 254.8026, 
    243.1539, 245.1255, 253.4012, 253.7848, 252.7683, 252.2895, 253.7347, 
    255.2827,
  266.8679, 265.2704, 263.126, 260.4117, 257.8018, 255.2841, 254.7065, 
    252.7946, 252.6556, 254.7213, 252.8936, 251.75, 251.0883, 253.1715, 
    254.3533,
  266.4552, 264.8209, 263.0825, 260.8705, 258.9745, 255.0035, 254.1512, 
    252.8276, 253.4408, 255.2797, 254.2885, 251.6493, 249.7871, 251.0855, 
    253.3806,
  265.5226, 263.9659, 261.8385, 259.901, 257.4732, 254.2024, 253.5017, 
    252.794, 252.8562, 254.5388, 254.762, 252.0531, 249.9114, 250.6672, 
    251.8414,
  264.9274, 262.8903, 260.5933, 257.656, 253.635, 251.6423, 252.3876, 
    252.6877, 252.3586, 253.7372, 254.5084, 253.4449, 250.2374, 250.3206, 
    251.0336,
  263.2221, 260.4486, 257.0421, 251.9881, 250.2667, 249.7409, 250.145, 
    252.5961, 251.1779, 251.4543, 252.7206, 254.7315, 252.6793, 250.4191, 
    250.5375,
  257.5096, 256.4904, 254.9157, 253.7497, 252.1938, 249.686, 249.2123, 
    248.4848, 248.8853, 247.452, 250.5477, 250.9885, 248.8837, 248.2347, 
    247.8729,
  257.2989, 256.1847, 256.1986, 254.952, 253.1131, 246.585, 247.5662, 
    247.7424, 248.2111, 250.4003, 251.2053, 252.1982, 252.3929, 249.4101, 
    246.5345,
  260.6709, 256, 256.3987, 256.1751, 255.0656, 246.0591, 248.6577, 248.2801, 
    247.9506, 249.9515, 252.079, 252.5382, 252.4292, 252.0003, 249.3355,
  265.4711, 263.6267, 260.0475, 255.7412, 257.2442, 254.6817, 245.2756, 
    249.7818, 250.5431, 251.8032, 253.2254, 254.0501, 253.7027, 253.4561, 
    252.0795,
  266.5616, 264.9236, 263.0957, 257.3597, 255.8289, 255.816, 254.5779, 
    242.0566, 244.8782, 253.4646, 254.4078, 253.8617, 253.7065, 253.9096, 
    254.4082,
  266.601, 265.2566, 263.3596, 259.5597, 257.3808, 255.0361, 254.6508, 
    253.6838, 252.9305, 253.4782, 251.9936, 251.9008, 252.2735, 253.0719, 
    253.756,
  266.9267, 265.6037, 263.9858, 261.7754, 259.7762, 254.5937, 253.208, 
    252.6735, 252.6579, 252.8024, 251.6703, 250.1073, 249.845, 251.1727, 
    252.7704,
  266.6733, 265.4044, 263.6756, 261.7723, 259.1795, 254.4437, 252.6246, 
    252.1361, 251.1632, 250.9367, 250.1812, 249.8935, 249.8587, 251.3046, 
    252.4534,
  266.7959, 265.1214, 263.2409, 260.6233, 256.2955, 253.3451, 252.0969, 
    252.3026, 251.1009, 250.2716, 249.2704, 249.965, 249.7458, 251.4332, 
    252.4563,
  266.5054, 264.4321, 261.7273, 257.3413, 254.2587, 253.0437, 251.8027, 
    254.0704, 251.4995, 247.9727, 246.2463, 248.6273, 249.76, 251.3884, 
    252.1016,
  255.5849, 254.3754, 252.6094, 252.1331, 249.5121, 246.0518, 247.6224, 
    248.2118, 249.0732, 247.3857, 249.0543, 250.9289, 250.0808, 250.6137, 
    251.1771,
  255.3855, 254.7768, 254.519, 254.2034, 252.2567, 248.4579, 249.1626, 
    248.952, 249.6724, 249.4713, 249.3003, 251.2552, 252.0654, 249.0869, 
    249.0202,
  261.5797, 257.3669, 256.2642, 256.9789, 256.4771, 249.677, 250.4342, 
    250.0371, 249.3774, 250.0929, 251.2487, 252.0484, 252.2091, 252.0944, 
    250.1472,
  267.6144, 266.7075, 264.4661, 259.9735, 260.4194, 258.1644, 251.2573, 
    251.8939, 251.6136, 252.0494, 252.665, 253.0987, 253.0086, 252.6806, 
    251.2375,
  269.3074, 269.0839, 268.725, 264.3362, 262.8246, 261.3437, 259.2994, 
    249.2265, 248.3356, 253.5517, 254.5389, 254.3094, 254.0201, 254.0206, 
    253.7468,
  270.1841, 270.215, 269.3965, 266.6416, 265.3495, 262.6059, 260.17, 
    257.7978, 255.2647, 254.0169, 253.5516, 253.7388, 253.646, 253.8499, 
    254.0776,
  271.286, 270.9958, 269.9152, 267.7828, 266.4301, 262.6122, 258.9761, 
    256.8761, 254.5478, 253.132, 251.9738, 252.004, 252.7434, 252.9899, 
    253.7367,
  271.952, 270.9496, 269.0649, 267.2964, 265.0164, 261.2866, 257.7823, 
    255.5515, 253.537, 252.0328, 250.981, 250.2229, 250.4645, 251.5866, 
    252.5968,
  271.9188, 270.2704, 268.2852, 265.7385, 261.8456, 258.7958, 255.944, 
    254.6371, 252.9165, 251.1662, 249.8905, 249.0987, 249.3038, 250.3775, 
    251.5421,
  271.2065, 269.0205, 266.4026, 262.4601, 259.3766, 256.8794, 253.7412, 
    253.3618, 252.0457, 249.8206, 248.2691, 248.2252, 248.1487, 249.1339, 
    250.3624,
  259.8616, 259.5746, 259.2329, 258.7689, 256.1921, 252.1507, 251.5468, 
    250.4335, 249.9993, 247.0077, 247.7906, 248.8228, 247.127, 247.7685, 
    246.6423,
  262.0175, 261.3744, 261.3781, 261.5707, 258.8966, 256.8044, 256.168, 
    255.4172, 253.7272, 252.6473, 252.2988, 252.5975, 251.9877, 248.9668, 
    248.135,
  267.786, 265.5675, 265.6422, 266.5313, 263.9372, 261.4029, 259.274, 
    256.7621, 255.7775, 255.0943, 254.095, 254.54, 253.5875, 252.5898, 
    251.0639,
  269.6788, 270.2161, 270.9695, 269.5682, 267.6479, 264.41, 257.7104, 
    257.0458, 257.002, 256.3714, 256.2147, 255.3088, 254.4449, 254.7082, 
    253.7466,
  270.1954, 271.4547, 272.0505, 269.7362, 266.2424, 263.492, 261.1705, 
    252.2839, 251.7184, 255.9931, 256.4636, 255.7561, 255.1601, 254.7514, 
    254.6664,
  271.943, 272.5737, 271.6406, 268.2107, 265.5989, 262.1802, 260.7899, 
    257.9402, 254.964, 252.075, 252.7018, 253.0324, 253.128, 253.5552, 
    254.0367,
  273.2203, 272.639, 270.4864, 267.5544, 265.7366, 261.4031, 257.9338, 
    255.067, 252.9132, 250.7482, 250.1295, 250.098, 250.4616, 251.0681, 
    251.983,
  273.0005, 271.1657, 268.8864, 266.2813, 262.9839, 256.5736, 252.4647, 
    250.7207, 250.214, 249.8741, 249.6827, 249.5167, 249.5921, 249.7016, 
    250.5706,
  271.6901, 269.7879, 266.8765, 262.603, 256.9727, 252.8485, 250.1803, 
    250.2451, 250.6575, 250.8588, 250.0305, 249.2517, 248.7882, 248.9355, 
    249.4997,
  270.0999, 267.0461, 262.9558, 256.6023, 253.065, 250.2594, 248.606, 
    249.9459, 250.1194, 248.7151, 248.7438, 248.5445, 246.8398, 246.9391, 
    248.2144,
  260.3281, 259.5408, 259.6886, 259.9312, 262.1812, 263.0345, 265.2867, 
    262.4818, 259.8904, 255.5782, 255.396, 254.9998, 251.479, 250.4115, 
    249.2194,
  260.4989, 260.3027, 260.4979, 261.69, 262.8518, 262.5755, 265.5222, 
    261.3629, 260.3007, 258.4505, 257.86, 258.3618, 257.4858, 255.1103, 
    254.1725,
  266.3875, 264.3669, 264.6211, 266.633, 267.3455, 264.3078, 261.3824, 
    258.6441, 256.8013, 255.8991, 255.4755, 256.7646, 256.7679, 256.5436, 
    255.1855,
  268.2099, 268.9401, 270.9488, 269.3682, 266.5643, 260.9926, 253.3891, 
    255.4336, 254.6958, 253.9571, 254.3222, 254.5735, 254.7905, 255.4626, 
    256.1434,
  269.2135, 270.9156, 271.7411, 265.8006, 259.7827, 258.2737, 256.4777, 
    249.0809, 249.6364, 253.2545, 254.2544, 254.1882, 253.961, 254.3854, 
    255.4449,
  271.4916, 272.3313, 269.1348, 262.4022, 259.2089, 254.4146, 252.9804, 
    251.7305, 250.8039, 249.0116, 250.3851, 252.0353, 252.2337, 252.8259, 
    253.5545,
  273.0277, 270.7624, 266.6505, 262.8032, 261.252, 254.0256, 251.4303, 
    250.2478, 249.5296, 248.8184, 248.5573, 248.7554, 249.1958, 249.3859, 
    249.7187,
  271.4679, 267.7845, 265.2321, 262.6452, 259.2704, 253.5726, 251.2321, 
    250.4424, 250.3107, 249.9503, 249.3456, 248.921, 248.841, 248.751, 
    249.1258,
  269.1959, 265.3027, 262.2197, 258.5278, 253.7182, 252.3605, 251.4009, 
    251.6971, 251.9569, 251.5273, 249.6653, 248.1611, 248.6197, 249.5672, 
    249.3339,
  266.0288, 261.9116, 258.1742, 253.3392, 252.1135, 251.868, 251.4262, 
    252.3003, 251.9936, 248.6676, 247.8537, 247.763, 248.4038, 249.8613, 
    248.7262,
  262.6249, 261.7228, 260.5368, 259.8324, 259.2, 258.9298, 260.9322, 
    261.8807, 260.2909, 256.0391, 253.8987, 252.0654, 250.1299, 250.5492, 
    249.9795,
  262.8154, 262.0115, 261.064, 260.5679, 258.9928, 258.857, 260.9557, 
    258.9621, 254.7884, 252.9451, 251.0459, 251.1684, 251.0063, 249.2097, 
    249.8017,
  266.2335, 263.4744, 262.2373, 261.9866, 262.2799, 260.072, 259.2162, 
    256.2766, 253.1477, 252.0364, 251.5462, 251.4139, 251.2768, 250.9109, 
    250.4321,
  268.2588, 268.3718, 268.2879, 266.8104, 265.6855, 263.9546, 254.5271, 
    253.095, 252.1576, 251.9121, 252.1783, 251.8858, 251.3874, 250.9871, 
    250.1394,
  268.9058, 269.172, 269.8785, 268.0032, 264.691, 263.2205, 259.2077, 249.23, 
    247.6039, 251.8001, 252.6304, 251.716, 250.8858, 250.5728, 250.5929,
  269.1295, 270.1182, 270.2815, 268.2254, 265.2611, 261.6187, 258.8678, 
    254.3828, 251.5803, 248.6288, 248.5553, 250.2149, 250.44, 250.2744, 
    249.8769,
  270.3699, 271.115, 270.6868, 268.3632, 267.2219, 261.1593, 254.7679, 
    251.2605, 250.4926, 250.0303, 250.8483, 250.6682, 250.3683, 249.4543, 
    249.1046,
  272.096, 271.8517, 270.484, 268.3803, 264.6243, 255.7281, 252.0773, 
    250.9341, 251.6458, 251.5573, 251.1917, 250.1381, 248.8247, 248.1579, 
    248.9167,
  273.7418, 272.0834, 269.2299, 264.6915, 257.6725, 253.9709, 252.1751, 
    252.3708, 253.2051, 252.5952, 249.6829, 247.3779, 247.1247, 248.2204, 
    249.1377,
  273.4352, 270.4937, 265.1088, 257.7252, 253.5901, 252.0739, 250.8921, 
    252.4789, 252.3069, 247.9309, 246.6499, 245.277, 245.8836, 248.8092, 
    249.4203,
  264.1085, 263.5738, 262.6701, 262.1118, 260.7938, 260.2758, 259.9751, 
    259.2936, 258.7941, 258.441, 258.9635, 259.4539, 258.0065, 257.1737, 
    255.3023,
  263.9617, 263.2163, 262.6763, 261.2297, 259.9296, 259.7979, 260.3766, 
    259.4715, 259.0451, 259.2609, 258.2003, 257.4734, 256.4928, 254.9149, 
    253.8071,
  266.214, 263.7169, 262.3736, 261.4766, 260.8496, 257.5872, 260.0909, 
    260.2978, 259.3114, 259.1976, 258.4403, 257.4927, 256.5363, 255.4267, 
    254.5708,
  268.2693, 267.6367, 266.3972, 263.5851, 261.8208, 262.0852, 257.0729, 
    259.9504, 260.1049, 259.5028, 258.7793, 257.9093, 256.709, 255.3308, 
    254.2075,
  269.1701, 269.2122, 269.021, 266.3702, 262.4041, 262.9141, 261.8328, 
    256.9082, 256.7983, 259.5151, 260.0579, 258.686, 256.8308, 255.3342, 
    254.1759,
  269.148, 269.8054, 269.6948, 268.2517, 264.6799, 262.9901, 262.7561, 
    261.534, 261.0642, 257.757, 255.9012, 256.2231, 254.9907, 253.6701, 
    252.5068,
  269.3416, 270.1636, 270.3017, 269.4721, 267.9227, 264.7131, 263.2137, 
    261.3116, 259.0639, 256.0936, 254.7804, 253.717, 253.0131, 251.1212, 
    249.9184,
  269.767, 270.277, 270.5426, 270.1884, 269.7643, 266.3537, 263.4532, 
    260.4557, 257.5641, 254.6996, 253.4687, 252.0609, 250.1258, 248.7911, 
    248.5784,
  271.1053, 270.9477, 270.9874, 270.5102, 268.6809, 265.8565, 262.8274, 
    258.9612, 256.4409, 254.2762, 251.2313, 248.735, 247.2753, 246.8034, 
    247.4709,
  271.7973, 271.7439, 270.3614, 267.9688, 265.644, 261.7882, 258.7163, 
    256.0143, 253.8864, 248.8159, 244.7192, 244.8022, 244.7503, 245.8912, 
    247.6402,
  265.1046, 264.8604, 264.4162, 264.0117, 263.2901, 262.435, 262.1464, 
    262.1738, 261.1385, 259.0708, 258.9162, 258.9685, 257.2688, 257.7341, 
    257.1408,
  265.9649, 265.5359, 265.1521, 264.2269, 262.9292, 262.144, 261.7533, 
    261.3592, 260.7855, 260.1455, 259.6675, 259.5837, 258.6643, 256.6213, 
    256.455,
  268.8769, 266.5381, 265.353, 264.7883, 263.7812, 260.5273, 261.5347, 
    260.9334, 260.7266, 260.0318, 259.5525, 259.1747, 258.5063, 257.9677, 
    257.4176,
  270.0833, 269.4612, 268.6646, 266.027, 264.3955, 263.2902, 258.1062, 
    259.9378, 260.0312, 259.5569, 259.2953, 258.9847, 258.5524, 257.881, 
    257.9089,
  270.0189, 269.5399, 269.1794, 266.0163, 263.4711, 263.5248, 261.6891, 
    256.2408, 255.6679, 258.5058, 259.9617, 259.5621, 258.7004, 258.0508, 
    258.1588,
  270.2755, 269.4785, 268.76, 266.203, 263.3892, 262.6773, 262.007, 260.3219, 
    258.6981, 256.9315, 257.7368, 258.5327, 258.0999, 258.1123, 258.0818,
  270.6106, 270.0366, 269.0805, 266.9989, 264.7021, 262.119, 260.7592, 
    259.2069, 257.7935, 257.2317, 257.0903, 256.6436, 256.8481, 256.3751, 
    256.4209,
  270.9945, 270.2034, 269.3554, 267.9388, 265.9341, 261.6455, 260.3725, 
    258.8466, 257.3682, 256.5326, 256.3009, 256.6177, 255.4746, 253.5842, 
    252.9201,
  270.6425, 269.9269, 268.5897, 266.8995, 263.9715, 261.7462, 260.3886, 
    258.6946, 256.5308, 254.067, 251.1056, 249.9561, 248.9091, 246.9854, 
    245.6797,
  266.6277, 266.2159, 263.7201, 260.8652, 259.3293, 257.51, 256.0814, 
    254.6786, 250.7836, 246.3189, 244.0554, 243.5666, 243.2949, 243.3884, 
    244.3948,
  267.6084, 266.9691, 267.0802, 266.5146, 265.2692, 264.5278, 264.4726, 
    264.6157, 264.5674, 262.9704, 261.9318, 262.0778, 260.7721, 260.0188, 
    259.5779,
  268.1689, 267.8887, 267.3336, 265.5326, 264.4478, 264.2155, 263.9936, 
    263.1516, 264.161, 263.8214, 262.8121, 262.6868, 262.0426, 259.2707, 
    258.0844,
  269.9838, 267.7683, 266.2504, 264.8803, 264.0294, 261.9178, 263.8343, 
    263.3454, 262.9077, 263.0024, 262.2186, 261.1738, 260.6226, 259.8131, 
    258.8387,
  269.9655, 268.9881, 267.6909, 264.677, 263.6775, 263.7333, 260.0292, 
    262.308, 261.4745, 260.9992, 260.2271, 260.0827, 259.7382, 259.8754, 
    258.9428,
  269.6132, 268.0133, 266.4898, 263.2527, 261.643, 262.5104, 262.5693, 
    256.6548, 257.2494, 259.8187, 260.2515, 259.8094, 259.2671, 258.9062, 
    258.7431,
  269.1329, 267.6628, 265.6617, 262.6676, 260.161, 259.2502, 260.2372, 
    260.2323, 259.5991, 259.4481, 259.4113, 259.6772, 259.188, 258.8231, 
    258.0808,
  268.3224, 267.1514, 265.3082, 262.4985, 259.8568, 256.5278, 256.4676, 
    257.086, 257.4504, 257.5536, 257.5506, 257.5372, 257.513, 257.218, 
    257.2763,
  267.3767, 266.1293, 264.2794, 262.1219, 259.2847, 254.8765, 254.152, 
    253.108, 252.9946, 252.712, 252.7716, 252.9638, 252.8158, 252.8748, 
    252.8205,
  266.4623, 264.6675, 262.2316, 258.5581, 254.0855, 253.054, 252.256, 
    251.2257, 249.2988, 247.8211, 246.6934, 247.2613, 247.3966, 247.2712, 
    246.3893,
  265.5391, 263.5019, 259.7071, 253.1944, 250.407, 249.8396, 250.9111, 
    251.9799, 248.2584, 245.085, 244.2222, 244.9364, 244.8931, 245.1689, 
    244.6903,
  264.1958, 263.1046, 263.4445, 262.6286, 260.2791, 259.396, 260.0201, 
    259.6591, 259.9722, 260.3364, 261.2834, 262.3866, 262.4122, 262.2635, 
    261.887,
  264.6204, 263.9976, 263.3359, 261.9946, 258.7855, 258.2239, 258.1224, 
    257.7527, 258.0529, 259.2126, 260.6906, 262.1419, 262.4745, 261.0883, 
    261.014,
  269.301, 266.102, 263.5819, 261.8464, 258.5533, 254.2997, 256.499, 
    256.5806, 257.3595, 258.652, 260.008, 260.4943, 260.5522, 260.9159, 
    260.5374,
  269.9899, 269.7261, 268.8541, 264.5125, 259.6897, 257.0087, 251.1074, 
    254.4034, 256.5051, 256.5436, 257.4827, 257.8953, 258.3174, 258.8405, 
    259.3431,
  270.4806, 269.9145, 269.2462, 265.0862, 259.7204, 257.1327, 256.2709, 
    246.9302, 249.931, 254.9465, 255.7403, 255.5611, 255.2887, 255.9613, 
    257.2476,
  271.1942, 270.5658, 269.3448, 265.4435, 259.3155, 255.3692, 254.4185, 
    252.9027, 252.4925, 252.5248, 251.9861, 253.0275, 253.3633, 254.2322, 
    255.1908,
  272.1313, 271.4685, 270.155, 265.9767, 259.381, 253.9861, 251.9374, 
    251.2931, 251.1075, 250.8587, 250.4615, 250.4796, 250.4194, 251.2531, 
    252.5242,
  272.7291, 272.1985, 270.1911, 265.5681, 258.7775, 252.545, 250.6832, 
    249.6845, 249.6263, 249.171, 248.6253, 249.1108, 248.045, 248.9651, 
    249.6156,
  272.2684, 271.2553, 268.9575, 263.2637, 255.1375, 251.7919, 250.7441, 
    250.7559, 249.6911, 248.434, 247.3539, 247.5147, 246.2905, 246.8292, 
    247.4393,
  270.6628, 269.1169, 265.7976, 258.088, 252.036, 250.5446, 250.7592, 
    251.5551, 249.2767, 246.7137, 245.9213, 246.1526, 244.9577, 245.4347, 
    245.5467,
  264.9844, 264.7872, 263.9718, 263.64, 262.4155, 262.3021, 263.3235, 
    261.3903, 259.797, 258.1283, 257.1756, 256.7762, 255.2154, 254.4133, 
    253.9581,
  262.8412, 263.0224, 263.3128, 262.8514, 261.9482, 262.0456, 261.5129, 
    260.1826, 259.0592, 257.5546, 256.8123, 257.2094, 255.7804, 253.196, 
    252.2772,
  267.7502, 264.8342, 262.8003, 262.4504, 261.163, 258.4918, 259.771, 
    259.1171, 257.4763, 257.7599, 257.8641, 257.0261, 255.8425, 254.2182, 
    252.6064,
  269.5055, 269.2475, 268.1754, 265.1679, 262.0551, 261.5016, 258.0817, 
    259.2177, 259.339, 257.7179, 256.4639, 254.9742, 254.1167, 253.1923, 
    251.5648,
  270.6508, 270.1759, 270.0399, 267.7603, 264.7855, 265.1495, 264.0784, 
    254.0997, 248.6205, 252.4397, 253.1896, 252.0437, 251.6737, 251.0839, 
    250.9707,
  271.6216, 270.2903, 268.316, 264.5144, 261.6046, 259.3094, 256.5829, 
    253.9296, 250.6626, 247.7231, 247.5244, 248.8681, 249.2998, 249.2625, 
    249.3883,
  269.5322, 267.5002, 264.8334, 260.2942, 256.7159, 253.2562, 251.9242, 
    249.8514, 248.0431, 247.636, 247.6457, 247.6392, 247.1417, 246.7631, 
    247.5185,
  268.163, 266.3192, 263.9169, 260.9388, 256.3725, 251.3255, 249.5175, 
    247.9163, 247.925, 247.5475, 246.3601, 246.1669, 244.8203, 245.1912, 
    246.4559,
  266.1207, 263.9581, 261.4662, 257.3589, 251.6328, 250.0107, 248.932, 
    248.636, 247.8692, 246.5075, 244.9929, 244.5103, 244.0275, 244.0306, 
    244.9491,
  263.6008, 261.0988, 256.8161, 250.9928, 249.2706, 248.6353, 248.3589, 
    249.3864, 247.7125, 245.4648, 244.413, 244.3039, 243.7369, 243.5134, 
    243.9035,
  266.0075, 265.3306, 264.4623, 264.3803, 265.712, 266.8681, 267.4736, 
    266.5365, 265.682, 265.1336, 264.8736, 264.703, 263.0586, 262.0876, 
    260.5386,
  265.4763, 264.7403, 264.2026, 263.9333, 263.6346, 263.7073, 264.437, 
    264.6353, 264.5316, 264.2456, 263.5653, 263.9528, 262.7668, 260.76, 
    259.6496,
  267.7509, 265.3011, 263.9514, 263.1729, 262.3932, 259.3918, 261.148, 
    261.4924, 262.0174, 263.2634, 263.4402, 262.8502, 262.1977, 261.7681, 
    260.5032,
  269.5247, 268.4467, 266.6231, 263.8161, 261.85, 261.6531, 259.0131, 
    260.0586, 260.1632, 259.923, 259.2787, 257.6853, 257.2791, 256.1469, 
    254.6422,
  269.774, 268.3408, 266.8737, 263.5049, 261.2617, 262.7821, 262.9268, 
    254.8303, 251.5083, 253.4676, 254.6541, 253.0245, 252.3462, 251.6921, 
    251.1826,
  267.6081, 265.6613, 262.8487, 258.4825, 256.8606, 256.093, 257.5678, 
    256.8958, 251.9301, 249.1657, 248.6241, 249.859, 249.4464, 249.0731, 
    248.3001,
  266.1237, 264.2092, 261.3466, 257.0979, 255.4071, 252.5726, 251.7996, 
    250.5934, 248.6009, 248.7417, 247.9728, 247.6194, 247.9996, 248.1326, 
    248.0551,
  267.4625, 265.5632, 263.5537, 261.4732, 257.2495, 251.065, 249.3134, 
    248.8433, 248.7811, 248.5964, 248.0193, 247.9883, 247.9647, 248.3094, 
    248.5229,
  268.0556, 266.7227, 265.2194, 263.173, 257.6427, 254.3595, 252.4907, 
    251.46, 250.8043, 250.5846, 250.3911, 250.0296, 249.7673, 249.5971, 
    249.2472,
  268.6853, 267.5596, 265.6898, 260.5868, 256.876, 255.2342, 253.2914, 
    253.2023, 253.3824, 253.1331, 253.4877, 252.7523, 251.9693, 251.8888, 
    251.3982,
  265.5267, 263.776, 263.3145, 263.7281, 267.1402, 268.5977, 269.4564, 
    268.5429, 269.2503, 268.3645, 268.1696, 268.6203, 267.7012, 266.5938, 
    266.4669,
  265.1514, 263.6686, 263.3424, 263.0969, 264.2009, 267.3761, 268.4844, 
    268.681, 269.1372, 268.8069, 268.3651, 268.4609, 267.3549, 265.1414, 
    265.0737,
  268.0522, 265.5853, 264.2036, 262.8294, 262.9707, 262.2265, 266.6717, 
    268.4567, 269.1057, 269.0307, 268.6347, 267.9517, 267.0207, 266.3625, 
    264.8222,
  268.6241, 267.6446, 266.1718, 262.0248, 261.9128, 263.5945, 262.8791, 
    265.7527, 267.3097, 267.8969, 267.9877, 267.157, 266.4459, 265.4339, 
    263.8492,
  268.6435, 267.3321, 266.0915, 261.0202, 260.1258, 261.6796, 263.9033, 
    260.3007, 259.3991, 265.0489, 266.2872, 265.4507, 264.9574, 264.2169, 
    262.8404,
  269.2795, 268.0987, 265.9766, 260.1359, 259.1363, 258.7858, 260.0608, 
    261.6033, 261.4027, 262.464, 263.1255, 263.047, 262.8111, 262.155, 
    260.5717,
  270.3647, 269.2632, 267.1534, 261.7816, 259.0929, 257.3275, 257.2538, 
    258.1627, 259.6406, 260.2861, 260.0762, 260.2022, 260.0416, 259.3656, 
    257.5966,
  271.7182, 271.3309, 270.1776, 267.838, 261.9518, 254.8701, 254.529, 
    254.7261, 255.4055, 256.9085, 257.507, 257.5045, 257.2087, 256.7368, 
    255.3604,
  272.7611, 272.5496, 271.9791, 270.2357, 264.9449, 257.335, 254.1931, 
    253.612, 253.6852, 254.2112, 254.8222, 255.056, 254.6705, 253.6786, 
    252.5154,
  272.2025, 271.742, 270.941, 268.9918, 266.8951, 260.3119, 254.8778, 
    252.9948, 252.6044, 252.1444, 253.9964, 253.3518, 252.9783, 252.9288, 
    252.3602,
  262.6177, 261.2606, 260.3084, 262.9781, 265.2805, 265.9273, 265.0523, 
    262.7865, 261.8495, 265.0705, 263.2204, 266.3047, 266.3536, 265.6611, 
    264.9645,
  263.9233, 262.9466, 262.629, 265.0127, 265.1281, 265.3366, 264.9592, 
    261.6591, 265.0707, 264.6544, 264.7993, 267.8855, 267.5646, 266.7458, 
    264.4258,
  270.008, 267.1339, 265.7697, 266.0448, 264.5065, 264.3981, 266.3134, 
    263.5618, 268.0069, 268.3698, 268.6886, 268.5079, 268.7559, 268.0069, 
    265.9281,
  270.8665, 270.6036, 270.5647, 267.2768, 264.5938, 265.7611, 264.3277, 
    265.2794, 268.5265, 268.6659, 268.5243, 267.7511, 267.6085, 266.366, 
    264.3384,
  271.4413, 271.1055, 270.9559, 265.8439, 263.993, 265.0854, 268.8517, 
    265.7887, 265.2649, 267.925, 268.1862, 266.7112, 266.4882, 264.6486, 
    263.8375,
  271.2425, 271.1089, 270.8, 266.036, 264.5854, 263.7158, 265.4845, 268.0544, 
    267.7275, 267.3738, 267.1658, 266.9398, 265.2734, 262.7923, 262.0848,
  270.5735, 270.5253, 270.6988, 268.7284, 265.9052, 262.9141, 264.6172, 
    266.0989, 267.1438, 267.4012, 266.6918, 266.5474, 264.3624, 262.4572, 
    260.569,
  269.4985, 269.4758, 269.8778, 270.7961, 267.7139, 261.2189, 261.52, 
    263.0694, 265.5092, 266.5239, 266.197, 266.1294, 263.9115, 261.6851, 
    259.0135,
  266.9987, 266.7855, 267.872, 269.7226, 269.2129, 264.258, 259.954, 
    262.1835, 263.2341, 264.6897, 266.0327, 265.7726, 263.3723, 260.4755, 
    258.0671,
  263.6013, 261.9778, 262.0442, 263.888, 268.1417, 265.251, 260.2065, 
    259.253, 261.1163, 262.7967, 264.795, 265.1758, 262.738, 259.8478, 
    258.7404,
  264.7237, 263.2468, 261.4502, 261.2719, 262.2553, 260.5101, 262.0896, 
    262.0519, 261.8418, 263.4354, 260.1734, 262.4189, 262.9143, 262.7676, 
    261.7337,
  266.4204, 265.0841, 263.901, 262.5008, 262.6677, 259.903, 260.9744, 
    261.1317, 262.7774, 259.029, 260.1601, 262.8534, 264.0066, 263.1476, 
    259.63,
  268.9849, 267.4018, 264.7761, 263.1648, 262.5419, 259.8814, 259.0965, 
    258.3568, 261.7921, 261.7571, 265.0577, 265.0083, 264.9883, 264.3824, 
    262.9162,
  268.506, 268.0995, 268.0135, 265.3619, 263.7762, 263.338, 260.2136, 
    260.0319, 265.2289, 265.6984, 262.9108, 264.2116, 265.1957, 265.7027, 
    265.1874,
  267.9683, 266.7575, 266.8395, 264.2223, 263.7031, 264.5502, 265.0541, 
    262.2757, 259.1964, 261.738, 264.5153, 265.7772, 266.3394, 266.6606, 
    266.0216,
  267.1299, 265.8044, 265.2554, 263.8622, 264.1501, 264.793, 265.1328, 
    264.7779, 263.9975, 264.8099, 263.1004, 265.8359, 266.5446, 266.1595, 
    263.6324,
  266.2793, 264.7461, 263.9437, 263.5611, 265.1896, 263.715, 266.1899, 
    261.597, 264.5575, 266.2352, 264.8317, 265.2428, 265.554, 263.578, 
    257.7875,
  265.2167, 263.4885, 262.5342, 262.8901, 265.551, 262.551, 261.3092, 
    263.3333, 264.263, 265.7123, 264.3077, 264.4929, 262.5527, 256.8329, 252.6,
  264.0918, 261.8886, 260.6028, 259.837, 264.5773, 264.8437, 261.7408, 
    262.786, 264.8506, 264.4569, 263.5524, 262.5278, 257.1712, 253.4907, 
    252.303,
  262.5131, 259.5269, 256.7862, 255.6919, 262.7204, 265.2732, 263.1993, 
    264.6916, 263.4396, 263.2282, 262.2086, 258.7674, 254.9019, 253.572, 
    253.1626,
  263.9331, 261.4456, 259.0991, 259.3966, 261.7411, 262.1843, 261.1423, 
    262.3753, 263.4173, 262.3512, 262.5096, 264.2699, 262.9178, 261.8381, 
    260.7384,
  265.5171, 262.4402, 260.6862, 260.1738, 261.3434, 261.3951, 262.1709, 
    262.206, 262.5945, 262.4983, 262.1232, 264.009, 263.4531, 259.8416, 
    258.3558,
  268.9861, 266.7584, 263.241, 260.9685, 260.0243, 260.3467, 260.8216, 
    260.1275, 258.8741, 260.048, 263.6034, 263.7798, 262.5776, 260.8036, 
    257.3455,
  269.1478, 268.601, 267.6523, 263.0482, 261.3376, 262.09, 260.222, 259.4887, 
    261.8671, 262.0482, 261.8191, 262.5134, 261.4167, 259.3107, 257.2043,
  268.9354, 268.269, 267.7112, 263.8644, 262.5573, 263.0081, 263.9779, 
    255.8109, 257.1703, 259.7351, 262.0226, 261.8784, 260.3486, 258.927, 
    257.089,
  268.3816, 268.1316, 267.5028, 265.6772, 264.6732, 263.4468, 264.0465, 
    263.7243, 261.2413, 261.9187, 260.5346, 261.1738, 259.0582, 257.3183, 
    255.3375,
  267.745, 267.2742, 267.2676, 266.7504, 265.765, 262.4339, 262.8179, 
    261.8285, 261.8032, 261.4952, 261.217, 259.4928, 256.7112, 253.9352, 
    252.2884,
  266.6113, 266.0708, 265.5343, 266.2048, 266.3891, 262.3924, 261.1248, 
    261.3578, 260.0715, 260.8604, 258.6296, 255.6302, 252.8093, 251.1698, 
    250.4847,
  265.0979, 264.0369, 263.2896, 261.7607, 263.1719, 263.0628, 260.4483, 
    260.622, 261.1738, 258.0977, 255.062, 252.6957, 251.1047, 250.8361, 
    250.5041,
  262.8036, 260.8516, 258.7797, 257.6986, 259.8112, 261.1179, 260.9357, 
    260.218, 259.5107, 255.8545, 252.7666, 251.1929, 250.8427, 250.8839, 
    251.1946,
  265.632, 262.7832, 261.0593, 262.291, 261.6665, 259.5823, 258.413, 
    259.9371, 260.3781, 259.4419, 259.1018, 260.3468, 259.5135, 258.362, 
    256.5512,
  267.3834, 263.9588, 263.1318, 262.3623, 260.8278, 257.926, 257.9044, 
    258.7045, 258.0074, 258.79, 258.2603, 260.0054, 260.1956, 256.9055, 
    256.3003,
  270.7654, 268.1355, 264.9392, 263.4101, 260.1199, 257.4345, 256.5615, 
    257.7103, 256.9238, 257.3454, 257.5605, 258.3427, 259.2176, 259.2729, 
    257.3394,
  271.0147, 269.9922, 268.1531, 263.7061, 261.543, 260.1498, 253.0791, 
    256.1591, 256.5692, 255.7993, 255.5309, 255.9753, 257.1119, 257.801, 
    258.0825,
  271.119, 269.9269, 268.2572, 262.8908, 261.0492, 260.6223, 259.1322, 
    251.6443, 252.1399, 254.6835, 254.6408, 254.1711, 254.9308, 255.5988, 
    256.6588,
  270.9141, 270.0347, 268.5847, 265.5617, 262.3151, 259.215, 258.3237, 
    257.6792, 254.5892, 255.029, 253.0563, 253.3069, 252.8692, 253.3062, 
    254.3204,
  270.4269, 269.222, 268.7777, 266.9156, 263.1198, 257.6895, 255.2387, 
    254.3287, 254.1041, 253.0487, 252.2499, 251.9758, 251.8446, 251.5366, 
    251.7754,
  270.2707, 268.9196, 267.0525, 266.9709, 265.4691, 258.6772, 254.5277, 
    252.7034, 251.4821, 251.0724, 250.3289, 250.5472, 250.5304, 250.7339, 
    250.5522,
  270.3608, 268.1175, 266.1805, 263.097, 263.4367, 262.0085, 255.1754, 
    252.8953, 250.7859, 249.4599, 249.0855, 249.4486, 249.2861, 249.9804, 
    250.5059,
  269.8008, 266.7819, 263.4643, 260.924, 260.8188, 260.314, 256.4965, 
    253.8922, 251.0769, 248.7731, 248.2712, 248.618, 248.2692, 249.0133, 
    250.3307,
  270.2751, 267.0952, 263.9043, 263.6691, 261.9125, 258.89, 257.1234, 
    256.2069, 255.8203, 255.3774, 255.5126, 257.672, 256.5197, 256.1386, 
    256.2067,
  270.5625, 268.9679, 265.9357, 264.3357, 263.1422, 260.0736, 258.3239, 
    256.8735, 256.1682, 256.433, 255.3858, 256.9509, 258.1102, 254.0054, 
    253.0205,
  272.1656, 271.0315, 268.3707, 265.8899, 262.8856, 258.6192, 258.8686, 
    257.0704, 256.4241, 255.8049, 255.5031, 256.1049, 257.2199, 257.3223, 
    254.1247,
  273.1179, 272.3477, 271.432, 267.3773, 264.2101, 261.5648, 256.5036, 
    256.8734, 256.5609, 255.6812, 254.94, 254.748, 255.5889, 256.2942, 
    255.8423,
  274.0513, 272.5921, 271.6447, 267.5652, 264.6485, 261.868, 259.9669, 
    252.8175, 251.895, 255.4166, 254.7483, 254.3068, 254.3656, 254.8943, 
    256.1702,
  274.2101, 272.7568, 271.0748, 267.9724, 265.3411, 261.9162, 259.5563, 
    259.226, 257.8851, 257.1151, 254.8296, 254.3287, 253.3964, 253.3322, 
    254.0159,
  274.1315, 272.84, 270.8599, 268.1208, 264.7967, 261.0617, 259.0971, 
    258.4222, 257.8464, 257.1292, 255.3255, 254.3896, 253.1244, 252.3065, 
    252.9198,
  273.5959, 272.1683, 269.8788, 266.9757, 263.7416, 260.4283, 258.8972, 
    258.8392, 258.1688, 257.2756, 256.3537, 254.7442, 252.7336, 251.5351, 
    251.4053,
  272.7427, 270.9045, 268.4538, 264.2149, 260.8527, 258.9106, 258.7055, 
    259.4952, 259.0355, 257.872, 256.6443, 255.1532, 252.843, 251.4293, 
    251.4202,
  271.2036, 268.6068, 265.1889, 261.5439, 258.7245, 257.3025, 258.0005, 
    259.8553, 260.0595, 258.0503, 256.7076, 254.8966, 252.5176, 251.4189, 
    251.3699,
  268.897, 267.7884, 265.4228, 263.7451, 262.6023, 261.4581, 260.9679, 
    259.9966, 259.2521, 257.6965, 257.549, 256.9197, 255.8191, 256.1967, 
    256.4607,
  269.0177, 267.7307, 265.2599, 262.7904, 261.456, 259.9886, 259.7523, 
    258.9976, 258.0599, 258.0553, 255.9466, 256.1498, 256.8393, 255.2383, 
    255.2753,
  270.5753, 269.0379, 266.2772, 262.4005, 260.1731, 257.363, 258.8354, 
    258.8058, 257.8947, 256.726, 256.2032, 256.5167, 256.9584, 257.8095, 
    257.3043,
  270.7048, 269.4504, 267.2438, 262.5098, 260.0602, 258.7295, 255.8349, 
    258.2823, 258.7442, 257.5012, 256.288, 257.6659, 257.3692, 258.655, 
    258.3414,
  270.5235, 268.7986, 266.4974, 261.5986, 260.052, 259.0318, 258.5955, 
    254.6436, 255.0067, 258.4428, 256.7301, 257.5071, 258.78, 258.7639, 
    258.7039,
  270.3265, 268.5209, 265.8172, 261.7228, 260.0067, 258.9923, 259.0655, 
    259.4846, 259.4285, 258.9066, 256.6594, 257.5325, 258.2584, 258.2672, 
    258.1667,
  270.1394, 268.1075, 265.7434, 262.8616, 259.6195, 257.696, 258.7007, 
    259.1302, 259.1168, 258.3225, 256.9548, 256.951, 257.0081, 256.6178, 
    256.1985,
  270.2605, 267.6928, 264.735, 262.0737, 259.58, 256.8834, 257.6047, 
    258.2669, 258.2642, 257.9835, 255.9448, 256.4783, 255.5662, 254.7377, 
    254.4561,
  270.5181, 267.1648, 264.0632, 259.3814, 257.2833, 256.1573, 256.9539, 
    257.601, 257.3025, 256.6281, 256.0573, 255.1397, 253.9348, 252.5665, 
    251.4081,
  269.9893, 265.8798, 261.4148, 257.9914, 256.8724, 255.698, 255.6217, 
    257.3235, 256.4894, 254.5397, 253.4185, 253.302, 252.102, 251.8595, 
    251.0217,
  266.8927, 265.3689, 262.6664, 261.2045, 260.9934, 259.0168, 258.3152, 
    257.9032, 257.3198, 256.1677, 257.5917, 257.0854, 254.4656, 253.7202, 
    253.8648,
  268.1292, 267.0724, 264.9631, 262.547, 261.6523, 259.6888, 259.7281, 
    258.8813, 258.0451, 257.2556, 255.2649, 257.9216, 257.7066, 255.7593, 
    251.6472,
  271.8011, 270.3274, 268.532, 265.0909, 262.0835, 258.761, 260.4168, 
    259.9127, 258.9431, 257.2355, 256.7721, 257.3619, 258.4526, 259.328, 
    255.3031,
  272.5768, 271.5881, 270.8204, 267.3152, 264.4105, 261.3971, 257.9792, 
    259.5579, 259.6416, 257.6414, 256.3398, 257.5054, 258.158, 257.9107, 
    257.2704,
  273.6472, 272.2362, 271.4803, 268.066, 266.3074, 263.9038, 260.6263, 
    255.3906, 255.1525, 258.3417, 256.287, 255.544, 256.3315, 257.3969, 
    258.0058,
  274.5097, 273.2814, 271.8492, 269.6006, 268.2616, 266.0313, 263.0166, 
    260.5912, 259.0133, 257.6, 255.3816, 254.7464, 254.3097, 254.8314, 
    255.9337,
  275.1927, 274.3097, 272.9424, 271.1606, 269.3384, 266.8146, 264.7163, 
    262.4503, 260.0918, 258.0433, 255.9113, 254.6969, 253.6308, 253.0329, 
    253.1455,
  275.5867, 274.895, 273.5887, 271.9485, 270.5927, 268.2332, 265.8051, 
    263.9941, 261.7319, 259.2404, 256.0796, 254.1788, 253.1087, 252.0378, 
    251.6296,
  275.374, 274.6199, 273.7314, 272.3315, 270.9368, 269.1617, 267.1279, 
    265.4166, 263.3877, 260.5364, 256.979, 254.2665, 252.4522, 251.4116, 
    250.9532,
  274.401, 273.4496, 272.6792, 272.1372, 271.1137, 269.726, 267.8839, 
    266.4628, 264.7591, 260.9219, 256.8103, 254.1626, 251.8132, 250.371, 
    251.1241,
  271.9366, 271.4437, 271.2425, 271.2599, 271.1078, 270.4268, 269.4467, 
    267.6982, 265.0865, 261.1568, 260.9335, 260.0952, 257.6732, 256.21, 
    254.6668,
  272.0014, 272.1754, 272.0706, 272.1181, 272.0601, 271.5038, 270.8323, 
    269.6709, 267.8587, 264.4091, 261.8475, 260.9583, 259.9809, 257.8003, 
    255.3999,
  272.9972, 272.3616, 272.0863, 272.2744, 272.4916, 270.9429, 271.7657, 
    271.2513, 269.6337, 267.6376, 264.735, 262.6214, 261.0547, 260.4157, 
    259.0742,
  273.5392, 272.7737, 272.283, 271.8214, 272.1873, 272.1005, 270.5296, 
    271.1373, 270.1205, 268.6988, 266.2121, 263.9149, 261.924, 260.6298, 
    259.5613,
  273.9524, 272.6522, 272.0712, 271.336, 271.5038, 271.5632, 271.339, 
    268.4868, 267.709, 270.3546, 269.169, 266.3518, 263.3831, 261.0782, 
    259.925,
  274.1603, 272.8455, 271.4586, 270.5963, 270.5518, 270.1727, 270.345, 
    270.047, 269.8742, 269.7379, 268.8098, 267.1437, 264.4343, 261.7231, 
    259.7749,
  274.0591, 272.9187, 271.407, 270.0484, 269.3188, 268.7712, 268.6205, 
    269.0708, 269.025, 269.1457, 268.3507, 266.7942, 263.7227, 260.873, 
    259.0712,
  273.7082, 272.5578, 270.8318, 268.9125, 267.8609, 267.373, 267.1177, 
    267.2604, 267.0164, 267.5185, 267.2807, 265.2162, 261.598, 259.0446, 
    257.8589,
  273.2844, 272.0259, 270.2368, 267.0546, 265.5563, 265.4641, 265.1936, 
    265.3315, 265.2797, 265.0563, 264.1775, 261.4699, 258.5492, 256.9291, 
    255.138,
  272.5977, 270.8949, 268.5391, 265.8902, 263.8737, 263.2638, 262.5757, 
    262.9442, 262.4513, 260.9878, 259.7608, 257.0771, 255.4645, 253.8749, 
    252.1203,
  272.6504, 271.7019, 270.9897, 269.7914, 268.0875, 266.8911, 266.3749, 
    266.1006, 268.6345, 268.453, 268.3967, 267.5565, 263.7055, 260.7423, 
    258.4379,
  272.6471, 272.0297, 271.2195, 269.6383, 267.0904, 265.0723, 264.6809, 
    264.0979, 264.8619, 266.3219, 266.9178, 267.5594, 265.7622, 261.514, 
    259.321,
  273.1517, 272.3561, 271.6154, 269.7972, 267.0786, 262.2551, 264.0671, 
    262.7055, 263.2195, 265.3781, 266.3755, 267.3325, 267.4156, 265.3322, 
    261.9284,
  274.0484, 273.3091, 272.4261, 270.036, 267.1527, 263.74, 259.1208, 
    261.7094, 261.549, 262.7001, 264.4883, 266.3866, 267.6505, 267.2307, 
    263.8671,
  274.8159, 273.6254, 272.8125, 270.0847, 267.4975, 263.9659, 261.3536, 
    255.7422, 257.0427, 260.9876, 263.0042, 265.3586, 267.205, 268.3046, 
    266.7631,
  275.3942, 274.3489, 272.7529, 270.5913, 268.6677, 265.1313, 261.6712, 
    260.3595, 258.0799, 258.8742, 260.9126, 264.0574, 266.249, 267.5503, 
    266.3207,
  275.7245, 274.9345, 273.4304, 271.5606, 269.4445, 266.3167, 262.853, 
    260.6981, 258.5756, 257.6669, 258.9764, 261.5045, 264.1349, 264.4638, 
    262.8464,
  275.9453, 275.1143, 273.7718, 272.0464, 270.1827, 267.3176, 264.1318, 
    261.1785, 258.1187, 256.2033, 257.3341, 256.972, 258.274, 258.8508, 
    258.3304,
  275.7357, 274.968, 273.8752, 272.1553, 270.0753, 267.6112, 264.6303, 
    261.9535, 258.9493, 256.286, 255.3479, 256.4237, 255.0029, 254.4992, 
    253.9353,
  274.7782, 273.9386, 273.0607, 271.934, 270.2349, 268.1858, 265.4933, 
    263.1667, 260.4736, 256.5764, 254.0598, 253.5872, 253.0436, 252.5332, 
    252.4276,
  273.5756, 273.0089, 272.6404, 272.6727, 272.2521, 269.4024, 267.7469, 
    264.673, 263.0334, 263.2177, 259.9388, 263.6459, 265.2689, 264.7664, 
    263.5536,
  273.3038, 272.8307, 272.4157, 272.2672, 272.2662, 270.0145, 268.1014, 
    264.852, 261.6737, 261.4069, 261.9336, 263.8882, 264.9697, 264.0139, 
    262.5377,
  273.653, 272.7792, 272.2199, 271.9357, 272.2295, 269.5679, 268.3518, 
    265.7971, 262.6765, 261.7978, 261.7735, 263.0921, 263.5045, 265.4704, 
    264.7947,
  274.576, 273.6155, 272.6592, 271.6602, 271.8372, 271.6924, 267.6852, 
    265.4418, 263.4622, 262.1776, 261.938, 261.2586, 262.2047, 264.3932, 
    265.7006,
  275.2405, 273.7649, 272.5321, 271.3548, 271.2834, 271.5467, 270.3519, 
    264.119, 261.5969, 264.9308, 263.1375, 261.552, 262.3596, 264.0356, 
    265.9848,
  275.7105, 274.1588, 272.122, 270.9344, 270.6493, 270.6961, 270.594, 
    269.1662, 266.9817, 264.173, 262.1605, 261.6241, 261.1057, 262.2996, 
    265.169,
  275.9142, 274.4727, 272.3835, 270.5007, 269.5919, 269.4797, 269.8715, 
    269.5436, 267.8425, 265.1534, 262.5946, 260.9104, 260.2719, 261.3333, 
    262.5834,
  275.8652, 274.3518, 272.2032, 269.6729, 268.0524, 267.637, 268.324, 
    268.6378, 267.755, 265.2553, 262.9476, 261.0646, 259.5714, 258.8164, 
    260.6634,
  275.5307, 273.8499, 271.6719, 268.0518, 265.9619, 265.6509, 266.2473, 
    266.6027, 266.2235, 264.591, 262.5021, 261.1488, 259.9703, 258.0945, 
    257.166,
  274.4767, 272.6379, 270.4479, 267.2427, 264.3957, 263.5989, 263.8311, 
    264.0704, 264.0862, 262.7982, 261.3522, 260.7676, 259.6934, 258.6194, 
    256.8831,
  273.5339, 272.4854, 271.4479, 269.8626, 268.4744, 268.6503, 268.827, 
    270.2994, 269.1062, 266.5273, 262.9303, 263.062, 261.1238, 263.6007, 
    265.4029,
  273.217, 272.4416, 270.9786, 268.9896, 266.5891, 266.1877, 267.6111, 
    269.0442, 269.08, 267.3432, 265.0477, 264.098, 262.6262, 260.854, 264.0326,
  273.5571, 272.4202, 270.9554, 268.2586, 266.14, 264.0927, 266.7234, 
    267.8465, 267.8651, 266.9218, 265.8144, 265.3167, 263.7204, 262.0952, 
    262.7521,
  274.1103, 272.75, 271.1338, 267.5421, 265.0051, 264.0101, 263.511, 265.435, 
    266.0274, 265.5197, 265.0577, 265.4661, 264.9159, 263.0726, 263.1973,
  274.3605, 272.2558, 270.5836, 266.8056, 263.886, 262.4054, 263.1059, 
    260.8998, 260.7584, 264.0165, 264.5323, 264.7766, 265.3956, 264.481, 
    263.3153,
  274.2457, 272.0694, 269.6607, 266.352, 263.0774, 260.3524, 260.9821, 
    260.8557, 260.9592, 261.3378, 261.1945, 262.2092, 263.3884, 264.368, 
    263.8764,
  273.7577, 271.7142, 269.1406, 265.9305, 261.82, 259.1618, 258.5693, 
    258.5487, 258.0361, 257.8132, 257.7466, 259.0458, 260.576, 261.9699, 
    263.4478,
  273.1357, 270.8911, 267.7609, 263.888, 260.2324, 257.7248, 256.9778, 
    256.2452, 255.6303, 255.1676, 254.9048, 255.8209, 257.7385, 259.8965, 
    262.0148,
  272.1047, 269.8445, 265.9542, 260.94, 257.6919, 256.8939, 256.0404, 
    255.6147, 254.3199, 253.9014, 253.046, 253.282, 254.4648, 257.417, 259.879,
  270.5673, 267.9622, 263.7626, 259.7704, 257.2922, 255.4404, 254.4208, 
    254.5607, 253.4971, 251.9581, 251.2889, 251.6913, 252.1681, 254.6428, 
    257.5073,
  266.1454, 261.9085, 259.4978, 258.972, 258.3875, 257.7444, 256.657, 
    257.273, 258.0886, 258.2909, 259.61, 262.4074, 263.4871, 263.1826, 
    262.0689,
  267.7915, 263.9268, 260.0213, 258.2931, 257.4963, 255.6059, 255.4443, 
    255.472, 255.7336, 255.757, 256.7686, 260.0968, 261.7647, 261.2556, 
    261.4392,
  269.1738, 267.2341, 264.2408, 258.864, 257.0254, 253.1942, 255.1342, 
    254.2781, 253.7682, 253.6259, 254.0654, 256.6277, 259.4729, 261.3931, 
    263.0446,
  269.3004, 267.6255, 265.4679, 259.6577, 257.5475, 255.3243, 251.2837, 
    253.5663, 253.8844, 252.8683, 252.5486, 253.7845, 256.592, 259.4481, 
    262.2334,
  269.577, 267.8334, 265.8902, 261.1189, 259.3131, 255.7811, 254.0642, 
    248.0499, 248.5345, 252.8452, 252.1364, 251.894, 253.4003, 256.5286, 
    260.6568,
  269.7973, 268.059, 266.0828, 262.9518, 260.9647, 256.2649, 254.3583, 
    253.1388, 251.4977, 249.9698, 249.3381, 250.3279, 251.6376, 253.4405, 
    257.6266,
  269.8225, 268.1896, 266.323, 263.8711, 260.606, 256.6864, 254.7416, 
    253.6072, 252.5589, 250.9524, 249.6144, 249.3782, 250.489, 251.5427, 
    254.7481,
  269.627, 267.9686, 266.0132, 262.7968, 260.1013, 257.085, 255.3113, 
    254.0417, 252.8962, 251.6127, 249.9426, 248.9571, 249.0504, 250.1868, 
    253.6171,
  269.2735, 267.5792, 265.3968, 260.8777, 258.3588, 257.3963, 255.0057, 
    253.9391, 252.9292, 252.0075, 249.9703, 248.5218, 247.8825, 249.2084, 
    252.4089,
  268.5077, 266.1537, 263.7839, 260.2437, 258.5033, 256.8735, 254.3288, 
    253.5717, 252.7085, 250.3371, 248.9609, 247.9261, 246.9056, 248.2149, 
    250.9693,
  267.8593, 266.0175, 264.1422, 263.0345, 262.2167, 260.0719, 256.8517, 
    253.2016, 252.131, 250.0462, 249.1954, 251.8487, 255.5269, 259.2943, 
    262.5532,
  270.3114, 268.5162, 266.3263, 264.1553, 262.5403, 259.5383, 256.2863, 
    253.3749, 252.5901, 252.0993, 249.0742, 251.2728, 253.1953, 254.2617, 
    258.4644,
  271.17, 270.2397, 269.2947, 265.1689, 263.4669, 257.7358, 257.2049, 
    254.8015, 253.8655, 252.4809, 251.7879, 250.618, 252.459, 254.649, 257.443,
  271.0068, 269.9183, 269.2499, 264.9904, 263.6909, 260.7135, 255.7112, 
    255.9679, 255.191, 254.3791, 253.1548, 250.9581, 250.6946, 252.5205, 
    255.5545,
  270.5937, 269.2144, 268.4038, 263.918, 263.3325, 262.0988, 258.9945, 
    253.5134, 251.7662, 255.7413, 255.0027, 252.1436, 249.877, 251.2633, 
    253.5891,
  269.9364, 268.3029, 266.9549, 264.4755, 263.5284, 260.4799, 259.5663, 
    257.5896, 255.5634, 253.1906, 252.6985, 251.7787, 249.9989, 249.8361, 
    252.4592,
  269.0079, 267.1571, 265.4862, 263.3392, 261.1782, 258.0735, 257.6633, 
    256.3822, 255.5045, 253.3023, 252.8707, 251.6877, 250.3836, 248.982, 
    251.4291,
  267.9682, 265.718, 263.588, 260.5223, 258.9753, 256.7677, 255.6597, 
    255.3343, 254.3795, 253.5538, 252.3198, 251.4542, 250.302, 248.6395, 
    251.121,
  266.7851, 264.1371, 261.4202, 257.9205, 256.6585, 255.749, 255.0697, 
    255.0159, 254.0634, 252.9424, 251.6548, 250.9237, 249.6892, 248.6071, 
    250.2869,
  265.4074, 261.6147, 259.1346, 256.9609, 256.0907, 255.2562, 254.3306, 
    254.7809, 253.9808, 252.3472, 250.8647, 250.2868, 248.822, 247.7436, 
    249.2869,
  266.6091, 264.2222, 262.1915, 261.1915, 261.2224, 262.6479, 263.0701, 
    260.9061, 258.2883, 255.854, 254.1857, 251.7507, 253.2388, 257.3641, 
    262.2993,
  267.8582, 265.8863, 263.4494, 261.1082, 261.779, 262.92, 261.3733, 
    258.8203, 256.9759, 254.7647, 252.5884, 252.0505, 254.4376, 257.0894, 
    261.448,
  267.7435, 266.4647, 265.4579, 261.8304, 261.9522, 259.1835, 259.2567, 
    256.8917, 255.0379, 253.4228, 252.7497, 252.0473, 254.6556, 258.6645, 
    262.6993,
  266.7485, 265.3857, 264.416, 261.0306, 260.7213, 259.9982, 254.677, 254.98, 
    253.9238, 253.1729, 252.5499, 252.0963, 255.1103, 258.3456, 261.8972,
  265.8233, 264.4158, 263.2141, 259.5446, 259.9963, 259.6755, 257.7093, 
    251.3793, 249.1042, 253.0355, 252.8471, 252.065, 254.2112, 257.7166, 
    260.9267,
  264.9319, 263.5932, 262.3421, 260.3066, 259.9397, 257.9959, 258.841, 
    257.8146, 254.8043, 253.062, 251.5646, 252.1362, 253.4432, 257.1599, 
    260.0888,
  264.1401, 263.0485, 262.0102, 260.5317, 259.6075, 257.8829, 258.9617, 
    257.4773, 255.352, 253.6731, 253.4808, 252.88, 253.9029, 257.1914, 
    260.0666,
  263.3056, 262.0659, 260.9491, 259.772, 259.2863, 258.3077, 257.8481, 
    256.1367, 254.3011, 253.7512, 253.0299, 253.0777, 254.1523, 257.0358, 
    259.642,
  262.3952, 260.8574, 258.9296, 257.3318, 257.7972, 257.2929, 256.6752, 
    254.718, 253.4934, 252.6713, 252.0077, 252.3787, 253.3943, 256.6562, 
    258.7784,
  260.7357, 258.2584, 257.1274, 256.3495, 256.1882, 256.105, 255.1712, 
    254.8509, 252.8077, 251.0445, 250.9964, 251.5767, 252.3647, 255.7562, 
    258.7146,
  264.6548, 261.737, 259.3122, 257.2602, 257.6242, 257.4892, 256.7143, 
    255.8104, 258.7423, 262.131, 263.5504, 261.6801, 259.5768, 258.0322, 
    255.7952,
  266.985, 264.3835, 260.8419, 257.5658, 258.1796, 258.1781, 258.5355, 
    257.6978, 259.8192, 262.5262, 262.4932, 260.7698, 259.3944, 255.5993, 
    255.027,
  267.739, 266.016, 263.2401, 258.3136, 257.9964, 255.8927, 258.9369, 
    259.2193, 260.3181, 261.7995, 261.1696, 259.8017, 258.7897, 257.2607, 
    256.712,
  267.7135, 265.9185, 263.4369, 258.597, 257.9501, 257.4503, 254.6115, 
    257.395, 258.8933, 259.5462, 258.5521, 258.1267, 258.5689, 257.8848, 
    258.1248,
  267.5824, 265.7769, 263.2332, 258.4442, 257.7973, 257.3927, 257.53, 
    250.8551, 250.2767, 256.2725, 256.5211, 254.7686, 257.1833, 259.1238, 
    259.3009,
  267.2548, 265.9386, 263.3867, 259.9725, 257.9025, 255.7923, 255.8071, 
    255.653, 252.4792, 251.9243, 251.4621, 253.8598, 258.5321, 260.3034, 
    260.3136,
  266.6119, 265.8097, 263.5729, 260.4275, 257.8047, 254.7982, 253.9992, 
    253.3852, 252.7188, 250.9012, 252.1752, 256.561, 260.9955, 262.5242, 
    262.2085,
  265.3577, 264.2994, 262.3271, 259.6171, 256.9927, 255.1051, 253.661, 
    252.9272, 251.882, 253.0745, 255.8376, 260.3652, 262.557, 263.1246, 
    263.2029,
  264.0219, 262.3784, 259.5445, 257.515, 255.9969, 254.9537, 254.5426, 
    254.2362, 254.0307, 255.2016, 258.4944, 262.0287, 262.7379, 262.4004, 
    262.1437,
  261.9854, 259.2388, 257.8523, 256.5927, 255.4976, 254.9378, 254.8789, 
    256.0986, 256.3141, 256.9814, 258.6972, 260.9973, 261.5504, 262.0824, 
    262.708,
  264.93, 259.7987, 258.0457, 257.0601, 258.2005, 259.4262, 260.9911, 
    261.3482, 261.7787, 261.1805, 261.062, 261.8116, 262.7497, 262.986, 
    262.5065,
  267.0902, 262.4737, 259.9731, 257.8004, 258.3785, 259.5837, 261.7665, 
    261.8405, 262.6752, 263.181, 263.9878, 265.1335, 264.8634, 262.5414, 
    262.7039,
  268.0116, 265.7513, 262.791, 258.3896, 258.2171, 257.4667, 261.3367, 
    261.6159, 261.6462, 261.8553, 261.9594, 262.7702, 263.3071, 263.6022, 
    263.3217,
  267.7025, 265.7539, 263.3168, 258.7297, 258.4741, 259.1445, 259.1496, 
    261.5093, 260.5457, 260.1978, 260.0546, 260.2579, 260.9701, 261.6818, 
    262.3804,
  267.4071, 265.4391, 263.098, 258.8793, 258.5592, 258.3149, 259.9065, 
    256.0552, 255.3797, 259.2847, 258.9222, 258.0691, 258.5354, 259.5722, 
    260.9389,
  267.0466, 265.2555, 263.2146, 260.369, 259.0901, 257.6991, 257.9439, 
    257.5509, 255.2195, 256.0881, 256.5976, 257.5457, 257.9251, 257.759, 
    258.9599,
  266.306, 264.835, 262.6082, 260.754, 258.8945, 257.84, 257.3914, 256.5273, 
    255.5968, 254.597, 255.0276, 256.6017, 258.028, 257.5565, 259.1049,
  265.5339, 263.9991, 261.3604, 259.3135, 258.4607, 258.214, 258.332, 
    258.3661, 257.3721, 255.7443, 255.8512, 255.3214, 256.6115, 259.4441, 
    260.7389,
  264.8247, 262.9546, 259.7076, 257.8872, 257.378, 257.5035, 259.2968, 
    259.5595, 259.5474, 258.5747, 259.195, 259.2529, 259.544, 259.7252, 
    261.9073,
  263.155, 260.0012, 258.2192, 257.0402, 257.0079, 257.2299, 259.3079, 
    262.1947, 262.0242, 262.0948, 262.7861, 262.9039, 262.6805, 262.1653, 
    262.4634,
  264.233, 262.3752, 260.5396, 260.254, 261.4189, 259.8481, 258.6284, 
    258.1313, 259.3589, 261.0743, 261.8169, 259.5576, 255.2877, 256.7964, 
    256.3045,
  267.4678, 265.094, 262.7737, 260.9155, 260.8071, 259.378, 258.9233, 
    258.0876, 258.2896, 260.0013, 261.0689, 262.2809, 259.1547, 254.9005, 
    255.6137,
  269.236, 268.2868, 266.2677, 261.5289, 259.6618, 257.1908, 259.31, 
    258.4855, 258.5732, 258.4086, 259.4246, 262.3977, 261.2336, 258.77, 
    257.0482,
  269.5071, 268.498, 266.9405, 262.0632, 260.5764, 259.2693, 256.7033, 
    258.2303, 259.0102, 258.5081, 257.8739, 260.5041, 263.5559, 261.6998, 
    258.6493,
  269.7415, 268.4231, 266.9559, 262.3975, 261.4364, 260.0876, 259.5093, 
    255.3773, 255.7172, 259.245, 257.9209, 258.825, 261.8913, 262.9095, 
    261.2867,
  269.986, 268.7345, 267.0914, 264.468, 262.0935, 260.0689, 259.5558, 
    260.2973, 260.4688, 259.4137, 257.4871, 258.1761, 260.4938, 262.6685, 
    262.8307,
  270.0692, 269.1264, 267.3361, 264.661, 261.6927, 259.9304, 259.235, 
    260.5973, 262.1213, 260.8362, 258.3251, 258.3387, 260.0128, 262.5263, 
    263.7325,
  270.5672, 269.8119, 267.4983, 263.963, 261.4612, 259.2839, 258.5577, 
    260.839, 263.0754, 262.6805, 259.8363, 258.9247, 259.5843, 261.9707, 
    263.065,
  271.6233, 270.3221, 267.1163, 263.6122, 260.9059, 258.5681, 257.9917, 
    260.5726, 263.0197, 263.6145, 261.7533, 260.74, 260.6034, 261.8361, 
    261.6152,
  271.8538, 269.0517, 266.0331, 263.2818, 261.2706, 257.8244, 257.2671, 
    260.0182, 262.6779, 264.0722, 263.3905, 262.4069, 262.4049, 262.6525, 
    262.1814,
  267.1902, 266.6334, 266.291, 265.0561, 264.1751, 263.7348, 262.7185, 
    260.7359, 258.7545, 260.3114, 260.4605, 259.288, 258.4857, 258.3192, 
    258.4275,
  270.4099, 269.388, 267.8432, 266.5227, 266.2763, 265.0081, 263.9671, 
    261.08, 258.1677, 261.043, 261.076, 260.1775, 259.8501, 256.6776, 257.5177,
  272.4998, 271.9823, 271.1466, 268.4067, 266.2166, 264.3927, 265.1131, 
    261.6838, 258.3999, 262.0446, 261.4222, 261.4996, 259.5601, 259.4868, 
    258.2078,
  273.3175, 272.8467, 272.3176, 269.748, 268.3607, 267.0824, 263.1399, 
    259.7308, 257.7347, 261.4434, 261.8707, 262.0338, 261.2751, 259.4617, 
    257.5325,
  274.2041, 273.1792, 272.5985, 270.3607, 268.8918, 266.6479, 264.0053, 
    253.8216, 254.2205, 260.7638, 262.0098, 262.1348, 262.931, 260.3235, 
    259.0662,
  274.7307, 273.5697, 272.173, 270.419, 268.231, 264.7089, 260.0392, 
    257.5594, 257.3531, 261.043, 261.7794, 262.0945, 263.4337, 262.4455, 
    261.343,
  274.6983, 273.6788, 271.9044, 269.3853, 266.2359, 261.8481, 258.9006, 
    259.2152, 259.9688, 263.047, 262.6077, 262.2369, 263.2193, 264.1888, 
    263.7099,
  274.344, 273.3081, 270.933, 267.2616, 263.804, 259.3073, 258.8409, 
    259.5076, 260.6839, 263.5439, 262.8084, 262.149, 262.7612, 263.4131, 
    264.1024,
  273.782, 272.2814, 269.4686, 264.3478, 261.0246, 258.149, 258.3192, 
    259.5803, 262.4647, 264.0154, 263.1958, 262.5535, 262.4857, 262.9082, 
    262.8861,
  272.5447, 270.7863, 267.6837, 264.048, 261.2245, 256.88, 257.6491, 
    260.1329, 262.7271, 263.0237, 262.8773, 262.8138, 263.1463, 263.4617, 
    263.09,
  269.4643, 269.1144, 269.2739, 268.5763, 268.3438, 268.6751, 268.4591, 
    268.0544, 266.225, 261.2173, 257.841, 261.337, 260.7775, 260.0804, 
    259.7284,
  271.4515, 270.8127, 269.0937, 267.6316, 266.4344, 266.9574, 267.6015, 
    266.3813, 263.5592, 259.1482, 258.1742, 262.2429, 261.6926, 259.1724, 
    259.506,
  272.5055, 271.0524, 269.0565, 265.445, 264.3543, 262.5692, 264.4679, 
    263.1255, 259.1586, 258.2541, 260.6825, 262.0151, 262.1763, 262.5757, 
    261.7433,
  272.8146, 270.9337, 268.8914, 263.8364, 262.4496, 261.4526, 258.9347, 
    259.8076, 257.6802, 258.4962, 259.6914, 261.8502, 262.628, 262.8448, 
    261.8253,
  272.8758, 270.2964, 268.2277, 262.7747, 261.7084, 259.278, 259.4064, 
    253.7329, 252.7744, 258.6472, 261.5703, 262.0703, 262.6812, 262.6844, 
    263.3712,
  273.255, 270.5442, 268.3647, 264.5291, 262.6657, 259.44, 258.5515, 
    259.3237, 258.9601, 259.0239, 261.8296, 261.383, 262.4247, 263.1871, 
    263.2446,
  273.7768, 271.4614, 269.5316, 265.6925, 263.387, 259.6313, 258.8413, 
    260.0929, 261.2668, 262.7122, 262.9821, 262.1047, 263.2045, 263.6657, 
    262.7958,
  274.2282, 272.6706, 270.5985, 266.4605, 264.2069, 259.4842, 258.7429, 
    260.6425, 262.6126, 263.4492, 263.5206, 262.8319, 264.0222, 263.9033, 
    262.7769,
  274.4732, 273.0913, 270.893, 267.4644, 264.9216, 260.4033, 258.3741, 
    260.9745, 263.0791, 263.9746, 263.9041, 263.8653, 264.8188, 264.5468, 
    263.7904,
  273.689, 272.139, 270.1712, 268.7618, 265.3033, 259.4227, 257.6109, 
    261.3698, 263.4109, 263.727, 264.3596, 265.0718, 265.4631, 264.5659, 
    262.9426,
  268.2651, 264.0588, 263.2116, 261.5948, 260.2274, 260.4765, 259.0799, 
    260.4388, 261.3661, 261.3905, 260.9057, 262.1464, 261.9961, 261.2665, 
    260.8185,
  269.8784, 266.856, 265.3857, 263.5419, 261.9787, 259.7937, 259.3201, 
    257.8517, 259.3829, 260.3821, 260.5251, 261.6436, 261.3065, 259.0103, 
    259.5717,
  271.6071, 270.8357, 269.5771, 265.6915, 263.8864, 259.9409, 259.0165, 
    258.9182, 260.2637, 260.2888, 260.6885, 262.2578, 262.1886, 262.022, 
    261.5752,
  273.0178, 272.2629, 271.3229, 267.4357, 266.6267, 263.8887, 258.4653, 
    258.1343, 260.9337, 262.0209, 262.5679, 263.415, 263.56, 263.9708, 
    263.9321,
  274.4101, 273.0027, 271.6719, 269.0598, 268.322, 265.6558, 260.3134, 
    256.7069, 257.9854, 263.2372, 263.8709, 263.6718, 263.9983, 263.8444, 
    264.0588,
  275.1147, 273.629, 271.5411, 270.4147, 268.1928, 265.34, 261.206, 261.6975, 
    262.4546, 263.5784, 263.472, 263.0806, 263.5114, 263.1309, 263.1,
  275.2271, 273.8262, 271.2518, 270.2942, 266.6931, 263.1376, 260.6338, 
    262.3727, 264.0269, 263.9341, 263.2346, 263.0751, 263.3218, 263.2774, 
    263.4377,
  275.137, 273.086, 270.1706, 268.9478, 264.6707, 261.5073, 260.8919, 
    263.6644, 263.864, 263.3511, 262.7611, 263.2074, 263.4621, 263.9122, 
    264.0376,
  274.999, 272.1684, 268.4761, 266.9046, 261.8219, 259.7162, 261.5113, 
    264.4559, 263.9478, 262.8399, 262.5566, 262.8425, 263.1753, 264.0266, 
    264.5606,
  273.8262, 270.865, 267.0406, 265.2418, 259.5867, 259.5549, 262.0022, 
    264.9378, 263.8637, 262.217, 261.913, 262.282, 262.6198, 263.0783, 
    263.9289,
  270.2596, 269.9516, 270.0226, 268.6472, 266.3797, 264.9185, 261.2017, 
    261.0907, 261.6088, 262.1042, 261.9132, 262.2983, 262.5744, 261.1701, 
    260.2258,
  271.2899, 271.4973, 270.1257, 267.8747, 266.1667, 262.9098, 262.1437, 
    259.9002, 260.0486, 260.5987, 261.8831, 262.7776, 263.1164, 261.8347, 
    261.0911,
  272.8908, 271.456, 269.8612, 267.3045, 264.8492, 262.2203, 261.5839, 
    261.6176, 261.6506, 262.561, 262.4851, 262.7502, 262.8694, 262.4094, 
    261.8777,
  273.4075, 271.6103, 269.5136, 266.814, 263.8842, 261.8271, 258.675, 
    261.4672, 262.5238, 262.535, 262.2848, 262.3526, 262.5563, 262.5871, 
    262.8038,
  272.981, 271.6674, 268.9492, 265.9669, 262.9498, 261.9397, 261.5218, 
    257.3104, 257.9999, 262.2677, 262.3997, 262.1203, 262.7711, 263.0943, 
    262.63,
  273.8806, 271.5112, 268.287, 265.6049, 262.9671, 261.495, 261.3922, 
    261.1192, 259.6722, 260.5274, 261.2893, 262.5227, 263.6497, 263.8307, 
    263.9634,
  274.5922, 271.482, 268.0668, 265.2299, 262.1632, 261.8076, 261.3353, 
    260.7992, 260.4007, 260.7895, 261.1568, 262.2605, 263.4153, 264.4865, 
    264.6256,
  274.8052, 271.3638, 267.5089, 263.7213, 261.7629, 263.129, 261.0613, 
    260.541, 260.7324, 261.0496, 261.1364, 261.695, 262.8958, 264.3154, 264.79,
  275.157, 271.8999, 266.5314, 262.5711, 261.9874, 262.2777, 260.7438, 
    261.1527, 261.2229, 261.3459, 260.8234, 260.8555, 262.0262, 263.6374, 
    265.0452,
  274.399, 271.3798, 267.0261, 263.3735, 261.826, 262.742, 260.9833, 262.386, 
    261.302, 259.6263, 259.4465, 260.3336, 261.2979, 263.0758, 264.6662,
  267.3489, 264.7579, 263.7476, 259.89, 258.296, 258.0068, 257.3409, 
    257.9401, 258.4245, 259.2721, 259.1343, 258.7734, 260.9328, 261.3932, 
    260.7517,
  269.4045, 266.6896, 264.8686, 261.4671, 260.0711, 258.8546, 258.649, 
    258.9424, 259.2523, 259.1982, 258.389, 259.3232, 259.892, 260.0403, 
    259.5458,
  271.8315, 270.088, 267.7486, 262.8961, 260.8853, 258.4828, 260.0219, 
    259.8638, 259.7465, 260.2838, 259.5645, 259.5229, 260.9005, 261.2612, 
    261.0596,
  273.1933, 271.7346, 269.8424, 265.8352, 262.7744, 260.9842, 258.3581, 
    260.436, 260.8551, 261.049, 260.3869, 259.8814, 260.6812, 261.2509, 
    260.991,
  274.6483, 272.709, 271.0602, 267.7965, 264.9916, 262.7684, 261.5337, 
    256.9418, 256.999, 261.7437, 261.1306, 260.247, 260.6718, 260.5964, 
    261.2603,
  275.614, 273.8341, 271.505, 269.0878, 267.1848, 264.9169, 262.5884, 
    261.6315, 260.5215, 260.3242, 260.2358, 260.3642, 260.883, 260.3905, 
    261.3536,
  275.8164, 274.5983, 272.4118, 270.2673, 267.8756, 266.0158, 263.9476, 
    262.9184, 262.1757, 261.691, 261.3456, 260.873, 260.225, 260.545, 262.0638,
  275.9245, 274.7977, 272.8532, 270.6558, 268.6453, 267.3315, 266.0509, 
    264.6796, 264.0554, 263.49, 262.4074, 261.0359, 259.9335, 260.8385, 
    262.3643,
  275.6501, 274.5679, 272.5442, 270.6142, 269.2864, 268.3708, 267.1428, 
    266.3188, 265.7294, 264.8285, 263.0589, 261.1873, 260.2999, 260.4386, 
    262.4598,
  274.3379, 273.0635, 272.6931, 271.9374, 270.2196, 269.6407, 268.3251, 
    267.9345, 267.0531, 265.1435, 262.1619, 260.5092, 259.0667, 260.098, 
    261.5261,
  270.6204, 269.4179, 268.5792, 267.2238, 265.7935, 263.7209, 262.1031, 
    260.4995, 260.9237, 260.4006, 260.5896, 258.6754, 258.2614, 257.7036, 
    255.4412,
  272.4157, 271.0936, 269.5469, 267.6964, 265.5432, 264.8337, 262.5788, 
    262.3628, 262.7642, 261.6199, 261.7164, 260.3065, 259.5696, 258.4951, 
    257.8242,
  274.204, 273.0383, 271.689, 268.6355, 267.4947, 264.7038, 266.1361, 
    265.5562, 264.9031, 264.4136, 264.0581, 263.0779, 262.2731, 261.4707, 
    260.7705,
  275.3382, 274.271, 273.2038, 271.0677, 269.7902, 267.4594, 265.4877, 
    267.2415, 266.7515, 266.4117, 265.6108, 264.5513, 263.8098, 263.2018, 
    261.8291,
  276.0525, 274.1257, 273.1562, 272.0076, 271.7005, 270.9648, 269.8989, 
    266.4958, 265.9594, 269.4246, 269.2005, 268.24, 267.1516, 265.7797, 
    264.0332,
  276.1969, 274.8064, 272.7407, 271.7943, 271.922, 272.1432, 271.8265, 
    271.4204, 271.009, 270.7443, 270.0074, 269.0271, 268.3887, 267.5564, 
    266.4038,
  275.6308, 274.8492, 273.3311, 271.9179, 272.0342, 272.2785, 272.2194, 
    271.5871, 270.2233, 269.151, 268.3281, 267.9061, 267.8296, 267.4664, 
    266.9565,
  276.424, 275.1542, 273.4064, 272.4293, 272.417, 272.1422, 270.994, 
    269.1442, 267.7336, 267.2632, 266.8453, 266.7376, 266.2245, 265.9715, 
    265.9588,
  276.4338, 274.9882, 272.7273, 272.3555, 271.464, 269.7853, 267.7525, 
    266.3424, 265.9087, 265.749, 264.2409, 264.0835, 264.3513, 264.2151, 
    264.9076,
  275.2657, 272.9807, 272.2334, 271.1721, 269.4182, 266.4548, 264.6425, 
    264.2202, 263.8239, 262.3957, 262.2152, 262.7209, 263.1959, 263.0921, 
    263.8165,
  272.1447, 271.4751, 272.2172, 271.3672, 270.4485, 270.0905, 269.0915, 
    267.0117, 265.935, 265.2677, 265.9422, 266.6743, 265.7579, 265.01, 
    263.7432,
  272.8898, 272.4826, 272.1141, 271.3221, 270.9199, 271.166, 269.87, 
    268.1256, 266.751, 266.3945, 266.9128, 267.4829, 267.3217, 265.3666, 
    264.2785,
  274.1069, 273.1724, 272.5347, 271.1988, 271.3394, 269.1417, 270.1128, 
    268.9848, 267.4601, 267.5041, 267.9395, 268.8862, 269.1901, 268.9147, 
    266.7717,
  274.7023, 273.5936, 272.3903, 270.6683, 270.3362, 268.9366, 266.8988, 
    267.334, 267.277, 267.3437, 267.356, 268.1081, 268.332, 268.2532, 267.4648,
  274.8674, 272.9093, 271.4296, 269.3858, 268.252, 267.5133, 266.9883, 
    263.5903, 263.6505, 265.434, 264.5335, 263.9443, 263.565, 263.5519, 
    264.7007,
  274.7841, 272.6512, 270.1115, 268.0126, 266.4514, 264.9717, 264.7332, 
    264.8199, 264.1855, 261.6878, 260.2079, 259.4048, 259.4401, 259.2477, 
    260.6758,
  274.2799, 272.0856, 269.2907, 266.4778, 264.2065, 262.3954, 261.3217, 
    261.6805, 261.3942, 260.897, 259.8129, 258.8398, 259.7471, 259.3862, 
    259.6942,
  273.6047, 271.0963, 267.428, 264.2512, 262.3223, 260.4829, 259.6647, 
    260.1551, 260.8318, 261.1738, 260.8897, 260.9122, 261.0294, 261.3008, 
    261.6951,
  272.3732, 269.1849, 264.7284, 261.5549, 261.3513, 259.8933, 259.5166, 
    260.7034, 261.3745, 261.7779, 261.4241, 260.9579, 261.0257, 261.1307, 
    261.8147,
  270.8119, 267.3148, 262.762, 261.3558, 260.4676, 259.6173, 259.6153, 
    260.5948, 261.8101, 261.4316, 261.3402, 260.9326, 260.5979, 261.0409, 
    261.3142,
  269.0364, 267.2206, 266.1548, 265.6266, 265.4963, 264.7079, 262.7419, 
    262.2208, 262.0627, 262.5691, 262.9968, 263.6166, 264.5054, 266.0144, 
    267.5821,
  269.054, 267.1052, 264.5534, 263.7627, 264.1226, 262.1498, 260.9377, 
    260.8267, 260.962, 260.8097, 261.8317, 262.9395, 263.6764, 264.069, 266.11,
  269.9368, 268.0943, 265.4974, 261.7906, 261.1899, 258.59, 260.0787, 
    260.3642, 261.0537, 260.3355, 259.9738, 260.8836, 261.5371, 262.7064, 
    265.2146,
  270.1396, 268.6663, 266.5048, 262.5229, 261.0776, 259.4691, 257.1383, 
    258.9717, 260.6044, 261.0823, 260.0727, 259.5817, 259.3958, 260.5587, 
    262.3063,
  270.8018, 269.1819, 267.3421, 263.5688, 261.601, 260.8369, 259.3876, 
    255.3704, 257.3726, 261.3294, 260.7104, 259.5608, 259.2288, 258.6414, 
    259.0049,
  271.9046, 270.3123, 267.966, 264.9968, 262.6606, 260.0813, 260.471, 
    261.2418, 261.687, 260.7741, 259.8353, 259.6276, 260.451, 258.9062, 
    258.3949,
  272.752, 271.4276, 268.8732, 265.584, 262.9081, 259.9782, 259.8554, 
    261.2517, 261.7276, 261.8251, 261.2511, 260.6538, 261.6692, 261.4149, 
    260.6325,
  273.644, 272.0563, 269.2601, 265.5718, 263.9164, 261.1353, 259.7887, 
    261.1295, 262.1288, 262.1843, 261.8522, 261.5657, 261.8601, 262.669, 
    262.7569,
  273.9534, 272.317, 269.0086, 264.8965, 264.5392, 261.8176, 260.1862, 
    261.4402, 262.4006, 263.195, 262.0778, 261.9924, 261.1843, 261.6887, 
    262.5706,
  274.1604, 271.6132, 269.2427, 266.628, 265.5262, 263.2173, 259.7638, 
    260.8155, 262.2512, 262.0676, 261.47, 261.5116, 260.724, 261.4331, 
    262.1452,
  269.086, 266.5672, 265.0927, 263.8658, 263.3246, 263.1218, 260.9416, 
    259.622, 259.4039, 259.7263, 260.4941, 258.2668, 258.7893, 260.7081, 
    262.3368,
  270.8596, 269.3852, 267.8452, 266.144, 265.3013, 263.5812, 262.3623, 
    261.1793, 260.3876, 259.6496, 259.0727, 257.4846, 257.5231, 259.7924, 
    259.5781,
  272.8316, 271.7643, 270.8459, 268.3157, 266.6501, 263.6658, 263.6864, 
    262.4297, 261.7128, 260.7697, 259.7483, 258.4756, 258.0871, 260.201, 
    259.7836,
  274.5441, 273.3671, 272.6542, 270.8219, 269.1385, 266.7631, 262.8304, 
    262.151, 261.8156, 261.1299, 260.5491, 258.6869, 258.2965, 260.3549, 
    259.6153,
  275.8396, 274.0042, 273.4817, 272.0937, 270.6974, 269.0513, 266.6435, 
    260.251, 258.8863, 261.9702, 260.8546, 258.7788, 258.5362, 260.1957, 
    260.727,
  276.2555, 275.0387, 273.37, 272.4686, 271.8242, 270.1702, 268.3011, 
    265.7316, 263.2816, 261.7756, 260.5829, 258.6678, 258.4917, 258.7715, 
    261.7944,
  276.406, 275.4234, 274.0531, 272.8156, 272.2255, 270.4789, 268.8444, 
    266.3226, 262.8329, 261.1627, 260.6639, 259.7743, 258.6096, 259.6232, 
    261.5787,
  276.5786, 275.318, 273.9857, 273.0137, 272.3008, 270.8054, 268.4252, 
    265.712, 262.6349, 261.73, 261.131, 259.9101, 258.8966, 260.4125, 261.2671,
  276.3051, 275.3934, 273.248, 272.9948, 271.9814, 270.2745, 268.4937, 
    265.4548, 263.1953, 262.4911, 259.7969, 258.7823, 258.2614, 259.0315, 
    261.571,
  275.4579, 273.5409, 272.9316, 272.4455, 271.219, 269.804, 267.9955, 
    265.3622, 263.569, 260.6036, 257.6863, 257.9485, 257.6846, 258.3194, 
    261.1895,
  272.5892, 271.7738, 271.4408, 270.502, 269.9445, 269.6552, 269.4925, 
    269.6932, 268.8223, 266.6412, 265.8646, 263.5471, 261.2234, 259.1777, 
    256.7918,
  272.9832, 272.3627, 271.9388, 271.4891, 271.0974, 270.5215, 269.7596, 
    269.7207, 269.3819, 267.5918, 266.3263, 263.9987, 260.8102, 258.9039, 
    257.0591,
  274.0335, 273.0909, 272.4033, 271.6401, 270.9882, 269.6621, 270.4885, 
    269.6954, 268.6714, 266.6992, 265.0718, 263.6271, 260.6675, 260.0635, 
    259.6622,
  274.8824, 273.7166, 272.7745, 271.1075, 270.1233, 270.0682, 268.2935, 
    268.1688, 267.0984, 265.5413, 264.0644, 261.8808, 259.9694, 260.0058, 
    260.0176,
  275.283, 273.2341, 272.346, 270.2378, 269.3245, 268.6907, 267.6699, 
    263.5474, 261.9965, 263.9766, 262.0836, 260.8062, 260.1747, 259.8465, 
    260.6737,
  275.3006, 273.2296, 271.3556, 269.3855, 268.4331, 267.1093, 265.9352, 
    264.5375, 262.9075, 262.187, 261.2786, 260.2746, 260.0048, 259.4413, 
    259.5405,
  275.0617, 272.9015, 271.0532, 268.9351, 267.2924, 265.477, 264.0339, 
    262.6993, 261.5714, 259.5414, 259.7124, 260.1628, 259.8702, 259.5643, 
    259.4483,
  274.6972, 272.5257, 269.996, 267.3968, 265.6775, 264.2981, 263.4433, 
    262.0448, 261.115, 259.8778, 259.1027, 259.3617, 260.1142, 260.219, 
    260.3001,
  273.7454, 271.576, 267.6852, 265.5891, 263.9542, 263.2187, 262.8809, 
    262.0507, 261.3212, 260.4747, 258.7449, 258.1561, 257.6123, 258.5103, 
    260.6004,
  272.0311, 269.0398, 265.8616, 263.2823, 261.5556, 260.4297, 260.2063, 
    260.6635, 259.9373, 258.0945, 256.3812, 256.4919, 256.2172, 256.9316, 
    259.4018,
  269.403, 267.4637, 266.7998, 266.6172, 265.613, 262.5879, 261.0197, 
    261.7608, 262.9716, 263.9622, 265.308, 266.4991, 266.8691, 266.5504, 
    264.6674,
  269.5456, 267.3624, 265.4101, 264.7772, 264.2968, 261.1261, 260.1141, 
    260.3481, 261.1501, 262.6207, 264.4621, 267.7153, 267.6117, 265.4653, 
    263.8897,
  270.1505, 268.1882, 265.8394, 263.1969, 262.1168, 259.7462, 260.1519, 
    260.1226, 260.808, 261.7582, 263.7161, 266.3436, 267.9802, 265.9098, 
    263.5892,
  270.3495, 268.3235, 266.075, 262.8588, 261.3376, 260.5962, 257.5781, 
    259.5334, 260.2214, 260.8386, 262.3777, 264.3734, 264.9616, 263.9091, 
    263.2738,
  270.512, 268.2575, 266.0992, 263.0341, 262.0026, 261.6282, 261.2571, 
    256.3289, 256.4743, 260.2644, 261.3174, 262.5579, 263.3815, 263.6924, 
    264.2803,
  270.6982, 268.3589, 265.6869, 263.8668, 262.0314, 261.3165, 261.3429, 
    261.1759, 259.7733, 259.4954, 260.0444, 261.3857, 262.249, 262.4402, 
    262.0873,
  270.7986, 268.4146, 265.6615, 263.3406, 261.5088, 261.2599, 261.1529, 
    261.2607, 260.9792, 259.024, 259.4026, 260.5094, 260.6665, 260.89, 
    260.6372,
  270.2549, 267.6338, 264.8726, 262.0835, 261.1133, 260.9495, 261.0305, 
    261.1197, 261.0703, 259.6034, 258.5832, 260.0481, 260.7498, 260.5468, 
    260.8895,
  269.5012, 266.9642, 263.41, 261.942, 260.9754, 260.4467, 260.9504, 
    261.5567, 261.5399, 260.6762, 259.1023, 258.5985, 258.985, 259.855, 
    259.8839,
  268.0254, 266.0018, 263.8706, 262.4009, 261.1588, 260.2192, 260.3877, 
    261.2491, 260.9355, 259.3611, 258.1467, 256.7473, 257.5387, 258.3767, 
    259.3232,
  268.1689, 266.8106, 265.8117, 264.9436, 263.6693, 260.5914, 259.0464, 
    257.7654, 257.7948, 259.3616, 260.6971, 262.7978, 264.0251, 265.3609, 
    265.514,
  270.2041, 269.109, 266.9404, 265.4511, 262.8903, 260.2225, 259.6049, 
    258.7608, 258.3703, 258.6781, 260.8434, 263.5048, 265.5284, 265.2923, 
    265.1112,
  271.3317, 270.6494, 268.9279, 265.3832, 262.4652, 259.6816, 259.7809, 
    260.1473, 259.52, 259.8654, 261.2219, 263.9017, 266.9247, 266.7741, 
    266.6082,
  271.7763, 270.8646, 269.3014, 266.0199, 262.867, 260.2761, 256.8122, 
    259.6664, 260.429, 260.4286, 260.8365, 263.3321, 266.4949, 267.4504, 
    267.017,
  272.2303, 270.764, 269.2025, 266.2141, 263.4436, 260.8819, 259.7185, 
    255.6405, 256.3806, 260.2257, 260.4974, 261.9352, 264.3579, 266.6429, 
    266.944,
  272.3991, 270.9527, 268.7233, 266.3269, 263.4569, 261.7292, 259.9482, 
    259.5706, 258.9465, 259.3267, 259.8234, 260.8127, 261.9082, 263.4494, 
    264.7715,
  272.5103, 270.9916, 268.5695, 265.5257, 263.3517, 261.9593, 260.1025, 
    260.2205, 259.4232, 259.0316, 259.5631, 260.3579, 261.2235, 261.7263, 
    262.2697,
  272.5105, 270.79, 267.7874, 264.7904, 263.1225, 261.7505, 260.7545, 
    260.763, 260.2049, 259.5513, 259.0887, 259.5107, 260.9173, 261.5241, 
    262.0576,
  272.4095, 270.4678, 267.0109, 264.301, 262.6234, 261.154, 261.155, 
    261.6485, 261.1553, 260.0804, 259.9076, 259.5065, 260.1147, 261.1485, 
    261.9484,
  272.1055, 269.6937, 266.3496, 264.0303, 262.3272, 260.8844, 260.5881, 
    261.5176, 261.2385, 259.9493, 259.1621, 259.5254, 260.0981, 260.9245, 
    261.9762,
  271.7288, 268.1551, 263.5078, 263.5694, 262.7525, 261.5359, 257.8589, 
    257.9079, 257.6686, 259.2029, 259.5362, 260.3482, 262.0464, 264.2514, 
    266.8683,
  271.8179, 268.4246, 264.1888, 262.5755, 262.1557, 260.5175, 258.4266, 
    258.6733, 258.7195, 258.0725, 259.1743, 261.9695, 263.1024, 263.244, 
    264.5304,
  272.2219, 269.1682, 266.1993, 262.1599, 260.7491, 259.0102, 259.0741, 
    259.957, 260.418, 260.0105, 259.5886, 262.5234, 263.88, 264.9399, 264.9958,
  272.3603, 268.9354, 266.647, 262.9471, 261.1374, 258.7857, 256.7949, 
    259.9915, 261.0438, 261.3091, 261.01, 261.871, 263.2149, 264.6081, 264.134,
  272.1626, 268.443, 266.313, 263.2021, 261.795, 260.8259, 258.8184, 
    255.8956, 256.7447, 261.3536, 261.8415, 262.3269, 262.9918, 264.4745, 
    266.8719,
  272.0524, 268.4844, 265.9597, 263.3864, 262.166, 261.9887, 260.8192, 
    260.5442, 260.6517, 261.1766, 261.7175, 262.8937, 263.1685, 262.651, 
    265.7882,
  271.922, 268.3162, 264.9962, 262.4519, 261.9185, 262.2045, 262.0143, 
    261.9745, 261.7945, 261.5113, 262.035, 263.201, 264.5136, 263.717, 
    263.9516,
  271.7729, 267.7939, 264.1687, 262.0171, 261.6521, 262.17, 262.7632, 
    262.8357, 262.4381, 261.7854, 262.0798, 263.4843, 265.0508, 265.6538, 
    264.8441,
  271.4079, 267.4129, 263.4026, 261.7586, 261.4398, 262.0309, 263.1886, 
    263.5572, 262.9794, 262.3209, 262.3464, 263.4718, 265.3284, 266.7243, 
    266.4077,
  270.9323, 266.7857, 262.6794, 262.1686, 261.5721, 261.9681, 263.1274, 
    263.9784, 263.2089, 262.0243, 262.1195, 263.2553, 264.8726, 266.9664, 
    268.0623,
  271.6234, 265.8669, 262.584, 260.8815, 258.5218, 258.9956, 260.189, 
    261.4783, 261.4774, 261.7437, 261.9089, 261.8585, 262.0981, 264.3721, 
    267.7609,
  268.7686, 264.3297, 261.9579, 260.2446, 260.0421, 259.5273, 261.6969, 
    261.8187, 261.902, 259.9052, 261.33, 263.0865, 262.0926, 262.9822, 
    266.1932,
  268.5889, 266.0939, 264.0024, 261.9637, 260.534, 258.4281, 261.9642, 
    263.3227, 263.7216, 263.0868, 261.3606, 263.303, 262.6071, 263.318, 
    266.5389,
  268.725, 266.926, 265.5059, 262.8702, 262.2198, 260.8583, 259.8922, 
    263.2645, 263.9724, 264.1348, 263.5172, 264.7801, 263.641, 261.5522, 
    265.9402,
  268.9853, 266.9997, 265.5782, 263.2062, 262.7887, 262.9271, 262.5408, 
    258.9157, 259.4615, 264.0749, 264.9968, 266.303, 264.6769, 260.6486, 
    265.2613,
  268.9878, 267.1304, 265.2989, 263.5133, 263.0806, 262.9004, 262.832, 
    262.5751, 262.5273, 263.7613, 265.5283, 267.4233, 266.0498, 263.436, 
    264.3372,
  269.105, 267.023, 264.5146, 262.9828, 263.0262, 262.8425, 262.5238, 
    262.5559, 262.6211, 263.8812, 265.782, 267.7209, 267.3311, 264.2491, 
    262.9429,
  269.5928, 266.7457, 263.7178, 262.6276, 263.016, 262.8434, 262.3911, 
    262.0119, 262.0302, 263.3509, 265.1876, 266.8792, 267.9844, 265.0257, 
    264.4084,
  269.7345, 265.9563, 262.6508, 262.338, 263.0494, 262.1934, 261.8737, 
    262.292, 262.1953, 263.1495, 264.4536, 266.1754, 267.4397, 265.9247, 
    264.8994,
  269.5924, 265.2956, 261.7368, 262.9872, 263.2486, 261.4512, 261.155, 
    261.7601, 261.6351, 261.8156, 263.4933, 265.1103, 267.1502, 268.7296, 
    265.52,
  266.9715, 264.3802, 262.4413, 260.2188, 259.9118, 258.8592, 260.2746, 
    261.4491, 263.2313, 264.0565, 265.1755, 265.4265, 264.7484, 264.7025, 
    264.6069,
  265.873, 263.8839, 262.3491, 261.2892, 260.9844, 260.5793, 262.03, 
    263.5017, 264.4438, 262.9994, 265.5496, 266.298, 265.9511, 263.9493, 
    264.494,
  267.5456, 266.4258, 264.7249, 262.5564, 261.3818, 259.2111, 262.8142, 
    263.9835, 265.143, 265.9218, 266.0018, 266.6654, 265.9888, 264.7648, 
    265.6706,
  268.3611, 267.1663, 266.2241, 263.0303, 261.641, 261.0155, 259.9987, 
    263.6234, 265.5284, 266.3273, 266.4982, 266.5367, 265.4674, 264.5837, 
    267.4203,
  268.5689, 266.9539, 266.3458, 263.709, 262.1542, 261.6152, 261.4016, 
    260.0526, 261.2455, 266.0823, 266.5928, 266.4748, 265.4021, 264.9384, 
    268.3478,
  268.7263, 267.1374, 265.8557, 264.1219, 262.1958, 261.3083, 261.7018, 
    262.4582, 263.9843, 265.4765, 266.5543, 266.9015, 265.5878, 265.1948, 
    267.9183,
  269.0573, 267.5758, 265.6168, 263.7455, 262.5421, 261.2387, 262.0012, 
    262.9364, 263.995, 265.2958, 266.1211, 267.3924, 266.2388, 265.4549, 
    267.1547,
  269.9062, 268.0288, 264.3766, 262.2862, 262.7859, 261.3007, 261.9094, 
    263.0168, 263.3975, 264.5099, 265.2687, 267.0643, 267.3783, 266.0455, 
    266.5787,
  270.9937, 268.6064, 263.8056, 261.5176, 261.9762, 260.9832, 261.5119, 
    263.7634, 264.1238, 264.6478, 264.212, 266.4765, 267.852, 267.1177, 
    266.1757,
  271.596, 269.058, 263.1549, 262.7276, 261.9448, 260.4334, 260.5683, 
    263.1638, 263.9373, 263.8138, 263.0915, 264.6403, 267.7993, 268.3198, 
    266.4289,
  265.3112, 263.828, 261.2449, 261.6547, 260.6727, 260.2648, 261.1242, 
    264.4094, 265.7972, 265.6702, 266.9361, 267.1805, 266.763, 266.5381, 
    266.2282,
  266.4032, 263.8776, 263.0836, 262.3542, 262.2015, 260.599, 261.0667, 
    264.5747, 265.6135, 266.403, 267.2948, 267.4158, 266.9963, 265.3853, 
    265.5143,
  269.2964, 267.8427, 265.5583, 262.6277, 261.5797, 259.6185, 261.5543, 
    263.2838, 265.6105, 266.6832, 267.2695, 267.6223, 267.1934, 266.7897, 
    266.2628,
  269.5122, 268.1224, 266.863, 263.0374, 261.7913, 260.4153, 260.007, 
    263.0444, 265.5967, 266.4184, 266.9609, 268.0322, 267.7553, 267.7329, 
    267.8107,
  269.9812, 268.1494, 267.0188, 263.8255, 262.2512, 262.2841, 263.4099, 
    260.6128, 261.4851, 266.0339, 266.6802, 268.168, 268.1894, 268.2321, 
    268.6509,
  270.4505, 268.8928, 266.8939, 264.0595, 262.4679, 262.3877, 263.8171, 
    264.4136, 264.7894, 265.3387, 266.2625, 268.1756, 268.5678, 268.3942, 
    268.9014,
  271.199, 269.6164, 267.2384, 263.0949, 262.7516, 262.4362, 263.8333, 
    264.5821, 264.9261, 265.1931, 265.813, 267.9719, 268.6593, 268.5701, 
    268.8381,
  271.6617, 270.2033, 266.4531, 261.1765, 263.0423, 262.2588, 263.8208, 
    264.612, 264.6631, 264.4856, 264.8861, 267.2604, 268.5743, 268.7123, 
    268.6757,
  272.5363, 271.7195, 267.3217, 261.6104, 262.0993, 262.2122, 263.474, 
    264.7915, 264.8131, 264.399, 264.0139, 266.214, 268.4704, 268.7104, 
    268.5913,
  272.7356, 271.658, 266.7013, 262.1061, 262.5886, 261.6313, 262.1974, 
    264.6348, 264.3588, 263.4245, 263.0258, 264.7607, 268.0474, 268.7595, 
    268.3933,
  265.2803, 264.0831, 263.0896, 262.6629, 262.112, 262.4583, 263.5826, 
    264.358, 264.9958, 265.7915, 266.0846, 267.4001, 268.0428, 267.9883, 
    267.9186,
  266.9985, 265.9199, 264.4737, 263.0945, 262.5588, 263.1675, 263.1501, 
    262.2062, 262.5176, 265.2849, 265.7456, 266.7488, 268.0193, 267.5487, 
    268.0163,
  269.1438, 267.7588, 266.2945, 263.523, 262.6819, 261.2344, 262.486, 
    261.9086, 263.8803, 265.0755, 265.1229, 266.2779, 267.8407, 268.6621, 
    268.918,
  270.5224, 268.8779, 267.0069, 263.9983, 263.4203, 262.9443, 261.4389, 
    261.8184, 263.0747, 264.3666, 264.4825, 265.5628, 267.6943, 268.3115, 
    268.767,
  270.7582, 269.0787, 267.3173, 264.3121, 263.5364, 263.9124, 264.1465, 
    259.7508, 260.167, 263.7841, 264.0311, 265.3066, 267.6254, 268.2022, 
    268.8875,
  270.8372, 269.6059, 267.3043, 264.4743, 263.4109, 263.7046, 264.1927, 
    264.1122, 263.1898, 262.9971, 263.5215, 265.2693, 267.674, 268.6266, 
    269.2458,
  271.2481, 270.3913, 267.3822, 263.2822, 263.2479, 263.5699, 264.2129, 
    264.1057, 263.4774, 262.8872, 263.4389, 265.3069, 267.8694, 268.7393, 
    268.442,
  271.515, 270.9691, 267.0758, 262.7998, 262.8193, 263.1445, 264.1462, 
    264.2988, 263.4728, 262.8203, 263.0461, 265.4177, 267.8836, 267.656, 
    268.3562,
  272.261, 271.6314, 267.2055, 264.2309, 263.6306, 262.9332, 263.7138, 
    264.4189, 263.6477, 262.8362, 262.8837, 265.4344, 267.6377, 266.3963, 
    266.9467,
  272.5126, 271.4689, 268.8676, 266.4259, 266.0907, 263.3111, 262.9134, 
    264.439, 263.3988, 261.8531, 262.2105, 265.3158, 267.0414, 266.0515, 
    266.4023,
  264.8061, 265.4756, 264.6414, 264.1221, 263.7631, 263.2567, 264.0441, 
    263.4663, 261.5735, 263.1907, 263.3822, 263.4685, 264.0029, 265.5303, 
    265.9951,
  266.5345, 267.6358, 266.2935, 265.1047, 264.3024, 263.7455, 263.7461, 
    260.6002, 259.9648, 261.6433, 262.603, 263.2456, 263.1705, 264.5829, 
    265.2718,
  269.2352, 269.5196, 268.676, 266.7362, 264.7475, 262.6712, 263.0657, 
    262.735, 261.332, 263.0913, 261.8513, 263.2924, 264.2716, 265.7297, 
    266.1042,
  270.7993, 270.5316, 270.0674, 267.9461, 266.7224, 265.2244, 262.0693, 
    262.4215, 262.1928, 262.4223, 262.8962, 263.0524, 264.2077, 265.7627, 
    266.5984,
  271.2378, 271.6255, 271.1566, 269.1435, 267.4094, 266.433, 264.909, 
    260.3469, 259.674, 263.0255, 263.0721, 262.7947, 264.3605, 265.3216, 
    265.4069,
  272.5374, 272.9356, 271.6249, 269.617, 267.5495, 266.208, 265.9117, 
    265.0457, 263.8213, 263.1037, 262.9624, 263.1015, 264.485, 264.8172, 
    265.298,
  273.2593, 273.3707, 271.9189, 269.2237, 267.2522, 265.8132, 266.096, 
    266.0047, 265.0201, 263.5609, 262.8743, 262.8135, 264.8896, 265.3535, 
    265.5382,
  273.5157, 273.0692, 271.019, 268.8671, 266.8383, 265.8476, 265.8605, 
    266.8156, 265.9889, 264.2045, 262.7965, 263.3819, 265.1952, 265.9568, 
    266.7746,
  273.2531, 272.1279, 269.8866, 268.3389, 267.3261, 266.3513, 265.6864, 
    266.3604, 265.286, 263.1094, 262.2281, 263.4755, 265.3746, 266.0261, 
    266.9129,
  272.4611, 270.7448, 269.1527, 267.8567, 266.5662, 264.9881, 264.0449, 
    265.1808, 263.8997, 262.9711, 262.3955, 264.7963, 265.8506, 267.1286, 
    267.7285,
  269.6454, 267.8345, 267.2623, 266.6038, 266.5326, 266.442, 265.3779, 
    264.8064, 264.783, 264.6132, 264.6928, 263.9186, 263.2847, 263.4576, 
    264.8427,
  270.0105, 268.5634, 268.8741, 268.4236, 268.0872, 267.9496, 266.8277, 
    265.9052, 264.8251, 264.1115, 263.4809, 263.2449, 261.6479, 262.369, 
    262.8666,
  271.6122, 271.0971, 270.2807, 269.3294, 269.1606, 267.5182, 269.2447, 
    268.5854, 267.1738, 265.8633, 264.0203, 263.3455, 261.9931, 263.2735, 
    263.4147,
  272.269, 271.2776, 270.4363, 268.6843, 267.7281, 267.9289, 266.2867, 
    268.5164, 267.7842, 267.4028, 266.1852, 264.4608, 262.4069, 263.2295, 
    263.0553,
  272.2345, 270.8994, 269.5444, 267.3693, 266.0602, 265.8514, 265.7922, 
    262.9403, 262.4373, 266.8685, 266.8517, 265.3154, 262.9264, 262.784, 
    262.378,
  271.6933, 270.3688, 268.3844, 265.9177, 264.8698, 264.5045, 264.3696, 
    264.933, 264.6147, 264.7656, 265.8643, 265.6953, 263.8116, 262.3361, 
    262.6478,
  271.0724, 269.8662, 267.7407, 265.0447, 264.5876, 264.4313, 264.2206, 
    264.9052, 265.3658, 264.8632, 266.5544, 265.6705, 263.7361, 262.5539, 
    263.4391,
  270.7125, 269.5618, 267.0021, 264.9626, 264.7624, 265.2998, 265.1876, 
    265.7614, 266.1434, 266.0248, 266.3937, 265.2138, 263.7976, 263.5775, 
    264.4114,
  270.5105, 269.2036, 266.5585, 265.3998, 265.466, 266.0339, 266.3168, 
    266.1932, 265.5748, 264.8445, 265.904, 264.4629, 263.7341, 264.2507, 
    264.9168,
  270.0935, 268.4898, 266.4831, 265.8163, 265.6723, 266.2439, 266.805, 
    267.3778, 265.786, 265.5974, 265.0702, 264.6544, 264.1355, 264.5846, 
    265.5391,
  269.9046, 266.6978, 268.2378, 265.492, 264.0614, 263.0312, 264.2359, 
    265.7923, 265.1054, 264.1618, 264.739, 264.8792, 263.7548, 263.5045, 
    264.0148,
  270.8164, 268.8135, 268.8965, 267.5236, 267.166, 267.1761, 267.1452, 
    266.9604, 266.1838, 264.8227, 264.7457, 265.3227, 264.2855, 262.7329, 
    263.3652,
  272.729, 272.1113, 270.8854, 268.3351, 267.1444, 265.2502, 266.1618, 
    265.6959, 267.1254, 266.7753, 265.2386, 265.5851, 264.2644, 264.3943, 
    263.6927,
  273.2535, 272.6401, 272.0594, 269.9448, 268.0573, 267.1152, 263.8291, 
    264.3217, 263.0158, 266.8673, 266.2795, 266.4754, 265.3121, 264.8767, 
    263.8213,
  273.5939, 272.7386, 271.9034, 270.0786, 267.4197, 266.9026, 266.067, 
    261.7311, 260.107, 263.6624, 267.3619, 267.2596, 265.7059, 265.503, 
    261.0834,
  273.3826, 272.4404, 270.8283, 268.1299, 266.4326, 265.3821, 266.2054, 
    265.7245, 264.0857, 262.7895, 266.903, 268.0881, 266.4055, 263.8984, 
    262.6547,
  272.8184, 271.7584, 269.366, 267.2566, 266.0583, 266.2455, 266.8586, 
    267.039, 265.7736, 262.5353, 265.4437, 268.4954, 266.3287, 263.5026, 
    264.6078,
  272.2193, 270.9793, 268.1735, 266.8086, 267.6585, 267.5086, 267.6336, 
    267.7007, 265.8097, 264.67, 265.448, 267.9622, 265.824, 263.7193, 265.4803,
  271.441, 270.2233, 267.8178, 267.0839, 267.1025, 266.6158, 268.5679, 
    268.2663, 266.3146, 265.2671, 265.4368, 267.4792, 264.8622, 264.1492, 
    265.3791,
  270.8488, 269.4196, 267.7061, 267.6652, 267.7679, 268.4017, 268.3466, 
    268.1516, 265.9646, 265.6369, 266.3869, 266.7515, 264.058, 264.2605, 
    264.9677,
  271.5689, 269.7354, 270.237, 269.8423, 268.1876, 266.1199, 266.5737, 
    266.4023, 266.0399, 267.5527, 266.5317, 264.6372, 264.1314, 263.6348, 
    265.7381,
  271.5932, 270.1001, 269.6207, 269.8832, 269.7318, 268.9031, 267.5355, 
    267.0356, 266.4836, 267.9014, 266.9601, 265.4942, 263.621, 261.6057, 
    264.0156,
  273.6076, 272.9834, 271.7059, 271.341, 270.9135, 268.8277, 269.0418, 
    267.8751, 266.9367, 267.8023, 266.6719, 265.5999, 264.6847, 263.0883, 
    264.3445,
  273.8966, 273.262, 272.3465, 270.0983, 269.119, 270.7462, 268.1785, 
    268.0429, 265.9611, 266.9308, 266.1838, 265.2498, 265.1248, 262.8929, 
    263.6526,
  273.6273, 272.7275, 271.5563, 269.5251, 266.9332, 267.6416, 266.7797, 
    265.1233, 262.6024, 265.4738, 266.4152, 265.1737, 264.455, 263.572, 
    262.684,
  272.9888, 272.2679, 271.0871, 269.463, 267.2051, 262.8131, 266.2378, 
    267.5578, 265.9383, 265.2844, 266.4847, 265.5394, 265.328, 263.0169, 
    263.0406,
  272.4638, 271.6803, 269.7851, 268.418, 267.4333, 263.317, 265.7585, 
    266.5424, 265.887, 265.1729, 266.3185, 265.4869, 265.1624, 263.2511, 
    266.0626,
  271.7378, 270.7314, 268.5529, 267.3296, 268.0981, 265.9528, 264.8277, 
    266.7809, 265.188, 265.4871, 266.2231, 265.5963, 264.586, 264.5316, 
    267.468,
  271.0748, 270.0233, 267.5017, 267.8969, 267.7413, 266.5483, 267.0359, 
    266.8867, 265.8375, 265.5935, 265.3205, 265.4035, 264.1615, 266.428, 
    267.2083,
  270.3352, 269.0535, 267.1094, 267.7905, 267.3067, 267.2509, 267.2236, 
    267.0944, 265.8342, 265.6057, 265.4542, 265.7162, 264.1602, 266.2573, 
    267.1163,
  272.6696, 268.8828, 268.6113, 269.1607, 269.5894, 268.593, 267.2669, 
    267.9061, 267.7377, 268.5689, 266.1571, 263.9958, 266.0862, 267.3134, 
    268.9189,
  271.8807, 270.4847, 269.3602, 270.4847, 270.6766, 268.8892, 268.1025, 
    267.8108, 266.2286, 266.1396, 267.5218, 264.5067, 265.9464, 266.2096, 
    268.4455,
  273.9823, 273.3867, 272.0166, 270.3533, 269.6935, 267.9912, 268.4344, 
    267.907, 266.4005, 267.4522, 266.7534, 264.9308, 266.0973, 266.4127, 
    268.2943,
  273.7611, 273.1231, 272.5692, 270.1944, 268.7678, 269.1521, 267.7619, 
    268.5881, 266.2324, 267.7326, 266.3176, 264.8063, 265.1317, 265.803, 
    267.6233,
  273.4034, 272.6768, 271.986, 270.074, 267.7965, 268.6838, 269.9597, 
    266.1708, 264.957, 266.9743, 266.2796, 266.0004, 265.291, 265.4701, 
    267.0977,
  272.5523, 272.0593, 270.8269, 269.3528, 267.2846, 265.1666, 268.072, 
    270.0434, 268.0474, 266.9167, 267.0379, 266.1096, 265.6944, 264.9442, 
    267.2097,
  272.0063, 271.284, 269.1336, 268.4101, 267.3603, 265.5924, 266.4204, 
    268.9118, 268.111, 266.6546, 267.0736, 266.1095, 266.1415, 265.8692, 
    267.7506,
  271.2574, 270.4019, 268.4327, 266.0053, 267.8046, 265.6118, 264.6769, 
    267.7999, 267.072, 265.9823, 266.3904, 265.6933, 265.0956, 266.1999, 
    268.0728,
  270.6664, 269.6646, 267.1385, 266.6569, 266.4922, 265.3384, 266.8046, 
    267.8632, 267.1272, 265.646, 266.0721, 265.1872, 264.5906, 266.8737, 
    267.9115,
  269.9839, 268.7881, 267.1522, 267.0207, 266.432, 266.8224, 267.5262, 
    267.738, 266.312, 265.4377, 265.4895, 265.2577, 264.6065, 267.0121, 
    267.4456,
  273.4251, 269.3577, 268.5622, 268.3617, 269.5255, 269.7434, 270.0497, 
    270.6273, 270.66, 270.2114, 268.6886, 267.1641, 266.8342, 266.6605, 
    268.3476,
  271.9102, 270.7154, 269.4194, 269.4139, 271.8332, 271.4596, 271.0842, 
    270.6354, 269.748, 268.5124, 268.6539, 266.9192, 266.5127, 266.6829, 
    269.2851,
  274.4603, 273.678, 272.5824, 269.2037, 271.3493, 268.5603, 269.6673, 
    268.3632, 269.0868, 268.0064, 267.3261, 266.2713, 266.3455, 267.8387, 
    270.6947,
  274.2629, 273.5654, 273.0313, 271.1833, 268.2957, 269.0764, 268.5078, 
    266.3878, 267.2364, 265.5678, 264.0538, 264.3332, 267.0526, 269.2993, 
    271.3074,
  273.6117, 272.9773, 272.2618, 270.5266, 269.5443, 269.7633, 270.0232, 
    264.7856, 262.9286, 266.9792, 265.3468, 266.7589, 268.5748, 270.1903, 
    270.7219,
  272.9937, 272.3392, 271.1874, 268.5595, 268.1866, 267.934, 268.4531, 
    267.0044, 266.6077, 266.1118, 267.1635, 268.1231, 269.5863, 270.3314, 
    270.2971,
  272.2468, 271.4457, 269.4442, 267.6734, 267.0234, 267.5898, 269.5766, 
    267.3973, 266.6335, 266.8629, 268.3245, 269.215, 269.6617, 269.9603, 
    269.5096,
  271.4191, 270.4995, 268.6151, 264.8893, 267.957, 267.0648, 268.8093, 
    268.1077, 266.7295, 267.3543, 268.5924, 269.1814, 269.2769, 269.0814, 
    268.8557,
  270.779, 269.7607, 267.2341, 267.2943, 267.9528, 267.4621, 268.6052, 
    267.7454, 266.7924, 266.9086, 268.121, 268.6729, 268.7118, 268.694, 
    268.4137,
  269.9867, 268.8384, 266.9693, 267.4666, 268.0558, 268.2604, 268.1895, 
    267.4117, 266.7111, 266.9966, 267.4799, 267.9586, 268.177, 268.091, 
    268.0591,
  272.7402, 270.514, 269.5293, 270.5396, 269.1861, 269.9055, 271.0406, 
    271.2702, 270.6507, 270.2557, 269.9507, 270.4825, 270.2042, 269.3719, 
    268.3847,
  271.7215, 269.914, 269.615, 269.3191, 270.7127, 271.5639, 271.6309, 
    271.2885, 270.4923, 270.4923, 269.721, 270.7465, 270.541, 268.8558, 
    268.4732,
  273.9233, 273.5615, 272.5242, 269.6158, 270.3498, 268.0483, 268.8651, 
    268.9881, 269.2746, 269.067, 269.2818, 270.3898, 269.4356, 268.0442, 
    267.4951,
  274.5492, 273.9636, 273.2105, 270.9964, 266.6612, 267.3484, 266.4435, 
    266.4435, 268.0956, 269.1635, 268.553, 268.2017, 267.1803, 267.0779, 
    267.6497,
  274.5682, 273.5345, 272.8056, 269.8252, 265.3307, 268.7379, 268.4347, 
    265.0039, 263.9424, 266.0427, 267.3051, 266.6239, 266.4421, 266.6754, 
    269.0672,
  273.7121, 272.8273, 271.442, 268.1852, 266.6494, 267.4126, 267.7333, 
    266.4947, 267.463, 265.0102, 265.3267, 266.5457, 267.1579, 269.0564, 
    269.5818,
  272.8674, 272.0409, 269.6378, 267.7454, 267.2464, 267.5143, 267.9506, 
    265.6509, 267.4636, 267.9281, 268.1658, 268.9747, 269.5135, 269.9409, 
    269.359,
  271.9616, 270.7874, 268.7626, 266.8362, 267.8181, 267.8896, 267.1927, 
    266.6537, 266.7614, 268.6746, 269.4646, 269.7105, 269.7682, 268.9854, 
    268.4061,
  271.1838, 269.935, 267.7062, 268.4073, 268.4509, 268.1072, 267.8643, 
    267.7896, 268.3455, 269.7695, 269.8489, 268.9801, 268.6355, 268.4017, 
    268.7213,
  270.4274, 269.3326, 267.9573, 267.962, 267.8315, 268.0091, 267.9895, 
    268.5251, 269.5028, 269.355, 268.998, 268.3813, 268.3676, 268.7727, 
    269.4207,
  275.2118, 272.1864, 270.7191, 269.7921, 269.7228, 270.1821, 269.6276, 
    269.1941, 268.3598, 268.7984, 270.27, 268.8913, 268.3119, 268.6052, 
    269.0904,
  272.5911, 271.0924, 270.5065, 270.1434, 269.6526, 270.9094, 269.8196, 
    268.9971, 268.1697, 268.5267, 269.6979, 269.4513, 268.1458, 268.7806, 
    267.4384,
  273.4501, 273.1699, 272.3345, 271.2816, 270.2266, 267.2368, 267.7602, 
    267.3446, 266.8782, 267.3441, 267.7274, 269.188, 268.6455, 267.611, 
    268.3508,
  273.9812, 273.5669, 273.1138, 271.9825, 268.8228, 268.6985, 264.3361, 
    265.0858, 265.0194, 267.9028, 269.3241, 269.2812, 269.3918, 268.9599, 
    269.013,
  274.4314, 273.7784, 273.4613, 271.4709, 267.0288, 267.1842, 266.5539, 
    264.0487, 262.2774, 266.8883, 268.6223, 269.1718, 269.8322, 268.0793, 
    268.0368,
  274.5956, 273.8564, 272.9486, 269.8749, 266.6622, 266.8625, 267.2624, 
    266.5046, 265.9846, 265.1366, 265.3577, 265.988, 267.5238, 268.6197, 
    269.2456,
  273.8293, 273.2793, 271.2926, 267.7977, 266.7716, 267.2182, 266.9968, 
    266.5907, 267.9277, 266.6483, 268.1631, 268.4864, 268.6731, 268.6917, 
    269.2352,
  272.9549, 272.3774, 269.144, 266.5467, 267.301, 267.3172, 266.2488, 
    266.7416, 264.8504, 265.5111, 266.9312, 268.3622, 268.8867, 268.9322, 
    268.86,
  271.9659, 271.5052, 268.0092, 267.5866, 268.3725, 266.2971, 265.7679, 
    265.4064, 267.0943, 267.7233, 265.9781, 267.7488, 269.0013, 269.0076, 
    269.0029,
  271.6692, 270.5404, 268.0835, 268.4977, 267.2979, 267.7321, 266.9811, 
    267.2314, 268.3269, 268.6145, 267.1061, 268.8941, 269.0366, 269.0442, 
    269.2634,
  280.0402, 277.2003, 275.0967, 274.8147, 274.2323, 273.5737, 272.8249, 
    272.1029, 271.2138, 270.5428, 270.4804, 269.8748, 269.6414, 269.6265, 
    269.7353,
  275.5172, 275.2701, 274.6891, 274.24, 274.2786, 273.0193, 272.3849, 
    271.6774, 270.8214, 269.6765, 269.6133, 268.9418, 268.1967, 269.0067, 
    268.4432,
  275.4808, 274.9286, 274.4454, 273.8323, 273.0527, 271.3433, 270.4696, 
    269.8883, 269.1962, 268.1196, 267.8227, 267.7603, 267.586, 267.3789, 
    268.7702,
  275.5625, 275.0135, 274.0491, 272.9577, 272.1241, 270.9931, 266.8963, 
    267.6273, 267.3722, 267.0803, 267.3948, 266.9204, 268.8213, 269.487, 
    268.0492,
  275.0649, 273.6199, 272.7327, 271.1618, 269.6246, 268.6659, 268.2319, 
    265.1888, 263.5461, 266.7873, 266.8665, 267.537, 268.351, 269.1431, 
    269.4193,
  272.9725, 272.2007, 271.1251, 269.5438, 268.0792, 267.2639, 266.7958, 
    267.1134, 266.6425, 265.6415, 265.6073, 265.5782, 268.2159, 269.004, 
    269.3116,
  272.8439, 272.1262, 270.3004, 267.7239, 266.8892, 266.5259, 266.0528, 
    266.0357, 267.0698, 267.4646, 268.1759, 267.6997, 268.5515, 269.0051, 
    269.322,
  272.7734, 271.687, 268.9134, 266.8595, 266.4408, 267.7152, 266.312, 
    266.9831, 266.5317, 267.243, 267.4211, 267.6343, 268.393, 269.5164, 
    269.5497,
  272.2003, 270.9473, 268.2585, 267.4473, 268.4472, 266.6414, 266.5497, 
    266.9858, 267.4607, 267.8029, 267.2192, 268.6794, 269.1733, 269.3723, 
    268.925,
  271.5306, 270.1452, 268.736, 268.6885, 267.3437, 267.4477, 267.1837, 
    267.2178, 267.4236, 268.2315, 267.2631, 268.5026, 268.8191, 268.7031, 
    268.4695,
  275.9587, 273.5919, 272.7467, 272.7362, 272.8138, 272.9278, 272.8337, 
    272.9706, 273.0632, 272.9836, 273.2405, 273.3774, 273.4384, 272.8276, 
    272.3005,
  273.3796, 272.7853, 272.4806, 272.433, 272.7166, 272.9152, 272.9522, 
    272.9432, 272.9781, 273.1159, 273.2565, 273.336, 273.0822, 272.0286, 
    271.5457,
  273.6729, 272.8823, 272.3192, 272.1476, 272.4626, 271.972, 272.568, 
    271.1447, 271.2781, 271.6763, 272.0818, 272.2928, 272.0559, 271.8025, 
    271.3607,
  273.1214, 272.2659, 271.8955, 271.5768, 271.6251, 271.7421, 268.1421, 
    269.3972, 269.5872, 269.9413, 270.2987, 270.6245, 270.8403, 270.5827, 
    270.3566,
  272.5788, 271.4202, 270.8946, 269.6038, 269.1443, 269.1154, 269.3033, 
    265.873, 264.8008, 268.7809, 269.0734, 269.3385, 269.6568, 269.8304, 
    270.0028,
  271.8062, 270.711, 269.7415, 268.0901, 267.4082, 267.0736, 267.0107, 
    267.6274, 268.0391, 268.3814, 268.4327, 268.5534, 268.8871, 269.1351, 
    269.179,
  271.5255, 270.3925, 268.8878, 267.1555, 266.7121, 266.3105, 266.1116, 
    266.2967, 266.9652, 268.0855, 268.3238, 268.2574, 268.4349, 268.5183, 
    268.386,
  270.8976, 269.8065, 268.1708, 267.3819, 266.8972, 266.9644, 266.5094, 
    266.3461, 266.3525, 266.9554, 267.6428, 267.8009, 268.1337, 268.3352, 
    268.1662,
  270.8748, 268.9648, 267.429, 267.3307, 267.3156, 267.4796, 266.9762, 
    267.2802, 267.3765, 267.1908, 267.3016, 267.6563, 267.8508, 267.8849, 
    268.9026,
  270.6447, 268.5718, 267.3926, 267.1156, 266.8977, 267.0359, 267.4662, 
    267.0186, 267.3417, 267.5358, 267.5009, 267.92, 268.0344, 268.3172, 
    268.8532,
  276.5476, 273.2044, 271.6925, 270.2451, 270.7134, 271.1063, 270.8304, 
    268.0519, 267.66, 268.2576, 269.5669, 270.2439, 270.754, 271.1121, 271.8,
  273.6931, 272.0811, 271.1425, 269.4948, 270.0832, 270.8315, 270.4029, 
    267.2578, 267.14, 267.6479, 268.7426, 270.0707, 270.5579, 270.8192, 
    271.9957,
  273.6572, 272.2238, 270.7823, 269.0594, 268.672, 268.2411, 269.9831, 
    266.6438, 266.5456, 267.0929, 267.6846, 269.0863, 270.4114, 271.6166, 
    272.5111,
  273.4778, 271.8422, 270.5208, 268.7752, 267.4282, 268.3853, 266.4569, 
    266.1418, 266.658, 267.2783, 267.2907, 268.4457, 270.2558, 271.7296, 
    272.5163,
  272.5284, 270.9244, 270.1253, 267.9313, 266.5457, 265.8649, 268.6686, 
    265.006, 264.5886, 267.4567, 267.2185, 267.8929, 269.9303, 271.6648, 
    272.5439,
  271.9085, 270.6039, 269.4868, 266.8635, 265.6293, 265.205, 268.1283, 
    268.1402, 267.7222, 267.3707, 266.6845, 268.0095, 269.4237, 270.6305, 
    271.7978,
  271.7209, 270.2449, 268.9129, 267.1866, 265.6109, 265.6119, 264.7269, 
    266.9818, 266.9804, 266.5031, 266.1662, 268.0417, 269.2332, 269.8984, 
    270.6642,
  271.6362, 270.3033, 268.1445, 267.3492, 266.7625, 266.7636, 265.3266, 
    265.3557, 266.4026, 265.3224, 266.3975, 268.2732, 269.3704, 269.802, 
    270.3517,
  271.9429, 269.8936, 267.4617, 267.2766, 267.2401, 267.4052, 266.1136, 
    265.7502, 265.4844, 265.4395, 266.2801, 268.5332, 269.6233, 270.1266, 
    270.4372,
  271.4802, 268.502, 267.7916, 268.0237, 268.0129, 266.5337, 266.937, 
    266.2082, 265.6012, 265.9572, 267.0934, 268.9267, 269.8802, 270.3801, 
    270.5771,
  273.6983, 272.2947, 271.858, 271.9996, 271.9482, 271.9229, 271.9415, 
    270.9763, 270.0172, 269.4996, 268.8998, 268.1833, 267.5038, 266.4113, 
    265.9363,
  272.3809, 271.8115, 271.9564, 271.6909, 271.9093, 271.7596, 271.501, 
    269.888, 268.8971, 268.4059, 268.3986, 267.6081, 265.8289, 264.8598, 
    265.5648,
  272.8058, 272.1594, 271.8546, 271.2721, 271.4337, 269.6143, 269.8039, 
    268.4256, 267.7608, 267.1959, 267.1175, 266.5667, 265.2231, 265.5928, 
    267.7617,
  272.6968, 271.7879, 271.2313, 270.3976, 269.9405, 269.6031, 266.282, 
    267.5169, 267.0767, 266.7151, 266.0085, 264.8053, 264.8979, 267.8376, 
    269.6853,
  272.3228, 270.7555, 269.9631, 268.6033, 268.5538, 268.501, 268.9274, 
    264.7715, 263.7539, 266.1912, 265.0871, 264.3249, 266.9731, 269.8371, 
    271.8254,
  272.2119, 270.2915, 268.7809, 267.4816, 267.3118, 267.4998, 268.1298, 
    268.0645, 266.9942, 266.7089, 266.4716, 266.6935, 269.396, 271.2858, 
    272.6407,
  272.2682, 270.1236, 268.0782, 266.9543, 266.9537, 267.1466, 266.6776, 
    266.7025, 266.7718, 266.7098, 265.3607, 268.7117, 270.5766, 271.6496, 
    272.6844,
  272.4914, 270.341, 267.5758, 267.36, 267.1719, 266.9023, 265.7717, 
    264.7001, 266.3231, 265.0329, 266.9535, 270.1161, 270.8008, 270.8788, 
    271.5188,
  272.7125, 270.654, 268.4756, 268.5087, 268.5793, 268.184, 267.4439, 
    264.164, 264.6031, 266.3106, 269.0212, 270.6893, 270.3486, 270.6585, 
    270.9207,
  272.4477, 270.7805, 269.7414, 269.1742, 269.332, 263.992, 264.1103, 
    264.7766, 264.8763, 267.8113, 269.7072, 270.4489, 269.9752, 270.053, 
    270.1526,
  277.5872, 274.2613, 272.4552, 269.252, 267.9254, 268.4004, 268.411, 
    269.1088, 270.2982, 271.1206, 271.2543, 270.1327, 269.6694, 269.3226, 
    269.3582,
  274.2061, 273.1342, 271.5886, 268.5089, 267.1692, 268.0865, 268.0876, 
    268.325, 269.2679, 269.7346, 269.6052, 269.1624, 269.0387, 267.8835, 
    267.965,
  274.6586, 273.3814, 271.5416, 267.8807, 266.3428, 266.4754, 267.8036, 
    267.7099, 267.979, 268.3601, 268.222, 267.9135, 267.4249, 267.3037, 
    268.1292,
  274.9908, 273.5862, 271.3262, 267.8134, 266.3063, 267.7468, 266.1543, 
    267.6304, 267.6187, 267.9939, 268.3241, 267.8659, 267.3106, 267.6906, 
    269.3372,
  275.1789, 273.2426, 271.1838, 267.3418, 266.5167, 267.8868, 267.9415, 
    264.1848, 263.7028, 268.2592, 268.7137, 269.1788, 270.1617, 271.1969, 
    271.9055,
  275.4407, 273.596, 271.166, 268.6569, 268.0242, 267.6169, 267.3503, 
    267.5756, 267.6479, 268.8751, 269.583, 270.4965, 271.7336, 272.3635, 
    272.4745,
  275.2947, 274.6275, 271.9599, 269.6848, 268.9377, 268.4061, 267.8221, 
    267.5016, 268.013, 269.1588, 270.1739, 271.2645, 272.133, 272.593, 
    272.8111,
  275.1897, 274.7262, 272.4932, 270.9569, 270.0518, 269.4008, 268.3783, 
    267.3198, 267.8792, 268.6097, 270.5168, 271.4197, 272.0411, 272.4451, 
    272.4035,
  274.711, 273.7362, 271.3799, 270.9081, 270.7574, 270.0315, 268.9181, 
    265.8608, 267.3816, 269.844, 270.5457, 270.9109, 271.1971, 271.3595, 
    271.3378,
  273.6414, 272.2924, 270.84, 269.8458, 270.2794, 269.381, 266.7941, 
    265.8921, 268.378, 270.0477, 269.8717, 269.9597, 270.1724, 270.5842, 
    270.5403,
  279.8343, 275.4482, 274.6396, 271.8266, 267.8536, 265.313, 263.4963, 
    265.5847, 269.0209, 270.5768, 271.5157, 271.6549, 271.391, 271.3077, 
    271.3838,
  275.1562, 273.7782, 272.8214, 270.1333, 267.6492, 265.2805, 263.6075, 
    265.7285, 267.914, 270.7264, 271.6964, 271.7785, 271.2396, 270.623, 
    271.3967,
  274.6138, 273.5538, 271.9644, 269.0963, 266.7821, 264.3517, 264.8807, 
    265.9292, 267.7248, 270.4026, 271.5222, 272.1389, 271.889, 271.7731, 
    272.0302,
  275.0117, 274.1287, 272.0797, 269.4409, 265.2964, 266.3736, 264.9438, 
    266.3217, 267.7676, 269.7601, 271.236, 272.2328, 272.2746, 272.1776, 
    271.9838,
  275.1479, 273.8185, 272.6351, 269.3044, 267.0779, 268.1563, 268.0981, 
    264.4371, 264.3386, 269.3712, 270.8629, 271.9957, 272.115, 271.7482, 
    271.6303,
  275.3317, 274.6096, 273.1461, 270.5906, 269.3265, 268.899, 268.8304, 
    268.676, 267.8006, 269.4946, 270.7724, 271.7724, 271.7427, 271.2435, 
    271.1154,
  274.8382, 274.3059, 272.7077, 271.8646, 270.799, 270.029, 269.6785, 
    269.1594, 267.607, 269.4844, 270.284, 271.3213, 271.2714, 270.8596, 
    270.6479,
  274.7903, 273.1557, 270.5624, 270.4276, 270.8073, 271.4139, 270.7121, 
    268.7139, 268.6885, 269.2099, 270.0669, 270.7895, 270.8322, 270.3927, 
    270.5195,
  273.0054, 271.635, 269.467, 268.9507, 271.1803, 271.1663, 270.0417, 
    267.2456, 268.8401, 269.0531, 269.9835, 270.5151, 270.5727, 270.356, 
    270.7235,
  272.0116, 270.4119, 269.5166, 268.9453, 268.4944, 270.4991, 268.9889, 
    266.7811, 268.944, 269.0128, 270.0414, 270.4258, 270.5861, 270.5961, 
    270.8645,
  275.8378, 272.3088, 271.1889, 268.7533, 267.0041, 265.6931, 264.1387, 
    264.153, 266.1978, 269.3612, 270.7805, 271.4871, 271.555, 271.4184, 
    270.9453,
  272.8766, 271.4842, 270.4701, 268.6778, 267.8814, 266.0775, 264.9366, 
    265.3042, 265.1385, 269.2418, 270.3854, 271.1488, 271.5063, 270.1661, 
    270.0449,
  273.0088, 271.9213, 271.0486, 269.1679, 268.2677, 265.7884, 266.9023, 
    268.228, 266.3586, 269.1194, 270.1594, 271.0498, 271.4407, 270.9403, 
    270.5846,
  273.2751, 272.21, 271.2964, 269.502, 266.9423, 268.126, 266.8046, 267.9963, 
    267.4901, 269.1195, 270.1189, 270.9527, 271.443, 271.3476, 271.0476,
  273.2458, 272.4657, 272.2006, 270.0675, 267.4996, 269.273, 269.4597, 
    265.7575, 264.906, 269.0338, 270.1648, 271.0187, 271.6414, 271.6006, 
    271.707,
  273.5725, 272.9067, 271.824, 271.188, 270.7832, 270.035, 268.817, 269.0858, 
    268.4768, 269.3622, 270.5119, 271.174, 271.8076, 271.9485, 272.1683,
  273.0944, 272.0687, 270.7116, 269.7244, 269.6465, 269.7813, 269.5174, 
    269.3298, 268.7358, 269.5946, 270.2457, 271.0516, 271.903, 272.1396, 
    272.4336,
  272.672, 271.3201, 269.8926, 269.5317, 269.343, 269.0322, 268.7763, 
    268.8911, 269.8405, 269.629, 270.689, 271.3824, 272.0448, 272.2903, 
    272.478,
  272.5063, 271.2676, 270.0242, 269.531, 268.9231, 268.5896, 268.4808, 
    269.0277, 269.8349, 270.0075, 270.7353, 271.5065, 272.2376, 272.2973, 
    272.3428,
  271.7274, 270.6314, 269.8952, 269.2407, 268.5342, 268.1548, 268.529, 
    269.3203, 269.6594, 270.0731, 270.7322, 271.7134, 272.376, 272.5013, 
    272.3604,
  272.8294, 270.2275, 269.2878, 268.1797, 268.3636, 267.3535, 266.7813, 
    267.2499, 268.4209, 269.8505, 270.7703, 271.7602, 272.0515, 271.9413, 
    272.0174,
  271.5712, 270.4889, 270.038, 269.1633, 269.1231, 268.9544, 268.3677, 
    268.874, 268.4186, 269.9802, 270.8802, 271.7942, 271.9715, 271.2938, 
    271.6445,
  272.1749, 271.2954, 270.3184, 268.9735, 268.1179, 266.6975, 269.3437, 
    269.5958, 269.5907, 270.1091, 270.7572, 271.5535, 271.9255, 271.878, 
    271.9284,
  272.7537, 271.5759, 270.1638, 269.2231, 268.4088, 268.6796, 266.9083, 
    268.6386, 269.549, 270.1541, 270.4615, 271.3251, 271.5626, 271.8336, 
    271.925,
  273.1848, 271.7441, 270.8043, 268.5632, 268.6254, 268.8029, 269.1145, 
    265.7087, 265.5729, 270.0956, 270.6256, 271.1033, 271.6739, 271.8731, 
    271.9713,
  273.1802, 271.6317, 269.9071, 268.5431, 268.5854, 268.9708, 269.1656, 
    269.0451, 269.2713, 270.0237, 270.9827, 271.2091, 271.7696, 271.9394, 
    272.1855,
  272.7726, 270.9354, 268.8112, 268.3292, 268.7503, 268.9783, 269.0654, 
    269.1713, 269.6071, 270.3237, 270.6333, 271.3969, 272.0387, 272.157, 
    272.2941,
  272.3357, 270.5997, 268.7921, 268.5757, 269.0623, 268.8734, 268.7791, 
    268.8689, 269.6349, 270.15, 270.6508, 271.5839, 272.0828, 272.1699, 
    272.2887,
  271.9027, 270.3448, 268.9868, 268.6736, 268.9953, 268.6543, 268.4269, 
    268.7661, 269.5775, 270.1137, 270.4117, 271.5294, 272.0802, 272.2133, 
    272.2284,
  271.3935, 270.0349, 269.6419, 268.8706, 268.8831, 268.4891, 268.2664, 
    268.5979, 269.4203, 269.8472, 270.4108, 271.4882, 272.0299, 272.3214, 
    272.3214,
  272.2301, 269.6943, 268.9328, 268.7048, 268.8351, 269.04, 268.8435, 
    269.1224, 269.5342, 269.854, 270.2108, 270.485, 270.809, 271.1988, 
    271.5752,
  270.5929, 269.5937, 269.2421, 269.0379, 269.0931, 269.3648, 269.1862, 
    269.2721, 269.6954, 270.0487, 270.2941, 270.5716, 270.8635, 270.5786, 
    271.4152,
  271.175, 270.1408, 269.7846, 269.1906, 268.8786, 266.9398, 268.9979, 
    269.4221, 269.6148, 269.9942, 270.1657, 270.7957, 271.3973, 271.6651, 
    271.9148,
  271.446, 270.4884, 270.027, 269.3596, 268.9205, 268.7929, 266.5722, 
    268.8098, 269.5621, 270.0728, 270.1073, 271.3151, 271.9201, 272.068, 
    272.3893,
  271.5995, 271.0596, 270.1721, 268.9259, 269.0693, 268.5567, 268.3737, 
    264.9239, 265.3001, 269.8087, 270.3904, 271.8252, 272.2955, 272.3079, 
    272.4082,
  271.9703, 271.0526, 269.6387, 268.8943, 268.9557, 268.4023, 268.1836, 
    268.2664, 268.9088, 269.4381, 271.0957, 272.4005, 272.6417, 272.3176, 
    272.1911,
  271.9507, 271.2905, 269.6948, 268.8097, 268.8843, 268.3991, 268.1606, 
    268.6462, 269.4413, 270.1825, 271.6595, 272.655, 272.5598, 272.2931, 
    272.096,
  271.8858, 271.4215, 269.7766, 269.1094, 268.8291, 268.3828, 268.4265, 
    269.0425, 269.8573, 270.6877, 271.9677, 272.6154, 272.5271, 272.2317, 
    271.8551,
  271.7946, 271.3845, 270.4444, 269.486, 268.8836, 268.5216, 268.7571, 
    269.5148, 270.1213, 271.0832, 272.1214, 272.5733, 272.4895, 272.2227, 
    271.834,
  271.7378, 271.5064, 271.2202, 269.8526, 269.1551, 268.7364, 269.0484, 
    269.8581, 270.6236, 271.6608, 272.3655, 272.5416, 272.4982, 272.3557, 
    271.8039,
  271.7108, 269.7189, 269.9846, 269.6474, 268.9859, 269.3711, 269.0564, 
    269.3357, 269.5747, 270.0405, 270.4775, 271.2704, 271.9066, 272.2535, 
    272.4711,
  270.1827, 270.4955, 270.4931, 269.9034, 269.6896, 269.5263, 269.416, 
    268.9555, 269.1141, 269.8922, 270.3975, 271.2082, 271.652, 271.4191, 
    272.2271,
  270.9186, 270.7484, 271.1062, 270.4334, 269.7366, 267.4945, 269.6169, 
    269.6681, 269.667, 269.8917, 270.3291, 270.8456, 271.3971, 271.7182, 
    272.1478,
  271.2402, 271.5432, 271.803, 270.8949, 269.9237, 269.4608, 267.4171, 
    270.0171, 270.3891, 270.239, 270.2249, 270.5774, 271.2807, 271.6938, 
    271.9766,
  271.2868, 272.3344, 272.2759, 271.0123, 270.1693, 270.071, 269.9167, 
    266.6778, 266.614, 270.7941, 270.5274, 270.3851, 271.0982, 271.5867, 
    272.0128,
  272.6797, 272.9781, 272.378, 271.1785, 270.5341, 270.4858, 270.6556, 
    270.5436, 270.4604, 270.4547, 270.5317, 270.6236, 271.0373, 271.5368, 
    271.9703,
  273.3421, 273.3947, 272.3164, 271.1631, 270.8894, 271.1505, 271.162, 
    271.21, 271.007, 271.0086, 271.0636, 271.0766, 271.2587, 271.6846, 
    271.9783,
  273.6135, 273.3474, 271.89, 271.2877, 271.1523, 271.5228, 271.4826, 
    271.401, 271.2524, 271.2861, 271.3914, 271.6037, 271.6281, 271.7493, 
    272.0109,
  273.6997, 272.993, 271.7625, 271.702, 271.4536, 271.777, 271.6414, 
    271.6232, 271.5188, 271.5894, 272.0458, 272.2953, 271.4474, 271.5839, 
    272.0724,
  273.6961, 272.8182, 271.9881, 271.782, 271.4556, 271.8744, 271.8593, 
    271.801, 271.8409, 272.0802, 272.4048, 272.4718, 272.4008, 272.1924, 
    272.2148,
  273.5461, 270.1051, 269.9682, 270.8123, 271.1071, 271.3067, 271.1884, 
    271.3279, 271.2601, 271.2623, 271.3016, 270.9456, 271.3774, 271.5002, 
    271.9263,
  270.6718, 269.8221, 271.0661, 271.411, 271.5458, 271.6028, 271.6874, 
    271.6909, 271.7256, 271.741, 271.8695, 271.3797, 271.0677, 270.5649, 
    271.6455,
  270.5819, 271.2152, 272.3585, 271.8779, 271.563, 269.6197, 271.9521, 
    272.0785, 272.3549, 272.1082, 271.8344, 271.6274, 271.125, 271.2748, 
    271.8206,
  271.6083, 272.625, 272.7171, 271.9635, 271.499, 271.6434, 270.0677, 
    272.0979, 272.7216, 272.5597, 272.0851, 271.8667, 271.3917, 271.1122, 
    271.5138,
  272.3788, 273.2607, 272.5576, 271.6829, 271.6939, 272.0454, 271.974, 
    269.2354, 269.1255, 272.6789, 272.4612, 272.0214, 271.5219, 271.0462, 
    271.2179,
  273.5916, 273.3783, 271.9952, 271.6856, 271.9023, 272.3021, 272.38, 
    272.3303, 272.4709, 272.5938, 272.6412, 272.1234, 271.7699, 271.1834, 
    271.2148,
  273.8044, 272.9858, 271.5952, 271.9065, 272.1346, 272.3922, 272.3671, 
    272.3348, 272.41, 272.483, 272.6539, 272.1037, 271.846, 271.1471, 271.1354,
  273.6789, 272.6642, 271.663, 272.0988, 272.2294, 272.3643, 272.3282, 
    272.2524, 272.3152, 272.5025, 272.6702, 272.5651, 272.0219, 271.1621, 
    271.1328,
  273.7664, 272.6096, 272.0633, 272.3286, 272.394, 272.4627, 272.367, 
    272.1689, 272.0675, 272.2381, 272.4825, 272.6499, 271.6018, 271.0832, 
    271.2251,
  273.1058, 272.1358, 272.3607, 272.4055, 272.4684, 272.486, 272.5253, 
    272.2251, 272.1699, 272.4558, 272.6617, 272.6369, 271.8851, 271.0074, 
    271.3845,
  273.0215, 270.8621, 271.009, 271.567, 271.57, 271.8269, 271.7128, 271.7213, 
    271.6081, 271.8907, 272.3903, 272.0025, 271.9135, 270.2545, 271.2593,
  271.0188, 271.5227, 271.8443, 271.4407, 271.7837, 272.1086, 272.0366, 
    271.7431, 271.5477, 271.9312, 271.9557, 271.4522, 272.0152, 271.4984, 
    271.4131,
  272.3925, 272.8564, 272.3359, 271.9403, 271.9471, 270.3045, 272.2287, 
    271.6804, 271.4815, 271.9025, 271.5581, 272.2926, 272.1256, 272.3838, 
    272.4342,
  273.0706, 273.1244, 272.4971, 272.0921, 272.1223, 272.1626, 270.5096, 
    271.7675, 271.2876, 271.9385, 272.0403, 272.3975, 271.9045, 271.6871, 
    271.6207,
  273.4665, 273.1162, 272.5255, 272.0376, 272.3571, 272.599, 272.4369, 
    269.2685, 268.7523, 271.9836, 272.5361, 272.3737, 271.9275, 271.3343, 
    270.779,
  273.3415, 273.1873, 272.3721, 272.1764, 272.5322, 272.727, 272.7503, 
    272.5274, 272.273, 272.6123, 272.7814, 272.2219, 271.826, 271.5788, 
    271.0932,
  273.25, 273.1357, 272.4248, 272.3924, 272.6148, 272.7606, 272.6006, 
    272.0317, 272.3094, 272.6821, 272.5705, 272.2209, 272.0068, 271.8712, 
    271.2849,
  273.3386, 273.1375, 272.3681, 272.495, 272.5717, 272.6814, 272.754, 
    272.7389, 272.7284, 272.7306, 272.6108, 272.2458, 271.9441, 271.9415, 
    271.739,
  273.2618, 272.9454, 272.3437, 272.6059, 272.6196, 272.5667, 272.5534, 
    272.4588, 272.5085, 272.532, 272.5582, 272.1734, 271.9325, 271.8755, 
    272.176,
  272.7982, 272.7402, 272.4507, 272.5623, 272.6719, 272.7025, 272.6356, 
    272.3501, 272.5258, 272.8094, 272.6323, 272.138, 271.8414, 271.9124, 
    272.3054,
  272.8405, 271.5182, 271.7273, 271.933, 271.677, 271.4772, 271.9707, 
    272.033, 271.251, 271.5028, 271.8116, 271.7142, 271.6758, 270.3506, 
    272.1483,
  271.879, 272.3862, 272.33, 271.8517, 272.108, 272.555, 272.438, 272.3173, 
    271.967, 271.6907, 271.6816, 271.3967, 269.5108, 271.3839, 272.0664,
  272.7101, 273.1784, 272.5871, 272.184, 271.8453, 271.5291, 272.4835, 
    272.3725, 272.0077, 271.813, 271.38, 271.5322, 269.136, 271.2399, 272.3629,
  273.4685, 273.1252, 272.6805, 272.5146, 272.4008, 272.4173, 271.283, 
    272.1083, 271.8528, 271.811, 271.4025, 271.8206, 272.1633, 272.0184, 
    272.299,
  273.4941, 272.9265, 272.8714, 272.5299, 272.713, 272.058, 273.0078, 
    269.3051, 267.9707, 271.8371, 271.6991, 272.0465, 271.2071, 271.3813, 
    272.0086,
  273.5731, 273.1185, 272.7321, 272.391, 272.5284, 272.579, 272.5929, 
    271.7448, 271.5901, 272.1447, 272.1198, 272.085, 271.9554, 271.6212, 
    272.1305,
  273.7881, 273.3144, 272.6595, 272.3463, 272.2632, 272.0812, 271.2947, 
    271.1643, 272.0436, 272.3127, 272.2304, 272.2108, 272.1025, 271.9655, 
    272.2064,
  273.9028, 273.518, 272.3841, 272.0585, 272.2865, 272.347, 272.3679, 
    272.2043, 272.1724, 272.2827, 272.1765, 272.1902, 272.151, 272.0744, 
    272.316,
  273.8706, 273.244, 272.1297, 272.1936, 272.277, 272.3062, 272.1449, 
    272.1771, 272.2545, 272.2211, 272.2025, 272.2263, 272.2904, 272.3448, 
    272.3859,
  273.6853, 272.9317, 272.3108, 272.4912, 272.5572, 272.493, 272.3812, 
    272.2055, 272.3826, 272.4828, 272.3968, 272.2175, 272.2222, 272.1903, 
    272.2564,
  277.5369, 273.3818, 273.2193, 272.0442, 271.5687, 271.1835, 271.05, 
    271.3865, 271.0708, 269.6523, 272.6482, 271.5807, 271.0027, 270.4098, 
    272.1257,
  272.9944, 272.5311, 272.403, 271.6505, 271.2977, 271.45, 271.6996, 
    271.9455, 271.7009, 271.7669, 272.2755, 271.6852, 267.7276, 270.6944, 
    271.6125,
  273.1082, 272.8756, 272.2185, 271.6359, 271.2899, 271.1037, 272.01, 
    272.1299, 272.1356, 271.9592, 271.7191, 271.5788, 268.185, 269.6037, 
    271.9675,
  273.3764, 272.8987, 272.2964, 272.0339, 271.6099, 272.0844, 269.7967, 
    272.2293, 272.0999, 271.5396, 271.8044, 271.6982, 269.7914, 270.8504, 
    272.6027,
  273.6176, 272.7348, 272.4293, 272.0965, 271.9533, 271.9644, 272.5992, 
    269.7699, 268.607, 270.5527, 271.6738, 270.6842, 270.3087, 271.8237, 
    272.9211,
  273.493, 272.6874, 272.234, 272.0264, 271.1972, 271.7314, 271.9822, 
    271.0581, 270.8687, 270.0444, 269.9283, 269.705, 271.5149, 272.7436, 
    273.0071,
  273.3467, 272.8869, 272.1279, 271.9428, 271.9701, 271.8357, 271.4931, 
    271.9234, 269.992, 269.8668, 271.3372, 271.6562, 272.4548, 272.9234, 
    273.0756,
  273.8453, 273.3476, 271.8872, 270.5163, 271.5374, 271.6595, 271.801, 
    271.7356, 271.5327, 271.7005, 271.7996, 272.4945, 272.7652, 272.9004, 
    272.9174,
  273.9779, 272.9256, 271.7874, 271.7921, 271.7695, 271.8332, 271.9807, 
    272.0326, 272.1987, 272.256, 272.5792, 272.7487, 272.8193, 272.8236, 
    272.7494,
  273.7538, 272.7844, 271.9732, 271.6991, 271.9905, 272.034, 271.6452, 
    271.9406, 272.3347, 272.6249, 272.7911, 272.7901, 272.7312, 272.6212, 
    272.4518,
  281.0288, 276.1098, 276.3989, 272.881, 272.3132, 271.4899, 270.5485, 
    270.3457, 270.2668, 271.2928, 271.8835, 271.7016, 269.1968, 271.3717, 
    271.7889,
  275.0149, 274.5425, 273.0891, 272.2146, 272.0809, 271.3105, 270.9218, 
    270.5905, 270.2885, 270.6082, 270.2749, 269.0166, 268.9295, 270.5964, 
    271.3201,
  274.5326, 273.7867, 272.932, 272.1864, 272.1079, 269.5319, 270.4854, 
    270.5632, 270.5991, 271.2644, 270.4787, 269.755, 270.8515, 270.6084, 
    271.875,
  274.2755, 273.6455, 272.9701, 272.3019, 271.9151, 271.6837, 268.5721, 
    270.6458, 270.9784, 271.1177, 269.8788, 270.8264, 270.6511, 271.3007, 
    272.5468,
  273.9117, 273.2037, 272.8111, 271.7886, 271.4673, 271.6198, 271.5668, 
    268.6836, 267.6341, 269.726, 271.8563, 270.6696, 270.6312, 272.0377, 
    272.9451,
  273.4172, 272.7686, 272.0349, 271.4853, 270.9172, 271.47, 271.8843, 
    271.128, 269.9649, 268.7127, 271.271, 270.196, 271.2336, 272.7235, 
    272.9499,
  273.0746, 272.6363, 271.8144, 271.449, 271.2352, 271.6495, 271.7286, 
    270.6496, 269.082, 268.8082, 270.2959, 270.7996, 272.4117, 272.8613, 
    273.0228,
  273.739, 273.1815, 271.256, 269.7458, 271.3252, 271.6678, 272.0882, 
    271.0208, 271.0141, 270.5094, 270.5166, 272.2144, 272.7587, 272.8776, 
    273.082,
  273.903, 273.087, 270.8241, 271.2002, 271.3706, 271.5659, 271.9076, 
    271.6109, 271.3497, 271.4117, 272.3145, 272.7691, 272.7763, 272.8676, 
    272.9301,
  273.4096, 272.6796, 271.5275, 271.5405, 271.6545, 271.6526, 271.3903, 
    271.7014, 271.3878, 272.2923, 272.8844, 272.8317, 272.7411, 272.699, 
    272.6203,
  282.7309, 278.1188, 279.108, 274.8434, 274.0837, 273.0396, 272.5157, 
    272.0844, 271.8811, 272.0907, 272.2159, 271.7269, 271.048, 270.8513, 
    270.9435,
  277.0132, 275.6672, 274.6312, 273.1424, 273.1927, 272.6594, 272.3847, 
    271.5756, 271.2877, 271.2432, 270.6449, 269.7143, 270.1881, 269.8603, 
    270.5463,
  275.6982, 274.882, 273.4871, 272.8357, 272.7927, 270.946, 271.7211, 
    271.6526, 271.013, 270.6717, 270.4205, 270.4028, 270.4203, 270.4835, 
    271.3938,
  275.6096, 274.6733, 273.4861, 272.923, 272.5483, 272.1609, 269.209, 
    270.3806, 270.297, 270.7643, 268.4195, 270.573, 270.747, 271.8339, 272.617,
  275.4379, 274.2098, 273.5381, 272.6261, 272.2711, 271.7278, 271.1944, 
    267.4675, 266.0978, 268.2342, 269.6168, 271.3636, 272.1933, 272.8176, 
    273.0662,
  275.0668, 273.9415, 272.9852, 272.08, 271.8893, 271.1914, 271.041, 
    270.5134, 269.7661, 269.0716, 270.5261, 271.6842, 272.7159, 272.9951, 
    273.0156,
  274.6217, 273.7133, 272.3721, 271.7884, 271.5911, 271.188, 270.7874, 269.2, 
    268.672, 269.0744, 271.2924, 272.7159, 272.9356, 272.9624, 273.1054,
  274.2798, 273.3391, 271.7034, 271.4043, 271.2224, 270.9768, 270.6438, 
    269.4478, 269.6439, 270.3224, 272.618, 272.8589, 272.84, 273.0241, 
    273.1502,
  273.9091, 272.7341, 271.3045, 271.2044, 271.0983, 270.9402, 270.7354, 
    269.1133, 270.0278, 270.8852, 272.8221, 272.8607, 272.8484, 272.9633, 
    273.0593,
  273.7704, 272.5889, 271.3076, 271.1165, 270.986, 271.0727, 270.7893, 
    270.6254, 270.475, 272.0567, 272.8834, 272.8818, 272.8395, 272.7728, 
    272.6827,
  278.944, 276.3396, 277.6743, 275.5344, 275.2468, 275.2078, 274.6311, 
    273.9219, 273.2587, 273.4155, 273.4726, 272.166, 271.5664, 271.1365, 
    270.0208,
  274.7561, 274.5406, 274.5931, 274.248, 274.7653, 273.6297, 273.6729, 
    273.229, 273.1292, 272.9653, 272.1819, 271.3701, 270.7388, 270.5808, 
    270.8585,
  275.2648, 274.7986, 274.2495, 274.2711, 273.5818, 272.9076, 272.9987, 
    272.9852, 272.4113, 271.6825, 271.2785, 270.538, 269.8232, 269.8928, 
    271.2902,
  275.5746, 274.7487, 274.0255, 273.6937, 273.2579, 273.384, 270.8593, 
    271.2538, 271.2258, 271.3025, 269.9304, 269.9939, 270.912, 271.4492, 
    271.8435,
  275.8243, 274.4418, 273.9829, 273.3959, 273.1856, 272.9036, 272.5986, 
    269.4361, 267.3468, 270.0028, 270.1671, 270.552, 271.3685, 272.2367, 
    272.5857,
  275.843, 274.4038, 273.3903, 272.9951, 272.7215, 272.4007, 272.1555, 
    272.0766, 270.5564, 269.9282, 270.049, 271.5396, 272.429, 272.856, 
    272.9937,
  275.6374, 274.3945, 273.015, 272.2196, 271.44, 270.4868, 270.3054, 
    270.2523, 270.4498, 270.9454, 271.9573, 272.7314, 272.9068, 272.8813, 
    272.8098,
  275.47, 274.0419, 272.1873, 271.2927, 270.4295, 270.1628, 270.5435, 
    270.9978, 271.4125, 272.452, 272.8543, 272.8928, 272.8483, 272.8657, 
    272.8421,
  274.6194, 272.8917, 271.2628, 270.6343, 270.3514, 270.3773, 270.4628, 
    270.7946, 271.7882, 272.8158, 272.9469, 272.899, 272.8713, 272.8636, 
    272.9106,
  273.7849, 272.5441, 271.3432, 270.4461, 270.4762, 270.5428, 270.6439, 
    271.491, 272.1606, 272.8917, 273.0034, 272.8817, 272.7635, 272.7015, 
    272.6738,
  278.6324, 276.2658, 277.5432, 274.8576, 274.6649, 274.5632, 273.7646, 
    273.7367, 274.2473, 274.2245, 274.6508, 273.643, 272.9178, 272.9035, 
    273.1302,
  275.2379, 274.5393, 274.8252, 274.5014, 274.5746, 273.5565, 273.4518, 
    273.7799, 273.9264, 273.8433, 273.7878, 273.3005, 273.0772, 272.3707, 
    272.3553,
  275.3192, 274.9968, 274.6817, 274.2684, 274.0468, 273.0491, 273.0623, 
    273.4755, 273.7189, 273.7581, 273.5247, 273.1714, 272.755, 272.4911, 
    272.2925,
  275.4486, 275.0459, 274.5351, 274.2305, 273.7321, 273.8129, 273.3104, 
    273.3692, 273.6378, 273.3766, 273.1405, 273.1144, 273.0438, 272.6674, 
    271.6602,
  275.5426, 274.7079, 274.4094, 273.8889, 273.7346, 272.7387, 273.1599, 
    272.8346, 271.9309, 272.971, 272.9501, 272.812, 272.3494, 271.8303, 
    271.7656,
  275.342, 274.5323, 273.7642, 273.4203, 273.4623, 273.522, 273.5121, 
    273.7884, 272.6073, 272.4, 272.3415, 272.0553, 271.8883, 271.7688, 
    271.9914,
  275.0542, 274.349, 273.2198, 272.9238, 272.7944, 272.571, 272.3906, 
    271.9634, 271.6845, 271.7928, 271.9175, 271.9078, 271.9889, 272.2472, 
    272.3087,
  274.6028, 273.6268, 272.1438, 271.8729, 271.9957, 272.0348, 271.9251, 
    271.8432, 271.8756, 272.1164, 272.2796, 272.3207, 272.4274, 272.5836, 
    272.5719,
  273.9849, 272.8727, 271.9373, 272.0546, 272.3486, 272.4149, 272.328, 
    272.3896, 272.701, 272.703, 272.6613, 272.7137, 272.7689, 272.72, 272.7439,
  273.5495, 272.6275, 272.0128, 272.1064, 272.5172, 272.7903, 272.9254, 
    272.9163, 273.0684, 273.0622, 273.0063, 272.815, 272.5548, 272.3902, 
    272.7242,
  277.4955, 274.8133, 276.4389, 273.8383, 273.5662, 274.1981, 274.2335, 
    273.8008, 273.4438, 273.4537, 274.7176, 274.2914, 273.9018, 274.3683, 
    274.0991,
  274.4497, 273.8282, 273.6263, 273.1153, 273.4453, 273.5237, 273.5961, 
    273.4364, 273.1277, 273.2837, 274.0858, 273.9008, 273.782, 273.6689, 
    273.5132,
  275.0403, 274.6062, 273.9139, 273.0731, 273.3177, 272.9004, 273.5211, 
    273.3196, 273.2816, 273.1227, 273.5695, 273.536, 273.3765, 273.7339, 
    273.3465,
  275.4576, 274.8904, 274.3109, 273.7395, 273.2124, 273.4856, 273.1484, 
    273.4802, 273.3564, 273.3295, 273.5305, 273.5916, 272.947, 273.4317, 
    273.32,
  275.8363, 274.7279, 274.1664, 273.3967, 273.3075, 273.1667, 273.9028, 
    273.2378, 272.7483, 273.4589, 273.4561, 273.3255, 273.251, 273.182, 
    273.0528,
  275.594, 274.5361, 273.528, 273.0288, 273.2546, 273.1744, 273.3857, 
    273.5379, 273.443, 273.3247, 273.5551, 273.3638, 273.1974, 272.9895, 
    272.7623,
  275.3983, 274.4842, 273.1443, 272.8033, 272.8862, 272.9408, 273.0008, 
    273.0951, 273.1431, 273.189, 273.3279, 273.1809, 272.9198, 272.5571, 
    272.3711,
  275.0287, 274.0763, 272.754, 272.5665, 272.6889, 272.7773, 272.8257, 
    272.9065, 272.963, 273.0466, 273.022, 272.7637, 272.4347, 272.1507, 
    272.1638,
  274.6178, 273.6413, 272.6914, 272.6391, 272.5831, 272.5634, 272.5993, 
    272.6435, 272.7437, 272.7475, 272.611, 272.5276, 272.3727, 272.4156, 
    272.5829,
  274.2483, 273.5837, 272.8918, 272.7803, 272.7425, 272.6864, 272.5065, 
    272.4428, 272.7018, 272.8384, 272.8128, 272.5431, 272.4807, 272.5222, 
    272.9637,
  276.9589, 274.3407, 275.5536, 274.1785, 274.1811, 275.5807, 275.2131, 
    274.7699, 275.3344, 273.5395, 273.7555, 274.6011, 274.8164, 275.1697, 
    274.6933,
  274.2654, 273.7094, 273.6034, 273.2421, 273.6009, 273.9825, 274.5695, 
    274.2477, 274.0902, 272.6083, 273.2726, 273.9842, 274.7683, 274.5193, 
    273.9285,
  274.9788, 274.6098, 274.1047, 273.0047, 273.2577, 273.1972, 273.8277, 
    273.8275, 273.8719, 272.3851, 273.0888, 273.5948, 274.2384, 274.6057, 
    273.9375,
  275.0158, 274.4498, 273.9164, 273.3796, 273.0275, 274.0497, 273.242, 
    273.1875, 273.2041, 272.4156, 273.2545, 273.4597, 273.6397, 274.101, 
    273.7557,
  274.7989, 274.0638, 273.5987, 273.0666, 272.9149, 273.4113, 274.574, 
    272.8716, 272.5757, 272.9471, 273.2838, 273.3586, 273.5347, 273.835, 
    274.2405,
  274.5071, 273.9286, 273.208, 272.5843, 272.8241, 273.2157, 274.1853, 
    274.5047, 274.3502, 273.5899, 273.4176, 273.3642, 273.3464, 273.6215, 
    273.8032,
  274.3107, 273.8628, 272.9013, 272.5696, 272.784, 273.2196, 273.9068, 
    274.163, 273.9167, 273.4315, 273.2923, 273.0418, 273.2227, 273.4998, 
    273.3776,
  274.0475, 273.54, 272.5601, 272.673, 272.8728, 273.2292, 273.5752, 
    273.8388, 273.5816, 273.1812, 273.013, 272.7692, 273.071, 273.1211, 
    272.9098,
  273.6457, 272.8924, 272.1774, 272.6223, 272.9869, 273.2417, 273.3745, 
    273.2084, 272.9489, 272.9286, 273.1309, 272.7584, 272.957, 272.983, 
    272.9675,
  273.0927, 272.3925, 271.8287, 272.169, 272.7497, 273.0387, 273.0473, 
    272.9753, 272.9719, 272.9648, 272.7475, 272.8554, 272.8304, 272.8514, 
    273.062,
  277.4546, 274.7606, 275.1194, 273.5916, 273.6753, 274.013, 273.6114, 
    273.33, 273.8259, 273.7924, 274.5927, 274.3599, 273.8692, 274.3101, 
    274.2171,
  275.0009, 274.1519, 274.0542, 273.3297, 273.4685, 273.3977, 273.357, 
    273.2118, 273.3311, 273.5352, 274.0901, 273.879, 273.8975, 273.8475, 
    273.9448,
  275.6708, 275.3092, 274.6026, 273.3728, 273.3048, 272.4861, 273.5543, 
    273.3758, 273.4002, 273.1779, 272.8582, 273.148, 273.7263, 274.1644, 
    274.2664,
  275.893, 275.2634, 274.5173, 273.9745, 273.1753, 273.3229, 272.685, 
    272.9717, 273.3472, 272.799, 273.0127, 273.3026, 273.6275, 273.8601, 
    273.774,
  275.5748, 274.8334, 274.5059, 273.6864, 273.3327, 273.015, 273.7086, 
    272.4108, 273.048, 273.1104, 272.8103, 273.2512, 273.5636, 273.8496, 
    274.4011,
  275.0954, 274.7539, 274.0483, 273.0954, 273.1239, 273.074, 273.3204, 
    274.0836, 274.1973, 273.0144, 273.1516, 273.2676, 273.5423, 273.7585, 
    274.0045,
  275.0429, 274.7777, 273.479, 272.5164, 272.7856, 273.0333, 273.2966, 
    273.6644, 273.2601, 272.7821, 273.0265, 273.2798, 273.4721, 273.4986, 
    273.3677,
  275.041, 274.4577, 272.7449, 272.3536, 272.7011, 273.0355, 273.2751, 
    273.3819, 273.1389, 272.9232, 273.0724, 273.1516, 273.3128, 273.1011, 
    272.963,
  274.8153, 273.8537, 272.7369, 272.7641, 272.9081, 273.1499, 273.2766, 
    273.0897, 273.0095, 272.9294, 273.1052, 273.0963, 273.1559, 273.036, 
    273.082,
  274.2951, 273.7269, 273.1513, 273.1003, 273.1305, 273.1568, 272.9449, 
    272.9086, 272.9796, 273.0786, 272.9685, 273.0342, 273.0871, 273.005, 
    273.1197,
  281.009, 276.977, 278.2149, 275.4567, 274.9714, 275.7317, 274.6318, 
    274.0632, 273.7052, 273.2777, 273.666, 273.949, 273.3545, 273.4802, 
    273.4173,
  276.6488, 275.0962, 274.9353, 273.7924, 274.2843, 274.6385, 274.1932, 
    273.8242, 273.4119, 273.2219, 273.4716, 273.4785, 273.3164, 273.1008, 
    273.463,
  276.1265, 275.7091, 275.0758, 273.7884, 273.8053, 273.2328, 274.0877, 
    273.8896, 273.575, 273.1487, 273.0287, 273.2434, 273.2256, 273.3368, 
    273.4317,
  276.1466, 275.5873, 274.8403, 274.3345, 273.5103, 273.6356, 272.7428, 
    273.7761, 273.316, 273.1743, 273.1215, 273.1835, 273.1617, 273.1238, 
    273.1835,
  276.041, 275.1831, 274.8289, 273.9243, 273.5846, 273.2273, 273.3379, 
    271.3948, 271.916, 273.8693, 273.1996, 273.2439, 273.2243, 273.1357, 
    273.359,
  275.8442, 275.0981, 274.3864, 273.2511, 273.2712, 273.2741, 273.16, 
    273.4402, 273.9274, 273.5415, 273.3747, 272.9967, 272.7715, 273.056, 
    273.3896,
  275.7198, 275.1604, 273.6759, 272.4245, 272.5834, 272.9337, 273.069, 
    273.118, 273.1864, 273.0937, 273.0437, 272.9247, 272.8802, 272.9373, 
    273.2114,
  275.5666, 274.625, 272.7487, 272.0607, 272.5142, 272.8561, 272.9747, 
    272.9394, 272.9675, 273.0066, 272.9745, 273.0015, 272.9786, 272.94, 
    273.1089,
  275.1314, 273.9211, 272.6658, 272.7249, 272.8095, 272.9454, 272.9468, 
    272.9261, 272.9949, 272.9841, 273.0712, 272.9705, 272.9328, 273.0157, 
    273.4224,
  274.5534, 273.7775, 273.0843, 272.9775, 272.9452, 272.8965, 272.7599, 
    272.7492, 272.9254, 273.0923, 273.1084, 272.9581, 272.9472, 273.0783, 
    273.4431,
  282.1683, 278.3808, 280.5246, 276.2599, 276.1852, 277.4785, 275.5445, 
    274.5119, 274.9568, 277.0871, 277.0802, 276.0242, 273.4752, 274.2448, 
    273.7897,
  277.3745, 276.4707, 276.4392, 274.8527, 276.2217, 276.6189, 274.0771, 
    273.8005, 274.1172, 275.1594, 274.7444, 273.5326, 273.2015, 272.379, 
    272.6863,
  276.1835, 275.8417, 274.9711, 273.9156, 274.7308, 274.1812, 273.7401, 
    273.6313, 273.6438, 273.5484, 272.726, 272.7992, 272.4384, 272.629, 
    272.8886,
  275.8271, 275.4258, 274.7216, 274.3307, 273.6127, 274.4351, 273.4335, 
    273.3424, 273.0116, 272.5842, 272.3643, 272.344, 272.1436, 272.5571, 
    272.9998,
  276.1131, 275.2761, 274.8516, 273.709, 273.412, 273.3187, 273.9759, 
    272.821, 272.485, 272.7937, 272.357, 271.9555, 272.3849, 272.6218, 
    272.7863,
  276.1784, 275.3741, 274.5025, 273.2789, 273.2731, 273.2746, 273.283, 
    274.0628, 274.4165, 273.5984, 272.5556, 272.2349, 271.3528, 272.5541, 
    272.9077,
  276.0933, 275.6526, 274.0593, 272.8406, 272.6356, 272.9683, 273.1223, 
    273.3735, 273.6835, 273.2835, 273.3287, 272.7433, 272.327, 272.53, 
    272.5329,
  276.4693, 275.6816, 273.6377, 272.824, 272.7157, 272.8079, 272.9108, 
    272.9951, 273.2118, 273.4784, 273.3509, 273.092, 272.7034, 272.3909, 
    272.2313,
  276.2486, 274.9833, 273.3385, 273.1068, 272.946, 272.8769, 272.8667, 
    272.9682, 273.1639, 273.3878, 273.4059, 273.1024, 272.614, 272.4471, 
    272.3772,
  275.4481, 274.5461, 273.4732, 273.1658, 272.9825, 272.8806, 272.7614, 
    272.8373, 273.1598, 273.4438, 273.3317, 272.8497, 272.7184, 272.5085, 
    272.3547,
  277.413, 275.8911, 278.1665, 274.9634, 276.1333, 277.151, 275.4233, 
    275.658, 276.6909, 279.6246, 278.2509, 276.8425, 274.0941, 273.7607, 
    274.3322,
  275.1944, 275.3004, 275.6065, 275.0565, 277.1445, 276.4376, 274.5208, 
    274.6865, 274.982, 275.8594, 276.2511, 272.7846, 271.5501, 272.0829, 
    272.9751,
  275.522, 275.6554, 274.9984, 274.5157, 275.2505, 273.5183, 273.8611, 
    273.5865, 273.672, 273.3853, 272.9673, 271.6731, 271.1793, 272.9483, 
    273.2946,
  275.3769, 275.2885, 274.9274, 274.6775, 274.2541, 274.656, 273.1189, 
    273.2126, 273.2504, 272.6383, 272.0256, 271.3706, 271.357, 273.0716, 
    273.4353,
  275.1689, 274.6419, 274.4815, 273.8854, 273.9259, 273.9996, 274.7205, 
    273.1236, 272.0209, 272.2861, 271.8468, 271.516, 271.7616, 272.8429, 
    272.8813,
  275.1631, 274.3968, 273.6047, 273.1022, 273.3781, 273.6914, 274.1055, 
    274.5197, 274.1824, 272.7156, 271.5113, 271.0296, 272.1683, 272.5926, 
    272.3904,
  275.296, 274.607, 273.1842, 272.5565, 272.7956, 273.4315, 273.6654, 
    273.9507, 273.2756, 272.2747, 271.8138, 272.0263, 271.9185, 271.7161, 
    271.5117,
  276.7786, 274.9331, 273.0212, 272.6048, 272.9062, 273.2895, 273.4166, 
    273.444, 272.8528, 272.7151, 272.1833, 272.1064, 271.6705, 271.4893, 
    271.3887,
  276.779, 275.0419, 273.202, 273.1982, 273.1614, 273.2826, 273.316, 
    273.3419, 273.2169, 273.1405, 272.5432, 272.0625, 271.6686, 271.472, 
    271.2442,
  276.0896, 275.1122, 273.6969, 273.5073, 273.3214, 273.3157, 273.1906, 
    273.2401, 273.371, 273.3163, 272.7639, 272.0296, 271.7393, 271.2808, 
    271.0758,
  277.4112, 274.4494, 275.3567, 273.5024, 274.7116, 275.2368, 273.8899, 
    274.463, 275.2202, 277.3068, 278.0158, 276.7703, 275.6353, 275.7907, 
    276.2288,
  274.8659, 274.4921, 274.362, 273.8831, 275.6784, 275.1119, 273.5754, 
    273.7552, 274.0969, 274.8022, 276.2263, 274.2322, 274.149, 273.5107, 
    273.9451,
  275.7017, 275.3299, 274.5617, 273.9886, 274.6007, 273.0482, 273.2981, 
    273.1017, 273.1031, 272.976, 272.9151, 272.8363, 273.3364, 273.7332, 
    273.5342,
  276.1435, 275.4959, 274.5964, 274.4769, 273.4797, 273.9174, 272.1546, 
    272.4022, 272.2809, 272.3095, 272.4443, 272.8432, 273.3869, 273.3798, 
    273.4716,
  276.3478, 275.2802, 274.3746, 273.8356, 273.5116, 273.701, 274.3492, 
    271.9216, 269.0336, 271.8892, 272.2876, 272.6071, 272.688, 272.4863, 
    272.2698,
  276.4842, 275.4043, 273.8997, 273.3466, 273.4536, 273.6348, 273.7519, 
    273.4372, 272.0142, 271.7346, 271.8148, 272.0474, 272.0302, 271.7119, 
    271.4056,
  276.7931, 275.7438, 273.4005, 272.8018, 273.0033, 273.3879, 273.1968, 
    272.4905, 271.5724, 271.4851, 271.7534, 271.7527, 271.2724, 270.5103, 
    270.3757,
  277.227, 275.7789, 272.5748, 272.4464, 272.71, 273.1785, 272.6087, 
    271.8315, 271.2904, 271.3972, 271.3982, 271.1816, 270.7794, 270.5501, 
    270.4578,
  277.0854, 274.9702, 272.629, 272.7923, 272.9152, 273.0551, 272.4835, 
    271.792, 271.5366, 271.4111, 271.3408, 270.9951, 270.8048, 270.5694, 
    270.635,
  276.3101, 274.7867, 273.0973, 273.1483, 273.1499, 273.0868, 272.298, 
    271.8279, 271.6194, 271.838, 271.2808, 270.8686, 270.6447, 270.36, 
    270.8501,
  282.0842, 275.9265, 276.287, 273.7544, 274.3206, 275.274, 273.9896, 
    274.6856, 275.5384, 278.889, 279.0223, 277.7117, 277.3534, 276.9318, 
    276.2442,
  276.2737, 274.8321, 274.7643, 274.0085, 275.9784, 275.0513, 273.7115, 
    273.9841, 273.9423, 275.331, 276.9421, 275.1049, 274.8508, 273.6274, 
    274.5994,
  276.2508, 275.2691, 274.6897, 274.0301, 275.7177, 273.0119, 273.4161, 
    273.2598, 273.3123, 273.7513, 274.3278, 273.2635, 272.9352, 272.7897, 
    272.6553,
  276.4895, 275.6251, 274.7517, 274.3788, 273.8321, 274.1756, 272.5236, 
    272.9071, 273.2513, 273.4554, 273.3165, 272.9435, 272.3779, 272.1848, 
    272.2784,
  276.3342, 275.2973, 274.6811, 273.8848, 273.2236, 273.3972, 273.9073, 
    270.9517, 270.2778, 273.1342, 272.895, 272.0456, 271.3727, 271.0631, 
    271.7614,
  276.1038, 275.1956, 274.2348, 273.0865, 272.8884, 273.1801, 273.4366, 
    273.5885, 273.3264, 272.7565, 272.2662, 271.1153, 270.7964, 270.5536, 
    271.8064,
  275.8905, 275.1158, 273.4742, 272.6044, 272.542, 272.8378, 273.0485, 
    272.6326, 272.4576, 271.9901, 271.6607, 270.564, 269.888, 270.2802, 
    271.233,
  275.7043, 274.6849, 272.5966, 272.2618, 272.3212, 272.7236, 272.5137, 
    272.1339, 271.9688, 271.3496, 271.1489, 270.3171, 270.5045, 271.0952, 
    272.0202,
  275.5763, 273.8698, 272.3278, 272.3851, 272.5379, 272.6595, 271.9705, 
    271.9675, 271.5638, 271.1299, 270.5864, 270.5448, 270.7853, 271.7282, 
    272.1042,
  275.4204, 274.0738, 272.7596, 272.8541, 272.8466, 272.6017, 271.6995, 
    271.5682, 271.1942, 270.9157, 270.5882, 270.522, 271.0446, 271.999, 
    272.5392,
  276.9368, 274.3329, 275.3098, 273.4884, 274.6053, 275.5488, 274.2768, 
    274.0498, 274.739, 279.6368, 279.7157, 277.7118, 276.8689, 276.1599, 
    276.0065,
  274.1651, 273.7573, 273.7599, 273.3907, 275.1487, 275.3448, 273.7095, 
    273.7926, 273.9164, 275.9174, 278.4282, 275.6581, 274.5002, 272.8832, 
    273.3025,
  274.6143, 274.1962, 273.8711, 273.4091, 273.9305, 272.2707, 273.8565, 
    273.6558, 273.7191, 274.069, 275.4803, 274.0091, 273.2191, 272.2075, 
    272.0099,
  275.157, 274.7852, 274.2828, 273.864, 273.0757, 273.4312, 272.3062, 
    273.3668, 273.443, 273.5783, 273.8318, 273.2191, 272.4145, 271.4621, 
    272.4754,
  275.3889, 274.8508, 274.64, 273.9501, 273.1641, 272.9428, 273.2311, 
    271.5993, 271.584, 273.5447, 273.3266, 272.7911, 272.0692, 271.6331, 
    272.2007,
  276.1528, 275.7614, 274.9773, 274.0243, 273.3266, 273.1398, 272.9191, 
    273.3265, 273.6198, 273.3458, 273.0314, 272.3684, 271.5469, 271.2687, 
    272.2278,
  276.8197, 276.2676, 274.6891, 273.6623, 273.1938, 272.8397, 273.0933, 
    273.1575, 273.0753, 272.7263, 272.3745, 271.6661, 270.8992, 271.3383, 
    271.7148,
  277.0385, 276.2597, 274.5065, 273.2837, 272.9041, 272.7525, 272.9854, 
    272.8385, 272.7157, 272.5098, 271.9606, 270.9127, 270.9584, 271.5185, 
    271.9979,
  276.881, 275.579, 273.5342, 272.8767, 272.5717, 272.565, 272.7337, 
    272.7655, 272.7185, 272.1998, 271.2338, 270.6813, 271.2487, 271.8035, 
    271.9283,
  276.0552, 274.9509, 273.1321, 272.597, 272.6143, 272.5839, 272.4412, 
    272.3734, 272.1136, 271.3981, 270.8187, 270.8296, 271.9537, 272.2411, 
    272.6148,
  281.1896, 277.581, 279.4959, 275.43, 275.1585, 275.3061, 274.3859, 
    274.3095, 275.1422, 278.3439, 280.5235, 279.6817, 279.5896, 277.6216, 
    276.5907,
  274.7824, 274.4923, 274.31, 273.6859, 274.2878, 273.3712, 272.962, 
    273.1745, 273.3574, 274.4145, 277.423, 276.3257, 276.5692, 275.5572, 
    275.7352,
  274.5222, 274.2043, 273.8306, 273.4759, 274.2712, 271.4646, 272.2473, 
    272.1533, 272.588, 272.7295, 273.7983, 274.015, 274.0844, 274.5166, 
    274.6463,
  274.4851, 274.0064, 273.4735, 273.2317, 272.7391, 273.0799, 270.596, 
    271.9374, 272.2136, 272.287, 272.7903, 273.1128, 273.3846, 273.4781, 
    273.3884,
  274.352, 274.0323, 273.9236, 273.4224, 272.8018, 272.4726, 272.5388, 
    269.8124, 270.1139, 272.9739, 272.375, 272.6015, 273.095, 272.9629, 
    272.803,
  275.2727, 275.2585, 274.7018, 273.9055, 273.1361, 273.185, 272.8919, 
    272.8892, 273.2592, 273.0665, 272.5016, 272.5095, 272.9106, 272.6808, 
    272.6289,
  276.5361, 276.0097, 274.267, 273.1989, 273.0511, 272.6727, 272.8978, 
    272.945, 272.8258, 272.5854, 272.3827, 272.5488, 272.7157, 272.4486, 
    272.4507,
  276.71, 275.9047, 273.867, 272.9135, 272.7563, 272.501, 272.6296, 272.6018, 
    272.5728, 272.6675, 272.6049, 272.5703, 272.5806, 272.1828, 271.8893,
  275.9953, 274.9725, 273.4719, 272.9148, 272.6599, 272.3677, 272.4032, 
    272.6108, 272.7248, 272.7635, 272.7617, 272.6846, 272.4259, 271.7821, 
    271.6832,
  275.1795, 274.5719, 273.5357, 272.7595, 272.7271, 272.6467, 272.3693, 
    272.6801, 272.8483, 272.8689, 272.7733, 272.5004, 272.0568, 271.6955, 
    272.0878,
  276.7419, 274.9318, 275.994, 274.8104, 274.7308, 275.8505, 275.2771, 
    274.9596, 275.168, 278.7115, 280.8768, 280.7196, 281.9099, 281.3122, 
    279.2043,
  274.5888, 274.3811, 274.5269, 273.9082, 275.0638, 275.2567, 274.2283, 
    274.1393, 274.1181, 275.3333, 277.8554, 276.609, 277.2746, 278.5142, 
    278.4261,
  274.8337, 274.569, 274.0688, 273.5686, 274.4419, 272.761, 273.7071, 
    273.4095, 273.3332, 273.5268, 274.4646, 274.1786, 274.2105, 275.2354, 
    276.3809,
  274.9285, 274.2709, 273.5161, 273.2402, 272.7986, 273.4925, 271.7552, 
    272.6807, 272.51, 272.6824, 272.8593, 272.945, 273.2643, 273.5198, 
    274.1386,
  275.1821, 274.2924, 273.5461, 272.717, 272.1406, 272.3395, 273.3091, 
    270.9355, 270.0109, 272.2296, 272.1721, 272.024, 272.828, 273.1056, 
    273.5254,
  275.4567, 274.5862, 273.5112, 272.6731, 272.1925, 272.2955, 272.4693, 
    272.7797, 272.9023, 272.2824, 272.0982, 271.9275, 272.4821, 272.9091, 
    273.0374,
  275.6043, 274.7491, 272.9835, 272.2781, 272.2048, 272.0386, 272.2779, 
    272.3637, 272.3348, 272.0918, 272.0964, 272.067, 272.3203, 272.6082, 
    272.9813,
  275.426, 274.6035, 272.7708, 272.2428, 272.2429, 272.0757, 272.2913, 
    272.3271, 272.2981, 272.2307, 272.3317, 272.454, 272.5209, 272.7209, 
    272.8076,
  274.9652, 273.9247, 272.6077, 272.4388, 272.4198, 272.2542, 272.4325, 
    272.6568, 272.6742, 272.6913, 272.6743, 272.6176, 272.6205, 272.4603, 
    272.3932,
  274.2934, 273.6971, 272.8148, 272.697, 272.6199, 272.5818, 272.5277, 
    272.8164, 272.9271, 272.834, 272.7696, 272.6042, 272.4783, 272.2133, 
    272.4498,
  274.7142, 273.5056, 273.8661, 272.6176, 273.3058, 274.0805, 272.8782, 
    272.7412, 272.8883, 274.262, 275.5575, 275.4681, 275.6734, 276.6014, 
    277.9768,
  273.7766, 273.4608, 273.4572, 273.0129, 273.7958, 274.1081, 272.9701, 
    272.9029, 272.9151, 273.4245, 274.8344, 274.6742, 274.2815, 274.11, 
    275.9662,
  274.7725, 274.3805, 274.0797, 273.4024, 273.4914, 271.3285, 273.4123, 
    273.0252, 273.0488, 272.8959, 273.323, 273.6103, 273.3092, 273.4398, 
    274.5141,
  275.544, 275.1896, 274.3606, 273.7307, 272.8489, 272.9918, 271.0444, 
    273.0097, 273.3656, 273.0434, 273.2071, 273.1971, 273.2082, 273.1887, 
    273.4861,
  276.2728, 275.3286, 274.6691, 273.6389, 272.5218, 272.4919, 272.7325, 
    269.9002, 269.5667, 273.3187, 273.2492, 273.2473, 273.2174, 273.0936, 
    273.2735,
  276.4297, 275.4028, 274.2609, 272.9234, 272.1574, 272.1151, 272.3514, 
    272.4737, 272.5771, 272.8388, 273.1634, 273.2939, 273.2377, 273.3227, 
    273.4555,
  276.2991, 275.5002, 273.4684, 272.3014, 272.1858, 272.0815, 272.1481, 
    272.4058, 272.5139, 272.61, 272.9449, 273.2032, 273.118, 273.0774, 
    273.2329,
  275.9574, 275.0152, 272.8762, 272.2182, 272.2765, 272.1836, 272.3334, 
    272.2849, 272.5204, 272.8311, 273.0626, 273.1085, 273.0362, 273.023, 
    273.0916,
  275.2373, 273.5213, 272.6164, 272.3488, 272.3819, 272.1677, 272.4636, 
    272.5726, 272.7849, 272.9449, 273.0013, 272.9629, 272.8802, 272.7711, 
    272.876,
  274.5822, 273.3768, 272.7934, 272.6258, 272.4845, 272.5315, 272.3034, 
    272.5941, 272.6964, 272.877, 272.869, 272.8023, 272.7026, 272.7461, 
    272.8948,
  278.5395, 276.479, 279.4326, 275.8873, 276.3543, 278.8189, 275.4162, 
    274.7484, 274.9689, 277.1114, 277.1844, 275.7746, 275.1554, 275.3896, 
    275.7722,
  273.8018, 274.2645, 274.9863, 274.5919, 276.6163, 275.7685, 273.7536, 
    273.5434, 273.5923, 274.5732, 275.7246, 274.4792, 273.6518, 273.4533, 
    274.3964,
  273.7671, 273.9109, 273.8863, 273.6882, 274.6126, 272.3395, 273.1249, 
    272.965, 273.0123, 273.0916, 273.5439, 273.341, 272.981, 273.1696, 
    274.1084,
  274.082, 273.5398, 273.1925, 273.1978, 273.0198, 273.7164, 271.5427, 
    272.3826, 272.8522, 272.9167, 273.0818, 273.0633, 272.6543, 272.8032, 
    273.7515,
  274.6781, 273.7856, 273.2716, 272.7065, 272.2558, 272.6691, 273.5049, 
    270.2296, 269.8669, 273.2649, 273.0387, 273.1996, 272.6686, 272.6997, 
    272.9314,
  275.3098, 274.3127, 273.3603, 272.4978, 272.0602, 272.0476, 272.5344, 
    273.2063, 273.3996, 272.9284, 272.5252, 273.1825, 272.7556, 272.694, 
    272.8004,
  275.5703, 274.4872, 272.8136, 272.1293, 272.117, 272.088, 272.0573, 
    272.3798, 272.4979, 272.4022, 272.5075, 272.562, 272.1577, 272.3042, 
    272.8752,
  275.7938, 274.4902, 272.5999, 271.852, 271.8177, 271.6949, 271.4396, 
    271.5421, 272.383, 272.5944, 272.653, 272.3648, 272.0517, 272.7735, 
    272.8151,
  275.0605, 273.4021, 272.5606, 272.231, 271.9593, 271.5803, 271.3965, 
    271.9166, 272.6527, 272.7816, 272.3068, 272.0781, 272.7968, 272.7122, 
    272.7988,
  274.4427, 273.5149, 272.6525, 272.435, 272.2116, 272.0909, 271.4458, 
    272.0365, 272.4533, 272.5714, 272.1851, 272.5099, 272.5778, 272.6424, 
    272.8147,
  275.7838, 274.4841, 276.2236, 274.2589, 274.9445, 279.1842, 277.7292, 
    277.7664, 278.6954, 286.8314, 285.981, 282.3589, 280.5448, 278.4476, 
    277.6192,
  274.0856, 273.9298, 274.2139, 273.9238, 277.5114, 279.9297, 275.5797, 
    275.9511, 276.5008, 279.7628, 284.2606, 278.7618, 276.9433, 276.8132, 
    276.5449,
  274.4229, 274.2975, 274.2622, 273.8722, 276.5, 275.5232, 275.104, 274.4415, 
    274.8102, 276.0905, 277.6263, 275.9025, 274.9469, 274.7162, 275.1866,
  274.588, 274.0179, 273.7543, 273.9963, 274.0177, 277.3329, 274.0831, 
    274.0082, 273.9797, 274.3484, 274.5722, 274.034, 273.6043, 273.3686, 
    274.4146,
  274.6616, 273.5708, 273.3923, 273.0911, 272.8734, 273.9818, 275.252, 
    274.1364, 274.213, 275.5619, 273.8004, 273.5905, 272.9954, 272.8294, 
    273.2809,
  274.8767, 273.462, 272.7469, 272.6418, 272.4726, 272.9081, 273.7901, 
    275.0489, 276.2475, 274.3457, 273.5322, 273.097, 272.7437, 272.5543, 
    272.6545,
  274.9429, 273.4691, 272.3105, 272.1155, 272.4459, 272.4561, 272.7656, 
    273.5305, 273.5143, 273.0587, 273.0153, 272.7537, 272.4153, 272.6008, 
    272.6761,
  274.8519, 273.3354, 272.1124, 271.9786, 272.1972, 272.3546, 272.4295, 
    272.8469, 272.8492, 272.7999, 272.6701, 272.399, 272.4277, 272.5606, 
    272.6886,
  274.606, 272.915, 271.9243, 271.6517, 271.7858, 271.9411, 272.501, 
    272.7742, 272.6926, 272.592, 272.2634, 272.2041, 272.6723, 272.6634, 
    272.8816,
  274.6513, 273.1498, 271.7807, 271.6589, 271.6659, 271.7884, 272.1548, 
    272.395, 272.4277, 272.2292, 271.8759, 272.0222, 272.3194, 272.7665, 
    273.0433,
  274.5531, 273.9082, 275.1693, 273.8772, 275.9049, 278.1309, 276.6096, 
    277.1342, 278.3835, 288.9897, 289.9384, 286.4744, 287.7094, 285.3973, 
    284.0612,
  273.7161, 273.5247, 273.5895, 273.792, 277.3328, 277.8493, 274.2485, 
    275.1209, 275.5088, 279.2035, 288.2575, 283.4916, 281.5548, 284.7459, 
    282.8891,
  274.0694, 273.8447, 273.6272, 273.17, 274.0638, 273.2681, 275.1169, 
    273.9768, 274.223, 275.2444, 278.5016, 278.0799, 277.0774, 278.6658, 
    279.934,
  274.5241, 273.701, 273.3506, 273.2589, 272.5341, 274.1667, 273.1835, 
    275.2141, 274.4514, 274.0536, 274.9124, 275.6161, 275.1883, 276.4946, 
    277.8085,
  274.9988, 273.6831, 273.224, 272.9958, 272.1016, 272.1936, 273.2354, 
    273.1579, 274.2109, 276.3767, 273.9178, 274.3756, 274.312, 274.7624, 
    275.2376,
  275.575, 274.1021, 272.6914, 272.7464, 271.9486, 271.9828, 272.2008, 
    272.8714, 274.7385, 274.4859, 275.3904, 274.0205, 273.8312, 273.8438, 
    274.2018,
  276.1656, 274.6571, 272.3309, 272.3885, 272.0833, 272.0826, 272.0546, 
    272.4389, 272.8131, 273.2111, 273.6204, 273.8609, 273.6297, 273.5282, 
    273.6291,
  276.584, 274.5716, 272.2996, 272.2624, 272.1088, 272.1835, 272.0663, 
    272.3079, 272.7226, 273.1684, 273.3856, 273.5156, 273.4786, 273.3389, 
    273.3329,
  276.6154, 273.9876, 272.1667, 272.3538, 271.9951, 272.1348, 272.203, 
    272.6364, 272.9994, 273.2644, 273.3204, 273.3343, 273.2621, 273.1588, 
    273.3308,
  275.9127, 273.5032, 272.2628, 272.4909, 272.3925, 272.2303, 272.1942, 
    272.5692, 272.9053, 273.2432, 273.3409, 273.174, 273.0774, 273.0759, 
    273.5084,
  273.7809, 274.0355, 277.0442, 276.5415, 278.0437, 280.3691, 277.4945, 
    277.7389, 280.8506, 289.7968, 290.9184, 287.5622, 290.0343, 288.698, 
    289.7201,
  273.4402, 273.332, 273.9945, 275.9846, 280.2321, 279.4054, 275.2039, 
    276.111, 277.7484, 281.4295, 288.8174, 283.5421, 282.4149, 288.8147, 
    288.7532,
  273.899, 273.5332, 273.3658, 273.7897, 276.5406, 274.237, 275.1461, 
    274.7285, 275.4494, 276.3775, 278.7334, 278.5443, 276.9135, 278.8646, 
    283.6092,
  274.4572, 273.6667, 272.9792, 272.9826, 273.4431, 276.2107, 273.7095, 
    275.0547, 274.3216, 274.239, 274.4819, 274.4791, 274.6179, 275.7387, 
    280.3794,
  275.1109, 273.742, 272.9169, 272.3802, 271.9664, 273.0064, 275.5161, 
    273.7761, 273.1091, 274.3734, 273.7654, 273.746, 273.8088, 273.9198, 
    275.4978,
  276.8725, 274.7108, 272.689, 272.088, 271.6681, 271.8171, 272.3686, 
    273.2455, 273.3953, 273.4096, 274.046, 273.2872, 273.435, 273.4079, 
    273.6755,
  277.4957, 276.3333, 273.0768, 271.9057, 271.4962, 271.6404, 271.5466, 
    271.9186, 271.9188, 272.2998, 272.406, 273.1212, 273.2289, 273.2085, 
    273.2613,
  277.5434, 276.5928, 274.0629, 272.087, 271.4383, 271.6776, 271.225, 
    271.6231, 271.7602, 272.2362, 272.3037, 272.8538, 273.0513, 273.0325, 
    273.2334,
  277.3312, 276.1072, 274.363, 272.3967, 271.6022, 271.4321, 271.4061, 
    271.6242, 271.6866, 272.0407, 272.4838, 272.7143, 272.7437, 272.7351, 
    273.0351,
  276.5887, 275.517, 274.0095, 273.3552, 272.5142, 271.4477, 271.4366, 
    271.5789, 271.8271, 272.1279, 271.9948, 272.1587, 272.2885, 272.3573, 
    272.8938,
  274.5247, 274.6476, 277.442, 276.2704, 277.3695, 279.6071, 277.3597, 
    277.7479, 280.804, 290.1337, 291.1661, 288.5938, 290.3933, 289.5814, 
    291.1012,
  273.5915, 274.0764, 275.4748, 275.5834, 281.6875, 280.4922, 275.5666, 
    276.8032, 278.7036, 282.7862, 289.9357, 284.561, 284.5905, 289.7946, 
    290.7503,
  273.8907, 274.2187, 275.0803, 275.6015, 280.5104, 275.2197, 275.9466, 
    275.5503, 276.8026, 278.4639, 281.9349, 281.7169, 279.3195, 280.2845, 
    285.9285,
  274.3279, 273.7446, 274.2936, 275.4389, 276.3253, 278.9213, 274.855, 
    276.8235, 275.8874, 276.1451, 277.1762, 277.4847, 276.5598, 277.5789, 
    281.908,
  274.739, 273.3783, 273.1774, 273.5917, 273.9858, 275.9106, 277.5263, 
    275.8462, 275.8873, 277.2892, 275.6602, 275.8955, 275.6228, 275.9045, 
    277.2696,
  275.2757, 273.5196, 272.6658, 272.3638, 272.8615, 273.9569, 275.6599, 
    277.0036, 279.8001, 277.1441, 276.8377, 275.314, 274.9204, 274.8157, 
    274.9974,
  276.1371, 274.1923, 272.3993, 271.8699, 272.3828, 272.9717, 273.7504, 
    274.8205, 275.6948, 274.8299, 274.9131, 274.4865, 274.3662, 274.2957, 
    274.2348,
  276.7063, 274.7953, 272.6791, 271.9428, 271.843, 272.4498, 272.6061, 
    273.5438, 274.1872, 274.1118, 274.1871, 273.8657, 273.7581, 273.6364, 
    274.0289,
  276.603, 275.1053, 273.223, 271.8369, 271.4982, 271.6743, 272.2534, 
    272.8817, 273.223, 273.3424, 273.4481, 273.3155, 273.1648, 273.0073, 
    273.4362,
  276.1302, 274.8147, 273.3179, 272.6562, 271.7615, 271.2753, 271.6653, 
    272.1588, 272.5324, 272.7141, 272.813, 272.7103, 272.6251, 272.4098, 
    272.6857,
  274.3205, 273.7538, 275.3074, 275.0832, 275.6113, 276.6422, 274.4219, 
    274.313, 275.3983, 288.9721, 290.2654, 287.6571, 288.9132, 288.2859, 
    289.0134,
  273.8648, 273.6681, 274.1505, 274.64, 277.1069, 277.4264, 274.7795, 
    274.4147, 274.9172, 280.0618, 289.2818, 284.6571, 285.0384, 288.6991, 
    289.1893,
  274.3449, 274.0681, 274.4464, 274.3987, 276.9021, 274.0747, 275.4093, 
    274.4444, 274.4677, 278.0689, 282.0342, 282.6995, 279.8193, 279.3183, 
    285.2096,
  274.857, 273.9345, 274.231, 274.6478, 275.4146, 277.8444, 274.448, 
    275.5832, 274.8846, 275.944, 277.4215, 277.3482, 276.9422, 277.7703, 
    281.9359,
  275.0547, 273.7126, 273.2216, 274.0543, 274.0929, 274.961, 277.2498, 
    274.8628, 275.0959, 277.0865, 275.7393, 276.0334, 276.1126, 275.8615, 
    277.0077,
  275.0601, 273.9559, 272.9501, 272.5718, 273.2722, 273.7809, 274.4124, 
    275.8034, 278.9718, 277.4937, 277.5245, 275.5296, 275.3726, 275.6805, 
    275.4252,
  275.8579, 274.4034, 272.6389, 272.1661, 272.6447, 273.2894, 273.9428, 
    274.4187, 275.1594, 274.926, 275.5084, 275.2621, 275.0464, 275.1752, 
    274.8623,
  276.3814, 274.6734, 272.9516, 272.1906, 272.2252, 272.6932, 273.0622, 
    273.801, 274.4569, 274.5837, 274.7257, 274.87, 274.6787, 275.0307, 
    274.9013,
  276.4386, 274.7051, 273.0668, 272.3188, 271.9469, 272.0896, 272.7482, 
    273.5523, 274.2332, 274.5147, 274.5074, 274.4529, 274.5715, 274.7471, 
    274.9001,
  276.3131, 275.0938, 273.2003, 272.641, 272.1716, 271.8417, 272.6503, 
    273.2197, 273.7603, 274.1801, 274.5378, 274.3485, 274.308, 274.1624, 
    274.7444,
  276.6397, 274.6842, 274.9878, 274.3778, 274.3826, 274.8456, 274.1597, 
    273.8038, 273.7263, 280.0927, 286.7118, 285.0305, 285.7111, 285.8818, 
    286.2967,
  274.6442, 274.1878, 274.337, 274.1039, 274.9421, 275.2175, 274.1999, 
    273.7697, 273.4861, 275.9173, 285.1715, 283.4779, 283.8561, 286.0367, 
    286.729,
  275.1971, 274.7285, 274.5112, 273.9995, 274.9564, 273.0215, 275.0164, 
    273.8958, 273.5832, 274.8429, 279.8831, 282.332, 278.7231, 277.489, 
    283.5872,
  275.7934, 274.7388, 274.0756, 274.1473, 274.4434, 276.2238, 273.4964, 
    275.031, 274.2304, 274.6784, 275.8551, 275.8321, 274.8311, 277.2173, 
    281.7436,
  275.8136, 274.2569, 273.6013, 274.1169, 273.69, 273.8812, 275.7913, 
    273.4701, 274.17, 276.0815, 274.4393, 274.4919, 274.0559, 275.5079, 
    276.6276,
  275.8491, 274.1984, 273.0703, 273.0722, 273.3139, 273.3098, 273.2905, 
    274.214, 277.3484, 277.1839, 276.3148, 274.3282, 274.0656, 274.6184, 
    274.8503,
  276.1337, 274.1661, 272.5877, 272.2791, 273.0652, 273.2964, 272.9611, 
    272.9555, 273.9397, 274.8614, 274.5004, 273.9606, 274.2551, 274.3926, 
    274.5143,
  276.286, 274.2063, 272.6055, 272.1642, 272.4835, 273.0552, 272.4721, 
    272.627, 273.5229, 274.0876, 274.1317, 274.2894, 274.3524, 274.1463, 
    273.9025,
  276.3472, 274.1661, 272.5839, 272.0308, 271.9842, 272.257, 272.1553, 
    272.7399, 273.4968, 273.9209, 273.8851, 274.2922, 274.2662, 274.333, 
    274.6259,
  276.3845, 274.6636, 272.7215, 272.1349, 272.0704, 272.0149, 272.4076, 
    272.7625, 273.3503, 273.7763, 274.1552, 274.1438, 274.085, 274.1841, 
    275.0553,
  280.228, 276.158, 277.0292, 275.0958, 274.5164, 274.5023, 273.4143, 
    273.0179, 272.7671, 275.9044, 279.1825, 282.0471, 285.2359, 286.0006, 
    286.7825,
  276.2313, 275.0549, 275.0924, 274.9356, 275.2894, 274.7659, 273.7014, 
    273.3601, 272.8995, 274.1918, 278.2304, 281.2496, 283.3365, 285.3447, 
    286.4841,
  275.697, 275.4762, 275.2044, 274.8151, 274.7785, 272.4272, 274.0489, 
    273.7095, 273.2378, 273.4424, 276.8824, 280.4738, 279.4489, 279.081, 
    283.5168,
  276.5867, 276.1032, 274.9707, 274.6646, 274.0318, 273.9138, 271.687, 
    274.2237, 273.9269, 273.8701, 273.6739, 274.6361, 275.4619, 277.9579, 
    281.5464,
  276.7172, 275.5916, 274.8883, 274.1902, 273.4985, 273.2108, 273.7038, 
    270.5483, 271.2081, 274.8319, 273.7573, 273.233, 274.6942, 276.617, 
    277.7971,
  277.0025, 275.5445, 274.5303, 273.5609, 273.117, 273.0138, 272.893, 
    273.2935, 273.692, 274.6916, 274.6134, 272.9009, 273.9519, 275.4697, 
    276.3329,
  277.0078, 275.7248, 273.9962, 273.0298, 272.9486, 273.0016, 272.6924, 
    272.67, 272.6725, 272.9532, 273.1016, 272.9278, 273.9176, 274.961, 
    275.3934,
  276.9443, 275.7437, 273.96, 272.9576, 272.7085, 272.9511, 272.7223, 
    272.3904, 272.4245, 272.8301, 272.9642, 273.0489, 273.8488, 274.5558, 
    274.8228,
  276.8228, 275.4141, 273.6183, 272.6306, 272.3048, 272.4331, 272.13, 
    272.406, 272.4653, 272.5935, 272.743, 273.0811, 273.5434, 274.2145, 
    275.0136,
  276.4318, 275.4108, 273.455, 272.4627, 272.3533, 272.0244, 272.0568, 
    272.2258, 272.4559, 273.1241, 273.1264, 273.1779, 273.4849, 273.9996, 
    275.4284,
  279.5537, 276.0513, 276.2969, 274.8032, 274.6701, 273.922, 272.9912, 
    273.0562, 273.176, 276.1557, 282.0968, 284.1177, 286.5718, 287.4813, 
    288.3843,
  276.8622, 275.3076, 275.6941, 275.5037, 275.781, 274.6056, 273.1127, 
    272.968, 272.9789, 274.2458, 280.5078, 282.6693, 283.3228, 286.632, 
    287.9527,
  276.2253, 275.6757, 275.8097, 275.6122, 275.8538, 272.26, 273.5135, 
    273.2714, 272.9943, 273.0518, 276.7778, 281.1913, 280.1033, 277.847, 
    283.507,
  276.6218, 276.1058, 275.6357, 275.61, 275.1893, 275.0056, 271.4959, 
    273.3204, 273.1355, 272.7706, 272.9976, 274.1657, 274.9229, 276.6784, 
    281.2416,
  276.9516, 275.9608, 275.5649, 275.1663, 274.619, 274.3671, 274.0111, 
    270.5891, 269.8162, 273.0264, 272.7892, 272.8417, 274.1772, 275.6644, 
    277.481,
  277.4215, 276.1537, 275.0679, 274.1702, 273.8027, 273.7726, 273.5369, 
    273.6893, 273.4607, 273.2122, 273.0724, 272.5325, 273.2957, 274.4413, 
    276.46,
  277.4268, 276.4431, 274.6637, 273.7454, 273.6943, 273.5764, 273.4876, 
    273.0287, 272.8712, 272.6483, 272.4188, 272.4343, 272.8736, 273.8675, 
    274.9314,
  277.1195, 276.2268, 274.5916, 273.718, 273.4853, 273.5304, 273.2634, 
    272.9736, 272.8828, 272.8166, 272.7474, 272.316, 272.6747, 273.402, 
    274.1528,
  276.2785, 275.4886, 274.0085, 273.421, 273.033, 273.0237, 272.8621, 
    272.8593, 273.0274, 272.9126, 272.7047, 272.2067, 272.4683, 273.1915, 
    274.202,
  275.8112, 275.1741, 273.9519, 273.3559, 273.1006, 272.6771, 272.6371, 
    272.838, 272.9285, 273.3214, 273.1114, 272.627, 272.4125, 273.1073, 
    274.6804 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;
}
