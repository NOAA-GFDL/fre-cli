netcdf atmos.1980-1981.alb_sfc.12 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:23 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.12.nc reduced/atmos.1980-1981.alb_sfc.12.nc\n",
			"Mon Aug 25 14:40:10 2025: cdo -O -s -select,month=12 merged_output.nc monthly_nc_files/all_years.12.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.10503, 76.10503, 76.10503, 76.10503, 76.10503, 76.10503, 76.10503, 
    76.08111, 76.08111, 76.08111, 76.08111, 76.08111, 76.08111, 76.08111, 
    76.0997, 76.0997, 76.0997, 76.0997, 76.0997, 76.0997, 76.0997, 76.11059, 
    76.11059, 76.11059, 76.11059, 76.11059, 76.11059, 76.11059, 76.10503,
  76.29614, 76.13136, 76.03885, 75.97415, 75.9507, 75.93606, 75.91145, 
    75.90384, 75.93697, 75.98314, 76.04004, 76.10185, 76.27303, 72.07031, 
    68.58884, 66.67876, 66.96962, 67.45403, 70.4799, 75.24809, 76.15636, 
    76.26704, 75.9642, 64.96976, 65.49171, 65.04669, 64.58506, 67.4993, 
    76.20941,
  46.87786, 39.96181, 64.39506, 66.27346, 75.86948, 76.18105, 55.03302, 
    76.14375, 75.89551, 75.77046, 75.85233, 75.91716, 72.28996, 70.72544, 
    59.35869, 46.08599, 42.78984, 61.48574, 57.78291, 61.92829, 56.04182, 
    46.98893, 62.13132, 63.71282, 63.57416, 61.41718, 45.91488, 50.13792, 
    55.66421,
  16.8133, 34.53127, 5.053813, 4.734261, 4.741735, 4.7216, 4.783731, 
    5.019849, 4.97082, 5.30272, 5.147202, 5.179983, 4.922304, 5.11463, 
    5.306605, 5.13544, 5.120944, 4.962682, 5.105036, 5.13433, 5.21972, 
    5.145105, 5.113221, 5.048722, 4.954862, 6.7939, 19.08561, 8.806641, 
    11.69949,
  4.279478, 4.443476, 4.287549, 4.443133, 4.395266, 4.343117, 4.45609, 
    4.392529, 4.348963, 4.415463, 4.569802, 4.435055, 4.449807, 4.427995, 
    4.543892, 4.518588, 4.367543, 4.524535, 4.392963, 4.63823, 4.468861, 
    4.473319, 4.473026, 8.907784, 5.150207, 4.617364, 4.425183, 4.311183, 
    4.342497,
  4.145757, 4.185833, 4.476629, 4.085831, 4.147009, 4.239552, 3.88379, 
    4.097924, 4.027151, 3.992097, 3.968961, 4.405072, 4.177349, 4.096833, 
    10.35499, 3.909516, 4.111835, 4.151862, 3.89616, 3.9253, 4.10831, 
    3.988275, 4.193695, 10.26426, 4.357756, 4.308887, 4.130498, 4.078637, 
    4.131315,
  3.802169, 4.166976, 13.13002, 3.700326, 3.919766, 4.071618, 3.718789, 
    4.005287, 3.860485, 4.156734, 10.4353, 16.16739, 10.9104, 4.065786, 
    3.951375, 3.790089, 4.054991, 3.733757, 3.501981, 3.711369, 4.074963, 
    3.999663, 3.962647, 4.880327, 9.682905, 3.896729, 3.785658, 3.857471, 
    3.856325,
  3.5819, 10.21433, 10.37079, 3.853421, 3.618266, 3.569721, 3.943085, 
    3.840947, 3.732431, 4.077193, 12.39938, 11.70889, 3.91102, 3.69136, 
    3.517444, 3.656796, 3.548066, 3.582819, 3.869015, 4.104854, 3.915275, 
    3.968794, 3.35065, 3.369767, 9.677103, 9.295023, 3.879828, 4.002501, 
    3.778033,
  3.283251, 6.729254, 8.97518, 9.309628, 3.391373, 3.468206, 3.432476, 
    3.41042, 3.64651, 3.323582, 4.918044, 3.414434, 4.531486, 3.515946, 
    3.478162, 3.662994, 3.553897, 3.859062, 3.635423, 3.985516, 3.735286, 
    3.714665, 3.370463, 8.979336, 8.593068, 9.004148, 3.942736, 3.602668, 
    3.73012,
  3.197361, 8.865829, 8.456902, 9.776688, 3.494531, 3.456484, 3.393553, 
    3.332913, 8.589512, 8.200069, 3.398462, 3.435102, 3.242892, 3.514468, 
    3.553082, 3.702202, 3.797708, 3.942632, 3.796981, 3.907762, 3.735628, 
    3.274373, 3.407699, 8.49506, 8.531149, 3.42116, 3.320045, 3.480578, 
    3.324142,
  10.11051, 10.34214, 10.31748, 9.427639, 14.11427, 3.485023, 5.617156, 
    3.862507, 3.442932, 3.518115, 4.111053, 3.377853, 3.455878, 3.545969, 
    3.406113, 3.495192, 3.777352, 3.279346, 3.604388, 3.329583, 3.361903, 
    3.549294, 8.49311, 7.21569, 3.516026, 3.676444, 3.156696, 3.611843, 
    9.082184,
  15.77451, 18.44079, 20.69578, 3.746661, 20.38319, 3.959573, 10.35046, 
    4.036091, 9.113181, 3.313825, 3.413391, 3.845028, 3.867935, 4.023733, 
    4.230939, 3.833264, 3.991562, 3.731984, 3.538241, 3.414243, 4.010314, 
    5.919721, 3.958119, 4.880523, 3.864221, 4.121014, 3.815927, 3.720226, 
    20.94269,
  20.05619, 16.51525, 17.01379, 16.10738, 10.76033, 12.31952, 11.08919, 
    21.27963, 13.78068, 9.569291, 3.448311, 3.771718, 4.110298, 3.894118, 
    3.717038, 3.743931, 3.651792, 3.89443, 3.63577, 3.887563, 8.502436, 
    10.1821, 8.058939, 3.561425, 3.862529, 3.696899, 4.047906, 3.937255, 
    9.66197,
  5.410643, 4.310389, 5.207832, 11.44706, 1.528826, 11.08989, 16.58542, 
    12.41909, 10.18968, 16.18176, 8.729153, 3.517613, 4.027048, 3.913574, 
    3.721427, 3.664709, 3.139412, 3.21302, 3.732711, 11.0225, 16.29063, 
    11.90427, 10.3259, 3.948894, 3.535845, 3.455247, 3.610365, 3.889568, 
    4.483768,
  4.025896, 7.95948, 11.29212, 15.24515, 13.80349, 16.54919, 9.917079, 
    24.06674, 12.42013, 6.424431, 8.225542, 13.37249, 3.493358, 3.886976, 
    3.788833, 3.28882, 3.47141, 3.444024, 3.784104, 11.80795, 12.13999, 
    17.39129, 12.57756, 20.22474, 5.366607, 3.385702, 3.327144, 3.428303, 
    3.309577,
  2.447707, 12.10244, 6.671196, 11.0071, 8.393936, 9.591779, 10.09949, 
    12.54754, 11.49754, 10.72755, 8.483713, 17.87166, 18.41294, 12.76131, 
    2.227526, 3.398121, 14.95881, 7.966526, 18.06502, 9.093077, 11.4062, 
    18.63674, 20.60293, 18.45658, 2.193076, 5.483738, 2.621521, 2.602271, 
    2.465904,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 average_DT = 730 ;

 average_T1 = 350.5 ;

 average_T2 = 1080.5 ;

 climatology_bounds =
  350.5, 1080.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
