netcdf atmos_tracer.pk {
dimensions:
	phalf = 50 ;
variables:
	double phalf(phalf) ;
		phalf:long_name = "ref half pressure level" ;
		phalf:units = "mb" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float pk(phalf) ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:units = "pascal" ;
		pk:missing_value = 1.e+20f ;
		pk:_FillValue = 1.e+20f ;
		pk:cell_methods = "time: point" ;

// global attributes:
		:filename = "00080101.atmos_tracer.tile1.nc" ;
		:title = "ESM4_piClim-NTCF" ;
		:associated_files = "area: 00080101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "19.1" ;
		:git_hash = "5a324f5f5c98dbb620b25cd98a6add9da8861ee5" ;
		:creationtime = "Mon Jun  6 22:26:34 2022" ;
		:hostname = "pp212" ;
		:history = "fregrid --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /xtmp/Luis.Sal-bey/ptmp/archive/oar.gfdl.bgrp-account/CMIP6/ESM4/AerChemMIP/ESM4_piClim-NTCF/gfdl.ncrc4-intel16-prod-openmp/history/00080101.nc --input_file 00080101.atmos_tracer --associated_file_dir /xtmp/Luis.Sal-bey/ptmp/archive/oar.gfdl.bgrp-account/CMIP6/ESM4/AerChemMIP/ESM4_piClim-NTCF/gfdl.ncrc4-intel16-prod-openmp/history/00080101.nc --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 00080101.atmos_tracer.nc" ;
data:

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;
}
