netcdf atmos.1980-1981.alb_sfc.02 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:16 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.02.nc reduced/atmos.1980-1981.alb_sfc.02.nc\n",
			"Mon Aug 25 14:40:03 2025: cdo -O -s -select,month=2 merged_output.nc monthly_nc_files/all_years.2.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  76.46632, 76.46632, 76.46632, 76.46632, 76.46632, 76.46632, 76.46632, 
    76.45107, 76.45107, 76.45107, 76.45107, 76.45107, 76.45107, 76.45107, 
    76.44231, 76.44231, 76.44231, 76.44231, 76.44231, 76.44231, 76.44231, 
    76.48018, 76.48018, 76.48018, 76.48018, 76.48018, 76.48018, 76.48018, 
    76.46632,
  73.33899, 73.05287, 72.96189, 73.0626, 72.84399, 72.94429, 72.894, 
    72.85896, 72.99685, 73.07772, 72.84206, 73.23705, 73.32324, 73.65193, 
    73.87918, 73.10371, 73.99498, 72.97849, 73.37125, 73.87116, 74.08426, 
    74.15184, 74.03844, 73.73395, 74.62515, 72.12745, 73.58112, 73.47295, 
    73.48403,
  29.96032, 29.15553, 7.876028, 47.24438, 55.84823, 55.81261, 42.92263, 
    55.7578, 55.84989, 56.08478, 55.68092, 55.5647, 55.35736, 23.60406, 
    5.641232, 5.47156, 5.572774, 5.154702, 5.114913, 9.704969, 17.25746, 
    15.24052, 45.39765, 47.7708, 47.69857, 26.88602, 5.29225, 5.234877, 
    5.939528,
  4.473701, 4.453276, 4.510859, 4.304663, 4.188403, 4.319375, 4.266176, 
    4.428085, 4.343897, 4.392703, 4.449575, 4.238505, 4.21286, 4.349861, 
    4.469809, 4.42102, 4.418945, 4.262979, 4.571476, 4.612138, 4.687686, 
    4.838447, 4.72905, 4.508259, 4.301525, 4.193824, 4.227023, 4.453783, 
    4.228896,
  4.023607, 3.954847, 3.970927, 4.019078, 4.06574, 4.042761, 3.945273, 
    4.098862, 4.089128, 4.082009, 4.085841, 4.054593, 4.048558, 4.085129, 
    4.080842, 3.924925, 3.995923, 3.896473, 4.07529, 4.063331, 4.304502, 
    4.104668, 4.207853, 7.891032, 4.54668, 4.271481, 4.038647, 4.055033, 
    3.819686,
  3.884533, 3.903846, 4.016439, 3.932561, 3.855958, 3.804621, 3.837975, 
    3.730464, 3.706554, 3.805989, 3.862039, 3.942483, 4.068407, 4.034425, 
    9.37828, 3.693163, 3.78522, 3.756308, 3.733602, 3.834393, 3.84114, 
    3.903701, 3.887255, 9.524237, 4.391875, 3.902371, 3.77731, 3.903416, 
    3.850276,
  3.878907, 4.175944, 11.95327, 3.890288, 3.726914, 3.568894, 3.939737, 
    3.771306, 3.826954, 3.914807, 9.765942, 14.66128, 10.35228, 3.71568, 
    3.651808, 3.748831, 3.55729, 3.544552, 3.50926, 3.754583, 3.83422, 
    3.96126, 3.71527, 4.206433, 9.428144, 3.438399, 3.792581, 3.787236, 
    4.089929,
  3.444427, 9.729572, 12.29994, 3.553975, 3.339023, 3.548722, 3.780568, 
    3.51337, 3.76131, 3.326385, 11.97927, 11.42973, 3.660969, 3.631499, 
    3.500576, 3.581405, 3.339772, 3.589286, 3.398526, 3.753402, 3.783792, 
    3.724665, 3.455577, 3.34839, 8.934858, 9.028818, 3.94543, 3.644099, 
    3.941237,
  3.321854, 6.36914, 8.458448, 9.155956, 3.347723, 3.238166, 3.569285, 
    3.372907, 3.303072, 3.233337, 4.50501, 3.140845, 4.320949, 3.197199, 
    3.155785, 3.572142, 3.423911, 3.521122, 3.531282, 3.813221, 3.539169, 
    3.835636, 3.423729, 8.32793, 8.435966, 8.834289, 3.520561, 3.538316, 
    3.755793,
  3.141441, 8.717727, 8.554625, 9.82284, 3.29614, 3.276848, 3.264101, 
    3.215625, 8.580481, 8.357949, 3.252137, 3.286335, 3.27492, 3.223899, 
    3.337106, 3.581286, 3.590884, 3.718259, 3.59503, 3.729609, 3.61101, 
    3.441164, 3.380523, 8.561865, 8.424257, 3.190678, 3.273814, 3.338884, 
    3.079715,
  9.946072, 10.1841, 10.84509, 9.350763, 14.29078, 3.501082, 5.316605, 
    3.571685, 3.77299, 3.446354, 3.980907, 3.464666, 3.205643, 3.35924, 
    3.559324, 3.386349, 3.55551, 3.53932, 3.451666, 3.287234, 3.430692, 
    3.394828, 8.533057, 7.632155, 3.325669, 3.466795, 3.173639, 3.28495, 
    8.979387,
  17.10796, 19.21441, 20.93988, 3.791083, 21.15709, 3.784735, 10.61384, 
    4.129487, 9.187893, 3.441311, 3.353195, 3.608513, 3.775432, 3.719488, 
    3.670495, 3.840092, 3.856375, 3.580884, 3.795105, 3.375807, 3.884954, 
    6.25952, 3.752212, 4.423144, 3.876687, 3.979011, 3.586429, 3.794988, 
    21.72717,
  21.32569, 16.66859, 17.84926, 17.25238, 11.9016, 13.44965, 12.30154, 
    25.51046, 9.955756, 10.62229, 3.280421, 3.656871, 3.781995, 3.80209, 
    3.762144, 3.512916, 3.766914, 3.442153, 3.675212, 3.957345, 11.9109, 
    12.36869, 12.25038, 3.561423, 3.706083, 3.826117, 3.761753, 3.793973, 
    10.19964,
  5.930854, 4.240141, 6.100352, 15.3324, 1.74908, 12.93776, 26.6163, 13.2911, 
    11.39474, 22.574, 9.517224, 3.666838, 3.59494, 3.841318, 3.884871, 
    3.753674, 3.306147, 3.470819, 3.76785, 11.4113, 26.02317, 18.61465, 
    19.25358, 4.699409, 3.402245, 3.452131, 3.533766, 3.722349, 4.799566,
  5.166562, 13.52938, 13.55248, 26.79116, 28.87493, 30.70369, 15.66949, 
    30.2417, 13.75195, 6.557472, 8.445839, 21.1758, 16.50112, 3.595986, 
    3.548397, 3.911432, 3.840993, 3.949238, 3.898877, 24.27809, 20.06975, 
    27.47622, 23.19306, 27.156, 12.59693, 3.484642, 3.845275, 3.871078, 
    3.830226,
  3.852965, 18.41452, 17.14652, 21.02898, 21.17858, 21.51122, 22.46184, 
    23.0162, 19.29049, 19.38416, 16.94293, 28.43177, 29.43278, 25.36406, 
    3.241355, 33.22471, 25.70556, 13.08142, 28.87255, 19.24388, 21.24431, 
    29.40742, 35.13428, 29.37322, 2.80198, 8.250795, 4.159647, 3.789786, 
    3.909448,
  3.054792, 2.94289, 14.87201, 2.484436, 13.20413, 25.8596, 22.16542, 
    22.18013, 21.86697, 21.71097, 14.80493, 12.79802, 21.76153, 26.20354, 
    25.96832, 26.68803, 23.74459, 23.90157, 25.76686, 25.88697, 22.02232, 
    24.59022, 22.82656, 22.61774, 26.60117, 22.47441, 22.54611, 24.55324, 
    3.044761,
  2.354074, 2.256808, 2.497179, 2.529313, 2.337799, 2.206168, 2.415388, 
    2.384713, 2.369056, 2.239275, 2.202894, 2.14653, 2.283909, 2.499045, 
    2.481931, 2.425821, 2.506456, 2.739497, 2.886353, 2.665874, 2.746998, 
    2.534967, 2.275367, 2.506107, 2.199348, 2.269395, 2.075997, 2.180186, 
    2.598958 ;

 average_DT = 731 ;

 average_T1 = 45 ;

 average_T2 = 776 ;

 climatology_bounds =
  45, 776 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
