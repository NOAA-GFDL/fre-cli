netcdf \20030101.grid_spec.tile6 {
dimensions:
	grid_x = 97 ;
	grid_y = 97 ;
	time = UNLIMITED ; // (1 currently)
	grid_xt = 96 ;
	grid_yt = 96 ;
	phalf = 50 ;
variables:
	double grid_x(grid_x) ;
		grid_x:units = "degrees_E" ;
		grid_x:long_name = "cell corner longitude" ;
		grid_x:axis = "X" ;
	double grid_y(grid_y) ;
		grid_y:units = "degrees_N" ;
		grid_y:long_name = "cell corner latitude" ;
		grid_y:axis = "Y" ;
	double time(time) ;
		time:units = "days since 1870-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "JULIAN" ;
		time:calendar = "julian" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	float grid_lon(grid_y, grid_x) ;
		grid_lon:_FillValue = 1.e+20f ;
		grid_lon:missing_value = 1.e+20f ;
		grid_lon:units = "degrees_E" ;
		grid_lon:long_name = "longitude" ;
		grid_lon:cell_methods = "time: point" ;
	float grid_lat(grid_y, grid_x) ;
		grid_lat:_FillValue = 1.e+20f ;
		grid_lat:missing_value = 1.e+20f ;
		grid_lat:units = "degrees_N" ;
		grid_lat:long_name = "latitude" ;
		grid_lat:cell_methods = "time: point" ;
	float grid_lont(grid_yt, grid_xt) ;
		grid_lont:_FillValue = 1.e+20f ;
		grid_lont:missing_value = 1.e+20f ;
		grid_lont:units = "degrees_E" ;
		grid_lont:long_name = "longitude" ;
		grid_lont:cell_methods = "time: point" ;
	float grid_latt(grid_yt, grid_xt) ;
		grid_latt:_FillValue = 1.e+20f ;
		grid_latt:missing_value = 1.e+20f ;
		grid_latt:units = "degrees_N" ;
		grid_latt:long_name = "latitude" ;
		grid_latt:cell_methods = "time: point" ;
	float area(grid_yt, grid_xt) ;
		area:_FillValue = 1.e+20f ;
		area:missing_value = 1.e+20f ;
		area:units = "m**2" ;
		area:long_name = "cell area" ;
		area:cell_methods = "time: point" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	float orog(grid_yt, grid_xt) ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:units = "m" ;
		orog:long_name = "Surface Altitude" ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:standard_name = "surface_altitude" ;
		orog:interp_method = "conserve_order1" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;

// global attributes:
		:title = "ESM4_longamip_D1_am4p2_proto7b_whiteCapsAlbedo_salt_SIS2" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
data:

 grid_x = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 grid_y = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97 ;

 time = 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96 ;

 phalf = 0.01, 0.0269722, 0.0517136, 0.0889455, 0.142479, 0.2207157, 
    0.3361283, 0.5048096, 0.7479993, 1.0940055, 1.580046, 2.2544108, 
    3.178956, 4.431935, 6.1111558, 8.3374392, 11.2583405, 15.0520759, 
    19.9315829, 26.1486254, 33.997842, 43.820624, 56.0087014, 71.0073115, 
    89.3178242, 111.4997021, 138.1716841, 170.012093, 207.7581856, 
    252.2033875, 304.1464563, 363.9522552, 430.6429622, 501.015122, 
    570.6113482, 635.806353, 694.8286462, 747.1992533, 793.0044191, 
    832.5750255, 866.4443202, 895.1917865, 919.4060705, 939.6860264, 
    956.4664631, 970.1833931, 981.1347983, 989.68, 995.9, 1000 ;

 grid_lon =
  215, 214.2172, 213.4273, 212.6302, 211.8259, 211.0143, 210.1953, 209.3691, 
    208.5354, 207.6944, 206.8459, 205.99, 205.1267, 204.256, 203.3779, 
    202.4925, 201.5998, 200.6998, 199.7926, 198.8784, 197.957, 197.0288, 
    196.0937, 195.1518, 194.2034, 193.2486, 192.2874, 191.3201, 190.3468, 
    189.3678, 188.3832, 187.3932, 186.3981, 185.3981, 184.3935, 183.3844, 
    182.3713, 181.3542, 180.3337, 179.3098, 178.283, 177.2535, 176.2217, 
    175.1878, 174.1523, 173.1154, 172.0775, 171.0389, 170, 168.9611, 
    167.9225, 166.8846, 165.8477, 164.8122, 163.7783, 162.7465, 161.717, 
    160.6902, 159.6663, 158.6458, 157.6287, 156.6156, 155.6065, 154.6019, 
    153.6019, 152.6068, 151.6168, 150.6322, 149.6532, 148.6799, 147.7126, 
    146.7514, 145.7966, 144.8482, 143.9063, 142.9712, 142.043, 141.1216, 
    140.2074, 139.3002, 138.4002, 137.5075, 136.6221, 135.744, 134.8733, 
    134.01, 133.1541, 132.3056, 131.4646, 130.6309, 129.8047, 128.9857, 
    128.1741, 127.3698, 126.5727, 125.7828, 125,
  215.7828, 215, 214.2095, 213.4112, 212.605, 211.791, 210.9689, 210.1388, 
    209.3007, 208.4544, 207.6001, 206.7375, 205.8669, 204.9881, 204.1011, 
    203.206, 202.3028, 201.3916, 200.4724, 199.5453, 198.6104, 197.6677, 
    196.7173, 195.7595, 194.7942, 193.8217, 192.8422, 191.8557, 190.8626, 
    189.8629, 188.8569, 187.8449, 186.8271, 185.8037, 184.775, 183.7414, 
    182.703, 181.6603, 180.6135, 179.563, 178.5091, 177.4522, 176.3926, 
    175.3307, 174.2669, 173.2016, 172.135, 171.0677, 170, 168.9323, 167.865, 
    166.7984, 165.7331, 164.6693, 163.6074, 162.5478, 161.4909, 160.437, 
    159.3865, 158.3397, 157.297, 156.2586, 155.225, 154.1963, 153.1729, 
    152.1551, 151.1431, 150.1371, 149.1374, 148.1443, 147.1578, 146.1783, 
    145.2058, 144.2405, 143.2827, 142.3323, 141.3896, 140.4547, 139.5276, 
    138.6084, 137.6972, 136.794, 135.8989, 135.0119, 134.1331, 133.2625, 
    132.3999, 131.5456, 130.6993, 129.8612, 129.0311, 128.209, 127.395, 
    126.5888, 125.7905, 125, 124.2172,
  216.5727, 215.7905, 215, 214.2011, 213.3937, 212.5777, 211.7531, 210.9198, 
    210.0777, 209.2268, 208.3671, 207.4984, 206.6208, 205.7343, 204.8389, 
    203.9345, 203.0212, 202.0991, 201.1681, 200.2284, 199.28, 198.323, 
    197.3575, 196.3837, 195.4016, 194.4114, 193.4133, 192.4075, 191.3942, 
    190.3736, 189.3458, 188.3113, 187.2702, 186.2229, 185.1696, 184.1107, 
    183.0465, 181.9773, 180.9035, 179.8255, 178.7436, 177.6583, 176.57, 
    175.479, 174.3859, 173.291, 172.1947, 171.0976, 170, 168.9024, 167.8053, 
    166.709, 165.6141, 164.521, 163.43, 162.3417, 161.2564, 160.1745, 
    159.0965, 158.0227, 156.9535, 155.8893, 154.8304, 153.7771, 152.7298, 
    151.6887, 150.6542, 149.6264, 148.6058, 147.5925, 146.5867, 145.5886, 
    144.5984, 143.6163, 142.6425, 141.677, 140.72, 139.7716, 138.8319, 
    137.9009, 136.9788, 136.0655, 135.1611, 134.2657, 133.3792, 132.5016, 
    131.6329, 130.7732, 129.9223, 129.0802, 128.2469, 127.4223, 126.6063, 
    125.7989, 125, 124.2095, 123.4273,
  217.3698, 216.5888, 215.7989, 215, 214.192, 213.3747, 212.5482, 211.7122, 
    210.8667, 210.0117, 209.1471, 208.2729, 207.3889, 206.4951, 205.5917, 
    204.6784, 203.7555, 202.8227, 201.8803, 200.9283, 199.9666, 198.9955, 
    198.015, 197.0252, 196.0262, 195.0183, 194.0016, 192.9762, 191.9425, 
    190.9006, 189.8508, 188.7933, 187.7285, 186.6567, 185.5781, 184.4932, 
    183.4023, 182.3059, 181.2042, 180.0977, 178.9869, 177.8722, 176.7541, 
    175.633, 174.5094, 173.3838, 172.2567, 171.1286, 170, 168.8714, 167.7433, 
    166.6162, 165.4906, 164.367, 163.2459, 162.1278, 161.0131, 159.9023, 
    158.7958, 157.6941, 156.5977, 155.5068, 154.4219, 153.3433, 152.2715, 
    151.2067, 150.1492, 149.0994, 148.0575, 147.0238, 145.9984, 144.9817, 
    143.9738, 142.9748, 141.985, 141.0045, 140.0334, 139.0717, 138.1197, 
    137.1773, 136.2445, 135.3216, 134.4083, 133.5049, 132.6111, 131.7271, 
    130.8529, 129.9883, 129.1333, 128.2878, 127.4518, 126.6253, 125.808, 125, 
    124.2011, 123.4112, 122.6302,
  218.1741, 217.395, 216.6063, 215.808, 215, 214.1821, 213.3542, 212.5162, 
    211.668, 210.8095, 209.9406, 209.0613, 208.1714, 207.271, 206.36, 
    205.4384, 204.5061, 203.5632, 202.6096, 201.6455, 200.6709, 199.6858, 
    198.6904, 197.6848, 196.669, 195.6433, 194.6078, 193.5628, 192.5084, 
    191.4449, 190.3726, 189.2918, 188.2027, 187.1058, 186.0013, 184.8897, 
    183.7714, 182.6468, 181.5163, 180.3804, 179.2397, 178.0945, 176.9455, 
    175.7931, 174.6379, 173.4804, 172.3212, 171.1609, 170, 168.8391, 
    167.6788, 166.5196, 165.3621, 164.2069, 163.0545, 161.9055, 160.7603, 
    159.6196, 158.4837, 157.3532, 156.2286, 155.1103, 153.9987, 152.8942, 
    151.7973, 150.7082, 149.6274, 148.5551, 147.4916, 146.4372, 145.3922, 
    144.3567, 143.331, 142.3152, 141.3096, 140.3142, 139.3291, 138.3545, 
    137.3904, 136.4368, 135.4939, 134.5616, 133.64, 132.729, 131.8286, 
    130.9387, 130.0594, 129.1905, 128.332, 127.4838, 126.6458, 125.8179, 125, 
    124.192, 123.3937, 122.605, 121.8259,
  218.9857, 218.209, 217.4223, 216.6253, 215.8179, 215, 214.1714, 213.332, 
    212.4817, 211.6204, 210.7478, 209.864, 208.9689, 208.0624, 207.1443, 
    206.2148, 205.2737, 204.321, 203.3567, 202.3809, 201.3936, 200.3948, 
    199.3847, 198.3633, 197.3308, 196.2873, 195.233, 194.1681, 193.0928, 
    192.0075, 190.9123, 189.8076, 188.6938, 187.5711, 186.4401, 185.301, 
    184.1545, 183.0008, 181.8406, 180.6743, 179.5025, 178.3257, 177.1446, 
    175.9597, 174.7716, 173.5809, 172.3884, 171.1945, 170, 168.8055, 
    167.6116, 166.4191, 165.2284, 164.0403, 162.8554, 161.6743, 160.4975, 
    159.3257, 158.1594, 156.9992, 155.8455, 154.699, 153.5599, 152.4289, 
    151.3062, 150.1924, 149.0877, 147.9925, 146.9072, 145.8319, 144.767, 
    143.7127, 142.6692, 141.6367, 140.6153, 139.6052, 138.6064, 137.6191, 
    136.6433, 135.679, 134.7263, 133.7852, 132.8557, 131.9376, 131.0311, 
    130.136, 129.2522, 128.3796, 127.5183, 126.668, 125.8286, 125, 124.1821, 
    123.3747, 122.5777, 121.791, 121.0143,
  219.8047, 219.0311, 218.2469, 217.4518, 216.6458, 215.8286, 215, 214.1599, 
    213.3082, 212.4446, 211.5691, 210.6815, 209.7817, 208.8696, 207.9451, 
    207.0082, 206.0587, 205.0967, 204.1222, 203.135, 202.1354, 201.1232, 
    200.0985, 199.0616, 198.0124, 196.9511, 195.878, 194.7931, 193.6968, 
    192.5893, 191.4709, 190.3419, 189.2028, 188.0538, 186.8955, 185.7282, 
    184.5525, 183.3689, 182.1779, 180.9801, 179.7761, 178.5665, 177.352, 
    176.1333, 174.911, 173.6858, 172.4584, 171.2296, 170, 168.7704, 167.5416, 
    166.3142, 165.089, 163.8667, 162.648, 161.4335, 160.2239, 159.0199, 
    157.8221, 156.6311, 155.4475, 154.2718, 153.1045, 151.9462, 150.7972, 
    149.6581, 148.5291, 147.4107, 146.3032, 145.2069, 144.122, 143.0489, 
    141.9876, 140.9384, 139.9015, 138.8768, 137.8646, 136.865, 135.8778, 
    134.9033, 133.9413, 132.9918, 132.0549, 131.1304, 130.2183, 129.3185, 
    128.4309, 127.5554, 126.6918, 125.8401, 125, 124.1714, 123.3542, 
    122.5482, 121.7531, 120.9689, 120.1954,
  220.6309, 219.8612, 219.0802, 218.2878, 217.4838, 216.668, 215.8401, 215, 
    214.1475, 213.2824, 212.4046, 211.5139, 210.61, 209.6931, 208.7628, 
    207.8191, 206.8618, 205.8911, 204.9067, 203.9087, 202.897, 201.8717, 
    200.8329, 199.7805, 198.7148, 197.6359, 196.5438, 195.4389, 194.3213, 
    193.1914, 192.0494, 190.8958, 189.7307, 188.5548, 187.3685, 186.1722, 
    184.9664, 183.7519, 182.529, 181.2986, 180.0612, 178.8175, 177.5684, 
    176.3144, 175.0564, 173.7952, 172.5315, 171.2661, 170, 168.7339, 
    167.4685, 166.2048, 164.9436, 163.6856, 162.4316, 161.1825, 159.9388, 
    158.7014, 157.471, 156.2481, 155.0336, 153.8278, 152.6315, 151.4452, 
    150.2693, 149.1042, 147.9506, 146.8086, 145.6787, 144.5611, 143.4562, 
    142.3641, 141.2852, 140.2195, 139.1671, 138.1283, 137.103, 136.0913, 
    135.0933, 134.1089, 133.1382, 132.1809, 131.2372, 130.3069, 129.39, 
    128.4861, 127.5954, 126.7176, 125.8525, 125, 124.1599, 123.332, 122.5162, 
    121.7122, 120.9198, 120.1388, 119.3691,
  221.4646, 220.6993, 219.9223, 219.1333, 218.332, 217.5183, 216.6918, 
    215.8525, 215, 214.1342, 213.2547, 212.3616, 211.4545, 210.5333, 
    209.5978, 208.648, 207.6836, 206.7046, 205.711, 204.7025, 203.6793, 
    202.6413, 201.5886, 200.5211, 199.4391, 198.3425, 197.2316, 196.1066, 
    194.9676, 193.815, 192.6491, 191.4703, 190.2789, 189.0754, 187.8603, 
    186.6341, 185.3974, 184.1508, 182.8951, 181.6307, 180.3586, 179.0795, 
    177.7942, 176.5035, 175.2083, 173.9094, 172.6078, 171.3044, 170, 
    168.6956, 167.3922, 166.0906, 164.7917, 163.4965, 162.2058, 160.9205, 
    159.6414, 158.3693, 157.1049, 155.8492, 154.6026, 153.3659, 152.1397, 
    150.9246, 149.7211, 148.5297, 147.3509, 146.185, 145.0324, 143.8934, 
    142.7684, 141.6575, 140.5609, 139.4789, 138.4114, 137.3587, 136.3207, 
    135.2975, 134.289, 133.2954, 132.3164, 131.352, 130.4022, 129.4667, 
    128.5455, 127.6384, 126.7453, 125.8659, 125, 124.1475, 123.3082, 
    122.4817, 121.668, 120.8667, 120.0777, 119.3007, 118.5354,
  222.3056, 221.5456, 220.7732, 219.9883, 219.1905, 218.3796, 217.5554, 
    216.7176, 215.8658, 215, 214.1198, 213.225, 212.3153, 211.3906, 210.4507, 
    209.4955, 208.5246, 207.538, 206.5357, 205.5174, 204.4831, 203.4329, 
    202.3666, 201.2843, 200.1862, 199.0721, 197.9424, 196.7972, 195.6368, 
    194.4613, 193.2712, 192.0667, 190.8484, 189.6167, 188.3721, 187.1152, 
    185.8465, 184.5669, 183.277, 181.9775, 180.6694, 179.3533, 178.0303, 
    176.7013, 175.3672, 174.029, 172.6877, 171.3444, 170, 168.6556, 167.3123, 
    165.971, 164.6328, 163.2987, 161.9697, 160.6467, 159.3306, 158.0225, 
    156.723, 155.4331, 154.1535, 152.8848, 151.6279, 150.3833, 149.1516, 
    147.9333, 146.7288, 145.5387, 144.3632, 143.2028, 142.0576, 140.9279, 
    139.8138, 138.7157, 137.6334, 136.5671, 135.5169, 134.4826, 133.4643, 
    132.462, 131.4754, 130.5045, 129.5493, 128.6094, 127.6847, 126.775, 
    125.8802, 125, 124.1341, 123.2824, 122.4446, 121.6204, 120.8095, 
    120.0117, 119.2268, 118.4544, 117.6944,
  223.1541, 222.3999, 221.6329, 220.8529, 220.0594, 219.2522, 218.4309, 
    217.5954, 216.7453, 215.8802, 215, 214.1043, 213.1929, 212.2656, 211.322, 
    210.362, 209.3854, 208.392, 207.3815, 206.354, 205.3093, 204.2473, 
    203.1679, 202.0712, 200.9572, 199.8259, 198.6775, 197.5122, 196.3302, 
    195.1316, 193.917, 192.6865, 191.4408, 190.1802, 188.9053, 187.6167, 
    186.3151, 185.0013, 183.676, 182.34, 180.9943, 179.6398, 178.2775, 
    176.9085, 175.5337, 174.1543, 172.7715, 171.3863, 170, 168.6137, 
    167.2285, 165.8457, 164.4663, 163.0915, 161.7225, 160.3602, 159.0057, 
    157.66, 156.324, 154.9987, 153.6849, 152.3833, 151.0947, 149.8198, 
    148.5592, 147.3135, 146.083, 144.8684, 143.6698, 142.4878, 141.3225, 
    140.1741, 139.0428, 137.9288, 136.8321, 135.7527, 134.6907, 133.646, 
    132.6185, 131.608, 130.6146, 129.638, 128.678, 127.7344, 126.8071, 
    125.8957, 125, 124.1198, 123.2547, 122.4046, 121.5691, 120.7478, 
    119.9406, 119.1471, 118.367, 117.6001, 116.8459,
  224.01, 223.2625, 222.5016, 221.7271, 220.9387, 220.136, 219.3185, 
    218.4861, 217.6384, 216.775, 215.8957, 215, 214.0877, 213.1585, 212.2121, 
    211.2482, 210.2666, 209.267, 208.2493, 207.2132, 206.1586, 205.0854, 
    203.9934, 202.8827, 201.7532, 200.605, 199.4382, 198.2528, 197.0491, 
    195.8274, 194.5879, 193.3311, 192.0573, 190.7672, 189.4613, 188.1401, 
    186.8046, 185.4553, 184.0933, 182.7194, 181.3346, 179.94, 178.5367, 
    177.1257, 175.7083, 174.2858, 172.8594, 171.4303, 170, 168.5697, 
    167.1406, 165.7142, 164.2917, 162.8743, 161.4633, 160.06, 158.6654, 
    157.2806, 155.9067, 154.5447, 153.1954, 151.8599, 150.5387, 149.2328, 
    147.9427, 146.6689, 145.4121, 144.1726, 142.9509, 141.7472, 140.5618, 
    139.395, 138.2468, 137.1173, 136.0066, 134.9146, 133.8414, 132.7868, 
    131.7507, 130.733, 129.7334, 128.7518, 127.7879, 126.8415, 125.9123, 125, 
    124.1043, 123.225, 122.3616, 121.5138, 120.6815, 119.8641, 119.0613, 
    118.2729, 117.4984, 116.7375, 115.99,
  224.8733, 224.1331, 223.3792, 222.6111, 221.8286, 221.0311, 220.2183, 
    219.39, 218.5455, 217.6847, 216.8071, 215.9123, 215, 214.0698, 213.1215, 
    212.1546, 211.1688, 210.164, 209.1397, 208.0958, 207.032, 205.9482, 
    204.8443, 203.7201, 202.5756, 201.4107, 200.2256, 199.0203, 197.7951, 
    196.55, 195.2856, 194.002, 192.6998, 191.3795, 190.0416, 188.687, 
    187.3164, 185.9305, 184.5304, 183.1171, 181.6915, 180.255, 178.8087, 
    177.3538, 175.8918, 174.424, 172.9518, 171.4766, 170, 168.5234, 167.0482, 
    165.576, 164.1082, 162.6462, 161.1913, 159.745, 158.3085, 156.8829, 
    155.4696, 154.0695, 152.6836, 151.313, 149.9584, 148.6205, 147.3002, 
    145.998, 144.7144, 143.45, 142.2049, 140.9797, 139.7744, 138.5893, 
    137.4244, 136.2799, 135.1557, 134.0518, 132.968, 131.9042, 130.8603, 
    129.836, 128.8312, 127.8454, 126.8785, 125.9302, 125, 124.0877, 123.1929, 
    122.3153, 121.4545, 120.6101, 119.7817, 118.9689, 118.1714, 117.3889, 
    116.6208, 115.8669, 115.1267,
  225.744, 225.0119, 224.2657, 223.5049, 222.729, 221.9376, 221.1304, 
    220.3069, 219.4667, 218.6094, 217.7344, 216.8415, 215.9302, 215, 
    214.0506, 213.0816, 212.0927, 211.0834, 210.0535, 209.0026, 207.9305, 
    206.8369, 205.7216, 204.5845, 203.4254, 202.2444, 201.0414, 199.8164, 
    198.5696, 197.3012, 196.0115, 194.7009, 193.3697, 192.0186, 190.6481, 
    189.259, 187.8522, 186.4284, 184.9888, 183.5343, 182.0663, 180.5859, 
    179.0946, 177.5938, 176.0848, 174.5694, 173.049, 171.5253, 170, 168.4747, 
    166.951, 165.4306, 163.9152, 162.4062, 160.9054, 159.4141, 157.9337, 
    156.4657, 155.0112, 153.5716, 152.1478, 150.741, 149.3519, 147.9814, 
    146.6303, 145.2991, 143.9885, 142.6988, 141.4304, 140.1836, 138.9586, 
    137.7556, 136.5746, 135.4155, 134.2784, 133.1631, 132.0695, 130.9974, 
    129.9465, 128.9166, 127.9073, 126.9184, 125.9494, 125, 124.0698, 
    123.1585, 122.2656, 121.3906, 120.5333, 119.6931, 118.8696, 118.0624, 
    117.271, 116.4951, 115.7343, 114.988, 114.256,
  226.6221, 225.8989, 225.1611, 224.4083, 223.64, 222.8557, 222.0549, 
    221.2372, 220.4022, 219.5493, 218.678, 217.7879, 216.8785, 215.9494, 215, 
    214.0299, 213.0388, 212.0261, 210.9914, 209.9344, 208.8548, 207.7522, 
    206.6264, 205.4771, 204.3041, 203.1074, 201.8868, 200.6424, 199.3743, 
    198.0826, 196.7676, 195.4296, 194.0691, 192.6865, 191.2826, 189.8581, 
    188.4138, 186.9508, 185.4701, 183.9728, 182.4604, 180.9342, 179.3957, 
    177.8465, 176.2883, 174.7227, 173.1516, 171.5767, 170, 168.4233, 
    166.8484, 165.2773, 163.7117, 162.1535, 160.6043, 159.0658, 157.5396, 
    156.0272, 154.5299, 153.0492, 151.5862, 150.1419, 148.7174, 147.3135, 
    145.9309, 144.5704, 143.2324, 141.9174, 140.6257, 139.3576, 138.1132, 
    136.8926, 135.6959, 134.5229, 133.3736, 132.2478, 131.1452, 130.0656, 
    129.0086, 127.9739, 126.9612, 125.9701, 125, 124.0506, 123.1215, 
    122.2121, 121.322, 120.4507, 119.5978, 118.7628, 117.9451, 117.1443, 
    116.36, 115.5917, 114.8389, 114.1011, 113.3779,
  227.5075, 226.794, 226.0655, 225.3216, 224.5616, 223.7852, 222.9918, 
    222.1809, 221.352, 220.5045, 219.638, 218.7518, 217.8454, 216.9184, 
    215.9701, 215, 214.0077, 212.9926, 211.9543, 210.8922, 209.8061, 
    208.6954, 207.5598, 206.3991, 205.213, 204.0012, 202.7636, 201.5002, 
    200.211, 198.8961, 197.5557, 196.1901, 194.7998, 193.3852, 191.9471, 
    190.4861, 189.0033, 187.4996, 185.9762, 184.4344, 182.8756, 181.3014, 
    179.7133, 178.1133, 176.5031, 174.8846, 173.2599, 171.631, 170, 168.369, 
    166.7401, 165.1154, 163.4969, 161.8867, 160.2867, 158.6986, 157.1244, 
    155.5656, 154.0238, 152.5004, 150.9967, 149.5139, 148.0529, 146.6148, 
    145.2002, 143.8099, 142.4443, 141.1039, 139.789, 138.4998, 137.2364, 
    135.9988, 134.787, 133.6009, 132.4402, 131.3046, 130.1939, 129.1078, 
    128.0457, 127.0074, 125.9923, 125, 124.0299, 123.0816, 122.1546, 
    121.2482, 120.362, 119.4954, 118.648, 117.8191, 117.0082, 116.2148, 
    115.4384, 114.6784, 113.9345, 113.206, 112.4925,
  228.4002, 227.6972, 226.9788, 226.2445, 225.4939, 224.7263, 223.9413, 
    223.1382, 222.3164, 221.4754, 220.6146, 219.7334, 218.8312, 217.9073, 
    216.9612, 215.9923, 215, 213.9837, 212.9428, 211.8768, 210.7852, 
    209.6675, 208.5232, 207.3519, 206.1534, 204.9273, 203.6733, 202.3914, 
    201.0815, 199.7436, 198.3779, 196.9846, 195.5641, 194.117, 192.6438, 
    191.1455, 189.6228, 188.077, 186.5092, 184.9209, 183.3136, 181.689, 
    180.0489, 178.3953, 176.7303, 175.0559, 173.3746, 171.6885, 170, 
    168.3115, 166.6254, 164.9441, 163.2697, 161.6047, 159.9511, 158.311, 
    156.6864, 155.0791, 153.4908, 151.923, 150.3772, 148.8545, 147.3562, 
    145.883, 144.4359, 143.0154, 141.6221, 140.2564, 138.9185, 137.6086, 
    136.3267, 135.0727, 133.8466, 132.6481, 131.4768, 130.3325, 129.2148, 
    128.1232, 127.0572, 126.0163, 125, 124.0077, 123.0388, 122.0927, 
    121.1688, 120.2666, 119.3854, 118.5246, 117.6836, 116.8618, 116.0587, 
    115.2737, 114.5061, 113.7555, 113.0212, 112.3028, 111.5998,
  229.3002, 228.6084, 227.9009, 227.1773, 226.4368, 225.679, 224.9033, 
    224.1089, 223.2954, 222.462, 221.608, 220.733, 219.836, 218.9166, 
    217.9739, 217.0074, 216.0163, 215, 213.9578, 212.8891, 211.7932, 
    210.6695, 209.5176, 208.3369, 207.1269, 205.8873, 204.6177, 203.3179, 
    201.9877, 200.6271, 199.2362, 197.8152, 196.3643, 194.8841, 193.3752, 
    191.8385, 190.2748, 188.6853, 187.0714, 185.4346, 183.7765, 182.099, 
    180.4041, 178.694, 176.971, 175.2375, 173.4962, 171.7494, 170, 168.2506, 
    166.5038, 164.7625, 163.029, 161.306, 159.5959, 157.901, 156.2235, 
    154.5654, 152.9286, 151.3147, 149.7252, 148.1615, 146.6248, 145.1159, 
    143.6357, 142.1848, 140.7638, 139.3729, 138.0123, 136.6821, 135.3823, 
    134.1127, 132.8731, 131.6631, 130.4824, 129.3305, 128.2068, 127.111, 
    126.0422, 125, 123.9837, 122.9926, 122.0261, 121.0834, 120.164, 119.267, 
    118.392, 117.538, 116.7046, 115.8911, 115.0967, 114.321, 113.5632, 
    112.8227, 112.0991, 111.3916, 110.6998,
  230.2074, 229.5276, 228.8319, 228.1197, 227.3904, 226.6433, 225.8778, 
    225.0933, 224.289, 223.4643, 222.6185, 221.7507, 220.8603, 219.9465, 
    219.0086, 218.0457, 217.0572, 216.0422, 215, 213.9298, 212.8309, 
    211.7027, 210.5443, 209.3553, 208.135, 206.8829, 205.5985, 204.2816, 
    202.9318, 201.549, 200.1331, 198.6844, 197.2029, 195.6893, 194.144, 
    192.5679, 190.9619, 189.3272, 187.6653, 185.9778, 184.2665, 182.5334, 
    180.7808, 179.011, 177.2267, 175.4305, 173.6254, 171.8142, 170, 168.1858, 
    166.3746, 164.5695, 162.7733, 160.989, 159.2192, 157.4666, 155.7335, 
    154.0222, 152.3347, 150.6728, 149.0381, 147.4321, 145.856, 144.3107, 
    142.7971, 141.3156, 139.8669, 138.451, 137.0682, 135.7184, 134.4015, 
    133.1171, 131.865, 130.6447, 129.4557, 128.2973, 127.169, 126.0702, 125, 
    123.9578, 122.9428, 121.9543, 120.9914, 120.0535, 119.1397, 118.2493, 
    117.3815, 116.5357, 115.711, 114.9067, 114.1222, 113.3567, 112.6096, 
    111.8803, 111.1681, 110.4724, 109.7927,
  231.1216, 230.4547, 229.7716, 229.0717, 228.3545, 227.6191, 226.865, 
    226.0913, 225.2975, 224.4826, 223.646, 222.7868, 221.9042, 220.9974, 
    220.0656, 219.1078, 218.1232, 217.1109, 216.0702, 215, 213.8996, 
    212.7681, 211.6047, 210.4086, 209.1792, 207.9158, 206.6177, 205.2846, 
    203.9159, 202.5115, 201.0711, 199.5948, 198.0828, 196.5353, 194.953, 
    193.3365, 191.687, 190.0056, 188.2939, 186.5534, 184.7863, 182.9947, 
    181.181, 179.3481, 177.4987, 175.6359, 173.763, 171.8832, 170, 168.1168, 
    166.237, 164.3641, 162.5013, 160.6519, 158.819, 157.0053, 155.2137, 
    153.4466, 151.7061, 149.9944, 148.313, 146.6635, 145.047, 143.4647, 
    141.9172, 140.4052, 138.9289, 137.4885, 136.0841, 134.7154, 133.3823, 
    132.0842, 130.8208, 129.5914, 128.3953, 127.2319, 126.1004, 125, 
    123.9298, 122.889, 121.8768, 120.8922, 119.9344, 119.0026, 118.0958, 
    117.2132, 116.354, 115.5174, 114.7025, 113.9087, 113.135, 112.3809, 
    111.6455, 110.9283, 110.2284, 109.5453, 108.8784,
  232.043, 231.3896, 230.72, 230.0334, 229.3291, 228.6064, 227.8646, 227.103, 
    226.3207, 225.5169, 224.6907, 223.8414, 222.968, 222.0695, 221.1452, 
    220.1939, 219.2148, 218.2068, 217.1691, 216.1004, 215, 213.8668, 
    212.6999, 211.4983, 210.2612, 208.9878, 207.6773, 206.329, 204.9425, 
    203.5172, 202.0529, 200.5494, 199.0068, 197.4253, 195.8054, 194.1478, 
    192.4535, 190.7238, 188.9601, 187.1643, 185.3386, 183.4854, 181.6073, 
    179.7074, 177.7889, 175.8552, 173.91, 171.9569, 170, 168.0431, 166.09, 
    164.1448, 162.2111, 160.2926, 158.3927, 156.5146, 154.6614, 152.8357, 
    151.0399, 149.2762, 147.5465, 145.8522, 144.1946, 142.5747, 140.9932, 
    139.4506, 137.9471, 136.4828, 135.0575, 133.671, 132.3227, 131.0122, 
    129.7388, 128.5017, 127.3001, 126.1332, 125, 123.8996, 122.831, 121.7932, 
    120.7852, 119.8061, 118.8548, 117.9305, 117.032, 116.1586, 115.3093, 
    114.4831, 113.6793, 112.897, 112.1354, 111.3936, 110.6709, 109.9666, 
    109.28, 108.6104, 107.957,
  232.9712, 232.3323, 231.677, 231.0045, 230.3142, 229.6052, 228.8768, 
    228.1283, 227.3587, 226.5671, 225.7527, 224.9146, 224.0518, 223.1631, 
    222.2478, 221.3046, 220.3325, 219.3305, 218.2973, 217.2319, 216.1332, 
    215, 213.8312, 212.6258, 211.3826, 210.1007, 208.7792, 207.4171, 
    206.0139, 204.5687, 203.0812, 201.551, 199.9781, 198.3625, 196.7047, 
    195.0052, 193.2649, 191.4852, 189.6676, 187.8141, 185.9268, 184.0086, 
    182.0623, 180.0913, 178.0992, 176.0898, 174.0672, 172.0359, 170, 
    167.9641, 165.9328, 163.9102, 161.9008, 159.9087, 157.9377, 155.9914, 
    154.0732, 152.1859, 150.3324, 148.5148, 146.7351, 144.9948, 143.2953, 
    141.6375, 140.0219, 138.449, 136.9188, 135.4313, 133.9861, 132.5829, 
    131.2208, 129.8993, 128.6174, 127.3742, 126.1688, 125, 123.8668, 
    122.7681, 121.7027, 120.6695, 119.6675, 118.6954, 117.7522, 116.8369, 
    115.9482, 115.0854, 114.2472, 113.4329, 112.6413, 111.8717, 111.1232, 
    110.3948, 109.6858, 108.9955, 108.323, 107.6677, 107.0288,
  233.9063, 233.2827, 232.6425, 231.985, 231.3096, 230.6153, 229.9015, 
    229.1671, 228.4114, 227.6334, 226.8321, 226.0066, 225.1557, 224.2784, 
    223.3736, 222.4402, 221.4768, 220.4824, 219.4557, 218.3953, 217.3001, 
    216.1688, 215, 213.7925, 212.5451, 211.2565, 209.9256, 208.5513, 
    207.1327, 205.6689, 204.1592, 202.6031, 201.0004, 199.3508, 197.6547, 
    195.9126, 194.1253, 192.294, 190.4204, 188.5065, 186.5546, 184.5678, 
    182.5491, 180.5025, 178.4318, 176.3414, 174.2361, 172.1206, 170, 
    167.8794, 165.7639, 163.6586, 161.5682, 159.4975, 157.4509, 155.4322, 
    153.4454, 151.4935, 149.5796, 147.706, 145.8747, 144.0874, 142.3453, 
    140.6492, 138.9996, 137.3969, 135.8408, 134.3311, 132.8673, 131.4487, 
    130.0744, 128.7435, 127.4549, 126.2075, 125, 123.8312, 122.6999, 
    121.6047, 120.5443, 119.5176, 118.5232, 117.5598, 116.6264, 115.7216, 
    114.8443, 113.9934, 113.1679, 112.3666, 111.5886, 110.8329, 110.0985, 
    109.3847, 108.6904, 108.015, 107.3575, 106.7173, 106.0937,
  234.8482, 234.2405, 233.6163, 232.9748, 232.3152, 231.6367, 230.9384, 
    230.2195, 229.4789, 228.7157, 227.9288, 227.1173, 226.2799, 225.4155, 
    224.5229, 223.6009, 222.6481, 221.6631, 220.6447, 219.5914, 218.5017, 
    217.3742, 216.2075, 215, 213.7503, 212.457, 211.1186, 209.7339, 208.3016, 
    206.8207, 205.2901, 203.7091, 202.0772, 200.394, 198.6597, 196.8744, 
    195.039, 193.1546, 191.2229, 189.2459, 187.2261, 185.1668, 183.0714, 
    180.944, 178.7893, 176.6121, 174.4178, 172.2118, 170, 167.7882, 165.5822, 
    163.3879, 161.2107, 159.056, 156.9286, 154.8332, 152.7739, 150.7541, 
    148.7771, 146.8454, 144.961, 143.1256, 141.3403, 139.606, 137.9228, 
    136.2909, 134.7099, 133.1793, 131.6984, 130.2661, 128.8814, 127.543, 
    126.2497, 125, 123.7925, 122.6258, 121.4983, 120.4086, 119.3553, 
    118.3369, 117.3519, 116.3991, 115.4771, 114.5845, 113.7201, 112.8827, 
    112.0712, 111.2843, 110.5211, 109.7805, 109.0616, 108.3633, 107.6848, 
    107.0252, 106.3837, 105.7595, 105.1518,
  235.7966, 235.2058, 234.5984, 233.9738, 233.331, 232.6692, 231.9876, 
    231.2852, 230.5609, 229.8138, 229.0428, 228.2468, 227.4244, 226.5746, 
    225.6959, 224.787, 223.8466, 222.8731, 221.865, 220.8208, 219.7388, 
    218.6174, 217.4549, 216.2497, 215, 213.7041, 212.3605, 210.9675, 
    209.5235, 208.0272, 206.4773, 204.8728, 203.2127, 201.4966, 199.7241, 
    197.8954, 196.0111, 194.0722, 192.0802, 190.0373, 187.9461, 185.8101, 
    183.6331, 181.4196, 179.1748, 176.9043, 174.614, 172.3103, 170, 167.6897, 
    165.386, 163.0957, 160.8252, 158.5804, 156.3669, 154.1899, 152.0539, 
    149.9627, 147.9198, 145.9278, 143.9889, 142.1046, 140.2759, 138.5034, 
    136.7873, 135.1272, 133.5227, 131.9728, 130.4765, 129.0325, 127.6395, 
    126.2958, 125, 123.7503, 122.5451, 121.3826, 120.2612, 119.1792, 118.135, 
    117.1269, 116.1534, 115.213, 114.3041, 113.4254, 112.5756, 111.7532, 
    110.9572, 110.1861, 109.4391, 108.7148, 108.0124, 107.3308, 106.669, 
    106.0262, 105.4016, 104.7942, 104.2034,
  236.7514, 236.1783, 235.5886, 234.9817, 234.3567, 233.7127, 233.0489, 
    232.3641, 231.6575, 230.9279, 230.1741, 229.395, 228.5893, 227.7556, 
    226.8926, 225.9988, 225.0727, 224.1127, 223.1171, 222.0842, 221.0122, 
    219.8993, 218.7435, 217.543, 216.2959, 215, 213.6535, 212.2546, 210.8012, 
    209.2917, 207.7245, 206.0981, 204.4113, 202.6631, 200.8531, 198.9809, 
    197.047, 195.0522, 192.9979, 190.8863, 188.7201, 186.5029, 184.239, 
    181.9334, 179.5918, 177.2205, 174.8266, 172.4172, 170, 167.5828, 
    165.1734, 162.7795, 160.4082, 158.0666, 155.761, 153.4971, 151.2799, 
    149.1137, 147.0021, 144.9478, 142.953, 141.0191, 139.1469, 137.3369, 
    135.5887, 133.9019, 132.2755, 130.7083, 129.1988, 127.7454, 126.3465, 
    125, 123.7042, 122.457, 121.2565, 120.1007, 118.9878, 117.9158, 116.8829, 
    115.8873, 114.9273, 114.0012, 113.1074, 112.2444, 111.4107, 110.605, 
    109.8259, 109.0721, 108.3425, 107.6359, 106.9511, 106.2873, 105.6433, 
    105.0183, 104.4114, 103.8217, 103.2486,
  237.7126, 237.1578, 236.5867, 235.9984, 235.3922, 234.767, 234.122, 
    233.4562, 232.7684, 232.0576, 231.3225, 230.5618, 229.7744, 228.9586, 
    228.1132, 227.2364, 226.3267, 225.3823, 224.4015, 223.3823, 222.3227, 
    221.2208, 220.0744, 218.8814, 217.6395, 216.3465, 215, 213.5979, 
    212.1378, 210.6177, 209.0356, 207.3894, 205.6776, 203.8988, 202.0521, 
    200.1368, 198.153, 196.1011, 193.9826, 191.7994, 189.5543, 187.2512, 
    184.8946, 182.4902, 180.0443, 177.5642, 175.0577, 172.5334, 170, 
    167.4666, 164.9423, 162.4358, 159.9557, 157.5098, 155.1054, 152.7488, 
    150.4457, 148.2006, 146.0174, 143.8989, 141.847, 139.8632, 137.9479, 
    136.1012, 134.3224, 132.6106, 130.9644, 129.3823, 127.8622, 126.4021, 
    125, 123.6535, 122.3605, 121.1186, 119.9256, 118.7792, 117.6773, 
    116.6177, 115.5985, 114.6177, 113.6733, 112.7636, 111.8868, 111.0414, 
    110.2256, 109.4382, 108.6775, 107.9424, 107.2316, 106.5438, 105.878, 
    105.233, 104.6078, 104.0016, 103.4133, 102.8422, 102.2874,
  238.6799, 238.1443, 237.5925, 237.0238, 236.4372, 235.8319, 235.2069, 
    234.5611, 233.8934, 233.2028, 232.4878, 231.7472, 230.9797, 230.1836, 
    229.3576, 228.4998, 227.6086, 226.6821, 225.7184, 224.7154, 223.671, 
    222.5829, 221.4487, 220.2661, 219.0325, 217.7454, 216.4021, 215, 
    213.5364, 212.0087, 210.4144, 208.7511, 207.0166, 205.2091, 203.3271, 
    201.3694, 199.3357, 197.226, 195.0414, 192.7838, 190.456, 188.0619, 
    185.6065, 183.0959, 180.5373, 177.9391, 175.3101, 172.6603, 170, 
    167.3397, 164.6899, 162.0609, 159.4627, 156.9041, 154.3935, 151.9381, 
    149.544, 147.2162, 144.9586, 142.774, 140.6643, 138.6306, 136.6729, 
    134.7909, 132.9834, 131.2489, 129.5856, 127.9913, 126.4636, 125, 
    123.5979, 122.2546, 120.9675, 119.7339, 118.5513, 117.4172, 116.329, 
    115.2846, 114.2816, 113.3179, 112.3914, 111.5002, 110.6424, 109.8164, 
    109.0203, 108.2528, 107.5122, 106.7972, 106.1066, 105.4389, 104.7931, 
    104.1681, 103.5628, 102.9762, 102.4075, 101.8557, 101.3201,
  239.6532, 239.1374, 238.6058, 238.0575, 237.4916, 236.9072, 236.3032, 
    235.6787, 235.0324, 234.3632, 233.6698, 232.9509, 232.2049, 231.4304, 
    230.6257, 229.789, 228.9185, 228.0123, 227.0682, 226.0841, 225.0575, 
    223.9861, 222.8673, 221.6984, 220.4765, 219.1988, 217.8622, 216.4636, 
    215, 213.4682, 211.8652, 210.188, 208.4338, 206.6, 204.6846, 202.6859, 
    200.6028, 198.4349, 196.1828, 193.8481, 191.4335, 188.943, 186.382, 
    183.7572, 181.0766, 178.3497, 175.5869, 172.7996, 170, 167.2004, 
    164.4131, 161.6503, 158.9234, 156.2428, 153.618, 151.057, 148.5665, 
    146.1519, 143.8172, 141.5651, 139.3972, 137.3141, 135.3154, 133.4, 
    131.5662, 129.812, 128.1348, 126.5318, 125, 123.5364, 122.1378, 120.8012, 
    119.5235, 118.3016, 117.1327, 116.0139, 114.9425, 113.9159, 112.9318, 
    111.9877, 111.0815, 110.211, 109.3743, 108.5696, 107.7951, 107.0491, 
    106.3302, 105.6368, 104.9676, 104.3213, 103.6968, 103.0928, 102.5084, 
    101.9425, 101.3942, 100.8626, 100.3468,
  240.6322, 240.1371, 239.6264, 239.0994, 238.5551, 237.9925, 237.4107, 
    236.8086, 236.185, 235.5387, 234.8684, 234.1726, 233.45, 232.6988, 
    231.9174, 231.1039, 230.2564, 229.3729, 228.451, 227.4885, 226.4828, 
    225.4313, 224.3311, 223.1793, 221.9728, 220.7083, 219.3823, 217.9913, 
    216.5318, 215, 213.3923, 211.705, 209.9346, 208.0779, 206.1319, 204.0941, 
    201.9628, 199.7368, 197.4161, 195.0019, 192.4965, 189.9041, 187.2302, 
    184.4821, 181.669, 178.8015, 175.8918, 172.9532, 170, 167.0468, 164.1082, 
    161.1985, 158.331, 155.5179, 152.7698, 150.0959, 147.5035, 144.9981, 
    142.5839, 140.2632, 138.0372, 135.9059, 133.8681, 131.9221, 130.0654, 
    128.295, 126.6077, 125, 123.4682, 122.0087, 120.6177, 119.2918, 118.0272, 
    116.8207, 115.6689, 114.5687, 113.5172, 112.5115, 111.549, 110.6271, 
    109.7436, 108.8961, 108.0826, 107.3012, 106.55, 105.8274, 105.1316, 
    104.4613, 103.815, 103.1914, 102.5893, 102.0075, 101.4449, 100.9006, 
    100.3735, 99.86288, 99.36778,
  241.6168, 241.1431, 240.6542, 240.1492, 239.6274, 239.0877, 238.5291, 
    237.9506, 237.3509, 236.7288, 236.083, 235.4121, 234.7144, 233.9885, 
    233.2324, 232.4443, 231.6221, 230.7638, 229.8669, 228.9289, 227.9471, 
    226.9188, 225.8408, 224.7099, 223.5227, 222.2755, 220.9644, 219.5856, 
    218.1348, 216.6077, 215, 213.3073, 211.5251, 209.6495, 207.6764, 
    205.6025, 203.4249, 201.1418, 198.7521, 196.2563, 193.6564, 190.9562, 
    188.1616, 185.2804, 182.3229, 179.3012, 176.2295, 173.1234, 170, 
    166.8766, 163.7705, 160.6988, 157.6771, 154.7196, 151.8384, 149.0438, 
    146.3436, 143.7437, 141.2479, 138.8582, 136.5751, 134.3975, 132.3236, 
    130.3505, 128.4749, 126.6928, 125, 123.3923, 121.8652, 120.4144, 
    119.0355, 117.7245, 116.4773, 115.2901, 114.1592, 113.0812, 112.0529, 
    111.0711, 110.1331, 109.2362, 108.3779, 107.5557, 106.7676, 106.0115, 
    105.2855, 104.5879, 103.917, 103.2712, 102.6491, 102.0494, 101.4709, 
    100.9123, 100.3726, 99.85078, 99.34584, 98.85692, 98.38318,
  242.6068, 242.1551, 241.6887, 241.2067, 240.7082, 240.1924, 239.6581, 
    239.1042, 238.5297, 237.9333, 237.3135, 236.6689, 235.998, 235.2991, 
    234.5704, 233.8099, 233.0154, 232.1848, 231.3156, 230.4052, 229.4506, 
    228.449, 227.3969, 226.2909, 225.1272, 223.9019, 222.6106, 221.2489, 
    219.812, 218.295, 216.6927, 215, 213.2115, 211.322, 209.3265, 207.2204, 
    204.9998, 202.6613, 200.2029, 197.6242, 194.9263, 192.1126, 189.1889, 
    186.1638, 183.0484, 179.8569, 176.6056, 173.3133, 170, 166.6867, 
    163.3944, 160.1431, 156.9516, 153.8362, 150.8111, 147.8874, 145.0737, 
    142.3758, 139.7971, 137.3387, 135.0002, 132.7796, 130.6735, 128.678, 
    126.7885, 125, 123.3072, 121.705, 120.188, 118.7511, 117.3894, 116.0981, 
    114.8728, 113.7091, 112.6031, 111.551, 110.5494, 109.5948, 108.6844, 
    107.8152, 106.9846, 106.1901, 105.4296, 104.7009, 104.002, 103.3311, 
    102.6865, 102.0667, 101.4703, 100.8958, 100.3419, 99.80763, 99.29177, 
    98.79331, 98.31132, 97.84489, 97.39321,
  243.6019, 243.1729, 242.7298, 242.2715, 241.7973, 241.3062, 240.7972, 
    240.2693, 239.7211, 239.1516, 238.5592, 237.9427, 237.3002, 236.6303, 
    235.9309, 235.2002, 234.4359, 233.6357, 232.7971, 231.9172, 230.9932, 
    230.0219, 228.9996, 227.9228, 226.7873, 225.5887, 224.3224, 222.9834, 
    221.5662, 220.0654, 218.4749, 216.7885, 215, 213.1029, 211.0909, 208.958, 
    206.6986, 204.308, 201.7826, 199.1205, 196.3217, 193.3888, 190.3274, 
    187.1464, 183.8581, 180.4786, 177.0273, 173.5263, 170, 166.4737, 
    162.9727, 159.5214, 156.1419, 152.8536, 149.6726, 146.6112, 143.6783, 
    140.8795, 138.2174, 135.692, 133.3014, 131.042, 128.9091, 126.8971, 125, 
    123.2115, 121.5251, 119.9346, 118.4338, 117.0166, 115.6776, 114.4113, 
    113.2127, 112.0772, 111.0003, 109.9781, 109.0068, 108.0828, 107.2029, 
    106.3643, 105.5641, 104.7998, 104.0691, 103.3697, 102.6998, 102.0574, 
    101.4408, 100.8484, 100.2789, 99.73074, 99.20277, 98.69379, 98.20271, 
    97.72851, 97.27025, 96.82706, 96.39812,
  244.6019, 244.1963, 243.7771, 243.3433, 242.8942, 242.4289, 241.9462, 
    241.4452, 240.9246, 240.3833, 239.8198, 239.2328, 238.6205, 237.9814, 
    237.3135, 236.6148, 235.883, 235.1159, 234.3107, 233.4647, 232.5747, 
    231.6375, 230.6492, 229.606, 228.5034, 227.3369, 226.1012, 224.7909, 
    223.4, 221.9221, 220.3505, 218.678, 216.8971, 215, 212.9789, 210.826, 
    208.534, 206.0961, 203.5069, 200.7623, 197.8607, 194.8035, 191.5955, 
    188.2456, 184.7673, 181.179, 177.5035, 173.7673, 170, 166.2327, 162.4965, 
    158.821, 155.2327, 151.7544, 148.4045, 145.1965, 142.1393, 139.2377, 
    136.4931, 133.9039, 131.466, 129.174, 127.0211, 125, 123.1029, 121.322, 
    119.6495, 118.0779, 116.6, 115.2091, 113.8988, 112.6631, 111.4966, 
    110.394, 109.3508, 108.3625, 107.4253, 106.5353, 105.6893, 104.8841, 
    104.117, 103.3852, 102.6865, 102.0186, 101.3794, 100.7672, 100.1802, 
    99.6167, 99.07538, 98.55483, 98.0538, 97.57114, 97.10576, 96.65666, 
    96.22292, 95.80368, 95.39812,
  245.6065, 245.225, 244.8304, 244.4219, 243.9987, 243.5599, 243.1045, 
    242.6315, 242.1397, 241.6279, 241.0947, 240.5387, 239.9584, 239.3519, 
    238.7174, 238.0529, 237.3562, 236.6248, 235.856, 235.047, 234.1946, 
    233.2953, 232.3453, 231.3403, 230.2759, 229.1469, 227.9479, 226.6729, 
    225.3154, 223.8681, 222.3236, 220.6735, 218.9091, 217.0211, 215, 212.836, 
    210.5196, 208.0415, 205.3936, 202.5694, 199.5649, 196.3791, 193.0156, 
    189.4829, 185.7955, 181.9741, 178.0455, 174.042, 170, 165.958, 161.9545, 
    158.0259, 154.2045, 150.5171, 146.9844, 143.6209, 140.4351, 137.4306, 
    134.6064, 131.9585, 129.4804, 127.164, 125, 122.9789, 121.0909, 119.3265, 
    117.6764, 116.1319, 114.6847, 113.3271, 112.0521, 110.8531, 109.7241, 
    108.6597, 107.6547, 106.7047, 105.8054, 104.953, 104.144, 103.3753, 
    102.6438, 101.9471, 101.2826, 100.6481, 100.0416, 99.46126, 98.90527, 
    98.37209, 97.86027, 97.36847, 96.89545, 96.44009, 96.0013, 95.57812, 
    95.16964, 94.77502, 94.39349,
  246.6156, 246.2586, 245.8893, 245.5068, 245.1103, 244.699, 244.2718, 
    243.8278, 243.3659, 242.8848, 242.3833, 241.8599, 241.313, 240.741, 
    240.1419, 239.5139, 238.8545, 238.1615, 237.4321, 236.6635, 235.8522, 
    234.9948, 234.0874, 233.1256, 232.1046, 231.0191, 229.8632, 228.6306, 
    227.3141, 225.9059, 224.3975, 222.7796, 221.042, 219.174, 217.164, 215, 
    212.6698, 210.1612, 207.4628, 204.5647, 201.4592, 198.1424, 194.6154, 
    190.8853, 186.9672, 182.8842, 178.6681, 174.3583, 170, 165.6417, 
    161.3319, 157.1158, 153.0328, 149.1147, 145.3846, 141.8576, 138.5408, 
    135.4353, 132.5372, 129.8388, 127.3302, 125, 122.836, 120.826, 118.958, 
    117.2204, 115.6025, 114.0941, 112.6859, 111.3694, 110.1368, 108.9809, 
    107.8954, 106.8744, 105.9126, 105.0052, 104.1478, 103.3366, 102.5679, 
    101.8385, 101.1455, 100.4862, 99.85809, 99.25905, 98.68702, 98.14013, 
    97.6167, 97.11516, 96.63409, 96.17216, 95.72819, 95.30104, 94.8897, 
    94.49322, 94.11072, 93.74137, 93.38445,
  247.6287, 247.297, 246.9535, 246.5977, 246.2286, 245.8455, 245.4475, 
    245.0336, 244.6026, 244.1535, 243.6849, 243.1954, 242.6836, 242.1478, 
    241.5862, 240.9967, 240.3772, 239.7252, 239.0381, 238.313, 237.5465, 
    236.7351, 235.8747, 234.961, 233.9889, 232.953, 231.847, 230.6643, 
    229.3972, 228.0372, 226.5751, 225.0002, 223.3014, 221.466, 219.4804, 
    217.3302, 215, 212.4741, 209.737, 206.7742, 203.5733, 200.1258, 196.4287, 
    192.4866, 188.314, 183.9362, 179.3909, 174.7264, 170, 165.2736, 160.6091, 
    156.0638, 151.686, 147.5134, 143.5713, 139.8742, 136.4267, 133.2258, 
    130.263, 127.5259, 125, 122.6698, 120.5196, 118.534, 116.6986, 114.9998, 
    113.4249, 111.9627, 110.6028, 109.3357, 108.153, 107.047, 106.0111, 
    105.039, 104.1253, 103.2649, 102.4535, 101.687, 100.9619, 100.2748, 
    99.62282, 99.0033, 98.41382, 97.85217, 97.31636, 96.80457, 96.31513, 
    95.84654, 95.3974, 94.96643, 94.55248, 94.15446, 93.77139, 93.40234, 
    93.04648, 92.70303, 92.37127,
  248.6458, 248.3397, 248.0227, 247.6941, 247.3532, 246.9992, 246.6311, 
    246.2481, 245.8492, 245.4331, 244.9987, 244.5447, 244.0695, 243.5716, 
    243.0492, 242.5004, 241.923, 241.3147, 240.6728, 239.9944, 239.2762, 
    238.5148, 237.706, 236.8454, 235.9278, 234.9478, 233.8989, 232.774, 
    231.5651, 230.2632, 228.8582, 227.3387, 225.692, 223.9039, 221.9585, 
    219.8388, 217.5259, 215, 212.2406, 209.2274, 205.9417, 202.3682, 
    198.4977, 194.33, 189.8769, 185.1656, 180.2401, 175.1604, 170, 164.8396, 
    159.7599, 154.8344, 150.1231, 145.67, 141.5023, 137.6318, 134.0583, 
    130.7726, 127.7594, 125, 122.4741, 120.1612, 118.0415, 116.0961, 114.308, 
    112.6613, 111.1418, 109.7368, 108.4349, 107.226, 106.1011, 105.0522, 
    104.0722, 103.1547, 102.294, 101.4852, 100.7238, 100.0056, 99.32724, 
    98.68533, 98.07699, 97.4996, 96.95078, 96.4284, 95.93051, 95.45535, 
    95.0013, 94.5669, 94.15083, 93.75185, 93.36886, 93.00081, 92.64677, 
    92.30585, 91.97729, 91.66032, 91.35426,
  249.6663, 249.3865, 249.0965, 248.7958, 248.4837, 248.1594, 247.8221, 
    247.471, 247.1049, 246.723, 246.324, 245.9067, 245.4696, 245.0112, 
    244.5299, 244.0238, 243.4908, 242.9286, 242.3347, 241.7061, 241.0399, 
    240.3324, 239.5796, 238.7771, 237.9198, 237.0021, 236.0174, 234.9586, 
    233.8172, 232.5839, 231.2479, 229.7971, 228.2174, 226.4931, 224.6064, 
    222.5372, 220.263, 217.7594, 215, 211.9573, 208.6043, 204.9164, 200.8747, 
    196.4705, 191.7102, 186.6204, 181.2519, 175.6798, 170, 164.3202, 
    158.7481, 153.3796, 148.2898, 143.5295, 139.1253, 135.0836, 131.3957, 
    128.0427, 125, 122.2406, 119.737, 117.4628, 115.3936, 113.5069, 111.7826, 
    110.2029, 108.7521, 107.4161, 106.1828, 105.0414, 103.9826, 102.9979, 
    102.0802, 101.2229, 100.4204, 99.66762, 98.96009, 98.29385, 97.66535, 
    97.07142, 96.50921, 95.97619, 95.47005, 94.98875, 94.5304, 94.09332, 
    93.67598, 93.27698, 92.89504, 92.52903, 92.17786, 91.84058, 91.5163, 
    91.20419, 90.9035, 90.61353, 90.33366,
  250.6902, 250.437, 250.1745, 249.9023, 249.6196, 249.3257, 249.0199, 
    248.7014, 248.3693, 248.0225, 247.66, 247.2806, 246.8829, 246.4657, 
    246.0272, 245.5656, 245.0791, 244.5654, 244.0222, 243.4466, 242.8357, 
    242.1859, 241.4935, 240.7541, 239.9627, 239.1137, 238.2006, 237.2162, 
    236.1519, 234.9981, 233.7437, 232.3758, 230.8795, 229.2377, 227.4306, 
    225.4353, 223.2258, 220.7726, 218.0427, 215, 211.6069, 207.826, 203.6246, 
    198.9797, 193.8866, 188.367, 182.4775, 176.3126, 170, 163.6874, 157.5225, 
    151.633, 146.1134, 141.0203, 136.3754, 132.174, 128.3931, 125, 121.9573, 
    119.2274, 116.7742, 114.5647, 112.5694, 110.7623, 109.1205, 107.6242, 
    106.2563, 105.0019, 103.8481, 102.7838, 101.7994, 100.8863, 100.0373, 
    99.24586, 98.50645, 97.81406, 97.16434, 96.55341, 95.97783, 95.43457, 
    94.92089, 94.43438, 93.97284, 93.53432, 93.11704, 92.71943, 92.34003, 
    91.97752, 91.63074, 91.29858, 90.98007, 90.6743, 90.38044, 90.09772, 
    89.82548, 89.56303, 89.30981,
  251.717, 251.4909, 251.2564, 251.0131, 250.7603, 250.4975, 250.2239, 
    249.9388, 249.6414, 249.3306, 249.0057, 248.6654, 248.3085, 247.9337, 
    247.5396, 247.1244, 246.6864, 246.2235, 245.7335, 245.2137, 244.6614, 
    244.0732, 243.4454, 242.7739, 242.0539, 241.2799, 240.4457, 239.544, 
    238.5665, 237.5035, 236.3436, 235.0737, 233.6783, 232.1393, 230.4351, 
    228.5408, 226.4267, 224.0583, 221.3957, 218.3931, 215, 211.1625, 
    206.8275, 201.9502, 196.5046, 190.4992, 183.9919, 177.1006, 170, 
    162.8994, 156.0081, 149.5008, 143.4954, 138.0498, 133.1725, 128.8375, 
    125, 121.6069, 118.6043, 115.9417, 113.5733, 111.4592, 109.5649, 
    107.8607, 106.3217, 104.9263, 103.6564, 102.4965, 101.4335, 100.456, 
    99.55431, 98.7201, 97.94613, 97.22612, 96.55462, 95.92685, 95.33863, 
    94.78626, 94.2665, 93.77647, 93.31358, 92.87559, 92.46043, 92.06629, 
    91.69152, 91.33465, 90.99432, 90.66936, 90.35864, 90.06119, 89.77608, 
    89.5025, 89.23968, 88.98693, 88.74361, 88.50915, 88.28298,
  252.7465, 252.5478, 252.3417, 252.1278, 251.9055, 251.6743, 251.4335, 
    251.1825, 250.9205, 250.6467, 250.3602, 250.06, 249.745, 249.4141, 
    249.0658, 248.6986, 248.311, 247.901, 247.4666, 247.0053, 246.5146, 
    245.9914, 245.4322, 244.8332, 244.1899, 243.4971, 242.7488, 241.9381, 
    241.057, 240.0959, 239.0438, 237.8874, 236.6112, 235.1965, 233.6209, 
    231.8576, 229.8742, 227.6318, 225.0836, 222.174, 218.8375, 215, 210.5811, 
    205.5019, 199.7001, 193.153, 185.908, 178.109, 170, 161.891, 154.092, 
    146.847, 140.2999, 134.4981, 129.4189, 125, 121.1625, 117.8261, 114.9164, 
    112.3682, 110.1258, 108.1424, 106.3791, 104.8035, 103.3888, 102.1126, 
    100.9562, 99.9041, 98.94302, 98.06187, 97.25119, 96.5029, 95.81008, 
    95.16676, 94.56776, 94.00861, 93.48539, 92.99465, 92.5334, 92.09896, 
    91.68898, 91.30136, 90.93423, 90.58595, 90.25499, 89.94002, 89.63983, 
    89.35334, 89.07954, 88.81754, 88.56652, 88.32574, 88.09452, 87.87224, 
    87.65831, 87.45223, 87.2535,
  253.7783, 253.6074, 253.43, 253.2459, 253.0545, 252.8554, 252.648, 
    252.4316, 252.2058, 251.9697, 251.7225, 251.4633, 251.1913, 250.9054, 
    250.6043, 250.2867, 249.9511, 249.5959, 249.2192, 248.819, 248.3927, 
    247.9377, 247.4509, 246.9286, 246.3669, 245.761, 245.1054, 244.3935, 
    243.618, 242.7698, 241.8384, 240.8111, 239.6726, 238.4045, 236.9844, 
    235.3846, 233.5713, 231.5023, 229.1253, 226.3754, 223.1725, 219.4189, 
    215, 209.7885, 203.661, 196.5311, 188.4048, 179.4445, 170, 160.5555, 
    151.5952, 143.4689, 136.339, 130.2115, 125, 120.5811, 116.8275, 113.6246, 
    110.8747, 108.4977, 106.4287, 104.6154, 103.0156, 101.5955, 100.3274, 
    99.18893, 98.1616, 97.23017, 96.382, 95.60646, 94.89464, 94.23899, 
    93.63306, 93.07137, 92.54916, 92.06232, 91.60732, 91.18104, 90.78075, 
    90.40408, 90.0489, 89.71334, 89.39574, 89.09463, 88.80865, 88.53665, 
    88.27754, 88.03036, 87.79422, 87.56836, 87.35204, 87.14461, 86.94548, 
    86.7541, 86.56998, 86.39264, 86.22168,
  254.8122, 254.6693, 254.521, 254.367, 254.2069, 254.0403, 253.8667, 
    253.6856, 253.4965, 253.2987, 253.0915, 252.8743, 252.6462, 252.4062, 
    252.1535, 251.8867, 251.6047, 251.306, 250.989, 250.6519, 250.2926, 
    249.9087, 249.4975, 249.056, 248.5804, 248.0666, 247.5098, 246.9041, 
    246.2428, 245.5179, 244.7196, 243.8362, 242.8536, 241.7544, 240.5171, 
    239.1147, 237.5134, 235.67, 233.5295, 231.0203, 228.0498, 224.4981, 
    220.2115, 215, 208.646, 200.9416, 191.7787, 181.2954, 170, 158.7046, 
    148.2213, 139.0584, 131.354, 125, 119.7885, 115.5019, 111.9502, 108.9797, 
    106.4705, 104.33, 102.4866, 100.8853, 99.48292, 98.24556, 97.14635, 
    96.16379, 95.28044, 94.48212, 93.75716, 93.09588, 92.49021, 91.93337, 
    91.41961, 90.94404, 90.50247, 90.0913, 89.70741, 89.3481, 89.01098, 
    88.69399, 88.3953, 88.1133, 87.84653, 87.59376, 87.35381, 87.12569, 
    86.90847, 86.70133, 86.50352, 86.31438, 86.13329, 85.95969, 85.79308, 
    85.633, 85.47902, 85.33075, 85.18784,
  255.8477, 255.7331, 255.6141, 255.4906, 255.3621, 255.2284, 255.089, 
    254.9436, 254.7917, 254.6328, 254.4663, 254.2917, 254.1082, 253.9152, 
    253.7117, 253.4969, 253.2697, 253.029, 252.7733, 252.5013, 252.2111, 
    251.9008, 251.5682, 251.2107, 250.8252, 250.4082, 249.9557, 249.4627, 
    248.9234, 248.331, 247.6771, 246.9516, 246.1419, 245.2327, 244.2045, 
    243.0328, 241.686, 240.1231, 238.2898, 236.1134, 233.4954, 230.2999, 
    226.339, 221.354, 215, 206.8593, 196.55, 184.0252, 170, 155.9748, 143.45, 
    133.1407, 125, 118.646, 113.661, 109.7001, 106.5046, 103.8865, 101.7102, 
    99.87689, 98.31396, 96.96719, 95.7955, 94.76733, 93.85809, 93.04843, 
    92.32288, 91.66899, 91.07659, 90.53735, 90.04433, 89.59177, 89.1748, 
    88.78931, 88.43176, 88.09916, 87.78889, 87.49871, 87.22665, 86.97101, 
    86.73026, 86.50307, 86.28828, 86.08483, 85.89179, 85.70834, 85.53371, 
    85.36723, 85.20831, 85.05639, 84.91096, 84.7716, 84.63787, 84.50941, 
    84.38586, 84.26693, 84.15231,
  256.8846, 256.7984, 256.709, 256.6162, 256.5196, 256.419, 256.3142, 
    256.2049, 256.0905, 255.971, 255.8457, 255.7142, 255.576, 255.4306, 
    255.2773, 255.1154, 254.9441, 254.7625, 254.5695, 254.3641, 254.1448, 
    253.9102, 253.6586, 253.3879, 253.0957, 252.7795, 252.4358, 252.0609, 
    251.6503, 251.1985, 250.6988, 250.1431, 249.5214, 248.821, 248.0259, 
    247.1158, 246.0638, 244.8344, 243.3796, 241.633, 239.5008, 236.847, 
    233.4689, 229.0584, 223.1407, 215, 203.6828, 188.4274, 170, 151.5726, 
    136.3172, 125, 116.8593, 110.9416, 106.5311, 103.153, 100.4992, 98.367, 
    96.62043, 95.16563, 93.93624, 92.88422, 91.97407, 91.17904, 90.47862, 
    89.85686, 89.30118, 88.80149, 88.34966, 87.93906, 87.5642, 87.22054, 
    86.90425, 86.61212, 86.34141, 86.08978, 85.8552, 85.63595, 85.4305, 
    85.23755, 85.05592, 84.88461, 84.72269, 84.56939, 84.42397, 84.28581, 
    84.15434, 84.02904, 83.90945, 83.79514, 83.68576, 83.58095, 83.48039, 
    83.38382, 83.29095, 83.20156, 83.11543,
  257.9225, 257.865, 257.8053, 257.7433, 257.6788, 257.6116, 257.5416, 
    257.4685, 257.3922, 257.3123, 257.2285, 257.1406, 257.0482, 256.951, 
    256.8484, 256.7401, 256.6254, 256.5038, 256.3746, 256.237, 256.0901, 
    255.9328, 255.7639, 255.5822, 255.386, 255.1734, 254.9423, 254.6899, 
    254.4131, 254.1082, 253.7705, 253.3944, 252.9727, 252.4965, 251.9545, 
    251.3319, 250.6091, 249.7599, 248.7481, 247.5225, 246.0081, 244.092, 
    241.5952, 238.2213, 233.45, 226.3172, 215, 196.5613, 170, 143.4387, 125, 
    113.6828, 106.55, 101.7787, 98.40478, 95.90804, 93.99186, 92.47754, 
    91.25187, 90.24007, 89.39088, 88.66811, 88.04547, 87.50346, 87.02731, 
    86.60561, 86.22946, 85.89178, 85.58688, 85.31013, 85.05774, 84.82656, 
    84.61398, 84.41776, 84.23605, 84.06725, 83.90996, 83.76301, 83.62537, 
    83.49615, 83.37456, 83.2599, 83.15157, 83.04901, 82.95177, 82.85939, 
    82.7715, 82.68775, 82.60783, 82.53146, 82.45838, 82.38837, 82.32121, 
    82.25671, 82.19471, 82.13503, 82.07752,
  258.9611, 258.9323, 258.9024, 258.8714, 258.8391, 258.8055, 258.7704, 
    258.7339, 258.6956, 258.6556, 258.6137, 258.5696, 258.5234, 258.4747, 
    258.4233, 258.369, 258.3115, 258.2506, 258.1858, 258.1168, 258.0431, 
    257.9641, 257.8794, 257.7882, 257.6896, 257.5828, 257.4666, 257.3397, 
    257.2004, 257.0468, 256.8766, 256.6867, 256.4737, 256.2327, 255.958, 
    255.6417, 255.2736, 254.8396, 254.3202, 253.6874, 252.8994, 251.891, 
    250.5555, 248.7046, 245.9748, 241.5726, 233.4387, 215, 170, 125, 
    106.5613, 98.42741, 94.02515, 91.29543, 89.44449, 88.10899, 87.10065, 
    86.31259, 85.67978, 85.16041, 84.72642, 84.35828, 84.042, 83.76727, 
    83.52634, 83.31327, 83.12345, 82.95321, 82.79963, 82.66034, 82.53339, 
    82.41718, 82.31036, 82.21181, 82.12057, 82.03585, 81.95693, 81.88322, 
    81.81421, 81.74942, 81.68847, 81.631, 81.57671, 81.52534, 81.47662, 
    81.43035, 81.38633, 81.34439, 81.30437, 81.26614, 81.22955, 81.19451, 
    81.16089, 81.12861, 81.09757, 81.0677, 81.03893,
  260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 
    260, 260, 260, 260, 260, 350, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 
    80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80,
  261.0389, 261.0677, 261.0976, 261.1286, 261.1609, 261.1945, 261.2296, 
    261.2661, 261.3044, 261.3444, 261.3863, 261.4304, 261.4766, 261.5253, 
    261.5767, 261.631, 261.6885, 261.7494, 261.8142, 261.8832, 261.9569, 
    262.0359, 262.1206, 262.2118, 262.3104, 262.4172, 262.5334, 262.6603, 
    262.7996, 262.9532, 263.1234, 263.3133, 263.5263, 263.7673, 264.042, 
    264.3583, 264.7264, 265.1604, 265.6798, 266.3126, 267.1006, 268.109, 
    269.4445, 271.2954, 274.0251, 278.4274, 286.5613, 305, 350, 35, 53.43872, 
    61.57259, 65.97485, 68.70457, 70.55551, 71.89101, 72.89935, 73.68741, 
    74.32022, 74.83959, 75.27358, 75.64172, 75.958, 76.23273, 76.47366, 
    76.68673, 76.87655, 77.04679, 77.20037, 77.33966, 77.46661, 77.58282, 
    77.68964, 77.78819, 77.87943, 77.96415, 78.04307, 78.11678, 78.18579, 
    78.25058, 78.31153, 78.369, 78.42329, 78.47466, 78.52338, 78.56965, 
    78.61367, 78.65561, 78.69563, 78.73386, 78.77045, 78.80549, 78.83911, 
    78.87139, 78.90243, 78.9323, 78.96107,
  262.0775, 262.135, 262.1947, 262.2567, 262.3212, 262.3884, 262.4584, 
    262.5315, 262.6078, 262.6877, 262.7715, 262.8594, 262.9518, 263.049, 
    263.1516, 263.2599, 263.3746, 263.4962, 263.6254, 263.763, 263.9099, 
    264.0672, 264.2361, 264.4178, 264.614, 264.8266, 265.0577, 265.3101, 
    265.5869, 265.8918, 266.2295, 266.6056, 267.0273, 267.5034, 268.0455, 
    268.6681, 269.3909, 270.2401, 271.2519, 272.4775, 273.9919, 275.908, 
    278.4048, 281.7787, 286.55, 293.6828, 305, 323.4387, 350, 16.56128, 35, 
    46.31718, 53.45003, 58.22134, 61.59522, 64.09196, 66.00814, 67.52246, 
    68.74813, 69.75993, 70.60912, 71.33189, 71.95453, 72.49654, 72.97269, 
    73.39439, 73.77054, 74.10822, 74.41312, 74.68987, 74.94226, 75.17344, 
    75.38602, 75.58224, 75.76395, 75.93275, 76.09004, 76.23699, 76.37463, 
    76.50385, 76.62544, 76.7401, 76.84843, 76.95099, 77.04823, 77.14061, 
    77.2285, 77.31225, 77.39217, 77.46854, 77.54162, 77.61163, 77.67879, 
    77.74329, 77.80529, 77.86497, 77.92248,
  263.1154, 263.2016, 263.291, 263.3838, 263.4804, 263.581, 263.6858, 
    263.7951, 263.9095, 264.029, 264.1543, 264.2858, 264.424, 264.5694, 
    264.7227, 264.8846, 265.0559, 265.2375, 265.4305, 265.636, 265.8552, 
    266.0898, 266.3414, 266.6121, 266.9043, 267.2206, 267.5642, 267.9391, 
    268.3497, 268.8015, 269.3012, 269.8569, 270.4786, 271.179, 271.9741, 
    272.8842, 273.9362, 275.1656, 276.6204, 278.367, 280.4992, 283.153, 
    286.5311, 290.9416, 296.8593, 305, 316.3172, 331.5726, 350, 8.427411, 
    23.68282, 35, 43.14066, 49.05843, 53.46891, 56.84695, 59.50083, 61.633, 
    63.37957, 64.83437, 66.06376, 67.11578, 68.02593, 68.82096, 69.52138, 
    70.14314, 70.69882, 71.19851, 71.65034, 72.06094, 72.4358, 72.77946, 
    73.09575, 73.38788, 73.65859, 73.91022, 74.1448, 74.36405, 74.5695, 
    74.76245, 74.94408, 75.11539, 75.27731, 75.43061, 75.57603, 75.71419, 
    75.84566, 75.97096, 76.09055, 76.20486, 76.31424, 76.41905, 76.51961, 
    76.61618, 76.70905, 76.79844, 76.88457,
  264.1523, 264.2669, 264.3859, 264.5094, 264.6379, 264.7716, 264.911, 
    265.0564, 265.2083, 265.3672, 265.5337, 265.7083, 265.8918, 266.0848, 
    266.2883, 266.5031, 266.7303, 266.971, 267.2267, 267.4987, 267.7889, 
    268.0992, 268.4318, 268.7893, 269.1748, 269.5918, 270.0443, 270.5374, 
    271.0766, 271.669, 272.3229, 273.0484, 273.8581, 274.7673, 275.7955, 
    276.9672, 278.314, 279.8769, 281.7102, 283.8865, 286.5046, 289.7002, 
    293.661, 298.646, 305, 313.1407, 323.45, 335.9749, 350, 4.025157, 
    16.54997, 26.85934, 35, 41.354, 46.33897, 50.29985, 53.49538, 56.11345, 
    58.2898, 60.12311, 61.68604, 63.03281, 64.2045, 65.23267, 66.14191, 
    66.95157, 67.67712, 68.33101, 68.92341, 69.46265, 69.95567, 70.40823, 
    70.8252, 71.21069, 71.56824, 71.90084, 72.21111, 72.50129, 72.77335, 
    73.02899, 73.26974, 73.49693, 73.71172, 73.91517, 74.10821, 74.29166, 
    74.46629, 74.63277, 74.79169, 74.94361, 75.08904, 75.2284, 75.36213, 
    75.49059, 75.61414, 75.73307, 75.84769,
  265.1878, 265.3307, 265.479, 265.633, 265.7931, 265.9597, 266.1333, 
    266.3144, 266.5035, 266.7013, 266.9085, 267.1257, 267.3538, 267.5938, 
    267.8465, 268.1133, 268.3953, 268.694, 269.011, 269.3481, 269.7074, 
    270.0913, 270.5025, 270.944, 271.4196, 271.9334, 272.4902, 273.0959, 
    273.7571, 274.4821, 275.2804, 276.1638, 277.1464, 278.2455, 279.4829, 
    280.8853, 282.4866, 284.33, 286.4705, 288.9797, 291.9502, 295.502, 
    299.7885, 305, 311.354, 319.0584, 328.2213, 338.7046, 350, 1.295434, 
    11.77866, 20.94157, 28.646, 35, 40.21146, 44.49806, 48.04982, 51.02029, 
    53.52949, 55.67005, 57.51336, 59.11468, 60.51708, 61.75444, 62.85364, 
    63.83621, 64.71956, 65.51788, 66.24284, 66.90412, 67.50979, 68.06663, 
    68.58039, 69.05596, 69.49753, 69.9087, 70.29259, 70.6519, 70.98902, 
    71.30601, 71.6047, 71.8867, 72.15347, 72.40624, 72.64619, 72.87431, 
    73.09153, 73.29867, 73.49648, 73.68562, 73.86671, 74.04031, 74.20692, 
    74.367, 74.52098, 74.66925, 74.81216,
  266.2217, 266.3926, 266.57, 266.7541, 266.9455, 267.1446, 267.3521, 
    267.5684, 267.7942, 268.0304, 268.2775, 268.5367, 268.8087, 269.0946, 
    269.3958, 269.7133, 270.0489, 270.4041, 270.7808, 271.181, 271.6073, 
    272.0623, 272.5492, 273.0714, 273.6331, 274.239, 274.8947, 275.6064, 
    276.382, 277.2302, 278.1616, 279.1889, 280.3274, 281.5955, 283.0156, 
    284.6154, 286.4287, 288.4977, 290.8747, 293.6246, 296.8275, 300.5811, 
    305, 310.2115, 316.339, 323.4689, 331.5952, 340.5555, 350, 359.4445, 
    8.404778, 16.53109, 23.66103, 29.78854, 35, 39.41894, 43.17246, 46.37541, 
    49.1253, 51.50228, 53.5713, 55.38464, 56.98439, 58.40453, 59.6726, 
    60.81107, 61.83841, 62.76982, 63.618, 64.39354, 65.10536, 65.76101, 
    66.36694, 66.92863, 67.45084, 67.93768, 68.39268, 68.81896, 69.21925, 
    69.59592, 69.9511, 70.28666, 70.60426, 70.90537, 71.19135, 71.46335, 
    71.72246, 71.96964, 72.20578, 72.43164, 72.64796, 72.85539, 73.05452, 
    73.2459, 73.43002, 73.60736, 73.77832,
  267.2535, 267.4522, 267.6583, 267.8722, 268.0945, 268.3257, 268.5665, 
    268.8175, 269.0795, 269.3533, 269.6398, 269.94, 270.255, 270.5859, 
    270.9342, 271.3014, 271.689, 272.099, 272.5334, 272.9947, 273.4854, 
    274.0086, 274.5677, 275.1667, 275.8101, 276.5029, 277.2512, 278.0619, 
    278.943, 279.9041, 280.9562, 282.1126, 283.3888, 284.8035, 286.3791, 
    288.1424, 290.1258, 292.3682, 294.9164, 297.826, 301.1625, 305, 309.4189, 
    314.498, 320.2998, 326.847, 334.092, 341.891, 350, 358.109, 5.908033, 
    13.15305, 19.70015, 25.50194, 30.58106, 35, 38.83752, 42.17395, 45.08361, 
    47.6318, 49.8742, 51.85757, 53.62088, 55.19647, 56.6112, 57.88741, 
    59.04377, 60.09591, 61.05698, 61.93813, 62.74881, 63.4971, 64.18992, 
    64.83324, 65.43224, 65.99139, 66.51461, 67.00535, 67.4666, 67.90104, 
    68.31102, 68.69864, 69.06577, 69.41405, 69.74501, 70.05998, 70.36017, 
    70.64666, 70.92046, 71.18246, 71.43348, 71.67426, 71.90548, 72.12776, 
    72.34169, 72.54777, 72.7465,
  268.283, 268.5092, 268.7436, 268.9869, 269.2397, 269.5025, 269.7761, 
    270.0612, 270.3586, 270.6694, 270.9943, 271.3347, 271.6915, 272.0663, 
    272.4604, 272.8756, 273.3136, 273.7765, 274.2665, 274.7863, 275.3386, 
    275.9268, 276.5546, 277.2261, 277.9461, 278.7201, 279.5543, 280.456, 
    281.4335, 282.4965, 283.6564, 284.9263, 286.3217, 287.8607, 289.5649, 
    291.4592, 293.5733, 295.9417, 298.6043, 301.6069, 305, 308.8375, 
    313.1725, 318.0498, 323.4954, 329.5008, 336.0081, 342.8994, 350, 
    357.1006, 3.991861, 10.49917, 16.50462, 21.95018, 26.82754, 31.16248, 35, 
    38.39312, 41.39567, 44.05833, 46.42671, 48.5408, 50.43513, 52.13926, 
    53.67833, 55.07372, 56.34361, 57.50347, 58.5665, 59.54401, 60.44569, 
    61.2799, 62.05387, 62.77388, 63.44538, 64.07315, 64.66137, 65.21374, 
    65.7335, 66.22353, 66.68642, 67.12441, 67.53957, 67.93371, 68.30848, 
    68.66535, 69.00568, 69.33064, 69.64136, 69.93881, 70.22392, 70.4975, 
    70.76032, 71.01307, 71.25639, 71.49085, 71.71702,
  269.3098, 269.563, 269.8255, 270.0977, 270.3804, 270.6743, 270.9801, 
    271.2986, 271.6307, 271.9775, 272.34, 272.7194, 273.117, 273.5343, 
    273.9728, 274.4344, 274.9209, 275.4346, 275.9778, 276.5534, 277.1643, 
    277.8141, 278.5064, 279.2459, 280.0373, 280.8863, 281.7993, 282.7838, 
    283.8481, 285.0019, 286.2563, 287.6242, 289.1205, 290.7623, 292.5694, 
    294.5647, 296.7742, 299.2274, 301.9573, 305, 308.3931, 312.174, 316.3754, 
    321.0203, 326.1135, 331.633, 337.5225, 343.6874, 350, 356.3126, 2.477536, 
    8.366995, 13.88655, 18.97971, 23.62459, 27.82605, 31.60689, 35, 38.04266, 
    40.77262, 43.22584, 45.43531, 47.43058, 49.23772, 50.87953, 52.37581, 
    53.74372, 54.99814, 56.15191, 57.21618, 58.20064, 59.11371, 59.96273, 
    60.75413, 61.49355, 62.18593, 62.83566, 63.4466, 64.02217, 64.56543, 
    65.07911, 65.56562, 66.02716, 66.46568, 66.88296, 67.28057, 67.65997, 
    68.02248, 68.36926, 68.70142, 69.01993, 69.3257, 69.61956, 69.90228, 
    70.17452, 70.43697, 70.69019,
  270.3337, 270.6135, 270.9035, 271.2042, 271.5163, 271.8406, 272.1779, 
    272.529, 272.8951, 273.277, 273.676, 274.0933, 274.5304, 274.9887, 
    275.4701, 275.9762, 276.5092, 277.0714, 277.6653, 278.2939, 278.9601, 
    279.6676, 280.4204, 281.2229, 282.0802, 282.9979, 283.9826, 285.0414, 
    286.1828, 287.4161, 288.7521, 290.2029, 291.7826, 293.5069, 295.3936, 
    297.4628, 299.737, 302.2406, 305, 308.0427, 311.3957, 315.0836, 319.1253, 
    323.5295, 328.2898, 333.3796, 338.7481, 344.3202, 350, 355.6798, 1.25187, 
    6.620432, 11.7102, 16.47051, 20.8747, 24.91639, 28.60433, 31.95734, 35, 
    37.75941, 40.263, 42.53716, 44.60641, 46.49313, 48.2174, 49.79707, 
    51.24794, 52.5839, 53.8172, 54.95856, 56.01741, 57.00206, 57.91981, 
    58.77709, 59.57961, 60.33239, 61.03991, 61.70615, 62.33465, 62.92859, 
    63.49079, 64.02381, 64.52995, 65.01125, 65.4696, 65.90668, 66.32402, 
    66.72302, 67.10496, 67.47097, 67.82214, 68.15942, 68.4837, 68.79581, 
    69.0965, 69.38647, 69.66634,
  271.3542, 271.6603, 271.9773, 272.3058, 272.6468, 273.0008, 273.3689, 
    273.7519, 274.1508, 274.5669, 275.0013, 275.4554, 275.9305, 276.4284, 
    276.9508, 277.4996, 278.077, 278.6853, 279.3272, 280.0056, 280.7238, 
    281.4852, 282.294, 283.1547, 284.0722, 285.0522, 286.1011, 287.226, 
    288.4349, 289.7368, 291.1418, 292.6613, 294.308, 296.0962, 298.0415, 
    300.1612, 302.4741, 305, 307.7594, 310.7726, 314.0583, 317.6318, 
    321.5023, 325.67, 330.1231, 334.8344, 339.7599, 344.8396, 350, 355.1604, 
    0.2400689, 5.165633, 9.876889, 14.32995, 18.49772, 22.3682, 25.94167, 
    29.22738, 32.24059, 35, 37.52589, 39.83878, 41.95853, 43.90385, 45.69201, 
    47.33874, 48.85823, 50.26324, 51.56511, 52.77399, 53.89887, 54.94778, 
    55.92782, 56.84534, 57.70599, 58.51479, 59.27624, 59.99436, 60.67276, 
    61.31467, 61.92302, 62.50041, 63.04922, 63.5716, 64.06949, 64.54465, 
    64.9987, 65.4331, 65.84917, 66.24815, 66.63114, 66.99919, 67.35323, 
    67.69415, 68.02271, 68.33968, 68.64574,
  272.3713, 272.703, 273.0465, 273.4023, 273.7714, 274.1544, 274.5525, 
    274.9664, 275.3974, 275.8465, 276.3151, 276.8046, 277.3163, 277.8522, 
    278.4138, 279.0033, 279.6228, 280.2748, 280.9619, 281.687, 282.4535, 
    283.2649, 284.1253, 285.039, 286.0111, 287.047, 288.153, 289.3357, 
    290.6028, 291.9627, 293.425, 294.9998, 296.6986, 298.534, 300.5196, 
    302.6698, 305, 307.5259, 310.263, 313.2258, 316.4267, 319.8742, 323.5713, 
    327.5134, 331.686, 336.0638, 340.6091, 345.2736, 350, 354.7264, 359.3909, 
    3.936238, 8.313965, 12.48664, 16.4287, 20.1258, 23.57329, 26.77416, 
    29.73699, 32.47411, 35, 37.33021, 39.48043, 41.46598, 43.30139, 45.00024, 
    46.57505, 48.03725, 49.39722, 50.66433, 51.84705, 52.95296, 53.98889, 
    54.96098, 55.87473, 56.73508, 57.54649, 58.31297, 59.03812, 59.72521, 
    60.37718, 60.9967, 61.58618, 62.14783, 62.68364, 63.19543, 63.68487, 
    64.15346, 64.6026, 65.03357, 65.44752, 65.84554, 66.22861, 66.59766, 
    66.95352, 67.29697, 67.62873,
  273.3844, 273.7414, 274.1107, 274.4932, 274.8897, 275.3011, 275.7282, 
    276.1721, 276.6341, 277.1151, 277.6167, 278.1401, 278.687, 279.2591, 
    279.8581, 280.4861, 281.1455, 281.8385, 282.5679, 283.3365, 284.1478, 
    285.0052, 285.9126, 286.8744, 287.8954, 288.981, 290.1368, 291.3694, 
    292.6859, 294.0941, 295.6025, 297.2205, 298.958, 300.826, 302.836, 305, 
    307.3302, 309.8388, 312.5372, 315.4353, 318.5408, 321.8576, 325.3846, 
    329.1147, 333.0328, 337.1158, 341.3319, 345.6417, 350, 354.3583, 
    358.6681, 2.884218, 6.967195, 10.88532, 14.61536, 18.14243, 21.4592, 
    24.56469, 27.46284, 30.16122, 32.66979, 35, 37.16397, 39.17396, 41.04199, 
    42.77955, 44.39749, 45.9059, 47.31408, 48.63058, 49.86321, 51.01906, 
    52.10457, 53.12559, 54.08742, 54.99484, 55.8522, 56.66345, 57.43214, 
    58.16152, 58.85453, 59.51385, 60.14192, 60.74095, 61.31298, 61.85987, 
    62.3833, 62.88484, 63.36592, 63.82784, 64.27181, 64.69896, 65.1103, 
    65.50678, 65.88928, 66.25863, 66.61555,
  274.3935, 274.775, 275.1696, 275.5781, 276.0013, 276.4401, 276.8954, 
    277.3685, 277.8603, 278.3721, 278.9053, 279.4612, 280.0416, 280.6481, 
    281.2826, 281.9471, 282.6438, 283.3752, 284.144, 284.953, 285.8054, 
    286.7047, 287.6547, 288.6597, 289.7241, 290.8531, 292.0521, 293.3271, 
    294.6847, 296.1319, 297.6764, 299.3265, 301.0909, 302.9789, 305, 307.164, 
    309.4804, 311.9585, 314.6064, 317.4306, 320.4351, 323.6209, 326.9844, 
    330.5171, 334.2045, 338.0259, 341.9545, 345.958, 350, 354.042, 358.0455, 
    1.974067, 5.795501, 9.482918, 13.01561, 16.37912, 19.56487, 22.56942, 
    25.39359, 28.04147, 30.51957, 32.83603, 35, 37.0211, 38.90907, 40.67348, 
    42.32358, 43.86813, 45.31535, 46.67292, 47.94793, 49.14692, 50.27589, 
    51.34034, 52.34529, 53.29532, 54.19463, 55.04703, 55.85601, 56.62475, 
    57.35616, 58.0529, 58.7174, 59.35187, 59.95836, 60.53875, 61.09473, 
    61.62791, 62.13973, 62.63153, 63.10454, 63.55991, 63.9987, 64.42188, 
    64.83036, 65.22498, 65.60651,
  275.3981, 275.8037, 276.2229, 276.6567, 277.1058, 277.5711, 278.0538, 
    278.5548, 279.0754, 279.6167, 280.1801, 280.7672, 281.3795, 282.0186, 
    282.6865, 283.3853, 284.117, 284.8841, 285.6893, 286.5353, 287.4253, 
    288.3625, 289.3508, 290.394, 291.4966, 292.6631, 293.8988, 295.2091, 
    296.6, 298.0779, 299.6495, 301.322, 303.1029, 305, 307.0211, 309.174, 
    311.466, 313.9038, 316.4931, 319.2377, 322.1393, 325.1965, 328.4045, 
    331.7545, 335.2327, 338.821, 342.4966, 346.2327, 350, 353.7673, 357.5034, 
    1.179037, 4.767325, 8.245557, 11.59547, 14.80353, 17.86074, 20.76228, 
    23.50687, 26.09615, 28.53402, 30.82604, 32.9789, 35, 36.89709, 38.67802, 
    40.35052, 41.92211, 43.39997, 44.79087, 46.10118, 47.33686, 48.50342, 
    49.60596, 50.64919, 51.63745, 52.57473, 53.4647, 54.31071, 55.11587, 
    55.88302, 56.61475, 57.31348, 57.9814, 58.62055, 59.23279, 59.81984, 
    60.3833, 60.92462, 61.44517, 61.94619, 62.42886, 62.89424, 63.34334, 
    63.77708, 64.19632, 64.60188,
  276.3981, 276.8271, 277.2703, 277.7285, 278.2027, 278.6938, 279.2028, 
    279.7307, 280.2789, 280.8484, 281.4408, 282.0573, 282.6998, 283.3697, 
    284.0691, 284.7998, 285.5641, 286.3643, 287.2029, 288.0828, 289.0067, 
    289.9781, 291.0003, 292.0772, 293.2127, 294.4113, 295.6776, 297.0166, 
    298.4337, 299.9346, 301.5251, 303.2115, 305, 306.8971, 308.9091, 311.042, 
    313.3014, 315.692, 318.2174, 320.8795, 323.6783, 326.6112, 329.6726, 
    332.8536, 336.1419, 339.5214, 342.9727, 346.4737, 350, 353.5263, 
    357.0273, 0.4786234, 3.858094, 7.146357, 10.3274, 13.3888, 16.32167, 
    19.12047, 21.7826, 24.30799, 26.69861, 28.95801, 31.09093, 33.10291, 35, 
    36.78852, 38.47487, 40.06539, 41.56625, 42.98337, 44.32241, 45.58871, 
    46.78728, 47.92281, 48.99965, 50.02188, 50.99324, 51.91722, 52.79705, 
    53.63569, 54.43589, 55.20019, 55.93093, 56.63028, 57.30024, 57.94265, 
    58.55923, 59.15157, 59.72112, 60.26925, 60.79723, 61.30621, 61.7973, 
    62.2715, 62.72975, 63.17294, 63.60188,
  277.3932, 277.8449, 278.3113, 278.7933, 279.2918, 279.8076, 280.3419, 
    280.8958, 281.4703, 282.0667, 282.6865, 283.3311, 284.002, 284.7009, 
    285.4296, 286.1902, 286.9846, 287.8152, 288.6844, 289.5948, 290.5494, 
    291.5511, 292.6031, 293.7091, 294.8728, 296.0981, 297.3894, 298.7511, 
    300.188, 301.705, 303.3073, 305, 306.7885, 308.678, 310.6735, 312.7795, 
    315.0002, 317.3387, 319.7971, 322.3758, 325.0737, 327.8874, 330.8111, 
    333.8362, 336.9516, 340.1431, 343.3944, 346.6867, 350, 353.3133, 
    356.6056, 359.8569, 3.048434, 6.163786, 9.188926, 12.11259, 14.92628, 
    17.62419, 20.20293, 22.66126, 24.99976, 27.22045, 29.32652, 31.32199, 
    33.21148, 35, 36.69275, 38.29502, 39.81203, 41.24892, 42.61062, 43.90189, 
    45.12722, 46.29089, 47.39688, 48.44895, 49.45062, 50.40517, 51.31562, 
    52.18483, 53.01543, 53.80986, 54.57038, 55.29913, 55.99803, 56.66891, 
    57.31347, 57.93325, 58.52973, 59.10424, 59.65807, 60.19236, 60.70823, 
    61.20669, 61.68868, 62.15511, 62.60678,
  278.3832, 278.8569, 279.3458, 279.8508, 280.3726, 280.9123, 281.4709, 
    282.0494, 282.6491, 283.2712, 283.917, 284.5879, 285.2856, 286.0115, 
    286.7676, 287.5557, 288.3778, 289.2362, 290.1331, 291.0711, 292.0529, 
    293.0812, 294.1592, 295.2901, 296.4773, 297.7245, 299.0356, 300.4144, 
    301.8652, 303.3923, 305, 306.6927, 308.4749, 310.3505, 312.3236, 
    314.3975, 316.575, 318.8582, 321.2479, 323.7437, 326.3436, 329.0438, 
    331.8384, 334.7196, 337.6771, 340.6988, 343.7705, 346.8766, 350, 
    353.1234, 356.2295, 359.3012, 2.322887, 5.280438, 8.161595, 10.95623, 
    13.65639, 16.25627, 18.75206, 21.14176, 23.42495, 25.60251, 27.67642, 
    29.64948, 31.52513, 33.30725, 35, 36.60772, 38.13481, 39.58562, 40.96445, 
    42.27547, 43.52268, 44.70991, 45.8408, 46.91879, 47.94713, 48.92886, 
    49.86686, 50.76379, 51.62215, 52.44429, 53.23239, 53.98848, 54.71445, 
    55.41209, 56.08303, 56.72881, 57.35088, 57.95056, 58.52911, 59.08768, 
    59.62738, 60.14923, 60.65416, 61.14308, 61.61683,
  279.3678, 279.8629, 280.3735, 280.9006, 281.4449, 282.0075, 282.5893, 
    283.1914, 283.815, 284.4613, 285.1317, 285.8274, 286.55, 287.3012, 
    288.0826, 288.8961, 289.7436, 290.6271, 291.549, 292.5115, 293.5172, 
    294.5687, 295.6689, 296.8207, 298.0272, 299.2917, 300.6177, 302.0087, 
    303.4682, 305, 306.6077, 308.295, 310.0654, 311.9221, 313.8681, 315.9059, 
    318.0373, 320.2632, 322.5839, 324.9981, 327.5035, 330.0959, 332.7698, 
    335.5179, 338.331, 341.1985, 344.1082, 347.0468, 350, 352.9532, 355.8918, 
    358.8015, 1.668989, 4.482118, 7.230175, 9.904095, 12.49653, 15.00186, 
    17.4161, 19.73676, 21.96275, 24.09411, 26.13187, 28.07789, 29.93461, 
    31.70498, 33.39228, 35, 36.53178, 37.99131, 39.38226, 40.70824, 41.9728, 
    43.17933, 44.33112, 45.43129, 46.48281, 47.48849, 48.45102, 49.37288, 
    50.25643, 51.1039, 51.91737, 52.69878, 53.44996, 54.17262, 54.86836, 
    55.53868, 56.18499, 56.80858, 57.41071, 57.99251, 58.55508, 59.09941, 
    59.62646, 60.13712, 60.63222,
  280.3468, 280.8625, 281.3942, 281.9425, 282.5084, 283.0928, 283.6968, 
    284.3214, 284.9676, 285.6368, 286.3302, 287.0491, 287.7951, 288.5696, 
    289.3743, 290.211, 291.0815, 291.9877, 292.9318, 293.916, 294.9425, 
    296.0139, 297.1327, 298.3016, 299.5235, 300.8012, 302.1378, 303.5364, 
    305, 306.5318, 308.1348, 309.812, 311.5663, 313.4, 315.3153, 317.3141, 
    319.3972, 321.5651, 323.8172, 326.1519, 328.5665, 331.057, 333.618, 
    336.2429, 338.9234, 341.6503, 344.4131, 347.2004, 350, 352.7996, 
    355.5869, 358.3497, 1.076589, 3.757156, 6.381995, 8.943019, 11.4335, 
    13.84809, 16.1828, 18.43489, 20.60278, 22.68592, 24.68465, 26.60003, 
    28.43375, 30.18797, 31.86519, 33.46822, 35, 36.46361, 37.86216, 39.19877, 
    40.47651, 41.69838, 42.86732, 43.98613, 45.05752, 46.08406, 47.06821, 
    48.0123, 48.91854, 49.78901, 50.62568, 51.4304, 52.20493, 52.95089, 
    53.66984, 54.36322, 55.0324, 55.67866, 56.3032, 56.90716, 57.49159, 
    58.0575, 58.60582, 59.13744, 59.65319,
  281.3201, 281.8557, 282.4075, 282.9762, 283.5628, 284.1681, 284.7931, 
    285.4389, 286.1065, 286.7972, 287.5122, 288.2528, 289.0204, 289.8164, 
    290.6424, 291.5002, 292.3914, 293.3179, 294.2816, 295.2846, 296.329, 
    297.4171, 298.5513, 299.7339, 300.9675, 302.2546, 303.5979, 305, 
    306.4636, 307.9913, 309.5856, 311.2489, 312.9834, 314.7909, 316.6729, 
    318.6306, 320.6643, 322.774, 324.9586, 327.2162, 329.544, 331.9381, 
    334.3936, 336.9041, 339.4626, 342.0609, 344.6899, 347.3397, 350, 
    352.6603, 355.3101, 357.9391, 0.5373426, 3.09588, 5.606458, 8.061871, 
    10.45599, 12.78382, 15.04144, 17.22602, 19.33566, 21.36942, 23.32708, 
    25.20913, 27.01663, 28.75108, 30.41438, 32.00869, 33.53639, 35, 36.40213, 
    37.74542, 39.03254, 40.26611, 41.44871, 42.58285, 43.67097, 44.7154, 
    45.71841, 46.68213, 47.60862, 48.49981, 49.35756, 50.18363, 50.97966, 
    51.74722, 52.48778, 53.20275, 53.89345, 54.5611, 55.20689, 55.83191, 
    56.43721, 57.02376, 57.59249, 58.14427, 58.67992,
  282.2874, 282.8422, 283.4133, 284.0016, 284.6078, 285.233, 285.878, 
    286.5438, 287.2316, 287.9424, 288.6776, 289.4381, 290.2256, 291.0414, 
    291.8868, 292.7636, 293.6733, 294.6177, 295.5985, 296.6177, 297.6773, 
    298.7792, 299.9256, 301.1186, 302.3605, 303.6535, 305, 306.4021, 
    307.8622, 309.3823, 310.9644, 312.6106, 314.3224, 316.1012, 317.9479, 
    319.8632, 321.847, 323.8989, 326.0174, 328.2007, 330.4457, 332.7488, 
    335.1053, 337.5098, 339.9557, 342.4358, 344.9423, 347.4666, 350, 
    352.5334, 355.0577, 357.5642, 0.04433093, 2.490215, 4.89464, 7.25119, 
    9.554314, 11.79936, 13.98259, 16.10113, 18.15295, 20.13679, 22.05207, 
    23.89882, 25.67759, 27.38938, 29.03555, 30.61774, 32.13784, 33.59787, 35, 
    36.34645, 37.6395, 38.8814, 40.07444, 41.22082, 42.32272, 43.38226, 
    44.40147, 45.38232, 46.3267, 47.23642, 48.11319, 48.95865, 49.77438, 
    50.56185, 51.32246, 52.05756, 52.7684, 53.45618, 54.12204, 54.76702, 
    55.39217, 55.99842, 56.58668, 57.15781, 57.71262,
  283.2486, 283.8217, 284.4114, 285.0183, 285.6433, 286.2873, 286.9511, 
    287.6359, 288.3425, 289.0721, 289.8259, 290.605, 291.4107, 292.2444, 
    293.1074, 294.0012, 294.9272, 295.8873, 296.8829, 297.9158, 298.9878, 
    300.1007, 301.2565, 302.457, 303.7042, 305, 306.3465, 307.7454, 309.1988, 
    310.7083, 312.2755, 313.9019, 315.5887, 317.3369, 319.1469, 321.019, 
    322.953, 324.9478, 327.0021, 329.1137, 331.2799, 333.4971, 335.761, 
    338.0666, 340.4082, 342.7794, 345.1734, 347.5828, 350, 352.4172, 
    354.8266, 357.2206, 359.5918, 1.933374, 4.238988, 6.502903, 8.720099, 
    10.88629, 12.99794, 15.05222, 17.04704, 18.98094, 20.85308, 22.66313, 
    24.41129, 26.09811, 27.72453, 29.29176, 30.80123, 32.25458, 33.65355, 35, 
    36.29585, 37.54304, 38.74353, 39.89928, 41.01221, 42.08421, 43.11712, 
    44.11272, 45.07275, 45.99885, 46.89263, 47.75561, 48.58926, 49.39498, 
    50.1741, 50.92786, 51.6575, 52.36414, 53.04887, 53.71273, 54.3567, 
    54.98169, 55.5886, 56.17825, 56.75144,
  284.2034, 284.7942, 285.4016, 286.0262, 286.669, 287.3307, 288.0124, 
    288.7148, 289.4391, 290.1862, 290.9572, 291.7532, 292.5756, 293.4254, 
    294.3041, 295.213, 296.1534, 297.1269, 298.135, 299.1792, 300.2612, 
    301.3826, 302.5451, 303.7503, 305, 306.2958, 307.6395, 309.0325, 
    310.4765, 311.9728, 313.5227, 315.1272, 316.7873, 318.5034, 320.2759, 
    322.1046, 323.9889, 325.9278, 327.9198, 329.9627, 332.0539, 334.1899, 
    336.3669, 338.5804, 340.8252, 343.0957, 345.386, 347.6896, 350, 352.3104, 
    354.614, 356.9043, 359.1748, 1.419612, 3.633067, 5.810081, 7.946126, 
    10.03727, 12.08019, 14.07218, 16.01111, 17.89543, 19.7241, 21.49658, 
    23.21272, 24.87277, 26.47732, 28.0272, 29.52349, 30.96746, 32.3605, 
    33.70415, 35, 36.2497, 37.45493, 38.6174, 39.73879, 40.82078, 41.86501, 
    42.8731, 43.8466, 44.78704, 45.6959, 46.57457, 47.42442, 48.24677, 
    49.04284, 49.81385, 50.56093, 51.28517, 51.98761, 52.66924, 53.33099, 
    53.97377, 54.59843, 55.20577, 55.79657,
  285.1519, 285.7595, 286.3837, 287.0252, 287.6848, 288.3633, 289.0616, 
    289.7805, 290.5211, 291.2843, 292.0712, 292.8827, 293.7201, 294.5845, 
    295.4771, 296.3991, 297.352, 298.3369, 299.3553, 300.4086, 301.4983, 
    302.6258, 303.7925, 305, 306.2497, 307.543, 308.8814, 310.2661, 311.6984, 
    313.1793, 314.7099, 316.2909, 317.9228, 319.606, 321.3403, 323.1256, 
    324.961, 326.8453, 328.7771, 330.7541, 332.7739, 334.8333, 336.9286, 
    339.056, 341.2107, 343.3879, 345.5822, 347.7882, 350, 352.2118, 354.4178, 
    356.6121, 358.7893, 0.9440413, 3.071369, 5.166756, 7.226121, 9.245869, 
    11.22291, 13.15465, 15.03902, 16.87441, 18.65966, 20.39404, 22.07719, 
    23.70911, 25.29009, 26.82067, 28.30161, 29.73389, 31.1186, 32.45696, 
    33.7503, 35, 36.20749, 37.37423, 38.50171, 39.59137, 40.6447, 41.66312, 
    42.64806, 43.60088, 44.52294, 45.41552, 46.2799, 47.11728, 47.92883, 
    48.71566, 49.47886, 50.21945, 50.93842, 51.63671, 52.31524, 52.97483, 
    53.61634, 54.24053, 54.84815,
  286.0937, 286.7173, 287.3575, 288.015, 288.6904, 289.3847, 290.0985, 
    290.8329, 291.5886, 292.3666, 293.1679, 293.9934, 294.8443, 295.7216, 
    296.6264, 297.5598, 298.5232, 299.5176, 300.5443, 301.6047, 302.6999, 
    303.8312, 305, 306.2075, 307.4549, 308.7435, 310.0744, 311.4487, 
    312.8673, 314.3311, 315.8408, 317.3969, 318.9997, 320.6492, 322.3453, 
    324.0874, 325.8747, 327.706, 329.5796, 331.4936, 333.4454, 335.4323, 
    337.4508, 339.4975, 341.5682, 343.6586, 345.7639, 347.8794, 350, 
    352.1206, 354.2361, 356.3414, 358.4318, 0.5024734, 2.549154, 4.567762, 
    6.554621, 8.506453, 10.42039, 12.29401, 14.12528, 15.91258, 17.65471, 
    19.35081, 21.00035, 22.60312, 24.1592, 25.66888, 27.13268, 28.55129, 
    29.92556, 31.25647, 32.54507, 33.79251, 35, 36.16879, 37.30013, 38.39533, 
    39.45566, 40.4824, 41.47682, 42.44015, 43.37363, 44.27842, 45.15569, 
    46.00657, 46.83212, 47.63339, 48.4114, 49.16711, 49.90145, 50.61533, 
    51.30958, 51.98503, 52.64248, 53.28267, 53.90633,
  287.0288, 287.6677, 288.323, 288.9955, 289.6859, 290.3948, 291.1232, 
    291.8717, 292.6414, 293.4329, 294.2473, 295.0854, 295.9482, 296.8369, 
    297.7522, 298.6954, 299.6674, 300.6695, 301.7027, 302.7681, 303.8668, 
    305, 306.1688, 307.3742, 308.6174, 309.8993, 311.2208, 312.5829, 
    313.9861, 315.4313, 316.9188, 318.4489, 320.0219, 321.6375, 323.2953, 
    324.9948, 326.7351, 328.5148, 330.3324, 332.1859, 334.0732, 335.9914, 
    337.9377, 339.9087, 341.9008, 343.9102, 345.9328, 347.9641, 350, 
    352.0359, 354.0672, 356.0898, 358.0992, 0.09130464, 2.062325, 4.008612, 
    5.926853, 7.814067, 9.667614, 11.48521, 13.26492, 15.00516, 16.70468, 
    18.36255, 19.97812, 21.55105, 23.08121, 24.56871, 26.01387, 27.41715, 
    28.77918, 30.10072, 31.3826, 32.62577, 33.83121, 35, 36.1332, 37.23193, 
    38.29732, 39.33048, 40.33253, 41.30461, 42.24778, 43.16315, 44.05175, 
    44.91462, 45.75275, 46.56712, 47.35865, 48.12827, 48.87683, 49.60519, 
    50.31416, 51.00451, 51.677, 52.33234, 52.97122,
  287.957, 288.6104, 289.28, 289.9666, 290.6709, 291.3936, 292.1353, 292.897, 
    293.6794, 294.4832, 295.3093, 296.1586, 297.032, 297.9305, 298.8548, 
    299.8061, 300.7852, 301.7932, 302.831, 303.8996, 305, 306.1332, 307.3001, 
    308.5017, 309.7388, 311.0122, 312.3227, 313.671, 315.0575, 316.4828, 
    317.9471, 319.4506, 320.9933, 322.5747, 324.1946, 325.8522, 327.5465, 
    329.2762, 331.0399, 332.8357, 334.6614, 336.5146, 338.3927, 340.2926, 
    342.2111, 344.1448, 346.0901, 348.0431, 350, 351.9569, 353.9099, 
    355.8552, 357.7889, 359.7074, 1.607323, 3.485386, 5.338629, 7.164339, 
    8.960093, 10.72376, 12.45351, 14.1478, 15.80537, 17.42527, 19.00676, 
    20.54938, 22.05287, 23.51719, 24.94248, 26.32903, 27.67728, 28.98779, 
    30.26121, 31.49829, 32.69987, 33.8668, 35, 36.10043, 37.16905, 38.20685, 
    39.21481, 40.19393, 41.14519, 42.06955, 42.96797, 43.84139, 44.69072, 
    45.51685, 46.32066, 47.10299, 47.86464, 48.60642, 49.32909, 50.03338, 
    50.72, 51.38964, 52.04295,
  288.8784, 289.5453, 290.2284, 290.9283, 291.6455, 292.3809, 293.135, 
    293.9087, 294.7025, 295.5174, 296.354, 297.2132, 298.0958, 299.0026, 
    299.9344, 300.8922, 301.8768, 302.889, 303.9298, 305, 306.1004, 307.2319, 
    308.3953, 309.5914, 310.8208, 312.0842, 313.3823, 314.7154, 316.084, 
    317.4885, 318.9289, 320.4052, 321.9172, 323.4647, 325.047, 326.6635, 
    328.313, 329.9944, 331.7061, 333.4466, 335.2137, 337.0053, 338.819, 
    340.6519, 342.5013, 344.364, 346.237, 348.1168, 350, 351.8832, 353.763, 
    355.636, 357.4987, 359.3481, 1.18104, 2.994655, 4.786263, 6.553403, 
    8.293855, 10.00564, 11.68703, 13.33655, 14.95297, 16.5353, 18.08277, 
    19.59484, 21.07113, 22.51151, 23.91594, 25.28459, 26.61774, 27.91578, 
    29.17922, 30.40863, 31.60467, 32.76807, 33.89957, 35, 36.07018, 37.11095, 
    38.1232, 39.10778, 40.06556, 40.99742, 41.90422, 42.78679, 43.64598, 
    44.4826, 45.29746, 46.09133, 46.86496, 47.6191, 48.35447, 49.07174, 
    49.7716, 50.45469, 51.12163,
  289.7927, 290.4724, 291.1681, 291.8803, 292.6096, 293.3567, 294.1222, 
    294.9067, 295.711, 296.5357, 297.3815, 298.2493, 299.1397, 300.0535, 
    300.9914, 301.9543, 302.9428, 303.9578, 305, 306.0702, 307.169, 308.2973, 
    309.4557, 310.6447, 311.865, 313.1171, 314.4015, 315.7184, 317.0682, 
    318.451, 319.8669, 321.3156, 322.7971, 324.3107, 325.856, 327.4321, 
    329.0381, 330.6728, 332.3347, 334.0222, 335.7335, 337.4666, 339.2192, 
    340.989, 342.7733, 344.5695, 346.3746, 348.1858, 350, 351.8142, 353.6254, 
    355.4305, 357.2267, 359.011, 0.7807565, 2.533401, 4.266501, 5.977829, 
    7.665351, 9.32724, 10.96188, 12.56786, 14.14399, 15.68929, 17.20295, 
    18.68438, 20.13314, 21.54898, 22.93179, 24.28159, 25.59853, 26.88288, 
    28.13499, 29.3553, 30.54434, 31.70268, 32.83095, 33.92982, 35, 36.04221, 
    37.05721, 38.04575, 39.00859, 39.94653, 40.86031, 41.7507, 42.61846, 
    43.46433, 44.28904, 45.0933, 45.87783, 46.64329, 47.39036, 48.11968, 
    48.83188, 49.52757, 50.20734,
  290.6998, 291.3916, 292.0991, 292.8227, 293.5632, 294.321, 295.0967, 
    295.8911, 296.7046, 297.538, 298.3919, 299.267, 300.164, 301.0834, 
    302.0261, 302.9926, 303.9837, 305, 306.0422, 307.111, 308.2068, 309.3305, 
    310.4824, 311.6631, 312.8731, 314.1127, 315.3823, 316.6821, 318.0123, 
    319.3729, 320.7638, 322.1848, 323.6357, 325.1159, 326.6248, 328.1615, 
    329.7252, 331.3147, 332.9286, 334.5654, 336.2235, 337.901, 339.5959, 
    341.306, 343.029, 344.7625, 346.5038, 348.2506, 350, 351.7494, 353.4962, 
    355.2375, 356.971, 358.694, 0.4040801, 2.098961, 3.776463, 5.434566, 
    7.071416, 8.685326, 10.27479, 11.83848, 13.37525, 14.88413, 16.36431, 
    17.81517, 19.23622, 20.62712, 21.9877, 23.31787, 24.61768, 25.88728, 
    27.1269, 28.33688, 29.5176, 30.66952, 31.79315, 32.88905, 33.95779, 35, 
    36.01632, 37.00741, 37.97394, 38.91659, 39.83604, 40.73296, 41.60805, 
    42.46196, 43.29537, 44.10892, 44.90327, 45.67903, 46.43683, 47.17727, 
    47.90092, 48.60838, 49.30018,
  291.5998, 292.3028, 293.0212, 293.7555, 294.5061, 295.2737, 296.0587, 
    296.8618, 297.6836, 298.5246, 299.3854, 300.2666, 301.1688, 302.0927, 
    303.0388, 304.0077, 305, 306.0163, 307.0572, 308.1232, 309.2148, 
    310.3326, 311.4768, 312.648, 313.8466, 315.0728, 316.3267, 317.6086, 
    318.9185, 320.2564, 321.6222, 323.0154, 324.4359, 325.883, 327.3562, 
    328.8545, 330.3772, 331.923, 333.4908, 335.0791, 336.6864, 338.311, 
    339.9511, 341.6047, 343.2697, 344.9441, 346.6254, 348.3115, 350, 
    351.6885, 353.3746, 355.0559, 356.7303, 358.3953, 0.04889843, 1.688978, 
    3.313586, 4.920894, 6.50921, 8.076985, 9.622821, 11.14547, 12.64384, 
    14.11698, 15.56411, 16.98457, 18.37785, 19.74357, 21.08146, 22.39138, 
    23.6733, 24.92726, 26.1534, 27.35194, 28.52318, 29.66747, 30.78519, 
    31.8768, 32.94279, 33.98368, 35, 35.99232, 36.96123, 37.90731, 38.83117, 
    39.73339, 40.61461, 41.47541, 42.31639, 43.13815, 43.94127, 44.72634, 
    45.49391, 46.24454, 46.97879, 47.69717, 48.40021,
  292.4925, 293.206, 293.9345, 294.6784, 295.4384, 296.2148, 297.0082, 
    297.8191, 298.648, 299.4955, 300.362, 301.2482, 302.1546, 303.0816, 
    304.0299, 305, 305.9923, 307.0074, 308.0457, 309.1078, 310.1939, 
    311.3046, 312.4402, 313.6009, 314.787, 315.9988, 317.2364, 318.4998, 
    319.789, 321.1039, 322.4443, 323.8098, 325.2002, 326.6147, 328.0529, 
    329.5139, 330.9967, 332.5004, 334.0238, 335.5656, 337.1244, 338.6986, 
    340.2867, 341.8867, 343.4969, 345.1154, 346.7401, 348.369, 350, 351.631, 
    353.2599, 354.8846, 356.5031, 358.1133, 359.7133, 1.301358, 2.875589, 
    4.434379, 5.976187, 7.499593, 9.003303, 10.48615, 11.9471, 13.38525, 
    14.79981, 16.19014, 17.55571, 18.8961, 20.21099, 21.50019, 22.76358, 
    24.00115, 25.21295, 26.39912, 27.55985, 28.69539, 29.80607, 30.89222, 
    31.95425, 32.99259, 34.00768, 35, 35.97005, 36.91836, 37.84542, 38.75179, 
    39.63799, 40.50455, 41.35203, 42.18094, 42.99183, 43.78522, 44.56163, 
    45.32156, 46.06552, 46.794, 47.50749,
  293.3779, 294.1011, 294.8388, 295.5917, 296.36, 297.1443, 297.9451, 
    298.7628, 299.5978, 300.4507, 301.322, 302.2121, 303.1215, 304.0506, 305, 
    305.9701, 306.9612, 307.9739, 309.0086, 310.0656, 311.1452, 312.2478, 
    313.3736, 314.5229, 315.6959, 316.8926, 318.1132, 319.3576, 320.6257, 
    321.9174, 323.2324, 324.5704, 325.9309, 327.3135, 328.7174, 330.1419, 
    331.5862, 333.0492, 334.5299, 336.0272, 337.5396, 339.0658, 340.6042, 
    342.1535, 343.7117, 345.2773, 346.8484, 348.4233, 350, 351.5767, 
    353.1516, 354.7227, 356.2883, 357.8465, 359.3958, 0.9342362, 2.460434, 
    3.97284, 5.470056, 6.950779, 8.413816, 9.858084, 11.28261, 12.68652, 
    14.06907, 15.42961, 16.76761, 18.08263, 19.37432, 20.64244, 21.88682, 
    23.10737, 24.3041, 25.47706, 26.62638, 27.75221, 28.85481, 29.93444, 
    30.9914, 32.02606, 33.03877, 34.02995, 35, 35.94938, 36.87852, 37.78791, 
    38.67799, 39.54926, 40.40218, 41.23724, 42.0549, 42.85566, 43.63998, 
    44.40832, 45.16115, 45.89892, 46.62207,
  294.256, 294.988, 295.7343, 296.4951, 297.271, 298.0624, 298.8696, 
    299.6931, 300.5333, 301.3906, 302.2656, 303.1585, 304.0699, 305, 
    305.9494, 306.9184, 307.9073, 308.9166, 309.9465, 310.9974, 312.0695, 
    313.1631, 314.2784, 315.4155, 316.5746, 317.7556, 318.9586, 320.1836, 
    321.4304, 322.6988, 323.9885, 325.2991, 326.6303, 327.9814, 329.3519, 
    330.7409, 332.1478, 333.5716, 335.0113, 336.4657, 337.9337, 339.4141, 
    340.9054, 342.4062, 343.9152, 345.4306, 346.951, 348.4747, 350, 351.5253, 
    353.049, 354.5694, 356.0848, 357.5938, 359.0946, 0.5859436, 2.066292, 
    3.534317, 4.988749, 6.428399, 7.852167, 9.259048, 10.64813, 12.01859, 
    13.36972, 14.70088, 16.01152, 17.30122, 18.5696, 19.81637, 21.04135, 
    22.24439, 23.42543, 24.58448, 25.72158, 26.83685, 27.93045, 29.00258, 
    30.05347, 31.08341, 32.09269, 33.08164, 34.05062, 35, 35.93016, 36.8415, 
    37.73442, 38.60936, 39.46672, 40.30694, 41.13043, 41.93763, 42.72896, 
    43.50485, 44.26571, 45.01196, 45.744,
  295.1267, 295.8669, 296.6208, 297.3889, 298.1714, 298.9689, 299.7816, 
    300.61, 301.4545, 302.3153, 303.1929, 304.0877, 305, 305.9301, 306.8785, 
    307.8454, 308.8312, 309.836, 310.8603, 311.9042, 312.968, 314.0518, 
    315.1557, 316.2799, 317.4244, 318.5893, 319.7744, 320.9796, 322.2049, 
    323.45, 324.7144, 325.998, 327.3002, 328.6205, 329.9584, 331.313, 
    332.6837, 334.0695, 335.4696, 336.883, 338.3085, 339.745, 341.1913, 
    342.6462, 344.1082, 345.576, 347.0482, 348.5234, 350, 351.4766, 352.9518, 
    354.424, 355.8918, 357.3538, 358.8087, 0.2549859, 1.691522, 3.117045, 
    4.530401, 5.930508, 7.316357, 8.687016, 10.04164, 11.37945, 12.69976, 
    14.00197, 15.28555, 16.55004, 17.79507, 19.02034, 20.22562, 21.41073, 
    22.57558, 23.7201, 24.84431, 25.94825, 27.03203, 28.09578, 29.13969, 
    30.16396, 31.16883, 32.15458, 33.12148, 34.06984, 35, 35.91229, 36.80707, 
    37.68469, 38.54552, 39.38995, 40.21834, 41.03108, 41.82855, 42.61113, 
    43.3792, 44.13313, 44.87331,
  295.99, 296.7375, 297.4984, 298.2729, 299.0613, 299.864, 300.6815, 
    301.5139, 302.3616, 303.2249, 304.1043, 305, 305.9123, 306.8415, 
    307.7879, 308.7518, 309.7334, 310.733, 311.7507, 312.7868, 313.8414, 
    314.9146, 316.0066, 317.1173, 318.2468, 319.395, 320.5619, 321.7472, 
    322.9509, 324.1726, 325.4121, 326.6689, 327.9427, 329.2328, 330.5388, 
    331.8599, 333.1954, 334.5446, 335.9067, 337.2806, 338.6653, 340.06, 
    341.4633, 342.8743, 344.2917, 345.7142, 347.1406, 348.5696, 350, 
    351.4304, 352.8594, 354.2858, 355.7083, 357.1257, 358.5367, 359.94, 
    1.334645, 2.719428, 4.093322, 5.455343, 6.804565, 8.140132, 9.461254, 
    10.76721, 12.05735, 13.33109, 14.58791, 15.82738, 17.04911, 18.25278, 
    19.43815, 20.60502, 21.75323, 22.88272, 23.99343, 25.08538, 26.15861, 
    27.21321, 28.2493, 29.26704, 30.2666, 31.24821, 32.21209, 33.1585, 
    34.08771, 35, 35.89568, 36.77504, 37.63843, 38.48615, 39.31855, 40.13595, 
    40.93871, 41.72715, 42.50162, 43.26246, 44.01001,
  296.8459, 297.6001, 298.367, 299.1471, 299.9406, 300.7478, 301.5691, 
    302.4046, 303.2547, 304.1198, 305, 305.8957, 306.8071, 307.7344, 308.678, 
    309.638, 310.6146, 311.6081, 312.6185, 313.646, 314.6907, 315.7527, 
    316.8321, 317.9288, 319.0428, 320.1741, 321.3224, 322.4878, 323.6698, 
    324.8683, 326.083, 327.3135, 328.5592, 329.8199, 331.0947, 332.3833, 
    333.6849, 334.9987, 336.324, 337.66, 339.0057, 340.3602, 341.7225, 
    343.0915, 344.4663, 345.8457, 347.2285, 348.6137, 350, 351.3863, 
    352.7715, 354.1543, 355.5337, 356.9085, 358.2775, 359.6398, 0.9943273, 
    2.340024, 3.675979, 5.001296, 6.315132, 7.616698, 8.905264, 10.18016, 
    11.44077, 12.68653, 13.91697, 15.13164, 16.33016, 17.51222, 18.67754, 
    19.82591, 20.95716, 22.07118, 23.16788, 24.24725, 25.30928, 26.35402, 
    27.38154, 28.39195, 29.38539, 30.36201, 31.32201, 32.26558, 33.19293, 
    34.10432, 35, 35.88022, 36.74526, 37.59541, 38.43094, 39.25217, 40.05937, 
    40.85287, 41.63295, 42.39994, 43.15412,
  297.6943, 298.4544, 299.2268, 300.0117, 300.8095, 301.6204, 302.4446, 
    303.2824, 304.1342, 305, 305.8802, 306.7751, 307.6847, 308.6094, 
    309.5493, 310.5045, 311.4754, 312.462, 313.4643, 314.4826, 315.5168, 
    316.5671, 317.6334, 318.7157, 319.8138, 320.9279, 322.0576, 323.2028, 
    324.3632, 325.5387, 326.7288, 327.9333, 329.1516, 330.3833, 331.6279, 
    332.8849, 334.1535, 335.4331, 336.723, 338.0225, 339.3306, 340.6467, 
    341.9696, 343.2987, 344.6328, 345.971, 347.3123, 348.6556, 350, 351.3444, 
    352.6877, 354.029, 355.3672, 356.7013, 358.0304, 359.3533, 0.6693593, 
    1.977523, 3.276976, 4.566904, 5.846539, 7.115158, 8.372087, 9.616703, 
    10.84843, 12.06675, 13.27118, 14.46132, 15.63678, 16.79724, 17.94244, 
    19.07214, 20.18615, 21.28434, 22.36661, 23.43288, 24.48314, 25.5174, 
    26.53567, 27.53804, 28.52459, 29.49545, 30.45074, 31.39064, 32.31531, 
    33.22496, 34.11978, 35, 35.86585, 36.71758, 37.55542, 38.37964, 39.19049, 
    39.98825, 40.77319, 41.54556, 42.30565,
  298.5354, 299.3007, 300.0777, 300.8667, 301.668, 302.4817, 303.3082, 
    304.1475, 305, 305.8658, 306.7453, 307.6384, 308.5455, 309.4667, 
    310.4022, 311.352, 312.3164, 313.2954, 314.289, 315.2975, 316.3206, 
    317.3586, 318.4114, 319.4789, 320.5609, 321.6575, 322.7684, 323.8935, 
    325.0324, 326.185, 327.3509, 328.5297, 329.7211, 330.9246, 332.1397, 
    333.3659, 334.6026, 335.8492, 337.1049, 338.3693, 339.6414, 340.9205, 
    342.2058, 343.4965, 344.7917, 346.0905, 347.3922, 348.6956, 350, 
    351.3044, 352.6078, 353.9095, 355.2083, 356.5035, 357.7942, 359.0795, 
    0.3586455, 1.630737, 2.895045, 4.150831, 5.397398, 6.634083, 7.86027, 
    9.075379, 10.27888, 11.47027, 12.64912, 13.81502, 14.9676, 16.10655, 
    17.2316, 18.3425, 19.43907, 20.52114, 21.5886, 22.64135, 23.67934, 
    24.70254, 25.71096, 26.70463, 27.68361, 28.64797, 29.59782, 30.53328, 
    31.45448, 32.36157, 33.25474, 34.13415, 35, 35.8525, 36.69184, 37.51827, 
    38.332, 39.13326, 39.92228, 40.69931, 41.46459,
  299.3691, 300.1388, 300.9198, 301.7122, 302.5162, 303.332, 304.1599, 305, 
    305.8525, 306.7176, 307.5954, 308.4861, 309.39, 310.3069, 311.2372, 
    312.1809, 313.1382, 314.1089, 315.0933, 316.0913, 317.103, 318.1283, 
    319.1671, 320.2195, 321.2852, 322.3641, 323.4562, 324.5611, 325.6786, 
    326.8086, 327.9506, 329.1042, 330.2693, 331.4452, 332.6315, 333.8279, 
    335.0336, 336.2481, 337.471, 338.7014, 339.9388, 341.1825, 342.4316, 
    343.6856, 344.9436, 346.2049, 347.4685, 348.7339, 350, 351.2661, 
    352.5315, 353.7951, 355.0564, 356.3144, 357.5684, 358.8175, 0.0611895, 
    1.298583, 2.529026, 3.751855, 4.966434, 6.172163, 7.368472, 8.554832, 
    9.730745, 10.89576, 12.04944, 13.19142, 14.32134, 15.4389, 16.54382, 
    17.63586, 18.71483, 19.78055, 20.83289, 21.87173, 22.89701, 23.90867, 
    24.90669, 25.89108, 26.86185, 27.81906, 28.76277, 29.69306, 30.61005, 
    31.51385, 32.40459, 33.28242, 34.1475, 35, 35.84009, 36.66796, 37.4838, 
    38.28781, 39.0802, 39.86116, 40.63093,
  300.1953, 300.9689, 301.7531, 302.5482, 303.3542, 304.1714, 305, 305.8401, 
    306.6918, 307.5554, 308.4309, 309.3185, 310.2184, 311.1304, 312.0549, 
    312.9918, 313.9413, 314.9033, 315.8778, 316.865, 317.8647, 318.8768, 
    319.9015, 320.9384, 321.9876, 323.0489, 324.122, 325.2069, 326.3032, 
    327.4107, 328.5291, 329.6581, 330.7972, 331.9462, 333.1046, 334.2718, 
    335.4475, 336.6311, 337.8221, 339.0199, 340.2239, 341.4335, 342.6479, 
    343.8667, 345.089, 346.3142, 347.5416, 348.7704, 350, 351.2296, 352.4584, 
    353.6858, 354.911, 356.1333, 357.3521, 358.5665, 359.7761, 0.9800709, 
    2.177862, 3.368856, 4.55248, 5.728187, 6.895458, 8.053806, 9.202773, 
    10.34193, 11.47089, 12.58929, 13.6968, 14.79311, 15.87796, 16.95113, 
    18.01239, 19.06158, 20.09855, 21.12317, 22.13536, 23.13504, 24.12217, 
    25.09674, 26.05873, 27.00817, 27.9451, 28.86957, 29.78166, 30.68145, 
    31.56906, 32.44458, 33.30816, 34.15991, 35, 35.82858, 36.6458, 37.45184, 
    38.24688, 39.03109, 39.80465,
  301.0143, 301.791, 302.5777, 303.3747, 304.1821, 305, 305.8286, 306.668, 
    307.5183, 308.3796, 309.2522, 310.136, 311.0311, 311.9376, 312.8557, 
    313.7852, 314.7263, 315.679, 316.6433, 317.6191, 318.6064, 319.6052, 
    320.6153, 321.6367, 322.6693, 323.7127, 324.767, 325.8319, 326.9072, 
    327.9925, 329.0877, 330.1924, 331.3062, 332.4289, 333.5599, 334.6989, 
    335.8456, 336.9992, 338.1594, 339.3257, 340.4975, 341.6743, 342.8554, 
    344.0403, 345.2284, 346.419, 347.6116, 348.8055, 350, 351.1945, 352.3884, 
    353.581, 354.7716, 355.9597, 357.1446, 358.3257, 359.5025, 0.6742983, 
    1.840581, 3.000807, 4.154459, 5.301043, 6.440085, 7.57114, 8.693789, 
    9.807635, 10.91231, 12.00749, 13.09284, 14.16809, 15.23297, 16.28727, 
    17.33076, 18.36328, 19.38468, 20.39481, 21.39358, 22.3809, 23.35671, 
    24.32097, 25.27366, 26.21478, 27.14434, 28.06237, 28.96892, 29.86405, 
    30.74784, 31.62036, 32.48173, 33.33204, 34.17142, 35, 35.8179, 36.62528, 
    37.42227, 38.20903, 38.98572,
  301.8259, 302.605, 303.3937, 304.192, 305, 305.8179, 306.6458, 307.4838, 
    308.332, 309.1905, 310.0594, 310.9387, 311.8286, 312.729, 313.64, 
    314.5616, 315.4939, 316.4368, 317.3904, 318.3545, 319.3291, 320.3141, 
    321.3096, 322.3152, 323.331, 324.3567, 325.3922, 326.4372, 327.4916, 
    328.5551, 329.6274, 330.7082, 331.7973, 332.8942, 333.9987, 335.1103, 
    336.2286, 337.3532, 338.4837, 339.6196, 340.7603, 341.9055, 343.0545, 
    344.2069, 345.3621, 346.5196, 347.6788, 348.8391, 350, 351.1609, 
    352.3212, 353.4804, 354.6379, 355.7931, 356.9455, 358.0945, 359.2397, 
    0.3804374, 1.516293, 2.646764, 3.771384, 4.889704, 6.001298, 7.105759, 
    8.202703, 9.291768, 10.37261, 11.44492, 12.50841, 13.56279, 14.60783, 
    15.6433, 16.66901, 17.68477, 18.69042, 19.68584, 20.67091, 21.64553, 
    22.60964, 23.56317, 24.50609, 25.43838, 26.36002, 27.27104, 28.17145, 
    29.0613, 29.94063, 30.8095, 31.668, 32.5162, 33.3542, 34.1821, 35, 
    35.80803, 36.6063, 37.39495, 38.17411,
  302.6302, 303.4112, 304.2011, 305, 305.808, 306.6253, 307.4518, 308.2878, 
    309.1333, 309.9883, 310.8529, 311.7271, 312.6111, 313.5049, 314.4083, 
    315.3216, 316.2445, 317.1773, 318.1197, 319.0717, 320.0334, 321.0045, 
    321.985, 322.9748, 323.9738, 324.9817, 325.9984, 327.0238, 328.0575, 
    329.0994, 330.1492, 331.2067, 332.2715, 333.3433, 334.4219, 335.5068, 
    336.5977, 337.6942, 338.7958, 339.9023, 341.0131, 342.1278, 343.2459, 
    344.367, 345.4906, 346.6162, 347.7433, 348.8714, 350, 351.1286, 352.2567, 
    353.3838, 354.5094, 355.633, 356.7541, 357.8722, 358.9869, 0.09772872, 
    1.204182, 2.305858, 3.402338, 4.49322, 5.578118, 6.656663, 7.728505, 
    8.793312, 9.850773, 10.90059, 11.9425, 12.97624, 14.00158, 15.01831, 
    16.02623, 17.02517, 18.01497, 18.99549, 19.96662, 20.92826, 21.88032, 
    22.82273, 23.75546, 24.67844, 25.59168, 26.49515, 27.38887, 28.27285, 
    29.14713, 30.01174, 30.86674, 31.71219, 32.54816, 33.37472, 34.19197, 35, 
    35.79891, 36.5888, 37.36979,
  303.4273, 304.2095, 305, 305.7989, 306.6063, 307.4223, 308.2469, 309.0802, 
    309.9223, 310.7732, 311.633, 312.5016, 313.3792, 314.2657, 315.1612, 
    316.0655, 316.9788, 317.9009, 318.8319, 319.7716, 320.72, 321.677, 
    322.6425, 323.6163, 324.5984, 325.5886, 326.5867, 327.5925, 328.6058, 
    329.6265, 330.6542, 331.6887, 332.7297, 333.7771, 334.8304, 335.8893, 
    336.9535, 338.0227, 339.0965, 340.1745, 341.2564, 342.3417, 343.43, 
    344.521, 345.6141, 346.709, 347.8053, 348.9024, 350, 351.0976, 352.1947, 
    353.291, 354.3859, 355.479, 356.57, 357.6583, 358.7436, 359.8255, 
    0.9034941, 1.977288, 3.046482, 4.110714, 5.16964, 6.222924, 7.270251, 
    8.311317, 9.345838, 10.37354, 11.39418, 12.40751, 13.41332, 14.4114, 
    15.40157, 16.38366, 17.35752, 18.323, 19.28, 20.2284, 21.16812, 22.09908, 
    23.02121, 23.93448, 24.83885, 25.73429, 26.6208, 27.49838, 28.36704, 
    29.22681, 30.07772, 30.91981, 31.75312, 32.57773, 33.3937, 34.20109, 35, 
    35.7905, 36.57269,
  304.2172, 305, 305.7905, 306.5888, 307.395, 308.209, 309.0311, 309.8612, 
    310.6993, 311.5456, 312.3999, 313.2625, 314.1331, 315.012, 315.8989, 
    316.794, 317.6972, 318.6084, 319.5276, 320.4547, 321.3896, 322.3323, 
    323.2827, 324.2405, 325.2058, 326.1783, 327.1578, 328.1443, 329.1375, 
    330.1371, 331.1431, 332.1551, 333.1729, 334.1963, 335.225, 336.2586, 
    337.297, 338.3397, 339.3865, 340.437, 341.4908, 342.5478, 343.6074, 
    344.6693, 345.7331, 346.7984, 347.865, 348.9323, 350, 351.0677, 352.135, 
    353.2016, 354.2669, 355.3307, 356.3926, 357.4522, 358.5092, 359.563, 
    0.6135356, 1.660314, 2.703033, 3.741373, 4.775022, 5.80368, 6.827063, 
    7.844895, 8.856917, 9.862885, 10.86256, 11.85573, 12.84219, 13.82175, 
    14.79423, 15.75947, 16.71733, 17.66766, 18.61036, 19.54531, 20.47243, 
    21.39162, 22.30283, 23.206, 24.10108, 24.98804, 25.86687, 26.73754, 
    27.60006, 28.45444, 29.30069, 30.13884, 30.96892, 31.79097, 32.60505, 
    33.4112, 34.2095, 35, 35.78278,
  305, 305.7828, 306.5727, 307.3698, 308.1741, 308.9857, 309.8047, 310.6309, 
    311.4646, 312.3057, 313.1541, 314.01, 314.8733, 315.744, 316.6221, 
    317.5075, 318.4002, 319.3002, 320.2073, 321.1216, 322.043, 322.9712, 
    323.9063, 324.8481, 325.7966, 326.7514, 327.7126, 328.6799, 329.6532, 
    330.6322, 331.6168, 332.6068, 333.6019, 334.6019, 335.6065, 336.6156, 
    337.6287, 338.6458, 339.6663, 340.6902, 341.717, 342.7465, 343.7783, 
    344.8122, 345.8477, 346.8846, 347.9225, 348.9611, 350, 351.0389, 
    352.0775, 353.1154, 354.1523, 355.1878, 356.2217, 357.2535, 358.283, 
    359.3098, 0.3336662, 1.354252, 2.371273, 3.384442, 4.393482, 5.398128, 
    6.39812, 7.393215, 8.383177, 9.367781, 10.34682, 11.32008, 12.28739, 
    13.24856, 14.20343, 15.15185, 16.09367, 17.02878, 17.95705, 18.87837, 
    19.79265, 20.69982, 21.59979, 22.49251, 23.37793, 24.256, 25.12669, 
    25.98999, 26.84588, 27.69435, 28.53541, 29.36907, 30.19535, 31.01428, 
    31.82589, 32.63021, 33.42731, 34.21722, 35 ;

 grid_lat =
  -35.26439, -35.62921, -35.98892, -36.34341, -36.69255, -37.03624, 
    -37.37434, -37.70675, -38.03334, -38.354, -38.66859, -38.977, -39.27911, 
    -39.57478, -39.8639, -40.14635, -40.42199, -40.69072, -40.9524, 
    -41.20691, -41.45414, -41.69396, -41.92625, -42.15091, -42.36781, 
    -42.57683, -42.77788, -42.97084, -43.1556, -43.33206, -43.50012, 
    -43.65969, -43.81068, -43.95298, -44.08652, -44.21122, -44.32701, 
    -44.4338, -44.53154, -44.62016, -44.6996, -44.76982, -44.83077, 
    -44.88241, -44.9247, -44.95763, -44.98116, -44.99529, -45, -44.99529, 
    -44.98116, -44.95763, -44.9247, -44.88241, -44.83077, -44.76982, 
    -44.6996, -44.62016, -44.53154, -44.4338, -44.32701, -44.21122, 
    -44.08652, -43.95298, -43.81068, -43.65969, -43.50012, -43.33206, 
    -43.1556, -42.97084, -42.77788, -42.57683, -42.36781, -42.15091, 
    -41.92625, -41.69396, -41.45414, -41.20691, -40.9524, -40.69072, 
    -40.42199, -40.14635, -39.8639, -39.57478, -39.27911, -38.977, -38.66859, 
    -38.354, -38.03334, -37.70675, -37.37434, -37.03624, -36.69255, 
    -36.34341, -35.98892, -35.62921, -35.26439,
  -35.62921, -36.00579, -36.37735, -36.74377, -37.10492, -37.46067, 
    -37.81089, -38.15546, -38.49422, -38.82706, -39.15382, -39.47439, 
    -39.78861, -40.09635, -40.39747, -40.69183, -40.97929, -41.25971, 
    -41.53295, -41.79888, -42.05735, -42.30823, -42.55138, -42.78666, 
    -43.01395, -43.23311, -43.44402, -43.64655, -43.84056, -44.02596, 
    -44.20261, -44.37041, -44.52925, -44.67902, -44.81961, -44.95095, 
    -45.07294, -45.18549, -45.28852, -45.38197, -45.46576, -45.53984, 
    -45.60415, -45.65865, -45.7033, -45.73805, -45.7629, -45.77781, 
    -45.78278, -45.77781, -45.7629, -45.73805, -45.7033, -45.65865, 
    -45.60415, -45.53984, -45.46576, -45.38197, -45.28852, -45.18549, 
    -45.07294, -44.95095, -44.81961, -44.67902, -44.52925, -44.37041, 
    -44.20261, -44.02596, -43.84056, -43.64655, -43.44402, -43.23311, 
    -43.01395, -42.78666, -42.55138, -42.30823, -42.05735, -41.79888, 
    -41.53295, -41.25971, -40.97929, -40.69183, -40.39747, -40.09635, 
    -39.78861, -39.47439, -39.15382, -38.82706, -38.49422, -38.15546, 
    -37.81089, -37.46067, -37.10492, -36.74377, -36.37735, -36.00579, 
    -35.62921,
  -35.98892, -36.37735, -36.76087, -37.13935, -37.51265, -37.88063, 
    -38.24314, -38.60004, -38.95119, -39.29642, -39.6356, -39.96857, 
    -40.29517, -40.61526, -40.92867, -41.23525, -41.53484, -41.82729, 
    -42.11243, -42.39012, -42.66019, -42.92249, -43.17686, -43.42315, 
    -43.66121, -43.89089, -44.11203, -44.3245, -44.52815, -44.72285, 
    -44.90845, -45.08484, -45.25187, -45.40944, -45.55742, -45.6957, 
    -45.82418, -45.94276, -46.05135, -46.14986, -46.23822, -46.31635, 
    -46.38419, -46.44169, -46.4888, -46.52548, -46.5517, -46.56744, 
    -46.57269, -46.56744, -46.5517, -46.52548, -46.4888, -46.44169, 
    -46.38419, -46.31635, -46.23822, -46.14986, -46.05135, -45.94276, 
    -45.82418, -45.6957, -45.55742, -45.40944, -45.25187, -45.08484, 
    -44.90845, -44.72285, -44.52815, -44.3245, -44.11203, -43.89089, 
    -43.66121, -43.42315, -43.17686, -42.92249, -42.66019, -42.39012, 
    -42.11243, -41.82729, -41.53484, -41.23525, -40.92867, -40.61526, 
    -40.29517, -39.96857, -39.6356, -39.29642, -38.95119, -38.60004, 
    -38.24314, -37.88063, -37.51265, -37.13935, -36.76087, -36.37735, 
    -35.98892,
  -36.34341, -36.74377, -37.13935, -37.53001, -37.91559, -38.29594, 
    -38.67091, -39.04033, -39.40405, -39.7619, -40.11372, -40.45934, 
    -40.79858, -41.13129, -41.45728, -41.77639, -42.08843, -42.39323, 
    -42.69062, -42.98042, -43.26245, -43.53653, -43.8025, -44.06018, 
    -44.30939, -44.54997, -44.78174, -45.00454, -45.21821, -45.42259, 
    -45.61752, -45.80286, -45.97845, -46.14417, -46.29986, -46.4454, 
    -46.58068, -46.70559, -46.82, -46.92382, -47.01697, -47.09935, -47.17091, 
    -47.23156, -47.28126, -47.31997, -47.34763, -47.36425, -47.36979, 
    -47.36425, -47.34763, -47.31997, -47.28126, -47.23156, -47.17091, 
    -47.09935, -47.01697, -46.92382, -46.82, -46.70559, -46.58068, -46.4454, 
    -46.29986, -46.14417, -45.97845, -45.80286, -45.61752, -45.42259, 
    -45.21821, -45.00454, -44.78174, -44.54997, -44.30939, -44.06018, 
    -43.8025, -43.53653, -43.26245, -42.98042, -42.69062, -42.39323, 
    -42.08843, -41.77639, -41.45728, -41.13129, -40.79858, -40.45934, 
    -40.11372, -39.7619, -39.40405, -39.04033, -38.67091, -38.29594, 
    -37.91559, -37.53001, -37.13935, -36.74377, -36.34341,
  -36.69255, -37.10492, -37.51265, -37.91559, -38.31358, -38.70644, 
    -39.09401, -39.47613, -39.85261, -40.22328, -40.58796, -40.94647, 
    -41.29861, -41.64421, -41.98307, -42.315, -42.6398, -42.95729, -43.26726, 
    -43.56952, -43.86388, -44.15013, -44.42807, -44.69753, -44.95829, 
    -45.21016, -45.45296, -45.68649, -45.91058, -46.12503, -46.32969, 
    -46.52436, -46.70888, -46.8831, -47.04686, -47.20001, -47.34241, 
    -47.47393, -47.59445, -47.70385, -47.80202, -47.88887, -47.96432, 
    -48.02829, -48.08072, -48.12155, -48.15074, -48.16827, -48.17411, 
    -48.16827, -48.15074, -48.12155, -48.08072, -48.02829, -47.96432, 
    -47.88887, -47.80202, -47.70385, -47.59445, -47.47393, -47.34241, 
    -47.20001, -47.04686, -46.8831, -46.70888, -46.52436, -46.32969, 
    -46.12503, -45.91058, -45.68649, -45.45296, -45.21016, -44.95829, 
    -44.69753, -44.42807, -44.15013, -43.86388, -43.56952, -43.26726, 
    -42.95729, -42.6398, -42.315, -41.98307, -41.64421, -41.29861, -40.94647, 
    -40.58796, -40.22328, -39.85261, -39.47613, -39.09401, -38.70644, 
    -38.31358, -37.91559, -37.51265, -37.10492, -36.69255,
  -37.03624, -37.46067, -37.88063, -38.29594, -38.70644, -39.11194, 
    -39.51227, -39.90724, -40.29666, -40.68035, -41.0581, -41.42973, 
    -41.79502, -42.15377, -42.50578, -42.85083, -43.18871, -43.51921, 
    -43.84211, -44.15719, -44.46423, -44.76302, -45.05334, -45.33495, 
    -45.60766, -45.87124, -46.12547, -46.37015, -46.60506, -46.83001, 
    -47.04478, -47.24918, -47.44304, -47.62614, -47.79833, -47.95944, 
    -48.10929, -48.24775, -48.37467, -48.48992, -48.59336, -48.68491, 
    -48.76445, -48.83191, -48.8872, -48.93027, -48.96106, -48.97956, 
    -48.98572, -48.97956, -48.96106, -48.93027, -48.8872, -48.83191, 
    -48.76445, -48.68491, -48.59336, -48.48992, -48.37467, -48.24775, 
    -48.10929, -47.95944, -47.79833, -47.62614, -47.44304, -47.24918, 
    -47.04478, -46.83001, -46.60506, -46.37015, -46.12547, -45.87124, 
    -45.60766, -45.33495, -45.05334, -44.76302, -44.46423, -44.15719, 
    -43.84211, -43.51921, -43.18871, -42.85083, -42.50578, -42.15377, 
    -41.79502, -41.42973, -41.0581, -40.68035, -40.29666, -39.90724, 
    -39.51227, -39.11194, -38.70644, -38.29594, -37.88063, -37.46067, 
    -37.03624,
  -37.37434, -37.81089, -38.24314, -38.67091, -39.09401, -39.51227, 
    -39.92548, -40.33345, -40.73598, -41.13287, -41.52391, -41.90887, 
    -42.28755, -42.65972, -43.02515, -43.38362, -43.73489, -44.07872, 
    -44.41489, -44.74314, -45.06325, -45.37495, -45.67802, -45.97221, 
    -46.25727, -46.53297, -46.79906, -47.05531, -47.30147, -47.53732, 
    -47.76263, -47.97718, -48.18076, -48.37315, -48.55416, -48.72359, 
    -48.88126, -49.02699, -49.16062, -49.282, -49.39099, -49.48746, 
    -49.57131, -49.64243, -49.70073, -49.74615, -49.77864, -49.79815, 
    -49.80465, -49.79815, -49.77864, -49.74615, -49.70073, -49.64243, 
    -49.57131, -49.48746, -49.39099, -49.282, -49.16062, -49.02699, 
    -48.88126, -48.72359, -48.55416, -48.37315, -48.18076, -47.97718, 
    -47.76263, -47.53732, -47.30147, -47.05531, -46.79906, -46.53297, 
    -46.25727, -45.97221, -45.67802, -45.37495, -45.06325, -44.74314, 
    -44.41489, -44.07872, -43.73489, -43.38362, -43.02515, -42.65972, 
    -42.28755, -41.90887, -41.52391, -41.13287, -40.73598, -40.33345, 
    -39.92548, -39.51227, -39.09401, -38.67091, -38.24314, -37.81089, 
    -37.37434,
  -37.70675, -38.15546, -38.60004, -39.04033, -39.47613, -39.90724, 
    -40.33345, -40.75457, -41.17037, -41.58063, -41.98514, -42.38366, 
    -42.77596, -43.16179, -43.54091, -43.91308, -44.27805, -44.63554, 
    -44.98531, -45.3271, -45.66063, -45.98564, -46.30186, -46.60902, 
    -46.90686, -47.1951, -47.47348, -47.74172, -47.99957, -48.24677, 
    -48.48305, -48.70818, -48.92191, -49.124, -49.31422, -49.49236, -49.6582, 
    -49.81155, -49.95222, -50.08005, -50.19486, -50.29652, -50.38489, 
    -50.45986, -50.52134, -50.56924, -50.6035, -50.62407, -50.63093, 
    -50.62407, -50.6035, -50.56924, -50.52134, -50.45986, -50.38489, 
    -50.29652, -50.19486, -50.08005, -49.95222, -49.81155, -49.6582, 
    -49.49236, -49.31422, -49.124, -48.92191, -48.70818, -48.48305, 
    -48.24677, -47.99957, -47.74172, -47.47348, -47.1951, -46.90686, 
    -46.60902, -46.30186, -45.98564, -45.66063, -45.3271, -44.98531, 
    -44.63554, -44.27805, -43.91308, -43.54091, -43.16179, -42.77596, 
    -42.38366, -41.98514, -41.58063, -41.17037, -40.75457, -40.33345, 
    -39.90724, -39.47613, -39.04033, -38.60004, -38.15546, -37.70675,
  -38.03334, -38.49422, -38.95119, -39.40405, -39.85261, -40.29666, 
    -40.73598, -41.17037, -41.59958, -42.02338, -42.44154, -42.85382, 
    -43.25996, -43.6597, -44.05278, -44.43893, -44.81789, -45.18936, 
    -45.55307, -45.90874, -46.25607, -46.59477, -46.92454, -47.24509, 
    -47.55613, -47.85734, -48.14844, -48.42913, -48.69912, -48.95811, 
    -49.20582, -49.44197, -49.66629, -49.8785, -50.07836, -50.26561, 
    -50.44002, -50.60136, -50.74942, -50.88401, -51.00494, -51.11204, 
    -51.20517, -51.2842, -51.34902, -51.39953, -51.43566, -51.45736, 
    -51.46459, -51.45736, -51.43566, -51.39953, -51.34902, -51.2842, 
    -51.20517, -51.11204, -51.00494, -50.88401, -50.74942, -50.60136, 
    -50.44002, -50.26561, -50.07836, -49.8785, -49.66629, -49.44197, 
    -49.20582, -48.95811, -48.69912, -48.42913, -48.14844, -47.85734, 
    -47.55613, -47.24509, -46.92454, -46.59477, -46.25607, -45.90874, 
    -45.55307, -45.18936, -44.81789, -44.43893, -44.05278, -43.6597, 
    -43.25996, -42.85382, -42.44154, -42.02338, -41.59958, -41.17037, 
    -40.73598, -40.29666, -39.85261, -39.40405, -38.95119, -38.49422, 
    -38.03334,
  -38.354, -38.82706, -39.29642, -39.7619, -40.22328, -40.68035, -41.13287, 
    -41.58063, -42.02338, -42.46088, -42.89287, -43.31909, -43.73928, 
    -44.15316, -44.56044, -44.96085, -45.35409, -45.73986, -46.11785, 
    -46.48775, -46.84925, -47.20202, -47.54575, -47.8801, -48.20476, 
    -48.51939, -48.82367, -49.11726, -49.39985, -49.6711, -49.9307, 
    -50.17833, -50.4137, -50.63649, -50.84642, -51.04321, -51.22659, 
    -51.39631, -51.55212, -51.69381, -51.82117, -51.934, -52.03214, 
    -52.11544, -52.18378, -52.23703, -52.27514, -52.29802, -52.30565, 
    -52.29802, -52.27514, -52.23703, -52.18378, -52.11544, -52.03214, 
    -51.934, -51.82117, -51.69381, -51.55212, -51.39631, -51.22659, 
    -51.04321, -50.84642, -50.63649, -50.4137, -50.17833, -49.9307, -49.6711, 
    -49.39985, -49.11726, -48.82367, -48.51939, -48.20476, -47.8801, 
    -47.54575, -47.20202, -46.84925, -46.48775, -46.11785, -45.73986, 
    -45.35409, -44.96085, -44.56044, -44.15316, -43.73928, -43.31909, 
    -42.89287, -42.46088, -42.02338, -41.58063, -41.13287, -40.68035, 
    -40.22328, -39.7619, -39.29642, -38.82706, -38.354,
  -38.66859, -39.15382, -39.6356, -40.11372, -40.58796, -41.0581, -41.52391, 
    -41.98514, -42.44154, -42.89287, -43.33884, -43.77919, -44.21362, 
    -44.64186, -45.0636, -45.47853, -45.88634, -46.28671, -46.67929, 
    -47.06378, -47.43981, -47.80704, -48.16513, -48.51371, -48.85243, 
    -49.18093, -49.49884, -49.8058, -50.10146, -50.38545, -50.65742, 
    -50.91702, -51.1639, -51.39774, -51.6182, -51.82498, -52.01776, 
    -52.19627, -52.36022, -52.50938, -52.64349, -52.76235, -52.86576, 
    -52.95356, -53.0256, -53.08176, -53.12194, -53.14607, -53.15412, 
    -53.14607, -53.12194, -53.08176, -53.0256, -52.95356, -52.86576, 
    -52.76235, -52.64349, -52.50938, -52.36022, -52.19627, -52.01776, 
    -51.82498, -51.6182, -51.39774, -51.1639, -50.91702, -50.65742, 
    -50.38545, -50.10146, -49.8058, -49.49884, -49.18093, -48.85243, 
    -48.51371, -48.16513, -47.80704, -47.43981, -47.06378, -46.67929, 
    -46.28671, -45.88634, -45.47853, -45.0636, -44.64186, -44.21362, 
    -43.77919, -43.33884, -42.89287, -42.44154, -41.98514, -41.52391, 
    -41.0581, -40.58796, -40.11372, -39.6356, -39.15382, -38.66859,
  -38.977, -39.47439, -39.96857, -40.45934, -40.94647, -41.42973, -41.90887, 
    -42.38366, -42.85382, -43.31909, -43.77919, -44.23382, -44.68269, 
    -45.1255, -45.56192, -45.99162, -46.41428, -46.82954, -47.23705, 
    -47.63646, -48.02739, -48.40947, -48.78232, -49.14555, -49.49877, 
    -49.84158, -50.1736, -50.49441, -50.80363, -51.10085, -51.38569, 
    -51.65775, -51.91666, -52.16203, -52.39351, -52.61073, -52.81337, 
    -53.00109, -53.17359, -53.33059, -53.47181, -53.59702, -53.70599, 
    -53.79853, -53.87448, -53.93369, -53.97606, -54.00152, -54.01001, 
    -54.00152, -53.97606, -53.93369, -53.87448, -53.79853, -53.70599, 
    -53.59702, -53.47181, -53.33059, -53.17359, -53.00109, -52.81337, 
    -52.61073, -52.39351, -52.16203, -51.91666, -51.65775, -51.38569, 
    -51.10085, -50.80363, -50.49441, -50.1736, -49.84158, -49.49877, 
    -49.14555, -48.78232, -48.40947, -48.02739, -47.63646, -47.23705, 
    -46.82954, -46.41428, -45.99162, -45.56192, -45.1255, -44.68269, 
    -44.23382, -43.77919, -43.31909, -42.85382, -42.38366, -41.90887, 
    -41.42973, -40.94647, -40.45934, -39.96857, -39.47439, -38.977,
  -39.27911, -39.78861, -40.29517, -40.79858, -41.29861, -41.79502, 
    -42.28755, -42.77596, -43.25996, -43.73928, -44.21362, -44.68269, 
    -45.14617, -45.60374, -46.05505, -46.49977, -46.93754, -47.36799, 
    -47.79074, -48.20541, -48.6116, -49.00891, -49.39692, -49.77522, 
    -50.14338, -50.50098, -50.84757, -51.18272, -51.506, -51.81697, 
    -52.11519, -52.40023, -52.67167, -52.92909, -53.17208, -53.40025, 
    -53.61321, -53.81061, -53.99209, -54.15733, -54.30604, -54.43793, 
    -54.55275, -54.6503, -54.73037, -54.79281, -54.8375, -54.86435, 
    -54.87331, -54.86435, -54.8375, -54.79281, -54.73037, -54.6503, 
    -54.55275, -54.43793, -54.30604, -54.15733, -53.99209, -53.81061, 
    -53.61321, -53.40025, -53.17208, -52.92909, -52.67167, -52.40023, 
    -52.11519, -51.81697, -51.506, -51.18272, -50.84757, -50.50098, 
    -50.14338, -49.77522, -49.39692, -49.00891, -48.6116, -48.20541, 
    -47.79074, -47.36799, -46.93754, -46.49977, -46.05505, -45.60374, 
    -45.14617, -44.68269, -44.21362, -43.73928, -43.25996, -42.77596, 
    -42.28755, -41.79502, -41.29861, -40.79858, -40.29517, -39.78861, 
    -39.27911,
  -39.57478, -40.09635, -40.61526, -41.13129, -41.64421, -42.15377, 
    -42.65972, -43.16179, -43.6597, -44.15316, -44.64186, -45.1255, 
    -45.60374, -46.07624, -46.54266, -47.00262, -47.45575, -47.90166, 
    -48.33995, -48.77021, -49.19202, -49.60493, -50.00851, -50.40231, 
    -50.78586, -51.1587, -51.52035, -51.87035, -52.2082, -52.53343, 
    -52.84557, -53.14412, -53.42863, -53.69863, -53.95366, -54.19329, 
    -54.41708, -54.62463, -54.81555, -54.98947, -55.14605, -55.28499, 
    -55.40599, -55.50881, -55.59324, -55.65909, -55.70623, -55.73455, 
    -55.744, -55.73455, -55.70623, -55.65909, -55.59324, -55.50881, 
    -55.40599, -55.28499, -55.14605, -54.98947, -54.81555, -54.62463, 
    -54.41708, -54.19329, -53.95366, -53.69863, -53.42863, -53.14412, 
    -52.84557, -52.53343, -52.2082, -51.87035, -51.52035, -51.1587, 
    -50.78586, -50.40231, -50.00851, -49.60493, -49.19202, -48.77021, 
    -48.33995, -47.90166, -47.45575, -47.00262, -46.54266, -46.07624, 
    -45.60374, -45.1255, -44.64186, -44.15316, -43.6597, -43.16179, 
    -42.65972, -42.15377, -41.64421, -41.13129, -40.61526, -40.09635, 
    -39.57478,
  -39.8639, -40.39747, -40.92867, -41.45728, -41.98307, -42.50578, -43.02515, 
    -43.54091, -44.05278, -44.56044, -45.0636, -45.56192, -46.05505, 
    -46.54266, -47.02436, -47.49977, -47.96851, -48.43015, -48.88427, 
    -49.33044, -49.7682, -50.19709, -50.61664, -51.02636, -51.42574, 
    -51.8143, -52.1915, -52.55685, -52.9098, -53.24984, -53.57643, -53.88906, 
    -54.18719, -54.47033, -54.73795, -54.98958, -55.22473, -55.44294, 
    -55.64378, -55.82684, -55.99172, -56.13808, -56.26561, -56.374, 
    -56.46303, -56.53249, -56.58222, -56.6121, -56.62207, -56.6121, 
    -56.58222, -56.53249, -56.46303, -56.374, -56.26561, -56.13808, 
    -55.99172, -55.82684, -55.64378, -55.44294, -55.22473, -54.98958, 
    -54.73795, -54.47033, -54.18719, -53.88906, -53.57643, -53.24984, 
    -52.9098, -52.55685, -52.1915, -51.8143, -51.42574, -51.02636, -50.61664, 
    -50.19709, -49.7682, -49.33044, -48.88427, -48.43015, -47.96851, 
    -47.49977, -47.02436, -46.54266, -46.05505, -45.56192, -45.0636, 
    -44.56044, -44.05278, -43.54091, -43.02515, -42.50578, -41.98307, 
    -41.45728, -40.92867, -40.39747, -39.8639,
  -40.14635, -40.69183, -41.23525, -41.77639, -42.315, -42.85083, -43.38362, 
    -43.91308, -44.43893, -44.96085, -45.47853, -45.99162, -46.49977, 
    -47.00262, -47.49977, -47.99084, -48.4754, -48.95301, -49.42325, 
    -49.88563, -50.33969, -50.78492, -51.22083, -51.64688, -52.06255, 
    -52.46729, -52.86054, -53.24175, -53.61034, -53.96573, -54.30735, 
    -54.63462, -54.94697, -55.24382, -55.52462, -55.78882, -56.03588, 
    -56.26529, -56.47657, -56.66924, -56.84288, -56.99708, -57.13149, 
    -57.24578, -57.33968, -57.41296, -57.46543, -57.49697, -57.50749, 
    -57.49697, -57.46543, -57.41296, -57.33968, -57.24578, -57.13149, 
    -56.99708, -56.84288, -56.66924, -56.47657, -56.26529, -56.03588, 
    -55.78882, -55.52462, -55.24382, -54.94697, -54.63462, -54.30735, 
    -53.96573, -53.61034, -53.24175, -52.86054, -52.46729, -52.06255, 
    -51.64688, -51.22083, -50.78492, -50.33969, -49.88563, -49.42325, 
    -48.95301, -48.4754, -47.99084, -47.49977, -47.00262, -46.49977, 
    -45.99162, -45.47853, -44.96085, -44.43893, -43.91308, -43.38362, 
    -42.85083, -42.315, -41.77639, -41.23525, -40.69183, -40.14635,
  -40.42199, -40.97929, -41.53484, -42.08843, -42.6398, -43.18871, -43.73489, 
    -44.27805, -44.81789, -45.35409, -45.88634, -46.41428, -46.93754, 
    -47.45575, -47.96851, -48.4754, -48.97598, -49.46981, -49.95642, 
    -50.43531, -50.90599, -51.36792, -51.82056, -52.26337, -52.69576, 
    -53.11716, -53.52696, -53.92455, -54.30932, -54.68064, -55.03786, 
    -55.38037, -55.70753, -56.01871, -56.31329, -56.59066, -56.85022, 
    -57.09141, -57.31367, -57.51648, -57.69935, -57.86184, -58.00352, 
    -58.12405, -58.22311, -58.30043, -58.35581, -58.3891, -58.40021, 
    -58.3891, -58.35581, -58.30043, -58.22311, -58.12405, -58.00352, 
    -57.86184, -57.69935, -57.51648, -57.31367, -57.09141, -56.85022, 
    -56.59066, -56.31329, -56.01871, -55.70753, -55.38037, -55.03786, 
    -54.68064, -54.30932, -53.92455, -53.52696, -53.11716, -52.69576, 
    -52.26337, -51.82056, -51.36792, -50.90599, -50.43531, -49.95642, 
    -49.46981, -48.97598, -48.4754, -47.96851, -47.45575, -46.93754, 
    -46.41428, -45.88634, -45.35409, -44.81789, -44.27805, -43.73489, 
    -43.18871, -42.6398, -42.08843, -41.53484, -40.97929, -40.42199,
  -40.69072, -41.25971, -41.82729, -42.39323, -42.95729, -43.51921, 
    -44.07872, -44.63554, -45.18936, -45.73986, -46.28671, -46.82954, 
    -47.36799, -47.90166, -48.43015, -48.95301, -49.46981, -49.98007, 
    -50.48329, -50.97897, -51.46657, -51.94554, -52.4153, -52.87527, 
    -53.32483, -53.76335, -54.1902, -54.60471, -55.00621, -55.39402, 
    -55.76746, -56.12582, -56.46842, -56.79456, -57.10355, -57.39472, 
    -57.66741, -57.92097, -58.1548, -58.36829, -58.56092, -58.73216, 
    -58.88156, -59.0087, -59.11322, -59.19484, -59.2533, -59.28845, 
    -59.30018, -59.28845, -59.2533, -59.19484, -59.11322, -59.0087, 
    -58.88156, -58.73216, -58.56092, -58.36829, -58.1548, -57.92097, 
    -57.66741, -57.39472, -57.10355, -56.79456, -56.46842, -56.12582, 
    -55.76746, -55.39402, -55.00621, -54.60471, -54.1902, -53.76335, 
    -53.32483, -52.87527, -52.4153, -51.94554, -51.46657, -50.97897, 
    -50.48329, -49.98007, -49.46981, -48.95301, -48.43015, -47.90166, 
    -47.36799, -46.82954, -46.28671, -45.73986, -45.18936, -44.63554, 
    -44.07872, -43.51921, -42.95729, -42.39323, -41.82729, -41.25971, 
    -40.69072,
  -40.9524, -41.53295, -42.11243, -42.69062, -43.26726, -43.84211, -44.41489, 
    -44.98531, -45.55307, -46.11785, -46.67929, -47.23705, -47.79074, 
    -48.33995, -48.88427, -49.42325, -49.95642, -50.48329, -51.00336, 
    -51.51608, -52.0209, -52.51723, -53.00447, -53.48199, -53.94915, 
    -54.40527, -54.84966, -55.28162, -55.70042, -56.10532, -56.49557, 
    -56.87043, -57.22911, -57.57087, -57.89494, -58.20058, -58.48705, 
    -58.75364, -58.99965, -59.22443, -59.42736, -59.60787, -59.76543, 
    -59.89958, -60.00991, -60.09608, -60.15783, -60.19496, -60.20734, 
    -60.19496, -60.15783, -60.09608, -60.00991, -59.89958, -59.76543, 
    -59.60787, -59.42736, -59.22443, -58.99965, -58.75364, -58.48705, 
    -58.20058, -57.89494, -57.57087, -57.22911, -56.87043, -56.49557, 
    -56.10532, -55.70042, -55.28162, -54.84966, -54.40527, -53.94915, 
    -53.48199, -53.00447, -52.51723, -52.0209, -51.51608, -51.00336, 
    -50.48329, -49.95642, -49.42325, -48.88427, -48.33995, -47.79074, 
    -47.23705, -46.67929, -46.11785, -45.55307, -44.98531, -44.41489, 
    -43.84211, -43.26726, -42.69062, -42.11243, -41.53295, -40.9524,
  -41.20691, -41.79888, -42.39012, -42.98042, -43.56952, -44.15719, 
    -44.74314, -45.3271, -45.90874, -46.48775, -47.06378, -47.63646, 
    -48.20541, -48.77021, -49.33044, -49.88563, -50.43531, -50.97897, 
    -51.51608, -52.04608, -52.56838, -53.08239, -53.58745, -54.08292, 
    -54.5681, -55.04227, -55.50471, -55.95465, -56.39131, -56.8139, -57.2216, 
    -57.61359, -57.98904, -58.34711, -58.68696, -59.00777, -59.30871, 
    -59.589, -59.84786, -60.08456, -60.29839, -60.48872, -60.65495, 
    -60.79654, -60.91304, -61.00407, -61.06931, -61.10854, -61.12163, 
    -61.10854, -61.06931, -61.00407, -60.91304, -60.79654, -60.65495, 
    -60.48872, -60.29839, -60.08456, -59.84786, -59.589, -59.30871, 
    -59.00777, -58.68696, -58.34711, -57.98904, -57.61359, -57.2216, 
    -56.8139, -56.39131, -55.95465, -55.50471, -55.04227, -54.5681, 
    -54.08292, -53.58745, -53.08239, -52.56838, -52.04608, -51.51608, 
    -50.97897, -50.43531, -49.88563, -49.33044, -48.77021, -48.20541, 
    -47.63646, -47.06378, -46.48775, -45.90874, -45.3271, -44.74314, 
    -44.15719, -43.56952, -42.98042, -42.39012, -41.79888, -41.20691,
  -41.45414, -42.05735, -42.66019, -43.26245, -43.86388, -44.46423, 
    -45.06325, -45.66063, -46.25607, -46.84925, -47.43981, -48.02739, 
    -48.6116, -49.19202, -49.7682, -50.33969, -50.90599, -51.46657, -52.0209, 
    -52.56838, -53.10843, -53.64039, -54.16361, -54.67738, -55.18099, 
    -55.67367, -56.15464, -56.62309, -57.07819, -57.51908, -57.94487, 
    -58.35467, -58.74758, -59.12267, -59.47903, -59.81574, -60.1319, 
    -60.42662, -60.69904, -60.94834, -61.17372, -61.37446, -61.54989, 
    -61.6994, -61.82248, -61.91867, -61.98763, -62.02911, -62.04295, 
    -62.02911, -61.98763, -61.91867, -61.82248, -61.6994, -61.54989, 
    -61.37446, -61.17372, -60.94834, -60.69904, -60.42662, -60.1319, 
    -59.81574, -59.47903, -59.12267, -58.74758, -58.35467, -57.94487, 
    -57.51908, -57.07819, -56.62309, -56.15464, -55.67367, -55.18099, 
    -54.67738, -54.16361, -53.64039, -53.10843, -52.56838, -52.0209, 
    -51.46657, -50.90599, -50.33969, -49.7682, -49.19202, -48.6116, 
    -48.02739, -47.43981, -46.84925, -46.25607, -45.66063, -45.06325, 
    -44.46423, -43.86388, -43.26245, -42.66019, -42.05735, -41.45414,
  -41.69396, -42.30823, -42.92249, -43.53653, -44.15013, -44.76302, 
    -45.37495, -45.98564, -46.59477, -47.20202, -47.80704, -48.40947, 
    -49.00891, -49.60493, -50.19709, -50.78492, -51.36792, -51.94554, 
    -52.51723, -53.08239, -53.64039, -54.19058, -54.73225, -55.26468, 
    -55.78711, -56.29873, -56.79872, -57.28621, -57.76032, -58.22011, 
    -58.66464, -59.09295, -59.50403, -59.89689, -60.27053, -60.62392, 
    -60.95608, -61.26601, -61.55275, -61.81537, -62.05299, -62.26479, 
    -62.45001, -62.60796, -62.73804, -62.83975, -62.91269, -62.95657, 
    -62.97122, -62.95657, -62.91269, -62.83975, -62.73804, -62.60796, 
    -62.45001, -62.26479, -62.05299, -61.81537, -61.55275, -61.26601, 
    -60.95608, -60.62392, -60.27053, -59.89689, -59.50403, -59.09295, 
    -58.66464, -58.22011, -57.76032, -57.28621, -56.79872, -56.29873, 
    -55.78711, -55.26468, -54.73225, -54.19058, -53.64039, -53.08239, 
    -52.51723, -51.94554, -51.36792, -50.78492, -50.19709, -49.60493, 
    -49.00891, -48.40947, -47.80704, -47.20202, -46.59477, -45.98564, 
    -45.37495, -44.76302, -44.15013, -43.53653, -42.92249, -42.30823, 
    -41.69396,
  -41.92625, -42.55138, -43.17686, -43.8025, -44.42807, -45.05334, -45.67802, 
    -46.30186, -46.92454, -47.54575, -48.16513, -48.78232, -49.39692, 
    -50.00851, -50.61664, -51.22083, -51.82056, -52.4153, -53.00447, 
    -53.58745, -54.16361, -54.73225, -55.29266, -55.84407, -56.38568, 
    -56.91667, -57.43615, -57.9432, -58.43688, -58.9162, -59.38013, 
    -59.82764, -60.25764, -60.66905, -61.06076, -61.43166, -61.78063, 
    -62.10659, -62.40846, -62.6852, -62.93583, -63.15939, -63.35503, 
    -63.52198, -63.65955, -63.76716, -63.84436, -63.89082, -63.90633, 
    -63.89082, -63.84436, -63.76716, -63.65955, -63.52198, -63.35503, 
    -63.15939, -62.93583, -62.6852, -62.40846, -62.10659, -61.78063, 
    -61.43166, -61.06076, -60.66905, -60.25764, -59.82764, -59.38013, 
    -58.9162, -58.43688, -57.9432, -57.43615, -56.91667, -56.38568, 
    -55.84407, -55.29266, -54.73225, -54.16361, -53.58745, -53.00447, 
    -52.4153, -51.82056, -51.22083, -50.61664, -50.00851, -49.39692, 
    -48.78232, -48.16513, -47.54575, -46.92454, -46.30186, -45.67802, 
    -45.05334, -44.42807, -43.8025, -43.17686, -42.55138, -41.92625,
  -42.15091, -42.78666, -43.42315, -44.06018, -44.69753, -45.33495, 
    -45.97221, -46.60902, -47.24509, -47.8801, -48.51371, -49.14555, 
    -49.77522, -50.40231, -51.02636, -51.64688, -52.26337, -52.87527, 
    -53.48199, -54.08292, -54.67738, -55.26468, -55.84407, -56.41476, 
    -56.97591, -57.52666, -58.06607, -58.59319, -59.10701, -59.60646, 
    -60.09047, -60.55789, -61.00757, -61.43833, -61.84895, -62.2382, 
    -62.60488, -62.94775, -63.26563, -63.55734, -63.82177, -64.05786, 
    -64.26463, -64.4412, -64.58678, -64.70073, -64.7825, -64.83172, 
    -64.84815, -64.83172, -64.7825, -64.70073, -64.58678, -64.4412, 
    -64.26463, -64.05786, -63.82177, -63.55734, -63.26563, -62.94775, 
    -62.60488, -62.2382, -61.84895, -61.43833, -61.00757, -60.55789, 
    -60.09047, -59.60646, -59.10701, -58.59319, -58.06607, -57.52666, 
    -56.97591, -56.41476, -55.84407, -55.26468, -54.67738, -54.08292, 
    -53.48199, -52.87527, -52.26337, -51.64688, -51.02636, -50.40231, 
    -49.77522, -49.14555, -48.51371, -47.8801, -47.24509, -46.60902, 
    -45.97221, -45.33495, -44.69753, -44.06018, -43.42315, -42.78666, 
    -42.15091,
  -42.36781, -43.01395, -43.66121, -44.30939, -44.95829, -45.60766, 
    -46.25727, -46.90686, -47.55613, -48.20476, -48.85243, -49.49877, 
    -50.14338, -50.78586, -51.42574, -52.06255, -52.69576, -53.32483, 
    -53.94915, -54.5681, -55.18099, -55.78711, -56.38568, -56.97591, 
    -57.55692, -58.1278, -58.68758, -59.23526, -59.76975, -60.28995, 
    -60.79469, -61.28276, -61.7529, -62.20383, -62.63423, -63.04275, 
    -63.42805, -63.78878, -64.1236, -64.4312, -64.71033, -64.95979, 
    -65.17846, -65.36533, -65.51952, -65.64027, -65.72695, -65.77914, 
    -65.79657, -65.77914, -65.72695, -65.64027, -65.51952, -65.36533, 
    -65.17846, -64.95979, -64.71033, -64.4312, -64.1236, -63.78878, 
    -63.42805, -63.04275, -62.63423, -62.20383, -61.7529, -61.28276, 
    -60.79469, -60.28995, -59.76975, -59.23526, -58.68758, -58.1278, 
    -57.55692, -56.97591, -56.38568, -55.78711, -55.18099, -54.5681, 
    -53.94915, -53.32483, -52.69576, -52.06255, -51.42574, -50.78586, 
    -50.14338, -49.49877, -48.85243, -48.20476, -47.55613, -46.90686, 
    -46.25727, -45.60766, -44.95829, -44.30939, -43.66121, -43.01395, 
    -42.36781,
  -42.57683, -43.23311, -43.89089, -44.54997, -45.21016, -45.87124, 
    -46.53297, -47.1951, -47.85734, -48.51939, -49.18093, -49.84158, 
    -50.50098, -51.1587, -51.8143, -52.46729, -53.11716, -53.76335, 
    -54.40527, -55.04227, -55.67367, -56.29873, -56.91667, -57.52666, 
    -58.1278, -58.71915, -59.2997, -59.86839, -60.4241, -60.96564, -61.49178, 
    -62.00122, -62.49262, -62.96457, -63.41565, -63.84439, -64.2493, 
    -64.62888, -64.98164, -65.30614, -65.60093, -65.86467, -66.09609, 
    -66.29404, -66.45748, -66.58555, -66.67754, -66.73294, -66.75144, 
    -66.73294, -66.67754, -66.58555, -66.45748, -66.29404, -66.09609, 
    -65.86467, -65.60093, -65.30614, -64.98164, -64.62888, -64.2493, 
    -63.84439, -63.41565, -62.96457, -62.49262, -62.00122, -61.49178, 
    -60.96564, -60.4241, -59.86839, -59.2997, -58.71915, -58.1278, -57.52666, 
    -56.91667, -56.29873, -55.67367, -55.04227, -54.40527, -53.76335, 
    -53.11716, -52.46729, -51.8143, -51.1587, -50.50098, -49.84158, 
    -49.18093, -48.51939, -47.85734, -47.1951, -46.53297, -45.87124, 
    -45.21016, -44.54997, -43.89089, -43.23311, -42.57683,
  -42.77788, -43.44402, -44.11203, -44.78174, -45.45296, -46.12547, 
    -46.79906, -47.47348, -48.14844, -48.82367, -49.49884, -50.1736, 
    -50.84757, -51.52035, -52.1915, -52.86054, -53.52696, -54.1902, 
    -54.84966, -55.50471, -56.15464, -56.79872, -57.43615, -58.06607, 
    -58.68758, -59.2997, -59.90138, -60.49152, -61.06895, -61.63241, 
    -62.18061, -62.71215, -63.2256, -63.71946, -64.19215, -64.6421, 
    -65.06765, -65.46716, -65.83895, -66.18141, -66.49293, -66.77197, 
    -67.01707, -67.22693, -67.40035, -67.53634, -67.63406, -67.69295, 
    -67.71262, -67.69295, -67.63406, -67.53634, -67.40035, -67.22693, 
    -67.01707, -66.77197, -66.49293, -66.18141, -65.83895, -65.46716, 
    -65.06765, -64.6421, -64.19215, -63.71946, -63.2256, -62.71215, 
    -62.18061, -61.63241, -61.06895, -60.49152, -59.90138, -59.2997, 
    -58.68758, -58.06607, -57.43615, -56.79872, -56.15464, -55.50471, 
    -54.84966, -54.1902, -53.52696, -52.86054, -52.1915, -51.52035, 
    -50.84757, -50.1736, -49.49884, -48.82367, -48.14844, -47.47348, 
    -46.79906, -46.12547, -45.45296, -44.78174, -44.11203, -43.44402, 
    -42.77788,
  -42.97084, -43.64655, -44.3245, -45.00454, -45.68649, -46.37015, -47.05531, 
    -47.74172, -48.42913, -49.11726, -49.8058, -50.49441, -51.18272, 
    -51.87035, -52.55685, -53.24175, -53.92455, -54.60471, -55.28162, 
    -55.95465, -56.62309, -57.28621, -57.9432, -58.59319, -59.23526, 
    -59.86839, -60.49152, -61.1035, -61.70312, -62.28906, -62.85994, 
    -63.41431, -63.95062, -64.46726, -64.96255, -65.43473, -65.88202, 
    -66.30258, -66.69459, -67.05619, -67.38558, -67.68102, -67.94086, 
    -68.16358, -68.3478, -68.49236, -68.59633, -68.65899, -68.67992, 
    -68.65899, -68.59633, -68.49236, -68.3478, -68.16358, -67.94086, 
    -67.68102, -67.38558, -67.05619, -66.69459, -66.30258, -65.88202, 
    -65.43473, -64.96255, -64.46726, -63.95062, -63.41431, -62.85994, 
    -62.28906, -61.70312, -61.1035, -60.49152, -59.86839, -59.23526, 
    -58.59319, -57.9432, -57.28621, -56.62309, -55.95465, -55.28162, 
    -54.60471, -53.92455, -53.24175, -52.55685, -51.87035, -51.18272, 
    -50.49441, -49.8058, -49.11726, -48.42913, -47.74172, -47.05531, 
    -46.37015, -45.68649, -45.00454, -44.3245, -43.64655, -42.97084,
  -43.1556, -43.84056, -44.52815, -45.21821, -45.91058, -46.60506, -47.30147, 
    -47.99957, -48.69912, -49.39985, -50.10146, -50.80363, -51.506, -52.2082, 
    -52.9098, -53.61034, -54.30932, -55.00621, -55.70042, -56.39131, 
    -57.07819, -57.76032, -58.43688, -59.10701, -59.76975, -60.4241, 
    -61.06895, -61.70312, -62.32535, -62.93428, -63.52847, -64.10636, 
    -64.66634, -65.20666, -65.72551, -66.22101, -66.69118, -67.13403, 
    -67.54749, -67.9295, -68.27805, -68.59113, -68.86686, -69.10349, 
    -69.29943, -69.45333, -69.56409, -69.63087, -69.65318, -69.63087, 
    -69.56409, -69.45333, -69.29943, -69.10349, -68.86686, -68.59113, 
    -68.27805, -67.9295, -67.54749, -67.13403, -66.69118, -66.22101, 
    -65.72551, -65.20666, -64.66634, -64.10636, -63.52847, -62.93428, 
    -62.32535, -61.70312, -61.06895, -60.4241, -59.76975, -59.10701, 
    -58.43688, -57.76032, -57.07819, -56.39131, -55.70042, -55.00621, 
    -54.30932, -53.61034, -52.9098, -52.2082, -51.506, -50.80363, -50.10146, 
    -49.39985, -48.69912, -47.99957, -47.30147, -46.60506, -45.91058, 
    -45.21821, -44.52815, -43.84056, -43.1556,
  -43.33206, -44.02596, -44.72285, -45.42259, -46.12503, -46.83001, 
    -47.53732, -48.24677, -48.95811, -49.6711, -50.38545, -51.10085, 
    -51.81697, -52.53343, -53.24984, -53.96573, -54.68064, -55.39402, 
    -56.10532, -56.8139, -57.51908, -58.22011, -58.9162, -59.60646, 
    -60.28995, -60.96564, -61.63241, -62.28906, -62.93428, -63.56667, 
    -64.18473, -64.78683, -65.37125, -65.93615, -66.47958, -66.9995, 
    -67.49377, -67.96017, -68.39644, -68.80025, -69.16933, -69.50142, 
    -69.79435, -70.04609, -70.2548, -70.4189, -70.53708, -70.60838, 
    -70.63222, -70.60838, -70.53708, -70.4189, -70.2548, -70.04609, 
    -69.79435, -69.50142, -69.16933, -68.80025, -68.39644, -67.96017, 
    -67.49377, -66.9995, -66.47958, -65.93615, -65.37125, -64.78683, 
    -64.18473, -63.56667, -62.93428, -62.28906, -61.63241, -60.96564, 
    -60.28995, -59.60646, -58.9162, -58.22011, -57.51908, -56.8139, 
    -56.10532, -55.39402, -54.68064, -53.96573, -53.24984, -52.53343, 
    -51.81697, -51.10085, -50.38545, -49.6711, -48.95811, -48.24677, 
    -47.53732, -46.83001, -46.12503, -45.42259, -44.72285, -44.02596, 
    -43.33206,
  -43.50012, -44.20261, -44.90845, -45.61752, -46.32969, -47.04478, 
    -47.76263, -48.48305, -49.20582, -49.9307, -50.65742, -51.38569, 
    -52.11519, -52.84557, -53.57643, -54.30735, -55.03786, -55.76746, 
    -56.49557, -57.2216, -57.94487, -58.66464, -59.38013, -60.09047, 
    -60.79469, -61.49178, -62.18061, -62.85994, -63.52847, -64.18473, 
    -64.82718, -65.45412, -66.06374, -66.65411, -67.22313, -67.76861, 
    -68.28822, -68.77954, -69.24005, -69.66718, -70.05833, -70.41093, 
    -70.72251, -70.99072, -71.21339, -71.38868, -71.51503, -71.59132, 
    -71.61682, -71.59132, -71.51503, -71.38868, -71.21339, -70.99072, 
    -70.72251, -70.41093, -70.05833, -69.66718, -69.24005, -68.77954, 
    -68.28822, -67.76861, -67.22313, -66.65411, -66.06374, -65.45412, 
    -64.82718, -64.18473, -63.52847, -62.85994, -62.18061, -61.49178, 
    -60.79469, -60.09047, -59.38013, -58.66464, -57.94487, -57.2216, 
    -56.49557, -55.76746, -55.03786, -54.30735, -53.57643, -52.84557, 
    -52.11519, -51.38569, -50.65742, -49.9307, -49.20582, -48.48305, 
    -47.76263, -47.04478, -46.32969, -45.61752, -44.90845, -44.20261, 
    -43.50012,
  -43.65969, -44.37041, -45.08484, -45.80286, -46.52436, -47.24918, 
    -47.97718, -48.70818, -49.44197, -50.17833, -50.91702, -51.65775, 
    -52.40023, -53.14412, -53.88906, -54.63462, -55.38037, -56.12582, 
    -56.87043, -57.61359, -58.35467, -59.09295, -59.82764, -60.55789, 
    -61.28276, -62.00122, -62.71215, -63.41431, -64.10636, -64.78683, 
    -65.45412, -66.10648, -66.74202, -67.3587, -67.95432, -68.5265, 
    -69.07276, -69.59042, -70.07672, -70.52879, -70.9437, -71.31852, 
    -71.6504, -71.9366, -72.17461, -72.36224, -72.49763, -72.57942, 
    -72.60679, -72.57942, -72.49763, -72.36224, -72.17461, -71.9366, 
    -71.6504, -71.31852, -70.9437, -70.52879, -70.07672, -69.59042, 
    -69.07276, -68.5265, -67.95432, -67.3587, -66.74202, -66.10648, 
    -65.45412, -64.78683, -64.10636, -63.41431, -62.71215, -62.00122, 
    -61.28276, -60.55789, -59.82764, -59.09295, -58.35467, -57.61359, 
    -56.87043, -56.12582, -55.38037, -54.63462, -53.88906, -53.14412, 
    -52.40023, -51.65775, -50.91702, -50.17833, -49.44197, -48.70818, 
    -47.97718, -47.24918, -46.52436, -45.80286, -45.08484, -44.37041, 
    -43.65969,
  -43.81068, -44.52925, -45.25187, -45.97845, -46.70888, -47.44304, 
    -48.18076, -48.92191, -49.66629, -50.4137, -51.1639, -51.91666, 
    -52.67167, -53.42863, -54.18719, -54.94697, -55.70753, -56.46842, 
    -57.22911, -57.98904, -58.74758, -59.50403, -60.25764, -61.00757, 
    -61.7529, -62.49262, -63.2256, -63.95062, -64.66634, -65.37125, 
    -66.06374, -66.74202, -67.40413, -68.04794, -68.67112, -69.27117, 
    -69.84539, -70.39089, -70.90462, -71.38338, -71.8239, -72.22283, 
    -72.57687, -72.88284, -73.13778, -73.33907, -73.4845, -73.57245, 
    -73.60188, -73.57245, -73.4845, -73.33907, -73.13778, -72.88284, 
    -72.57687, -72.22283, -71.8239, -71.38338, -70.90462, -70.39089, 
    -69.84539, -69.27117, -68.67112, -68.04794, -67.40413, -66.74202, 
    -66.06374, -65.37125, -64.66634, -63.95062, -63.2256, -62.49262, 
    -61.7529, -61.00757, -60.25764, -59.50403, -58.74758, -57.98904, 
    -57.22911, -56.46842, -55.70753, -54.94697, -54.18719, -53.42863, 
    -52.67167, -51.91666, -51.1639, -50.4137, -49.66629, -48.92191, 
    -48.18076, -47.44304, -46.70888, -45.97845, -45.25187, -44.52925, 
    -43.81068,
  -43.95298, -44.67902, -45.40944, -46.14417, -46.8831, -47.62614, -48.37315, 
    -49.124, -49.8785, -50.63649, -51.39774, -52.16203, -52.92909, -53.69863, 
    -54.47033, -55.24382, -56.01871, -56.79456, -57.57087, -58.34711, 
    -59.12267, -59.89689, -60.66905, -61.43833, -62.20383, -62.96457, 
    -63.71946, -64.46726, -65.20666, -65.93615, -66.65411, -67.3587, 
    -68.04794, -68.7196, -69.37128, -70.00032, -70.60384, -71.17871, 
    -71.7216, -72.22897, -72.69713, -73.12227, -73.50058, -73.82835, 
    -74.10206, -74.31858, -74.47527, -74.57011, -74.60188, -74.57011, 
    -74.47527, -74.31858, -74.10206, -73.82835, -73.50058, -73.12227, 
    -72.69713, -72.22897, -71.7216, -71.17871, -70.60384, -70.00032, 
    -69.37128, -68.7196, -68.04794, -67.3587, -66.65411, -65.93615, 
    -65.20666, -64.46726, -63.71946, -62.96457, -62.20383, -61.43833, 
    -60.66905, -59.89689, -59.12267, -58.34711, -57.57087, -56.79456, 
    -56.01871, -55.24382, -54.47033, -53.69863, -52.92909, -52.16203, 
    -51.39774, -50.63649, -49.8785, -49.124, -48.37315, -47.62614, -46.8831, 
    -46.14417, -45.40944, -44.67902, -43.95298,
  -44.08652, -44.81961, -45.55742, -46.29986, -47.04686, -47.79833, 
    -48.55416, -49.31422, -50.07836, -50.84642, -51.6182, -52.39351, 
    -53.17208, -53.95366, -54.73795, -55.52462, -56.31329, -57.10355, 
    -57.89494, -58.68696, -59.47903, -60.27053, -61.06076, -61.84895, 
    -62.63423, -63.41565, -64.19215, -64.96255, -65.72551, -66.47958, 
    -67.22313, -67.95432, -68.67112, -69.37128, -70.0523, -70.7114, 
    -71.34553, -71.95134, -72.5252, -73.06321, -73.56123, -74.01492, 
    -74.41991, -74.77181, -75.06647, -75.30009, -75.46947, -75.57212, 
    -75.60651, -75.57212, -75.46947, -75.30009, -75.06647, -74.77181, 
    -74.41991, -74.01492, -73.56123, -73.06321, -72.5252, -71.95134, 
    -71.34553, -70.7114, -70.0523, -69.37128, -68.67112, -67.95432, 
    -67.22313, -66.47958, -65.72551, -64.96255, -64.19215, -63.41565, 
    -62.63423, -61.84895, -61.06076, -60.27053, -59.47903, -58.68696, 
    -57.89494, -57.10355, -56.31329, -55.52462, -54.73795, -53.95366, 
    -53.17208, -52.39351, -51.6182, -50.84642, -50.07836, -49.31422, 
    -48.55416, -47.79833, -47.04686, -46.29986, -45.55742, -44.81961, 
    -44.08652,
  -44.21122, -44.95095, -45.6957, -46.4454, -47.20001, -47.95944, -48.72359, 
    -49.49236, -50.26561, -51.04321, -51.82498, -52.61073, -53.40025, 
    -54.19329, -54.98958, -55.78882, -56.59066, -57.39472, -58.20058, 
    -59.00777, -59.81574, -60.62392, -61.43166, -62.2382, -63.04275, 
    -63.84439, -64.6421, -65.43473, -66.22101, -66.9995, -67.76861, -68.5265, 
    -69.27117, -70.00032, -70.7114, -71.40154, -72.06753, -72.70583, 
    -73.31252, -73.88333, -74.41362, -74.8985, -75.33289, -75.71165, 
    -76.02982, -76.28278, -76.46657, -76.57815, -76.61555, -76.57815, 
    -76.46657, -76.28278, -76.02982, -75.71165, -75.33289, -74.8985, 
    -74.41362, -73.88333, -73.31252, -72.70583, -72.06753, -71.40154, 
    -70.7114, -70.00032, -69.27117, -68.5265, -67.76861, -66.9995, -66.22101, 
    -65.43473, -64.6421, -63.84439, -63.04275, -62.2382, -61.43166, 
    -60.62392, -59.81574, -59.00777, -58.20058, -57.39472, -56.59066, 
    -55.78882, -54.98958, -54.19329, -53.40025, -52.61073, -51.82498, 
    -51.04321, -50.26561, -49.49236, -48.72359, -47.95944, -47.20001, 
    -46.4454, -45.6957, -44.95095, -44.21122,
  -44.32701, -45.07294, -45.82418, -46.58068, -47.34241, -48.10929, 
    -48.88126, -49.6582, -50.44002, -51.22659, -52.01776, -52.81337, 
    -53.61321, -54.41708, -55.22473, -56.03588, -56.85022, -57.66741, 
    -58.48705, -59.30871, -60.1319, -60.95608, -61.78063, -62.60488, 
    -63.42805, -64.2493, -65.06765, -65.88202, -66.69118, -67.49377, 
    -68.28822, -69.07276, -69.84539, -70.60384, -71.34553, -72.06753, 
    -72.76654, -73.43884, -74.08022, -74.68606, -75.25123, -75.77019, 
    -76.23708, -76.64588, -76.99059, -77.26559, -77.46595, -77.58782, 
    -77.62873, -77.58782, -77.46595, -77.26559, -76.99059, -76.64588, 
    -76.23708, -75.77019, -75.25123, -74.68606, -74.08022, -73.43884, 
    -72.76654, -72.06753, -71.34553, -70.60384, -69.84539, -69.07276, 
    -68.28822, -67.49377, -66.69118, -65.88202, -65.06765, -64.2493, 
    -63.42805, -62.60488, -61.78063, -60.95608, -60.1319, -59.30871, 
    -58.48705, -57.66741, -56.85022, -56.03588, -55.22473, -54.41708, 
    -53.61321, -52.81337, -52.01776, -51.22659, -50.44002, -49.6582, 
    -48.88126, -48.10929, -47.34241, -46.58068, -45.82418, -45.07294, 
    -44.32701,
  -44.4338, -45.18549, -45.94276, -46.70559, -47.47393, -48.24775, -49.02699, 
    -49.81155, -50.60136, -51.39631, -52.19627, -53.00109, -53.81061, 
    -54.62463, -55.44294, -56.26529, -57.09141, -57.92097, -58.75364, 
    -59.589, -60.42662, -61.26601, -62.10659, -62.94775, -63.78878, 
    -64.62888, -65.46716, -66.30258, -67.13403, -67.96017, -68.77954, 
    -69.59042, -70.39089, -71.17871, -71.95134, -72.70583, -73.43884, 
    -74.14648, -74.82438, -75.46753, -76.07032, -76.62655, -77.12947, 
    -77.572, -77.94691, -78.24726, -78.46685, -78.60075, -78.64574, 
    -78.60075, -78.46685, -78.24726, -77.94691, -77.572, -77.12947, 
    -76.62655, -76.07032, -75.46753, -74.82438, -74.14648, -73.43884, 
    -72.70583, -71.95134, -71.17871, -70.39089, -69.59042, -68.77954, 
    -67.96017, -67.13403, -66.30258, -65.46716, -64.62888, -63.78878, 
    -62.94775, -62.10659, -61.26601, -60.42662, -59.589, -58.75364, 
    -57.92097, -57.09141, -56.26529, -55.44294, -54.62463, -53.81061, 
    -53.00109, -52.19627, -51.39631, -50.60136, -49.81155, -49.02699, 
    -48.24775, -47.47393, -46.70559, -45.94276, -45.18549, -44.4338,
  -44.53154, -45.28852, -46.05135, -46.82, -47.59445, -48.37467, -49.16062, 
    -49.95222, -50.74942, -51.55212, -52.36022, -53.17359, -53.99209, 
    -54.81555, -55.64378, -56.47657, -57.31367, -58.1548, -58.99965, 
    -59.84786, -60.69904, -61.55275, -62.40846, -63.26563, -64.1236, 
    -64.98164, -65.83895, -66.69459, -67.54749, -68.39644, -69.24005, 
    -70.07672, -70.90462, -71.7216, -72.5252, -73.31252, -74.08022, 
    -74.82438, -75.54044, -76.22314, -76.86639, -77.46332, -78.00623, 
    -78.4868, -78.89631, -79.22611, -79.46831, -79.61646, -79.66634, 
    -79.61646, -79.46831, -79.22611, -78.89631, -78.4868, -78.00623, 
    -77.46332, -76.86639, -76.22314, -75.54044, -74.82438, -74.08022, 
    -73.31252, -72.5252, -71.7216, -70.90462, -70.07672, -69.24005, 
    -68.39644, -67.54749, -66.69459, -65.83895, -64.98164, -64.1236, 
    -63.26563, -62.40846, -61.55275, -60.69904, -59.84786, -58.99965, 
    -58.1548, -57.31367, -56.47657, -55.64378, -54.81555, -53.99209, 
    -53.17359, -52.36022, -51.55212, -50.74942, -49.95222, -49.16062, 
    -48.37467, -47.59445, -46.82, -46.05135, -45.28852, -44.53154,
  -44.62016, -45.38197, -46.14986, -46.92382, -47.70385, -48.48992, -49.282, 
    -50.08005, -50.88401, -51.69381, -52.50938, -53.33059, -54.15733, 
    -54.98947, -55.82684, -56.66924, -57.51648, -58.36829, -59.22443, 
    -60.08456, -60.94834, -61.81537, -62.6852, -63.55734, -64.4312, 
    -65.30614, -66.18141, -67.05619, -67.9295, -68.80025, -69.66718, 
    -70.52879, -71.38338, -72.22897, -73.06321, -73.88333, -74.68606, 
    -75.46753, -76.22314, -76.94742, -77.63395, -78.2752, -78.8625, 
    -79.38612, -79.83553, -80.19992, -80.46906, -80.6344, -80.69019, 
    -80.6344, -80.46906, -80.19992, -79.83553, -79.38612, -78.8625, -78.2752, 
    -77.63395, -76.94742, -76.22314, -75.46753, -74.68606, -73.88333, 
    -73.06321, -72.22897, -71.38338, -70.52879, -69.66718, -68.80025, 
    -67.9295, -67.05619, -66.18141, -65.30614, -64.4312, -63.55734, -62.6852, 
    -61.81537, -60.94834, -60.08456, -59.22443, -58.36829, -57.51648, 
    -56.66924, -55.82684, -54.98947, -54.15733, -53.33059, -52.50938, 
    -51.69381, -50.88401, -50.08005, -49.282, -48.48992, -47.70385, 
    -46.92382, -46.14986, -45.38197, -44.62016,
  -44.6996, -45.46576, -46.23822, -47.01697, -47.80202, -48.59336, -49.39099, 
    -50.19486, -51.00494, -51.82117, -52.64349, -53.47181, -54.30604, 
    -55.14605, -55.99172, -56.84288, -57.69935, -58.56092, -59.42736, 
    -60.29839, -61.17372, -62.05299, -62.93583, -63.82177, -64.71033, 
    -65.60093, -66.49293, -67.38558, -68.27805, -69.16933, -70.05833, 
    -70.9437, -71.8239, -72.69713, -73.56123, -74.41362, -75.25123, 
    -76.07032, -76.86639, -77.63395, -78.36636, -79.05556, -79.69198, 
    -80.2644, -80.76014, -81.16562, -81.46742, -81.65389, -81.71702, 
    -81.65389, -81.46742, -81.16562, -80.76014, -80.2644, -79.69198, 
    -79.05556, -78.36636, -77.63395, -76.86639, -76.07032, -75.25123, 
    -74.41362, -73.56123, -72.69713, -71.8239, -70.9437, -70.05833, 
    -69.16933, -68.27805, -67.38558, -66.49293, -65.60093, -64.71033, 
    -63.82177, -62.93583, -62.05299, -61.17372, -60.29839, -59.42736, 
    -58.56092, -57.69935, -56.84288, -55.99172, -55.14605, -54.30604, 
    -53.47181, -52.64349, -51.82117, -51.00494, -50.19486, -49.39099, 
    -48.59336, -47.80202, -47.01697, -46.23822, -45.46576, -44.6996,
  -44.76982, -45.53984, -46.31635, -47.09935, -47.88887, -48.68491, 
    -49.48746, -50.29652, -51.11204, -51.934, -52.76235, -53.59702, 
    -54.43793, -55.28499, -56.13808, -56.99708, -57.86184, -58.73216, 
    -59.60787, -60.48872, -61.37446, -62.26479, -63.15939, -64.05786, 
    -64.95979, -65.86467, -66.77197, -67.68102, -68.59113, -69.50142, 
    -70.41093, -71.31852, -72.22283, -73.12227, -74.01492, -74.8985, 
    -75.77019, -76.62655, -77.46332, -78.2752, -79.05556, -79.7961, 
    -80.48651, -81.11414, -81.66392, -82.11877, -82.46091, -82.67403, 
    -82.7465, -82.67403, -82.46091, -82.11877, -81.66392, -81.11414, 
    -80.48651, -79.7961, -79.05556, -78.2752, -77.46332, -76.62655, 
    -75.77019, -74.8985, -74.01492, -73.12227, -72.22283, -71.31852, 
    -70.41093, -69.50142, -68.59113, -67.68102, -66.77197, -65.86467, 
    -64.95979, -64.05786, -63.15939, -62.26479, -61.37446, -60.48872, 
    -59.60787, -58.73216, -57.86184, -56.99708, -56.13808, -55.28499, 
    -54.43793, -53.59702, -52.76235, -51.934, -51.11204, -50.29652, 
    -49.48746, -48.68491, -47.88887, -47.09935, -46.31635, -45.53984, 
    -44.76982,
  -44.83077, -45.60415, -46.38419, -47.17091, -47.96432, -48.76445, 
    -49.57131, -50.38489, -51.20517, -52.03214, -52.86576, -53.70599, 
    -54.55275, -55.40599, -56.26561, -57.13149, -58.00352, -58.88156, 
    -59.76543, -60.65495, -61.54989, -62.45001, -63.35503, -64.26463, 
    -65.17846, -66.09609, -67.01707, -67.94086, -68.86686, -69.79435, 
    -70.72251, -71.6504, -72.57687, -73.50058, -74.41991, -75.33289, 
    -76.23708, -77.12947, -78.00623, -78.8625, -79.69198, -80.48651, 
    -81.23547, -81.92511, -82.53796, -83.0528, -83.44577, -83.69351, 
    -83.77832, -83.69351, -83.44577, -83.0528, -82.53796, -81.92511, 
    -81.23547, -80.48651, -79.69198, -78.8625, -78.00623, -77.12947, 
    -76.23708, -75.33289, -74.41991, -73.50058, -72.57687, -71.6504, 
    -70.72251, -69.79435, -68.86686, -67.94086, -67.01707, -66.09609, 
    -65.17846, -64.26463, -63.35503, -62.45001, -61.54989, -60.65495, 
    -59.76543, -58.88156, -58.00352, -57.13149, -56.26561, -55.40599, 
    -54.55275, -53.70599, -52.86576, -52.03214, -51.20517, -50.38489, 
    -49.57131, -48.76445, -47.96432, -47.17091, -46.38419, -45.60415, 
    -44.83077,
  -44.88241, -45.65865, -46.44169, -47.23156, -48.02829, -48.83191, 
    -49.64243, -50.45986, -51.2842, -52.11544, -52.95356, -53.79853, 
    -54.6503, -55.50881, -56.374, -57.24578, -58.12405, -59.0087, -59.89958, 
    -60.79654, -61.6994, -62.60796, -63.52198, -64.4412, -65.36533, 
    -66.29404, -67.22693, -68.16358, -69.10349, -70.04609, -70.99072, 
    -71.9366, -72.88284, -73.82835, -74.77181, -75.71165, -76.64588, -77.572, 
    -78.4868, -79.38612, -80.2644, -81.11414, -81.92511, -82.6832, -83.36916, 
    -83.95731, -84.41584, -84.71027, -84.81216, -84.71027, -84.41584, 
    -83.95731, -83.36916, -82.6832, -81.92511, -81.11414, -80.2644, 
    -79.38612, -78.4868, -77.572, -76.64588, -75.71165, -74.77181, -73.82835, 
    -72.88284, -71.9366, -70.99072, -70.04609, -69.10349, -68.16358, 
    -67.22693, -66.29404, -65.36533, -64.4412, -63.52198, -62.60796, 
    -61.6994, -60.79654, -59.89958, -59.0087, -58.12405, -57.24578, -56.374, 
    -55.50881, -54.6503, -53.79853, -52.95356, -52.11544, -51.2842, 
    -50.45986, -49.64243, -48.83191, -48.02829, -47.23156, -46.44169, 
    -45.65865, -44.88241,
  -44.9247, -45.7033, -46.4888, -47.28126, -48.08072, -48.8872, -49.70073, 
    -50.52134, -51.34902, -52.18378, -53.0256, -53.87448, -54.73037, 
    -55.59324, -56.46303, -57.33968, -58.22311, -59.11322, -60.00991, 
    -60.91304, -61.82248, -62.73804, -63.65955, -64.58678, -65.51952, 
    -66.45748, -67.40035, -68.3478, -69.29943, -70.2548, -71.21339, 
    -72.17461, -73.13778, -74.10206, -75.06647, -76.02982, -76.99059, 
    -77.94691, -78.89631, -79.83553, -80.76014, -81.66392, -82.53796, 
    -83.36916, -84.13799, -84.81542, -85.36021, -85.72057, -85.84769, 
    -85.72057, -85.36021, -84.81542, -84.13799, -83.36916, -82.53796, 
    -81.66392, -80.76014, -79.83553, -78.89631, -77.94691, -76.99059, 
    -76.02982, -75.06647, -74.10206, -73.13778, -72.17461, -71.21339, 
    -70.2548, -69.29943, -68.3478, -67.40035, -66.45748, -65.51952, 
    -64.58678, -63.65955, -62.73804, -61.82248, -60.91304, -60.00991, 
    -59.11322, -58.22311, -57.33968, -56.46303, -55.59324, -54.73037, 
    -53.87448, -53.0256, -52.18378, -51.34902, -50.52134, -49.70073, 
    -48.8872, -48.08072, -47.28126, -46.4888, -45.7033, -44.9247,
  -44.95763, -45.73805, -46.52548, -47.31997, -48.12155, -48.93027, 
    -49.74615, -50.56924, -51.39953, -52.23703, -53.08176, -53.93369, 
    -54.79281, -55.65909, -56.53249, -57.41296, -58.30043, -59.19484, 
    -60.09608, -61.00407, -61.91867, -62.83975, -63.76716, -64.70073, 
    -65.64027, -66.58555, -67.53634, -68.49236, -69.45333, -70.4189, 
    -71.38868, -72.36224, -73.33907, -74.31858, -75.30009, -76.28278, 
    -77.26559, -78.24726, -79.22611, -80.19992, -81.16562, -82.11877, 
    -83.0528, -83.95731, -84.81542, -85.59846, -86.25768, -86.71655, 
    -86.88457, -86.71655, -86.25768, -85.59846, -84.81542, -83.95731, 
    -83.0528, -82.11877, -81.16562, -80.19992, -79.22611, -78.24726, 
    -77.26559, -76.28278, -75.30009, -74.31858, -73.33907, -72.36224, 
    -71.38868, -70.4189, -69.45333, -68.49236, -67.53634, -66.58555, 
    -65.64027, -64.70073, -63.76716, -62.83975, -61.91867, -61.00407, 
    -60.09608, -59.19484, -58.30043, -57.41296, -56.53249, -55.65909, 
    -54.79281, -53.93369, -53.08176, -52.23703, -51.39953, -50.56924, 
    -49.74615, -48.93027, -48.12155, -47.31997, -46.52548, -45.73805, 
    -44.95763,
  -44.98116, -45.7629, -46.5517, -47.34763, -48.15074, -48.96106, -49.77864, 
    -50.6035, -51.43566, -52.27514, -53.12194, -53.97606, -54.8375, 
    -55.70623, -56.58222, -57.46543, -58.35581, -59.2533, -60.15783, 
    -61.06931, -61.98763, -62.91269, -63.84436, -64.7825, -65.72695, 
    -66.67754, -67.63406, -68.59633, -69.56409, -70.53708, -71.51503, 
    -72.49763, -73.4845, -74.47527, -75.46947, -76.46657, -77.46595, 
    -78.46685, -79.46831, -80.46906, -81.46742, -82.46091, -83.44577, 
    -84.41584, -85.36021, -86.25768, -87.06323, -87.6776, -87.92248, 
    -87.6776, -87.06323, -86.25768, -85.36021, -84.41584, -83.44577, 
    -82.46091, -81.46742, -80.46906, -79.46831, -78.46685, -77.46595, 
    -76.46657, -75.46947, -74.47527, -73.4845, -72.49763, -71.51503, 
    -70.53708, -69.56409, -68.59633, -67.63406, -66.67754, -65.72695, 
    -64.7825, -63.84436, -62.91269, -61.98763, -61.06931, -60.15783, 
    -59.2533, -58.35581, -57.46543, -56.58222, -55.70623, -54.8375, 
    -53.97606, -53.12194, -52.27514, -51.43566, -50.6035, -49.77864, 
    -48.96106, -48.15074, -47.34763, -46.5517, -45.7629, -44.98116,
  -44.99529, -45.77781, -46.56744, -47.36425, -48.16827, -48.97956, 
    -49.79815, -50.62407, -51.45736, -52.29802, -53.14607, -54.00152, 
    -54.86435, -55.73455, -56.6121, -57.49697, -58.3891, -59.28845, 
    -60.19496, -61.10854, -62.02911, -62.95657, -63.89082, -64.83172, 
    -65.77914, -66.73294, -67.69295, -68.65899, -69.63087, -70.60838, 
    -71.59132, -72.57942, -73.57245, -74.57011, -75.57212, -76.57815, 
    -77.58782, -78.60075, -79.61646, -80.6344, -81.65389, -82.67403, 
    -83.69351, -84.71027, -85.72057, -86.71655, -87.6776, -88.53089, 
    -88.96107, -88.53089, -87.6776, -86.71655, -85.72057, -84.71027, 
    -83.69351, -82.67403, -81.65389, -80.6344, -79.61646, -78.60075, 
    -77.58782, -76.57815, -75.57212, -74.57011, -73.57245, -72.57942, 
    -71.59132, -70.60838, -69.63087, -68.65899, -67.69295, -66.73294, 
    -65.77914, -64.83172, -63.89082, -62.95657, -62.02911, -61.10854, 
    -60.19496, -59.28845, -58.3891, -57.49697, -56.6121, -55.73455, 
    -54.86435, -54.00152, -53.14607, -52.29802, -51.45736, -50.62407, 
    -49.79815, -48.97956, -48.16827, -47.36425, -46.56744, -45.77781, 
    -44.99529,
  -45, -45.78278, -46.57269, -47.36979, -48.17411, -48.98572, -49.80465, 
    -50.63093, -51.46459, -52.30565, -53.15412, -54.01001, -54.87331, 
    -55.744, -56.62207, -57.50749, -58.40021, -59.30018, -60.20734, 
    -61.12163, -62.04295, -62.97122, -63.90633, -64.84815, -65.79657, 
    -66.75144, -67.71262, -68.67992, -69.65318, -70.63222, -71.61682, 
    -72.60679, -73.60188, -74.60188, -75.60651, -76.61555, -77.62873, 
    -78.64574, -79.66634, -80.69019, -81.71702, -82.7465, -83.77832, 
    -84.81216, -85.84769, -86.88457, -87.92248, -88.96107, -90, -88.96107, 
    -87.92248, -86.88457, -85.84769, -84.81216, -83.77832, -82.7465, 
    -81.71702, -80.69019, -79.66634, -78.64574, -77.62873, -76.61555, 
    -75.60651, -74.60188, -73.60188, -72.60679, -71.61682, -70.63222, 
    -69.65318, -68.67992, -67.71262, -66.75144, -65.79657, -64.84815, 
    -63.90633, -62.97122, -62.04295, -61.12163, -60.20734, -59.30018, 
    -58.40021, -57.50749, -56.62207, -55.744, -54.87331, -54.01001, 
    -53.15412, -52.30565, -51.46459, -50.63093, -49.80465, -48.98572, 
    -48.17411, -47.36979, -46.57269, -45.78278, -45,
  -44.99529, -45.77781, -46.56744, -47.36425, -48.16827, -48.97956, 
    -49.79815, -50.62407, -51.45736, -52.29802, -53.14607, -54.00152, 
    -54.86435, -55.73455, -56.6121, -57.49697, -58.3891, -59.28845, 
    -60.19496, -61.10854, -62.02911, -62.95657, -63.89082, -64.83172, 
    -65.77914, -66.73294, -67.69295, -68.65899, -69.63087, -70.60838, 
    -71.59132, -72.57942, -73.57245, -74.57011, -75.57212, -76.57815, 
    -77.58782, -78.60075, -79.61646, -80.6344, -81.65389, -82.67403, 
    -83.69351, -84.71027, -85.72057, -86.71655, -87.6776, -88.53089, 
    -88.96107, -88.53089, -87.6776, -86.71655, -85.72057, -84.71027, 
    -83.69351, -82.67403, -81.65389, -80.6344, -79.61646, -78.60075, 
    -77.58782, -76.57815, -75.57212, -74.57011, -73.57245, -72.57942, 
    -71.59132, -70.60838, -69.63087, -68.65899, -67.69295, -66.73294, 
    -65.77914, -64.83172, -63.89082, -62.95657, -62.02911, -61.10854, 
    -60.19496, -59.28845, -58.3891, -57.49697, -56.6121, -55.73455, 
    -54.86435, -54.00152, -53.14607, -52.29802, -51.45736, -50.62407, 
    -49.79815, -48.97956, -48.16827, -47.36425, -46.56744, -45.77781, 
    -44.99529,
  -44.98116, -45.7629, -46.5517, -47.34763, -48.15074, -48.96106, -49.77864, 
    -50.6035, -51.43566, -52.27514, -53.12194, -53.97606, -54.8375, 
    -55.70623, -56.58222, -57.46543, -58.35581, -59.2533, -60.15783, 
    -61.06931, -61.98763, -62.91269, -63.84436, -64.7825, -65.72695, 
    -66.67754, -67.63406, -68.59633, -69.56409, -70.53708, -71.51503, 
    -72.49763, -73.4845, -74.47527, -75.46947, -76.46657, -77.46595, 
    -78.46685, -79.46831, -80.46906, -81.46742, -82.46091, -83.44577, 
    -84.41584, -85.36021, -86.25768, -87.06323, -87.6776, -87.92248, 
    -87.6776, -87.06323, -86.25768, -85.36021, -84.41584, -83.44577, 
    -82.46091, -81.46742, -80.46906, -79.46831, -78.46685, -77.46595, 
    -76.46657, -75.46947, -74.47527, -73.4845, -72.49763, -71.51503, 
    -70.53708, -69.56409, -68.59633, -67.63406, -66.67754, -65.72695, 
    -64.7825, -63.84436, -62.91269, -61.98763, -61.06931, -60.15783, 
    -59.2533, -58.35581, -57.46543, -56.58222, -55.70623, -54.8375, 
    -53.97606, -53.12194, -52.27514, -51.43566, -50.6035, -49.77864, 
    -48.96106, -48.15074, -47.34763, -46.5517, -45.7629, -44.98116,
  -44.95763, -45.73805, -46.52548, -47.31997, -48.12155, -48.93027, 
    -49.74615, -50.56924, -51.39953, -52.23703, -53.08176, -53.93369, 
    -54.79281, -55.65909, -56.53249, -57.41296, -58.30043, -59.19484, 
    -60.09608, -61.00407, -61.91867, -62.83975, -63.76716, -64.70073, 
    -65.64027, -66.58555, -67.53634, -68.49236, -69.45333, -70.4189, 
    -71.38868, -72.36224, -73.33907, -74.31858, -75.30009, -76.28278, 
    -77.26559, -78.24726, -79.22611, -80.19992, -81.16562, -82.11877, 
    -83.0528, -83.95731, -84.81542, -85.59846, -86.25768, -86.71655, 
    -86.88457, -86.71655, -86.25768, -85.59846, -84.81542, -83.95731, 
    -83.0528, -82.11877, -81.16562, -80.19992, -79.22611, -78.24726, 
    -77.26559, -76.28278, -75.30009, -74.31858, -73.33907, -72.36224, 
    -71.38868, -70.4189, -69.45333, -68.49236, -67.53634, -66.58555, 
    -65.64027, -64.70073, -63.76716, -62.83975, -61.91867, -61.00407, 
    -60.09608, -59.19484, -58.30043, -57.41296, -56.53249, -55.65909, 
    -54.79281, -53.93369, -53.08176, -52.23703, -51.39953, -50.56924, 
    -49.74615, -48.93027, -48.12155, -47.31997, -46.52548, -45.73805, 
    -44.95763,
  -44.9247, -45.7033, -46.4888, -47.28126, -48.08072, -48.8872, -49.70073, 
    -50.52134, -51.34902, -52.18378, -53.0256, -53.87448, -54.73037, 
    -55.59324, -56.46303, -57.33968, -58.22311, -59.11322, -60.00991, 
    -60.91304, -61.82248, -62.73804, -63.65955, -64.58678, -65.51952, 
    -66.45748, -67.40035, -68.3478, -69.29943, -70.2548, -71.21339, 
    -72.17461, -73.13778, -74.10206, -75.06647, -76.02982, -76.99059, 
    -77.94691, -78.89631, -79.83553, -80.76014, -81.66392, -82.53796, 
    -83.36916, -84.13799, -84.81542, -85.36021, -85.72057, -85.84769, 
    -85.72057, -85.36021, -84.81542, -84.13799, -83.36916, -82.53796, 
    -81.66392, -80.76014, -79.83553, -78.89631, -77.94691, -76.99059, 
    -76.02982, -75.06647, -74.10206, -73.13778, -72.17461, -71.21339, 
    -70.2548, -69.29943, -68.3478, -67.40035, -66.45748, -65.51952, 
    -64.58678, -63.65955, -62.73804, -61.82248, -60.91304, -60.00991, 
    -59.11322, -58.22311, -57.33968, -56.46303, -55.59324, -54.73037, 
    -53.87448, -53.0256, -52.18378, -51.34902, -50.52134, -49.70073, 
    -48.8872, -48.08072, -47.28126, -46.4888, -45.7033, -44.9247,
  -44.88241, -45.65865, -46.44169, -47.23156, -48.02829, -48.83191, 
    -49.64243, -50.45986, -51.2842, -52.11544, -52.95356, -53.79853, 
    -54.6503, -55.50881, -56.374, -57.24578, -58.12405, -59.0087, -59.89958, 
    -60.79654, -61.6994, -62.60796, -63.52198, -64.4412, -65.36533, 
    -66.29404, -67.22693, -68.16358, -69.10349, -70.04609, -70.99072, 
    -71.9366, -72.88284, -73.82835, -74.77181, -75.71165, -76.64588, -77.572, 
    -78.4868, -79.38612, -80.2644, -81.11414, -81.92511, -82.6832, -83.36916, 
    -83.95731, -84.41584, -84.71027, -84.81216, -84.71027, -84.41584, 
    -83.95731, -83.36916, -82.6832, -81.92511, -81.11414, -80.2644, 
    -79.38612, -78.4868, -77.572, -76.64588, -75.71165, -74.77181, -73.82835, 
    -72.88284, -71.9366, -70.99072, -70.04609, -69.10349, -68.16358, 
    -67.22693, -66.29404, -65.36533, -64.4412, -63.52198, -62.60796, 
    -61.6994, -60.79654, -59.89958, -59.0087, -58.12405, -57.24578, -56.374, 
    -55.50881, -54.6503, -53.79853, -52.95356, -52.11544, -51.2842, 
    -50.45986, -49.64243, -48.83191, -48.02829, -47.23156, -46.44169, 
    -45.65865, -44.88241,
  -44.83077, -45.60415, -46.38419, -47.17091, -47.96432, -48.76445, 
    -49.57131, -50.38489, -51.20517, -52.03214, -52.86576, -53.70599, 
    -54.55275, -55.40599, -56.26561, -57.13149, -58.00352, -58.88156, 
    -59.76543, -60.65495, -61.54989, -62.45001, -63.35503, -64.26463, 
    -65.17846, -66.09609, -67.01707, -67.94086, -68.86686, -69.79435, 
    -70.72251, -71.6504, -72.57687, -73.50058, -74.41991, -75.33289, 
    -76.23708, -77.12947, -78.00623, -78.8625, -79.69198, -80.48651, 
    -81.23547, -81.92511, -82.53796, -83.0528, -83.44577, -83.69351, 
    -83.77832, -83.69351, -83.44577, -83.0528, -82.53796, -81.92511, 
    -81.23547, -80.48651, -79.69198, -78.8625, -78.00623, -77.12947, 
    -76.23708, -75.33289, -74.41991, -73.50058, -72.57687, -71.6504, 
    -70.72251, -69.79435, -68.86686, -67.94086, -67.01707, -66.09609, 
    -65.17846, -64.26463, -63.35503, -62.45001, -61.54989, -60.65495, 
    -59.76543, -58.88156, -58.00352, -57.13149, -56.26561, -55.40599, 
    -54.55275, -53.70599, -52.86576, -52.03214, -51.20517, -50.38489, 
    -49.57131, -48.76445, -47.96432, -47.17091, -46.38419, -45.60415, 
    -44.83077,
  -44.76982, -45.53984, -46.31635, -47.09935, -47.88887, -48.68491, 
    -49.48746, -50.29652, -51.11204, -51.934, -52.76235, -53.59702, 
    -54.43793, -55.28499, -56.13808, -56.99708, -57.86184, -58.73216, 
    -59.60787, -60.48872, -61.37446, -62.26479, -63.15939, -64.05786, 
    -64.95979, -65.86467, -66.77197, -67.68102, -68.59113, -69.50142, 
    -70.41093, -71.31852, -72.22283, -73.12227, -74.01492, -74.8985, 
    -75.77019, -76.62655, -77.46332, -78.2752, -79.05556, -79.7961, 
    -80.48651, -81.11414, -81.66392, -82.11877, -82.46091, -82.67403, 
    -82.7465, -82.67403, -82.46091, -82.11877, -81.66392, -81.11414, 
    -80.48651, -79.7961, -79.05556, -78.2752, -77.46332, -76.62655, 
    -75.77019, -74.8985, -74.01492, -73.12227, -72.22283, -71.31852, 
    -70.41093, -69.50142, -68.59113, -67.68102, -66.77197, -65.86467, 
    -64.95979, -64.05786, -63.15939, -62.26479, -61.37446, -60.48872, 
    -59.60787, -58.73216, -57.86184, -56.99708, -56.13808, -55.28499, 
    -54.43793, -53.59702, -52.76235, -51.934, -51.11204, -50.29652, 
    -49.48746, -48.68491, -47.88887, -47.09935, -46.31635, -45.53984, 
    -44.76982,
  -44.6996, -45.46576, -46.23822, -47.01697, -47.80202, -48.59336, -49.39099, 
    -50.19486, -51.00494, -51.82117, -52.64349, -53.47181, -54.30604, 
    -55.14605, -55.99172, -56.84288, -57.69935, -58.56092, -59.42736, 
    -60.29839, -61.17372, -62.05299, -62.93583, -63.82177, -64.71033, 
    -65.60093, -66.49293, -67.38558, -68.27805, -69.16933, -70.05833, 
    -70.9437, -71.8239, -72.69713, -73.56123, -74.41362, -75.25123, 
    -76.07032, -76.86639, -77.63395, -78.36636, -79.05556, -79.69198, 
    -80.2644, -80.76014, -81.16562, -81.46742, -81.65389, -81.71702, 
    -81.65389, -81.46742, -81.16562, -80.76014, -80.2644, -79.69198, 
    -79.05556, -78.36636, -77.63395, -76.86639, -76.07032, -75.25123, 
    -74.41362, -73.56123, -72.69713, -71.8239, -70.9437, -70.05833, 
    -69.16933, -68.27805, -67.38558, -66.49293, -65.60093, -64.71033, 
    -63.82177, -62.93583, -62.05299, -61.17372, -60.29839, -59.42736, 
    -58.56092, -57.69935, -56.84288, -55.99172, -55.14605, -54.30604, 
    -53.47181, -52.64349, -51.82117, -51.00494, -50.19486, -49.39099, 
    -48.59336, -47.80202, -47.01697, -46.23822, -45.46576, -44.6996,
  -44.62016, -45.38197, -46.14986, -46.92382, -47.70385, -48.48992, -49.282, 
    -50.08005, -50.88401, -51.69381, -52.50938, -53.33059, -54.15733, 
    -54.98947, -55.82684, -56.66924, -57.51648, -58.36829, -59.22443, 
    -60.08456, -60.94834, -61.81537, -62.6852, -63.55734, -64.4312, 
    -65.30614, -66.18141, -67.05619, -67.9295, -68.80025, -69.66718, 
    -70.52879, -71.38338, -72.22897, -73.06321, -73.88333, -74.68606, 
    -75.46753, -76.22314, -76.94742, -77.63395, -78.2752, -78.8625, 
    -79.38612, -79.83553, -80.19992, -80.46906, -80.6344, -80.69019, 
    -80.6344, -80.46906, -80.19992, -79.83553, -79.38612, -78.8625, -78.2752, 
    -77.63395, -76.94742, -76.22314, -75.46753, -74.68606, -73.88333, 
    -73.06321, -72.22897, -71.38338, -70.52879, -69.66718, -68.80025, 
    -67.9295, -67.05619, -66.18141, -65.30614, -64.4312, -63.55734, -62.6852, 
    -61.81537, -60.94834, -60.08456, -59.22443, -58.36829, -57.51648, 
    -56.66924, -55.82684, -54.98947, -54.15733, -53.33059, -52.50938, 
    -51.69381, -50.88401, -50.08005, -49.282, -48.48992, -47.70385, 
    -46.92382, -46.14986, -45.38197, -44.62016,
  -44.53154, -45.28852, -46.05135, -46.82, -47.59445, -48.37467, -49.16062, 
    -49.95222, -50.74942, -51.55212, -52.36022, -53.17359, -53.99209, 
    -54.81555, -55.64378, -56.47657, -57.31367, -58.1548, -58.99965, 
    -59.84786, -60.69904, -61.55275, -62.40846, -63.26563, -64.1236, 
    -64.98164, -65.83895, -66.69459, -67.54749, -68.39644, -69.24005, 
    -70.07672, -70.90462, -71.7216, -72.5252, -73.31252, -74.08022, 
    -74.82438, -75.54044, -76.22314, -76.86639, -77.46332, -78.00623, 
    -78.4868, -78.89631, -79.22611, -79.46831, -79.61646, -79.66634, 
    -79.61646, -79.46831, -79.22611, -78.89631, -78.4868, -78.00623, 
    -77.46332, -76.86639, -76.22314, -75.54044, -74.82438, -74.08022, 
    -73.31252, -72.5252, -71.7216, -70.90462, -70.07672, -69.24005, 
    -68.39644, -67.54749, -66.69459, -65.83895, -64.98164, -64.1236, 
    -63.26563, -62.40846, -61.55275, -60.69904, -59.84786, -58.99965, 
    -58.1548, -57.31367, -56.47657, -55.64378, -54.81555, -53.99209, 
    -53.17359, -52.36022, -51.55212, -50.74942, -49.95222, -49.16062, 
    -48.37467, -47.59445, -46.82, -46.05135, -45.28852, -44.53154,
  -44.4338, -45.18549, -45.94276, -46.70559, -47.47393, -48.24775, -49.02699, 
    -49.81155, -50.60136, -51.39631, -52.19627, -53.00109, -53.81061, 
    -54.62463, -55.44294, -56.26529, -57.09141, -57.92097, -58.75364, 
    -59.589, -60.42662, -61.26601, -62.10659, -62.94775, -63.78878, 
    -64.62888, -65.46716, -66.30258, -67.13403, -67.96017, -68.77954, 
    -69.59042, -70.39089, -71.17871, -71.95134, -72.70583, -73.43884, 
    -74.14648, -74.82438, -75.46753, -76.07032, -76.62655, -77.12947, 
    -77.572, -77.94691, -78.24726, -78.46685, -78.60075, -78.64574, 
    -78.60075, -78.46685, -78.24726, -77.94691, -77.572, -77.12947, 
    -76.62655, -76.07032, -75.46753, -74.82438, -74.14648, -73.43884, 
    -72.70583, -71.95134, -71.17871, -70.39089, -69.59042, -68.77954, 
    -67.96017, -67.13403, -66.30258, -65.46716, -64.62888, -63.78878, 
    -62.94775, -62.10659, -61.26601, -60.42662, -59.589, -58.75364, 
    -57.92097, -57.09141, -56.26529, -55.44294, -54.62463, -53.81061, 
    -53.00109, -52.19627, -51.39631, -50.60136, -49.81155, -49.02699, 
    -48.24775, -47.47393, -46.70559, -45.94276, -45.18549, -44.4338,
  -44.32701, -45.07294, -45.82418, -46.58068, -47.34241, -48.10929, 
    -48.88126, -49.6582, -50.44002, -51.22659, -52.01776, -52.81337, 
    -53.61321, -54.41708, -55.22473, -56.03588, -56.85022, -57.66741, 
    -58.48705, -59.30871, -60.1319, -60.95608, -61.78063, -62.60488, 
    -63.42805, -64.2493, -65.06765, -65.88202, -66.69118, -67.49377, 
    -68.28822, -69.07276, -69.84539, -70.60384, -71.34553, -72.06753, 
    -72.76654, -73.43884, -74.08022, -74.68606, -75.25123, -75.77019, 
    -76.23708, -76.64588, -76.99059, -77.26559, -77.46595, -77.58782, 
    -77.62873, -77.58782, -77.46595, -77.26559, -76.99059, -76.64588, 
    -76.23708, -75.77019, -75.25123, -74.68606, -74.08022, -73.43884, 
    -72.76654, -72.06753, -71.34553, -70.60384, -69.84539, -69.07276, 
    -68.28822, -67.49377, -66.69118, -65.88202, -65.06765, -64.2493, 
    -63.42805, -62.60488, -61.78063, -60.95608, -60.1319, -59.30871, 
    -58.48705, -57.66741, -56.85022, -56.03588, -55.22473, -54.41708, 
    -53.61321, -52.81337, -52.01776, -51.22659, -50.44002, -49.6582, 
    -48.88126, -48.10929, -47.34241, -46.58068, -45.82418, -45.07294, 
    -44.32701,
  -44.21122, -44.95095, -45.6957, -46.4454, -47.20001, -47.95944, -48.72359, 
    -49.49236, -50.26561, -51.04321, -51.82498, -52.61073, -53.40025, 
    -54.19329, -54.98958, -55.78882, -56.59066, -57.39472, -58.20058, 
    -59.00777, -59.81574, -60.62392, -61.43166, -62.2382, -63.04275, 
    -63.84439, -64.6421, -65.43473, -66.22101, -66.9995, -67.76861, -68.5265, 
    -69.27117, -70.00032, -70.7114, -71.40154, -72.06753, -72.70583, 
    -73.31252, -73.88333, -74.41362, -74.8985, -75.33289, -75.71165, 
    -76.02982, -76.28278, -76.46657, -76.57815, -76.61555, -76.57815, 
    -76.46657, -76.28278, -76.02982, -75.71165, -75.33289, -74.8985, 
    -74.41362, -73.88333, -73.31252, -72.70583, -72.06753, -71.40154, 
    -70.7114, -70.00032, -69.27117, -68.5265, -67.76861, -66.9995, -66.22101, 
    -65.43473, -64.6421, -63.84439, -63.04275, -62.2382, -61.43166, 
    -60.62392, -59.81574, -59.00777, -58.20058, -57.39472, -56.59066, 
    -55.78882, -54.98958, -54.19329, -53.40025, -52.61073, -51.82498, 
    -51.04321, -50.26561, -49.49236, -48.72359, -47.95944, -47.20001, 
    -46.4454, -45.6957, -44.95095, -44.21122,
  -44.08652, -44.81961, -45.55742, -46.29986, -47.04686, -47.79833, 
    -48.55416, -49.31422, -50.07836, -50.84642, -51.6182, -52.39351, 
    -53.17208, -53.95366, -54.73795, -55.52462, -56.31329, -57.10355, 
    -57.89494, -58.68696, -59.47903, -60.27053, -61.06076, -61.84895, 
    -62.63423, -63.41565, -64.19215, -64.96255, -65.72551, -66.47958, 
    -67.22313, -67.95432, -68.67112, -69.37128, -70.0523, -70.7114, 
    -71.34553, -71.95134, -72.5252, -73.06321, -73.56123, -74.01492, 
    -74.41991, -74.77181, -75.06647, -75.30009, -75.46947, -75.57212, 
    -75.60651, -75.57212, -75.46947, -75.30009, -75.06647, -74.77181, 
    -74.41991, -74.01492, -73.56123, -73.06321, -72.5252, -71.95134, 
    -71.34553, -70.7114, -70.0523, -69.37128, -68.67112, -67.95432, 
    -67.22313, -66.47958, -65.72551, -64.96255, -64.19215, -63.41565, 
    -62.63423, -61.84895, -61.06076, -60.27053, -59.47903, -58.68696, 
    -57.89494, -57.10355, -56.31329, -55.52462, -54.73795, -53.95366, 
    -53.17208, -52.39351, -51.6182, -50.84642, -50.07836, -49.31422, 
    -48.55416, -47.79833, -47.04686, -46.29986, -45.55742, -44.81961, 
    -44.08652,
  -43.95298, -44.67902, -45.40944, -46.14417, -46.8831, -47.62614, -48.37315, 
    -49.124, -49.8785, -50.63649, -51.39774, -52.16203, -52.92909, -53.69863, 
    -54.47033, -55.24382, -56.01871, -56.79456, -57.57087, -58.34711, 
    -59.12267, -59.89689, -60.66905, -61.43833, -62.20383, -62.96457, 
    -63.71946, -64.46726, -65.20666, -65.93615, -66.65411, -67.3587, 
    -68.04794, -68.7196, -69.37128, -70.00032, -70.60384, -71.17871, 
    -71.7216, -72.22897, -72.69713, -73.12227, -73.50058, -73.82835, 
    -74.10206, -74.31858, -74.47527, -74.57011, -74.60188, -74.57011, 
    -74.47527, -74.31858, -74.10206, -73.82835, -73.50058, -73.12227, 
    -72.69713, -72.22897, -71.7216, -71.17871, -70.60384, -70.00032, 
    -69.37128, -68.7196, -68.04794, -67.3587, -66.65411, -65.93615, 
    -65.20666, -64.46726, -63.71946, -62.96457, -62.20383, -61.43833, 
    -60.66905, -59.89689, -59.12267, -58.34711, -57.57087, -56.79456, 
    -56.01871, -55.24382, -54.47033, -53.69863, -52.92909, -52.16203, 
    -51.39774, -50.63649, -49.8785, -49.124, -48.37315, -47.62614, -46.8831, 
    -46.14417, -45.40944, -44.67902, -43.95298,
  -43.81068, -44.52925, -45.25187, -45.97845, -46.70888, -47.44304, 
    -48.18076, -48.92191, -49.66629, -50.4137, -51.1639, -51.91666, 
    -52.67167, -53.42863, -54.18719, -54.94697, -55.70753, -56.46842, 
    -57.22911, -57.98904, -58.74758, -59.50403, -60.25764, -61.00757, 
    -61.7529, -62.49262, -63.2256, -63.95062, -64.66634, -65.37125, 
    -66.06374, -66.74202, -67.40413, -68.04794, -68.67112, -69.27117, 
    -69.84539, -70.39089, -70.90462, -71.38338, -71.8239, -72.22283, 
    -72.57687, -72.88284, -73.13778, -73.33907, -73.4845, -73.57245, 
    -73.60188, -73.57245, -73.4845, -73.33907, -73.13778, -72.88284, 
    -72.57687, -72.22283, -71.8239, -71.38338, -70.90462, -70.39089, 
    -69.84539, -69.27117, -68.67112, -68.04794, -67.40413, -66.74202, 
    -66.06374, -65.37125, -64.66634, -63.95062, -63.2256, -62.49262, 
    -61.7529, -61.00757, -60.25764, -59.50403, -58.74758, -57.98904, 
    -57.22911, -56.46842, -55.70753, -54.94697, -54.18719, -53.42863, 
    -52.67167, -51.91666, -51.1639, -50.4137, -49.66629, -48.92191, 
    -48.18076, -47.44304, -46.70888, -45.97845, -45.25187, -44.52925, 
    -43.81068,
  -43.65969, -44.37041, -45.08484, -45.80286, -46.52436, -47.24918, 
    -47.97718, -48.70818, -49.44197, -50.17833, -50.91702, -51.65775, 
    -52.40023, -53.14412, -53.88906, -54.63462, -55.38037, -56.12582, 
    -56.87043, -57.61359, -58.35467, -59.09295, -59.82764, -60.55789, 
    -61.28276, -62.00122, -62.71215, -63.41431, -64.10636, -64.78683, 
    -65.45412, -66.10648, -66.74202, -67.3587, -67.95432, -68.5265, 
    -69.07276, -69.59042, -70.07672, -70.52879, -70.9437, -71.31852, 
    -71.6504, -71.9366, -72.17461, -72.36224, -72.49763, -72.57942, 
    -72.60679, -72.57942, -72.49763, -72.36224, -72.17461, -71.9366, 
    -71.6504, -71.31852, -70.9437, -70.52879, -70.07672, -69.59042, 
    -69.07276, -68.5265, -67.95432, -67.3587, -66.74202, -66.10648, 
    -65.45412, -64.78683, -64.10636, -63.41431, -62.71215, -62.00122, 
    -61.28276, -60.55789, -59.82764, -59.09295, -58.35467, -57.61359, 
    -56.87043, -56.12582, -55.38037, -54.63462, -53.88906, -53.14412, 
    -52.40023, -51.65775, -50.91702, -50.17833, -49.44197, -48.70818, 
    -47.97718, -47.24918, -46.52436, -45.80286, -45.08484, -44.37041, 
    -43.65969,
  -43.50012, -44.20261, -44.90845, -45.61752, -46.32969, -47.04478, 
    -47.76263, -48.48305, -49.20582, -49.9307, -50.65742, -51.38569, 
    -52.11519, -52.84557, -53.57643, -54.30735, -55.03786, -55.76746, 
    -56.49557, -57.2216, -57.94487, -58.66464, -59.38013, -60.09047, 
    -60.79469, -61.49178, -62.18061, -62.85994, -63.52847, -64.18473, 
    -64.82718, -65.45412, -66.06374, -66.65411, -67.22313, -67.76861, 
    -68.28822, -68.77954, -69.24005, -69.66718, -70.05833, -70.41093, 
    -70.72251, -70.99072, -71.21339, -71.38868, -71.51503, -71.59132, 
    -71.61682, -71.59132, -71.51503, -71.38868, -71.21339, -70.99072, 
    -70.72251, -70.41093, -70.05833, -69.66718, -69.24005, -68.77954, 
    -68.28822, -67.76861, -67.22313, -66.65411, -66.06374, -65.45412, 
    -64.82718, -64.18473, -63.52847, -62.85994, -62.18061, -61.49178, 
    -60.79469, -60.09047, -59.38013, -58.66464, -57.94487, -57.2216, 
    -56.49557, -55.76746, -55.03786, -54.30735, -53.57643, -52.84557, 
    -52.11519, -51.38569, -50.65742, -49.9307, -49.20582, -48.48305, 
    -47.76263, -47.04478, -46.32969, -45.61752, -44.90845, -44.20261, 
    -43.50012,
  -43.33206, -44.02596, -44.72285, -45.42259, -46.12503, -46.83001, 
    -47.53732, -48.24677, -48.95811, -49.6711, -50.38545, -51.10085, 
    -51.81697, -52.53343, -53.24984, -53.96573, -54.68064, -55.39402, 
    -56.10532, -56.8139, -57.51908, -58.22011, -58.9162, -59.60646, 
    -60.28995, -60.96564, -61.63241, -62.28906, -62.93428, -63.56667, 
    -64.18473, -64.78683, -65.37125, -65.93615, -66.47958, -66.9995, 
    -67.49377, -67.96017, -68.39644, -68.80025, -69.16933, -69.50142, 
    -69.79435, -70.04609, -70.2548, -70.4189, -70.53708, -70.60838, 
    -70.63222, -70.60838, -70.53708, -70.4189, -70.2548, -70.04609, 
    -69.79435, -69.50142, -69.16933, -68.80025, -68.39644, -67.96017, 
    -67.49377, -66.9995, -66.47958, -65.93615, -65.37125, -64.78683, 
    -64.18473, -63.56667, -62.93428, -62.28906, -61.63241, -60.96564, 
    -60.28995, -59.60646, -58.9162, -58.22011, -57.51908, -56.8139, 
    -56.10532, -55.39402, -54.68064, -53.96573, -53.24984, -52.53343, 
    -51.81697, -51.10085, -50.38545, -49.6711, -48.95811, -48.24677, 
    -47.53732, -46.83001, -46.12503, -45.42259, -44.72285, -44.02596, 
    -43.33206,
  -43.1556, -43.84056, -44.52815, -45.21821, -45.91058, -46.60506, -47.30147, 
    -47.99957, -48.69912, -49.39985, -50.10146, -50.80363, -51.506, -52.2082, 
    -52.9098, -53.61034, -54.30932, -55.00621, -55.70042, -56.39131, 
    -57.07819, -57.76032, -58.43688, -59.10701, -59.76975, -60.4241, 
    -61.06895, -61.70312, -62.32535, -62.93428, -63.52847, -64.10636, 
    -64.66634, -65.20666, -65.72551, -66.22101, -66.69118, -67.13403, 
    -67.54749, -67.9295, -68.27805, -68.59113, -68.86686, -69.10349, 
    -69.29943, -69.45333, -69.56409, -69.63087, -69.65318, -69.63087, 
    -69.56409, -69.45333, -69.29943, -69.10349, -68.86686, -68.59113, 
    -68.27805, -67.9295, -67.54749, -67.13403, -66.69118, -66.22101, 
    -65.72551, -65.20666, -64.66634, -64.10636, -63.52847, -62.93428, 
    -62.32535, -61.70312, -61.06895, -60.4241, -59.76975, -59.10701, 
    -58.43688, -57.76032, -57.07819, -56.39131, -55.70042, -55.00621, 
    -54.30932, -53.61034, -52.9098, -52.2082, -51.506, -50.80363, -50.10146, 
    -49.39985, -48.69912, -47.99957, -47.30147, -46.60506, -45.91058, 
    -45.21821, -44.52815, -43.84056, -43.1556,
  -42.97084, -43.64655, -44.3245, -45.00454, -45.68649, -46.37015, -47.05531, 
    -47.74172, -48.42913, -49.11726, -49.8058, -50.49441, -51.18272, 
    -51.87035, -52.55685, -53.24175, -53.92455, -54.60471, -55.28162, 
    -55.95465, -56.62309, -57.28621, -57.9432, -58.59319, -59.23526, 
    -59.86839, -60.49152, -61.1035, -61.70312, -62.28906, -62.85994, 
    -63.41431, -63.95062, -64.46726, -64.96255, -65.43473, -65.88202, 
    -66.30258, -66.69459, -67.05619, -67.38558, -67.68102, -67.94086, 
    -68.16358, -68.3478, -68.49236, -68.59633, -68.65899, -68.67992, 
    -68.65899, -68.59633, -68.49236, -68.3478, -68.16358, -67.94086, 
    -67.68102, -67.38558, -67.05619, -66.69459, -66.30258, -65.88202, 
    -65.43473, -64.96255, -64.46726, -63.95062, -63.41431, -62.85994, 
    -62.28906, -61.70312, -61.1035, -60.49152, -59.86839, -59.23526, 
    -58.59319, -57.9432, -57.28621, -56.62309, -55.95465, -55.28162, 
    -54.60471, -53.92455, -53.24175, -52.55685, -51.87035, -51.18272, 
    -50.49441, -49.8058, -49.11726, -48.42913, -47.74172, -47.05531, 
    -46.37015, -45.68649, -45.00454, -44.3245, -43.64655, -42.97084,
  -42.77788, -43.44402, -44.11203, -44.78174, -45.45296, -46.12547, 
    -46.79906, -47.47348, -48.14844, -48.82367, -49.49884, -50.1736, 
    -50.84757, -51.52035, -52.1915, -52.86054, -53.52696, -54.1902, 
    -54.84966, -55.50471, -56.15464, -56.79872, -57.43615, -58.06607, 
    -58.68758, -59.2997, -59.90138, -60.49152, -61.06895, -61.63241, 
    -62.18061, -62.71215, -63.2256, -63.71946, -64.19215, -64.6421, 
    -65.06765, -65.46716, -65.83895, -66.18141, -66.49293, -66.77197, 
    -67.01707, -67.22693, -67.40035, -67.53634, -67.63406, -67.69295, 
    -67.71262, -67.69295, -67.63406, -67.53634, -67.40035, -67.22693, 
    -67.01707, -66.77197, -66.49293, -66.18141, -65.83895, -65.46716, 
    -65.06765, -64.6421, -64.19215, -63.71946, -63.2256, -62.71215, 
    -62.18061, -61.63241, -61.06895, -60.49152, -59.90138, -59.2997, 
    -58.68758, -58.06607, -57.43615, -56.79872, -56.15464, -55.50471, 
    -54.84966, -54.1902, -53.52696, -52.86054, -52.1915, -51.52035, 
    -50.84757, -50.1736, -49.49884, -48.82367, -48.14844, -47.47348, 
    -46.79906, -46.12547, -45.45296, -44.78174, -44.11203, -43.44402, 
    -42.77788,
  -42.57683, -43.23311, -43.89089, -44.54997, -45.21016, -45.87124, 
    -46.53297, -47.1951, -47.85734, -48.51939, -49.18093, -49.84158, 
    -50.50098, -51.1587, -51.8143, -52.46729, -53.11716, -53.76335, 
    -54.40527, -55.04227, -55.67367, -56.29873, -56.91667, -57.52666, 
    -58.1278, -58.71915, -59.2997, -59.86839, -60.4241, -60.96564, -61.49178, 
    -62.00122, -62.49262, -62.96457, -63.41565, -63.84439, -64.2493, 
    -64.62888, -64.98164, -65.30614, -65.60093, -65.86467, -66.09609, 
    -66.29404, -66.45748, -66.58555, -66.67754, -66.73294, -66.75144, 
    -66.73294, -66.67754, -66.58555, -66.45748, -66.29404, -66.09609, 
    -65.86467, -65.60093, -65.30614, -64.98164, -64.62888, -64.2493, 
    -63.84439, -63.41565, -62.96457, -62.49262, -62.00122, -61.49178, 
    -60.96564, -60.4241, -59.86839, -59.2997, -58.71915, -58.1278, -57.52666, 
    -56.91667, -56.29873, -55.67367, -55.04227, -54.40527, -53.76335, 
    -53.11716, -52.46729, -51.8143, -51.1587, -50.50098, -49.84158, 
    -49.18093, -48.51939, -47.85734, -47.1951, -46.53297, -45.87124, 
    -45.21016, -44.54997, -43.89089, -43.23311, -42.57683,
  -42.36781, -43.01395, -43.66121, -44.30939, -44.95829, -45.60766, 
    -46.25727, -46.90686, -47.55613, -48.20476, -48.85243, -49.49877, 
    -50.14338, -50.78586, -51.42574, -52.06255, -52.69576, -53.32483, 
    -53.94915, -54.5681, -55.18099, -55.78711, -56.38568, -56.97591, 
    -57.55692, -58.1278, -58.68758, -59.23526, -59.76975, -60.28995, 
    -60.79469, -61.28276, -61.7529, -62.20383, -62.63423, -63.04275, 
    -63.42805, -63.78878, -64.1236, -64.4312, -64.71033, -64.95979, 
    -65.17846, -65.36533, -65.51952, -65.64027, -65.72695, -65.77914, 
    -65.79657, -65.77914, -65.72695, -65.64027, -65.51952, -65.36533, 
    -65.17846, -64.95979, -64.71033, -64.4312, -64.1236, -63.78878, 
    -63.42805, -63.04275, -62.63423, -62.20383, -61.7529, -61.28276, 
    -60.79469, -60.28995, -59.76975, -59.23526, -58.68758, -58.1278, 
    -57.55692, -56.97591, -56.38568, -55.78711, -55.18099, -54.5681, 
    -53.94915, -53.32483, -52.69576, -52.06255, -51.42574, -50.78586, 
    -50.14338, -49.49877, -48.85243, -48.20476, -47.55613, -46.90686, 
    -46.25727, -45.60766, -44.95829, -44.30939, -43.66121, -43.01395, 
    -42.36781,
  -42.15091, -42.78666, -43.42315, -44.06018, -44.69753, -45.33495, 
    -45.97221, -46.60902, -47.24509, -47.8801, -48.51371, -49.14555, 
    -49.77522, -50.40231, -51.02636, -51.64688, -52.26337, -52.87527, 
    -53.48199, -54.08292, -54.67738, -55.26468, -55.84407, -56.41476, 
    -56.97591, -57.52666, -58.06607, -58.59319, -59.10701, -59.60646, 
    -60.09047, -60.55789, -61.00757, -61.43833, -61.84895, -62.2382, 
    -62.60488, -62.94775, -63.26563, -63.55734, -63.82177, -64.05786, 
    -64.26463, -64.4412, -64.58678, -64.70073, -64.7825, -64.83172, 
    -64.84815, -64.83172, -64.7825, -64.70073, -64.58678, -64.4412, 
    -64.26463, -64.05786, -63.82177, -63.55734, -63.26563, -62.94775, 
    -62.60488, -62.2382, -61.84895, -61.43833, -61.00757, -60.55789, 
    -60.09047, -59.60646, -59.10701, -58.59319, -58.06607, -57.52666, 
    -56.97591, -56.41476, -55.84407, -55.26468, -54.67738, -54.08292, 
    -53.48199, -52.87527, -52.26337, -51.64688, -51.02636, -50.40231, 
    -49.77522, -49.14555, -48.51371, -47.8801, -47.24509, -46.60902, 
    -45.97221, -45.33495, -44.69753, -44.06018, -43.42315, -42.78666, 
    -42.15091,
  -41.92625, -42.55138, -43.17686, -43.8025, -44.42807, -45.05334, -45.67802, 
    -46.30186, -46.92454, -47.54575, -48.16513, -48.78232, -49.39692, 
    -50.00851, -50.61664, -51.22083, -51.82056, -52.4153, -53.00447, 
    -53.58745, -54.16361, -54.73225, -55.29266, -55.84407, -56.38568, 
    -56.91667, -57.43615, -57.9432, -58.43688, -58.9162, -59.38013, 
    -59.82764, -60.25764, -60.66905, -61.06076, -61.43166, -61.78063, 
    -62.10659, -62.40846, -62.6852, -62.93583, -63.15939, -63.35503, 
    -63.52198, -63.65955, -63.76716, -63.84436, -63.89082, -63.90633, 
    -63.89082, -63.84436, -63.76716, -63.65955, -63.52198, -63.35503, 
    -63.15939, -62.93583, -62.6852, -62.40846, -62.10659, -61.78063, 
    -61.43166, -61.06076, -60.66905, -60.25764, -59.82764, -59.38013, 
    -58.9162, -58.43688, -57.9432, -57.43615, -56.91667, -56.38568, 
    -55.84407, -55.29266, -54.73225, -54.16361, -53.58745, -53.00447, 
    -52.4153, -51.82056, -51.22083, -50.61664, -50.00851, -49.39692, 
    -48.78232, -48.16513, -47.54575, -46.92454, -46.30186, -45.67802, 
    -45.05334, -44.42807, -43.8025, -43.17686, -42.55138, -41.92625,
  -41.69396, -42.30823, -42.92249, -43.53653, -44.15013, -44.76302, 
    -45.37495, -45.98564, -46.59477, -47.20202, -47.80704, -48.40947, 
    -49.00891, -49.60493, -50.19709, -50.78492, -51.36792, -51.94554, 
    -52.51723, -53.08239, -53.64039, -54.19058, -54.73225, -55.26468, 
    -55.78711, -56.29873, -56.79872, -57.28621, -57.76032, -58.22011, 
    -58.66464, -59.09295, -59.50403, -59.89689, -60.27053, -60.62392, 
    -60.95608, -61.26601, -61.55275, -61.81537, -62.05299, -62.26479, 
    -62.45001, -62.60796, -62.73804, -62.83975, -62.91269, -62.95657, 
    -62.97122, -62.95657, -62.91269, -62.83975, -62.73804, -62.60796, 
    -62.45001, -62.26479, -62.05299, -61.81537, -61.55275, -61.26601, 
    -60.95608, -60.62392, -60.27053, -59.89689, -59.50403, -59.09295, 
    -58.66464, -58.22011, -57.76032, -57.28621, -56.79872, -56.29873, 
    -55.78711, -55.26468, -54.73225, -54.19058, -53.64039, -53.08239, 
    -52.51723, -51.94554, -51.36792, -50.78492, -50.19709, -49.60493, 
    -49.00891, -48.40947, -47.80704, -47.20202, -46.59477, -45.98564, 
    -45.37495, -44.76302, -44.15013, -43.53653, -42.92249, -42.30823, 
    -41.69396,
  -41.45414, -42.05735, -42.66019, -43.26245, -43.86388, -44.46423, 
    -45.06325, -45.66063, -46.25607, -46.84925, -47.43981, -48.02739, 
    -48.6116, -49.19202, -49.7682, -50.33969, -50.90599, -51.46657, -52.0209, 
    -52.56838, -53.10843, -53.64039, -54.16361, -54.67738, -55.18099, 
    -55.67367, -56.15464, -56.62309, -57.07819, -57.51908, -57.94487, 
    -58.35467, -58.74758, -59.12267, -59.47903, -59.81574, -60.1319, 
    -60.42662, -60.69904, -60.94834, -61.17372, -61.37446, -61.54989, 
    -61.6994, -61.82248, -61.91867, -61.98763, -62.02911, -62.04295, 
    -62.02911, -61.98763, -61.91867, -61.82248, -61.6994, -61.54989, 
    -61.37446, -61.17372, -60.94834, -60.69904, -60.42662, -60.1319, 
    -59.81574, -59.47903, -59.12267, -58.74758, -58.35467, -57.94487, 
    -57.51908, -57.07819, -56.62309, -56.15464, -55.67367, -55.18099, 
    -54.67738, -54.16361, -53.64039, -53.10843, -52.56838, -52.0209, 
    -51.46657, -50.90599, -50.33969, -49.7682, -49.19202, -48.6116, 
    -48.02739, -47.43981, -46.84925, -46.25607, -45.66063, -45.06325, 
    -44.46423, -43.86388, -43.26245, -42.66019, -42.05735, -41.45414,
  -41.20691, -41.79888, -42.39012, -42.98042, -43.56952, -44.15719, 
    -44.74314, -45.3271, -45.90874, -46.48775, -47.06378, -47.63646, 
    -48.20541, -48.77021, -49.33044, -49.88563, -50.43531, -50.97897, 
    -51.51608, -52.04608, -52.56838, -53.08239, -53.58745, -54.08292, 
    -54.5681, -55.04227, -55.50471, -55.95465, -56.39131, -56.8139, -57.2216, 
    -57.61359, -57.98904, -58.34711, -58.68696, -59.00777, -59.30871, 
    -59.589, -59.84786, -60.08456, -60.29839, -60.48872, -60.65495, 
    -60.79654, -60.91304, -61.00407, -61.06931, -61.10854, -61.12163, 
    -61.10854, -61.06931, -61.00407, -60.91304, -60.79654, -60.65495, 
    -60.48872, -60.29839, -60.08456, -59.84786, -59.589, -59.30871, 
    -59.00777, -58.68696, -58.34711, -57.98904, -57.61359, -57.2216, 
    -56.8139, -56.39131, -55.95465, -55.50471, -55.04227, -54.5681, 
    -54.08292, -53.58745, -53.08239, -52.56838, -52.04608, -51.51608, 
    -50.97897, -50.43531, -49.88563, -49.33044, -48.77021, -48.20541, 
    -47.63646, -47.06378, -46.48775, -45.90874, -45.3271, -44.74314, 
    -44.15719, -43.56952, -42.98042, -42.39012, -41.79888, -41.20691,
  -40.9524, -41.53295, -42.11243, -42.69062, -43.26726, -43.84211, -44.41489, 
    -44.98531, -45.55307, -46.11785, -46.67929, -47.23705, -47.79074, 
    -48.33995, -48.88427, -49.42325, -49.95642, -50.48329, -51.00336, 
    -51.51608, -52.0209, -52.51723, -53.00447, -53.48199, -53.94915, 
    -54.40527, -54.84966, -55.28162, -55.70042, -56.10532, -56.49557, 
    -56.87043, -57.22911, -57.57087, -57.89494, -58.20058, -58.48705, 
    -58.75364, -58.99965, -59.22443, -59.42736, -59.60787, -59.76543, 
    -59.89958, -60.00991, -60.09608, -60.15783, -60.19496, -60.20734, 
    -60.19496, -60.15783, -60.09608, -60.00991, -59.89958, -59.76543, 
    -59.60787, -59.42736, -59.22443, -58.99965, -58.75364, -58.48705, 
    -58.20058, -57.89494, -57.57087, -57.22911, -56.87043, -56.49557, 
    -56.10532, -55.70042, -55.28162, -54.84966, -54.40527, -53.94915, 
    -53.48199, -53.00447, -52.51723, -52.0209, -51.51608, -51.00336, 
    -50.48329, -49.95642, -49.42325, -48.88427, -48.33995, -47.79074, 
    -47.23705, -46.67929, -46.11785, -45.55307, -44.98531, -44.41489, 
    -43.84211, -43.26726, -42.69062, -42.11243, -41.53295, -40.9524,
  -40.69072, -41.25971, -41.82729, -42.39323, -42.95729, -43.51921, 
    -44.07872, -44.63554, -45.18936, -45.73986, -46.28671, -46.82954, 
    -47.36799, -47.90166, -48.43015, -48.95301, -49.46981, -49.98007, 
    -50.48329, -50.97897, -51.46657, -51.94554, -52.4153, -52.87527, 
    -53.32483, -53.76335, -54.1902, -54.60471, -55.00621, -55.39402, 
    -55.76746, -56.12582, -56.46842, -56.79456, -57.10355, -57.39472, 
    -57.66741, -57.92097, -58.1548, -58.36829, -58.56092, -58.73216, 
    -58.88156, -59.0087, -59.11322, -59.19484, -59.2533, -59.28845, 
    -59.30018, -59.28845, -59.2533, -59.19484, -59.11322, -59.0087, 
    -58.88156, -58.73216, -58.56092, -58.36829, -58.1548, -57.92097, 
    -57.66741, -57.39472, -57.10355, -56.79456, -56.46842, -56.12582, 
    -55.76746, -55.39402, -55.00621, -54.60471, -54.1902, -53.76335, 
    -53.32483, -52.87527, -52.4153, -51.94554, -51.46657, -50.97897, 
    -50.48329, -49.98007, -49.46981, -48.95301, -48.43015, -47.90166, 
    -47.36799, -46.82954, -46.28671, -45.73986, -45.18936, -44.63554, 
    -44.07872, -43.51921, -42.95729, -42.39323, -41.82729, -41.25971, 
    -40.69072,
  -40.42199, -40.97929, -41.53484, -42.08843, -42.6398, -43.18871, -43.73489, 
    -44.27805, -44.81789, -45.35409, -45.88634, -46.41428, -46.93754, 
    -47.45575, -47.96851, -48.4754, -48.97598, -49.46981, -49.95642, 
    -50.43531, -50.90599, -51.36792, -51.82056, -52.26337, -52.69576, 
    -53.11716, -53.52696, -53.92455, -54.30932, -54.68064, -55.03786, 
    -55.38037, -55.70753, -56.01871, -56.31329, -56.59066, -56.85022, 
    -57.09141, -57.31367, -57.51648, -57.69935, -57.86184, -58.00352, 
    -58.12405, -58.22311, -58.30043, -58.35581, -58.3891, -58.40021, 
    -58.3891, -58.35581, -58.30043, -58.22311, -58.12405, -58.00352, 
    -57.86184, -57.69935, -57.51648, -57.31367, -57.09141, -56.85022, 
    -56.59066, -56.31329, -56.01871, -55.70753, -55.38037, -55.03786, 
    -54.68064, -54.30932, -53.92455, -53.52696, -53.11716, -52.69576, 
    -52.26337, -51.82056, -51.36792, -50.90599, -50.43531, -49.95642, 
    -49.46981, -48.97598, -48.4754, -47.96851, -47.45575, -46.93754, 
    -46.41428, -45.88634, -45.35409, -44.81789, -44.27805, -43.73489, 
    -43.18871, -42.6398, -42.08843, -41.53484, -40.97929, -40.42199,
  -40.14635, -40.69183, -41.23525, -41.77639, -42.315, -42.85083, -43.38362, 
    -43.91308, -44.43893, -44.96085, -45.47853, -45.99162, -46.49977, 
    -47.00262, -47.49977, -47.99084, -48.4754, -48.95301, -49.42325, 
    -49.88563, -50.33969, -50.78492, -51.22083, -51.64688, -52.06255, 
    -52.46729, -52.86054, -53.24175, -53.61034, -53.96573, -54.30735, 
    -54.63462, -54.94697, -55.24382, -55.52462, -55.78882, -56.03588, 
    -56.26529, -56.47657, -56.66924, -56.84288, -56.99708, -57.13149, 
    -57.24578, -57.33968, -57.41296, -57.46543, -57.49697, -57.50749, 
    -57.49697, -57.46543, -57.41296, -57.33968, -57.24578, -57.13149, 
    -56.99708, -56.84288, -56.66924, -56.47657, -56.26529, -56.03588, 
    -55.78882, -55.52462, -55.24382, -54.94697, -54.63462, -54.30735, 
    -53.96573, -53.61034, -53.24175, -52.86054, -52.46729, -52.06255, 
    -51.64688, -51.22083, -50.78492, -50.33969, -49.88563, -49.42325, 
    -48.95301, -48.4754, -47.99084, -47.49977, -47.00262, -46.49977, 
    -45.99162, -45.47853, -44.96085, -44.43893, -43.91308, -43.38362, 
    -42.85083, -42.315, -41.77639, -41.23525, -40.69183, -40.14635,
  -39.8639, -40.39747, -40.92867, -41.45728, -41.98307, -42.50578, -43.02515, 
    -43.54091, -44.05278, -44.56044, -45.0636, -45.56192, -46.05505, 
    -46.54266, -47.02436, -47.49977, -47.96851, -48.43015, -48.88427, 
    -49.33044, -49.7682, -50.19709, -50.61664, -51.02636, -51.42574, 
    -51.8143, -52.1915, -52.55685, -52.9098, -53.24984, -53.57643, -53.88906, 
    -54.18719, -54.47033, -54.73795, -54.98958, -55.22473, -55.44294, 
    -55.64378, -55.82684, -55.99172, -56.13808, -56.26561, -56.374, 
    -56.46303, -56.53249, -56.58222, -56.6121, -56.62207, -56.6121, 
    -56.58222, -56.53249, -56.46303, -56.374, -56.26561, -56.13808, 
    -55.99172, -55.82684, -55.64378, -55.44294, -55.22473, -54.98958, 
    -54.73795, -54.47033, -54.18719, -53.88906, -53.57643, -53.24984, 
    -52.9098, -52.55685, -52.1915, -51.8143, -51.42574, -51.02636, -50.61664, 
    -50.19709, -49.7682, -49.33044, -48.88427, -48.43015, -47.96851, 
    -47.49977, -47.02436, -46.54266, -46.05505, -45.56192, -45.0636, 
    -44.56044, -44.05278, -43.54091, -43.02515, -42.50578, -41.98307, 
    -41.45728, -40.92867, -40.39747, -39.8639,
  -39.57478, -40.09635, -40.61526, -41.13129, -41.64421, -42.15377, 
    -42.65972, -43.16179, -43.6597, -44.15316, -44.64186, -45.1255, 
    -45.60374, -46.07624, -46.54266, -47.00262, -47.45575, -47.90166, 
    -48.33995, -48.77021, -49.19202, -49.60493, -50.00851, -50.40231, 
    -50.78586, -51.1587, -51.52035, -51.87035, -52.2082, -52.53343, 
    -52.84557, -53.14412, -53.42863, -53.69863, -53.95366, -54.19329, 
    -54.41708, -54.62463, -54.81555, -54.98947, -55.14605, -55.28499, 
    -55.40599, -55.50881, -55.59324, -55.65909, -55.70623, -55.73455, 
    -55.744, -55.73455, -55.70623, -55.65909, -55.59324, -55.50881, 
    -55.40599, -55.28499, -55.14605, -54.98947, -54.81555, -54.62463, 
    -54.41708, -54.19329, -53.95366, -53.69863, -53.42863, -53.14412, 
    -52.84557, -52.53343, -52.2082, -51.87035, -51.52035, -51.1587, 
    -50.78586, -50.40231, -50.00851, -49.60493, -49.19202, -48.77021, 
    -48.33995, -47.90166, -47.45575, -47.00262, -46.54266, -46.07624, 
    -45.60374, -45.1255, -44.64186, -44.15316, -43.6597, -43.16179, 
    -42.65972, -42.15377, -41.64421, -41.13129, -40.61526, -40.09635, 
    -39.57478,
  -39.27911, -39.78861, -40.29517, -40.79858, -41.29861, -41.79502, 
    -42.28755, -42.77596, -43.25996, -43.73928, -44.21362, -44.68269, 
    -45.14617, -45.60374, -46.05505, -46.49977, -46.93754, -47.36799, 
    -47.79074, -48.20541, -48.6116, -49.00891, -49.39692, -49.77522, 
    -50.14338, -50.50098, -50.84757, -51.18272, -51.506, -51.81697, 
    -52.11519, -52.40023, -52.67167, -52.92909, -53.17208, -53.40025, 
    -53.61321, -53.81061, -53.99209, -54.15733, -54.30604, -54.43793, 
    -54.55275, -54.6503, -54.73037, -54.79281, -54.8375, -54.86435, 
    -54.87331, -54.86435, -54.8375, -54.79281, -54.73037, -54.6503, 
    -54.55275, -54.43793, -54.30604, -54.15733, -53.99209, -53.81061, 
    -53.61321, -53.40025, -53.17208, -52.92909, -52.67167, -52.40023, 
    -52.11519, -51.81697, -51.506, -51.18272, -50.84757, -50.50098, 
    -50.14338, -49.77522, -49.39692, -49.00891, -48.6116, -48.20541, 
    -47.79074, -47.36799, -46.93754, -46.49977, -46.05505, -45.60374, 
    -45.14617, -44.68269, -44.21362, -43.73928, -43.25996, -42.77596, 
    -42.28755, -41.79502, -41.29861, -40.79858, -40.29517, -39.78861, 
    -39.27911,
  -38.977, -39.47439, -39.96857, -40.45934, -40.94647, -41.42973, -41.90887, 
    -42.38366, -42.85382, -43.31909, -43.77919, -44.23382, -44.68269, 
    -45.1255, -45.56192, -45.99162, -46.41428, -46.82954, -47.23705, 
    -47.63646, -48.02739, -48.40947, -48.78232, -49.14555, -49.49877, 
    -49.84158, -50.1736, -50.49441, -50.80363, -51.10085, -51.38569, 
    -51.65775, -51.91666, -52.16203, -52.39351, -52.61073, -52.81337, 
    -53.00109, -53.17359, -53.33059, -53.47181, -53.59702, -53.70599, 
    -53.79853, -53.87448, -53.93369, -53.97606, -54.00152, -54.01001, 
    -54.00152, -53.97606, -53.93369, -53.87448, -53.79853, -53.70599, 
    -53.59702, -53.47181, -53.33059, -53.17359, -53.00109, -52.81337, 
    -52.61073, -52.39351, -52.16203, -51.91666, -51.65775, -51.38569, 
    -51.10085, -50.80363, -50.49441, -50.1736, -49.84158, -49.49877, 
    -49.14555, -48.78232, -48.40947, -48.02739, -47.63646, -47.23705, 
    -46.82954, -46.41428, -45.99162, -45.56192, -45.1255, -44.68269, 
    -44.23382, -43.77919, -43.31909, -42.85382, -42.38366, -41.90887, 
    -41.42973, -40.94647, -40.45934, -39.96857, -39.47439, -38.977,
  -38.66859, -39.15382, -39.6356, -40.11372, -40.58796, -41.0581, -41.52391, 
    -41.98514, -42.44154, -42.89287, -43.33884, -43.77919, -44.21362, 
    -44.64186, -45.0636, -45.47853, -45.88634, -46.28671, -46.67929, 
    -47.06378, -47.43981, -47.80704, -48.16513, -48.51371, -48.85243, 
    -49.18093, -49.49884, -49.8058, -50.10146, -50.38545, -50.65742, 
    -50.91702, -51.1639, -51.39774, -51.6182, -51.82498, -52.01776, 
    -52.19627, -52.36022, -52.50938, -52.64349, -52.76235, -52.86576, 
    -52.95356, -53.0256, -53.08176, -53.12194, -53.14607, -53.15412, 
    -53.14607, -53.12194, -53.08176, -53.0256, -52.95356, -52.86576, 
    -52.76235, -52.64349, -52.50938, -52.36022, -52.19627, -52.01776, 
    -51.82498, -51.6182, -51.39774, -51.1639, -50.91702, -50.65742, 
    -50.38545, -50.10146, -49.8058, -49.49884, -49.18093, -48.85243, 
    -48.51371, -48.16513, -47.80704, -47.43981, -47.06378, -46.67929, 
    -46.28671, -45.88634, -45.47853, -45.0636, -44.64186, -44.21362, 
    -43.77919, -43.33884, -42.89287, -42.44154, -41.98514, -41.52391, 
    -41.0581, -40.58796, -40.11372, -39.6356, -39.15382, -38.66859,
  -38.354, -38.82706, -39.29642, -39.7619, -40.22328, -40.68035, -41.13287, 
    -41.58063, -42.02338, -42.46088, -42.89287, -43.31909, -43.73928, 
    -44.15316, -44.56044, -44.96085, -45.35409, -45.73986, -46.11785, 
    -46.48775, -46.84925, -47.20202, -47.54575, -47.8801, -48.20476, 
    -48.51939, -48.82367, -49.11726, -49.39985, -49.6711, -49.9307, 
    -50.17833, -50.4137, -50.63649, -50.84642, -51.04321, -51.22659, 
    -51.39631, -51.55212, -51.69381, -51.82117, -51.934, -52.03214, 
    -52.11544, -52.18378, -52.23703, -52.27514, -52.29802, -52.30565, 
    -52.29802, -52.27514, -52.23703, -52.18378, -52.11544, -52.03214, 
    -51.934, -51.82117, -51.69381, -51.55212, -51.39631, -51.22659, 
    -51.04321, -50.84642, -50.63649, -50.4137, -50.17833, -49.9307, -49.6711, 
    -49.39985, -49.11726, -48.82367, -48.51939, -48.20476, -47.8801, 
    -47.54575, -47.20202, -46.84925, -46.48775, -46.11785, -45.73986, 
    -45.35409, -44.96085, -44.56044, -44.15316, -43.73928, -43.31909, 
    -42.89287, -42.46088, -42.02338, -41.58063, -41.13287, -40.68035, 
    -40.22328, -39.7619, -39.29642, -38.82706, -38.354,
  -38.03334, -38.49422, -38.95119, -39.40405, -39.85261, -40.29666, 
    -40.73598, -41.17037, -41.59958, -42.02338, -42.44154, -42.85382, 
    -43.25996, -43.6597, -44.05278, -44.43893, -44.81789, -45.18936, 
    -45.55307, -45.90874, -46.25607, -46.59477, -46.92454, -47.24509, 
    -47.55613, -47.85734, -48.14844, -48.42913, -48.69912, -48.95811, 
    -49.20582, -49.44197, -49.66629, -49.8785, -50.07836, -50.26561, 
    -50.44002, -50.60136, -50.74942, -50.88401, -51.00494, -51.11204, 
    -51.20517, -51.2842, -51.34902, -51.39953, -51.43566, -51.45736, 
    -51.46459, -51.45736, -51.43566, -51.39953, -51.34902, -51.2842, 
    -51.20517, -51.11204, -51.00494, -50.88401, -50.74942, -50.60136, 
    -50.44002, -50.26561, -50.07836, -49.8785, -49.66629, -49.44197, 
    -49.20582, -48.95811, -48.69912, -48.42913, -48.14844, -47.85734, 
    -47.55613, -47.24509, -46.92454, -46.59477, -46.25607, -45.90874, 
    -45.55307, -45.18936, -44.81789, -44.43893, -44.05278, -43.6597, 
    -43.25996, -42.85382, -42.44154, -42.02338, -41.59958, -41.17037, 
    -40.73598, -40.29666, -39.85261, -39.40405, -38.95119, -38.49422, 
    -38.03334,
  -37.70675, -38.15546, -38.60004, -39.04033, -39.47613, -39.90724, 
    -40.33345, -40.75457, -41.17037, -41.58063, -41.98514, -42.38366, 
    -42.77596, -43.16179, -43.54091, -43.91308, -44.27805, -44.63554, 
    -44.98531, -45.3271, -45.66063, -45.98564, -46.30186, -46.60902, 
    -46.90686, -47.1951, -47.47348, -47.74172, -47.99957, -48.24677, 
    -48.48305, -48.70818, -48.92191, -49.124, -49.31422, -49.49236, -49.6582, 
    -49.81155, -49.95222, -50.08005, -50.19486, -50.29652, -50.38489, 
    -50.45986, -50.52134, -50.56924, -50.6035, -50.62407, -50.63093, 
    -50.62407, -50.6035, -50.56924, -50.52134, -50.45986, -50.38489, 
    -50.29652, -50.19486, -50.08005, -49.95222, -49.81155, -49.6582, 
    -49.49236, -49.31422, -49.124, -48.92191, -48.70818, -48.48305, 
    -48.24677, -47.99957, -47.74172, -47.47348, -47.1951, -46.90686, 
    -46.60902, -46.30186, -45.98564, -45.66063, -45.3271, -44.98531, 
    -44.63554, -44.27805, -43.91308, -43.54091, -43.16179, -42.77596, 
    -42.38366, -41.98514, -41.58063, -41.17037, -40.75457, -40.33345, 
    -39.90724, -39.47613, -39.04033, -38.60004, -38.15546, -37.70675,
  -37.37434, -37.81089, -38.24314, -38.67091, -39.09401, -39.51227, 
    -39.92548, -40.33345, -40.73598, -41.13287, -41.52391, -41.90887, 
    -42.28755, -42.65972, -43.02515, -43.38362, -43.73489, -44.07872, 
    -44.41489, -44.74314, -45.06325, -45.37495, -45.67802, -45.97221, 
    -46.25727, -46.53297, -46.79906, -47.05531, -47.30147, -47.53732, 
    -47.76263, -47.97718, -48.18076, -48.37315, -48.55416, -48.72359, 
    -48.88126, -49.02699, -49.16062, -49.282, -49.39099, -49.48746, 
    -49.57131, -49.64243, -49.70073, -49.74615, -49.77864, -49.79815, 
    -49.80465, -49.79815, -49.77864, -49.74615, -49.70073, -49.64243, 
    -49.57131, -49.48746, -49.39099, -49.282, -49.16062, -49.02699, 
    -48.88126, -48.72359, -48.55416, -48.37315, -48.18076, -47.97718, 
    -47.76263, -47.53732, -47.30147, -47.05531, -46.79906, -46.53297, 
    -46.25727, -45.97221, -45.67802, -45.37495, -45.06325, -44.74314, 
    -44.41489, -44.07872, -43.73489, -43.38362, -43.02515, -42.65972, 
    -42.28755, -41.90887, -41.52391, -41.13287, -40.73598, -40.33345, 
    -39.92548, -39.51227, -39.09401, -38.67091, -38.24314, -37.81089, 
    -37.37434,
  -37.03624, -37.46067, -37.88063, -38.29594, -38.70644, -39.11194, 
    -39.51227, -39.90724, -40.29666, -40.68035, -41.0581, -41.42973, 
    -41.79502, -42.15377, -42.50578, -42.85083, -43.18871, -43.51921, 
    -43.84211, -44.15719, -44.46423, -44.76302, -45.05334, -45.33495, 
    -45.60766, -45.87124, -46.12547, -46.37015, -46.60506, -46.83001, 
    -47.04478, -47.24918, -47.44304, -47.62614, -47.79833, -47.95944, 
    -48.10929, -48.24775, -48.37467, -48.48992, -48.59336, -48.68491, 
    -48.76445, -48.83191, -48.8872, -48.93027, -48.96106, -48.97956, 
    -48.98572, -48.97956, -48.96106, -48.93027, -48.8872, -48.83191, 
    -48.76445, -48.68491, -48.59336, -48.48992, -48.37467, -48.24775, 
    -48.10929, -47.95944, -47.79833, -47.62614, -47.44304, -47.24918, 
    -47.04478, -46.83001, -46.60506, -46.37015, -46.12547, -45.87124, 
    -45.60766, -45.33495, -45.05334, -44.76302, -44.46423, -44.15719, 
    -43.84211, -43.51921, -43.18871, -42.85083, -42.50578, -42.15377, 
    -41.79502, -41.42973, -41.0581, -40.68035, -40.29666, -39.90724, 
    -39.51227, -39.11194, -38.70644, -38.29594, -37.88063, -37.46067, 
    -37.03624,
  -36.69255, -37.10492, -37.51265, -37.91559, -38.31358, -38.70644, 
    -39.09401, -39.47613, -39.85261, -40.22328, -40.58796, -40.94647, 
    -41.29861, -41.64421, -41.98307, -42.315, -42.6398, -42.95729, -43.26726, 
    -43.56952, -43.86388, -44.15013, -44.42807, -44.69753, -44.95829, 
    -45.21016, -45.45296, -45.68649, -45.91058, -46.12503, -46.32969, 
    -46.52436, -46.70888, -46.8831, -47.04686, -47.20001, -47.34241, 
    -47.47393, -47.59445, -47.70385, -47.80202, -47.88887, -47.96432, 
    -48.02829, -48.08072, -48.12155, -48.15074, -48.16827, -48.17411, 
    -48.16827, -48.15074, -48.12155, -48.08072, -48.02829, -47.96432, 
    -47.88887, -47.80202, -47.70385, -47.59445, -47.47393, -47.34241, 
    -47.20001, -47.04686, -46.8831, -46.70888, -46.52436, -46.32969, 
    -46.12503, -45.91058, -45.68649, -45.45296, -45.21016, -44.95829, 
    -44.69753, -44.42807, -44.15013, -43.86388, -43.56952, -43.26726, 
    -42.95729, -42.6398, -42.315, -41.98307, -41.64421, -41.29861, -40.94647, 
    -40.58796, -40.22328, -39.85261, -39.47613, -39.09401, -38.70644, 
    -38.31358, -37.91559, -37.51265, -37.10492, -36.69255,
  -36.34341, -36.74377, -37.13935, -37.53001, -37.91559, -38.29594, 
    -38.67091, -39.04033, -39.40405, -39.7619, -40.11372, -40.45934, 
    -40.79858, -41.13129, -41.45728, -41.77639, -42.08843, -42.39323, 
    -42.69062, -42.98042, -43.26245, -43.53653, -43.8025, -44.06018, 
    -44.30939, -44.54997, -44.78174, -45.00454, -45.21821, -45.42259, 
    -45.61752, -45.80286, -45.97845, -46.14417, -46.29986, -46.4454, 
    -46.58068, -46.70559, -46.82, -46.92382, -47.01697, -47.09935, -47.17091, 
    -47.23156, -47.28126, -47.31997, -47.34763, -47.36425, -47.36979, 
    -47.36425, -47.34763, -47.31997, -47.28126, -47.23156, -47.17091, 
    -47.09935, -47.01697, -46.92382, -46.82, -46.70559, -46.58068, -46.4454, 
    -46.29986, -46.14417, -45.97845, -45.80286, -45.61752, -45.42259, 
    -45.21821, -45.00454, -44.78174, -44.54997, -44.30939, -44.06018, 
    -43.8025, -43.53653, -43.26245, -42.98042, -42.69062, -42.39323, 
    -42.08843, -41.77639, -41.45728, -41.13129, -40.79858, -40.45934, 
    -40.11372, -39.7619, -39.40405, -39.04033, -38.67091, -38.29594, 
    -37.91559, -37.53001, -37.13935, -36.74377, -36.34341,
  -35.98892, -36.37735, -36.76087, -37.13935, -37.51265, -37.88063, 
    -38.24314, -38.60004, -38.95119, -39.29642, -39.6356, -39.96857, 
    -40.29517, -40.61526, -40.92867, -41.23525, -41.53484, -41.82729, 
    -42.11243, -42.39012, -42.66019, -42.92249, -43.17686, -43.42315, 
    -43.66121, -43.89089, -44.11203, -44.3245, -44.52815, -44.72285, 
    -44.90845, -45.08484, -45.25187, -45.40944, -45.55742, -45.6957, 
    -45.82418, -45.94276, -46.05135, -46.14986, -46.23822, -46.31635, 
    -46.38419, -46.44169, -46.4888, -46.52548, -46.5517, -46.56744, 
    -46.57269, -46.56744, -46.5517, -46.52548, -46.4888, -46.44169, 
    -46.38419, -46.31635, -46.23822, -46.14986, -46.05135, -45.94276, 
    -45.82418, -45.6957, -45.55742, -45.40944, -45.25187, -45.08484, 
    -44.90845, -44.72285, -44.52815, -44.3245, -44.11203, -43.89089, 
    -43.66121, -43.42315, -43.17686, -42.92249, -42.66019, -42.39012, 
    -42.11243, -41.82729, -41.53484, -41.23525, -40.92867, -40.61526, 
    -40.29517, -39.96857, -39.6356, -39.29642, -38.95119, -38.60004, 
    -38.24314, -37.88063, -37.51265, -37.13935, -36.76087, -36.37735, 
    -35.98892,
  -35.62921, -36.00579, -36.37735, -36.74377, -37.10492, -37.46067, 
    -37.81089, -38.15546, -38.49422, -38.82706, -39.15382, -39.47439, 
    -39.78861, -40.09635, -40.39747, -40.69183, -40.97929, -41.25971, 
    -41.53295, -41.79888, -42.05735, -42.30823, -42.55138, -42.78666, 
    -43.01395, -43.23311, -43.44402, -43.64655, -43.84056, -44.02596, 
    -44.20261, -44.37041, -44.52925, -44.67902, -44.81961, -44.95095, 
    -45.07294, -45.18549, -45.28852, -45.38197, -45.46576, -45.53984, 
    -45.60415, -45.65865, -45.7033, -45.73805, -45.7629, -45.77781, 
    -45.78278, -45.77781, -45.7629, -45.73805, -45.7033, -45.65865, 
    -45.60415, -45.53984, -45.46576, -45.38197, -45.28852, -45.18549, 
    -45.07294, -44.95095, -44.81961, -44.67902, -44.52925, -44.37041, 
    -44.20261, -44.02596, -43.84056, -43.64655, -43.44402, -43.23311, 
    -43.01395, -42.78666, -42.55138, -42.30823, -42.05735, -41.79888, 
    -41.53295, -41.25971, -40.97929, -40.69183, -40.39747, -40.09635, 
    -39.78861, -39.47439, -39.15382, -38.82706, -38.49422, -38.15546, 
    -37.81089, -37.46067, -37.10492, -36.74377, -36.37735, -36.00579, 
    -35.62921,
  -35.26439, -35.62921, -35.98892, -36.34341, -36.69255, -37.03624, 
    -37.37434, -37.70675, -38.03334, -38.354, -38.66859, -38.977, -39.27911, 
    -39.57478, -39.8639, -40.14635, -40.42199, -40.69072, -40.9524, 
    -41.20691, -41.45414, -41.69396, -41.92625, -42.15091, -42.36781, 
    -42.57683, -42.77788, -42.97084, -43.1556, -43.33206, -43.50012, 
    -43.65969, -43.81068, -43.95298, -44.08652, -44.21122, -44.32701, 
    -44.4338, -44.53154, -44.62016, -44.6996, -44.76982, -44.83077, 
    -44.88241, -44.9247, -44.95763, -44.98116, -44.99529, -45, -44.99529, 
    -44.98116, -44.95763, -44.9247, -44.88241, -44.83077, -44.76982, 
    -44.6996, -44.62016, -44.53154, -44.4338, -44.32701, -44.21122, 
    -44.08652, -43.95298, -43.81068, -43.65969, -43.50012, -43.33206, 
    -43.1556, -42.97084, -42.77788, -42.57683, -42.36781, -42.15091, 
    -41.92625, -41.69396, -41.45414, -41.20691, -40.9524, -40.69072, 
    -40.42199, -40.14635, -39.8639, -39.57478, -39.27911, -38.977, -38.66859, 
    -38.354, -38.03334, -37.70675, -37.37434, -37.03624, -36.69255, 
    -36.34341, -35.98892, -35.62921, -35.26439 ;

 grid_lont =
  215, 214.2135, 213.4195, 212.618, 211.8089, 210.9922, 210.1678, 209.3358, 
    208.4959, 207.6484, 206.793, 205.9299, 205.059, 204.1803, 203.2939, 
    202.3998, 201.498, 200.5886, 199.6716, 198.7471, 197.8153, 196.8762, 
    195.9299, 194.9766, 194.0163, 193.0493, 192.0756, 191.0956, 190.1093, 
    189.117, 188.1189, 187.1152, 186.1061, 185.0919, 184.073, 183.0495, 
    182.0217, 180.9899, 179.9545, 178.9158, 177.8741, 176.8297, 175.7829, 
    174.7342, 173.6839, 172.6322, 171.5797, 170.5266, 169.4734, 168.4203, 
    167.3678, 166.3161, 165.2658, 164.2171, 163.1703, 162.1259, 161.0842, 
    160.0455, 159.0101, 157.9783, 156.9505, 155.927, 154.9081, 153.8939, 
    152.8848, 151.8811, 150.883, 149.8907, 148.9044, 147.9244, 146.9507, 
    145.9837, 145.0234, 144.0701, 143.1238, 142.1847, 141.2529, 140.3284, 
    139.4114, 138.502, 137.6002, 136.7061, 135.8197, 134.941, 134.0701, 
    133.207, 132.3516, 131.5041, 130.6642, 129.8322, 129.0078, 128.1911, 
    127.382, 126.5805, 125.7865, 125,
  215.7865, 215, 214.2054, 213.4027, 212.5918, 211.7726, 210.945, 210.1091, 
    209.2647, 208.4118, 207.5504, 206.6805, 205.8021, 204.9151, 204.0196, 
    203.1156, 202.2032, 201.2823, 200.353, 199.4154, 198.4696, 197.5157, 
    196.5538, 195.584, 194.6065, 193.6215, 192.629, 191.6293, 190.6226, 
    189.6091, 188.589, 187.5627, 186.5303, 185.4922, 184.4486, 183.3998, 
    182.3462, 181.2881, 180.2259, 179.1599, 178.0904, 177.0179, 175.9428, 
    174.8654, 173.7861, 172.7054, 171.6237, 170.5413, 169.4587, 168.3763, 
    167.2946, 166.2139, 165.1346, 164.0572, 162.9821, 161.9096, 160.8401, 
    159.7741, 158.7119, 157.6538, 156.6002, 155.5514, 154.5078, 153.4697, 
    152.4373, 151.411, 150.3909, 149.3774, 148.3707, 147.371, 146.3785, 
    145.3935, 144.416, 143.4462, 142.4843, 141.5304, 140.5846, 139.647, 
    138.7177, 137.7968, 136.8844, 135.9804, 135.0849, 134.1979, 133.3195, 
    132.4496, 131.5882, 130.7353, 129.8909, 129.055, 128.2274, 127.4082, 
    126.5973, 125.7946, 125, 124.2135,
  216.5805, 215.7946, 215, 214.1967, 213.3845, 212.5633, 211.7332, 210.8939, 
    210.0455, 209.1879, 208.3211, 207.4449, 206.5594, 205.6646, 204.7604, 
    203.8469, 202.9241, 201.992, 201.0507, 200.1002, 199.1406, 198.1721, 
    197.1947, 196.2085, 195.2137, 194.2104, 193.1989, 192.1794, 191.152, 
    190.117, 189.0746, 188.0251, 186.9689, 185.9062, 184.8373, 183.7626, 
    182.6824, 181.5972, 180.5072, 179.413, 178.3148, 177.2133, 176.1087, 
    175.0016, 173.8923, 172.7814, 171.6693, 170.5565, 169.4435, 168.3307, 
    167.2186, 166.1077, 164.9984, 163.8913, 162.7867, 161.6852, 160.587, 
    159.4928, 158.4028, 157.3176, 156.2374, 155.1627, 154.0938, 153.0311, 
    151.9749, 150.9254, 149.883, 148.848, 147.8206, 146.8011, 145.7896, 
    144.7863, 143.7915, 142.8053, 141.8279, 140.8594, 139.8998, 138.9493, 
    138.008, 137.0759, 136.1531, 135.2396, 134.3354, 133.4406, 132.5551, 
    131.6789, 130.8121, 129.9545, 129.1061, 128.2668, 127.4367, 126.6155, 
    125.8033, 125, 124.2054, 123.4195,
  217.382, 216.5973, 215.8033, 215, 214.1872, 213.3647, 212.5326, 211.6906, 
    210.8388, 209.977, 209.1052, 208.2233, 207.3313, 206.4291, 205.5167, 
    204.5941, 203.6614, 202.7184, 201.7654, 200.8022, 199.8291, 198.846, 
    197.8531, 196.8506, 195.8385, 194.817, 193.7864, 192.7467, 191.6984, 
    190.6415, 189.5764, 188.5033, 187.4227, 186.3348, 185.2399, 184.1385, 
    183.031, 181.9177, 180.7991, 179.6757, 178.5479, 177.4162, 176.2811, 
    175.1431, 174.0027, 172.8604, 171.7168, 170.5723, 169.4277, 168.2832, 
    167.1396, 165.9973, 164.8569, 163.7189, 162.5838, 161.4521, 160.3243, 
    159.2009, 158.0823, 156.969, 155.8615, 154.7601, 153.6652, 152.5773, 
    151.4967, 150.4236, 149.3585, 148.3016, 147.2533, 146.2136, 145.183, 
    144.1615, 143.1494, 142.1469, 141.154, 140.1709, 139.1978, 138.2346, 
    137.2816, 136.3386, 135.4059, 134.4833, 133.5709, 132.6687, 131.7767, 
    130.8948, 130.023, 129.1612, 128.3094, 127.4674, 126.6353, 125.8128, 125, 
    124.1967, 123.4027, 122.618,
  218.1911, 217.4082, 216.6155, 215.8128, 215, 214.1769, 213.3434, 212.4994, 
    211.6447, 210.7794, 209.9032, 209.0162, 208.1181, 207.2091, 206.289, 
    205.3578, 204.4155, 203.4621, 202.4977, 201.5221, 200.5357, 199.5383, 
    198.5301, 197.5113, 196.4819, 195.4421, 194.3922, 193.3323, 192.2627, 
    191.1836, 190.0953, 188.9982, 187.8926, 186.7789, 185.6573, 184.5285, 
    183.3927, 182.2505, 181.1024, 179.9487, 178.7902, 177.6272, 176.4604, 
    175.2903, 174.1175, 172.9426, 171.7661, 170.5888, 169.4112, 168.2339, 
    167.0574, 165.8825, 164.7097, 163.5396, 162.3728, 161.2098, 160.0513, 
    158.8976, 157.7495, 156.6073, 155.4715, 154.3427, 153.2211, 152.1074, 
    151.0018, 149.9047, 148.8164, 147.7373, 146.6677, 145.6078, 144.5579, 
    143.5181, 142.4887, 141.4699, 140.4617, 139.4643, 138.4779, 137.5023, 
    136.5379, 135.5845, 134.6422, 133.711, 132.7909, 131.8819, 130.9838, 
    130.0968, 129.2206, 128.3553, 127.5006, 126.6566, 125.8231, 125, 
    124.1872, 123.3845, 122.5918, 121.8089,
  219.0078, 218.2274, 217.4367, 216.6353, 215.8231, 215, 214.1658, 213.3204, 
    212.4636, 211.5953, 210.7154, 209.8238, 208.9203, 208.005, 207.0777, 
    206.1384, 205.1871, 204.2236, 203.2482, 202.2607, 201.2611, 200.2497, 
    199.2264, 198.1913, 197.1447, 196.0866, 195.0173, 193.937, 192.8458, 
    191.7442, 190.6324, 189.5108, 188.3796, 187.2394, 186.0905, 184.9334, 
    183.7685, 182.5964, 181.4176, 180.2327, 179.0422, 177.8468, 176.647, 
    175.4436, 174.2371, 173.0282, 171.8176, 170.606, 169.394, 168.1824, 
    166.9718, 165.7629, 164.5564, 163.353, 162.1532, 160.9578, 159.7673, 
    158.5824, 157.4036, 156.2315, 155.0666, 153.9095, 152.7606, 151.6204, 
    150.4892, 149.3676, 148.2558, 147.1542, 146.063, 144.9827, 143.9134, 
    142.8553, 141.8087, 140.7736, 139.7503, 138.7389, 137.7393, 136.7518, 
    135.7764, 134.8129, 133.8616, 132.9223, 131.995, 131.0797, 130.1762, 
    129.2846, 128.4047, 127.5364, 126.6796, 125.8342, 125, 124.1769, 
    123.3647, 122.5633, 121.7725, 120.9922,
  219.8322, 219.055, 218.2668, 217.4674, 216.6566, 215.8342, 215, 214.1539, 
    213.2956, 212.425, 211.5421, 210.6465, 209.7383, 208.8173, 207.8834, 
    206.9366, 205.9767, 205.0037, 204.0176, 203.0185, 202.0062, 200.981, 
    199.9427, 198.8916, 197.8278, 196.7515, 195.6627, 194.5618, 193.4489, 
    192.3245, 191.1887, 190.042, 188.8848, 187.7174, 186.5403, 185.3541, 
    184.1592, 182.9563, 181.7458, 180.5284, 179.3048, 178.0757, 176.8416, 
    175.6034, 174.3618, 173.1175, 171.8713, 170.6239, 169.3761, 168.1287, 
    166.8825, 165.6382, 164.3966, 163.1584, 161.9243, 160.6952, 159.4716, 
    158.2542, 157.0437, 155.8408, 154.6459, 153.4597, 152.2826, 151.1152, 
    149.958, 148.8113, 147.6755, 146.5511, 145.4382, 144.3373, 143.2485, 
    142.1722, 141.1084, 140.0573, 139.019, 137.9938, 136.9815, 135.9824, 
    134.9963, 134.0233, 133.0634, 132.1166, 131.1827, 130.2617, 129.3535, 
    128.4579, 127.575, 126.7044, 125.8461, 125, 124.1658, 123.3434, 122.5326, 
    121.7332, 120.945, 120.1678,
  220.6642, 219.8909, 219.1061, 218.3094, 217.5006, 216.6796, 215.8461, 215, 
    214.141, 213.2689, 212.3836, 211.4848, 210.5725, 209.6465, 208.7066, 
    207.7528, 206.7849, 205.8029, 204.8067, 203.7964, 202.7718, 201.733, 
    200.6802, 199.6132, 198.5324, 197.4377, 196.3295, 195.2078, 194.0731, 
    192.9255, 191.7654, 190.5931, 189.4092, 188.214, 187.008, 185.7918, 
    184.5659, 183.331, 182.0877, 180.8367, 179.5787, 178.3145, 177.0447, 
    175.7703, 174.4921, 173.2108, 171.9273, 170.6426, 169.3574, 168.0727, 
    166.7892, 165.5079, 164.2297, 162.9553, 161.6855, 160.4213, 159.1633, 
    157.9123, 156.669, 155.4341, 154.2082, 152.992, 151.786, 150.5908, 
    149.4069, 148.2346, 147.0745, 145.9269, 144.7922, 143.6705, 142.5623, 
    141.4676, 140.3868, 139.3198, 138.267, 137.2282, 136.2036, 135.1933, 
    134.1971, 133.2151, 132.2472, 131.2934, 130.3535, 129.4275, 128.5152, 
    127.6164, 126.7311, 125.859, 125, 124.1539, 123.3204, 122.4994, 121.6906, 
    120.8939, 120.109, 119.3358,
  221.5041, 220.7353, 219.9545, 219.1612, 218.3553, 217.5364, 216.7044, 
    215.859, 215, 214.1271, 213.2402, 212.3389, 211.4232, 210.4929, 209.5477, 
    208.5876, 207.6124, 206.6219, 205.6162, 204.5951, 203.5586, 202.5068, 
    201.4395, 200.357, 199.2593, 198.1464, 197.0187, 195.8763, 194.7194, 
    193.5484, 192.3635, 191.1653, 189.954, 188.7303, 187.4946, 186.2475, 
    184.9897, 183.7218, 182.4444, 181.1585, 179.8647, 178.5639, 177.257, 
    175.9448, 174.6282, 173.3083, 171.986, 170.6622, 169.3378, 168.014, 
    166.6917, 165.3718, 164.0552, 162.743, 161.4361, 160.1353, 158.8415, 
    157.5556, 156.2782, 155.0103, 153.7525, 152.5054, 151.2697, 150.046, 
    148.8347, 147.6365, 146.4516, 145.2806, 144.1237, 142.9813, 141.8536, 
    140.7407, 139.643, 138.5605, 137.4932, 136.4414, 135.4049, 134.3838, 
    133.3781, 132.3876, 131.4124, 130.4523, 129.5071, 128.5768, 127.661, 
    126.7598, 125.8729, 125, 124.141, 123.2956, 122.4636, 121.6447, 120.8388, 
    120.0455, 119.2647, 118.4959,
  222.3516, 221.5882, 220.8121, 220.023, 219.2206, 218.4047, 217.575, 
    216.7311, 215.8729, 215, 214.1122, 213.2093, 212.291, 211.3571, 210.4073, 
    209.4416, 208.4597, 207.4614, 206.4467, 205.4155, 204.3676, 203.3031, 
    202.2219, 201.1241, 200.0097, 198.8788, 197.7316, 196.5683, 195.3892, 
    194.1945, 192.9845, 191.7598, 190.5207, 189.2677, 188.0015, 186.7226, 
    185.4317, 184.1296, 182.817, 181.4947, 180.1637, 178.8248, 177.479, 
    176.1273, 174.7708, 173.4105, 172.0474, 170.6826, 169.3174, 167.9526, 
    166.5895, 165.2292, 163.8727, 162.521, 161.1752, 159.8363, 158.5053, 
    157.183, 155.8704, 154.5683, 153.2774, 151.9985, 150.7323, 149.4793, 
    148.2402, 147.0155, 145.8055, 144.6108, 143.4317, 142.2684, 141.1212, 
    139.9903, 138.8759, 137.7781, 136.6969, 135.6324, 134.5845, 133.5533, 
    132.5386, 131.5403, 130.5584, 129.5927, 128.6429, 127.709, 126.7907, 
    125.8878, 125, 124.1271, 123.2689, 122.425, 121.5953, 120.7794, 119.977, 
    119.1879, 118.4118, 117.6484,
  223.207, 222.4496, 221.6789, 220.8948, 220.0968, 219.2846, 218.4579, 
    217.6164, 216.7598, 215.8878, 215, 214.0962, 213.1761, 212.2394, 
    211.2859, 210.3153, 209.3275, 208.3221, 207.2991, 206.2583, 205.1996, 
    204.1229, 203.0282, 201.9154, 200.7847, 199.6359, 198.4694, 197.2853, 
    196.0838, 194.8652, 193.6298, 192.3781, 191.1105, 189.8277, 188.53, 
    187.2183, 185.8933, 184.5558, 183.2065, 181.8465, 180.4766, 179.098, 
    177.7117, 176.3187, 174.9203, 173.5175, 172.1118, 170.7041, 169.2959, 
    167.8882, 166.4825, 165.0797, 163.6813, 162.2883, 160.902, 159.5234, 
    158.1535, 156.7935, 155.4442, 154.1067, 152.7817, 151.47, 150.1723, 
    148.8895, 147.6219, 146.3702, 145.1348, 143.9162, 142.7147, 141.5306, 
    140.3641, 139.2153, 138.0846, 136.9718, 135.8771, 134.8004, 133.7417, 
    132.7009, 131.6779, 130.6725, 129.6847, 128.7141, 127.7606, 126.8239, 
    125.9038, 125, 124.1122, 123.2402, 122.3836, 121.5421, 120.7154, 
    119.9032, 119.1052, 118.3211, 117.5504, 116.793,
  224.0701, 223.3195, 222.5551, 221.7767, 220.9838, 220.1762, 219.3535, 
    218.5152, 217.6611, 216.7907, 215.9038, 215, 214.079, 213.1404, 212.1839, 
    211.2094, 210.2164, 209.2047, 208.1741, 207.1245, 206.0556, 204.9673, 
    203.8596, 202.7323, 201.5855, 200.4192, 199.2335, 198.0286, 196.8046, 
    195.5619, 194.3008, 193.0217, 191.7251, 190.4115, 189.0817, 187.7362, 
    186.3759, 185.0016, 183.6143, 182.215, 180.8047, 179.3846, 177.9557, 
    176.5195, 175.0772, 173.63, 172.1794, 170.7267, 169.2733, 167.8206, 
    166.37, 164.9228, 163.4805, 162.0443, 160.6154, 159.1953, 157.785, 
    156.3857, 154.9984, 153.6241, 152.2638, 150.9183, 149.5885, 148.2749, 
    146.9783, 145.6992, 144.4381, 143.1954, 141.9714, 140.7665, 139.5808, 
    138.4145, 137.2677, 136.1404, 135.0327, 133.9444, 132.8755, 131.8259, 
    130.7953, 129.7836, 128.7906, 127.8161, 126.8596, 125.921, 125, 124.0962, 
    123.2093, 122.339, 121.4848, 120.6465, 119.8238, 119.0162, 118.2233, 
    117.4449, 116.6805, 115.9299,
  224.941, 224.1979, 223.4406, 222.6687, 221.8819, 221.0797, 220.2617, 
    219.4275, 218.5768, 217.709, 216.8239, 215.921, 215, 214.0604, 213.102, 
    212.1243, 211.127, 210.1099, 209.0726, 208.0148, 206.9365, 205.8373, 
    204.7171, 203.5758, 202.4134, 201.2298, 200.0252, 198.7996, 197.5532, 
    196.2863, 194.9991, 193.6922, 192.366, 191.0211, 189.6581, 188.2778, 
    186.8811, 185.4688, 184.0419, 182.6016, 181.1491, 179.6855, 178.2122, 
    176.7307, 175.2422, 173.7483, 172.2505, 170.7504, 169.2496, 167.7495, 
    166.2517, 164.7578, 163.2693, 161.7878, 160.3145, 158.8509, 157.3984, 
    155.9581, 154.5312, 153.1189, 151.7222, 150.3419, 148.9789, 147.634, 
    146.3078, 145.0009, 143.7137, 142.4468, 141.2004, 139.9748, 138.7702, 
    137.5866, 136.4242, 135.2829, 134.1627, 133.0635, 131.9852, 130.9274, 
    129.8901, 128.873, 127.8757, 126.898, 125.9396, 125, 124.079, 123.1761, 
    122.291, 121.4232, 120.5725, 119.7383, 118.9203, 118.1181, 117.3313, 
    116.5594, 115.8021, 115.059,
  225.8197, 225.0849, 224.3354, 223.5709, 222.7909, 221.995, 221.1827, 
    220.3535, 219.5071, 218.6429, 217.7606, 216.8596, 215.9396, 215, 
    214.0405, 213.0607, 212.0601, 211.0384, 209.9952, 208.9302, 207.8432, 
    206.7338, 205.6019, 204.4472, 203.2697, 202.0693, 200.846, 199.5999, 
    198.3312, 197.0399, 195.7266, 194.3915, 193.0351, 191.6581, 190.2611, 
    188.8449, 187.4105, 185.9587, 184.4907, 183.0078, 181.5111, 180.0021, 
    178.4822, 176.9529, 175.416, 173.8729, 172.3255, 170.7755, 169.2245, 
    167.6745, 166.1271, 164.584, 163.0471, 161.5178, 159.9979, 158.4889, 
    156.9922, 155.5093, 154.0413, 152.5895, 151.1551, 149.7389, 148.3419, 
    146.9649, 145.6085, 144.2734, 142.9601, 141.6688, 140.4001, 139.154, 
    137.9307, 136.7303, 135.5528, 134.3981, 133.2662, 132.1568, 131.0698, 
    130.0048, 128.9616, 127.9399, 126.9393, 125.9595, 125, 124.0604, 
    123.1404, 122.2394, 121.3571, 120.4929, 119.6465, 118.8173, 118.005, 
    117.2091, 116.4291, 115.6646, 114.9151, 114.1803,
  226.7061, 225.9804, 225.2396, 224.4833, 223.711, 222.9223, 222.1166, 
    221.2934, 220.4523, 219.5927, 218.7141, 217.8161, 216.898, 215.9595, 215, 
    214.019, 213.0162, 211.9909, 210.9429, 209.8716, 208.7768, 207.6581, 
    206.5151, 205.3478, 204.1558, 202.9391, 201.6976, 200.4313, 199.1402, 
    197.8247, 196.4849, 195.1213, 193.7343, 192.3245, 190.8926, 189.4395, 
    187.966, 186.4733, 184.9626, 183.4351, 181.8922, 180.3356, 178.7667, 
    177.1874, 175.5993, 174.0044, 172.4046, 170.8019, 169.1981, 167.5954, 
    165.9956, 164.4007, 162.8126, 161.2333, 159.6644, 158.1078, 156.5649, 
    155.0374, 153.5267, 152.034, 150.5605, 149.1074, 147.6755, 146.2657, 
    144.8787, 143.5151, 142.1753, 140.8598, 139.5687, 138.3024, 137.0609, 
    135.8442, 134.6522, 133.4849, 132.3419, 131.2232, 130.1284, 129.0571, 
    128.0091, 126.9838, 125.981, 125, 124.0405, 123.102, 122.1839, 121.2859, 
    120.4073, 119.5477, 118.7066, 117.8834, 117.0777, 116.289, 115.5167, 
    114.7604, 114.0196, 113.2939,
  227.6002, 226.8844, 226.1531, 225.4059, 224.6422, 223.8616, 223.0634, 
    222.2472, 221.4124, 220.5584, 219.6847, 218.7906, 217.8757, 216.9393, 
    215.981, 215, 213.9959, 212.9682, 211.9164, 210.8398, 209.7382, 208.6111, 
    207.4581, 206.2789, 205.0732, 203.8407, 202.5815, 201.2953, 199.9823, 
    198.6425, 197.2762, 195.8838, 194.4657, 193.0224, 191.5547, 190.0636, 
    188.5498, 187.0146, 185.4594, 183.8854, 182.2942, 180.6875, 179.0672, 
    177.435, 175.7931, 174.1435, 172.4883, 170.8298, 169.1702, 167.5117, 
    165.8565, 164.2069, 162.565, 160.9328, 159.3125, 157.7058, 156.1146, 
    154.5406, 152.9854, 151.4502, 149.9364, 148.4453, 146.9776, 145.5343, 
    144.1162, 142.7238, 141.3575, 140.0177, 138.7047, 137.4185, 136.1593, 
    134.9268, 133.7211, 132.5419, 131.3889, 130.2618, 129.1602, 128.0836, 
    127.0318, 126.0041, 125, 124.019, 123.0607, 122.1243, 121.2094, 120.3153, 
    119.4416, 118.5876, 117.7528, 116.9366, 116.1384, 115.3578, 114.5941, 
    113.8469, 113.1156, 112.3998,
  228.502, 227.7968, 227.0759, 226.3386, 225.5845, 224.8129, 224.0233, 
    223.2151, 222.3876, 221.5403, 220.6725, 219.7836, 218.873, 217.9399, 
    216.9838, 216.0041, 215, 213.971, 212.9165, 211.8359, 210.7286, 209.5941, 
    208.432, 207.2418, 206.0232, 204.7758, 203.4994, 202.1939, 200.8592, 
    199.4954, 198.1026, 196.6812, 195.2315, 193.7542, 192.2498, 190.7195, 
    189.1641, 187.5849, 185.9832, 184.3606, 182.7188, 181.0596, 179.385, 
    177.6972, 175.9983, 174.2908, 172.577, 170.8594, 169.1406, 167.423, 
    165.7092, 164.0017, 162.3028, 160.615, 158.9404, 157.2812, 155.6394, 
    154.0168, 152.4151, 150.8359, 149.2805, 147.7502, 146.2458, 144.7685, 
    143.3188, 141.8974, 140.5046, 139.1408, 137.8061, 136.5006, 135.2242, 
    133.9768, 132.7582, 131.568, 130.4059, 129.2714, 128.1641, 127.0835, 
    126.029, 125, 123.9959, 123.0162, 122.0601, 121.127, 120.2164, 119.3275, 
    118.4597, 117.6124, 116.7849, 115.9767, 115.1871, 114.4155, 113.6614, 
    112.9241, 112.2032, 111.498,
  229.4114, 228.7177, 228.008, 227.2816, 226.5379, 225.7764, 224.9963, 
    224.1971, 223.3781, 222.5386, 221.6779, 220.7953, 219.8901, 218.9616, 
    218.0091, 217.0318, 216.029, 215, 213.9441, 212.8606, 211.7489, 210.6083, 
    209.4382, 208.2381, 207.0076, 205.7461, 204.4533, 203.1291, 201.7732, 
    200.3856, 198.9664, 197.5159, 196.0343, 194.5223, 192.9805, 191.4098, 
    189.8114, 188.1864, 186.5364, 184.863, 183.1681, 181.4536, 179.7219, 
    177.9752, 176.216, 174.4471, 172.6711, 170.8909, 169.1091, 167.3289, 
    165.5529, 163.784, 162.0248, 160.2781, 158.5464, 156.8319, 155.137, 
    153.4636, 151.8136, 150.1886, 148.5902, 147.0195, 145.4777, 143.9657, 
    142.4841, 141.0336, 139.6144, 138.2268, 136.8709, 135.5467, 134.2539, 
    132.9924, 131.7619, 130.5618, 129.3917, 128.2511, 127.1394, 126.0559, 
    125, 123.971, 122.9682, 121.9909, 121.0384, 120.1099, 119.2047, 118.3221, 
    117.4614, 116.6219, 115.8029, 115.0037, 114.2237, 113.4621, 112.7184, 
    111.992, 111.2822, 110.5886,
  230.3284, 229.647, 228.9493, 228.2346, 227.5023, 226.7518, 225.9824, 
    225.1933, 224.3838, 223.5533, 222.7009, 221.8259, 220.9274, 220.0048, 
    219.0571, 218.0836, 217.0835, 216.0559, 215, 213.915, 212.8002, 211.6547, 
    210.478, 209.2692, 208.0278, 206.7533, 205.4451, 204.1029, 202.7264, 
    201.3154, 199.8701, 198.3904, 196.8767, 195.3295, 193.7494, 192.1374, 
    190.4945, 188.8221, 187.1217, 185.3952, 183.6444, 181.8718, 180.0796, 
    178.2706, 176.4475, 174.6134, 172.7713, 170.9243, 169.0757, 167.2287, 
    165.3866, 163.5525, 161.7294, 159.9204, 158.1282, 156.3556, 154.6048, 
    152.8783, 151.1779, 149.5055, 147.8626, 146.2506, 144.6705, 143.1233, 
    141.6096, 140.1299, 138.6846, 137.2736, 135.8971, 134.5549, 133.2467, 
    131.9722, 130.7308, 129.522, 128.3453, 127.1998, 126.085, 125, 123.9441, 
    122.9165, 121.9163, 120.9429, 119.9952, 119.0726, 118.1741, 117.2991, 
    116.4467, 115.6162, 114.8067, 114.0176, 113.2482, 112.4977, 111.7654, 
    111.0507, 110.353, 109.6716,
  231.2529, 230.5846, 229.8998, 229.1978, 228.4779, 227.7393, 226.9815, 
    226.2036, 225.4049, 224.5845, 223.7417, 222.8755, 221.9852, 221.0698, 
    220.1284, 219.1602, 218.1641, 217.1394, 216.085, 215, 213.8835, 212.7347, 
    211.5527, 210.3366, 209.0856, 207.7992, 206.4767, 205.1174, 203.7211, 
    202.2875, 200.8163, 199.3076, 197.7617, 196.1788, 194.5597, 192.9053, 
    191.2165, 189.4949, 187.742, 185.9598, 184.1504, 182.3164, 180.4603, 
    178.5852, 176.6942, 174.7907, 172.8781, 170.96, 169.04, 167.1219, 
    165.2093, 163.3058, 161.4148, 159.5397, 157.6836, 155.8496, 154.0402, 
    152.258, 150.5051, 148.7835, 147.0947, 145.4403, 143.8212, 142.2383, 
    140.6924, 139.1837, 137.7125, 136.2789, 134.8826, 133.5233, 132.2008, 
    130.9144, 129.6634, 128.4473, 127.2653, 126.1165, 125, 123.915, 122.8606, 
    121.8359, 120.8398, 119.8716, 118.9302, 118.0148, 117.1245, 116.2583, 
    115.4155, 114.5951, 113.7964, 113.0185, 112.2607, 111.5221, 110.8022, 
    110.1002, 109.4154, 108.7472,
  232.1847, 231.5304, 230.8594, 230.1709, 229.4643, 228.7389, 227.9938, 
    227.2282, 226.4414, 225.6324, 224.8004, 223.9444, 223.0635, 222.1568, 
    221.2232, 220.2618, 219.2714, 218.2511, 217.1998, 216.1165, 215, 
    213.8494, 212.6637, 211.4417, 210.1828, 208.8859, 207.5502, 206.1751, 
    204.76, 203.3043, 201.8079, 200.2705, 198.6923, 197.0736, 195.4148, 
    193.7169, 191.9809, 190.2082, 188.4006, 186.5601, 184.689, 182.7901, 
    180.8664, 178.9211, 176.9578, 174.9802, 172.9923, 170.9981, 169.0019, 
    167.0077, 165.0198, 163.0422, 161.0789, 159.1336, 157.2099, 155.311, 
    153.4399, 151.5994, 149.7918, 148.0191, 146.2831, 144.5852, 142.9264, 
    141.3077, 139.7295, 138.1921, 136.6957, 135.24, 133.8249, 132.4498, 
    131.1141, 129.8172, 128.5583, 127.3364, 126.1506, 125, 123.8835, 
    122.8002, 121.7489, 120.7286, 119.7382, 118.7768, 117.8432, 116.9365, 
    116.0556, 115.1996, 114.3676, 113.5586, 112.7718, 112.0062, 111.2611, 
    110.5357, 109.8291, 109.1406, 108.4696, 107.8153,
  233.1238, 232.4843, 231.8279, 231.154, 230.4617, 229.7503, 229.019, 
    228.267, 227.4932, 226.6969, 225.8771, 225.0327, 224.1627, 223.2662, 
    222.3419, 221.3889, 220.4059, 219.3917, 218.3453, 217.2653, 216.1506, 
    215, 213.8123, 212.5863, 211.321, 210.0152, 208.6679, 207.2783, 205.8455, 
    204.3689, 202.8479, 201.2824, 199.6721, 198.0173, 196.3184, 194.576, 
    192.7914, 190.9658, 189.1012, 187.1996, 185.2636, 183.2962, 181.3006, 
    179.2806, 177.2401, 175.1833, 173.1147, 171.039, 168.961, 166.8853, 
    164.8167, 162.7599, 160.7194, 158.6994, 156.7038, 154.7364, 152.8004, 
    150.8988, 149.0342, 147.2086, 145.424, 143.6816, 141.9827, 140.3279, 
    138.7176, 137.1521, 135.6311, 134.1545, 132.7217, 131.3321, 129.9848, 
    128.679, 127.4137, 126.1877, 125, 123.8494, 122.7347, 121.6547, 120.6083, 
    119.5941, 118.6111, 117.6581, 116.7338, 115.8373, 114.9673, 114.1229, 
    113.3031, 112.5068, 111.733, 110.981, 110.2497, 109.5383, 108.846, 
    108.1721, 107.5157, 106.8762,
  234.0701, 233.4462, 232.8053, 232.1469, 231.4699, 230.7736, 230.0573, 
    229.3198, 228.5605, 227.7781, 226.9718, 226.1404, 225.2829, 224.3981, 
    223.4849, 222.5419, 221.568, 220.5618, 219.522, 218.4473, 217.3363, 
    216.1877, 215, 213.7719, 212.502, 211.1892, 209.832, 208.4295, 206.9805, 
    205.4841, 203.9397, 202.3467, 200.7048, 199.0139, 197.2744, 195.4869, 
    193.6523, 191.772, 189.8479, 187.8823, 185.8779, 183.8379, 181.766, 
    179.6663, 177.5432, 175.4015, 173.2463, 171.083, 168.917, 166.7537, 
    164.5985, 162.4568, 160.3337, 158.234, 156.1621, 154.1221, 152.1177, 
    150.1521, 148.228, 146.3477, 144.5131, 142.7256, 140.9861, 139.2952, 
    137.6533, 136.0603, 134.5159, 133.0195, 131.5705, 130.168, 128.8108, 
    127.498, 126.2281, 125, 123.8123, 122.6636, 121.5527, 120.478, 119.4382, 
    118.432, 117.4581, 116.5151, 115.6019, 114.7171, 113.8596, 113.0282, 
    112.2219, 111.4395, 110.6802, 109.9427, 109.2264, 108.5301, 107.8532, 
    107.1946, 106.5538, 105.9299,
  235.0234, 234.416, 233.7915, 233.1494, 232.4887, 231.8087, 231.1084, 
    230.3868, 229.643, 228.8759, 228.0846, 227.2677, 226.4242, 225.5528, 
    224.6522, 223.7211, 222.7582, 221.7619, 220.7308, 219.6634, 218.5583, 
    217.4137, 216.2281, 215, 213.7278, 212.4099, 211.0449, 209.6313, 
    208.1678, 206.6533, 205.0867, 203.4673, 201.7944, 200.0677, 198.2875, 
    196.454, 194.5683, 192.6315, 190.6456, 188.6129, 186.5363, 184.4195, 
    182.2663, 180.0813, 177.8696, 175.6366, 173.3882, 171.1305, 168.8695, 
    166.6118, 164.3634, 162.1304, 159.9187, 157.7337, 155.5805, 153.4637, 
    151.3871, 149.3544, 147.3685, 145.4317, 143.546, 141.7125, 139.9323, 
    138.2056, 136.5327, 134.9133, 133.3467, 131.8322, 130.3687, 128.9551, 
    127.5901, 126.2722, 125, 123.7719, 122.5863, 121.4417, 120.3366, 
    119.2692, 118.2381, 117.2418, 116.2789, 115.3478, 114.4472, 113.5758, 
    112.7323, 111.9154, 111.1241, 110.357, 109.6132, 108.8917, 108.1913, 
    107.5113, 106.8506, 106.2085, 105.584, 104.9766,
  235.9837, 235.3935, 234.7863, 234.1615, 233.5181, 232.8553, 232.1722, 
    231.4676, 230.7407, 229.9903, 229.2153, 228.4145, 227.5866, 226.7303, 
    225.8442, 224.9268, 223.9768, 222.9924, 221.9722, 220.9144, 219.8172, 
    218.679, 217.498, 216.2722, 215, 213.6795, 212.3089, 210.8864, 209.4106, 
    207.8797, 206.2926, 204.6481, 202.9452, 201.1834, 199.3625, 197.4827, 
    195.5447, 193.5496, 191.4994, 189.3965, 187.2439, 185.0454, 182.8055, 
    180.5292, 178.2223, 175.8909, 173.5418, 171.1818, 168.8182, 166.4582, 
    164.1091, 161.7777, 159.4708, 157.1945, 154.9546, 152.7561, 150.6035, 
    148.5006, 146.4504, 144.4553, 142.5173, 140.6375, 138.8166, 137.0548, 
    135.3519, 133.7074, 132.1203, 130.5894, 129.1136, 127.6912, 126.3205, 
    125, 123.7278, 122.502, 121.321, 120.1828, 119.0856, 118.0278, 117.0076, 
    116.0232, 115.0732, 114.1558, 113.2697, 112.4134, 111.5855, 110.7847, 
    110.0097, 109.2593, 108.5324, 107.8278, 107.1447, 106.4819, 105.8385, 
    105.2137, 104.6065, 104.0163,
  236.9507, 236.3785, 235.7896, 235.183, 234.5579, 233.9134, 233.2485, 
    232.5623, 231.8536, 231.1212, 230.3641, 229.5808, 228.7702, 227.9307, 
    227.0609, 226.1593, 225.2242, 224.2539, 223.2467, 222.2008, 221.1141, 
    219.9848, 218.8108, 217.5901, 216.3205, 215, 213.6264, 212.1977, 
    210.7119, 209.167, 207.5614, 205.8935, 204.162, 202.366, 200.5049, 
    198.5785, 196.5874, 194.5325, 192.4155, 190.239, 188.0061, 185.721, 
    183.3885, 181.0142, 178.6046, 176.1668, 173.7085, 171.2375, 168.7625, 
    166.2915, 163.8332, 161.3954, 158.9858, 156.6115, 154.279, 151.9939, 
    149.761, 147.5845, 145.4675, 143.4126, 141.4215, 139.4951, 137.634, 
    135.838, 134.1065, 132.4386, 130.833, 129.2881, 127.8023, 126.3736, 125, 
    123.6795, 122.4099, 121.1892, 120.0152, 118.8859, 117.7992, 116.7533, 
    115.7461, 114.7758, 113.8407, 112.9391, 112.0693, 111.2298, 110.4192, 
    109.6359, 108.8788, 108.1464, 107.4377, 106.7515, 106.0866, 105.4421, 
    104.817, 104.2104, 103.6215, 103.0493,
  237.9244, 237.371, 236.8011, 236.2136, 235.6078, 234.9827, 234.3373, 
    233.6705, 232.9813, 232.2684, 231.5306, 230.7665, 229.9748, 229.154, 
    228.3024, 227.4185, 226.5006, 225.5467, 224.5549, 223.5233, 222.4498, 
    221.3321, 220.168, 218.9551, 217.6911, 216.3736, 215, 213.5679, 212.075, 
    210.5188, 208.8972, 207.2082, 205.4499, 203.6211, 201.7205, 199.7478, 
    197.703, 195.5868, 193.4008, 191.1474, 188.8298, 186.4526, 184.0209, 
    181.5412, 179.0206, 176.4673, 173.8901, 171.2983, 168.7017, 166.1099, 
    163.5327, 160.9794, 158.4588, 155.9791, 153.5474, 151.1702, 148.8526, 
    146.5992, 144.4132, 142.297, 140.2522, 138.2795, 136.3789, 134.5501, 
    132.7918, 131.1028, 129.4812, 127.925, 126.4321, 125, 123.6264, 122.3088, 
    121.0449, 119.832, 118.6679, 117.5502, 116.4767, 115.4451, 114.4533, 
    113.4994, 112.5815, 111.6976, 110.846, 110.0252, 109.2335, 108.4694, 
    107.7316, 107.0187, 106.3295, 105.6627, 105.0173, 104.3922, 103.7864, 
    103.1989, 102.629, 102.0756,
  238.9044, 238.3707, 237.8206, 237.2533, 236.6677, 236.063, 235.4382, 
    234.7922, 234.1237, 233.4317, 232.7147, 231.9714, 231.2004, 230.4001, 
    229.5687, 228.7047, 227.8061, 226.8709, 225.8971, 224.8826, 223.8249, 
    222.7217, 221.5705, 220.3687, 219.1136, 217.8023, 216.4321, 215, 
    213.5032, 211.9389, 210.3043, 208.5969, 206.8143, 204.9546, 203.016, 
    200.9976, 198.8989, 196.7203, 194.463, 192.1293, 189.7226, 187.2474, 
    184.7095, 182.116, 179.475, 176.796, 174.0889, 171.3649, 168.6351, 
    165.9111, 163.204, 160.525, 157.884, 155.2905, 152.7526, 150.2774, 
    147.8707, 145.537, 143.2797, 141.1011, 139.0024, 136.984, 135.0454, 
    133.1857, 131.4031, 129.6957, 128.0611, 126.4968, 125, 123.5679, 
    122.1977, 120.8864, 119.6313, 118.4295, 117.2783, 116.1751, 115.1174, 
    114.1029, 113.1291, 112.1939, 111.2953, 110.4313, 109.5999, 108.7996, 
    108.0286, 107.2853, 106.5683, 105.8763, 105.2078, 104.5618, 103.937, 
    103.3323, 102.7467, 102.1794, 101.6293, 101.0956,
  239.8907, 239.3774, 238.848, 238.3016, 237.7373, 237.1542, 236.5511, 
    235.9269, 235.2806, 234.6108, 233.9162, 233.1954, 232.4468, 231.6688, 
    230.8598, 230.0177, 229.1408, 228.2268, 227.2736, 226.2789, 225.24, 
    224.1545, 223.0195, 221.8322, 220.5894, 219.2881, 217.925, 216.4968, 215, 
    213.4313, 211.7874, 210.065, 208.2611, 206.373, 204.3985, 202.3356, 
    200.1834, 197.9417, 195.6112, 193.194, 190.6933, 188.1138, 185.4619, 
    182.7454, 179.9735, 177.157, 174.3076, 171.4381, 168.5619, 165.6924, 
    162.843, 160.0265, 157.2546, 154.5381, 151.8862, 149.3067, 146.806, 
    144.3888, 142.0583, 139.8166, 137.6644, 135.6015, 133.627, 131.7389, 
    129.935, 128.2126, 126.5687, 125, 123.5032, 122.075, 120.7119, 119.4106, 
    118.1678, 116.9805, 115.8455, 114.76, 113.7211, 112.7264, 111.7732, 
    110.8592, 109.9823, 109.1402, 108.3312, 107.5532, 106.8046, 106.0838, 
    105.3892, 104.7194, 104.0731, 103.4489, 102.8458, 102.2627, 101.6984, 
    101.152, 100.6226, 100.1093,
  240.883, 240.3909, 239.883, 239.3585, 238.8164, 238.2558, 237.6755, 
    237.0745, 236.4516, 235.8055, 235.1348, 234.4381, 233.7137, 232.9601, 
    232.1753, 231.3575, 230.5046, 229.6144, 228.6846, 227.7125, 226.6957, 
    225.6311, 224.5159, 223.3467, 222.1203, 220.833, 219.4812, 218.0611, 
    216.5687, 215, 213.351, 211.6178, 209.7964, 207.8834, 205.8756, 203.7704, 
    201.5657, 199.2607, 196.8556, 194.3517, 191.7523, 189.062, 186.2876, 
    183.4378, 180.5229, 177.5555, 174.5491, 171.5191, 168.4809, 165.4509, 
    162.4445, 159.4771, 156.5622, 153.7124, 150.938, 148.2477, 145.6483, 
    143.1444, 140.7393, 138.4343, 136.2296, 134.1244, 132.1166, 130.2036, 
    128.3822, 126.649, 125, 123.4313, 121.9389, 120.5188, 119.167, 117.8797, 
    116.6533, 115.4841, 114.3689, 113.3043, 112.2875, 111.3155, 110.3856, 
    109.4954, 108.6425, 107.8247, 107.0399, 106.2863, 105.5619, 104.8652, 
    104.1945, 103.5484, 102.9255, 102.3245, 101.7442, 101.1836, 100.6415, 
    100.117, 99.60909, 99.117,
  241.8811, 241.411, 240.9254, 240.4236, 239.9047, 239.3676, 238.8113, 
    238.2346, 237.6365, 237.0155, 236.3702, 235.6992, 235.0009, 234.2734, 
    233.5151, 232.7238, 231.8974, 231.0336, 230.1299, 229.1837, 228.1921, 
    227.1521, 226.0603, 224.9133, 223.7074, 222.4386, 221.1028, 219.6957, 
    218.2126, 216.649, 215, 213.2608, 211.4268, 209.4932, 207.4559, 205.3113, 
    203.0562, 200.6886, 198.2079, 195.6148, 192.9118, 190.1038, 187.1977, 
    184.203, 181.1316, 177.9977, 174.8176, 171.6091, 168.3909, 165.1824, 
    162.0023, 158.8684, 155.797, 152.8023, 149.8962, 147.0882, 144.3852, 
    141.7921, 139.3114, 136.9438, 134.6887, 132.5441, 130.5068, 128.5732, 
    126.7392, 125, 123.351, 121.7874, 120.3043, 118.8972, 117.5614, 116.2926, 
    115.0867, 113.9397, 112.8479, 111.8079, 110.8163, 109.8701, 108.9664, 
    108.1026, 107.2762, 106.4849, 105.7266, 104.9991, 104.3008, 103.6298, 
    102.9845, 102.3635, 101.7654, 101.1887, 100.6324, 100.0953, 99.57638, 
    99.07459, 98.58904, 98.11887,
  242.8848, 242.4373, 241.9749, 241.4967, 241.0018, 240.4892, 239.958, 
    239.4069, 238.8347, 238.2402, 237.6219, 236.9783, 236.3078, 235.6085, 
    234.8787, 234.1162, 233.3188, 232.4841, 231.6096, 230.6924, 229.7295, 
    228.7176, 227.6533, 226.5327, 225.3519, 224.1065, 222.7918, 221.4031, 
    219.935, 218.3822, 216.7392, 215, 213.159, 211.2103, 209.1486, 206.9686, 
    204.6662, 202.2379, 199.6816, 196.9971, 194.1863, 191.2534, 188.2056, 
    185.0533, 181.8097, 178.4915, 175.1178, 171.7098, 168.2902, 164.8822, 
    161.5085, 158.1903, 154.9467, 151.7944, 148.7466, 145.8137, 143.0029, 
    140.3184, 137.7621, 135.3338, 133.0314, 130.8514, 128.7897, 126.841, 125, 
    123.2608, 121.6178, 120.065, 118.5969, 117.2082, 115.8935, 114.6481, 
    113.4673, 112.3467, 111.2824, 110.2705, 109.3076, 108.3904, 107.5158, 
    106.6812, 105.8838, 105.1213, 104.3915, 103.6922, 103.0217, 102.3781, 
    101.7598, 101.1653, 100.5931, 100.042, 99.51077, 98.99823, 98.50335, 
    98.02514, 97.56269, 97.11515,
  243.8939, 243.4697, 243.0311, 242.5773, 242.1074, 241.6204, 241.1152, 
    240.5908, 240.046, 239.4793, 238.8895, 238.2749, 237.634, 236.9649, 
    236.2657, 235.5343, 234.7685, 233.9657, 233.1233, 232.2383, 231.3077, 
    230.3279, 229.2952, 228.2056, 227.0548, 225.838, 224.5501, 223.1857, 
    221.7389, 220.2036, 218.5732, 216.841, 215, 213.043, 210.9632, 208.7537, 
    206.4086, 203.9227, 201.2922, 198.5153, 195.5927, 192.5277, 189.3277, 
    186.0034, 182.57, 179.0465, 175.4557, 171.8233, 168.1767, 164.5443, 
    160.9535, 157.43, 153.9966, 150.6723, 147.4723, 144.4073, 141.4847, 
    138.7078, 136.0773, 133.5914, 131.2463, 129.0368, 126.957, 125, 123.159, 
    121.4268, 119.7964, 118.2611, 116.8143, 115.4499, 114.162, 112.9452, 
    111.7944, 110.7048, 109.6721, 108.6923, 107.7617, 106.8767, 106.0343, 
    105.2315, 104.4657, 103.7343, 103.0351, 102.366, 101.7251, 101.1105, 
    100.5207, 99.95405, 99.40917, 98.88477, 98.37963, 97.89262, 97.4227, 
    96.96889, 96.5303, 96.10609,
  244.9081, 244.5078, 244.0938, 243.6652, 243.2211, 242.7606, 242.2826, 
    241.786, 241.2697, 240.7323, 240.1723, 239.5885, 238.9789, 238.3419, 
    237.6755, 236.9776, 236.2458, 235.4777, 234.6705, 233.8212, 232.9264, 
    231.9827, 230.9861, 229.9323, 228.8166, 227.634, 226.3789, 225.0454, 
    223.627, 222.1166, 220.5068, 218.7897, 216.957, 215, 212.9101, 210.6786, 
    208.2973, 205.7589, 203.0573, 200.1884, 197.1511, 193.9474, 190.5838, 
    187.0719, 183.4281, 179.6749, 175.8391, 171.9522, 168.0478, 164.1609, 
    160.3251, 156.5719, 152.9281, 149.4162, 146.0526, 142.8489, 139.8116, 
    136.9427, 134.2411, 131.7027, 129.3214, 127.0899, 125, 123.043, 121.2103, 
    119.4932, 117.8834, 116.373, 114.9546, 113.6211, 112.366, 111.1834, 
    110.0677, 109.0139, 108.0173, 107.0736, 106.1788, 105.3295, 104.5223, 
    103.7541, 103.0224, 102.3245, 101.6581, 101.0211, 100.4115, 99.82764, 
    99.26775, 98.73032, 98.21397, 97.71739, 97.2394, 96.77886, 96.33477, 
    95.90617, 95.49216, 95.09195,
  245.927, 245.5514, 245.1627, 244.7601, 244.3427, 243.9095, 243.4597, 
    242.992, 242.5054, 241.9985, 241.47, 240.9183, 240.3419, 239.7389, 
    239.1074, 238.4453, 237.7502, 237.0195, 236.2506, 235.4403, 234.5852, 
    233.6816, 232.7256, 231.7125, 230.6375, 229.4951, 228.2795, 226.984, 
    225.6015, 224.1244, 222.5441, 220.8514, 219.0368, 217.0899, 215, 
    212.7562, 210.3477, 207.7643, 204.997, 202.0387, 198.8855, 195.5371, 
    191.9988, 188.2818, 184.4044, 180.3923, 176.278, 172.0999, 167.9001, 
    163.722, 159.6077, 155.5956, 151.7182, 148.0012, 144.4629, 141.1145, 
    137.9613, 135.003, 132.2357, 129.6523, 127.2438, 125, 122.9101, 120.9632, 
    119.1486, 117.4559, 115.8756, 114.3984, 113.016, 111.7205, 110.5049, 
    109.3625, 108.2875, 107.2744, 106.3184, 105.4148, 104.5597, 103.7494, 
    102.9805, 102.2498, 101.5547, 100.8926, 100.2611, 99.65811, 99.08168, 
    98.53003, 98.00151, 97.49463, 97.008, 96.54034, 96.09048, 95.65735, 
    95.23992, 94.83728, 94.44856, 94.07298,
  246.9505, 246.6002, 246.2374, 245.8615, 245.4715, 245.0666, 244.6459, 
    244.2082, 243.7525, 243.2774, 242.7817, 242.2638, 241.7222, 241.1551, 
    240.5605, 239.9364, 239.2805, 238.5902, 237.8626, 237.0947, 236.2831, 
    235.424, 234.5131, 233.546, 232.5173, 231.4215, 230.2522, 229.0024, 
    227.6644, 226.2296, 224.6887, 223.0314, 221.2463, 219.3214, 217.2438, 
    215, 212.5761, 209.9584, 207.1341, 204.0921, 200.8243, 197.3271, 193.603, 
    189.6623, 185.5245, 181.2192, 176.7855, 172.271, 167.729, 163.2145, 
    158.7808, 154.4755, 150.3377, 146.397, 142.6729, 139.1757, 135.9079, 
    132.8659, 130.0416, 127.4239, 125, 122.7562, 120.6786, 118.7537, 
    116.9687, 115.3113, 113.7703, 112.3356, 110.9976, 109.7478, 108.5785, 
    107.4827, 106.454, 105.4869, 104.576, 103.7169, 102.9053, 102.1374, 
    101.4098, 100.7195, 100.0635, 99.43947, 98.84492, 98.27782, 97.73621, 
    97.21835, 96.72261, 96.24755, 95.79179, 95.35411, 94.93336, 94.52849, 
    94.13853, 93.76257, 93.3998, 93.04945,
  247.9783, 247.6538, 247.3176, 246.969, 246.6073, 246.2315, 245.8408, 
    245.4341, 245.0103, 244.5683, 244.1067, 243.6241, 243.1189, 242.5895, 
    242.034, 241.4502, 240.8359, 240.1886, 239.5055, 238.7835, 238.0191, 
    237.2086, 236.3477, 235.4317, 234.4553, 233.4126, 232.297, 231.1011, 
    229.8166, 228.4343, 226.9438, 225.3338, 223.5914, 221.7027, 219.6523, 
    217.4239, 215, 212.3627, 209.4944, 206.3785, 203.0015, 199.3542, 
    195.4348, 191.2509, 186.8223, 182.1825, 177.379, 172.4715, 167.5285, 
    162.621, 157.8175, 153.1777, 148.7491, 144.5652, 140.6458, 136.9985, 
    133.6215, 130.5056, 127.6373, 125, 122.5761, 120.3477, 118.2973, 
    116.4086, 114.6662, 113.0562, 111.5657, 110.1834, 108.8989, 107.703, 
    106.5874, 105.5447, 104.5683, 103.6523, 102.7914, 101.9809, 101.2165, 
    100.4945, 99.81139, 99.16409, 98.5498, 97.96602, 97.41046, 96.88105, 
    96.37591, 95.89333, 95.43173, 94.9897, 94.56594, 94.15924, 93.7685, 
    93.39273, 93.03098, 92.6824, 92.34621, 92.02168,
  249.0101, 248.7119, 248.4028, 248.0823, 247.7495, 247.4036, 247.0437, 
    246.669, 246.2782, 245.8704, 245.4442, 244.9984, 244.5312, 244.0413, 
    243.5267, 242.9854, 242.4151, 241.8136, 241.1779, 240.5051, 239.7918, 
    239.0342, 238.228, 237.3685, 236.4504, 235.4675, 234.4132, 233.2797, 
    232.0583, 230.7393, 229.3114, 227.7621, 226.0773, 224.2411, 222.2357, 
    220.0416, 217.6373, 215, 212.1061, 208.9323, 205.457, 201.6635, 197.5423, 
    193.096, 188.3424, 183.3188, 178.0826, 172.7099, 167.2901, 161.9174, 
    156.6812, 151.6576, 146.904, 142.4577, 138.3365, 134.543, 131.0677, 
    127.8939, 125, 122.3627, 119.9584, 117.7643, 115.7589, 113.9227, 
    112.2379, 110.6886, 109.2607, 107.9417, 106.7203, 105.5868, 104.5325, 
    103.5496, 102.6315, 101.772, 100.9658, 100.2082, 99.4949, 98.82211, 
    98.18644, 97.58487, 97.01465, 96.47334, 95.9587, 95.46874, 95.00165, 
    94.55576, 94.12959, 93.72176, 93.33103, 92.95627, 92.59641, 92.25053, 
    91.91771, 91.59716, 91.28813, 90.98993,
  250.0455, 249.7741, 249.4928, 249.2009, 248.8976, 248.5824, 248.2542, 
    247.9123, 247.5556, 247.183, 246.7935, 246.3857, 245.9581, 245.5093, 
    245.0374, 244.5406, 244.0168, 243.4636, 242.8783, 242.258, 241.5994, 
    240.8988, 240.1521, 239.3544, 238.5006, 237.5845, 236.5992, 235.537, 
    234.3888, 233.1444, 231.7921, 230.3184, 228.7078, 226.9427, 225.003, 
    222.8659, 220.5056, 217.8939, 215, 211.7919, 208.238, 204.3098, 199.9866, 
    195.2609, 190.1452, 184.6786, 178.93, 172.9979, 167.0021, 161.07, 
    155.3214, 149.8548, 144.7391, 140.0134, 135.6902, 131.762, 128.2081, 125, 
    122.1061, 119.4944, 117.1341, 114.997, 113.0573, 111.2922, 109.6816, 
    108.2079, 106.8556, 105.6112, 104.463, 103.4008, 102.4155, 101.4994, 
    100.6456, 99.84793, 99.10118, 98.4006, 97.74202, 97.12173, 96.53644, 
    95.98319, 95.45937, 94.96259, 94.49074, 94.0419, 93.61434, 93.2065, 
    92.81697, 92.44444, 92.08774, 91.7458, 91.41763, 91.10236, 90.79913, 
    90.50721, 90.2259, 89.95454,
  251.0842, 250.8401, 250.587, 250.3243, 250.0513, 249.7673, 249.4716, 
    249.1633, 248.8415, 248.5053, 248.1535, 247.785, 247.3984, 246.9922, 
    246.5649, 246.1146, 245.6394, 245.137, 244.6048, 244.0402, 243.4399, 
    242.8004, 242.1177, 241.3871, 240.6035, 239.761, 238.8526, 237.8707, 
    236.806, 235.6483, 234.3852, 233.0029, 231.4847, 229.8116, 227.9613, 
    225.9079, 223.6215, 221.0677, 218.2081, 215, 211.3986, 207.3597, 
    202.8449, 197.8296, 192.3137, 186.3334, 179.9703, 173.3532, 166.6468, 
    160.0297, 153.6666, 147.6863, 142.1704, 137.1551, 132.6403, 128.6014, 
    125, 121.7919, 118.9323, 116.3785, 114.0921, 112.0387, 110.1884, 
    108.5153, 106.9972, 105.6148, 104.3517, 103.194, 102.1293, 101.1473, 
    100.239, 99.39646, 98.61288, 97.88232, 97.19958, 96.56008, 95.95979, 
    95.39516, 94.86303, 94.3606, 93.88536, 93.43508, 93.00777, 92.60162, 
    92.215, 91.84647, 91.49471, 91.15849, 90.83672, 90.52844, 90.23272, 
    89.94873, 89.67571, 89.41297, 89.15987, 88.91582,
  252.1259, 251.9096, 251.6852, 251.4521, 251.2098, 250.9578, 250.6952, 
    250.4213, 250.1353, 249.8363, 249.5234, 249.1953, 248.8509, 248.4889, 
    248.1078, 247.7058, 247.2812, 246.8319, 246.3556, 245.8496, 245.311, 
    244.7364, 244.1221, 243.4637, 242.7561, 241.9939, 241.1702, 240.2774, 
    239.3067, 238.2477, 237.0882, 235.8137, 234.4073, 232.8489, 231.1145, 
    229.1757, 226.9985, 224.543, 221.762, 218.6014, 215, 210.8925, 206.2148, 
    200.9138, 194.9639, 188.3878, 181.2773, 173.8024, 166.1976, 158.7227, 
    151.6122, 145.0361, 139.0862, 133.7852, 129.1075, 125, 121.3986, 118.238, 
    115.457, 113.0015, 110.8243, 108.8855, 107.1511, 105.5927, 104.1863, 
    102.9118, 101.7523, 100.6933, 99.72258, 98.82985, 98.00616, 97.24386, 
    96.53635, 95.87792, 95.2636, 94.68904, 94.15043, 93.64443, 93.16808, 
    92.71877, 92.29418, 91.89223, 91.51109, 91.14906, 90.8047, 90.47663, 
    90.16367, 89.86469, 89.57872, 89.30485, 89.04224, 88.79016, 88.5479, 
    88.31486, 88.09042, 87.87408,
  253.1703, 252.9821, 252.7867, 252.5838, 252.3728, 252.1532, 251.9243, 
    251.6855, 251.4361, 251.1752, 250.902, 250.6154, 250.3145, 249.9979, 
    249.6644, 249.3125, 248.9404, 248.5464, 248.1282, 247.6836, 247.2099, 
    246.7038, 246.1621, 245.5805, 244.9546, 244.279, 243.5474, 242.7526, 
    241.8862, 240.938, 239.8962, 238.7466, 237.4723, 236.0526, 234.4629, 
    232.6729, 230.6458, 228.3365, 225.6902, 222.6403, 219.1075, 215, 
    210.2177, 204.6628, 198.2614, 190.9996, 182.9671, 174.3886, 165.6114, 
    157.0329, 149.0004, 141.7386, 135.3372, 129.7823, 125, 120.8926, 
    117.3597, 114.3098, 111.6635, 109.3542, 107.3271, 105.5371, 103.9474, 
    102.5277, 101.2534, 100.1038, 99.062, 98.11382, 97.24737, 96.4526, 
    95.72102, 95.04538, 94.41947, 93.83794, 93.29617, 92.79015, 92.31637, 
    91.87176, 91.45362, 91.05958, 90.68752, 90.33557, 90.00206, 89.6855, 
    89.38454, 89.098, 88.82478, 88.5639, 88.31446, 88.07568, 87.84682, 
    87.62719, 87.4162, 87.21329, 87.01794, 86.82967,
  254.2171, 254.0572, 253.8913, 253.7189, 253.5396, 253.353, 253.1584, 
    252.9553, 252.743, 252.521, 252.2883, 252.0443, 251.7878, 251.5178, 
    251.2333, 250.9328, 250.615, 250.2781, 249.9204, 249.5397, 249.1336, 
    248.6994, 248.234, 247.7337, 247.1945, 246.6115, 245.9791, 245.2905, 
    244.5381, 243.7124, 242.8023, 241.7944, 240.6723, 239.4162, 238.0012, 
    236.397, 234.5652, 232.4577, 230.0134, 227.1551, 223.7852, 219.7823, 215, 
    209.274, 202.4456, 194.4155, 185.2328, 175.1859, 164.8141, 154.7672, 
    145.5845, 137.5544, 130.726, 125, 120.2177, 116.2148, 112.8449, 109.9866, 
    107.5423, 105.4348, 103.603, 101.9988, 100.5838, 99.32767, 98.20561, 
    97.1977, 96.28763, 95.46194, 94.70948, 94.02094, 93.38848, 92.80547, 
    92.26626, 91.76603, 91.30061, 90.86642, 90.46033, 90.0796, 89.72186, 
    89.385, 89.06716, 88.76671, 88.48216, 88.21223, 87.95574, 87.71165, 
    87.479, 87.25695, 87.04473, 86.84164, 86.64705, 86.46037, 86.28109, 
    86.10871, 85.94279, 85.78294,
  255.2658, 255.1346, 254.9984, 254.8569, 254.7097, 254.5564, 254.3966, 
    254.2297, 254.0552, 253.8727, 253.6813, 253.4805, 253.2693, 253.0471, 
    252.8126, 252.565, 252.3028, 252.0248, 251.7294, 251.4148, 251.0789, 
    250.7194, 250.3337, 249.9187, 249.4708, 248.9858, 248.4588, 247.884, 
    247.2546, 246.5622, 245.797, 244.9467, 243.9966, 242.9281, 241.7182, 
    240.3377, 238.7491, 236.904, 234.7391, 232.1704, 229.0862, 225.3372, 
    220.726, 215, 207.8628, 199.0359, 188.418, 176.3333, 163.6667, 151.582, 
    140.9641, 132.1372, 125, 119.274, 114.6628, 110.9138, 107.8296, 105.2609, 
    103.096, 101.2509, 99.66229, 98.28175, 97.07185, 96.00339, 95.05325, 
    94.203, 93.43776, 92.7454, 92.11596, 91.5412, 91.01421, 90.52921, 
    90.08129, 89.66628, 89.28058, 88.92112, 88.58524, 88.27059, 87.97516, 
    87.69716, 87.43502, 87.18736, 86.95293, 86.73065, 86.51952, 86.31868, 
    86.12733, 85.94476, 85.77032, 85.60345, 85.44359, 85.29028, 85.14307, 
    85.00156, 84.86539, 84.73421,
  256.3161, 256.2139, 256.1077, 255.9973, 255.8825, 255.7629, 255.6382, 
    255.5079, 255.3718, 255.2292, 255.0797, 254.9228, 254.7578, 254.584, 
    254.4007, 254.2069, 254.0017, 253.784, 253.5525, 253.3058, 253.0422, 
    252.7599, 252.4568, 252.1304, 251.7777, 251.3954, 250.9794, 250.525, 
    250.0265, 249.4771, 248.8684, 248.1903, 247.43, 246.5719, 245.5956, 
    244.4755, 243.1777, 241.6576, 239.8548, 237.6863, 235.0361, 231.7386, 
    227.5544, 222.1372, 215, 205.5288, 193.1872, 178.1248, 161.8752, 
    146.8128, 134.4712, 125, 117.8628, 112.4456, 108.2614, 104.9639, 
    102.3137, 100.1452, 98.34243, 96.8223, 95.52452, 94.40438, 93.42815, 
    92.56996, 91.80973, 91.1316, 90.52293, 89.97351, 89.47502, 89.02062, 
    88.60463, 88.22229, 87.8696, 87.54314, 87.24004, 86.9578, 86.69425, 
    86.44754, 86.21603, 85.99831, 85.7931, 85.59932, 85.41596, 85.24218, 
    85.07717, 84.92026, 84.7708, 84.62823, 84.49207, 84.36182, 84.23708, 
    84.11748, 84.00266, 83.8923, 83.78613, 83.68387,
  257.3678, 257.2946, 257.2186, 257.1396, 257.0574, 256.9718, 256.8825, 
    256.7892, 256.6917, 256.5895, 256.4825, 256.37, 256.2517, 256.1271, 
    255.9956, 255.8565, 255.7092, 255.5529, 255.3866, 255.2093, 255.0198, 
    254.8167, 254.5985, 254.3634, 254.1091, 253.8332, 253.5327, 253.204, 
    252.843, 252.4445, 252.0023, 251.5085, 250.9535, 250.3251, 249.6077, 
    248.7808, 247.8175, 246.6812, 245.3214, 243.6666, 241.6122, 239.0004, 
    235.5845, 230.9641, 224.4712, 215, 200.9582, 181.3063, 158.6937, 
    139.0418, 125, 115.5288, 109.0359, 104.4156, 100.9996, 98.3878, 96.33337, 
    94.67856, 93.3188, 92.1825, 91.21916, 90.39229, 89.67486, 89.04649, 
    88.49151, 87.99772, 87.55544, 87.15694, 86.79595, 86.46733, 86.16683, 
    85.89092, 85.63664, 85.40147, 85.18327, 84.98021, 84.79071, 84.6134, 
    84.44711, 84.29077, 84.14349, 84.00444, 83.87292, 83.74831, 83.63001, 
    83.51755, 83.41045, 83.30832, 83.21078, 83.11752, 83.0282, 82.94257, 
    82.86038, 82.7814, 82.70542, 82.63225,
  258.4203, 258.3763, 258.3307, 258.2832, 258.2339, 258.1824, 258.1287, 
    258.0727, 258.014, 257.9526, 257.8882, 257.8206, 257.7495, 257.6745, 
    257.5954, 257.5117, 257.423, 257.3289, 257.2287, 257.1219, 257.0077, 
    256.8853, 256.7537, 256.6118, 256.4582, 256.2915, 256.1099, 255.9111, 
    255.6924, 255.4509, 255.1824, 254.8822, 254.5443, 254.1609, 253.722, 
    253.2145, 252.621, 251.9174, 251.07, 250.0297, 248.7227, 247.0329, 
    244.7672, 241.582, 236.8128, 229.0418, 215, 188.4331, 151.5669, 125, 
    110.9582, 103.1872, 98.41799, 95.2328, 92.96709, 91.27731, 89.97034, 
    88.93002, 88.08257, 87.37898, 86.78548, 86.27804, 85.83914, 85.4557, 
    85.11776, 84.8176, 84.54914, 84.30756, 84.08895, 83.89012, 83.70845, 
    83.54176, 83.38824, 83.24632, 83.11472, 82.99229, 82.87809, 82.77127, 
    82.67111, 82.57698, 82.48832, 82.40464, 82.32552, 82.25054, 82.1794, 
    82.11176, 82.04737, 81.98597, 81.92734, 81.87128, 81.8176, 81.76615, 
    81.71677, 81.66931, 81.62366, 81.57971,
  259.4734, 259.4587, 259.4435, 259.4276, 259.4112, 259.394, 259.3761, 
    259.3574, 259.3379, 259.3174, 259.2959, 259.2733, 259.2495, 259.2245, 
    259.1981, 259.1702, 259.1406, 259.1092, 259.0757, 259.04, 259.0019, 
    258.961, 258.917, 258.8695, 258.8182, 258.7625, 258.7017, 258.6351, 
    258.5619, 258.481, 258.3909, 258.2902, 258.1767, 258.0478, 257.9001, 
    257.729, 257.5284, 257.2901, 257.002, 256.6468, 256.1976, 255.6114, 
    254.8141, 253.6667, 251.8752, 248.6937, 241.5669, 215, 125, 98.43307, 
    91.30631, 88.12482, 86.3333, 85.18594, 84.38862, 83.8024, 83.3532, 
    82.99795, 82.70988, 82.47154, 82.27102, 82.09992, 81.95218, 81.82327, 
    81.70978, 81.60906, 81.51905, 81.4381, 81.36489, 81.29834, 81.23755, 
    81.1818, 81.13046, 81.08302, 81.03903, 80.99813, 80.95998, 80.92429, 
    80.89085, 80.85941, 80.82981, 80.80188, 80.77547, 80.75044, 80.7267, 
    80.70412, 80.68264, 80.66216, 80.64259, 80.62389, 80.60598, 80.58882, 
    80.57234, 80.55652, 80.54129, 80.52663,
  260.5266, 260.5413, 260.5565, 260.5724, 260.5888, 260.606, 260.6239, 
    260.6426, 260.6621, 260.6826, 260.7041, 260.7267, 260.7505, 260.7755, 
    260.8019, 260.8298, 260.8594, 260.8908, 260.9243, 260.96, 260.9981, 
    261.039, 261.083, 261.1305, 261.1818, 261.2375, 261.2983, 261.3649, 
    261.4381, 261.519, 261.6091, 261.7098, 261.8233, 261.9522, 262.0999, 
    262.271, 262.4716, 262.7099, 262.998, 263.3532, 263.8024, 264.3886, 
    265.1859, 266.3333, 268.1248, 271.3063, 278.4331, 305, 35, 61.56694, 
    68.69369, 71.87518, 73.6667, 74.81406, 75.61138, 76.1976, 76.6468, 
    77.00205, 77.29012, 77.52846, 77.72898, 77.90008, 78.04782, 78.17673, 
    78.29022, 78.39094, 78.48095, 78.5619, 78.63511, 78.70166, 78.76245, 
    78.8182, 78.86954, 78.91698, 78.96097, 79.00187, 79.04002, 79.07571, 
    79.10915, 79.14059, 79.17019, 79.19812, 79.22453, 79.24956, 79.2733, 
    79.29588, 79.31736, 79.33784, 79.35741, 79.37611, 79.39402, 79.41118, 
    79.42766, 79.44348, 79.45871, 79.47337,
  261.5797, 261.6237, 261.6693, 261.7168, 261.7661, 261.8176, 261.8713, 
    261.9273, 261.986, 262.0474, 262.1118, 262.1794, 262.2505, 262.3255, 
    262.4046, 262.4883, 262.577, 262.6711, 262.7713, 262.8781, 262.9923, 
    263.1147, 263.2463, 263.3882, 263.5418, 263.7085, 263.8901, 264.089, 
    264.3076, 264.5491, 264.8176, 265.1178, 265.4557, 265.8391, 266.278, 
    266.7855, 267.379, 268.0826, 268.93, 269.9703, 271.2773, 272.9671, 
    275.2328, 278.418, 283.1872, 290.9582, 305, 331.5669, 8.433065, 35, 
    49.04179, 56.81278, 61.58201, 64.7672, 67.03291, 68.72269, 70.02966, 
    71.06998, 71.91743, 72.62102, 73.21452, 73.72196, 74.16086, 74.5443, 
    74.88224, 75.1824, 75.45086, 75.69244, 75.91105, 76.10988, 76.29155, 
    76.45824, 76.61176, 76.75368, 76.88528, 77.00771, 77.12191, 77.22873, 
    77.32889, 77.42302, 77.51168, 77.59536, 77.67448, 77.74946, 77.8206, 
    77.88824, 77.95263, 78.01403, 78.07266, 78.12872, 78.1824, 78.23385, 
    78.28323, 78.33069, 78.37634, 78.42029,
  262.6322, 262.7054, 262.7814, 262.8604, 262.9426, 263.0282, 263.1175, 
    263.2108, 263.3083, 263.4105, 263.5175, 263.63, 263.7483, 263.8729, 
    264.0044, 264.1435, 264.2908, 264.4471, 264.6134, 264.7907, 264.9802, 
    265.1833, 265.4015, 265.6366, 265.8909, 266.1668, 266.4673, 266.796, 
    267.157, 267.5555, 267.9977, 268.4915, 269.0465, 269.6749, 270.3923, 
    271.2192, 272.1825, 273.3188, 274.6786, 276.3334, 278.3878, 280.9996, 
    284.4156, 289.0359, 295.5288, 305, 319.0418, 338.6937, 1.30631, 20.95822, 
    35, 44.47124, 50.96407, 55.58445, 59.00039, 61.6122, 63.66663, 65.32144, 
    66.6812, 67.8175, 68.78084, 69.60771, 70.32514, 70.95351, 71.50849, 
    72.00228, 72.44456, 72.84306, 73.20405, 73.53267, 73.83317, 74.10908, 
    74.36336, 74.59853, 74.81673, 75.01979, 75.20929, 75.3866, 75.55289, 
    75.70923, 75.85651, 75.99556, 76.12708, 76.25169, 76.36999, 76.48245, 
    76.58955, 76.69168, 76.78922, 76.88248, 76.9718, 77.05743, 77.13962, 
    77.2186, 77.29458, 77.36775,
  263.6839, 263.7861, 263.8923, 264.0027, 264.1175, 264.2371, 264.3618, 
    264.4921, 264.6282, 264.7708, 264.9203, 265.0772, 265.2422, 265.416, 
    265.5993, 265.7931, 265.9983, 266.216, 266.4475, 266.6942, 266.9578, 
    267.2401, 267.5432, 267.8696, 268.2223, 268.6046, 269.0206, 269.475, 
    269.9735, 270.5229, 271.1316, 271.8097, 272.57, 273.4281, 274.4044, 
    275.5245, 276.8223, 278.3424, 280.1453, 282.3137, 284.9639, 288.2614, 
    292.4456, 297.8628, 305, 314.4712, 326.8128, 341.8752, 358.1248, 
    13.18722, 25.52876, 35, 42.1372, 47.55444, 51.73862, 55.03613, 57.68631, 
    59.85475, 61.65757, 63.17771, 64.47548, 65.59562, 66.57185, 67.43004, 
    68.19027, 68.8684, 69.47707, 70.02649, 70.52498, 70.97938, 71.39537, 
    71.77771, 72.1304, 72.45686, 72.75996, 73.0422, 73.30575, 73.55246, 
    73.78397, 74.00169, 74.2069, 74.40068, 74.58404, 74.75782, 74.92283, 
    75.07974, 75.2292, 75.37177, 75.50793, 75.63818, 75.76292, 75.88252, 
    75.99734, 76.1077, 76.21387, 76.31613,
  264.7342, 264.8654, 265.0016, 265.1431, 265.2903, 265.4436, 265.6035, 
    265.7703, 265.9448, 266.1273, 266.3187, 266.5195, 266.7307, 266.9529, 
    267.1873, 267.435, 267.6972, 267.9752, 268.2706, 268.5852, 268.9211, 
    269.2806, 269.6663, 270.0813, 270.5292, 271.0142, 271.5412, 272.116, 
    272.7454, 273.4378, 274.203, 275.0533, 276.0034, 277.0719, 278.2817, 
    279.6623, 281.2509, 283.096, 285.2609, 287.8296, 290.9138, 294.6628, 
    299.274, 305, 312.1372, 320.9641, 331.582, 343.6667, 356.3333, 8.417991, 
    19.03593, 27.8628, 35, 40.72601, 45.33723, 49.08622, 52.17041, 54.73909, 
    56.90404, 58.74911, 60.33771, 61.71825, 62.92815, 63.99661, 64.94675, 
    65.797, 66.56224, 67.2546, 67.88404, 68.4588, 68.98579, 69.47079, 
    69.91871, 70.33372, 70.71942, 71.07888, 71.41476, 71.72941, 72.02484, 
    72.30284, 72.56498, 72.81264, 73.04707, 73.26935, 73.48048, 73.68132, 
    73.87267, 74.05524, 74.22968, 74.39655, 74.55641, 74.70972, 74.85693, 
    74.99844, 75.13461, 75.26579,
  265.7829, 265.9428, 266.1087, 266.2811, 266.4604, 266.6471, 266.8416, 
    267.0447, 267.257, 267.479, 267.7116, 267.9557, 268.2122, 268.4822, 
    268.7667, 269.0672, 269.385, 269.7219, 270.0796, 270.4603, 270.8664, 
    271.3006, 271.766, 272.2663, 272.8055, 273.3885, 274.0209, 274.7095, 
    275.4619, 276.2876, 277.1977, 278.2056, 279.3277, 280.5839, 281.9988, 
    283.603, 285.4348, 287.5423, 289.9866, 292.8449, 296.2148, 300.2177, 305, 
    310.726, 317.5544, 325.5844, 334.7672, 344.8141, 355.1859, 5.232795, 
    14.41555, 22.44556, 29.27399, 35, 39.78226, 43.7852, 47.1551, 50.01339, 
    52.45767, 54.56522, 56.39701, 58.00124, 59.41615, 60.67233, 61.79439, 
    62.8023, 63.71237, 64.53806, 65.29052, 65.97906, 66.61152, 67.19453, 
    67.73374, 68.23397, 68.69939, 69.13358, 69.53967, 69.9204, 70.27814, 
    70.615, 70.93284, 71.23329, 71.51784, 71.78777, 72.04426, 72.28835, 
    72.521, 72.74305, 72.95527, 73.15836, 73.35295, 73.53963, 73.71891, 
    73.89129, 74.05721, 74.21706,
  266.8297, 267.0179, 267.2133, 267.4162, 267.6272, 267.8468, 268.0757, 
    268.3145, 268.5639, 268.8248, 269.098, 269.3846, 269.6855, 270.0021, 
    270.3356, 270.6875, 271.0596, 271.4536, 271.8718, 272.3164, 272.7902, 
    273.2962, 273.838, 274.4195, 275.0454, 275.721, 276.4526, 277.2474, 
    278.1138, 279.062, 280.1038, 281.2534, 282.5277, 283.9474, 285.5371, 
    287.3271, 289.3542, 291.6635, 294.3098, 297.3597, 300.8925, 305, 
    309.7823, 315.3372, 321.7386, 329.0004, 337.0329, 345.6114, 354.3886, 
    2.967087, 10.99961, 18.26138, 24.66276, 30.21773, 35, 39.10745, 42.64027, 
    45.6902, 48.33653, 50.64579, 52.6729, 54.46289, 56.05262, 57.47225, 
    58.74662, 59.8962, 60.938, 61.88618, 62.75264, 63.5474, 64.27898, 
    64.95462, 65.58053, 66.16206, 66.70383, 67.20985, 67.68363, 68.12824, 
    68.54638, 68.94042, 69.31248, 69.66443, 69.99794, 70.3145, 70.61546, 
    70.902, 71.17522, 71.4361, 71.68554, 71.92432, 72.15318, 72.37281, 
    72.5838, 72.78671, 72.98206, 73.17033,
  267.8741, 268.0904, 268.3148, 268.5479, 268.7902, 269.0422, 269.3048, 
    269.5787, 269.8647, 270.1637, 270.4766, 270.8047, 271.1491, 271.5111, 
    271.8922, 272.2942, 272.7188, 273.1681, 273.6444, 274.1504, 274.689, 
    275.2636, 275.8779, 276.5363, 277.2439, 278.0062, 278.8298, 279.7226, 
    280.6932, 281.7523, 282.9118, 284.1863, 285.5927, 287.1511, 288.8855, 
    290.8243, 293.0015, 295.457, 298.238, 301.3986, 305, 309.1075, 313.7852, 
    319.0862, 325.0361, 331.6122, 338.7227, 346.1976, 353.8024, 1.277307, 
    8.387803, 14.96387, 20.91378, 26.2148, 30.89255, 35, 38.60137, 41.76202, 
    44.54297, 46.99852, 49.17569, 51.11454, 52.84893, 54.40734, 55.81371, 
    57.08818, 58.24773, 59.30675, 60.27742, 61.17015, 61.99385, 62.75614, 
    63.46365, 64.12208, 64.7364, 65.31096, 65.84957, 66.35557, 66.83192, 
    67.28123, 67.70582, 68.10777, 68.48891, 68.85094, 69.1953, 69.52337, 
    69.83633, 70.13531, 70.42128, 70.69515, 70.95776, 71.20984, 71.4521, 
    71.68514, 71.90958, 72.12592,
  268.9158, 269.1599, 269.413, 269.6757, 269.9487, 270.2327, 270.5284, 
    270.8367, 271.1585, 271.4947, 271.8465, 272.215, 272.6016, 273.0078, 
    273.4351, 273.8853, 274.3606, 274.863, 275.3952, 275.9598, 276.5601, 
    277.1996, 277.8823, 278.6129, 279.3965, 280.239, 281.1473, 282.1293, 
    283.194, 284.3517, 285.6147, 286.9972, 288.5153, 290.1884, 292.0387, 
    294.0921, 296.3785, 298.9323, 301.7919, 305, 308.6014, 312.6403, 
    317.1551, 322.1704, 327.6863, 333.6666, 340.0297, 346.6468, 353.3532, 
    359.9703, 6.333375, 12.31369, 17.82959, 22.8449, 27.35973, 31.39863, 35, 
    38.20808, 41.06774, 43.62146, 45.90788, 47.96128, 49.81158, 51.48467, 
    53.00285, 54.38524, 55.64827, 56.80604, 57.87068, 58.85265, 59.76099, 
    60.60354, 61.38712, 62.11768, 62.80042, 63.43991, 64.04021, 64.60484, 
    65.13697, 65.6394, 66.11464, 66.56492, 66.99223, 67.39838, 67.785, 
    68.15353, 68.50529, 68.84151, 69.16328, 69.47156, 69.76728, 70.05127, 
    70.32429, 70.58703, 70.84013, 71.08418,
  269.9545, 270.2259, 270.5072, 270.7991, 271.1024, 271.4176, 271.7458, 
    272.0877, 272.4444, 272.817, 273.2065, 273.6143, 274.0419, 274.4907, 
    274.9626, 275.4594, 275.9832, 276.5364, 277.1217, 277.742, 278.4006, 
    279.1012, 279.8479, 280.6456, 281.4994, 282.4155, 283.4008, 284.463, 
    285.6112, 286.8556, 288.2079, 289.6816, 291.2922, 293.0573, 294.9969, 
    297.1341, 299.4944, 302.1061, 305, 308.2081, 311.762, 315.6902, 320.0134, 
    324.7391, 329.8547, 335.3214, 341.07, 347.002, 352.998, 358.93, 4.678558, 
    10.14525, 15.26091, 19.9866, 24.3098, 28.23798, 31.79192, 35, 37.89388, 
    40.50561, 42.86588, 45.00304, 46.94274, 48.70781, 50.31837, 51.7921, 
    53.14442, 54.3888, 55.53698, 56.59922, 57.58447, 58.50058, 59.35443, 
    60.15207, 60.89882, 61.5994, 62.25798, 62.87827, 63.46357, 64.01681, 
    64.54063, 65.03741, 65.50926, 65.9581, 66.38566, 66.7935, 67.18303, 
    67.55556, 67.91226, 68.2542, 68.58237, 68.89764, 69.20087, 69.49279, 
    69.7741, 70.04546,
  270.9899, 271.2881, 271.5972, 271.9177, 272.2505, 272.5964, 272.9563, 
    273.331, 273.7218, 274.1296, 274.5558, 275.0016, 275.4688, 275.9587, 
    276.4733, 277.0146, 277.5849, 278.1864, 278.8221, 279.4949, 280.2082, 
    280.9659, 281.772, 282.6315, 283.5496, 284.5325, 285.5868, 286.7203, 
    287.9417, 289.2607, 290.6886, 292.2379, 293.9227, 295.7589, 297.7643, 
    299.9584, 302.3627, 305, 307.8939, 311.0677, 314.543, 318.3365, 322.4577, 
    326.904, 331.6576, 336.6812, 341.9174, 347.2901, 352.7099, 358.0826, 
    3.318798, 8.342426, 13.09596, 17.54233, 21.66347, 25.45703, 28.93226, 
    32.10612, 35, 37.63727, 40.04157, 42.23573, 44.24112, 46.07734, 47.76212, 
    49.31137, 50.73925, 52.05832, 53.2797, 54.4132, 55.46753, 56.45037, 
    57.36851, 58.22799, 59.03416, 59.79178, 60.5051, 61.17789, 61.81356, 
    62.41513, 62.98535, 63.52666, 64.0413, 64.53126, 64.99835, 65.44424, 
    65.87041, 66.27824, 66.66897, 67.04373, 67.40359, 67.74947, 68.08229, 
    68.40284, 68.71187, 69.01007,
  272.0217, 272.3462, 272.6824, 273.031, 273.3927, 273.7685, 274.1592, 
    274.5659, 274.9897, 275.4317, 275.8933, 276.3759, 276.881, 277.4105, 
    277.966, 278.5498, 279.1641, 279.8114, 280.4945, 281.2166, 281.9809, 
    282.7914, 283.6523, 284.5683, 285.5446, 286.5874, 287.703, 288.8989, 
    290.1834, 291.5657, 293.0562, 294.6662, 296.4086, 298.2973, 300.3477, 
    302.5761, 305, 307.6373, 310.5056, 313.6215, 316.9985, 320.6458, 
    324.5652, 328.7491, 333.1777, 337.8175, 342.621, 347.5284, 352.4716, 
    357.379, 2.182494, 6.822294, 11.25089, 15.43478, 19.35421, 23.00148, 
    26.37854, 29.49439, 32.36273, 35, 37.4239, 39.65233, 41.70267, 43.5914, 
    45.33379, 46.94384, 48.43428, 49.81659, 51.10109, 52.29701, 53.41263, 
    54.45534, 55.43174, 56.34774, 57.20862, 58.01911, 58.78346, 59.50549, 
    60.1886, 60.83591, 61.4502, 62.03398, 62.58954, 63.11895, 63.62409, 
    64.10667, 64.56827, 65.0103, 65.43406, 65.84076, 66.2315, 66.60727, 
    66.96902, 67.3176, 67.65379, 67.97832,
  273.0494, 273.3998, 273.7626, 274.1385, 274.5285, 274.9333, 275.3541, 
    275.7918, 276.2476, 276.7226, 277.2184, 277.7362, 278.2778, 278.8449, 
    279.4395, 280.0635, 280.7195, 281.4098, 282.1374, 282.9053, 283.7169, 
    284.576, 285.4869, 286.454, 287.4827, 288.5785, 289.7478, 290.9976, 
    292.3356, 293.7704, 295.3112, 296.9687, 298.7537, 300.6786, 302.7562, 
    305, 307.4239, 310.0416, 312.8659, 315.9079, 319.1757, 322.6729, 326.397, 
    330.3377, 334.4755, 338.7808, 343.2145, 347.729, 352.271, 356.7855, 
    1.219163, 5.524519, 9.662291, 13.60299, 17.3271, 20.82431, 24.09212, 
    27.13412, 29.95843, 32.5761, 35, 37.24382, 39.3214, 41.24627, 43.03135, 
    44.68874, 46.22965, 47.66441, 49.0024, 50.25218, 51.42148, 52.5173, 
    53.54596, 54.51313, 55.42397, 56.28311, 57.09473, 57.86261, 58.59017, 
    59.28052, 59.93645, 60.56054, 61.15507, 61.72218, 62.26379, 62.78166, 
    63.27739, 63.75245, 64.20821, 64.64589, 65.06664, 65.47151, 65.86147, 
    66.23743, 66.6002, 66.95055,
  274.073, 274.4485, 274.8373, 275.2399, 275.6573, 276.0905, 276.5403, 
    277.008, 277.4946, 278.0015, 278.53, 279.0817, 279.6581, 280.2611, 
    280.8926, 281.5547, 282.2498, 282.9805, 283.7494, 284.5598, 285.4148, 
    286.3184, 287.2744, 288.2875, 289.3625, 290.5049, 291.7205, 293.016, 
    294.3984, 295.8756, 297.456, 299.1486, 300.9632, 302.9101, 305, 307.2438, 
    309.6523, 312.2357, 315.0031, 317.9613, 321.1145, 324.4629, 328.0012, 
    331.7183, 335.5956, 339.6077, 343.722, 347.9001, 352.0999, 356.278, 
    0.3922898, 4.404378, 8.281747, 11.99876, 15.53711, 18.88546, 22.03872, 
    24.99696, 27.76427, 30.34767, 32.75618, 35, 37.08991, 39.03682, 40.85144, 
    42.54405, 44.12439, 45.60155, 46.98399, 48.27946, 49.49513, 50.63749, 
    51.7125, 52.72558, 53.68164, 54.58518, 55.44026, 56.25058, 57.01952, 
    57.75015, 58.44526, 59.1074, 59.7389, 60.34189, 60.91832, 61.46997, 
    61.99849, 62.50537, 62.992, 63.45966, 63.90952, 64.34265, 64.76008, 
    65.16272, 65.55144, 65.92702,
  275.0919, 275.4922, 275.9062, 276.3348, 276.7789, 277.2394, 277.7174, 
    278.214, 278.7303, 279.2677, 279.8276, 280.4116, 281.0211, 281.6581, 
    282.3245, 283.0224, 283.7542, 284.5222, 285.3295, 286.1788, 287.0736, 
    288.0173, 289.0139, 290.0677, 291.1834, 292.366, 293.6211, 294.9546, 
    296.373, 297.8834, 299.4932, 301.2103, 303.043, 305, 307.0899, 309.3214, 
    311.7027, 314.2411, 316.9427, 319.8116, 322.8489, 326.0526, 329.4161, 
    332.9281, 336.5719, 340.3251, 344.1609, 348.0478, 351.9522, 355.8391, 
    359.6749, 3.428143, 7.071855, 10.58385, 13.94739, 17.15107, 20.18842, 
    23.05726, 25.75888, 28.29732, 30.6786, 32.91009, 35, 36.95695, 38.78968, 
    40.50679, 42.11657, 43.62696, 45.04543, 46.37894, 47.634, 48.81659, 
    49.93225, 50.98606, 51.9827, 52.92643, 53.82118, 54.67052, 55.47775, 
    56.24585, 56.9776, 57.67552, 58.34191, 58.9789, 59.58846, 60.17235, 
    60.73225, 61.26968, 61.78603, 62.28261, 62.76061, 63.22114, 63.66523, 
    64.09383, 64.50784, 64.90805,
  276.1061, 276.5303, 276.9689, 277.4227, 277.8926, 278.3796, 278.8848, 
    279.4092, 279.954, 280.5207, 281.1105, 281.7251, 282.366, 283.0351, 
    283.7343, 284.4657, 285.2315, 286.0343, 286.8767, 287.7617, 288.6923, 
    289.6721, 290.7048, 291.7943, 292.9452, 294.162, 295.4499, 296.8143, 
    298.2611, 299.7964, 301.4268, 303.159, 305, 306.957, 309.0368, 311.2463, 
    313.5914, 316.0773, 318.7078, 321.4847, 324.4073, 327.4723, 330.6723, 
    333.9966, 337.43, 340.9535, 344.5443, 348.1767, 351.8233, 355.4557, 
    359.0465, 2.569962, 6.003388, 9.32767, 12.52775, 15.59266, 18.51533, 
    21.29219, 23.92266, 26.4086, 28.75373, 30.96318, 33.04305, 35, 36.84104, 
    38.57323, 40.20359, 41.73889, 43.18566, 44.55008, 45.83797, 47.0548, 
    48.20564, 49.29521, 50.32788, 51.30768, 52.23835, 53.1233, 53.96572, 
    54.76851, 55.53435, 56.26572, 56.96489, 57.63398, 58.2749, 58.88946, 
    59.4793, 60.04595, 60.59082, 61.11523, 61.62037, 62.10738, 62.5773, 
    63.03111, 63.46969, 63.89391,
  277.1151, 277.5627, 278.0251, 278.5034, 278.9982, 279.5108, 280.042, 
    280.5931, 281.1653, 281.7598, 282.3781, 283.0217, 283.6922, 284.3914, 
    285.1213, 285.8838, 286.6812, 287.5158, 288.3904, 289.3076, 290.2705, 
    291.2824, 292.3467, 293.4673, 294.6481, 295.8935, 297.2082, 298.5969, 
    300.065, 301.6178, 303.2608, 305, 306.841, 308.7897, 310.8514, 313.0313, 
    315.3338, 317.7621, 320.3184, 323.0028, 325.8137, 328.7466, 331.7944, 
    334.9467, 338.1903, 341.5085, 344.8822, 348.2902, 351.7098, 355.1178, 
    358.4915, 1.809731, 5.053253, 8.20561, 11.25338, 14.18629, 16.99715, 
    19.68163, 22.23788, 24.66621, 26.96865, 29.14856, 31.21031, 33.15896, 35, 
    36.73916, 38.38225, 39.93501, 41.40307, 42.79184, 44.10649, 45.35192, 
    46.53275, 47.65329, 48.71761, 49.72948, 50.69239, 51.60961, 52.48415, 
    53.31882, 54.1162, 54.8787, 55.60854, 56.30777, 56.9783, 57.6219, 
    58.2402, 58.83472, 59.40688, 59.95797, 60.48923, 61.00177, 61.49665, 
    61.97486, 62.43731, 62.88485,
  278.1189, 278.5891, 279.0746, 279.5764, 280.0953, 280.6324, 281.1887, 
    281.7654, 282.3635, 282.9845, 283.6298, 284.3008, 284.9991, 285.7266, 
    286.4849, 287.2762, 288.1026, 288.9664, 289.8701, 290.8163, 291.8079, 
    292.8479, 293.9397, 295.0867, 296.2926, 297.5614, 298.8972, 300.3043, 
    301.7874, 303.351, 305, 306.7392, 308.5732, 310.5068, 312.544, 314.6888, 
    316.9438, 319.3114, 321.7921, 324.3853, 327.0882, 329.8962, 332.8023, 
    335.797, 338.8684, 342.0023, 345.1824, 348.3909, 351.6091, 354.8176, 
    357.9977, 1.131602, 4.203004, 7.197704, 10.1038, 12.91182, 15.61476, 
    18.2079, 20.68863, 23.05616, 25.31126, 27.45595, 29.49321, 31.42676, 
    33.26084, 35, 36.64899, 38.21262, 39.69566, 41.10281, 42.43859, 43.70737, 
    44.91329, 46.06028, 47.15206, 48.19212, 49.18372, 50.12992, 51.03359, 
    51.89737, 52.72377, 53.51507, 54.27343, 55.00086, 55.6992, 56.3702, 
    57.01546, 57.63647, 58.23465, 58.81128, 59.36757, 59.90467, 60.42362, 
    60.92541, 61.41096, 61.88113,
  279.117, 279.6091, 280.117, 280.6415, 281.1836, 281.7442, 282.3245, 
    282.9254, 283.5484, 284.1945, 284.8652, 285.5619, 286.2863, 287.0399, 
    287.8247, 288.6425, 289.4954, 290.3856, 291.3155, 292.2875, 293.3043, 
    294.3689, 295.4841, 296.6533, 297.8797, 299.167, 300.5188, 301.9389, 
    303.4313, 305, 306.649, 308.3822, 310.2036, 312.1166, 314.1244, 316.2296, 
    318.4343, 320.7393, 323.1444, 325.6483, 328.2477, 330.938, 333.7124, 
    336.5622, 339.4771, 342.4445, 345.4509, 348.481, 351.519, 354.5491, 
    357.5555, 0.5229301, 3.43776, 6.287628, 9.062004, 11.75227, 14.35173, 
    16.85558, 19.26074, 21.56572, 23.77035, 25.87561, 27.88343, 29.79641, 
    31.61775, 33.35101, 35, 36.56869, 38.06109, 39.48121, 40.83299, 42.12026, 
    43.34671, 44.51587, 45.63113, 46.69568, 47.71254, 48.68455, 49.6144, 
    50.50459, 51.35749, 52.1753, 52.96007, 53.71373, 54.4381, 55.13484, 
    55.80553, 56.45164, 57.07454, 57.67552, 58.25577, 58.81642, 59.35852, 
    59.88304, 60.39091, 60.88301,
  280.1093, 280.6226, 281.152, 281.6984, 282.2627, 282.8458, 283.4489, 
    284.0731, 284.7194, 285.3892, 286.0838, 286.8046, 287.5532, 288.3311, 
    289.1402, 289.9823, 290.8592, 291.7732, 292.7264, 293.7211, 294.7599, 
    295.8455, 296.9805, 298.1678, 299.4106, 300.7119, 302.075, 303.5032, 305, 
    306.5687, 308.2126, 309.935, 311.7389, 313.627, 315.6016, 317.6644, 
    319.8166, 322.0583, 324.3888, 326.806, 329.3068, 331.8862, 334.5381, 
    337.2546, 340.0265, 342.843, 345.6924, 348.5619, 351.4381, 354.3076, 
    357.157, 359.9735, 2.745399, 5.461938, 8.113825, 10.69325, 13.19396, 
    15.6112, 17.94168, 20.18341, 22.3356, 24.39845, 26.37304, 28.26111, 
    30.06499, 31.78738, 33.43131, 35, 36.49678, 37.92503, 39.28814, 40.58944, 
    41.83219, 43.01954, 44.15452, 45.24004, 46.27887, 47.27363, 48.22681, 
    49.14077, 50.01773, 50.85976, 51.66884, 52.44681, 53.19539, 53.91622, 
    54.61082, 55.28061, 55.92694, 56.55107, 57.15416, 57.73734, 58.30164, 
    58.84803, 59.37743, 59.89069,
  281.0956, 281.6293, 282.1794, 282.7467, 283.3323, 283.937, 284.5618, 
    285.2078, 285.8763, 286.5683, 287.2853, 288.0286, 288.7996, 289.5999, 
    290.4312, 291.2953, 292.1939, 293.1291, 294.1029, 295.1174, 296.1751, 
    297.2783, 298.4294, 299.6313, 300.8864, 302.1977, 303.5679, 305, 
    306.4968, 308.0611, 309.6957, 311.4031, 313.1857, 315.0454, 316.984, 
    319.0024, 321.1011, 323.2797, 325.537, 327.8707, 330.2774, 332.7526, 
    335.2905, 337.884, 340.525, 343.204, 345.911, 348.6351, 351.3649, 
    354.089, 356.796, 359.475, 2.115962, 4.709482, 7.247366, 9.722579, 
    12.12932, 14.46302, 16.7203, 18.89891, 20.9976, 23.01601, 24.95457, 
    26.81434, 28.59693, 30.30434, 31.93891, 33.50322, 35, 36.43207, 37.80231, 
    39.11358, 40.36873, 41.57055, 42.72173, 43.82489, 44.88256, 45.89714, 
    46.87091, 47.80608, 48.7047, 49.56874, 50.40006, 51.20041, 51.97144, 
    52.7147, 53.43167, 54.12373, 54.79218, 55.43823, 56.06305, 56.66772, 
    57.25326, 57.82062, 58.37072, 58.90441,
  282.0757, 282.629, 283.1989, 283.7864, 284.3922, 285.0173, 285.6627, 
    286.3295, 287.0187, 287.7316, 288.4694, 289.2335, 290.0252, 290.846, 
    291.6976, 292.5815, 293.4994, 294.4533, 295.4451, 296.4767, 297.5502, 
    298.6679, 299.832, 301.0449, 302.3088, 303.6264, 305, 306.4321, 307.925, 
    309.4812, 311.1028, 312.7918, 314.5501, 316.3789, 318.2795, 320.2522, 
    322.297, 324.4132, 326.5992, 328.8527, 331.1702, 333.5474, 335.9791, 
    338.4588, 340.9794, 343.5327, 346.1099, 348.7017, 351.2983, 353.8901, 
    356.4673, 359.0206, 1.541195, 4.02094, 6.452599, 8.829846, 11.14735, 
    13.40078, 15.5868, 17.70299, 19.74782, 21.72053, 23.62106, 25.44992, 
    27.20815, 28.89719, 30.51879, 32.07497, 33.56793, 35, 36.37359, 37.69115, 
    38.95514, 40.16799, 41.3321, 42.44979, 43.52334, 44.55494, 45.54667, 
    46.50057, 47.41854, 48.30243, 49.15396, 49.9748, 50.76651, 51.53057, 
    52.26839, 52.98129, 53.67054, 54.33731, 54.98272, 55.60782, 56.21362, 
    56.80106, 57.37103, 57.92436,
  283.0493, 283.6215, 284.2104, 284.817, 285.4421, 286.0866, 286.7515, 
    287.4377, 288.1465, 288.8788, 289.636, 290.4192, 291.2299, 292.0693, 
    292.9391, 293.8407, 294.7758, 295.7461, 296.7533, 297.7992, 298.8859, 
    300.0152, 301.1891, 302.4099, 303.6795, 305, 306.3736, 307.8023, 
    309.2881, 310.833, 312.4386, 314.1065, 315.838, 317.634, 319.4951, 
    321.4215, 323.4126, 325.4675, 327.5845, 329.761, 331.9938, 334.279, 
    336.6115, 338.9858, 341.3954, 343.8332, 346.2915, 348.7625, 351.2375, 
    353.7085, 356.1668, 358.6046, 1.014209, 3.388479, 5.721019, 8.006155, 
    10.23901, 12.41553, 14.53247, 16.58737, 18.57852, 20.50487, 22.366, 
    24.16203, 25.89351, 27.56141, 29.16701, 30.71186, 32.19769, 33.62641, 35, 
    36.32053, 37.59011, 38.81084, 39.98483, 41.11413, 42.20078, 43.24675, 
    44.25394, 45.22419, 46.15928, 47.0609, 47.93068, 48.77015, 49.58081, 
    50.36406, 51.12122, 51.85356, 52.56229, 53.24854, 53.9134, 54.55788, 
    55.18297, 55.78957, 56.37855, 56.95073,
  284.0163, 284.6065, 285.2137, 285.8385, 286.4819, 287.1447, 287.8279, 
    288.5323, 289.2593, 290.0096, 290.7847, 291.5855, 292.4134, 293.2697, 
    294.1558, 295.0732, 296.0232, 297.0075, 298.0278, 299.0856, 300.1828, 
    301.321, 302.502, 303.7278, 305, 306.3205, 307.6912, 309.1136, 310.5894, 
    312.1203, 313.7074, 315.3519, 317.0548, 318.8166, 320.6375, 322.5173, 
    324.4554, 326.4504, 328.5006, 330.6035, 332.7561, 334.9546, 337.1945, 
    339.4708, 341.7777, 344.1091, 346.4582, 348.8182, 351.1818, 353.5418, 
    355.8909, 358.2223, 0.5292088, 2.805467, 5.045379, 7.243857, 9.396461, 
    11.49942, 13.54963, 15.54466, 17.48269, 19.36251, 21.18341, 22.9452, 
    24.64808, 26.29263, 27.87974, 29.41056, 30.88642, 32.30885, 33.67947, 35, 
    36.27223, 37.49796, 38.67902, 39.81722, 40.91436, 41.97219, 42.99245, 
    43.9768, 44.92685, 45.84418, 46.73028, 47.5866, 48.41451, 49.21534, 
    49.99035, 50.74073, 51.46764, 52.17216, 52.85532, 53.51813, 54.1615, 
    54.78633, 55.39347, 55.98371,
  284.9766, 285.584, 286.2085, 286.8506, 287.5113, 288.1913, 288.8917, 
    289.6132, 290.357, 291.1241, 291.9154, 292.7323, 293.5758, 294.4472, 
    295.3478, 296.2789, 297.2419, 298.2381, 299.2692, 300.3365, 301.4417, 
    302.5863, 303.7719, 305, 306.2722, 307.5901, 308.9551, 310.3687, 
    311.8322, 313.3467, 314.9133, 316.5327, 318.2057, 319.9323, 321.7125, 
    323.546, 325.4317, 327.3685, 329.3544, 331.3871, 333.4637, 335.5805, 
    337.7337, 339.9187, 342.1304, 344.3634, 346.6118, 348.8695, 351.1305, 
    353.3882, 355.6366, 357.8696, 0.08128966, 2.266261, 4.419468, 6.536353, 
    8.612883, 10.64557, 12.63149, 14.56826, 16.45404, 18.2875, 20.06775, 
    21.79436, 23.46725, 25.08671, 26.65329, 28.16781, 29.63127, 31.04486, 
    32.40989, 33.72777, 35, 36.22811, 37.41367, 38.55825, 39.66344, 40.7308, 
    41.76188, 42.75816, 43.72113, 44.65221, 45.55278, 46.42419, 47.2677, 
    48.08456, 48.87594, 49.64299, 50.38678, 51.10835, 51.80869, 52.48874, 
    53.1494, 53.79154, 54.41596, 55.02345,
  285.9299, 286.5538, 287.1946, 287.8531, 288.5301, 289.2263, 289.9427, 
    290.6801, 291.4395, 292.2219, 293.0282, 293.8596, 294.7171, 295.6019, 
    296.5151, 297.4581, 298.432, 299.4382, 300.478, 301.5526, 302.6636, 
    303.8123, 305, 306.2281, 307.498, 308.8109, 310.168, 311.5706, 313.0195, 
    314.5159, 316.0603, 317.6533, 319.2952, 320.9861, 322.7256, 324.5131, 
    326.3477, 328.228, 330.1521, 332.1177, 334.1221, 336.162, 338.234, 
    340.3337, 342.4568, 344.5985, 346.7537, 348.917, 351.083, 353.2463, 
    355.4015, 357.5432, 359.6663, 1.766029, 3.837941, 5.877925, 7.882326, 
    9.847935, 11.77201, 13.65226, 15.48687, 17.27442, 19.01393, 20.70479, 
    22.3467, 23.93972, 25.48413, 26.98046, 28.42946, 29.83201, 31.18916, 
    32.50204, 33.77189, 35, 36.1877, 37.33636, 38.44734, 39.52203, 40.56179, 
    41.56797, 42.5419, 43.48486, 44.39812, 45.28292, 46.14042, 46.97178, 
    47.77811, 48.56046, 49.31985, 50.05726, 50.77364, 51.46988, 52.14684, 
    52.80535, 53.44618, 54.0701,
  286.8762, 287.5157, 288.1721, 288.846, 289.5383, 290.2497, 290.981, 
    291.733, 292.5068, 293.3031, 294.123, 294.9673, 295.8373, 296.7338, 
    297.6581, 298.6111, 299.5941, 300.6083, 301.6548, 302.7347, 303.8494, 
    305, 306.1877, 307.4137, 308.679, 309.9848, 311.3321, 312.7217, 314.1545, 
    315.6311, 317.1521, 318.7176, 320.3279, 321.9827, 323.6816, 325.424, 
    327.2086, 329.0341, 330.8988, 332.8004, 334.7364, 336.7038, 338.6994, 
    340.7194, 342.7599, 344.8167, 346.8853, 348.961, 351.039, 353.1147, 
    355.1833, 357.2401, 359.2806, 1.300613, 3.296174, 5.263601, 7.199584, 
    9.101182, 10.96584, 12.79138, 14.57603, 16.31836, 18.0173, 19.67212, 
    21.28238, 22.84794, 24.36887, 25.84548, 27.27827, 28.66791, 30.01517, 
    31.32098, 32.58633, 33.8123, 35, 36.1506, 37.26529, 38.34526, 39.39172, 
    40.40586, 41.38889, 42.34195, 43.26619, 44.16273, 45.03267, 45.87705, 
    46.69691, 47.49323, 48.26696, 49.01904, 49.75033, 50.4617, 51.15397, 
    51.82791, 52.48428, 53.1238,
  287.8153, 288.4696, 289.1407, 289.8291, 290.5357, 291.2611, 292.0062, 
    292.7718, 293.5586, 294.3676, 295.1996, 296.0556, 296.9365, 297.8432, 
    298.7768, 299.7382, 300.7286, 301.7489, 302.8002, 303.8835, 305, 
    306.1506, 307.3364, 308.5583, 309.8172, 311.1141, 312.4498, 313.8249, 
    315.2401, 316.6957, 318.1921, 319.7295, 321.3077, 322.9264, 324.5852, 
    326.2831, 328.0191, 329.7918, 331.5994, 333.4399, 335.311, 337.2098, 
    339.1336, 341.0789, 343.0422, 345.0198, 347.0077, 349.0019, 350.9981, 
    352.9923, 354.9802, 356.9578, 358.9211, 0.8664198, 2.790152, 4.689038, 
    6.560083, 8.4006, 10.20822, 11.98089, 13.71689, 15.41482, 17.07357, 
    18.69232, 20.27052, 21.80788, 23.30432, 24.75996, 26.1751, 27.55021, 
    28.88587, 30.18278, 31.44175, 32.66364, 33.8494, 35, 36.11646, 37.19981, 
    38.25111, 39.27141, 40.26177, 41.22322, 42.1568, 43.06353, 43.94439, 
    44.80036, 45.63238, 46.44137, 47.22821, 47.99377, 48.73887, 49.46433, 
    50.17091, 50.85935, 51.53038, 52.18468,
  288.7472, 289.4154, 290.1002, 290.8022, 291.5222, 292.2607, 293.0185, 
    293.7964, 294.5951, 295.4155, 296.2583, 297.1245, 298.0148, 298.9302, 
    299.8716, 300.8398, 301.8359, 302.8606, 303.915, 305, 306.1165, 307.2653, 
    308.4474, 309.6635, 310.9144, 312.2008, 313.5233, 314.8826, 316.2789, 
    317.7125, 319.1837, 320.6924, 322.2383, 323.8212, 325.4402, 327.0947, 
    328.7834, 330.5051, 332.258, 334.0402, 335.8496, 337.6836, 339.5397, 
    341.4148, 343.3058, 345.2093, 347.1219, 349.04, 350.96, 352.8781, 
    354.7907, 356.6942, 358.5852, 0.4603243, 2.31637, 4.15043, 5.959797, 
    7.742018, 9.494904, 11.21654, 12.90528, 14.55974, 16.17882, 17.76165, 
    19.30761, 20.81628, 22.28746, 23.72113, 25.11744, 26.47666, 27.79922, 
    29.08564, 30.33656, 31.55266, 32.73471, 33.88354, 35, 36.08498, 37.13938, 
    38.16413, 39.16016, 40.1284, 41.06976, 41.98516, 42.8755, 43.74166, 
    44.58451, 45.4049, 46.20364, 46.98153, 47.73935, 48.47785, 49.19776, 
    49.89978, 50.58459, 51.25285,
  289.6716, 290.353, 291.0507, 291.7654, 292.4977, 293.2482, 294.0176, 
    294.8067, 295.6162, 296.4467, 297.2991, 298.1741, 299.0726, 299.9952, 
    300.9429, 301.9164, 302.9165, 303.9441, 305, 306.085, 307.1998, 308.3452, 
    309.522, 310.7308, 311.9722, 313.2467, 314.5549, 315.8971, 317.2736, 
    318.6845, 320.1299, 321.6096, 323.1233, 324.6705, 326.2506, 327.8626, 
    329.5055, 331.1779, 332.8783, 334.6048, 336.3556, 338.1282, 339.9204, 
    341.7294, 343.5525, 345.3866, 347.2287, 349.0757, 350.9243, 352.7713, 
    354.6134, 356.4475, 358.2706, 0.07960072, 1.87176, 3.644429, 5.395164, 
    7.121729, 8.822109, 10.49452, 12.13739, 13.74942, 15.32948, 16.8767, 
    18.39039, 19.87008, 21.31545, 22.72637, 24.10286, 25.44506, 26.75325, 
    28.02781, 29.2692, 30.47797, 31.65474, 32.80019, 33.91502, 35, 36.0559, 
    37.08351, 38.08365, 39.05714, 40.0048, 40.92743, 41.82586, 42.70088, 
    43.55327, 44.38382, 45.19327, 45.98236, 46.75183, 47.50235, 48.23462, 
    48.9493, 49.64702, 50.32841,
  290.5886, 291.2823, 291.992, 292.7184, 293.4621, 294.2237, 295.0037, 
    295.8029, 296.6219, 297.4614, 298.3221, 299.2047, 300.1099, 301.0384, 
    301.9909, 302.9682, 303.971, 305, 306.0559, 307.1394, 308.2511, 309.3917, 
    310.5618, 311.7619, 312.9925, 314.2539, 315.5467, 316.8709, 318.2268, 
    319.6144, 321.0336, 322.4842, 323.9657, 325.4778, 327.0195, 328.5902, 
    330.1886, 331.8136, 333.4636, 335.137, 336.8319, 338.5464, 340.2781, 
    342.0248, 343.784, 345.5529, 347.3289, 349.1092, 350.8908, 352.6711, 
    354.4471, 356.216, 357.9752, 359.7219, 1.453624, 3.168084, 4.863032, 
    6.536436, 8.186443, 9.811396, 11.40983, 12.98048, 14.52226, 16.03428, 
    17.51585, 18.96641, 20.3856, 21.77319, 23.12908, 24.45333, 25.74607, 
    27.00755, 28.23813, 29.43821, 30.60828, 31.74889, 32.86062, 33.9441, 35, 
    36.02899, 37.03178, 38.00909, 38.96163, 39.89013, 40.79531, 41.67789, 
    42.53858, 43.37809, 44.1971, 44.9963, 45.77634, 46.53789, 47.28156, 
    48.00798, 48.71775, 49.41144,
  291.498, 292.2032, 292.9241, 293.6614, 294.4155, 295.1871, 295.9767, 
    296.7849, 297.6124, 298.4597, 299.3275, 300.2164, 301.127, 302.0601, 
    303.0162, 303.9959, 305, 306.029, 307.0835, 308.1641, 309.2714, 310.4059, 
    311.568, 312.7581, 313.9768, 315.2242, 316.5006, 317.8061, 319.1408, 
    320.5046, 321.8974, 323.3188, 324.7685, 326.2458, 327.7502, 329.2805, 
    330.8359, 332.4151, 334.0168, 335.6394, 337.2812, 338.9404, 340.615, 
    342.3028, 344.0017, 345.7092, 347.423, 349.1406, 350.8594, 352.577, 
    354.2908, 355.9983, 357.6972, 359.385, 1.05958, 2.718776, 4.360597, 
    5.983191, 7.584867, 9.164087, 10.71948, 12.24985, 13.75415, 15.2315, 
    16.68118, 18.10262, 19.49541, 20.85923, 22.19392, 23.49943, 24.77581, 
    26.0232, 27.24184, 28.43203, 29.59413, 30.72859, 31.83587, 32.91649, 
    33.97101, 35, 36.00407, 36.98384, 37.93993, 38.87298, 39.78364, 40.67255, 
    41.54034, 42.38765, 43.2151, 44.02333, 44.81293, 45.5845, 46.33863, 
    47.07589, 47.79684, 48.50203,
  292.3998, 293.1156, 293.8469, 294.5941, 295.3578, 296.1384, 296.9366, 
    297.7528, 298.5876, 299.4416, 300.3153, 301.2094, 302.1243, 303.0607, 
    304.019, 305, 306.0041, 307.0318, 308.0836, 309.1602, 310.2618, 311.3889, 
    312.5419, 313.7211, 314.9268, 316.1593, 317.4185, 318.7047, 320.0177, 
    321.3575, 322.7238, 324.1162, 325.5343, 326.9776, 328.4453, 329.9365, 
    331.4502, 332.9854, 334.5406, 336.1147, 337.7058, 339.3125, 340.9328, 
    342.565, 344.2069, 345.8565, 347.5117, 349.1702, 350.8298, 352.4883, 
    354.1435, 355.7931, 357.435, 359.0672, 0.6875198, 2.294184, 3.885358, 
    5.459363, 7.01465, 8.549803, 10.06355, 11.55474, 13.0224, 14.46565, 
    15.8838, 17.27624, 18.64251, 19.98227, 21.2953, 22.58146, 23.84072, 
    25.07315, 26.27887, 27.4581, 28.61111, 29.73823, 30.83984, 31.91635, 
    32.96822, 33.99593, 35, 35.98096, 36.93934, 37.87572, 38.79064, 39.68468, 
    40.55842, 41.41241, 42.24723, 43.06343, 43.86158, 44.64221, 45.40587, 
    46.15308, 46.88437, 47.60023,
  293.2939, 294.0196, 294.7604, 295.5167, 296.289, 297.0777, 297.8834, 
    298.7066, 299.5477, 300.4073, 301.2859, 302.1839, 303.102, 304.0405, 305, 
    305.981, 306.9838, 308.0091, 309.0571, 310.1284, 311.2232, 312.3419, 
    313.4849, 314.6522, 315.8442, 317.0609, 318.3024, 319.5688, 320.8598, 
    322.1753, 323.5151, 324.8787, 326.2657, 327.6755, 329.1074, 330.5605, 
    332.034, 333.5267, 335.0374, 336.5649, 338.1078, 339.6644, 341.2333, 
    342.8127, 344.4007, 345.9956, 347.5954, 349.1981, 350.8019, 352.4046, 
    354.0044, 355.5993, 357.1873, 358.7667, 0.3355702, 1.892236, 3.435082, 
    4.962586, 6.473334, 7.966022, 9.439466, 10.8926, 12.32448, 13.73428, 
    15.1213, 16.48493, 17.8247, 19.14024, 20.43126, 21.69757, 22.9391, 
    24.15582, 25.34779, 26.51514, 27.65805, 28.77678, 29.8716, 30.94286, 
    31.99091, 33.01616, 34.01904, 35, 35.9595, 36.89802, 37.81606, 38.71411, 
    39.59268, 40.45227, 41.2934, 42.11657, 42.92228, 43.71102, 44.4833, 
    45.23958, 45.98036, 46.7061,
  294.1803, 294.9151, 295.6646, 296.4291, 297.2091, 298.005, 298.8173, 
    299.6465, 300.4929, 301.3571, 302.2394, 303.1404, 304.0604, 305, 
    305.9595, 306.9393, 307.9399, 308.9616, 310.0048, 311.0698, 312.1568, 
    313.2662, 314.3981, 315.5528, 316.7303, 317.9307, 319.154, 320.4001, 
    321.6689, 322.9601, 324.2734, 325.6086, 326.9649, 328.3419, 329.7389, 
    331.1551, 332.5895, 334.0413, 335.5093, 336.9922, 338.4889, 339.9979, 
    341.5178, 343.0471, 344.584, 346.1271, 347.6745, 349.2245, 350.7755, 
    352.3255, 353.8729, 355.416, 356.9529, 358.4822, 0.002061171, 1.511083, 
    3.007768, 4.490737, 5.9587, 7.410462, 8.844927, 10.2611, 11.65809, 
    13.03511, 14.39146, 15.72657, 17.03993, 18.33116, 19.59994, 20.84604, 
    22.06932, 23.26972, 24.44721, 25.60187, 26.73381, 27.8432, 28.93024, 
    29.9952, 31.03837, 32.06007, 33.06066, 34.0405, 35, 35.93956, 36.85962, 
    37.7606, 38.64294, 39.5071, 40.35353, 41.18267, 41.99498, 42.79092, 
    43.57091, 44.33541, 45.08487, 45.81969,
  295.059, 295.8021, 296.5594, 297.3313, 298.1181, 298.9203, 299.7383, 
    300.5725, 301.4232, 302.291, 303.1761, 304.079, 305, 305.9396, 306.898, 
    307.8757, 308.873, 309.8901, 310.9274, 311.9852, 313.0635, 314.1627, 
    315.2829, 316.4242, 317.5866, 318.7701, 319.9748, 321.2004, 322.4468, 
    323.7137, 325.0009, 326.3078, 327.634, 328.9789, 330.3419, 331.7222, 
    333.119, 334.5312, 335.9581, 337.3984, 338.8509, 340.3145, 341.7878, 
    343.2693, 344.7578, 346.2517, 347.7495, 349.2495, 350.7505, 352.2505, 
    353.7483, 355.2422, 356.7307, 358.2122, 359.6855, 1.149067, 2.601616, 
    4.041899, 5.468743, 6.881052, 8.277816, 9.65811, 11.0211, 12.36602, 
    13.69223, 14.99914, 16.28627, 17.55319, 18.79959, 20.0252, 21.22985, 
    22.4134, 23.57581, 24.71708, 25.83727, 26.93647, 28.01484, 29.07257, 
    30.10987, 31.12702, 32.12428, 33.10198, 34.06044, 35, 35.92104, 36.82391, 
    37.70902, 38.57675, 39.4275, 40.26167, 41.07965, 41.88187, 42.66872, 
    43.44059, 44.1979, 44.94102,
  295.9299, 296.6805, 297.4449, 298.2233, 299.0161, 299.8238, 300.6465, 
    301.4848, 302.339, 303.2093, 304.0962, 305, 305.921, 306.8596, 307.8161, 
    308.7906, 309.7836, 310.7953, 311.8259, 312.8755, 313.9444, 315.0327, 
    316.1404, 317.2677, 318.4145, 319.5808, 320.7665, 321.9714, 323.1954, 
    324.4381, 325.6992, 326.9783, 328.2749, 329.5884, 330.9183, 332.2638, 
    333.6241, 334.9984, 336.3857, 337.785, 339.1953, 340.6154, 342.0443, 
    343.4805, 344.9228, 346.37, 347.8206, 349.2733, 350.7267, 352.1794, 
    353.63, 355.0772, 356.5195, 357.9557, 359.3846, 0.8046976, 2.215007, 
    3.614345, 5.001646, 6.37591, 7.736207, 9.08168, 10.41155, 11.7251, 
    13.0217, 14.3008, 15.5619, 16.80461, 18.02856, 19.23349, 20.41919, 
    21.58549, 22.7323, 23.85958, 24.96733, 26.05561, 27.1245, 28.17414, 
    29.20469, 30.21636, 31.20936, 32.18394, 33.14038, 34.07896, 35, 35.9038, 
    36.79071, 37.66105, 38.51518, 39.35345, 40.17622, 40.98385, 41.77669, 
    42.55511, 43.31946, 44.07011,
  296.793, 297.5504, 298.321, 299.1052, 299.9032, 300.7154, 301.5421, 
    302.3836, 303.2402, 304.1122, 305, 305.9038, 306.8239, 307.7606, 
    308.7141, 309.6847, 310.6725, 311.6779, 312.7009, 313.7417, 314.8004, 
    315.877, 316.9718, 318.0846, 319.2153, 320.364, 321.5306, 322.7147, 
    323.9162, 325.1348, 326.3702, 327.6219, 328.8895, 330.1724, 331.47, 
    332.7816, 334.1067, 335.4442, 336.7935, 338.1535, 339.5234, 340.902, 
    342.2884, 343.6813, 345.0797, 346.4825, 347.8882, 349.2959, 350.7041, 
    352.1118, 353.5175, 354.9203, 356.3187, 357.7116, 359.098, 0.4766341, 
    1.846476, 3.206508, 4.555761, 5.893324, 7.218343, 8.530026, 9.827646, 
    11.11054, 12.3781, 13.6298, 14.86516, 16.08378, 17.2853, 18.46943, 
    19.63594, 20.78466, 21.91544, 23.02822, 24.12295, 25.19964, 26.25834, 
    27.29912, 28.32211, 29.32745, 30.31532, 31.28589, 32.2394, 33.17609, 
    34.0962, 35, 35.88778, 36.75983, 37.61644, 38.45793, 39.2846, 40.09678, 
    40.89479, 41.67894, 42.44957, 43.20698,
  297.6484, 298.4118, 299.1879, 299.977, 300.7794, 301.5953, 302.425, 
    303.2689, 304.1271, 305, 305.8878, 306.7907, 307.709, 308.6429, 309.5927, 
    310.5584, 311.5403, 312.5386, 313.5533, 314.5845, 315.6324, 316.6969, 
    317.7781, 318.8759, 319.9904, 321.1212, 322.2684, 323.4317, 324.6108, 
    325.8055, 327.0155, 328.2402, 329.4793, 330.7323, 331.9985, 333.2774, 
    334.5683, 335.8704, 337.183, 338.5053, 339.8363, 341.1752, 342.521, 
    343.8727, 345.2292, 346.5895, 347.9526, 349.3174, 350.6826, 352.0474, 
    353.4105, 354.7708, 356.1273, 357.479, 358.8248, 0.1636643, 1.494702, 
    2.816969, 4.129589, 5.43173, 6.722614, 8.001512, 9.267746, 10.5207, 
    11.7598, 12.98454, 14.19447, 15.38918, 16.56833, 17.73161, 18.87879, 
    20.00965, 21.12406, 22.22189, 23.30309, 24.36762, 25.41549, 26.44673, 
    27.46142, 28.45966, 29.44158, 30.40732, 31.35706, 32.29098, 33.20929, 
    34.11222, 35, 35.87288, 36.73111, 37.57496, 38.4047, 39.22061, 40.02298, 
    40.81208, 41.5882, 42.35163,
  298.4959, 299.2647, 300.0455, 300.8388, 301.6447, 302.4636, 303.2956, 
    304.141, 305, 305.8729, 306.7598, 307.661, 308.5768, 309.5071, 310.4523, 
    311.4124, 312.3876, 313.3781, 314.3838, 315.4049, 316.4414, 317.4932, 
    318.5605, 319.643, 320.7407, 321.8535, 322.9813, 324.1237, 325.2806, 
    326.4516, 327.6365, 328.8347, 330.046, 331.2697, 332.5054, 333.7524, 
    335.0103, 336.2782, 337.5556, 338.8415, 340.1353, 341.4361, 342.743, 
    344.0552, 345.3718, 346.6917, 348.014, 349.3379, 350.6621, 351.986, 
    353.3083, 354.6282, 355.9448, 357.257, 358.5639, 359.8647, 1.158482, 
    2.444437, 3.721762, 4.989704, 6.247549, 7.494629, 8.730321, 9.954047, 
    11.16528, 12.36353, 13.54836, 14.71939, 15.87627, 17.01871, 18.14644, 
    19.25927, 20.35701, 21.43955, 22.50677, 23.55863, 24.5951, 25.61618, 
    26.62191, 27.61235, 28.58759, 29.54773, 30.4929, 31.42325, 32.33895, 
    33.24017, 34.12712, 35, 35.85902, 36.70441, 37.53641, 38.35526, 39.16119, 
    39.95446, 40.73534, 41.50406,
  299.3358, 300.109, 300.8939, 301.6906, 302.4994, 303.3204, 304.1538, 305, 
    305.859, 306.7311, 307.6164, 308.5152, 309.4275, 310.3535, 311.2934, 
    312.2472, 313.2151, 314.1971, 315.1933, 316.2036, 317.2282, 318.267, 
    319.3199, 320.3868, 321.4677, 322.5623, 323.6705, 324.7922, 325.9269, 
    327.0746, 328.2346, 329.4069, 330.5908, 331.786, 332.992, 334.2082, 
    335.4341, 336.669, 337.9123, 339.1633, 340.4213, 341.6855, 342.9553, 
    344.2297, 345.5079, 346.7892, 348.0727, 349.3574, 350.6426, 351.9273, 
    353.2108, 354.4921, 355.7703, 357.0447, 358.3145, 359.5787, 0.8367262, 
    2.087737, 3.331035, 4.565938, 5.791796, 7.007998, 8.213969, 9.409175, 
    10.59312, 11.76535, 12.92546, 14.07306, 15.20782, 16.32946, 17.43771, 
    18.53236, 19.61322, 20.68015, 21.73304, 22.77179, 23.79636, 24.80673, 
    25.8029, 26.7849, 27.75277, 28.7066, 29.64647, 30.5725, 31.48482, 
    32.38356, 33.26889, 34.14098, 35, 35.84615, 36.67962, 37.50062, 38.30936, 
    39.10607, 39.89095, 40.66424,
  300.1678, 300.945, 301.7332, 302.5326, 303.3434, 304.1658, 305, 305.8462, 
    306.7044, 307.575, 308.4579, 309.3535, 310.2617, 311.1827, 312.1166, 
    313.0634, 314.0233, 314.9963, 315.9824, 316.9815, 317.9938, 319.019, 
    320.0573, 321.1083, 322.1721, 323.2485, 324.3373, 325.4382, 326.5511, 
    327.6755, 328.8113, 329.958, 331.1152, 332.2826, 333.4597, 334.6459, 
    335.8408, 337.0437, 338.2542, 339.4716, 340.6952, 341.9243, 343.1584, 
    344.3965, 345.6382, 346.8825, 348.1287, 349.3761, 350.6239, 351.8713, 
    353.1175, 354.3618, 355.6035, 356.8416, 358.0757, 359.3048, 0.5284402, 
    1.745796, 2.956268, 4.159237, 5.354114, 6.540341, 7.717392, 8.884773, 
    10.04203, 11.18872, 12.32448, 13.44893, 14.56177, 15.66269, 16.75146, 
    17.82784, 18.89165, 19.94274, 20.98096, 22.00623, 23.01847, 24.01764, 
    25.0037, 25.97667, 26.93657, 27.88343, 28.81733, 29.73833, 30.64655, 
    31.54207, 32.42504, 33.29559, 34.15385, 35, 35.83419, 36.65661, 37.46742, 
    38.26682, 39.05501, 39.83216,
  300.9922, 301.7726, 302.5633, 303.3647, 304.1769, 305, 305.8342, 306.6796, 
    307.5364, 308.4047, 309.2846, 310.1762, 311.0797, 311.995, 312.9223, 
    313.8616, 314.8129, 315.7763, 316.7518, 317.7393, 318.7389, 319.7503, 
    320.7737, 321.8087, 322.8553, 323.9134, 324.9827, 326.063, 327.1542, 
    328.2558, 329.3676, 330.4892, 331.6204, 332.7606, 333.9095, 335.0667, 
    336.2315, 337.4036, 338.5824, 339.7673, 340.9578, 342.1532, 343.3529, 
    344.5564, 345.7629, 346.9718, 348.1824, 349.394, 350.606, 351.8176, 
    353.0282, 354.2371, 355.4436, 356.6471, 357.8468, 359.0422, 0.2327171, 
    1.417635, 2.596416, 3.768503, 4.933362, 6.090485, 7.239392, 8.379629, 
    9.510773, 10.63243, 11.74423, 12.84584, 13.93695, 15.01729, 16.0866, 
    17.14467, 18.19131, 19.22636, 20.24967, 21.26113, 22.26065, 23.24817, 
    24.22366, 25.18707, 26.13842, 27.07773, 28.00501, 28.92034, 29.82378, 
    30.7154, 31.5953, 32.46359, 33.32038, 34.16581, 35, 35.8231, 36.63528, 
    37.43667, 38.22746, 39.00779,
  301.8089, 302.5918, 303.3845, 304.1872, 305, 305.8231, 306.6566, 307.5006, 
    308.3553, 309.2206, 310.0968, 310.9839, 311.8819, 312.7909, 313.711, 
    314.6422, 315.5845, 316.5379, 317.5023, 318.4778, 319.4643, 320.4617, 
    321.4699, 322.4887, 323.5181, 324.5579, 325.6078, 326.6677, 327.7373, 
    328.8164, 329.9047, 331.0018, 332.1074, 333.2211, 334.3427, 335.4715, 
    336.6073, 337.7495, 338.8976, 340.0513, 341.2098, 342.3728, 343.5396, 
    344.7097, 345.8825, 347.0574, 348.2339, 349.4112, 350.5888, 351.7661, 
    352.9426, 354.1175, 355.2903, 356.4604, 357.6272, 358.7902, 359.9487, 
    1.102355, 2.250523, 3.392728, 4.528489, 5.657345, 6.77886, 7.892619, 
    8.998231, 10.09533, 11.18358, 12.26266, 13.33228, 14.39218, 15.44211, 
    16.48187, 17.51126, 18.53012, 19.53829, 20.53567, 21.52215, 22.49765, 
    23.46211, 24.4155, 25.35779, 26.28898, 27.20908, 28.11813, 29.01615, 
    29.90322, 30.77939, 31.64474, 32.49938, 33.34339, 34.1769, 35, 35.81284, 
    36.61554, 37.40824, 38.19109,
  302.618, 303.4027, 304.1967, 305, 305.8128, 306.6353, 307.4674, 308.3094, 
    309.1612, 310.023, 310.8948, 311.7767, 312.6687, 313.5709, 314.4833, 
    315.4059, 316.3386, 317.2816, 318.2346, 319.1978, 320.1709, 321.154, 
    322.1469, 323.1494, 324.1615, 325.183, 326.2136, 327.2533, 328.3016, 
    329.3585, 330.4236, 331.4966, 332.5773, 333.6652, 334.7601, 335.8615, 
    336.969, 338.0823, 339.2009, 340.3243, 341.4521, 342.5838, 343.7189, 
    344.8569, 345.9973, 347.1396, 348.2832, 349.4276, 350.5724, 351.7168, 
    352.8604, 354.0027, 355.1431, 356.2811, 357.4162, 358.5479, 359.6757, 
    0.7991334, 1.917706, 3.030981, 4.138524, 5.239919, 6.334769, 7.422698, 
    8.503347, 9.576381, 10.64148, 11.69836, 12.74674, 13.78638, 14.81703, 
    15.8385, 16.8506, 17.85316, 18.84603, 19.82909, 20.80224, 21.76538, 
    22.71844, 23.66137, 24.59413, 25.51671, 26.42909, 27.33128, 28.22331, 
    29.10521, 29.97702, 30.83881, 31.69064, 32.53258, 33.36472, 34.18716, 35, 
    35.80334, 36.59731, 37.38202,
  303.4195, 304.2054, 305, 305.8033, 306.6155, 307.4367, 308.2668, 309.1061, 
    309.9545, 310.8121, 311.679, 312.5551, 313.4406, 314.3354, 315.2396, 
    316.1531, 317.0759, 318.008, 318.9493, 319.8998, 320.8593, 321.8279, 
    322.8054, 323.7915, 324.7863, 325.7896, 326.8011, 327.8206, 328.848, 
    329.883, 330.9254, 331.9749, 333.0311, 334.0938, 335.1627, 336.2374, 
    337.3176, 338.4028, 339.4928, 340.587, 341.6852, 342.7867, 343.8913, 
    344.9984, 346.1077, 347.2186, 348.3307, 349.4435, 350.5565, 351.6693, 
    352.7814, 353.8923, 355.0016, 356.1087, 357.2133, 358.3148, 359.413, 
    0.5072123, 1.597158, 2.682407, 3.762572, 4.837277, 5.906166, 6.968895, 
    8.025139, 9.074591, 10.11696, 11.15197, 12.17938, 13.19894, 14.21043, 
    15.21367, 16.20846, 17.19465, 18.17209, 19.14065, 20.10022, 21.0507, 
    21.99202, 22.9241, 23.84692, 24.76042, 25.66458, 26.55941, 27.44489, 
    28.32106, 29.18793, 30.04553, 30.89393, 31.73318, 32.56333, 33.38446, 
    34.19666, 35, 35.79459, 36.58051,
  304.2135, 305, 305.7946, 306.5973, 307.4082, 308.2274, 309.055, 309.891, 
    310.7353, 311.5882, 312.4496, 313.3195, 314.1979, 315.0849, 315.9804, 
    316.8844, 317.7968, 318.7177, 319.647, 320.5846, 321.5304, 322.4843, 
    323.4462, 324.416, 325.3935, 326.3785, 327.371, 328.3707, 329.3774, 
    330.3909, 331.4109, 332.4373, 333.4697, 334.5078, 335.5515, 336.6002, 
    337.6538, 338.7119, 339.7741, 340.8401, 341.9096, 342.9821, 344.0572, 
    345.1346, 346.2139, 347.2946, 348.3763, 349.4587, 350.5413, 351.6237, 
    352.7054, 353.7861, 354.8654, 355.9428, 357.0179, 358.0904, 359.1599, 
    0.2258954, 1.28813, 2.346215, 3.399804, 4.448562, 5.492166, 6.530308, 
    7.562692, 8.589039, 9.609083, 10.62257, 11.62928, 12.62897, 13.62145, 
    14.60653, 15.58404, 16.55382, 17.51572, 18.46962, 19.41541, 20.35298, 
    21.28225, 22.20316, 23.11563, 24.01964, 24.91513, 25.8021, 26.68054, 
    27.55043, 28.4118, 29.26466, 30.10905, 30.94499, 31.77254, 32.59176, 
    33.40269, 34.20541, 35, 35.78653,
  305, 305.7865, 306.5805, 307.382, 308.1911, 309.0078, 309.8322, 310.6642, 
    311.5041, 312.3516, 313.207, 314.0701, 314.941, 315.8197, 316.7061, 
    317.6002, 318.502, 319.4114, 320.3284, 321.2528, 322.1847, 323.1238, 
    324.0701, 325.0234, 325.9837, 326.9507, 327.9243, 328.9044, 329.8907, 
    330.883, 331.8811, 332.8849, 333.8939, 334.9081, 335.927, 336.9506, 
    337.9783, 339.0101, 340.0455, 341.0842, 342.1259, 343.1703, 344.2171, 
    345.2658, 346.3161, 347.3678, 348.4203, 349.4734, 350.5266, 351.5797, 
    352.6322, 353.6839, 354.7342, 355.7829, 356.8297, 357.8741, 358.9158, 
    359.9545, 0.989933, 2.021674, 3.049454, 4.072974, 5.091947, 6.106095, 
    7.115152, 8.118866, 9.116993, 10.10931, 11.09559, 12.07564, 13.04927, 
    14.01629, 14.97656, 15.9299, 16.8762, 17.81532, 18.74715, 19.67159, 
    20.58856, 21.49797, 22.39977, 23.2939, 24.18031, 25.05898, 25.92989, 
    26.79302, 27.64837, 28.49594, 29.33576, 30.16784, 30.99221, 31.80891, 
    32.61798, 33.41949, 34.21347, 35 ;

 grid_latt =
  -35.63342, -36.0016, -36.36466, -36.72248, -37.07492, -37.42188, -37.76321, 
    -38.09881, -38.42853, -38.75225, -39.06984, -39.38117, -39.68611, 
    -39.98453, -40.27629, -40.56128, -40.83934, -41.11036, -41.37419, 
    -41.63073, -41.87982, -42.12135, -42.35519, -42.58122, -42.7993, 
    -43.00933, -43.21118, -43.40474, -43.58989, -43.76653, -43.93454, 
    -44.09382, -44.24429, -44.38583, -44.51836, -44.64181, -44.75608, 
    -44.8611, -44.9568, -45.04311, -45.11999, -45.18737, -45.24522, 
    -45.29348, -45.33213, -45.36115, -45.3805, -45.39018, -45.39018, 
    -45.3805, -45.36115, -45.33213, -45.29348, -45.24522, -45.18737, 
    -45.11999, -45.04311, -44.9568, -44.8611, -44.75608, -44.64181, 
    -44.51836, -44.38583, -44.24429, -44.09382, -43.93454, -43.76653, 
    -43.58989, -43.40474, -43.21118, -43.00933, -42.7993, -42.58122, 
    -42.35519, -42.12135, -41.87982, -41.63073, -41.37419, -41.11036, 
    -40.83934, -40.56128, -40.27629, -39.98453, -39.68611, -39.38117, 
    -39.06984, -38.75225, -38.42853, -38.09881, -37.76321, -37.42188, 
    -37.07492, -36.72248, -36.36466, -36.0016, -35.63342,
  -36.0016, -36.38164, -36.75665, -37.12651, -37.49107, -37.8502, -38.20377, 
    -38.55162, -38.89363, -39.22964, -39.55952, -39.88312, -40.20029, 
    -40.51088, -40.81476, -41.11176, -41.40174, -41.68456, -41.96006, 
    -42.2281, -42.48852, -42.74119, -42.98596, -43.22269, -43.45123, 
    -43.67144, -43.8832, -44.08636, -44.28079, -44.46637, -44.64297, 
    -44.81047, -44.96877, -45.11773, -45.25727, -45.38729, -45.50768, 
    -45.61835, -45.71924, -45.81026, -45.89135, -45.96243, -46.02346, 
    -46.07439, -46.11519, -46.14581, -46.16624, -46.17646, -46.17646, 
    -46.16624, -46.14581, -46.11519, -46.07439, -46.02346, -45.96243, 
    -45.89135, -45.81026, -45.71924, -45.61835, -45.50768, -45.38729, 
    -45.25727, -45.11773, -44.96877, -44.81047, -44.64297, -44.46637, 
    -44.28079, -44.08636, -43.8832, -43.67144, -43.45123, -43.22269, 
    -42.98596, -42.74119, -42.48852, -42.2281, -41.96006, -41.68456, 
    -41.40174, -41.11176, -40.81476, -40.51088, -40.20029, -39.88312, 
    -39.55952, -39.22964, -38.89363, -38.55162, -38.20377, -37.8502, 
    -37.49107, -37.12651, -36.75665, -36.38164, -36.0016,
  -36.36466, -36.75665, -37.14373, -37.52576, -37.90258, -38.27405, 
    -38.64002, -39.00033, -39.35483, -39.70337, -40.04577, -40.38189, 
    -40.71156, -41.03462, -41.35089, -41.66023, -41.96246, -42.2574, 
    -42.54491, -42.82481, -43.09693, -43.36111, -43.61718, -43.86499, 
    -44.10437, -44.33515, -44.55719, -44.77034, -44.97443, -45.16932, 
    -45.35488, -45.53096, -45.69742, -45.85415, -46.00101, -46.13791, 
    -46.26471, -46.38132, -46.48764, -46.5836, -46.66909, -46.74407, 
    -46.80845, -46.86219, -46.90523, -46.93755, -46.95911, -46.96989, 
    -46.96989, -46.95911, -46.93755, -46.90523, -46.86219, -46.80845, 
    -46.74407, -46.66909, -46.5836, -46.48764, -46.38132, -46.26471, 
    -46.13791, -46.00101, -45.85415, -45.69742, -45.53096, -45.35488, 
    -45.16932, -44.97443, -44.77034, -44.55719, -44.33515, -44.10437, 
    -43.86499, -43.61718, -43.36111, -43.09693, -42.82481, -42.54491, 
    -42.2574, -41.96246, -41.66023, -41.35089, -41.03462, -40.71156, 
    -40.38189, -40.04577, -39.70337, -39.35483, -39.00033, -38.64002, 
    -38.27405, -37.90258, -37.52576, -37.14373, -36.75665, -36.36466,
  -36.72248, -37.12651, -37.52576, -37.92007, -38.30929, -38.69325, 
    -39.07178, -39.44474, -39.81194, -40.17321, -40.52837, -40.87727, 
    -41.2197, -41.5555, -41.88448, -42.20646, -42.52125, -42.82867, 
    -43.12852, -43.42064, -43.70482, -43.98088, -44.24864, -44.50792, 
    -44.75852, -45.00027, -45.23299, -45.45651, -45.67065, -45.87524, 
    -46.07014, -46.25516, -46.43016, -46.595, -46.74953, -46.89362, 
    -47.02713, -47.14996, -47.26199, -47.36312, -47.45325, -47.53231, 
    -47.6002, -47.65689, -47.7023, -47.7364, -47.75915, -47.77053, -47.77053, 
    -47.75915, -47.7364, -47.7023, -47.65689, -47.6002, -47.53231, -47.45325, 
    -47.36312, -47.26199, -47.14996, -47.02713, -46.89362, -46.74953, 
    -46.595, -46.43016, -46.25516, -46.07014, -45.87524, -45.67065, 
    -45.45651, -45.23299, -45.00027, -44.75852, -44.50792, -44.24864, 
    -43.98088, -43.70482, -43.42064, -43.12852, -42.82867, -42.52125, 
    -42.20646, -41.88448, -41.5555, -41.2197, -40.87727, -40.52837, 
    -40.17321, -39.81194, -39.44474, -39.07178, -38.69325, -38.30929, 
    -37.92007, -37.52576, -37.12651, -36.72248,
  -37.07492, -37.49107, -37.90258, -38.30929, -38.71102, -39.10761, 
    -39.49888, -39.88465, -40.26473, -40.63895, -41.00711, -41.36901, 
    -41.72447, -42.07329, -42.41526, -42.75019, -43.07787, -43.39809, 
    -43.71065, -44.01534, -44.31195, -44.60027, -44.88011, -45.15124, 
    -45.41347, -45.66659, -45.91039, -46.14469, -46.36929, -46.58398, 
    -46.7886, -46.98296, -47.16688, -47.34019, -47.50273, -47.65435, 
    -47.79491, -47.92425, -48.04226, -48.14882, -48.24382, -48.32716, 
    -48.39876, -48.45854, -48.50644, -48.54241, -48.56641, -48.57842, 
    -48.57842, -48.56641, -48.54241, -48.50644, -48.45854, -48.39876, 
    -48.32716, -48.24382, -48.14882, -48.04226, -47.92425, -47.79491, 
    -47.65435, -47.50273, -47.34019, -47.16688, -46.98296, -46.7886, 
    -46.58398, -46.36929, -46.14469, -45.91039, -45.66659, -45.41347, 
    -45.15124, -44.88011, -44.60027, -44.31195, -44.01534, -43.71065, 
    -43.39809, -43.07787, -42.75019, -42.41526, -42.07329, -41.72447, 
    -41.36901, -41.00711, -40.63895, -40.26473, -39.88465, -39.49888, 
    -39.10761, -38.71102, -38.30929, -37.90258, -37.49107, -37.07492,
  -37.42188, -37.8502, -38.27405, -38.69325, -39.10761, -39.51696, -39.9211, 
    -40.31985, -40.71301, -41.10036, -41.48173, -41.85689, -42.22562, 
    -42.58773, -42.94299, -43.29116, -43.63205, -43.9654, -44.29101, 
    -44.60864, -44.91806, -45.21903, -45.51133, -45.79473, -46.06899, 
    -46.33389, -46.5892, -46.83469, -47.07016, -47.29537, -47.51012, 
    -47.71421, -47.90744, -48.08961, -48.26053, -48.42004, -48.56796, 
    -48.70414, -48.82842, -48.94068, -49.04079, -49.12864, -49.20412, 
    -49.26716, -49.31768, -49.35562, -49.38094, -49.3936, -49.3936, 
    -49.38094, -49.35562, -49.31768, -49.26716, -49.20412, -49.12864, 
    -49.04079, -48.94068, -48.82842, -48.70414, -48.56796, -48.42004, 
    -48.26053, -48.08961, -47.90744, -47.71421, -47.51012, -47.29537, 
    -47.07016, -46.83469, -46.5892, -46.33389, -46.06899, -45.79473, 
    -45.51133, -45.21903, -44.91806, -44.60864, -44.29101, -43.9654, 
    -43.63205, -43.29116, -42.94299, -42.58773, -42.22562, -41.85689, 
    -41.48173, -41.10036, -40.71301, -40.31985, -39.9211, -39.51696, 
    -39.10761, -38.69325, -38.27405, -37.8502, -37.42188,
  -37.76321, -38.20377, -38.64002, -39.07178, -39.49888, -39.9211, -40.33826, 
    -40.75014, -41.15653, -41.55723, -41.95201, -42.34064, -42.7229, 
    -43.09856, -43.46738, -43.82911, -44.18351, -44.53034, -44.86935, 
    -45.20028, -45.52287, -45.83688, -46.14204, -46.43811, -46.72482, 
    -47.00192, -47.26916, -47.52629, -47.77305, -48.0092, -48.23452, 
    -48.44876, -48.6517, -48.84312, -49.02282, -49.19058, -49.34622, 
    -49.48956, -49.62043, -49.73867, -49.84415, -49.93674, -50.01631, 
    -50.08277, -50.13604, -50.17606, -50.20276, -50.21612, -50.21612, 
    -50.20276, -50.17606, -50.13604, -50.08277, -50.01631, -49.93674, 
    -49.84415, -49.73867, -49.62043, -49.48956, -49.34622, -49.19058, 
    -49.02282, -48.84312, -48.6517, -48.44876, -48.23452, -48.0092, 
    -47.77305, -47.52629, -47.26916, -47.00192, -46.72482, -46.43811, 
    -46.14204, -45.83688, -45.52287, -45.20028, -44.86935, -44.53034, 
    -44.18351, -43.82911, -43.46738, -43.09856, -42.7229, -42.34064, 
    -41.95201, -41.55723, -41.15653, -40.75014, -40.33826, -39.9211, 
    -39.49888, -39.07178, -38.64002, -38.20377, -37.76321,
  -38.09881, -38.55162, -39.00033, -39.44474, -39.88465, -40.31985, 
    -40.75014, -41.17529, -41.59509, -42.0093, -42.41769, -42.82002, 
    -43.21604, -43.60551, -43.98816, -44.36374, -44.73198, -45.0926, 
    -45.44535, -45.78994, -46.12609, -46.45353, -46.77196, -47.08112, 
    -47.3807, -47.67044, -47.95004, -48.21923, -48.47774, -48.72528, 
    -48.9616, -49.18642, -49.39951, -49.6006, -49.78946, -49.96586, 
    -50.12959, -50.28045, -50.41822, -50.54276, -50.65387, -50.75143, 
    -50.83531, -50.90538, -50.96155, -51.00375, -51.03191, -51.046, -51.046, 
    -51.03191, -51.00375, -50.96155, -50.90538, -50.83531, -50.75143, 
    -50.65387, -50.54276, -50.41822, -50.28045, -50.12959, -49.96586, 
    -49.78946, -49.6006, -49.39951, -49.18642, -48.9616, -48.72528, 
    -48.47774, -48.21923, -47.95004, -47.67044, -47.3807, -47.08112, 
    -46.77196, -46.45353, -46.12609, -45.78994, -45.44535, -45.0926, 
    -44.73198, -44.36374, -43.98816, -43.60551, -43.21604, -42.82002, 
    -42.41769, -42.0093, -41.59509, -41.17529, -40.75014, -40.31985, 
    -39.88465, -39.44474, -39.00033, -38.55162, -38.09881,
  -38.42853, -38.89363, -39.35483, -39.81194, -40.26473, -40.71301, 
    -41.15653, -41.59509, -42.02843, -42.45632, -42.87851, -43.29474, 
    -43.70475, -44.10828, -44.50503, -44.89474, -45.27712, -45.65187, 
    -46.0187, -46.37732, -46.72741, -47.06866, -47.40077, -47.72343, 
    -48.03632, -48.33913, -48.63155, -48.91327, -49.18397, -49.44336, 
    -49.69113, -49.927, -50.15067, -50.36186, -50.56031, -50.74577, 
    -50.91797, -51.0767, -51.22174, -51.35287, -51.46992, -51.57272, 
    -51.66111, -51.73498, -51.7942, -51.8387, -51.8684, -51.88326, -51.88326, 
    -51.8684, -51.8387, -51.7942, -51.73498, -51.66111, -51.57272, -51.46992, 
    -51.35287, -51.22174, -51.0767, -50.91797, -50.74577, -50.56031, 
    -50.36186, -50.15067, -49.927, -49.69113, -49.44336, -49.18397, 
    -48.91327, -48.63155, -48.33913, -48.03632, -47.72343, -47.40077, 
    -47.06866, -46.72741, -46.37732, -46.0187, -45.65187, -45.27712, 
    -44.89474, -44.50503, -44.10828, -43.70475, -43.29474, -42.87851, 
    -42.45632, -42.02843, -41.59509, -41.15653, -40.71301, -40.26473, 
    -39.81194, -39.35483, -38.89363, -38.42853,
  -38.75225, -39.22964, -39.70337, -40.17321, -40.63895, -41.10036, 
    -41.55723, -42.0093, -42.45632, -42.89805, -43.33421, -43.76454, 
    -44.18875, -44.60656, -45.01768, -45.4218, -45.81862, -46.20782, 
    -46.58908, -46.96207, -47.32647, -47.68195, -48.02814, -48.36473, 
    -48.69137, -49.00771, -49.3134, -49.6081, -49.89148, -50.16318, 
    -50.42288, -50.67025, -50.90497, -51.12672, -51.33521, -51.53014, 
    -51.71123, -51.87823, -52.03088, -52.16895, -52.29223, -52.40054, 
    -52.4937, -52.57156, -52.63401, -52.68093, -52.71225, -52.72793, 
    -52.72793, -52.71225, -52.68093, -52.63401, -52.57156, -52.4937, 
    -52.40054, -52.29223, -52.16895, -52.03088, -51.87823, -51.71123, 
    -51.53014, -51.33521, -51.12672, -50.90497, -50.67025, -50.42288, 
    -50.16318, -49.89148, -49.6081, -49.3134, -49.00771, -48.69137, 
    -48.36473, -48.02814, -47.68195, -47.32647, -46.96207, -46.58908, 
    -46.20782, -45.81862, -45.4218, -45.01768, -44.60656, -44.18875, 
    -43.76454, -43.33421, -42.89805, -42.45632, -42.0093, -41.55723, 
    -41.10036, -40.63895, -40.17321, -39.70337, -39.22964, -38.75225,
  -39.06984, -39.55952, -40.04577, -40.52837, -41.00711, -41.48173, 
    -41.95201, -42.41769, -42.87851, -43.33421, -43.7845, -44.22911, 
    -44.66773, -45.10006, -45.52579, -45.94459, -46.35614, -46.76009, 
    -47.15612, -47.54385, -47.92294, -48.29302, -48.65372, -49.00467, 
    -49.3455, -49.67582, -49.99525, -50.30342, -50.59995, -50.88446, 
    -51.15658, -51.41594, -51.66219, -51.89498, -52.11396, -52.31881, 
    -52.50922, -52.68489, -52.84554, -52.99091, -53.12075, -53.23486, 
    -53.33304, -53.41512, -53.48095, -53.53043, -53.56347, -53.58, -53.58, 
    -53.56347, -53.53043, -53.48095, -53.41512, -53.33304, -53.23486, 
    -53.12075, -52.99091, -52.84554, -52.68489, -52.50922, -52.31881, 
    -52.11396, -51.89498, -51.66219, -51.41594, -51.15658, -50.88446, 
    -50.59995, -50.30342, -49.99525, -49.67582, -49.3455, -49.00467, 
    -48.65372, -48.29302, -47.92294, -47.54385, -47.15612, -46.76009, 
    -46.35614, -45.94459, -45.52579, -45.10006, -44.66773, -44.22911, 
    -43.7845, -43.33421, -42.87851, -42.41769, -41.95201, -41.48173, 
    -41.00711, -40.52837, -40.04577, -39.55952, -39.06984,
  -39.38117, -39.88312, -40.38189, -40.87727, -41.36901, -41.85689, 
    -42.34064, -42.82002, -43.29474, -43.76454, -44.22911, -44.68816, 
    -45.14137, -45.58843, -46.029, -46.46275, -46.88931, -47.30833, 
    -47.71944, -48.12227, -48.51642, -48.9015, -49.27712, -49.64286, 
    -49.99833, -50.34309, -50.67675, -50.99888, -51.30906, -51.60688, 
    -51.89192, -52.16379, -52.42207, -52.66639, -52.89635, -53.1116, 
    -53.31178, -53.49655, -53.6656, -53.81864, -53.95539, -54.07561, 
    -54.17908, -54.26561, -54.33502, -54.3872, -54.42204, -54.43948, 
    -54.43948, -54.42204, -54.3872, -54.33502, -54.26561, -54.17908, 
    -54.07561, -53.95539, -53.81864, -53.6656, -53.49655, -53.31178, 
    -53.1116, -52.89635, -52.66639, -52.42207, -52.16379, -51.89192, 
    -51.60688, -51.30906, -50.99888, -50.67675, -50.34309, -49.99833, 
    -49.64286, -49.27712, -48.9015, -48.51642, -48.12227, -47.71944, 
    -47.30833, -46.88931, -46.46275, -46.029, -45.58843, -45.14137, 
    -44.68816, -44.22911, -43.76454, -43.29474, -42.82002, -42.34064, 
    -41.85689, -41.36901, -40.87727, -40.38189, -39.88312, -39.38117,
  -39.68611, -40.20029, -40.71156, -41.2197, -41.72447, -42.22562, -42.7229, 
    -43.21604, -43.70475, -44.18875, -44.66773, -45.14137, -45.60936, 
    -46.07135, -46.52699, -46.97591, -47.41776, -47.85214, -48.27867, 
    -48.69693, -49.10651, -49.50698, -49.89793, -50.2789, -50.64946, 
    -51.00915, -51.35751, -51.6941, -52.01844, -52.33009, -52.62858, 
    -52.91348, -53.18432, -53.44069, -53.68214, -53.90828, -54.1187, 
    -54.31304, -54.49093, -54.65204, -54.79607, -54.92273, -55.03177, 
    -55.12299, -55.19618, -55.25121, -55.28796, -55.30635, -55.30635, 
    -55.28796, -55.25121, -55.19618, -55.12299, -55.03177, -54.92273, 
    -54.79607, -54.65204, -54.49093, -54.31304, -54.1187, -53.90828, 
    -53.68214, -53.44069, -53.18432, -52.91348, -52.62858, -52.33009, 
    -52.01844, -51.6941, -51.35751, -51.00915, -50.64946, -50.2789, 
    -49.89793, -49.50698, -49.10651, -48.69693, -48.27867, -47.85214, 
    -47.41776, -46.97591, -46.52699, -46.07135, -45.60936, -45.14137, 
    -44.66773, -44.18875, -43.70475, -43.21604, -42.7229, -42.22562, 
    -41.72447, -41.2197, -40.71156, -40.20029, -39.68611,
  -39.98453, -40.51088, -41.03462, -41.5555, -42.07329, -42.58773, -43.09856, 
    -43.60551, -44.10828, -44.60656, -45.10006, -45.58843, -46.07135, 
    -46.54844, -47.01936, -47.4837, -47.94109, -48.39112, -48.83337, 
    -49.2674, -49.69277, -50.10903, -50.51572, -50.91235, -51.29846, 
    -51.67355, -52.03711, -52.38867, -52.7277, -53.05371, -53.3662, 
    -53.66467, -53.94862, -54.21758, -54.47105, -54.70861, -54.92978, 
    -55.13416, -55.32135, -55.49096, -55.64265, -55.7761, -55.89104, 
    -55.9872, -56.06439, -56.12244, -56.1612, -56.18061, -56.18061, -56.1612, 
    -56.12244, -56.06439, -55.9872, -55.89104, -55.7761, -55.64265, 
    -55.49096, -55.32135, -55.13416, -54.92978, -54.70861, -54.47105, 
    -54.21758, -53.94862, -53.66467, -53.3662, -53.05371, -52.7277, 
    -52.38867, -52.03711, -51.67355, -51.29846, -50.91235, -50.51572, 
    -50.10903, -49.69277, -49.2674, -48.83337, -48.39112, -47.94109, 
    -47.4837, -47.01936, -46.54844, -46.07135, -45.58843, -45.10006, 
    -44.60656, -44.10828, -43.60551, -43.09856, -42.58773, -42.07329, 
    -41.5555, -41.03462, -40.51088, -39.98453,
  -40.27629, -40.81476, -41.35089, -41.88448, -42.41526, -42.94299, 
    -43.46738, -43.98816, -44.50503, -45.01768, -45.52579, -46.029, 
    -46.52699, -47.01936, -47.50573, -47.98571, -48.45889, -48.92484, 
    -49.3831, -49.83323, -50.27475, -50.70718, -51.13002, -51.54275, 
    -51.94487, -52.33583, -52.7151, -53.08215, -53.43641, -53.77734, 
    -54.10438, -54.41699, -54.71461, -54.99673, -55.2628, -55.51231, 
    -55.74477, -55.95971, -56.15667, -56.33524, -56.49501, -56.63563, 
    -56.75679, -56.85819, -56.93961, -57.00084, -57.04174, -57.06222, 
    -57.06222, -57.04174, -57.00084, -56.93961, -56.85819, -56.75679, 
    -56.63563, -56.49501, -56.33524, -56.15667, -55.95971, -55.74477, 
    -55.51231, -55.2628, -54.99673, -54.71461, -54.41699, -54.10438, 
    -53.77734, -53.43641, -53.08215, -52.7151, -52.33583, -51.94487, 
    -51.54275, -51.13002, -50.70718, -50.27475, -49.83323, -49.3831, 
    -48.92484, -48.45889, -47.98571, -47.50573, -47.01936, -46.52699, 
    -46.029, -45.52579, -45.01768, -44.50503, -43.98816, -43.46738, 
    -42.94299, -42.41526, -41.88448, -41.35089, -40.81476, -40.27629,
  -40.56128, -41.11176, -41.66023, -42.20646, -42.75019, -43.29116, 
    -43.82911, -44.36374, -44.89474, -45.4218, -45.94459, -46.46275, 
    -46.97591, -47.4837, -47.98571, -48.48154, -48.97073, -49.45285, 
    -49.92742, -50.39396, -50.85197, -51.30094, -51.74033, -52.16959, 
    -52.58817, -52.9955, -53.39099, -53.77406, -54.14409, -54.5005, 
    -54.84268, -55.17002, -55.48191, -55.77778, -56.05703, -56.31908, 
    -56.56339, -56.78943, -56.99669, -57.18469, -57.35299, -57.50119, 
    -57.62892, -57.73586, -57.82175, -57.88636, -57.92953, -57.95115, 
    -57.95115, -57.92953, -57.88636, -57.82175, -57.73586, -57.62892, 
    -57.50119, -57.35299, -57.18469, -56.99669, -56.78943, -56.56339, 
    -56.31908, -56.05703, -55.77778, -55.48191, -55.17002, -54.84268, 
    -54.5005, -54.14409, -53.77406, -53.39099, -52.9955, -52.58817, 
    -52.16959, -51.74033, -51.30094, -50.85197, -50.39396, -49.92742, 
    -49.45285, -48.97073, -48.48154, -47.98571, -47.4837, -46.97591, 
    -46.46275, -45.94459, -45.4218, -44.89474, -44.36374, -43.82911, 
    -43.29116, -42.75019, -42.20646, -41.66023, -41.11176, -40.56128,
  -40.83934, -41.40174, -41.96246, -42.52125, -43.07787, -43.63205, 
    -44.18351, -44.73198, -45.27712, -45.81862, -46.35614, -46.88931, 
    -47.41776, -47.94109, -48.45889, -48.97073, -49.47615, -49.97467, 
    -50.46582, -50.94908, -51.42391, -51.88978, -52.34612, -52.79234, 
    -53.22784, -53.65202, -54.06424, -54.46386, -54.85024, -55.22271, 
    -55.58062, -55.9233, -56.25008, -56.56032, -56.85336, -57.12857, 
    -57.38533, -57.62305, -57.84115, -58.0391, -58.21642, -58.37262, 
    -58.50731, -58.62013, -58.71076, -58.77895, -58.82452, -58.84734, 
    -58.84734, -58.82452, -58.77895, -58.71076, -58.62013, -58.50731, 
    -58.37262, -58.21642, -58.0391, -57.84115, -57.62305, -57.38533, 
    -57.12857, -56.85336, -56.56032, -56.25008, -55.9233, -55.58062, 
    -55.22271, -54.85024, -54.46386, -54.06424, -53.65202, -53.22784, 
    -52.79234, -52.34612, -51.88978, -51.42391, -50.94908, -50.46582, 
    -49.97467, -49.47615, -48.97073, -48.45889, -47.94109, -47.41776, 
    -46.88931, -46.35614, -45.81862, -45.27712, -44.73198, -44.18351, 
    -43.63205, -43.07787, -42.52125, -41.96246, -41.40174, -40.83934,
  -41.11036, -41.68456, -42.2574, -42.82867, -43.39809, -43.9654, -44.53034, 
    -45.0926, -45.65187, -46.20782, -46.76009, -47.30833, -47.85214, 
    -48.39112, -48.92484, -49.45285, -49.97467, -50.48983, -50.9978, 
    -51.49806, -51.99004, -52.47316, -52.94683, -53.41042, -53.8633, 
    -54.30482, -54.73428, -55.15101, -55.55429, -55.94343, -56.31768, 
    -56.67633, -57.01865, -57.34391, -57.65139, -57.9404, -58.21024, 
    -58.46024, -58.68978, -58.89825, -59.08508, -59.24976, -59.39183, 
    -59.51086, -59.60653, -59.67853, -59.72665, -59.75075, -59.75075, 
    -59.72665, -59.67853, -59.60653, -59.51086, -59.39183, -59.24976, 
    -59.08508, -58.89825, -58.68978, -58.46024, -58.21024, -57.9404, 
    -57.65139, -57.34391, -57.01865, -56.67633, -56.31768, -55.94343, 
    -55.55429, -55.15101, -54.73428, -54.30482, -53.8633, -53.41042, 
    -52.94683, -52.47316, -51.99004, -51.49806, -50.9978, -50.48983, 
    -49.97467, -49.45285, -48.92484, -48.39112, -47.85214, -47.30833, 
    -46.76009, -46.20782, -45.65187, -45.0926, -44.53034, -43.9654, 
    -43.39809, -42.82867, -42.2574, -41.68456, -41.11036,
  -41.37419, -41.96006, -42.54491, -43.12852, -43.71065, -44.29101, 
    -44.86935, -45.44535, -46.0187, -46.58908, -47.15612, -47.71944, 
    -48.27867, -48.83337, -49.3831, -49.92742, -50.46582, -50.9978, 
    -51.52283, -52.04035, -52.54977, -53.05048, -53.54185, -54.02324, 
    -54.49394, -54.95327, -55.40049, -55.83487, -56.25565, -56.66205, 
    -57.05328, -57.42855, -57.78707, -58.12803, -58.45065, -58.75413, 
    -59.03772, -59.30067, -59.54227, -59.76184, -59.95875, -60.13241, 
    -60.2823, -60.40795, -60.50896, -60.58501, -60.63584, -60.6613, -60.6613, 
    -60.63584, -60.58501, -60.50896, -60.40795, -60.2823, -60.13241, 
    -59.95875, -59.76184, -59.54227, -59.30067, -59.03772, -58.75413, 
    -58.45065, -58.12803, -57.78707, -57.42855, -57.05328, -56.66205, 
    -56.25565, -55.83487, -55.40049, -54.95327, -54.49394, -54.02324, 
    -53.54185, -53.05048, -52.54977, -52.04035, -51.52283, -50.9978, 
    -50.46582, -49.92742, -49.3831, -48.83337, -48.27867, -47.71944, 
    -47.15612, -46.58908, -46.0187, -45.44535, -44.86935, -44.29101, 
    -43.71065, -43.12852, -42.54491, -41.96006, -41.37419,
  -41.63073, -42.2281, -42.82481, -43.42064, -44.01534, -44.60864, -45.20028, 
    -45.78994, -46.37732, -46.96207, -47.54385, -48.12227, -48.69693, 
    -49.2674, -49.83323, -50.39396, -50.94908, -51.49806, -52.04035, 
    -52.57537, -53.10251, -53.62113, -54.13057, -54.63013, -55.11909, 
    -55.59671, -56.06221, -56.51479, -56.95364, -57.37793, -57.78679, 
    -58.17936, -58.55478, -58.91215, -59.25061, -59.56929, -59.86734, 
    -60.14393, -60.39826, -60.62958, -60.83716, -61.02035, -61.17855, 
    -61.31122, -61.41792, -61.49828, -61.55201, -61.57893, -61.57893, 
    -61.55201, -61.49828, -61.41792, -61.31122, -61.17855, -61.02035, 
    -60.83716, -60.62958, -60.39826, -60.14393, -59.86734, -59.56929, 
    -59.25061, -58.91215, -58.55478, -58.17936, -57.78679, -57.37793, 
    -56.95364, -56.51479, -56.06221, -55.59671, -55.11909, -54.63013, 
    -54.13057, -53.62113, -53.10251, -52.57537, -52.04035, -51.49806, 
    -50.94908, -50.39396, -49.83323, -49.2674, -48.69693, -48.12227, 
    -47.54385, -46.96207, -46.37732, -45.78994, -45.20028, -44.60864, 
    -44.01534, -43.42064, -42.82481, -42.2281, -41.63073,
  -41.87982, -42.48852, -43.09693, -43.70482, -44.31195, -44.91806, 
    -45.52287, -46.12609, -46.72741, -47.32647, -47.92294, -48.51642, 
    -49.10651, -49.69277, -50.27475, -50.85197, -51.42391, -51.99004, 
    -52.54977, -53.10251, -53.64762, -54.18444, -54.71228, -55.2304, 
    -55.73805, -56.23442, -56.7187, -57.19004, -57.64757, -58.09037, 
    -58.51752, -58.92809, -59.32111, -59.69563, -60.05069, -60.38533, 
    -60.6986, -60.98957, -61.25736, -61.50111, -61.72001, -61.91332, 
    -62.08035, -62.22052, -62.33329, -62.41824, -62.47506, -62.50353, 
    -62.50353, -62.47506, -62.41824, -62.33329, -62.22052, -62.08035, 
    -61.91332, -61.72001, -61.50111, -61.25736, -60.98957, -60.6986, 
    -60.38533, -60.05069, -59.69563, -59.32111, -58.92809, -58.51752, 
    -58.09037, -57.64757, -57.19004, -56.7187, -56.23442, -55.73805, 
    -55.2304, -54.71228, -54.18444, -53.64762, -53.10251, -52.54977, 
    -51.99004, -51.42391, -50.85197, -50.27475, -49.69277, -49.10651, 
    -48.51642, -47.92294, -47.32647, -46.72741, -46.12609, -45.52287, 
    -44.91806, -44.31195, -43.70482, -43.09693, -42.48852, -41.87982,
  -42.12135, -42.74119, -43.36111, -43.98088, -44.60027, -45.21903, 
    -45.83688, -46.45353, -47.06866, -47.68195, -48.29302, -48.9015, 
    -49.50698, -50.10903, -50.70718, -51.30094, -51.88978, -52.47316, 
    -53.05048, -53.62113, -54.18444, -54.73974, -55.28629, -55.82333, 
    -56.35006, -56.86565, -57.36921, -57.85986, -58.33664, -58.79859, 
    -59.24471, -59.67398, -60.08537, -60.47782, -60.85027, -61.20166, 
    -61.53094, -61.8371, -62.11912, -62.37604, -62.60696, -62.81103, 
    -62.98748, -63.13563, -63.25488, -63.34475, -63.40488, -63.43501, 
    -63.43501, -63.40488, -63.34475, -63.25488, -63.13563, -62.98748, 
    -62.81103, -62.60696, -62.37604, -62.11912, -61.8371, -61.53094, 
    -61.20166, -60.85027, -60.47782, -60.08537, -59.67398, -59.24471, 
    -58.79859, -58.33664, -57.85986, -57.36921, -56.86565, -56.35006, 
    -55.82333, -55.28629, -54.73974, -54.18444, -53.62113, -53.05048, 
    -52.47316, -51.88978, -51.30094, -50.70718, -50.10903, -49.50698, 
    -48.9015, -48.29302, -47.68195, -47.06866, -46.45353, -45.83688, 
    -45.21903, -44.60027, -43.98088, -43.36111, -42.74119, -42.12135,
  -42.35519, -42.98596, -43.61718, -44.24864, -44.88011, -45.51133, 
    -46.14204, -46.77196, -47.40077, -48.02814, -48.65372, -49.27712, 
    -49.89793, -50.51572, -51.13002, -51.74033, -52.34612, -52.94683, 
    -53.54185, -54.13057, -54.71228, -55.28629, -55.85184, -56.40814, 
    -56.95434, -57.48957, -58.01291, -58.52339, -59.02002, -59.50176, 
    -59.96754, -60.41625, -60.84677, -61.25794, -61.64861, -62.0176, 
    -62.36376, -62.68594, -62.98302, -63.25393, -63.49763, -63.71317, 
    -63.89967, -64.05634, -64.18253, -64.27767, -64.34134, -64.37325, 
    -64.37325, -64.34134, -64.27767, -64.18253, -64.05634, -63.89967, 
    -63.71317, -63.49763, -63.25393, -62.98302, -62.68594, -62.36376, 
    -62.0176, -61.64861, -61.25794, -60.84677, -60.41625, -59.96754, 
    -59.50176, -59.02002, -58.52339, -58.01291, -57.48957, -56.95434, 
    -56.40814, -55.85184, -55.28629, -54.71228, -54.13057, -53.54185, 
    -52.94683, -52.34612, -51.74033, -51.13002, -50.51572, -49.89793, 
    -49.27712, -48.65372, -48.02814, -47.40077, -46.77196, -46.14204, 
    -45.51133, -44.88011, -44.24864, -43.61718, -42.98596, -42.35519,
  -42.58122, -43.22269, -43.86499, -44.50792, -45.15124, -45.79473, 
    -46.43811, -47.08112, -47.72343, -48.36473, -49.00467, -49.64286, 
    -50.2789, -50.91235, -51.54275, -52.16959, -52.79234, -53.41042, 
    -54.02324, -54.63013, -55.2304, -55.82333, -56.40814, -56.98399, 
    -57.55002, -58.1053, -58.64888, -59.17973, -59.6968, -60.19897, -60.6851, 
    -61.154, -61.60444, -62.03517, -62.44493, -62.83242, -63.19636, 
    -63.53547, -63.84851, -64.13426, -64.39157, -64.61935, -64.81659, 
    -64.98241, -65.11604, -65.21684, -65.28431, -65.31813, -65.31813, 
    -65.28431, -65.21684, -65.11604, -64.98241, -64.81659, -64.61935, 
    -64.39157, -64.13426, -63.84851, -63.53547, -63.19636, -62.83242, 
    -62.44493, -62.03517, -61.60444, -61.154, -60.6851, -60.19897, -59.6968, 
    -59.17973, -58.64888, -58.1053, -57.55002, -56.98399, -56.40814, 
    -55.82333, -55.2304, -54.63013, -54.02324, -53.41042, -52.79234, 
    -52.16959, -51.54275, -50.91235, -50.2789, -49.64286, -49.00467, 
    -48.36473, -47.72343, -47.08112, -46.43811, -45.79473, -45.15124, 
    -44.50792, -43.86499, -43.22269, -42.58122,
  -42.7993, -43.45123, -44.10437, -44.75852, -45.41347, -46.06899, -46.72482, 
    -47.3807, -48.03632, -48.69137, -49.3455, -49.99833, -50.64946, 
    -51.29846, -51.94487, -52.58817, -53.22784, -53.8633, -54.49394, 
    -55.11909, -55.73805, -56.35006, -56.95434, -57.55002, -58.1362, 
    -58.71193, -59.2762, -59.82792, -60.36599, -60.88923, -61.39641, 
    -61.88625, -62.35743, -62.80859, -63.23833, -63.64526, -64.02795, 
    -64.38497, -64.71494, -65.01648, -65.2883, -65.52915, -65.73791, 
    -65.91354, -66.05517, -66.16206, -66.23363, -66.26952, -66.26952, 
    -66.23363, -66.16206, -66.05517, -65.91354, -65.73791, -65.52915, 
    -65.2883, -65.01648, -64.71494, -64.38497, -64.02795, -63.64526, 
    -63.23833, -62.80859, -62.35743, -61.88625, -61.39641, -60.88923, 
    -60.36599, -59.82792, -59.2762, -58.71193, -58.1362, -57.55002, 
    -56.95434, -56.35006, -55.73805, -55.11909, -54.49394, -53.8633, 
    -53.22784, -52.58817, -51.94487, -51.29846, -50.64946, -49.99833, 
    -49.3455, -48.69137, -48.03632, -47.3807, -46.72482, -46.06899, 
    -45.41347, -44.75852, -44.10437, -43.45123, -42.7993,
  -43.00933, -43.67144, -44.33515, -45.00027, -45.66659, -46.33389, 
    -47.00192, -47.67044, -48.33913, -49.00771, -49.67582, -50.34309, 
    -51.00915, -51.67355, -52.33583, -52.9955, -53.65202, -54.30482, 
    -54.95327, -55.59671, -56.23442, -56.86565, -57.48957, -58.1053, 
    -58.71193, -59.30845, -59.89382, -60.4669, -61.02654, -61.57146, 
    -62.10038, -62.61193, -63.10468, -63.57715, -64.02785, -64.4552, 
    -64.85765, -65.23363, -65.58157, -65.89993, -66.18724, -66.44211, 
    -66.66322, -66.84942, -66.99967, -67.11313, -67.18914, -67.22726, 
    -67.22726, -67.18914, -67.11313, -66.99967, -66.84942, -66.66322, 
    -66.44211, -66.18724, -65.89993, -65.58157, -65.23363, -64.85765, 
    -64.4552, -64.02785, -63.57715, -63.10468, -62.61193, -62.10038, 
    -61.57146, -61.02654, -60.4669, -59.89382, -59.30845, -58.71193, 
    -58.1053, -57.48957, -56.86565, -56.23442, -55.59671, -54.95327, 
    -54.30482, -53.65202, -52.9955, -52.33583, -51.67355, -51.00915, 
    -50.34309, -49.67582, -49.00771, -48.33913, -47.67044, -47.00192, 
    -46.33389, -45.66659, -45.00027, -44.33515, -43.67144, -43.00933,
  -43.21118, -43.8832, -44.55719, -45.23299, -45.91039, -46.5892, -47.26916, 
    -47.95004, -48.63155, -49.3134, -49.99525, -50.67675, -51.35751, 
    -52.03711, -52.7151, -53.39099, -54.06424, -54.73428, -55.40049, 
    -56.06221, -56.7187, -57.36921, -58.01291, -58.64888, -59.2762, 
    -59.89382, -60.50066, -61.09555, -61.67727, -62.2445, -62.79585, 
    -63.32987, -63.84503, -64.33974, -64.81236, -65.26118, -65.68449, 
    -66.08053, -66.44756, -66.78387, -67.08776, -67.35767, -67.59209, 
    -67.78967, -67.94925, -68.06983, -68.15065, -68.19119, -68.19119, 
    -68.15065, -68.06983, -67.94925, -67.78967, -67.59209, -67.35767, 
    -67.08776, -66.78387, -66.44756, -66.08053, -65.68449, -65.26118, 
    -64.81236, -64.33974, -63.84503, -63.32987, -62.79585, -62.2445, 
    -61.67727, -61.09555, -60.50066, -59.89382, -59.2762, -58.64888, 
    -58.01291, -57.36921, -56.7187, -56.06221, -55.40049, -54.73428, 
    -54.06424, -53.39099, -52.7151, -52.03711, -51.35751, -50.67675, 
    -49.99525, -49.3134, -48.63155, -47.95004, -47.26916, -46.5892, 
    -45.91039, -45.23299, -44.55719, -43.8832, -43.21118,
  -43.40474, -44.08636, -44.77034, -45.45651, -46.14469, -46.83469, 
    -47.52629, -48.21923, -48.91327, -49.6081, -50.30342, -50.99888, 
    -51.6941, -52.38867, -53.08215, -53.77406, -54.46386, -55.15101, 
    -55.83487, -56.51479, -57.19004, -57.85986, -58.52339, -59.17973, 
    -59.82792, -60.4669, -61.09555, -61.71267, -62.31697, -62.90707, 
    -63.48152, -64.03877, -64.57719, -65.09508, -65.59063, -66.06201, 
    -66.50732, -66.92463, -67.31198, -67.66744, -67.98912, -68.2752, 
    -68.52398, -68.7339, -68.90359, -69.03191, -69.11797, -69.16115, 
    -69.16115, -69.11797, -69.03191, -68.90359, -68.7339, -68.52398, 
    -68.2752, -67.98912, -67.66744, -67.31198, -66.92463, -66.50732, 
    -66.06201, -65.59063, -65.09508, -64.57719, -64.03877, -63.48152, 
    -62.90707, -62.31697, -61.71267, -61.09555, -60.4669, -59.82792, 
    -59.17973, -58.52339, -57.85986, -57.19004, -56.51479, -55.83487, 
    -55.15101, -54.46386, -53.77406, -53.08215, -52.38867, -51.6941, 
    -50.99888, -50.30342, -49.6081, -48.91327, -48.21923, -47.52629, 
    -46.83469, -46.14469, -45.45651, -44.77034, -44.08636, -43.40474,
  -43.58989, -44.28079, -44.97443, -45.67065, -46.36929, -47.07016, 
    -47.77305, -48.47774, -49.18397, -49.89148, -50.59995, -51.30906, 
    -52.01844, -52.7277, -53.43641, -54.14409, -54.85024, -55.55429, 
    -56.25565, -56.95364, -57.64757, -58.33664, -59.02002, -59.6968, 
    -60.36599, -61.02654, -61.67727, -62.31697, -62.94429, -63.55782, 
    -64.15601, -64.73723, -65.29976, -65.84176, -66.36131, -66.85638, 
    -67.32491, -67.76476, -68.17374, -68.54969, -68.89046, -69.19399, 
    -69.45831, -69.68162, -69.86233, -69.99909, -70.09087, -70.13693, 
    -70.13693, -70.09087, -69.99909, -69.86233, -69.68162, -69.45831, 
    -69.19399, -68.89046, -68.54969, -68.17374, -67.76476, -67.32491, 
    -66.85638, -66.36131, -65.84176, -65.29976, -64.73723, -64.15601, 
    -63.55782, -62.94429, -62.31697, -61.67727, -61.02654, -60.36599, 
    -59.6968, -59.02002, -58.33664, -57.64757, -56.95364, -56.25565, 
    -55.55429, -54.85024, -54.14409, -53.43641, -52.7277, -52.01844, 
    -51.30906, -50.59995, -49.89148, -49.18397, -48.47774, -47.77305, 
    -47.07016, -46.36929, -45.67065, -44.97443, -44.28079, -43.58989,
  -43.76653, -44.46637, -45.16932, -45.87524, -46.58398, -47.29537, -48.0092, 
    -48.72528, -49.44336, -50.16318, -50.88446, -51.60688, -52.33009, 
    -53.05371, -53.77734, -54.5005, -55.22271, -55.94343, -56.66205, 
    -57.37793, -58.09037, -58.79859, -59.50176, -60.19897, -60.88923, 
    -61.57146, -62.2445, -62.90707, -63.55782, -64.19525, -64.81778, 
    -65.42369, -66.01116, -66.57823, -67.12283, -67.64278, -68.13581, 
    -68.59956, -69.03159, -69.4295, -69.79082, -70.1132, -70.39439, 
    -70.63229, -70.82504, -70.97105, -71.06911, -71.11835, -71.11835, 
    -71.06911, -70.97105, -70.82504, -70.63229, -70.39439, -70.1132, 
    -69.79082, -69.4295, -69.03159, -68.59956, -68.13581, -67.64278, 
    -67.12283, -66.57823, -66.01116, -65.42369, -64.81778, -64.19525, 
    -63.55782, -62.90707, -62.2445, -61.57146, -60.88923, -60.19897, 
    -59.50176, -58.79859, -58.09037, -57.37793, -56.66205, -55.94343, 
    -55.22271, -54.5005, -53.77734, -53.05371, -52.33009, -51.60688, 
    -50.88446, -50.16318, -49.44336, -48.72528, -48.0092, -47.29537, 
    -46.58398, -45.87524, -45.16932, -44.46637, -43.76653,
  -43.93454, -44.64297, -45.35488, -46.07014, -46.7886, -47.51012, -48.23452, 
    -48.9616, -49.69113, -50.42288, -51.15658, -51.89192, -52.62858, 
    -53.3662, -54.10438, -54.84268, -55.58062, -56.31768, -57.05328, 
    -57.78679, -58.51752, -59.24471, -59.96754, -60.6851, -61.39641, 
    -62.10038, -62.79585, -63.48152, -64.15601, -64.81778, -65.46519, 
    -66.09647, -66.70969, -67.30276, -67.8735, -68.41954, -68.9384, 
    -69.42749, -69.88412, -70.30556, -70.68905, -71.03188, -71.33143, 
    -71.58528, -71.79124, -71.94746, -72.05244, -72.10519, -72.10519, 
    -72.05244, -71.94746, -71.79124, -71.58528, -71.33143, -71.03188, 
    -70.68905, -70.30556, -69.88412, -69.42749, -68.9384, -68.41954, 
    -67.8735, -67.30276, -66.70969, -66.09647, -65.46519, -64.81778, 
    -64.15601, -63.48152, -62.79585, -62.10038, -61.39641, -60.6851, 
    -59.96754, -59.24471, -58.51752, -57.78679, -57.05328, -56.31768, 
    -55.58062, -54.84268, -54.10438, -53.3662, -52.62858, -51.89192, 
    -51.15658, -50.42288, -49.69113, -48.9616, -48.23452, -47.51012, 
    -46.7886, -46.07014, -45.35488, -44.64297, -43.93454,
  -44.09382, -44.81047, -45.53096, -46.25516, -46.98296, -47.71421, 
    -48.44876, -49.18642, -49.927, -50.67025, -51.41594, -52.16379, 
    -52.91348, -53.66467, -54.41699, -55.17002, -55.9233, -56.67633, 
    -57.42855, -58.17936, -58.92809, -59.67398, -60.41625, -61.154, 
    -61.88625, -62.61193, -63.32987, -64.03877, -64.73723, -65.42369, 
    -66.09647, -66.75372, -67.39344, -68.01344, -68.61138, -69.18474, 
    -69.73082, -70.24678, -70.72966, -71.17637, -71.5838, -71.94884, 
    -72.26848, -72.53986, -72.76041, -72.92789, -73.04058, -73.09724, 
    -73.09724, -73.04058, -72.92789, -72.76041, -72.53986, -72.26848, 
    -71.94884, -71.5838, -71.17637, -70.72966, -70.24678, -69.73082, 
    -69.18474, -68.61138, -68.01344, -67.39344, -66.75372, -66.09647, 
    -65.42369, -64.73723, -64.03877, -63.32987, -62.61193, -61.88625, 
    -61.154, -60.41625, -59.67398, -58.92809, -58.17936, -57.42855, 
    -56.67633, -55.9233, -55.17002, -54.41699, -53.66467, -52.91348, 
    -52.16379, -51.41594, -50.67025, -49.927, -49.18642, -48.44876, 
    -47.71421, -46.98296, -46.25516, -45.53096, -44.81047, -44.09382,
  -44.24429, -44.96877, -45.69742, -46.43016, -47.16688, -47.90744, -48.6517, 
    -49.39951, -50.15067, -50.90497, -51.66219, -52.42207, -53.18432, 
    -53.94862, -54.71461, -55.48191, -56.25008, -57.01865, -57.78707, 
    -58.55478, -59.32111, -60.08537, -60.84677, -61.60444, -62.35743, 
    -63.10468, -63.84503, -64.57719, -65.29976, -66.01116, -66.70969, 
    -67.39344, -68.06035, -68.70814, -69.33433, -69.93623, -70.51096, 
    -71.0554, -71.56628, -72.04017, -72.47352, -72.86278, -73.20444, 
    -73.49516, -73.73187, -73.91193, -74.03321, -74.09423, -74.09423, 
    -74.03321, -73.91193, -73.73187, -73.49516, -73.20444, -72.86278, 
    -72.47352, -72.04017, -71.56628, -71.0554, -70.51096, -69.93623, 
    -69.33433, -68.70814, -68.06035, -67.39344, -66.70969, -66.01116, 
    -65.29976, -64.57719, -63.84503, -63.10468, -62.35743, -61.60444, 
    -60.84677, -60.08537, -59.32111, -58.55478, -57.78707, -57.01865, 
    -56.25008, -55.48191, -54.71461, -53.94862, -53.18432, -52.42207, 
    -51.66219, -50.90497, -50.15067, -49.39951, -48.6517, -47.90744, 
    -47.16688, -46.43016, -45.69742, -44.96877, -44.24429,
  -44.38583, -45.11773, -45.85415, -46.595, -47.34019, -48.08961, -48.84312, 
    -49.6006, -50.36186, -51.12672, -51.89498, -52.66639, -53.44069, 
    -54.21758, -54.99673, -55.77778, -56.56032, -57.34391, -58.12803, 
    -58.91215, -59.69563, -60.47782, -61.25794, -62.03517, -62.80859, 
    -63.57715, -64.33974, -65.09508, -65.84176, -66.57823, -67.30276, 
    -68.01344, -68.70814, -69.38449, -70.03993, -70.67162, -71.27643, 
    -71.85101, -72.39178, -72.89487, -73.35633, -73.77206, -74.13797, 
    -74.45013, -74.70488, -74.89902, -75.02998, -75.09593, -75.09593, 
    -75.02998, -74.89902, -74.70488, -74.45013, -74.13797, -73.77206, 
    -73.35633, -72.89487, -72.39178, -71.85101, -71.27643, -70.67162, 
    -70.03993, -69.38449, -68.70814, -68.01344, -67.30276, -66.57823, 
    -65.84176, -65.09508, -64.33974, -63.57715, -62.80859, -62.03517, 
    -61.25794, -60.47782, -59.69563, -58.91215, -58.12803, -57.34391, 
    -56.56032, -55.77778, -54.99673, -54.21758, -53.44069, -52.66639, 
    -51.89498, -51.12672, -50.36186, -49.6006, -48.84312, -48.08961, 
    -47.34019, -46.595, -45.85415, -45.11773, -44.38583,
  -44.51836, -45.25727, -46.00101, -46.74953, -47.50273, -48.26053, 
    -49.02282, -49.78946, -50.56031, -51.33521, -52.11396, -52.89635, 
    -53.68214, -54.47105, -55.2628, -56.05703, -56.85336, -57.65139, 
    -58.45065, -59.25061, -60.05069, -60.85027, -61.64861, -62.44493, 
    -63.23833, -64.02785, -64.81236, -65.59063, -66.36131, -67.12283, 
    -67.8735, -68.61138, -69.33433, -70.03993, -70.72552, -71.38813, 
    -72.02446, -72.6309, -73.20351, -73.73804, -74.23001, -74.67474, 
    -75.06745, -75.40351, -75.67852, -75.88858, -76.03052, -76.10207, 
    -76.10207, -76.03052, -75.88858, -75.67852, -75.40351, -75.06745, 
    -74.67474, -74.23001, -73.73804, -73.20351, -72.6309, -72.02446, 
    -71.38813, -70.72552, -70.03993, -69.33433, -68.61138, -67.8735, 
    -67.12283, -66.36131, -65.59063, -64.81236, -64.02785, -63.23833, 
    -62.44493, -61.64861, -60.85027, -60.05069, -59.25061, -58.45065, 
    -57.65139, -56.85336, -56.05703, -55.2628, -54.47105, -53.68214, 
    -52.89635, -52.11396, -51.33521, -50.56031, -49.78946, -49.02282, 
    -48.26053, -47.50273, -46.74953, -46.00101, -45.25727, -44.51836,
  -44.64181, -45.38729, -46.13791, -46.89362, -47.65435, -48.42004, 
    -49.19058, -49.96586, -50.74577, -51.53014, -52.31881, -53.1116, 
    -53.90828, -54.70861, -55.51231, -56.31908, -57.12857, -57.9404, 
    -58.75413, -59.56929, -60.38533, -61.20166, -62.0176, -62.83242, 
    -63.64526, -64.4552, -65.26118, -66.06201, -66.85638, -67.64278, 
    -68.41954, -69.18474, -69.93623, -70.67162, -71.38813, -72.08273, 
    -72.75193, -73.39191, -73.99841, -74.56674, -75.09187, -75.56844, 
    -75.99091, -76.35376, -76.65166, -76.87985, -77.03436, -77.11236, 
    -77.11236, -77.03436, -76.87985, -76.65166, -76.35376, -75.99091, 
    -75.56844, -75.09187, -74.56674, -73.99841, -73.39191, -72.75193, 
    -72.08273, -71.38813, -70.67162, -69.93623, -69.18474, -68.41954, 
    -67.64278, -66.85638, -66.06201, -65.26118, -64.4552, -63.64526, 
    -62.83242, -62.0176, -61.20166, -60.38533, -59.56929, -58.75413, 
    -57.9404, -57.12857, -56.31908, -55.51231, -54.70861, -53.90828, 
    -53.1116, -52.31881, -51.53014, -50.74577, -49.96586, -49.19058, 
    -48.42004, -47.65435, -46.89362, -46.13791, -45.38729, -44.64181,
  -44.75608, -45.50768, -46.26471, -47.02713, -47.79491, -48.56796, 
    -49.34622, -50.12959, -50.91797, -51.71123, -52.50922, -53.31178, 
    -54.1187, -54.92978, -55.74477, -56.56339, -57.38533, -58.21024, 
    -59.03772, -59.86734, -60.6986, -61.53094, -62.36376, -63.19636, 
    -64.02795, -64.85765, -65.68449, -66.50732, -67.32491, -68.13581, 
    -68.9384, -69.73082, -70.51096, -71.27643, -72.02446, -72.75193, 
    -73.45528, -74.13045, -74.77289, -75.37749, -75.93864, -76.45026, 
    -76.90587, -77.2989, -77.62291, -77.87194, -78.04102, -78.1265, -78.1265, 
    -78.04102, -77.87194, -77.62291, -77.2989, -76.90587, -76.45026, 
    -75.93864, -75.37749, -74.77289, -74.13045, -73.45528, -72.75193, 
    -72.02446, -71.27643, -70.51096, -69.73082, -68.9384, -68.13581, 
    -67.32491, -66.50732, -65.68449, -64.85765, -64.02795, -63.19636, 
    -62.36376, -61.53094, -60.6986, -59.86734, -59.03772, -58.21024, 
    -57.38533, -56.56339, -55.74477, -54.92978, -54.1187, -53.31178, 
    -52.50922, -51.71123, -50.91797, -50.12959, -49.34622, -48.56796, 
    -47.79491, -47.02713, -46.26471, -45.50768, -44.75608,
  -44.8611, -45.61835, -46.38132, -47.14996, -47.92425, -48.70414, -49.48956, 
    -50.28045, -51.0767, -51.87823, -52.68489, -53.49655, -54.31304, 
    -55.13416, -55.95971, -56.78943, -57.62305, -58.46024, -59.30067, 
    -60.14393, -60.98957, -61.8371, -62.68594, -63.53547, -64.38497, 
    -65.23363, -66.08053, -66.92463, -67.76476, -68.59956, -69.42749, 
    -70.24678, -71.0554, -71.85101, -72.6309, -73.39191, -74.13045, 
    -74.84232, -75.5227, -76.16611, -76.76637, -77.31655, -77.8092, 
    -78.23647, -78.59045, -78.86371, -79.04986, -79.14419, -79.14419, 
    -79.04986, -78.86371, -78.59045, -78.23647, -77.8092, -77.31655, 
    -76.76637, -76.16611, -75.5227, -74.84232, -74.13045, -73.39191, 
    -72.6309, -71.85101, -71.0554, -70.24678, -69.42749, -68.59956, 
    -67.76476, -66.92463, -66.08053, -65.23363, -64.38497, -63.53547, 
    -62.68594, -61.8371, -60.98957, -60.14393, -59.30067, -58.46024, 
    -57.62305, -56.78943, -55.95971, -55.13416, -54.31304, -53.49655, 
    -52.68489, -51.87823, -51.0767, -50.28045, -49.48956, -48.70414, 
    -47.92425, -47.14996, -46.38132, -45.61835, -44.8611,
  -44.9568, -45.71924, -46.48764, -47.26199, -48.04226, -48.82842, -49.62043, 
    -50.41822, -51.22174, -52.03088, -52.84554, -53.6656, -54.49093, 
    -55.32135, -56.15667, -56.99669, -57.84115, -58.68978, -59.54227, 
    -60.39826, -61.25736, -62.11912, -62.98302, -63.84851, -64.71494, 
    -65.58157, -66.44756, -67.31198, -68.17374, -69.03159, -69.88412, 
    -70.72966, -71.56628, -72.39178, -73.20351, -73.99841, -74.77289, 
    -75.5227, -76.24287, -76.9276, -77.57013, -78.16277, -78.69691, 
    -79.16319, -79.55191, -79.85367, -80.06013, -80.16506, -80.16506, 
    -80.06013, -79.85367, -79.55191, -79.16319, -78.69691, -78.16277, 
    -77.57013, -76.9276, -76.24287, -75.5227, -74.77289, -73.99841, 
    -73.20351, -72.39178, -71.56628, -70.72966, -69.88412, -69.03159, 
    -68.17374, -67.31198, -66.44756, -65.58157, -64.71494, -63.84851, 
    -62.98302, -62.11912, -61.25736, -60.39826, -59.54227, -58.68978, 
    -57.84115, -56.99669, -56.15667, -55.32135, -54.49093, -53.6656, 
    -52.84554, -52.03088, -51.22174, -50.41822, -49.62043, -48.82842, 
    -48.04226, -47.26199, -46.48764, -45.71924, -44.9568,
  -45.04311, -45.81026, -46.5836, -47.36312, -48.14882, -48.94068, -49.73867, 
    -50.54276, -51.35287, -52.16895, -52.99091, -53.81864, -54.65204, 
    -55.49096, -56.33524, -57.18469, -58.0391, -58.89825, -59.76184, 
    -60.62958, -61.50111, -62.37604, -63.25393, -64.13426, -65.01648, 
    -65.89993, -66.78387, -67.66744, -68.54969, -69.4295, -70.30556, 
    -71.17637, -72.04017, -72.89487, -73.73804, -74.56674, -75.37749, 
    -76.16611, -76.9276, -77.65593, -78.34393, -78.98316, -79.56378, 
    -80.07474, -80.5041, -80.83981, -81.07088, -81.18875, -81.18875, 
    -81.07088, -80.83981, -80.5041, -80.07474, -79.56378, -78.98316, 
    -78.34393, -77.65593, -76.9276, -76.16611, -75.37749, -74.56674, 
    -73.73804, -72.89487, -72.04017, -71.17637, -70.30556, -69.4295, 
    -68.54969, -67.66744, -66.78387, -65.89993, -65.01648, -64.13426, 
    -63.25393, -62.37604, -61.50111, -60.62958, -59.76184, -58.89825, 
    -58.0391, -57.18469, -56.33524, -55.49096, -54.65204, -53.81864, 
    -52.99091, -52.16895, -51.35287, -50.54276, -49.73867, -48.94068, 
    -48.14882, -47.36312, -46.5836, -45.81026, -45.04311,
  -45.11999, -45.89135, -46.66909, -47.45325, -48.24382, -49.04079, 
    -49.84415, -50.65387, -51.46992, -52.29223, -53.12075, -53.95539, 
    -54.79607, -55.64265, -56.49501, -57.35299, -58.21642, -59.08508, 
    -59.95875, -60.83716, -61.72001, -62.60696, -63.49763, -64.39157, 
    -65.2883, -66.18724, -67.08776, -67.98912, -68.89046, -69.79082, 
    -70.68905, -71.5838, -72.47352, -73.35633, -74.23001, -75.09187, 
    -75.93864, -76.76637, -77.57013, -78.34393, -79.08037, -79.77036, 
    -80.40296, -80.96523, -81.44252, -81.81931, -82.08073, -82.21483, 
    -82.21483, -82.08073, -81.81931, -81.44252, -80.96523, -80.40296, 
    -79.77036, -79.08037, -78.34393, -77.57013, -76.76637, -75.93864, 
    -75.09187, -74.23001, -73.35633, -72.47352, -71.5838, -70.68905, 
    -69.79082, -68.89046, -67.98912, -67.08776, -66.18724, -65.2883, 
    -64.39157, -63.49763, -62.60696, -61.72001, -60.83716, -59.95875, 
    -59.08508, -58.21642, -57.35299, -56.49501, -55.64265, -54.79607, 
    -53.95539, -53.12075, -52.29223, -51.46992, -50.65387, -49.84415, 
    -49.04079, -48.24382, -47.45325, -46.66909, -45.89135, -45.11999,
  -45.18737, -45.96243, -46.74407, -47.53231, -48.32716, -49.12864, 
    -49.93674, -50.75143, -51.57272, -52.40054, -53.23486, -54.07561, 
    -54.92273, -55.7761, -56.63563, -57.50119, -58.37262, -59.24976, 
    -60.13241, -61.02035, -61.91332, -62.81103, -63.71317, -64.61935, 
    -65.52915, -66.44211, -67.35767, -68.2752, -69.19399, -70.1132, 
    -71.03188, -71.94884, -72.86278, -73.77206, -74.67474, -75.56844, 
    -76.45026, -77.31655, -78.16277, -78.98316, -79.77036, -80.51504, 
    -81.20532, -81.82646, -82.3607, -82.78796, -83.08778, -83.24277, 
    -83.24277, -83.08778, -82.78796, -82.3607, -81.82646, -81.20532, 
    -80.51504, -79.77036, -78.98316, -78.16277, -77.31655, -76.45026, 
    -75.56844, -74.67474, -73.77206, -72.86278, -71.94884, -71.03188, 
    -70.1132, -69.19399, -68.2752, -67.35767, -66.44211, -65.52915, 
    -64.61935, -63.71317, -62.81103, -61.91332, -61.02035, -60.13241, 
    -59.24976, -58.37262, -57.50119, -56.63563, -55.7761, -54.92273, 
    -54.07561, -53.23486, -52.40054, -51.57272, -50.75143, -49.93674, 
    -49.12864, -48.32716, -47.53231, -46.74407, -45.96243, -45.18737,
  -45.24522, -46.02346, -46.80845, -47.6002, -48.39876, -49.20412, -50.01631, 
    -50.83531, -51.66111, -52.4937, -53.33304, -54.17908, -55.03177, 
    -55.89104, -56.75679, -57.62892, -58.50731, -59.39183, -60.2823, 
    -61.17855, -62.08035, -62.98748, -63.89967, -64.81659, -65.73791, 
    -66.66322, -67.59209, -68.52398, -69.45831, -70.39439, -71.33143, 
    -72.26848, -73.20444, -74.13797, -75.06745, -75.99091, -76.90587, 
    -77.8092, -78.69691, -79.56378, -80.40296, -81.20532, -81.95869, 
    -82.6469, -83.249, -83.73922, -84.08896, -84.27195, -84.27195, -84.08896, 
    -83.73922, -83.249, -82.6469, -81.95869, -81.20532, -80.40296, -79.56378, 
    -78.69691, -77.8092, -76.90587, -75.99091, -75.06745, -74.13797, 
    -73.20444, -72.26848, -71.33143, -70.39439, -69.45831, -68.52398, 
    -67.59209, -66.66322, -65.73791, -64.81659, -63.89967, -62.98748, 
    -62.08035, -61.17855, -60.2823, -59.39183, -58.50731, -57.62892, 
    -56.75679, -55.89104, -55.03177, -54.17908, -53.33304, -52.4937, 
    -51.66111, -50.83531, -50.01631, -49.20412, -48.39876, -47.6002, 
    -46.80845, -46.02346, -45.24522,
  -45.29348, -46.07439, -46.86219, -47.65689, -48.45854, -49.26716, 
    -50.08277, -50.90538, -51.73498, -52.57156, -53.41512, -54.26561, 
    -55.12299, -55.9872, -56.85819, -57.73586, -58.62013, -59.51086, 
    -60.40795, -61.31122, -62.22052, -63.13563, -64.05634, -64.98241, 
    -65.91354, -66.84942, -67.78967, -68.7339, -69.68162, -70.63229, 
    -71.58528, -72.53986, -73.49516, -74.45013, -75.40351, -76.35376, 
    -77.2989, -78.23647, -79.16319, -80.07474, -80.96523, -81.82646, 
    -82.6469, -83.41006, -84.09252, -84.66222, -85.079, -85.30138, -85.30138, 
    -85.079, -84.66222, -84.09252, -83.41006, -82.6469, -81.82646, -80.96523, 
    -80.07474, -79.16319, -78.23647, -77.2989, -76.35376, -75.40351, 
    -74.45013, -73.49516, -72.53986, -71.58528, -70.63229, -69.68162, 
    -68.7339, -67.78967, -66.84942, -65.91354, -64.98241, -64.05634, 
    -63.13563, -62.22052, -61.31122, -60.40795, -59.51086, -58.62013, 
    -57.73586, -56.85819, -55.9872, -55.12299, -54.26561, -53.41512, 
    -52.57156, -51.73498, -50.90538, -50.08277, -49.26716, -48.45854, 
    -47.65689, -46.86219, -46.07439, -45.29348,
  -45.33213, -46.11519, -46.90523, -47.7023, -48.50644, -49.31768, -50.13604, 
    -50.96155, -51.7942, -52.63401, -53.48095, -54.33502, -55.19618, 
    -56.06439, -56.93961, -57.82175, -58.71076, -59.60653, -60.50896, 
    -61.41792, -62.33329, -63.25488, -64.18253, -65.11604, -66.05517, 
    -66.99967, -67.94925, -68.90359, -69.86233, -70.82504, -71.79124, 
    -72.76041, -73.73187, -74.70488, -75.67852, -76.65166, -77.62291, 
    -78.59045, -79.55191, -80.5041, -81.44252, -82.3607, -83.249, -84.09252, 
    -84.8678, -85.53786, -86.04778, -86.32938, -86.32938, -86.04778, 
    -85.53786, -84.8678, -84.09252, -83.249, -82.3607, -81.44252, -80.5041, 
    -79.55191, -78.59045, -77.62291, -76.65166, -75.67852, -74.70488, 
    -73.73187, -72.76041, -71.79124, -70.82504, -69.86233, -68.90359, 
    -67.94925, -66.99967, -66.05517, -65.11604, -64.18253, -63.25488, 
    -62.33329, -61.41792, -60.50896, -59.60653, -58.71076, -57.82175, 
    -56.93961, -56.06439, -55.19618, -54.33502, -53.48095, -52.63401, 
    -51.7942, -50.96155, -50.13604, -49.31768, -48.50644, -47.7023, 
    -46.90523, -46.11519, -45.33213,
  -45.36115, -46.14581, -46.93755, -47.7364, -48.54241, -49.35562, -50.17606, 
    -51.00375, -51.8387, -52.68093, -53.53043, -54.3872, -55.25121, 
    -56.12244, -57.00084, -57.88636, -58.77895, -59.67853, -60.58501, 
    -61.49828, -62.41824, -63.34475, -64.27767, -65.21684, -66.16206, 
    -67.11313, -68.06983, -69.03191, -69.99909, -70.97105, -71.94746, 
    -72.92789, -73.91193, -74.89902, -75.88858, -76.87985, -77.87194, 
    -78.86371, -79.85367, -80.83981, -81.81931, -82.78796, -83.73922, 
    -84.66222, -85.53786, -86.33054, -86.97294, -87.35221, -87.35221, 
    -86.97294, -86.33054, -85.53786, -84.66222, -83.73922, -82.78796, 
    -81.81931, -80.83981, -79.85367, -78.86371, -77.87194, -76.87985, 
    -75.88858, -74.89902, -73.91193, -72.92789, -71.94746, -70.97105, 
    -69.99909, -69.03191, -68.06983, -67.11313, -66.16206, -65.21684, 
    -64.27767, -63.34475, -62.41824, -61.49828, -60.58501, -59.67853, 
    -58.77895, -57.88636, -57.00084, -56.12244, -55.25121, -54.3872, 
    -53.53043, -52.68093, -51.8387, -51.00375, -50.17606, -49.35562, 
    -48.54241, -47.7364, -46.93755, -46.14581, -45.36115,
  -45.3805, -46.16624, -46.95911, -47.75915, -48.56641, -49.38094, -50.20276, 
    -51.03191, -51.8684, -52.71225, -53.56347, -54.42204, -55.28796, 
    -56.1612, -57.04174, -57.92953, -58.82452, -59.72665, -60.63584, 
    -61.55201, -62.47506, -63.40488, -64.34134, -65.28431, -66.23363, 
    -67.18914, -68.15065, -69.11797, -70.09087, -71.06911, -72.05244, 
    -73.04058, -74.03321, -75.02998, -76.03052, -77.03436, -78.04102, 
    -79.04986, -80.06013, -81.07088, -82.08073, -83.08778, -84.08896, 
    -85.079, -86.04778, -86.97294, -87.79688, -88.35755, -88.35755, 
    -87.79688, -86.97294, -86.04778, -85.079, -84.08896, -83.08778, 
    -82.08073, -81.07088, -80.06013, -79.04986, -78.04102, -77.03436, 
    -76.03052, -75.02998, -74.03321, -73.04058, -72.05244, -71.06911, 
    -70.09087, -69.11797, -68.15065, -67.18914, -66.23363, -65.28431, 
    -64.34134, -63.40488, -62.47506, -61.55201, -60.63584, -59.72665, 
    -58.82452, -57.92953, -57.04174, -56.1612, -55.28796, -54.42204, 
    -53.56347, -52.71225, -51.8684, -51.03191, -50.20276, -49.38094, 
    -48.56641, -47.75915, -46.95911, -46.16624, -45.3805,
  -45.39018, -46.17646, -46.96989, -47.77053, -48.57842, -49.3936, -50.21612, 
    -51.046, -51.88326, -52.72793, -53.58, -54.43948, -55.30635, -56.18061, 
    -57.06222, -57.95115, -58.84734, -59.75075, -60.6613, -61.57893, 
    -62.50353, -63.43501, -64.37325, -65.31813, -66.26952, -67.22726, 
    -68.19119, -69.16115, -70.13693, -71.11835, -72.10519, -73.09724, 
    -74.09423, -75.09593, -76.10207, -77.11236, -78.1265, -79.14419, 
    -80.16506, -81.18875, -82.21483, -83.24277, -84.27195, -85.30138, 
    -86.32938, -87.35221, -88.35755, -89.26539, -89.26539, -88.35755, 
    -87.35221, -86.32938, -85.30138, -84.27195, -83.24277, -82.21483, 
    -81.18875, -80.16506, -79.14419, -78.1265, -77.11236, -76.10207, 
    -75.09593, -74.09423, -73.09724, -72.10519, -71.11835, -70.13693, 
    -69.16115, -68.19119, -67.22726, -66.26952, -65.31813, -64.37325, 
    -63.43501, -62.50353, -61.57893, -60.6613, -59.75075, -58.84734, 
    -57.95115, -57.06222, -56.18061, -55.30635, -54.43948, -53.58, -52.72793, 
    -51.88326, -51.046, -50.21612, -49.3936, -48.57842, -47.77053, -46.96989, 
    -46.17646, -45.39018,
  -45.39018, -46.17646, -46.96989, -47.77053, -48.57842, -49.3936, -50.21612, 
    -51.046, -51.88326, -52.72793, -53.58, -54.43948, -55.30635, -56.18061, 
    -57.06222, -57.95115, -58.84734, -59.75075, -60.6613, -61.57893, 
    -62.50353, -63.43501, -64.37325, -65.31813, -66.26952, -67.22726, 
    -68.19119, -69.16115, -70.13693, -71.11835, -72.10519, -73.09724, 
    -74.09423, -75.09593, -76.10207, -77.11236, -78.1265, -79.14419, 
    -80.16506, -81.18875, -82.21483, -83.24277, -84.27195, -85.30138, 
    -86.32938, -87.35221, -88.35755, -89.26539, -89.26539, -88.35755, 
    -87.35221, -86.32938, -85.30138, -84.27195, -83.24277, -82.21483, 
    -81.18875, -80.16506, -79.14419, -78.1265, -77.11236, -76.10207, 
    -75.09593, -74.09423, -73.09724, -72.10519, -71.11835, -70.13693, 
    -69.16115, -68.19119, -67.22726, -66.26952, -65.31813, -64.37325, 
    -63.43501, -62.50353, -61.57893, -60.6613, -59.75075, -58.84734, 
    -57.95115, -57.06222, -56.18061, -55.30635, -54.43948, -53.58, -52.72793, 
    -51.88326, -51.046, -50.21612, -49.3936, -48.57842, -47.77053, -46.96989, 
    -46.17646, -45.39018,
  -45.3805, -46.16624, -46.95911, -47.75915, -48.56641, -49.38094, -50.20276, 
    -51.03191, -51.8684, -52.71225, -53.56347, -54.42204, -55.28796, 
    -56.1612, -57.04174, -57.92953, -58.82452, -59.72665, -60.63584, 
    -61.55201, -62.47506, -63.40488, -64.34134, -65.28431, -66.23363, 
    -67.18914, -68.15065, -69.11797, -70.09087, -71.06911, -72.05244, 
    -73.04058, -74.03321, -75.02998, -76.03052, -77.03436, -78.04102, 
    -79.04986, -80.06013, -81.07088, -82.08073, -83.08778, -84.08896, 
    -85.079, -86.04778, -86.97294, -87.79688, -88.35755, -88.35755, 
    -87.79688, -86.97294, -86.04778, -85.079, -84.08896, -83.08778, 
    -82.08073, -81.07088, -80.06013, -79.04986, -78.04102, -77.03436, 
    -76.03052, -75.02998, -74.03321, -73.04058, -72.05244, -71.06911, 
    -70.09087, -69.11797, -68.15065, -67.18914, -66.23363, -65.28431, 
    -64.34134, -63.40488, -62.47506, -61.55201, -60.63584, -59.72665, 
    -58.82452, -57.92953, -57.04174, -56.1612, -55.28796, -54.42204, 
    -53.56347, -52.71225, -51.8684, -51.03191, -50.20276, -49.38094, 
    -48.56641, -47.75915, -46.95911, -46.16624, -45.3805,
  -45.36115, -46.14581, -46.93755, -47.7364, -48.54241, -49.35562, -50.17606, 
    -51.00375, -51.8387, -52.68093, -53.53043, -54.3872, -55.25121, 
    -56.12244, -57.00084, -57.88636, -58.77895, -59.67853, -60.58501, 
    -61.49828, -62.41824, -63.34475, -64.27767, -65.21684, -66.16206, 
    -67.11313, -68.06983, -69.03191, -69.99909, -70.97105, -71.94746, 
    -72.92789, -73.91193, -74.89902, -75.88858, -76.87985, -77.87194, 
    -78.86371, -79.85367, -80.83981, -81.81931, -82.78796, -83.73922, 
    -84.66222, -85.53786, -86.33054, -86.97294, -87.35221, -87.35221, 
    -86.97294, -86.33054, -85.53786, -84.66222, -83.73922, -82.78796, 
    -81.81931, -80.83981, -79.85367, -78.86371, -77.87194, -76.87985, 
    -75.88858, -74.89902, -73.91193, -72.92789, -71.94746, -70.97105, 
    -69.99909, -69.03191, -68.06983, -67.11313, -66.16206, -65.21684, 
    -64.27767, -63.34475, -62.41824, -61.49828, -60.58501, -59.67853, 
    -58.77895, -57.88636, -57.00084, -56.12244, -55.25121, -54.3872, 
    -53.53043, -52.68093, -51.8387, -51.00375, -50.17606, -49.35562, 
    -48.54241, -47.7364, -46.93755, -46.14581, -45.36115,
  -45.33213, -46.11519, -46.90523, -47.7023, -48.50644, -49.31768, -50.13604, 
    -50.96155, -51.7942, -52.63401, -53.48095, -54.33502, -55.19618, 
    -56.06439, -56.93961, -57.82175, -58.71076, -59.60653, -60.50896, 
    -61.41792, -62.33329, -63.25488, -64.18253, -65.11604, -66.05517, 
    -66.99967, -67.94925, -68.90359, -69.86233, -70.82504, -71.79124, 
    -72.76041, -73.73187, -74.70488, -75.67852, -76.65166, -77.62291, 
    -78.59045, -79.55191, -80.5041, -81.44252, -82.3607, -83.249, -84.09252, 
    -84.8678, -85.53786, -86.04778, -86.32938, -86.32938, -86.04778, 
    -85.53786, -84.8678, -84.09252, -83.249, -82.3607, -81.44252, -80.5041, 
    -79.55191, -78.59045, -77.62291, -76.65166, -75.67852, -74.70488, 
    -73.73187, -72.76041, -71.79124, -70.82504, -69.86233, -68.90359, 
    -67.94925, -66.99967, -66.05517, -65.11604, -64.18253, -63.25488, 
    -62.33329, -61.41792, -60.50896, -59.60653, -58.71076, -57.82175, 
    -56.93961, -56.06439, -55.19618, -54.33502, -53.48095, -52.63401, 
    -51.7942, -50.96155, -50.13604, -49.31768, -48.50644, -47.7023, 
    -46.90523, -46.11519, -45.33213,
  -45.29348, -46.07439, -46.86219, -47.65689, -48.45854, -49.26716, 
    -50.08277, -50.90538, -51.73498, -52.57156, -53.41512, -54.26561, 
    -55.12299, -55.9872, -56.85819, -57.73586, -58.62013, -59.51086, 
    -60.40795, -61.31122, -62.22052, -63.13563, -64.05634, -64.98241, 
    -65.91354, -66.84942, -67.78967, -68.7339, -69.68162, -70.63229, 
    -71.58528, -72.53986, -73.49516, -74.45013, -75.40351, -76.35376, 
    -77.2989, -78.23647, -79.16319, -80.07474, -80.96523, -81.82646, 
    -82.6469, -83.41006, -84.09252, -84.66222, -85.079, -85.30138, -85.30138, 
    -85.079, -84.66222, -84.09252, -83.41006, -82.6469, -81.82646, -80.96523, 
    -80.07474, -79.16319, -78.23647, -77.2989, -76.35376, -75.40351, 
    -74.45013, -73.49516, -72.53986, -71.58528, -70.63229, -69.68162, 
    -68.7339, -67.78967, -66.84942, -65.91354, -64.98241, -64.05634, 
    -63.13563, -62.22052, -61.31122, -60.40795, -59.51086, -58.62013, 
    -57.73586, -56.85819, -55.9872, -55.12299, -54.26561, -53.41512, 
    -52.57156, -51.73498, -50.90538, -50.08277, -49.26716, -48.45854, 
    -47.65689, -46.86219, -46.07439, -45.29348,
  -45.24522, -46.02346, -46.80845, -47.6002, -48.39876, -49.20412, -50.01631, 
    -50.83531, -51.66111, -52.4937, -53.33304, -54.17908, -55.03177, 
    -55.89104, -56.75679, -57.62892, -58.50731, -59.39183, -60.2823, 
    -61.17855, -62.08035, -62.98748, -63.89967, -64.81659, -65.73791, 
    -66.66322, -67.59209, -68.52398, -69.45831, -70.39439, -71.33143, 
    -72.26848, -73.20444, -74.13797, -75.06745, -75.99091, -76.90587, 
    -77.8092, -78.69691, -79.56378, -80.40296, -81.20532, -81.95869, 
    -82.6469, -83.249, -83.73922, -84.08896, -84.27195, -84.27195, -84.08896, 
    -83.73922, -83.249, -82.6469, -81.95869, -81.20532, -80.40296, -79.56378, 
    -78.69691, -77.8092, -76.90587, -75.99091, -75.06745, -74.13797, 
    -73.20444, -72.26848, -71.33143, -70.39439, -69.45831, -68.52398, 
    -67.59209, -66.66322, -65.73791, -64.81659, -63.89967, -62.98748, 
    -62.08035, -61.17855, -60.2823, -59.39183, -58.50731, -57.62892, 
    -56.75679, -55.89104, -55.03177, -54.17908, -53.33304, -52.4937, 
    -51.66111, -50.83531, -50.01631, -49.20412, -48.39876, -47.6002, 
    -46.80845, -46.02346, -45.24522,
  -45.18737, -45.96243, -46.74407, -47.53231, -48.32716, -49.12864, 
    -49.93674, -50.75143, -51.57272, -52.40054, -53.23486, -54.07561, 
    -54.92273, -55.7761, -56.63563, -57.50119, -58.37262, -59.24976, 
    -60.13241, -61.02035, -61.91332, -62.81103, -63.71317, -64.61935, 
    -65.52915, -66.44211, -67.35767, -68.2752, -69.19399, -70.1132, 
    -71.03188, -71.94884, -72.86278, -73.77206, -74.67474, -75.56844, 
    -76.45026, -77.31655, -78.16277, -78.98316, -79.77036, -80.51504, 
    -81.20532, -81.82646, -82.3607, -82.78796, -83.08778, -83.24277, 
    -83.24277, -83.08778, -82.78796, -82.3607, -81.82646, -81.20532, 
    -80.51504, -79.77036, -78.98316, -78.16277, -77.31655, -76.45026, 
    -75.56844, -74.67474, -73.77206, -72.86278, -71.94884, -71.03188, 
    -70.1132, -69.19399, -68.2752, -67.35767, -66.44211, -65.52915, 
    -64.61935, -63.71317, -62.81103, -61.91332, -61.02035, -60.13241, 
    -59.24976, -58.37262, -57.50119, -56.63563, -55.7761, -54.92273, 
    -54.07561, -53.23486, -52.40054, -51.57272, -50.75143, -49.93674, 
    -49.12864, -48.32716, -47.53231, -46.74407, -45.96243, -45.18737,
  -45.11999, -45.89135, -46.66909, -47.45325, -48.24382, -49.04079, 
    -49.84415, -50.65387, -51.46992, -52.29223, -53.12075, -53.95539, 
    -54.79607, -55.64265, -56.49501, -57.35299, -58.21642, -59.08508, 
    -59.95875, -60.83716, -61.72001, -62.60696, -63.49763, -64.39157, 
    -65.2883, -66.18724, -67.08776, -67.98912, -68.89046, -69.79082, 
    -70.68905, -71.5838, -72.47352, -73.35633, -74.23001, -75.09187, 
    -75.93864, -76.76637, -77.57013, -78.34393, -79.08037, -79.77036, 
    -80.40296, -80.96523, -81.44252, -81.81931, -82.08073, -82.21483, 
    -82.21483, -82.08073, -81.81931, -81.44252, -80.96523, -80.40296, 
    -79.77036, -79.08037, -78.34393, -77.57013, -76.76637, -75.93864, 
    -75.09187, -74.23001, -73.35633, -72.47352, -71.5838, -70.68905, 
    -69.79082, -68.89046, -67.98912, -67.08776, -66.18724, -65.2883, 
    -64.39157, -63.49763, -62.60696, -61.72001, -60.83716, -59.95875, 
    -59.08508, -58.21642, -57.35299, -56.49501, -55.64265, -54.79607, 
    -53.95539, -53.12075, -52.29223, -51.46992, -50.65387, -49.84415, 
    -49.04079, -48.24382, -47.45325, -46.66909, -45.89135, -45.11999,
  -45.04311, -45.81026, -46.5836, -47.36312, -48.14882, -48.94068, -49.73867, 
    -50.54276, -51.35287, -52.16895, -52.99091, -53.81864, -54.65204, 
    -55.49096, -56.33524, -57.18469, -58.0391, -58.89825, -59.76184, 
    -60.62958, -61.50111, -62.37604, -63.25393, -64.13426, -65.01648, 
    -65.89993, -66.78387, -67.66744, -68.54969, -69.4295, -70.30556, 
    -71.17637, -72.04017, -72.89487, -73.73804, -74.56674, -75.37749, 
    -76.16611, -76.9276, -77.65593, -78.34393, -78.98316, -79.56378, 
    -80.07474, -80.5041, -80.83981, -81.07088, -81.18875, -81.18875, 
    -81.07088, -80.83981, -80.5041, -80.07474, -79.56378, -78.98316, 
    -78.34393, -77.65593, -76.9276, -76.16611, -75.37749, -74.56674, 
    -73.73804, -72.89487, -72.04017, -71.17637, -70.30556, -69.4295, 
    -68.54969, -67.66744, -66.78387, -65.89993, -65.01648, -64.13426, 
    -63.25393, -62.37604, -61.50111, -60.62958, -59.76184, -58.89825, 
    -58.0391, -57.18469, -56.33524, -55.49096, -54.65204, -53.81864, 
    -52.99091, -52.16895, -51.35287, -50.54276, -49.73867, -48.94068, 
    -48.14882, -47.36312, -46.5836, -45.81026, -45.04311,
  -44.9568, -45.71924, -46.48764, -47.26199, -48.04226, -48.82842, -49.62043, 
    -50.41822, -51.22174, -52.03088, -52.84554, -53.6656, -54.49093, 
    -55.32135, -56.15667, -56.99669, -57.84115, -58.68978, -59.54227, 
    -60.39826, -61.25736, -62.11912, -62.98302, -63.84851, -64.71494, 
    -65.58157, -66.44756, -67.31198, -68.17374, -69.03159, -69.88412, 
    -70.72966, -71.56628, -72.39178, -73.20351, -73.99841, -74.77289, 
    -75.5227, -76.24287, -76.9276, -77.57013, -78.16277, -78.69691, 
    -79.16319, -79.55191, -79.85367, -80.06013, -80.16506, -80.16506, 
    -80.06013, -79.85367, -79.55191, -79.16319, -78.69691, -78.16277, 
    -77.57013, -76.9276, -76.24287, -75.5227, -74.77289, -73.99841, 
    -73.20351, -72.39178, -71.56628, -70.72966, -69.88412, -69.03159, 
    -68.17374, -67.31198, -66.44756, -65.58157, -64.71494, -63.84851, 
    -62.98302, -62.11912, -61.25736, -60.39826, -59.54227, -58.68978, 
    -57.84115, -56.99669, -56.15667, -55.32135, -54.49093, -53.6656, 
    -52.84554, -52.03088, -51.22174, -50.41822, -49.62043, -48.82842, 
    -48.04226, -47.26199, -46.48764, -45.71924, -44.9568,
  -44.8611, -45.61835, -46.38132, -47.14996, -47.92425, -48.70414, -49.48956, 
    -50.28045, -51.0767, -51.87823, -52.68489, -53.49655, -54.31304, 
    -55.13416, -55.95971, -56.78943, -57.62305, -58.46024, -59.30067, 
    -60.14393, -60.98957, -61.8371, -62.68594, -63.53547, -64.38497, 
    -65.23363, -66.08053, -66.92463, -67.76476, -68.59956, -69.42749, 
    -70.24678, -71.0554, -71.85101, -72.6309, -73.39191, -74.13045, 
    -74.84232, -75.5227, -76.16611, -76.76637, -77.31655, -77.8092, 
    -78.23647, -78.59045, -78.86371, -79.04986, -79.14419, -79.14419, 
    -79.04986, -78.86371, -78.59045, -78.23647, -77.8092, -77.31655, 
    -76.76637, -76.16611, -75.5227, -74.84232, -74.13045, -73.39191, 
    -72.6309, -71.85101, -71.0554, -70.24678, -69.42749, -68.59956, 
    -67.76476, -66.92463, -66.08053, -65.23363, -64.38497, -63.53547, 
    -62.68594, -61.8371, -60.98957, -60.14393, -59.30067, -58.46024, 
    -57.62305, -56.78943, -55.95971, -55.13416, -54.31304, -53.49655, 
    -52.68489, -51.87823, -51.0767, -50.28045, -49.48956, -48.70414, 
    -47.92425, -47.14996, -46.38132, -45.61835, -44.8611,
  -44.75608, -45.50768, -46.26471, -47.02713, -47.79491, -48.56796, 
    -49.34622, -50.12959, -50.91797, -51.71123, -52.50922, -53.31178, 
    -54.1187, -54.92978, -55.74477, -56.56339, -57.38533, -58.21024, 
    -59.03772, -59.86734, -60.6986, -61.53094, -62.36376, -63.19636, 
    -64.02795, -64.85765, -65.68449, -66.50732, -67.32491, -68.13581, 
    -68.9384, -69.73082, -70.51096, -71.27643, -72.02446, -72.75193, 
    -73.45528, -74.13045, -74.77289, -75.37749, -75.93864, -76.45026, 
    -76.90587, -77.2989, -77.62291, -77.87194, -78.04102, -78.1265, -78.1265, 
    -78.04102, -77.87194, -77.62291, -77.2989, -76.90587, -76.45026, 
    -75.93864, -75.37749, -74.77289, -74.13045, -73.45528, -72.75193, 
    -72.02446, -71.27643, -70.51096, -69.73082, -68.9384, -68.13581, 
    -67.32491, -66.50732, -65.68449, -64.85765, -64.02795, -63.19636, 
    -62.36376, -61.53094, -60.6986, -59.86734, -59.03772, -58.21024, 
    -57.38533, -56.56339, -55.74477, -54.92978, -54.1187, -53.31178, 
    -52.50922, -51.71123, -50.91797, -50.12959, -49.34622, -48.56796, 
    -47.79491, -47.02713, -46.26471, -45.50768, -44.75608,
  -44.64181, -45.38729, -46.13791, -46.89362, -47.65435, -48.42004, 
    -49.19058, -49.96586, -50.74577, -51.53014, -52.31881, -53.1116, 
    -53.90828, -54.70861, -55.51231, -56.31908, -57.12857, -57.9404, 
    -58.75413, -59.56929, -60.38533, -61.20166, -62.0176, -62.83242, 
    -63.64526, -64.4552, -65.26118, -66.06201, -66.85638, -67.64278, 
    -68.41954, -69.18474, -69.93623, -70.67162, -71.38813, -72.08273, 
    -72.75193, -73.39191, -73.99841, -74.56674, -75.09187, -75.56844, 
    -75.99091, -76.35376, -76.65166, -76.87985, -77.03436, -77.11236, 
    -77.11236, -77.03436, -76.87985, -76.65166, -76.35376, -75.99091, 
    -75.56844, -75.09187, -74.56674, -73.99841, -73.39191, -72.75193, 
    -72.08273, -71.38813, -70.67162, -69.93623, -69.18474, -68.41954, 
    -67.64278, -66.85638, -66.06201, -65.26118, -64.4552, -63.64526, 
    -62.83242, -62.0176, -61.20166, -60.38533, -59.56929, -58.75413, 
    -57.9404, -57.12857, -56.31908, -55.51231, -54.70861, -53.90828, 
    -53.1116, -52.31881, -51.53014, -50.74577, -49.96586, -49.19058, 
    -48.42004, -47.65435, -46.89362, -46.13791, -45.38729, -44.64181,
  -44.51836, -45.25727, -46.00101, -46.74953, -47.50273, -48.26053, 
    -49.02282, -49.78946, -50.56031, -51.33521, -52.11396, -52.89635, 
    -53.68214, -54.47105, -55.2628, -56.05703, -56.85336, -57.65139, 
    -58.45065, -59.25061, -60.05069, -60.85027, -61.64861, -62.44493, 
    -63.23833, -64.02785, -64.81236, -65.59063, -66.36131, -67.12283, 
    -67.8735, -68.61138, -69.33433, -70.03993, -70.72552, -71.38813, 
    -72.02446, -72.6309, -73.20351, -73.73804, -74.23001, -74.67474, 
    -75.06745, -75.40351, -75.67852, -75.88858, -76.03052, -76.10207, 
    -76.10207, -76.03052, -75.88858, -75.67852, -75.40351, -75.06745, 
    -74.67474, -74.23001, -73.73804, -73.20351, -72.6309, -72.02446, 
    -71.38813, -70.72552, -70.03993, -69.33433, -68.61138, -67.8735, 
    -67.12283, -66.36131, -65.59063, -64.81236, -64.02785, -63.23833, 
    -62.44493, -61.64861, -60.85027, -60.05069, -59.25061, -58.45065, 
    -57.65139, -56.85336, -56.05703, -55.2628, -54.47105, -53.68214, 
    -52.89635, -52.11396, -51.33521, -50.56031, -49.78946, -49.02282, 
    -48.26053, -47.50273, -46.74953, -46.00101, -45.25727, -44.51836,
  -44.38583, -45.11773, -45.85415, -46.595, -47.34019, -48.08961, -48.84312, 
    -49.6006, -50.36186, -51.12672, -51.89498, -52.66639, -53.44069, 
    -54.21758, -54.99673, -55.77778, -56.56032, -57.34391, -58.12803, 
    -58.91215, -59.69563, -60.47782, -61.25794, -62.03517, -62.80859, 
    -63.57715, -64.33974, -65.09508, -65.84176, -66.57823, -67.30276, 
    -68.01344, -68.70814, -69.38449, -70.03993, -70.67162, -71.27643, 
    -71.85101, -72.39178, -72.89487, -73.35633, -73.77206, -74.13797, 
    -74.45013, -74.70488, -74.89902, -75.02998, -75.09593, -75.09593, 
    -75.02998, -74.89902, -74.70488, -74.45013, -74.13797, -73.77206, 
    -73.35633, -72.89487, -72.39178, -71.85101, -71.27643, -70.67162, 
    -70.03993, -69.38449, -68.70814, -68.01344, -67.30276, -66.57823, 
    -65.84176, -65.09508, -64.33974, -63.57715, -62.80859, -62.03517, 
    -61.25794, -60.47782, -59.69563, -58.91215, -58.12803, -57.34391, 
    -56.56032, -55.77778, -54.99673, -54.21758, -53.44069, -52.66639, 
    -51.89498, -51.12672, -50.36186, -49.6006, -48.84312, -48.08961, 
    -47.34019, -46.595, -45.85415, -45.11773, -44.38583,
  -44.24429, -44.96877, -45.69742, -46.43016, -47.16688, -47.90744, -48.6517, 
    -49.39951, -50.15067, -50.90497, -51.66219, -52.42207, -53.18432, 
    -53.94862, -54.71461, -55.48191, -56.25008, -57.01865, -57.78707, 
    -58.55478, -59.32111, -60.08537, -60.84677, -61.60444, -62.35743, 
    -63.10468, -63.84503, -64.57719, -65.29976, -66.01116, -66.70969, 
    -67.39344, -68.06035, -68.70814, -69.33433, -69.93623, -70.51096, 
    -71.0554, -71.56628, -72.04017, -72.47352, -72.86278, -73.20444, 
    -73.49516, -73.73187, -73.91193, -74.03321, -74.09423, -74.09423, 
    -74.03321, -73.91193, -73.73187, -73.49516, -73.20444, -72.86278, 
    -72.47352, -72.04017, -71.56628, -71.0554, -70.51096, -69.93623, 
    -69.33433, -68.70814, -68.06035, -67.39344, -66.70969, -66.01116, 
    -65.29976, -64.57719, -63.84503, -63.10468, -62.35743, -61.60444, 
    -60.84677, -60.08537, -59.32111, -58.55478, -57.78707, -57.01865, 
    -56.25008, -55.48191, -54.71461, -53.94862, -53.18432, -52.42207, 
    -51.66219, -50.90497, -50.15067, -49.39951, -48.6517, -47.90744, 
    -47.16688, -46.43016, -45.69742, -44.96877, -44.24429,
  -44.09382, -44.81047, -45.53096, -46.25516, -46.98296, -47.71421, 
    -48.44876, -49.18642, -49.927, -50.67025, -51.41594, -52.16379, 
    -52.91348, -53.66467, -54.41699, -55.17002, -55.9233, -56.67633, 
    -57.42855, -58.17936, -58.92809, -59.67398, -60.41625, -61.154, 
    -61.88625, -62.61193, -63.32987, -64.03877, -64.73723, -65.42369, 
    -66.09647, -66.75372, -67.39344, -68.01344, -68.61138, -69.18474, 
    -69.73082, -70.24678, -70.72966, -71.17637, -71.5838, -71.94884, 
    -72.26848, -72.53986, -72.76041, -72.92789, -73.04058, -73.09724, 
    -73.09724, -73.04058, -72.92789, -72.76041, -72.53986, -72.26848, 
    -71.94884, -71.5838, -71.17637, -70.72966, -70.24678, -69.73082, 
    -69.18474, -68.61138, -68.01344, -67.39344, -66.75372, -66.09647, 
    -65.42369, -64.73723, -64.03877, -63.32987, -62.61193, -61.88625, 
    -61.154, -60.41625, -59.67398, -58.92809, -58.17936, -57.42855, 
    -56.67633, -55.9233, -55.17002, -54.41699, -53.66467, -52.91348, 
    -52.16379, -51.41594, -50.67025, -49.927, -49.18642, -48.44876, 
    -47.71421, -46.98296, -46.25516, -45.53096, -44.81047, -44.09382,
  -43.93454, -44.64297, -45.35488, -46.07014, -46.7886, -47.51012, -48.23452, 
    -48.9616, -49.69113, -50.42288, -51.15658, -51.89192, -52.62858, 
    -53.3662, -54.10438, -54.84268, -55.58062, -56.31768, -57.05328, 
    -57.78679, -58.51752, -59.24471, -59.96754, -60.6851, -61.39641, 
    -62.10038, -62.79585, -63.48152, -64.15601, -64.81778, -65.46519, 
    -66.09647, -66.70969, -67.30276, -67.8735, -68.41954, -68.9384, 
    -69.42749, -69.88412, -70.30556, -70.68905, -71.03188, -71.33143, 
    -71.58528, -71.79124, -71.94746, -72.05244, -72.10519, -72.10519, 
    -72.05244, -71.94746, -71.79124, -71.58528, -71.33143, -71.03188, 
    -70.68905, -70.30556, -69.88412, -69.42749, -68.9384, -68.41954, 
    -67.8735, -67.30276, -66.70969, -66.09647, -65.46519, -64.81778, 
    -64.15601, -63.48152, -62.79585, -62.10038, -61.39641, -60.6851, 
    -59.96754, -59.24471, -58.51752, -57.78679, -57.05328, -56.31768, 
    -55.58062, -54.84268, -54.10438, -53.3662, -52.62858, -51.89192, 
    -51.15658, -50.42288, -49.69113, -48.9616, -48.23452, -47.51012, 
    -46.7886, -46.07014, -45.35488, -44.64297, -43.93454,
  -43.76653, -44.46637, -45.16932, -45.87524, -46.58398, -47.29537, -48.0092, 
    -48.72528, -49.44336, -50.16318, -50.88446, -51.60688, -52.33009, 
    -53.05371, -53.77734, -54.5005, -55.22271, -55.94343, -56.66205, 
    -57.37793, -58.09037, -58.79859, -59.50176, -60.19897, -60.88923, 
    -61.57146, -62.2445, -62.90707, -63.55782, -64.19525, -64.81778, 
    -65.42369, -66.01116, -66.57823, -67.12283, -67.64278, -68.13581, 
    -68.59956, -69.03159, -69.4295, -69.79082, -70.1132, -70.39439, 
    -70.63229, -70.82504, -70.97105, -71.06911, -71.11835, -71.11835, 
    -71.06911, -70.97105, -70.82504, -70.63229, -70.39439, -70.1132, 
    -69.79082, -69.4295, -69.03159, -68.59956, -68.13581, -67.64278, 
    -67.12283, -66.57823, -66.01116, -65.42369, -64.81778, -64.19525, 
    -63.55782, -62.90707, -62.2445, -61.57146, -60.88923, -60.19897, 
    -59.50176, -58.79859, -58.09037, -57.37793, -56.66205, -55.94343, 
    -55.22271, -54.5005, -53.77734, -53.05371, -52.33009, -51.60688, 
    -50.88446, -50.16318, -49.44336, -48.72528, -48.0092, -47.29537, 
    -46.58398, -45.87524, -45.16932, -44.46637, -43.76653,
  -43.58989, -44.28079, -44.97443, -45.67065, -46.36929, -47.07016, 
    -47.77305, -48.47774, -49.18397, -49.89148, -50.59995, -51.30906, 
    -52.01844, -52.7277, -53.43641, -54.14409, -54.85024, -55.55429, 
    -56.25565, -56.95364, -57.64757, -58.33664, -59.02002, -59.6968, 
    -60.36599, -61.02654, -61.67727, -62.31697, -62.94429, -63.55782, 
    -64.15601, -64.73723, -65.29976, -65.84176, -66.36131, -66.85638, 
    -67.32491, -67.76476, -68.17374, -68.54969, -68.89046, -69.19399, 
    -69.45831, -69.68162, -69.86233, -69.99909, -70.09087, -70.13693, 
    -70.13693, -70.09087, -69.99909, -69.86233, -69.68162, -69.45831, 
    -69.19399, -68.89046, -68.54969, -68.17374, -67.76476, -67.32491, 
    -66.85638, -66.36131, -65.84176, -65.29976, -64.73723, -64.15601, 
    -63.55782, -62.94429, -62.31697, -61.67727, -61.02654, -60.36599, 
    -59.6968, -59.02002, -58.33664, -57.64757, -56.95364, -56.25565, 
    -55.55429, -54.85024, -54.14409, -53.43641, -52.7277, -52.01844, 
    -51.30906, -50.59995, -49.89148, -49.18397, -48.47774, -47.77305, 
    -47.07016, -46.36929, -45.67065, -44.97443, -44.28079, -43.58989,
  -43.40474, -44.08636, -44.77034, -45.45651, -46.14469, -46.83469, 
    -47.52629, -48.21923, -48.91327, -49.6081, -50.30342, -50.99888, 
    -51.6941, -52.38867, -53.08215, -53.77406, -54.46386, -55.15101, 
    -55.83487, -56.51479, -57.19004, -57.85986, -58.52339, -59.17973, 
    -59.82792, -60.4669, -61.09555, -61.71267, -62.31697, -62.90707, 
    -63.48152, -64.03877, -64.57719, -65.09508, -65.59063, -66.06201, 
    -66.50732, -66.92463, -67.31198, -67.66744, -67.98912, -68.2752, 
    -68.52398, -68.7339, -68.90359, -69.03191, -69.11797, -69.16115, 
    -69.16115, -69.11797, -69.03191, -68.90359, -68.7339, -68.52398, 
    -68.2752, -67.98912, -67.66744, -67.31198, -66.92463, -66.50732, 
    -66.06201, -65.59063, -65.09508, -64.57719, -64.03877, -63.48152, 
    -62.90707, -62.31697, -61.71267, -61.09555, -60.4669, -59.82792, 
    -59.17973, -58.52339, -57.85986, -57.19004, -56.51479, -55.83487, 
    -55.15101, -54.46386, -53.77406, -53.08215, -52.38867, -51.6941, 
    -50.99888, -50.30342, -49.6081, -48.91327, -48.21923, -47.52629, 
    -46.83469, -46.14469, -45.45651, -44.77034, -44.08636, -43.40474,
  -43.21118, -43.8832, -44.55719, -45.23299, -45.91039, -46.5892, -47.26916, 
    -47.95004, -48.63155, -49.3134, -49.99525, -50.67675, -51.35751, 
    -52.03711, -52.7151, -53.39099, -54.06424, -54.73428, -55.40049, 
    -56.06221, -56.7187, -57.36921, -58.01291, -58.64888, -59.2762, 
    -59.89382, -60.50066, -61.09555, -61.67727, -62.2445, -62.79585, 
    -63.32987, -63.84503, -64.33974, -64.81236, -65.26118, -65.68449, 
    -66.08053, -66.44756, -66.78387, -67.08776, -67.35767, -67.59209, 
    -67.78967, -67.94925, -68.06983, -68.15065, -68.19119, -68.19119, 
    -68.15065, -68.06983, -67.94925, -67.78967, -67.59209, -67.35767, 
    -67.08776, -66.78387, -66.44756, -66.08053, -65.68449, -65.26118, 
    -64.81236, -64.33974, -63.84503, -63.32987, -62.79585, -62.2445, 
    -61.67727, -61.09555, -60.50066, -59.89382, -59.2762, -58.64888, 
    -58.01291, -57.36921, -56.7187, -56.06221, -55.40049, -54.73428, 
    -54.06424, -53.39099, -52.7151, -52.03711, -51.35751, -50.67675, 
    -49.99525, -49.3134, -48.63155, -47.95004, -47.26916, -46.5892, 
    -45.91039, -45.23299, -44.55719, -43.8832, -43.21118,
  -43.00933, -43.67144, -44.33515, -45.00027, -45.66659, -46.33389, 
    -47.00192, -47.67044, -48.33913, -49.00771, -49.67582, -50.34309, 
    -51.00915, -51.67355, -52.33583, -52.9955, -53.65202, -54.30482, 
    -54.95327, -55.59671, -56.23442, -56.86565, -57.48957, -58.1053, 
    -58.71193, -59.30845, -59.89382, -60.4669, -61.02654, -61.57146, 
    -62.10038, -62.61193, -63.10468, -63.57715, -64.02785, -64.4552, 
    -64.85765, -65.23363, -65.58157, -65.89993, -66.18724, -66.44211, 
    -66.66322, -66.84942, -66.99967, -67.11313, -67.18914, -67.22726, 
    -67.22726, -67.18914, -67.11313, -66.99967, -66.84942, -66.66322, 
    -66.44211, -66.18724, -65.89993, -65.58157, -65.23363, -64.85765, 
    -64.4552, -64.02785, -63.57715, -63.10468, -62.61193, -62.10038, 
    -61.57146, -61.02654, -60.4669, -59.89382, -59.30845, -58.71193, 
    -58.1053, -57.48957, -56.86565, -56.23442, -55.59671, -54.95327, 
    -54.30482, -53.65202, -52.9955, -52.33583, -51.67355, -51.00915, 
    -50.34309, -49.67582, -49.00771, -48.33913, -47.67044, -47.00192, 
    -46.33389, -45.66659, -45.00027, -44.33515, -43.67144, -43.00933,
  -42.7993, -43.45123, -44.10437, -44.75852, -45.41347, -46.06899, -46.72482, 
    -47.3807, -48.03632, -48.69137, -49.3455, -49.99833, -50.64946, 
    -51.29846, -51.94487, -52.58817, -53.22784, -53.8633, -54.49394, 
    -55.11909, -55.73805, -56.35006, -56.95434, -57.55002, -58.1362, 
    -58.71193, -59.2762, -59.82792, -60.36599, -60.88923, -61.39641, 
    -61.88625, -62.35743, -62.80859, -63.23833, -63.64526, -64.02795, 
    -64.38497, -64.71494, -65.01648, -65.2883, -65.52915, -65.73791, 
    -65.91354, -66.05517, -66.16206, -66.23363, -66.26952, -66.26952, 
    -66.23363, -66.16206, -66.05517, -65.91354, -65.73791, -65.52915, 
    -65.2883, -65.01648, -64.71494, -64.38497, -64.02795, -63.64526, 
    -63.23833, -62.80859, -62.35743, -61.88625, -61.39641, -60.88923, 
    -60.36599, -59.82792, -59.2762, -58.71193, -58.1362, -57.55002, 
    -56.95434, -56.35006, -55.73805, -55.11909, -54.49394, -53.8633, 
    -53.22784, -52.58817, -51.94487, -51.29846, -50.64946, -49.99833, 
    -49.3455, -48.69137, -48.03632, -47.3807, -46.72482, -46.06899, 
    -45.41347, -44.75852, -44.10437, -43.45123, -42.7993,
  -42.58122, -43.22269, -43.86499, -44.50792, -45.15124, -45.79473, 
    -46.43811, -47.08112, -47.72343, -48.36473, -49.00467, -49.64286, 
    -50.2789, -50.91235, -51.54275, -52.16959, -52.79234, -53.41042, 
    -54.02324, -54.63013, -55.2304, -55.82333, -56.40814, -56.98399, 
    -57.55002, -58.1053, -58.64888, -59.17973, -59.6968, -60.19897, -60.6851, 
    -61.154, -61.60444, -62.03517, -62.44493, -62.83242, -63.19636, 
    -63.53547, -63.84851, -64.13426, -64.39157, -64.61935, -64.81659, 
    -64.98241, -65.11604, -65.21684, -65.28431, -65.31813, -65.31813, 
    -65.28431, -65.21684, -65.11604, -64.98241, -64.81659, -64.61935, 
    -64.39157, -64.13426, -63.84851, -63.53547, -63.19636, -62.83242, 
    -62.44493, -62.03517, -61.60444, -61.154, -60.6851, -60.19897, -59.6968, 
    -59.17973, -58.64888, -58.1053, -57.55002, -56.98399, -56.40814, 
    -55.82333, -55.2304, -54.63013, -54.02324, -53.41042, -52.79234, 
    -52.16959, -51.54275, -50.91235, -50.2789, -49.64286, -49.00467, 
    -48.36473, -47.72343, -47.08112, -46.43811, -45.79473, -45.15124, 
    -44.50792, -43.86499, -43.22269, -42.58122,
  -42.35519, -42.98596, -43.61718, -44.24864, -44.88011, -45.51133, 
    -46.14204, -46.77196, -47.40077, -48.02814, -48.65372, -49.27712, 
    -49.89793, -50.51572, -51.13002, -51.74033, -52.34612, -52.94683, 
    -53.54185, -54.13057, -54.71228, -55.28629, -55.85184, -56.40814, 
    -56.95434, -57.48957, -58.01291, -58.52339, -59.02002, -59.50176, 
    -59.96754, -60.41625, -60.84677, -61.25794, -61.64861, -62.0176, 
    -62.36376, -62.68594, -62.98302, -63.25393, -63.49763, -63.71317, 
    -63.89967, -64.05634, -64.18253, -64.27767, -64.34134, -64.37325, 
    -64.37325, -64.34134, -64.27767, -64.18253, -64.05634, -63.89967, 
    -63.71317, -63.49763, -63.25393, -62.98302, -62.68594, -62.36376, 
    -62.0176, -61.64861, -61.25794, -60.84677, -60.41625, -59.96754, 
    -59.50176, -59.02002, -58.52339, -58.01291, -57.48957, -56.95434, 
    -56.40814, -55.85184, -55.28629, -54.71228, -54.13057, -53.54185, 
    -52.94683, -52.34612, -51.74033, -51.13002, -50.51572, -49.89793, 
    -49.27712, -48.65372, -48.02814, -47.40077, -46.77196, -46.14204, 
    -45.51133, -44.88011, -44.24864, -43.61718, -42.98596, -42.35519,
  -42.12135, -42.74119, -43.36111, -43.98088, -44.60027, -45.21903, 
    -45.83688, -46.45353, -47.06866, -47.68195, -48.29302, -48.9015, 
    -49.50698, -50.10903, -50.70718, -51.30094, -51.88978, -52.47316, 
    -53.05048, -53.62113, -54.18444, -54.73974, -55.28629, -55.82333, 
    -56.35006, -56.86565, -57.36921, -57.85986, -58.33664, -58.79859, 
    -59.24471, -59.67398, -60.08537, -60.47782, -60.85027, -61.20166, 
    -61.53094, -61.8371, -62.11912, -62.37604, -62.60696, -62.81103, 
    -62.98748, -63.13563, -63.25488, -63.34475, -63.40488, -63.43501, 
    -63.43501, -63.40488, -63.34475, -63.25488, -63.13563, -62.98748, 
    -62.81103, -62.60696, -62.37604, -62.11912, -61.8371, -61.53094, 
    -61.20166, -60.85027, -60.47782, -60.08537, -59.67398, -59.24471, 
    -58.79859, -58.33664, -57.85986, -57.36921, -56.86565, -56.35006, 
    -55.82333, -55.28629, -54.73974, -54.18444, -53.62113, -53.05048, 
    -52.47316, -51.88978, -51.30094, -50.70718, -50.10903, -49.50698, 
    -48.9015, -48.29302, -47.68195, -47.06866, -46.45353, -45.83688, 
    -45.21903, -44.60027, -43.98088, -43.36111, -42.74119, -42.12135,
  -41.87982, -42.48852, -43.09693, -43.70482, -44.31195, -44.91806, 
    -45.52287, -46.12609, -46.72741, -47.32647, -47.92294, -48.51642, 
    -49.10651, -49.69277, -50.27475, -50.85197, -51.42391, -51.99004, 
    -52.54977, -53.10251, -53.64762, -54.18444, -54.71228, -55.2304, 
    -55.73805, -56.23442, -56.7187, -57.19004, -57.64757, -58.09037, 
    -58.51752, -58.92809, -59.32111, -59.69563, -60.05069, -60.38533, 
    -60.6986, -60.98957, -61.25736, -61.50111, -61.72001, -61.91332, 
    -62.08035, -62.22052, -62.33329, -62.41824, -62.47506, -62.50353, 
    -62.50353, -62.47506, -62.41824, -62.33329, -62.22052, -62.08035, 
    -61.91332, -61.72001, -61.50111, -61.25736, -60.98957, -60.6986, 
    -60.38533, -60.05069, -59.69563, -59.32111, -58.92809, -58.51752, 
    -58.09037, -57.64757, -57.19004, -56.7187, -56.23442, -55.73805, 
    -55.2304, -54.71228, -54.18444, -53.64762, -53.10251, -52.54977, 
    -51.99004, -51.42391, -50.85197, -50.27475, -49.69277, -49.10651, 
    -48.51642, -47.92294, -47.32647, -46.72741, -46.12609, -45.52287, 
    -44.91806, -44.31195, -43.70482, -43.09693, -42.48852, -41.87982,
  -41.63073, -42.2281, -42.82481, -43.42064, -44.01534, -44.60864, -45.20028, 
    -45.78994, -46.37732, -46.96207, -47.54385, -48.12227, -48.69693, 
    -49.2674, -49.83323, -50.39396, -50.94908, -51.49806, -52.04035, 
    -52.57537, -53.10251, -53.62113, -54.13057, -54.63013, -55.11909, 
    -55.59671, -56.06221, -56.51479, -56.95364, -57.37793, -57.78679, 
    -58.17936, -58.55478, -58.91215, -59.25061, -59.56929, -59.86734, 
    -60.14393, -60.39826, -60.62958, -60.83716, -61.02035, -61.17855, 
    -61.31122, -61.41792, -61.49828, -61.55201, -61.57893, -61.57893, 
    -61.55201, -61.49828, -61.41792, -61.31122, -61.17855, -61.02035, 
    -60.83716, -60.62958, -60.39826, -60.14393, -59.86734, -59.56929, 
    -59.25061, -58.91215, -58.55478, -58.17936, -57.78679, -57.37793, 
    -56.95364, -56.51479, -56.06221, -55.59671, -55.11909, -54.63013, 
    -54.13057, -53.62113, -53.10251, -52.57537, -52.04035, -51.49806, 
    -50.94908, -50.39396, -49.83323, -49.2674, -48.69693, -48.12227, 
    -47.54385, -46.96207, -46.37732, -45.78994, -45.20028, -44.60864, 
    -44.01534, -43.42064, -42.82481, -42.2281, -41.63073,
  -41.37419, -41.96006, -42.54491, -43.12852, -43.71065, -44.29101, 
    -44.86935, -45.44535, -46.0187, -46.58908, -47.15612, -47.71944, 
    -48.27867, -48.83337, -49.3831, -49.92742, -50.46582, -50.9978, 
    -51.52283, -52.04035, -52.54977, -53.05048, -53.54185, -54.02324, 
    -54.49394, -54.95327, -55.40049, -55.83487, -56.25565, -56.66205, 
    -57.05328, -57.42855, -57.78707, -58.12803, -58.45065, -58.75413, 
    -59.03772, -59.30067, -59.54227, -59.76184, -59.95875, -60.13241, 
    -60.2823, -60.40795, -60.50896, -60.58501, -60.63584, -60.6613, -60.6613, 
    -60.63584, -60.58501, -60.50896, -60.40795, -60.2823, -60.13241, 
    -59.95875, -59.76184, -59.54227, -59.30067, -59.03772, -58.75413, 
    -58.45065, -58.12803, -57.78707, -57.42855, -57.05328, -56.66205, 
    -56.25565, -55.83487, -55.40049, -54.95327, -54.49394, -54.02324, 
    -53.54185, -53.05048, -52.54977, -52.04035, -51.52283, -50.9978, 
    -50.46582, -49.92742, -49.3831, -48.83337, -48.27867, -47.71944, 
    -47.15612, -46.58908, -46.0187, -45.44535, -44.86935, -44.29101, 
    -43.71065, -43.12852, -42.54491, -41.96006, -41.37419,
  -41.11036, -41.68456, -42.2574, -42.82867, -43.39809, -43.9654, -44.53034, 
    -45.0926, -45.65187, -46.20782, -46.76009, -47.30833, -47.85214, 
    -48.39112, -48.92484, -49.45285, -49.97467, -50.48983, -50.9978, 
    -51.49806, -51.99004, -52.47316, -52.94683, -53.41042, -53.8633, 
    -54.30482, -54.73428, -55.15101, -55.55429, -55.94343, -56.31768, 
    -56.67633, -57.01865, -57.34391, -57.65139, -57.9404, -58.21024, 
    -58.46024, -58.68978, -58.89825, -59.08508, -59.24976, -59.39183, 
    -59.51086, -59.60653, -59.67853, -59.72665, -59.75075, -59.75075, 
    -59.72665, -59.67853, -59.60653, -59.51086, -59.39183, -59.24976, 
    -59.08508, -58.89825, -58.68978, -58.46024, -58.21024, -57.9404, 
    -57.65139, -57.34391, -57.01865, -56.67633, -56.31768, -55.94343, 
    -55.55429, -55.15101, -54.73428, -54.30482, -53.8633, -53.41042, 
    -52.94683, -52.47316, -51.99004, -51.49806, -50.9978, -50.48983, 
    -49.97467, -49.45285, -48.92484, -48.39112, -47.85214, -47.30833, 
    -46.76009, -46.20782, -45.65187, -45.0926, -44.53034, -43.9654, 
    -43.39809, -42.82867, -42.2574, -41.68456, -41.11036,
  -40.83934, -41.40174, -41.96246, -42.52125, -43.07787, -43.63205, 
    -44.18351, -44.73198, -45.27712, -45.81862, -46.35614, -46.88931, 
    -47.41776, -47.94109, -48.45889, -48.97073, -49.47615, -49.97467, 
    -50.46582, -50.94908, -51.42391, -51.88978, -52.34612, -52.79234, 
    -53.22784, -53.65202, -54.06424, -54.46386, -54.85024, -55.22271, 
    -55.58062, -55.9233, -56.25008, -56.56032, -56.85336, -57.12857, 
    -57.38533, -57.62305, -57.84115, -58.0391, -58.21642, -58.37262, 
    -58.50731, -58.62013, -58.71076, -58.77895, -58.82452, -58.84734, 
    -58.84734, -58.82452, -58.77895, -58.71076, -58.62013, -58.50731, 
    -58.37262, -58.21642, -58.0391, -57.84115, -57.62305, -57.38533, 
    -57.12857, -56.85336, -56.56032, -56.25008, -55.9233, -55.58062, 
    -55.22271, -54.85024, -54.46386, -54.06424, -53.65202, -53.22784, 
    -52.79234, -52.34612, -51.88978, -51.42391, -50.94908, -50.46582, 
    -49.97467, -49.47615, -48.97073, -48.45889, -47.94109, -47.41776, 
    -46.88931, -46.35614, -45.81862, -45.27712, -44.73198, -44.18351, 
    -43.63205, -43.07787, -42.52125, -41.96246, -41.40174, -40.83934,
  -40.56128, -41.11176, -41.66023, -42.20646, -42.75019, -43.29116, 
    -43.82911, -44.36374, -44.89474, -45.4218, -45.94459, -46.46275, 
    -46.97591, -47.4837, -47.98571, -48.48154, -48.97073, -49.45285, 
    -49.92742, -50.39396, -50.85197, -51.30094, -51.74033, -52.16959, 
    -52.58817, -52.9955, -53.39099, -53.77406, -54.14409, -54.5005, 
    -54.84268, -55.17002, -55.48191, -55.77778, -56.05703, -56.31908, 
    -56.56339, -56.78943, -56.99669, -57.18469, -57.35299, -57.50119, 
    -57.62892, -57.73586, -57.82175, -57.88636, -57.92953, -57.95115, 
    -57.95115, -57.92953, -57.88636, -57.82175, -57.73586, -57.62892, 
    -57.50119, -57.35299, -57.18469, -56.99669, -56.78943, -56.56339, 
    -56.31908, -56.05703, -55.77778, -55.48191, -55.17002, -54.84268, 
    -54.5005, -54.14409, -53.77406, -53.39099, -52.9955, -52.58817, 
    -52.16959, -51.74033, -51.30094, -50.85197, -50.39396, -49.92742, 
    -49.45285, -48.97073, -48.48154, -47.98571, -47.4837, -46.97591, 
    -46.46275, -45.94459, -45.4218, -44.89474, -44.36374, -43.82911, 
    -43.29116, -42.75019, -42.20646, -41.66023, -41.11176, -40.56128,
  -40.27629, -40.81476, -41.35089, -41.88448, -42.41526, -42.94299, 
    -43.46738, -43.98816, -44.50503, -45.01768, -45.52579, -46.029, 
    -46.52699, -47.01936, -47.50573, -47.98571, -48.45889, -48.92484, 
    -49.3831, -49.83323, -50.27475, -50.70718, -51.13002, -51.54275, 
    -51.94487, -52.33583, -52.7151, -53.08215, -53.43641, -53.77734, 
    -54.10438, -54.41699, -54.71461, -54.99673, -55.2628, -55.51231, 
    -55.74477, -55.95971, -56.15667, -56.33524, -56.49501, -56.63563, 
    -56.75679, -56.85819, -56.93961, -57.00084, -57.04174, -57.06222, 
    -57.06222, -57.04174, -57.00084, -56.93961, -56.85819, -56.75679, 
    -56.63563, -56.49501, -56.33524, -56.15667, -55.95971, -55.74477, 
    -55.51231, -55.2628, -54.99673, -54.71461, -54.41699, -54.10438, 
    -53.77734, -53.43641, -53.08215, -52.7151, -52.33583, -51.94487, 
    -51.54275, -51.13002, -50.70718, -50.27475, -49.83323, -49.3831, 
    -48.92484, -48.45889, -47.98571, -47.50573, -47.01936, -46.52699, 
    -46.029, -45.52579, -45.01768, -44.50503, -43.98816, -43.46738, 
    -42.94299, -42.41526, -41.88448, -41.35089, -40.81476, -40.27629,
  -39.98453, -40.51088, -41.03462, -41.5555, -42.07329, -42.58773, -43.09856, 
    -43.60551, -44.10828, -44.60656, -45.10006, -45.58843, -46.07135, 
    -46.54844, -47.01936, -47.4837, -47.94109, -48.39112, -48.83337, 
    -49.2674, -49.69277, -50.10903, -50.51572, -50.91235, -51.29846, 
    -51.67355, -52.03711, -52.38867, -52.7277, -53.05371, -53.3662, 
    -53.66467, -53.94862, -54.21758, -54.47105, -54.70861, -54.92978, 
    -55.13416, -55.32135, -55.49096, -55.64265, -55.7761, -55.89104, 
    -55.9872, -56.06439, -56.12244, -56.1612, -56.18061, -56.18061, -56.1612, 
    -56.12244, -56.06439, -55.9872, -55.89104, -55.7761, -55.64265, 
    -55.49096, -55.32135, -55.13416, -54.92978, -54.70861, -54.47105, 
    -54.21758, -53.94862, -53.66467, -53.3662, -53.05371, -52.7277, 
    -52.38867, -52.03711, -51.67355, -51.29846, -50.91235, -50.51572, 
    -50.10903, -49.69277, -49.2674, -48.83337, -48.39112, -47.94109, 
    -47.4837, -47.01936, -46.54844, -46.07135, -45.58843, -45.10006, 
    -44.60656, -44.10828, -43.60551, -43.09856, -42.58773, -42.07329, 
    -41.5555, -41.03462, -40.51088, -39.98453,
  -39.68611, -40.20029, -40.71156, -41.2197, -41.72447, -42.22562, -42.7229, 
    -43.21604, -43.70475, -44.18875, -44.66773, -45.14137, -45.60936, 
    -46.07135, -46.52699, -46.97591, -47.41776, -47.85214, -48.27867, 
    -48.69693, -49.10651, -49.50698, -49.89793, -50.2789, -50.64946, 
    -51.00915, -51.35751, -51.6941, -52.01844, -52.33009, -52.62858, 
    -52.91348, -53.18432, -53.44069, -53.68214, -53.90828, -54.1187, 
    -54.31304, -54.49093, -54.65204, -54.79607, -54.92273, -55.03177, 
    -55.12299, -55.19618, -55.25121, -55.28796, -55.30635, -55.30635, 
    -55.28796, -55.25121, -55.19618, -55.12299, -55.03177, -54.92273, 
    -54.79607, -54.65204, -54.49093, -54.31304, -54.1187, -53.90828, 
    -53.68214, -53.44069, -53.18432, -52.91348, -52.62858, -52.33009, 
    -52.01844, -51.6941, -51.35751, -51.00915, -50.64946, -50.2789, 
    -49.89793, -49.50698, -49.10651, -48.69693, -48.27867, -47.85214, 
    -47.41776, -46.97591, -46.52699, -46.07135, -45.60936, -45.14137, 
    -44.66773, -44.18875, -43.70475, -43.21604, -42.7229, -42.22562, 
    -41.72447, -41.2197, -40.71156, -40.20029, -39.68611,
  -39.38117, -39.88312, -40.38189, -40.87727, -41.36901, -41.85689, 
    -42.34064, -42.82002, -43.29474, -43.76454, -44.22911, -44.68816, 
    -45.14137, -45.58843, -46.029, -46.46275, -46.88931, -47.30833, 
    -47.71944, -48.12227, -48.51642, -48.9015, -49.27712, -49.64286, 
    -49.99833, -50.34309, -50.67675, -50.99888, -51.30906, -51.60688, 
    -51.89192, -52.16379, -52.42207, -52.66639, -52.89635, -53.1116, 
    -53.31178, -53.49655, -53.6656, -53.81864, -53.95539, -54.07561, 
    -54.17908, -54.26561, -54.33502, -54.3872, -54.42204, -54.43948, 
    -54.43948, -54.42204, -54.3872, -54.33502, -54.26561, -54.17908, 
    -54.07561, -53.95539, -53.81864, -53.6656, -53.49655, -53.31178, 
    -53.1116, -52.89635, -52.66639, -52.42207, -52.16379, -51.89192, 
    -51.60688, -51.30906, -50.99888, -50.67675, -50.34309, -49.99833, 
    -49.64286, -49.27712, -48.9015, -48.51642, -48.12227, -47.71944, 
    -47.30833, -46.88931, -46.46275, -46.029, -45.58843, -45.14137, 
    -44.68816, -44.22911, -43.76454, -43.29474, -42.82002, -42.34064, 
    -41.85689, -41.36901, -40.87727, -40.38189, -39.88312, -39.38117,
  -39.06984, -39.55952, -40.04577, -40.52837, -41.00711, -41.48173, 
    -41.95201, -42.41769, -42.87851, -43.33421, -43.7845, -44.22911, 
    -44.66773, -45.10006, -45.52579, -45.94459, -46.35614, -46.76009, 
    -47.15612, -47.54385, -47.92294, -48.29302, -48.65372, -49.00467, 
    -49.3455, -49.67582, -49.99525, -50.30342, -50.59995, -50.88446, 
    -51.15658, -51.41594, -51.66219, -51.89498, -52.11396, -52.31881, 
    -52.50922, -52.68489, -52.84554, -52.99091, -53.12075, -53.23486, 
    -53.33304, -53.41512, -53.48095, -53.53043, -53.56347, -53.58, -53.58, 
    -53.56347, -53.53043, -53.48095, -53.41512, -53.33304, -53.23486, 
    -53.12075, -52.99091, -52.84554, -52.68489, -52.50922, -52.31881, 
    -52.11396, -51.89498, -51.66219, -51.41594, -51.15658, -50.88446, 
    -50.59995, -50.30342, -49.99525, -49.67582, -49.3455, -49.00467, 
    -48.65372, -48.29302, -47.92294, -47.54385, -47.15612, -46.76009, 
    -46.35614, -45.94459, -45.52579, -45.10006, -44.66773, -44.22911, 
    -43.7845, -43.33421, -42.87851, -42.41769, -41.95201, -41.48173, 
    -41.00711, -40.52837, -40.04577, -39.55952, -39.06984,
  -38.75225, -39.22964, -39.70337, -40.17321, -40.63895, -41.10036, 
    -41.55723, -42.0093, -42.45632, -42.89805, -43.33421, -43.76454, 
    -44.18875, -44.60656, -45.01768, -45.4218, -45.81862, -46.20782, 
    -46.58908, -46.96207, -47.32647, -47.68195, -48.02814, -48.36473, 
    -48.69137, -49.00771, -49.3134, -49.6081, -49.89148, -50.16318, 
    -50.42288, -50.67025, -50.90497, -51.12672, -51.33521, -51.53014, 
    -51.71123, -51.87823, -52.03088, -52.16895, -52.29223, -52.40054, 
    -52.4937, -52.57156, -52.63401, -52.68093, -52.71225, -52.72793, 
    -52.72793, -52.71225, -52.68093, -52.63401, -52.57156, -52.4937, 
    -52.40054, -52.29223, -52.16895, -52.03088, -51.87823, -51.71123, 
    -51.53014, -51.33521, -51.12672, -50.90497, -50.67025, -50.42288, 
    -50.16318, -49.89148, -49.6081, -49.3134, -49.00771, -48.69137, 
    -48.36473, -48.02814, -47.68195, -47.32647, -46.96207, -46.58908, 
    -46.20782, -45.81862, -45.4218, -45.01768, -44.60656, -44.18875, 
    -43.76454, -43.33421, -42.89805, -42.45632, -42.0093, -41.55723, 
    -41.10036, -40.63895, -40.17321, -39.70337, -39.22964, -38.75225,
  -38.42853, -38.89363, -39.35483, -39.81194, -40.26473, -40.71301, 
    -41.15653, -41.59509, -42.02843, -42.45632, -42.87851, -43.29474, 
    -43.70475, -44.10828, -44.50503, -44.89474, -45.27712, -45.65187, 
    -46.0187, -46.37732, -46.72741, -47.06866, -47.40077, -47.72343, 
    -48.03632, -48.33913, -48.63155, -48.91327, -49.18397, -49.44336, 
    -49.69113, -49.927, -50.15067, -50.36186, -50.56031, -50.74577, 
    -50.91797, -51.0767, -51.22174, -51.35287, -51.46992, -51.57272, 
    -51.66111, -51.73498, -51.7942, -51.8387, -51.8684, -51.88326, -51.88326, 
    -51.8684, -51.8387, -51.7942, -51.73498, -51.66111, -51.57272, -51.46992, 
    -51.35287, -51.22174, -51.0767, -50.91797, -50.74577, -50.56031, 
    -50.36186, -50.15067, -49.927, -49.69113, -49.44336, -49.18397, 
    -48.91327, -48.63155, -48.33913, -48.03632, -47.72343, -47.40077, 
    -47.06866, -46.72741, -46.37732, -46.0187, -45.65187, -45.27712, 
    -44.89474, -44.50503, -44.10828, -43.70475, -43.29474, -42.87851, 
    -42.45632, -42.02843, -41.59509, -41.15653, -40.71301, -40.26473, 
    -39.81194, -39.35483, -38.89363, -38.42853,
  -38.09881, -38.55162, -39.00033, -39.44474, -39.88465, -40.31985, 
    -40.75014, -41.17529, -41.59509, -42.0093, -42.41769, -42.82002, 
    -43.21604, -43.60551, -43.98816, -44.36374, -44.73198, -45.0926, 
    -45.44535, -45.78994, -46.12609, -46.45353, -46.77196, -47.08112, 
    -47.3807, -47.67044, -47.95004, -48.21923, -48.47774, -48.72528, 
    -48.9616, -49.18642, -49.39951, -49.6006, -49.78946, -49.96586, 
    -50.12959, -50.28045, -50.41822, -50.54276, -50.65387, -50.75143, 
    -50.83531, -50.90538, -50.96155, -51.00375, -51.03191, -51.046, -51.046, 
    -51.03191, -51.00375, -50.96155, -50.90538, -50.83531, -50.75143, 
    -50.65387, -50.54276, -50.41822, -50.28045, -50.12959, -49.96586, 
    -49.78946, -49.6006, -49.39951, -49.18642, -48.9616, -48.72528, 
    -48.47774, -48.21923, -47.95004, -47.67044, -47.3807, -47.08112, 
    -46.77196, -46.45353, -46.12609, -45.78994, -45.44535, -45.0926, 
    -44.73198, -44.36374, -43.98816, -43.60551, -43.21604, -42.82002, 
    -42.41769, -42.0093, -41.59509, -41.17529, -40.75014, -40.31985, 
    -39.88465, -39.44474, -39.00033, -38.55162, -38.09881,
  -37.76321, -38.20377, -38.64002, -39.07178, -39.49888, -39.9211, -40.33826, 
    -40.75014, -41.15653, -41.55723, -41.95201, -42.34064, -42.7229, 
    -43.09856, -43.46738, -43.82911, -44.18351, -44.53034, -44.86935, 
    -45.20028, -45.52287, -45.83688, -46.14204, -46.43811, -46.72482, 
    -47.00192, -47.26916, -47.52629, -47.77305, -48.0092, -48.23452, 
    -48.44876, -48.6517, -48.84312, -49.02282, -49.19058, -49.34622, 
    -49.48956, -49.62043, -49.73867, -49.84415, -49.93674, -50.01631, 
    -50.08277, -50.13604, -50.17606, -50.20276, -50.21612, -50.21612, 
    -50.20276, -50.17606, -50.13604, -50.08277, -50.01631, -49.93674, 
    -49.84415, -49.73867, -49.62043, -49.48956, -49.34622, -49.19058, 
    -49.02282, -48.84312, -48.6517, -48.44876, -48.23452, -48.0092, 
    -47.77305, -47.52629, -47.26916, -47.00192, -46.72482, -46.43811, 
    -46.14204, -45.83688, -45.52287, -45.20028, -44.86935, -44.53034, 
    -44.18351, -43.82911, -43.46738, -43.09856, -42.7229, -42.34064, 
    -41.95201, -41.55723, -41.15653, -40.75014, -40.33826, -39.9211, 
    -39.49888, -39.07178, -38.64002, -38.20377, -37.76321,
  -37.42188, -37.8502, -38.27405, -38.69325, -39.10761, -39.51696, -39.9211, 
    -40.31985, -40.71301, -41.10036, -41.48173, -41.85689, -42.22562, 
    -42.58773, -42.94299, -43.29116, -43.63205, -43.9654, -44.29101, 
    -44.60864, -44.91806, -45.21903, -45.51133, -45.79473, -46.06899, 
    -46.33389, -46.5892, -46.83469, -47.07016, -47.29537, -47.51012, 
    -47.71421, -47.90744, -48.08961, -48.26053, -48.42004, -48.56796, 
    -48.70414, -48.82842, -48.94068, -49.04079, -49.12864, -49.20412, 
    -49.26716, -49.31768, -49.35562, -49.38094, -49.3936, -49.3936, 
    -49.38094, -49.35562, -49.31768, -49.26716, -49.20412, -49.12864, 
    -49.04079, -48.94068, -48.82842, -48.70414, -48.56796, -48.42004, 
    -48.26053, -48.08961, -47.90744, -47.71421, -47.51012, -47.29537, 
    -47.07016, -46.83469, -46.5892, -46.33389, -46.06899, -45.79473, 
    -45.51133, -45.21903, -44.91806, -44.60864, -44.29101, -43.9654, 
    -43.63205, -43.29116, -42.94299, -42.58773, -42.22562, -41.85689, 
    -41.48173, -41.10036, -40.71301, -40.31985, -39.9211, -39.51696, 
    -39.10761, -38.69325, -38.27405, -37.8502, -37.42188,
  -37.07492, -37.49107, -37.90258, -38.30929, -38.71102, -39.10761, 
    -39.49888, -39.88465, -40.26473, -40.63895, -41.00711, -41.36901, 
    -41.72447, -42.07329, -42.41526, -42.75019, -43.07787, -43.39809, 
    -43.71065, -44.01534, -44.31195, -44.60027, -44.88011, -45.15124, 
    -45.41347, -45.66659, -45.91039, -46.14469, -46.36929, -46.58398, 
    -46.7886, -46.98296, -47.16688, -47.34019, -47.50273, -47.65435, 
    -47.79491, -47.92425, -48.04226, -48.14882, -48.24382, -48.32716, 
    -48.39876, -48.45854, -48.50644, -48.54241, -48.56641, -48.57842, 
    -48.57842, -48.56641, -48.54241, -48.50644, -48.45854, -48.39876, 
    -48.32716, -48.24382, -48.14882, -48.04226, -47.92425, -47.79491, 
    -47.65435, -47.50273, -47.34019, -47.16688, -46.98296, -46.7886, 
    -46.58398, -46.36929, -46.14469, -45.91039, -45.66659, -45.41347, 
    -45.15124, -44.88011, -44.60027, -44.31195, -44.01534, -43.71065, 
    -43.39809, -43.07787, -42.75019, -42.41526, -42.07329, -41.72447, 
    -41.36901, -41.00711, -40.63895, -40.26473, -39.88465, -39.49888, 
    -39.10761, -38.71102, -38.30929, -37.90258, -37.49107, -37.07492,
  -36.72248, -37.12651, -37.52576, -37.92007, -38.30929, -38.69325, 
    -39.07178, -39.44474, -39.81194, -40.17321, -40.52837, -40.87727, 
    -41.2197, -41.5555, -41.88448, -42.20646, -42.52125, -42.82867, 
    -43.12852, -43.42064, -43.70482, -43.98088, -44.24864, -44.50792, 
    -44.75852, -45.00027, -45.23299, -45.45651, -45.67065, -45.87524, 
    -46.07014, -46.25516, -46.43016, -46.595, -46.74953, -46.89362, 
    -47.02713, -47.14996, -47.26199, -47.36312, -47.45325, -47.53231, 
    -47.6002, -47.65689, -47.7023, -47.7364, -47.75915, -47.77053, -47.77053, 
    -47.75915, -47.7364, -47.7023, -47.65689, -47.6002, -47.53231, -47.45325, 
    -47.36312, -47.26199, -47.14996, -47.02713, -46.89362, -46.74953, 
    -46.595, -46.43016, -46.25516, -46.07014, -45.87524, -45.67065, 
    -45.45651, -45.23299, -45.00027, -44.75852, -44.50792, -44.24864, 
    -43.98088, -43.70482, -43.42064, -43.12852, -42.82867, -42.52125, 
    -42.20646, -41.88448, -41.5555, -41.2197, -40.87727, -40.52837, 
    -40.17321, -39.81194, -39.44474, -39.07178, -38.69325, -38.30929, 
    -37.92007, -37.52576, -37.12651, -36.72248,
  -36.36466, -36.75665, -37.14373, -37.52576, -37.90258, -38.27405, 
    -38.64002, -39.00033, -39.35483, -39.70337, -40.04577, -40.38189, 
    -40.71156, -41.03462, -41.35089, -41.66023, -41.96246, -42.2574, 
    -42.54491, -42.82481, -43.09693, -43.36111, -43.61718, -43.86499, 
    -44.10437, -44.33515, -44.55719, -44.77034, -44.97443, -45.16932, 
    -45.35488, -45.53096, -45.69742, -45.85415, -46.00101, -46.13791, 
    -46.26471, -46.38132, -46.48764, -46.5836, -46.66909, -46.74407, 
    -46.80845, -46.86219, -46.90523, -46.93755, -46.95911, -46.96989, 
    -46.96989, -46.95911, -46.93755, -46.90523, -46.86219, -46.80845, 
    -46.74407, -46.66909, -46.5836, -46.48764, -46.38132, -46.26471, 
    -46.13791, -46.00101, -45.85415, -45.69742, -45.53096, -45.35488, 
    -45.16932, -44.97443, -44.77034, -44.55719, -44.33515, -44.10437, 
    -43.86499, -43.61718, -43.36111, -43.09693, -42.82481, -42.54491, 
    -42.2574, -41.96246, -41.66023, -41.35089, -41.03462, -40.71156, 
    -40.38189, -40.04577, -39.70337, -39.35483, -39.00033, -38.64002, 
    -38.27405, -37.90258, -37.52576, -37.14373, -36.75665, -36.36466,
  -36.0016, -36.38164, -36.75665, -37.12651, -37.49107, -37.8502, -38.20377, 
    -38.55162, -38.89363, -39.22964, -39.55952, -39.88312, -40.20029, 
    -40.51088, -40.81476, -41.11176, -41.40174, -41.68456, -41.96006, 
    -42.2281, -42.48852, -42.74119, -42.98596, -43.22269, -43.45123, 
    -43.67144, -43.8832, -44.08636, -44.28079, -44.46637, -44.64297, 
    -44.81047, -44.96877, -45.11773, -45.25727, -45.38729, -45.50768, 
    -45.61835, -45.71924, -45.81026, -45.89135, -45.96243, -46.02346, 
    -46.07439, -46.11519, -46.14581, -46.16624, -46.17646, -46.17646, 
    -46.16624, -46.14581, -46.11519, -46.07439, -46.02346, -45.96243, 
    -45.89135, -45.81026, -45.71924, -45.61835, -45.50768, -45.38729, 
    -45.25727, -45.11773, -44.96877, -44.81047, -44.64297, -44.46637, 
    -44.28079, -44.08636, -43.8832, -43.67144, -43.45123, -43.22269, 
    -42.98596, -42.74119, -42.48852, -42.2281, -41.96006, -41.68456, 
    -41.40174, -41.11176, -40.81476, -40.51088, -40.20029, -39.88312, 
    -39.55952, -39.22964, -38.89363, -38.55162, -38.20377, -37.8502, 
    -37.49107, -37.12651, -36.75665, -36.38164, -36.0016,
  -35.63342, -36.0016, -36.36466, -36.72248, -37.07492, -37.42188, -37.76321, 
    -38.09881, -38.42853, -38.75225, -39.06984, -39.38117, -39.68611, 
    -39.98453, -40.27629, -40.56128, -40.83934, -41.11036, -41.37419, 
    -41.63073, -41.87982, -42.12135, -42.35519, -42.58122, -42.7993, 
    -43.00933, -43.21118, -43.40474, -43.58989, -43.76653, -43.93454, 
    -44.09382, -44.24429, -44.38583, -44.51836, -44.64181, -44.75608, 
    -44.8611, -44.9568, -45.04311, -45.11999, -45.18737, -45.24522, 
    -45.29348, -45.33213, -45.36115, -45.3805, -45.39018, -45.39018, 
    -45.3805, -45.36115, -45.33213, -45.29348, -45.24522, -45.18737, 
    -45.11999, -45.04311, -44.9568, -44.8611, -44.75608, -44.64181, 
    -44.51836, -44.38583, -44.24429, -44.09382, -43.93454, -43.76653, 
    -43.58989, -43.40474, -43.21118, -43.00933, -42.7993, -42.58122, 
    -42.35519, -42.12135, -41.87982, -41.63073, -41.37419, -41.11036, 
    -40.83934, -40.56128, -40.27629, -39.98453, -39.68611, -39.38117, 
    -39.06984, -38.75225, -38.42853, -38.09881, -37.76321, -37.42188, 
    -37.07492, -36.72248, -36.36466, -36.0016, -35.63342 ;

 area =
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.158754e+09, 7.321026e+09, 7.485062e+09, 7.650767e+09, 7.818037e+09, 
    7.986756e+09, 8.156796e+09, 8.32802e+09, 8.500278e+09, 8.673409e+09, 
    8.84724e+09, 9.021585e+09, 9.196247e+09, 9.371016e+09, 9.54567e+09, 
    9.719975e+09, 9.893683e+09, 1.006654e+10, 1.023827e+10, 1.040861e+10, 
    1.057725e+10, 1.07439e+10, 1.090825e+10, 1.106999e+10, 1.122879e+10, 
    1.138432e+10, 1.153626e+10, 1.168427e+10, 1.1828e+10, 1.196713e+10, 
    1.210132e+10, 1.223023e+10, 1.235355e+10, 1.247093e+10, 1.258209e+10, 
    1.268671e+10, 1.27845e+10, 1.287519e+10, 1.295852e+10, 1.303425e+10, 
    1.310215e+10, 1.316203e+10, 1.32137e+10, 1.3257e+10, 1.32918e+10, 
    1.3318e+10, 1.333551e+10, 1.334428e+10, 1.334428e+10, 1.333551e+10, 
    1.3318e+10, 1.32918e+10, 1.3257e+10, 1.32137e+10, 1.316203e+10, 
    1.310215e+10, 1.303425e+10, 1.295852e+10, 1.287519e+10, 1.27845e+10, 
    1.268671e+10, 1.258209e+10, 1.247093e+10, 1.235355e+10, 1.223023e+10, 
    1.210132e+10, 1.196713e+10, 1.1828e+10, 1.168427e+10, 1.153626e+10, 
    1.138432e+10, 1.122879e+10, 1.106999e+10, 1.090825e+10, 1.07439e+10, 
    1.057725e+10, 1.040861e+10, 1.023827e+10, 1.006654e+10, 9.893683e+09, 
    9.719975e+09, 9.54567e+09, 9.371016e+09, 9.196247e+09, 9.021585e+09, 
    8.84724e+09, 8.673409e+09, 8.500278e+09, 8.32802e+09, 8.156796e+09, 
    7.986756e+09, 7.818037e+09, 7.650767e+09, 7.485062e+09, 7.321026e+09, 
    7.158754e+09,
  7.157529e+09, 7.319673e+09, 7.483577e+09, 7.649145e+09, 7.816271e+09, 
    7.984841e+09, 8.154726e+09, 8.32579e+09, 8.497883e+09, 8.670843e+09, 
    8.844498e+09, 9.018663e+09, 9.193139e+09, 9.367718e+09, 9.542177e+09, 
    9.716282e+09, 9.88979e+09, 1.006244e+10, 1.023397e+10, 1.040409e+10, 
    1.057252e+10, 1.073895e+10, 1.090309e+10, 1.106461e+10, 1.12232e+10, 
    1.137852e+10, 1.153025e+10, 1.167804e+10, 1.182158e+10, 1.19605e+10, 
    1.209449e+10, 1.222321e+10, 1.234634e+10, 1.246355e+10, 1.257453e+10, 
    1.267899e+10, 1.277663e+10, 1.286718e+10, 1.295038e+10, 1.302599e+10, 
    1.309378e+10, 1.315356e+10, 1.320514e+10, 1.324837e+10, 1.328312e+10, 
    1.330927e+10, 1.332675e+10, 1.333551e+10, 1.333551e+10, 1.332675e+10, 
    1.330927e+10, 1.328312e+10, 1.324837e+10, 1.320514e+10, 1.315356e+10, 
    1.309378e+10, 1.302599e+10, 1.295038e+10, 1.286718e+10, 1.277663e+10, 
    1.267899e+10, 1.257453e+10, 1.246355e+10, 1.234634e+10, 1.222321e+10, 
    1.209449e+10, 1.19605e+10, 1.182158e+10, 1.167804e+10, 1.153025e+10, 
    1.137852e+10, 1.12232e+10, 1.106461e+10, 1.090309e+10, 1.073895e+10, 
    1.057252e+10, 1.040409e+10, 1.023397e+10, 1.006244e+10, 9.88979e+09, 
    9.716282e+09, 9.542177e+09, 9.367718e+09, 9.193139e+09, 9.018663e+09, 
    8.844498e+09, 8.670843e+09, 8.497883e+09, 8.32579e+09, 8.154726e+09, 
    7.984841e+09, 7.816271e+09, 7.649145e+09, 7.483577e+09, 7.319673e+09, 
    7.157529e+09,
  7.155078e+09, 7.316969e+09, 7.480609e+09, 7.645901e+09, 7.812741e+09, 
    7.981012e+09, 8.150589e+09, 8.321333e+09, 8.493095e+09, 8.665715e+09, 
    8.839017e+09, 9.012821e+09, 9.186927e+09, 9.361125e+09, 9.535196e+09, 
    9.708905e+09, 9.882009e+09, 1.005425e+10, 1.022536e+10, 1.039506e+10, 
    1.056306e+10, 1.072907e+10, 1.089278e+10, 1.105388e+10, 1.121203e+10, 
    1.136693e+10, 1.151823e+10, 1.166561e+10, 1.180873e+10, 1.194726e+10, 
    1.208085e+10, 1.220919e+10, 1.233195e+10, 1.24488e+10, 1.255944e+10, 
    1.266358e+10, 1.276091e+10, 1.285118e+10, 1.293411e+10, 1.300948e+10, 
    1.307706e+10, 1.313664e+10, 1.318806e+10, 1.323115e+10, 1.326578e+10, 
    1.329185e+10, 1.330927e+10, 1.3318e+10, 1.3318e+10, 1.330927e+10, 
    1.329185e+10, 1.326578e+10, 1.323115e+10, 1.318806e+10, 1.313664e+10, 
    1.307706e+10, 1.300948e+10, 1.293411e+10, 1.285118e+10, 1.276091e+10, 
    1.266358e+10, 1.255944e+10, 1.24488e+10, 1.233195e+10, 1.220919e+10, 
    1.208085e+10, 1.194726e+10, 1.180873e+10, 1.166561e+10, 1.151823e+10, 
    1.136693e+10, 1.121203e+10, 1.105388e+10, 1.089278e+10, 1.072907e+10, 
    1.056306e+10, 1.039506e+10, 1.022536e+10, 1.005425e+10, 9.882009e+09, 
    9.708905e+09, 9.535196e+09, 9.361125e+09, 9.186927e+09, 9.012821e+09, 
    8.839017e+09, 8.665715e+09, 8.493095e+09, 8.321333e+09, 8.150589e+09, 
    7.981012e+09, 7.812741e+09, 7.645901e+09, 7.480609e+09, 7.316969e+09, 
    7.155078e+09,
  7.151404e+09, 7.312915e+09, 7.476158e+09, 7.641037e+09, 7.807448e+09, 
    7.975273e+09, 8.144387e+09, 8.314652e+09, 8.485919e+09, 8.658028e+09, 
    8.830806e+09, 9.004068e+09, 9.177618e+09, 9.351248e+09, 9.524738e+09, 
    9.697854e+09, 9.870353e+09, 1.004198e+10, 1.021247e+10, 1.038154e+10, 
    1.054891e+10, 1.071428e+10, 1.087735e+10, 1.10378e+10, 1.119532e+10, 
    1.134958e+10, 1.150025e+10, 1.164701e+10, 1.178951e+10, 1.192743e+10, 
    1.206044e+10, 1.218821e+10, 1.231041e+10, 1.242673e+10, 1.253687e+10, 
    1.264052e+10, 1.273739e+10, 1.282723e+10, 1.290977e+10, 1.298478e+10, 
    1.305203e+10, 1.311133e+10, 1.316249e+10, 1.320537e+10, 1.323984e+10, 
    1.326578e+10, 1.328312e+10, 1.32918e+10, 1.32918e+10, 1.328312e+10, 
    1.326578e+10, 1.323984e+10, 1.320537e+10, 1.316249e+10, 1.311133e+10, 
    1.305203e+10, 1.298478e+10, 1.290977e+10, 1.282723e+10, 1.273739e+10, 
    1.264052e+10, 1.253687e+10, 1.242673e+10, 1.231041e+10, 1.218821e+10, 
    1.206044e+10, 1.192743e+10, 1.178951e+10, 1.164701e+10, 1.150025e+10, 
    1.134958e+10, 1.119532e+10, 1.10378e+10, 1.087735e+10, 1.071428e+10, 
    1.054891e+10, 1.038154e+10, 1.021247e+10, 1.004198e+10, 9.870353e+09, 
    9.697854e+09, 9.524738e+09, 9.351248e+09, 9.177618e+09, 9.004068e+09, 
    8.830806e+09, 8.658028e+09, 8.485919e+09, 8.314652e+09, 8.144387e+09, 
    7.975273e+09, 7.807448e+09, 7.641037e+09, 7.476158e+09, 7.312915e+09, 
    7.151404e+09,
  7.146505e+09, 7.307511e+09, 7.470226e+09, 7.634556e+09, 7.800395e+09, 
    7.967627e+09, 8.136126e+09, 8.305754e+09, 8.476363e+09, 8.647793e+09, 
    8.819871e+09, 8.992415e+09, 9.165227e+09, 9.338102e+09, 9.510819e+09, 
    9.683147e+09, 9.854844e+09, 1.002566e+10, 1.019532e+10, 1.036355e+10, 
    1.053008e+10, 1.06946e+10, 1.085682e+10, 1.101642e+10, 1.117309e+10, 
    1.13265e+10, 1.147634e+10, 1.162227e+10, 1.176396e+10, 1.190108e+10, 
    1.203331e+10, 1.216031e+10, 1.228178e+10, 1.23974e+10, 1.250686e+10, 
    1.260987e+10, 1.270614e+10, 1.279542e+10, 1.287743e+10, 1.295196e+10, 
    1.301878e+10, 1.30777e+10, 1.312854e+10, 1.317114e+10, 1.320537e+10, 
    1.323115e+10, 1.324837e+10, 1.3257e+10, 1.3257e+10, 1.324837e+10, 
    1.323115e+10, 1.320537e+10, 1.317114e+10, 1.312854e+10, 1.30777e+10, 
    1.301878e+10, 1.295196e+10, 1.287743e+10, 1.279542e+10, 1.270614e+10, 
    1.260987e+10, 1.250686e+10, 1.23974e+10, 1.228178e+10, 1.216031e+10, 
    1.203331e+10, 1.190108e+10, 1.176396e+10, 1.162227e+10, 1.147634e+10, 
    1.13265e+10, 1.117309e+10, 1.101642e+10, 1.085682e+10, 1.06946e+10, 
    1.053008e+10, 1.036355e+10, 1.019532e+10, 1.002566e+10, 9.854844e+09, 
    9.683147e+09, 9.510819e+09, 9.338102e+09, 9.165227e+09, 8.992415e+09, 
    8.819871e+09, 8.647793e+09, 8.476363e+09, 8.305754e+09, 8.136126e+09, 
    7.967627e+09, 7.800395e+09, 7.634556e+09, 7.470226e+09, 7.307511e+09, 
    7.146505e+09,
  7.140384e+09, 7.30076e+09, 7.462817e+09, 7.626462e+09, 7.791588e+09, 
    7.958081e+09, 8.125813e+09, 8.294647e+09, 8.464436e+09, 8.63502e+09, 
    8.806228e+09, 8.977876e+09, 9.14977e+09, 9.321703e+09, 9.49346e+09, 
    9.664807e+09, 9.835507e+09, 1.00053e+10, 1.017394e+10, 1.034114e+10, 
    1.050662e+10, 1.067009e+10, 1.083124e+10, 1.098979e+10, 1.11454e+10, 
    1.129776e+10, 1.144656e+10, 1.159146e+10, 1.173213e+10, 1.186826e+10, 
    1.199952e+10, 1.212559e+10, 1.224615e+10, 1.236089e+10, 1.246951e+10, 
    1.257172e+10, 1.266725e+10, 1.275582e+10, 1.283719e+10, 1.291113e+10, 
    1.297741e+10, 1.303585e+10, 1.308628e+10, 1.312854e+10, 1.316249e+10, 
    1.318806e+10, 1.320514e+10, 1.32137e+10, 1.32137e+10, 1.320514e+10, 
    1.318806e+10, 1.316249e+10, 1.312854e+10, 1.308628e+10, 1.303585e+10, 
    1.297741e+10, 1.291113e+10, 1.283719e+10, 1.275582e+10, 1.266725e+10, 
    1.257172e+10, 1.246951e+10, 1.236089e+10, 1.224615e+10, 1.212559e+10, 
    1.199952e+10, 1.186826e+10, 1.173213e+10, 1.159146e+10, 1.144656e+10, 
    1.129776e+10, 1.11454e+10, 1.098979e+10, 1.083124e+10, 1.067009e+10, 
    1.050662e+10, 1.034114e+10, 1.017394e+10, 1.00053e+10, 9.835507e+09, 
    9.664807e+09, 9.49346e+09, 9.321703e+09, 9.14977e+09, 8.977876e+09, 
    8.806228e+09, 8.63502e+09, 8.464436e+09, 8.294647e+09, 8.125813e+09, 
    7.958081e+09, 7.791588e+09, 7.626462e+09, 7.462817e+09, 7.30076e+09, 
    7.140384e+09,
  7.133041e+09, 7.292662e+09, 7.453934e+09, 7.616759e+09, 7.781033e+09, 
    7.946641e+09, 8.113456e+09, 8.281342e+09, 8.450151e+09, 8.619724e+09, 
    8.789891e+09, 8.96047e+09, 9.131267e+09, 9.302078e+09, 9.472687e+09, 
    9.642865e+09, 9.812372e+09, 9.980962e+09, 1.014837e+10, 1.031433e+10, 
    1.047856e+10, 1.064077e+10, 1.080067e+10, 1.095795e+10, 1.111231e+10, 
    1.126342e+10, 1.141097e+10, 1.155465e+10, 1.169412e+10, 1.182907e+10, 
    1.195917e+10, 1.208412e+10, 1.220359e+10, 1.231729e+10, 1.242492e+10, 
    1.252618e+10, 1.262082e+10, 1.270856e+10, 1.278916e+10, 1.286239e+10, 
    1.292804e+10, 1.298592e+10, 1.303585e+10, 1.30777e+10, 1.311133e+10, 
    1.313664e+10, 1.315356e+10, 1.316203e+10, 1.316203e+10, 1.315356e+10, 
    1.313664e+10, 1.311133e+10, 1.30777e+10, 1.303585e+10, 1.298592e+10, 
    1.292804e+10, 1.286239e+10, 1.278916e+10, 1.270856e+10, 1.262082e+10, 
    1.252618e+10, 1.242492e+10, 1.231729e+10, 1.220359e+10, 1.208412e+10, 
    1.195917e+10, 1.182907e+10, 1.169412e+10, 1.155465e+10, 1.141097e+10, 
    1.126342e+10, 1.111231e+10, 1.095795e+10, 1.080067e+10, 1.064077e+10, 
    1.047856e+10, 1.031433e+10, 1.014837e+10, 9.980962e+09, 9.812372e+09, 
    9.642865e+09, 9.472687e+09, 9.302078e+09, 9.131267e+09, 8.96047e+09, 
    8.789891e+09, 8.619724e+09, 8.450151e+09, 8.281342e+09, 8.113456e+09, 
    7.946641e+09, 7.781033e+09, 7.616759e+09, 7.453934e+09, 7.292662e+09, 
    7.133041e+09,
  7.124479e+09, 7.283223e+09, 7.443579e+09, 7.605452e+09, 7.768736e+09, 
    7.933316e+09, 8.099066e+09, 8.26585e+09, 8.433522e+09, 8.601922e+09, 
    8.770882e+09, 8.940219e+09, 9.109745e+09, 9.279254e+09, 9.448532e+09, 
    9.617354e+09, 9.785482e+09, 9.95267e+09, 1.011866e+10, 1.028319e+10, 
    1.044597e+10, 1.060673e+10, 1.076517e+10, 1.092099e+10, 1.107389e+10, 
    1.122356e+10, 1.136968e+10, 1.151193e+10, 1.165001e+10, 1.17836e+10, 
    1.191237e+10, 1.203602e+10, 1.215424e+10, 1.226673e+10, 1.237321e+10, 
    1.247338e+10, 1.256699e+10, 1.265377e+10, 1.273348e+10, 1.280589e+10, 
    1.287081e+10, 1.292804e+10, 1.297741e+10, 1.301878e+10, 1.305203e+10, 
    1.307706e+10, 1.309378e+10, 1.310215e+10, 1.310215e+10, 1.309378e+10, 
    1.307706e+10, 1.305203e+10, 1.301878e+10, 1.297741e+10, 1.292804e+10, 
    1.287081e+10, 1.280589e+10, 1.273348e+10, 1.265377e+10, 1.256699e+10, 
    1.247338e+10, 1.237321e+10, 1.226673e+10, 1.215424e+10, 1.203602e+10, 
    1.191237e+10, 1.17836e+10, 1.165001e+10, 1.151193e+10, 1.136968e+10, 
    1.122356e+10, 1.107389e+10, 1.092099e+10, 1.076517e+10, 1.060673e+10, 
    1.044597e+10, 1.028319e+10, 1.011866e+10, 9.95267e+09, 9.785482e+09, 
    9.617354e+09, 9.448532e+09, 9.279254e+09, 9.109745e+09, 8.940219e+09, 
    8.770882e+09, 8.601922e+09, 8.433522e+09, 8.26585e+09, 8.099066e+09, 
    7.933316e+09, 7.768736e+09, 7.605452e+09, 7.443579e+09, 7.283223e+09, 
    7.124479e+09,
  7.1147e+09, 7.272444e+09, 7.431758e+09, 7.592547e+09, 7.754704e+09, 
    7.918115e+09, 8.082655e+09, 8.248187e+09, 8.414565e+09, 8.581632e+09, 
    8.749221e+09, 8.917151e+09, 9.085231e+09, 9.253263e+09, 9.421031e+09, 
    9.588315e+09, 9.754878e+09, 9.920478e+09, 1.008486e+10, 1.024776e+10, 
    1.040891e+10, 1.056802e+10, 1.07248e+10, 1.087898e+10, 1.103023e+10, 
    1.117826e+10, 1.132276e+10, 1.146341e+10, 1.159992e+10, 1.173195e+10, 
    1.185922e+10, 1.198141e+10, 1.209821e+10, 1.220935e+10, 1.231452e+10, 
    1.241347e+10, 1.250591e+10, 1.25916e+10, 1.267031e+10, 1.27418e+10, 
    1.280589e+10, 1.286239e+10, 1.291113e+10, 1.295196e+10, 1.298478e+10, 
    1.300948e+10, 1.302599e+10, 1.303425e+10, 1.303425e+10, 1.302599e+10, 
    1.300948e+10, 1.298478e+10, 1.295196e+10, 1.291113e+10, 1.286239e+10, 
    1.280589e+10, 1.27418e+10, 1.267031e+10, 1.25916e+10, 1.250591e+10, 
    1.241347e+10, 1.231452e+10, 1.220935e+10, 1.209821e+10, 1.198141e+10, 
    1.185922e+10, 1.173195e+10, 1.159992e+10, 1.146341e+10, 1.132276e+10, 
    1.117826e+10, 1.103023e+10, 1.087898e+10, 1.07248e+10, 1.056802e+10, 
    1.040891e+10, 1.024776e+10, 1.008486e+10, 9.920478e+09, 9.754878e+09, 
    9.588315e+09, 9.421031e+09, 9.253263e+09, 9.085231e+09, 8.917151e+09, 
    8.749221e+09, 8.581632e+09, 8.414565e+09, 8.248187e+09, 8.082655e+09, 
    7.918115e+09, 7.754704e+09, 7.592547e+09, 7.431758e+09, 7.272444e+09, 
    7.1147e+09,
  7.103705e+09, 7.260329e+09, 7.418477e+09, 7.578052e+09, 7.738948e+09, 
    7.901051e+09, 8.064236e+09, 8.228367e+09, 8.3933e+09, 8.558878e+09, 
    8.724934e+09, 8.891291e+09, 9.05776e+09, 9.224142e+09, 9.390226e+09, 
    9.555794e+09, 9.720613e+09, 9.884442e+09, 1.004703e+10, 1.020812e+10, 
    1.036744e+10, 1.052472e+10, 1.067967e+10, 1.0832e+10, 1.098142e+10, 
    1.112763e+10, 1.127033e+10, 1.14092e+10, 1.154395e+10, 1.167428e+10, 
    1.179987e+10, 1.192043e+10, 1.203567e+10, 1.214529e+10, 1.224902e+10, 
    1.234659e+10, 1.243775e+10, 1.252223e+10, 1.259983e+10, 1.267031e+10, 
    1.273348e+10, 1.278916e+10, 1.283719e+10, 1.287743e+10, 1.290977e+10, 
    1.293411e+10, 1.295038e+10, 1.295852e+10, 1.295852e+10, 1.295038e+10, 
    1.293411e+10, 1.290977e+10, 1.287743e+10, 1.283719e+10, 1.278916e+10, 
    1.273348e+10, 1.267031e+10, 1.259983e+10, 1.252223e+10, 1.243775e+10, 
    1.234659e+10, 1.224902e+10, 1.214529e+10, 1.203567e+10, 1.192043e+10, 
    1.179987e+10, 1.167428e+10, 1.154395e+10, 1.14092e+10, 1.127033e+10, 
    1.112763e+10, 1.098142e+10, 1.0832e+10, 1.067967e+10, 1.052472e+10, 
    1.036744e+10, 1.020812e+10, 1.004703e+10, 9.884442e+09, 9.720613e+09, 
    9.555794e+09, 9.390226e+09, 9.224142e+09, 9.05776e+09, 8.891291e+09, 
    8.724934e+09, 8.558878e+09, 8.3933e+09, 8.228367e+09, 8.064236e+09, 
    7.901051e+09, 7.738948e+09, 7.578052e+09, 7.418477e+09, 7.260329e+09, 
    7.103705e+09,
  7.091497e+09, 7.246883e+09, 7.403741e+09, 7.561974e+09, 7.721477e+09, 
    7.882135e+09, 8.043825e+09, 8.20641e+09, 8.369748e+09, 8.533684e+09, 
    8.698051e+09, 8.862674e+09, 9.027367e+09, 9.191932e+09, 9.356163e+09, 
    9.519842e+09, 9.68274e+09, 9.844622e+09, 1.000524e+10, 1.016434e+10, 
    1.032166e+10, 1.047692e+10, 1.062985e+10, 1.078017e+10, 1.092757e+10, 
    1.107179e+10, 1.12125e+10, 1.134943e+10, 1.148226e+10, 1.16107e+10, 
    1.173446e+10, 1.185324e+10, 1.196675e+10, 1.207473e+10, 1.217688e+10, 
    1.227295e+10, 1.236269e+10, 1.244586e+10, 1.252223e+10, 1.25916e+10, 
    1.265377e+10, 1.270856e+10, 1.275582e+10, 1.279542e+10, 1.282723e+10, 
    1.285118e+10, 1.286718e+10, 1.287519e+10, 1.287519e+10, 1.286718e+10, 
    1.285118e+10, 1.282723e+10, 1.279542e+10, 1.275582e+10, 1.270856e+10, 
    1.265377e+10, 1.25916e+10, 1.252223e+10, 1.244586e+10, 1.236269e+10, 
    1.227295e+10, 1.217688e+10, 1.207473e+10, 1.196675e+10, 1.185324e+10, 
    1.173446e+10, 1.16107e+10, 1.148226e+10, 1.134943e+10, 1.12125e+10, 
    1.107179e+10, 1.092757e+10, 1.078017e+10, 1.062985e+10, 1.047692e+10, 
    1.032166e+10, 1.016434e+10, 1.000524e+10, 9.844622e+09, 9.68274e+09, 
    9.519842e+09, 9.356163e+09, 9.191932e+09, 9.027367e+09, 8.862674e+09, 
    8.698051e+09, 8.533684e+09, 8.369748e+09, 8.20641e+09, 8.043825e+09, 
    7.882135e+09, 7.721477e+09, 7.561974e+09, 7.403741e+09, 7.246883e+09, 
    7.091497e+09,
  7.078078e+09, 7.23211e+09, 7.387556e+09, 7.544322e+09, 7.702302e+09, 
    7.861382e+09, 8.021437e+09, 8.182336e+09, 8.343933e+09, 8.506077e+09, 
    8.668601e+09, 8.831335e+09, 8.994092e+09, 9.156679e+09, 9.318892e+09, 
    9.480515e+09, 9.641325e+09, 9.801088e+09, 9.959563e+09, 1.01165e+10, 
    1.027164e+10, 1.042471e+10, 1.057545e+10, 1.072358e+10, 1.08688e+10, 
    1.101085e+10, 1.114942e+10, 1.128423e+10, 1.141498e+10, 1.154138e+10, 
    1.166315e+10, 1.178001e+10, 1.189166e+10, 1.199784e+10, 1.209829e+10, 
    1.219274e+10, 1.228095e+10, 1.236269e+10, 1.243775e+10, 1.250591e+10, 
    1.256699e+10, 1.262082e+10, 1.266725e+10, 1.270614e+10, 1.273739e+10, 
    1.276091e+10, 1.277663e+10, 1.27845e+10, 1.27845e+10, 1.277663e+10, 
    1.276091e+10, 1.273739e+10, 1.270614e+10, 1.266725e+10, 1.262082e+10, 
    1.256699e+10, 1.250591e+10, 1.243775e+10, 1.236269e+10, 1.228095e+10, 
    1.219274e+10, 1.209829e+10, 1.199784e+10, 1.189166e+10, 1.178001e+10, 
    1.166315e+10, 1.154138e+10, 1.141498e+10, 1.128423e+10, 1.114942e+10, 
    1.101085e+10, 1.08688e+10, 1.072358e+10, 1.057545e+10, 1.042471e+10, 
    1.027164e+10, 1.01165e+10, 9.959563e+09, 9.801088e+09, 9.641325e+09, 
    9.480515e+09, 9.318892e+09, 9.156679e+09, 8.994092e+09, 8.831335e+09, 
    8.668601e+09, 8.506077e+09, 8.343933e+09, 8.182336e+09, 8.021437e+09, 
    7.861382e+09, 7.702302e+09, 7.544322e+09, 7.387556e+09, 7.23211e+09, 
    7.078078e+09,
  7.063453e+09, 7.216014e+09, 7.36993e+09, 7.525106e+09, 7.681435e+09, 
    7.838806e+09, 7.997093e+09, 8.156166e+09, 8.31588e+09, 8.476086e+09, 
    8.636621e+09, 8.797313e+09, 8.95798e+09, 9.118431e+09, 9.278465e+09, 
    9.437871e+09, 9.596429e+09, 9.753911e+09, 9.910078e+09, 1.006469e+10, 
    1.021748e+10, 1.03682e+10, 1.051658e+10, 1.066235e+10, 1.080523e+10, 
    1.094495e+10, 1.108122e+10, 1.121375e+10, 1.134227e+10, 1.146649e+10, 
    1.158613e+10, 1.170091e+10, 1.181057e+10, 1.191483e+10, 1.201345e+10, 
    1.210616e+10, 1.219274e+10, 1.227295e+10, 1.234659e+10, 1.241347e+10, 
    1.247338e+10, 1.252618e+10, 1.257172e+10, 1.260987e+10, 1.264052e+10, 
    1.266358e+10, 1.267899e+10, 1.268671e+10, 1.268671e+10, 1.267899e+10, 
    1.266358e+10, 1.264052e+10, 1.260987e+10, 1.257172e+10, 1.252618e+10, 
    1.247338e+10, 1.241347e+10, 1.234659e+10, 1.227295e+10, 1.219274e+10, 
    1.210616e+10, 1.201345e+10, 1.191483e+10, 1.181057e+10, 1.170091e+10, 
    1.158613e+10, 1.146649e+10, 1.134227e+10, 1.121375e+10, 1.108122e+10, 
    1.094495e+10, 1.080523e+10, 1.066235e+10, 1.051658e+10, 1.03682e+10, 
    1.021748e+10, 1.006469e+10, 9.910078e+09, 9.753911e+09, 9.596429e+09, 
    9.437871e+09, 9.278465e+09, 9.118431e+09, 8.95798e+09, 8.797313e+09, 
    8.636621e+09, 8.476086e+09, 8.31588e+09, 8.156166e+09, 7.997093e+09, 
    7.838806e+09, 7.681435e+09, 7.525106e+09, 7.36993e+09, 7.216014e+09, 
    7.063453e+09,
  7.047623e+09, 7.198601e+09, 7.350871e+09, 7.504335e+09, 7.65889e+09, 
    7.814423e+09, 7.970811e+09, 8.127923e+09, 8.285618e+09, 8.443745e+09, 
    8.602145e+09, 8.760649e+09, 8.919077e+09, 9.077242e+09, 9.234944e+09, 
    9.391978e+09, 9.548129e+09, 9.703171e+09, 9.856871e+09, 1.000899e+10, 
    1.015928e+10, 1.030749e+10, 1.045336e+10, 1.059662e+10, 1.0737e+10, 
    1.087423e+10, 1.100805e+10, 1.113816e+10, 1.12643e+10, 1.13862e+10, 
    1.150357e+10, 1.161615e+10, 1.172369e+10, 1.182591e+10, 1.192258e+10, 
    1.201345e+10, 1.209829e+10, 1.217688e+10, 1.224902e+10, 1.231452e+10, 
    1.237321e+10, 1.242492e+10, 1.246951e+10, 1.250686e+10, 1.253687e+10, 
    1.255944e+10, 1.257453e+10, 1.258209e+10, 1.258209e+10, 1.257453e+10, 
    1.255944e+10, 1.253687e+10, 1.250686e+10, 1.246951e+10, 1.242492e+10, 
    1.237321e+10, 1.231452e+10, 1.224902e+10, 1.217688e+10, 1.209829e+10, 
    1.201345e+10, 1.192258e+10, 1.182591e+10, 1.172369e+10, 1.161615e+10, 
    1.150357e+10, 1.13862e+10, 1.12643e+10, 1.113816e+10, 1.100805e+10, 
    1.087423e+10, 1.0737e+10, 1.059662e+10, 1.045336e+10, 1.030749e+10, 
    1.015928e+10, 1.000899e+10, 9.856871e+09, 9.703171e+09, 9.548129e+09, 
    9.391978e+09, 9.234944e+09, 9.077242e+09, 8.919077e+09, 8.760649e+09, 
    8.602145e+09, 8.443745e+09, 8.285618e+09, 8.127923e+09, 7.970811e+09, 
    7.814423e+09, 7.65889e+09, 7.504335e+09, 7.350871e+09, 7.198601e+09, 
    7.047623e+09,
  7.030593e+09, 7.179877e+09, 7.330385e+09, 7.482021e+09, 7.634681e+09, 
    7.788252e+09, 7.942612e+09, 8.097633e+09, 8.253174e+09, 8.409087e+09, 
    8.565214e+09, 8.721389e+09, 8.877434e+09, 9.033167e+09, 9.188391e+09, 
    9.342905e+09, 9.496498e+09, 9.64895e+09, 9.800034e+09, 9.949515e+09, 
    1.009715e+10, 1.02427e+10, 1.03859e+10, 1.05265e+10, 1.066424e+10, 
    1.079885e+10, 1.093007e+10, 1.105763e+10, 1.118125e+10, 1.130069e+10, 
    1.141567e+10, 1.152593e+10, 1.163122e+10, 1.17313e+10, 1.182591e+10, 
    1.191483e+10, 1.199784e+10, 1.207473e+10, 1.214529e+10, 1.220935e+10, 
    1.226673e+10, 1.231729e+10, 1.236089e+10, 1.23974e+10, 1.242673e+10, 
    1.24488e+10, 1.246355e+10, 1.247093e+10, 1.247093e+10, 1.246355e+10, 
    1.24488e+10, 1.242673e+10, 1.23974e+10, 1.236089e+10, 1.231729e+10, 
    1.226673e+10, 1.220935e+10, 1.214529e+10, 1.207473e+10, 1.199784e+10, 
    1.191483e+10, 1.182591e+10, 1.17313e+10, 1.163122e+10, 1.152593e+10, 
    1.141567e+10, 1.130069e+10, 1.118125e+10, 1.105763e+10, 1.093007e+10, 
    1.079885e+10, 1.066424e+10, 1.05265e+10, 1.03859e+10, 1.02427e+10, 
    1.009715e+10, 9.949515e+09, 9.800034e+09, 9.64895e+09, 9.496498e+09, 
    9.342905e+09, 9.188391e+09, 9.033167e+09, 8.877434e+09, 8.721389e+09, 
    8.565214e+09, 8.409087e+09, 8.253174e+09, 8.097633e+09, 7.942612e+09, 
    7.788252e+09, 7.634681e+09, 7.482021e+09, 7.330385e+09, 7.179877e+09, 
    7.030593e+09,
  7.012366e+09, 7.159848e+09, 7.308484e+09, 7.458176e+09, 7.608822e+09, 
    7.760311e+09, 7.912521e+09, 8.065324e+09, 8.218582e+09, 8.372148e+09, 
    8.525868e+09, 8.679578e+09, 8.833104e+09, 8.986266e+09, 9.138871e+09, 
    9.290724e+09, 9.441618e+09, 9.591338e+09, 9.739662e+09, 9.886363e+09, 
    1.00312e+10, 1.017395e+10, 1.031435e+10, 1.045215e+10, 1.058711e+10, 
    1.071896e+10, 1.084745e+10, 1.097232e+10, 1.109331e+10, 1.121017e+10, 
    1.132264e+10, 1.143046e+10, 1.153341e+10, 1.163122e+10, 1.172369e+10, 
    1.181057e+10, 1.189166e+10, 1.196675e+10, 1.203567e+10, 1.209821e+10, 
    1.215424e+10, 1.220359e+10, 1.224615e+10, 1.228178e+10, 1.231041e+10, 
    1.233195e+10, 1.234634e+10, 1.235355e+10, 1.235355e+10, 1.234634e+10, 
    1.233195e+10, 1.231041e+10, 1.228178e+10, 1.224615e+10, 1.220359e+10, 
    1.215424e+10, 1.209821e+10, 1.203567e+10, 1.196675e+10, 1.189166e+10, 
    1.181057e+10, 1.172369e+10, 1.163122e+10, 1.153341e+10, 1.143046e+10, 
    1.132264e+10, 1.121017e+10, 1.109331e+10, 1.097232e+10, 1.084745e+10, 
    1.071896e+10, 1.058711e+10, 1.045215e+10, 1.031435e+10, 1.017395e+10, 
    1.00312e+10, 9.886363e+09, 9.739662e+09, 9.591338e+09, 9.441618e+09, 
    9.290724e+09, 9.138871e+09, 8.986266e+09, 8.833104e+09, 8.679578e+09, 
    8.525868e+09, 8.372148e+09, 8.218582e+09, 8.065324e+09, 7.912521e+09, 
    7.760311e+09, 7.608822e+09, 7.458176e+09, 7.308484e+09, 7.159848e+09, 
    7.012366e+09,
  6.992947e+09, 7.138521e+09, 7.285175e+09, 7.432813e+09, 7.581331e+09, 
    7.73062e+09, 7.880559e+09, 8.031022e+09, 8.181873e+09, 8.332967e+09, 
    8.484152e+09, 8.635267e+09, 8.786142e+09, 8.936601e+09, 9.086456e+09, 
    9.235513e+09, 9.383574e+09, 9.530426e+09, 9.675857e+09, 9.819643e+09, 
    9.961556e+09, 1.010136e+10, 1.023883e+10, 1.037371e+10, 1.050575e+10, 
    1.063472e+10, 1.076036e+10, 1.088243e+10, 1.100067e+10, 1.111483e+10, 
    1.122468e+10, 1.132997e+10, 1.143046e+10, 1.152593e+10, 1.161615e+10, 
    1.170091e+10, 1.178001e+10, 1.185324e+10, 1.192043e+10, 1.198141e+10, 
    1.203602e+10, 1.208412e+10, 1.212559e+10, 1.216031e+10, 1.218821e+10, 
    1.220919e+10, 1.222321e+10, 1.223023e+10, 1.223023e+10, 1.222321e+10, 
    1.220919e+10, 1.218821e+10, 1.216031e+10, 1.212559e+10, 1.208412e+10, 
    1.203602e+10, 1.198141e+10, 1.192043e+10, 1.185324e+10, 1.178001e+10, 
    1.170091e+10, 1.161615e+10, 1.152593e+10, 1.143046e+10, 1.132997e+10, 
    1.122468e+10, 1.111483e+10, 1.100067e+10, 1.088243e+10, 1.076036e+10, 
    1.063472e+10, 1.050575e+10, 1.037371e+10, 1.023883e+10, 1.010136e+10, 
    9.961556e+09, 9.819643e+09, 9.675857e+09, 9.530426e+09, 9.383574e+09, 
    9.235513e+09, 9.086456e+09, 8.936601e+09, 8.786142e+09, 8.635267e+09, 
    8.484152e+09, 8.332967e+09, 8.181873e+09, 8.031022e+09, 7.880559e+09, 
    7.73062e+09, 7.581331e+09, 7.432813e+09, 7.285175e+09, 7.138521e+09, 
    6.992947e+09,
  6.972339e+09, 7.115902e+09, 7.260469e+09, 7.405943e+09, 7.552224e+09, 
    7.699199e+09, 7.846753e+09, 7.994759e+09, 8.143084e+09, 8.291585e+09, 
    8.440113e+09, 8.58851e+09, 8.736609e+09, 8.884238e+09, 9.031216e+09, 
    9.177352e+09, 9.322452e+09, 9.466312e+09, 9.608722e+09, 9.749469e+09, 
    9.88833e+09, 1.002508e+10, 1.015949e+10, 1.029132e+10, 1.042034e+10, 
    1.054631e+10, 1.066899e+10, 1.078814e+10, 1.090352e+10, 1.10149e+10, 
    1.112203e+10, 1.122468e+10, 1.132264e+10, 1.141567e+10, 1.150357e+10, 
    1.158613e+10, 1.166315e+10, 1.173446e+10, 1.179987e+10, 1.185922e+10, 
    1.191237e+10, 1.195917e+10, 1.199952e+10, 1.203331e+10, 1.206044e+10, 
    1.208085e+10, 1.209449e+10, 1.210132e+10, 1.210132e+10, 1.209449e+10, 
    1.208085e+10, 1.206044e+10, 1.203331e+10, 1.199952e+10, 1.195917e+10, 
    1.191237e+10, 1.185922e+10, 1.179987e+10, 1.173446e+10, 1.166315e+10, 
    1.158613e+10, 1.150357e+10, 1.141567e+10, 1.132264e+10, 1.122468e+10, 
    1.112203e+10, 1.10149e+10, 1.090352e+10, 1.078814e+10, 1.066899e+10, 
    1.054631e+10, 1.042034e+10, 1.029132e+10, 1.015949e+10, 1.002508e+10, 
    9.88833e+09, 9.749469e+09, 9.608722e+09, 9.466312e+09, 9.322452e+09, 
    9.177352e+09, 9.031216e+09, 8.884238e+09, 8.736609e+09, 8.58851e+09, 
    8.440113e+09, 8.291585e+09, 8.143084e+09, 7.994759e+09, 7.846753e+09, 
    7.699199e+09, 7.552224e+09, 7.405943e+09, 7.260469e+09, 7.115902e+09, 
    6.972339e+09,
  6.950547e+09, 7.092e+09, 7.234377e+09, 7.377583e+09, 7.521518e+09, 
    7.666072e+09, 7.811129e+09, 7.956566e+09, 8.10225e+09, 8.248043e+09, 
    8.393798e+09, 8.539359e+09, 8.684566e+09, 8.829247e+09, 8.973229e+09, 
    9.116325e+09, 9.258346e+09, 9.399095e+09, 9.53837e+09, 9.67596e+09, 
    9.811654e+09, 9.945231e+09, 1.007647e+10, 1.020515e+10, 1.033104e+10, 
    1.045391e+10, 1.057352e+10, 1.068966e+10, 1.080209e+10, 1.091057e+10, 
    1.10149e+10, 1.111483e+10, 1.121017e+10, 1.130069e+10, 1.13862e+10, 
    1.146649e+10, 1.154138e+10, 1.16107e+10, 1.167428e+10, 1.173195e+10, 
    1.17836e+10, 1.182907e+10, 1.186826e+10, 1.190108e+10, 1.192743e+10, 
    1.194726e+10, 1.19605e+10, 1.196713e+10, 1.196713e+10, 1.19605e+10, 
    1.194726e+10, 1.192743e+10, 1.190108e+10, 1.186826e+10, 1.182907e+10, 
    1.17836e+10, 1.173195e+10, 1.167428e+10, 1.16107e+10, 1.154138e+10, 
    1.146649e+10, 1.13862e+10, 1.130069e+10, 1.121017e+10, 1.111483e+10, 
    1.10149e+10, 1.091057e+10, 1.080209e+10, 1.068966e+10, 1.057352e+10, 
    1.045391e+10, 1.033104e+10, 1.020515e+10, 1.007647e+10, 9.945231e+09, 
    9.811654e+09, 9.67596e+09, 9.53837e+09, 9.399095e+09, 9.258346e+09, 
    9.116325e+09, 8.973229e+09, 8.829247e+09, 8.684566e+09, 8.539359e+09, 
    8.393798e+09, 8.248043e+09, 8.10225e+09, 7.956566e+09, 7.811129e+09, 
    7.666072e+09, 7.521518e+09, 7.377583e+09, 7.234377e+09, 7.092e+09, 
    6.950547e+09,
  6.927576e+09, 7.066821e+09, 7.206909e+09, 7.347746e+09, 7.489233e+09, 
    7.631261e+09, 7.773715e+09, 7.916475e+09, 8.059411e+09, 8.202386e+09, 
    8.345257e+09, 8.487873e+09, 8.630074e+09, 8.771699e+09, 8.912572e+09, 
    9.052518e+09, 9.191351e+09, 9.32888e+09, 9.464909e+09, 9.599237e+09, 
    9.731658e+09, 9.861961e+09, 9.989933e+09, 1.011536e+10, 1.023802e+10, 
    1.035769e+10, 1.047415e+10, 1.058718e+10, 1.069657e+10, 1.080209e+10, 
    1.090352e+10, 1.100067e+10, 1.109331e+10, 1.118125e+10, 1.12643e+10, 
    1.134227e+10, 1.141498e+10, 1.148226e+10, 1.154395e+10, 1.159992e+10, 
    1.165001e+10, 1.169412e+10, 1.173213e+10, 1.176396e+10, 1.178951e+10, 
    1.180873e+10, 1.182158e+10, 1.1828e+10, 1.1828e+10, 1.182158e+10, 
    1.180873e+10, 1.178951e+10, 1.176396e+10, 1.173213e+10, 1.169412e+10, 
    1.165001e+10, 1.159992e+10, 1.154395e+10, 1.148226e+10, 1.141498e+10, 
    1.134227e+10, 1.12643e+10, 1.118125e+10, 1.109331e+10, 1.100067e+10, 
    1.090352e+10, 1.080209e+10, 1.069657e+10, 1.058718e+10, 1.047415e+10, 
    1.035769e+10, 1.023802e+10, 1.011536e+10, 9.989933e+09, 9.861961e+09, 
    9.731658e+09, 9.599237e+09, 9.464909e+09, 9.32888e+09, 9.191351e+09, 
    9.052518e+09, 8.912572e+09, 8.771699e+09, 8.630074e+09, 8.487873e+09, 
    8.345257e+09, 8.202386e+09, 8.059411e+09, 7.916475e+09, 7.773715e+09, 
    7.631261e+09, 7.489233e+09, 7.347746e+09, 7.206909e+09, 7.066821e+09, 
    6.927576e+09,
  6.903431e+09, 7.040374e+09, 7.178077e+09, 7.316448e+09, 7.455388e+09, 
    7.594789e+09, 7.734541e+09, 7.874522e+09, 8.014606e+09, 8.15466e+09, 
    8.294543e+09, 8.434108e+09, 8.573202e+09, 8.711665e+09, 8.849328e+09, 
    8.986021e+09, 9.121564e+09, 9.255772e+09, 9.388457e+09, 9.519426e+09, 
    9.648477e+09, 9.775411e+09, 9.900023e+09, 1.00221e+10, 1.014144e+10, 
    1.025783e+10, 1.037106e+10, 1.048091e+10, 1.058718e+10, 1.068966e+10, 
    1.078814e+10, 1.088243e+10, 1.097232e+10, 1.105763e+10, 1.113816e+10, 
    1.121375e+10, 1.128423e+10, 1.134943e+10, 1.14092e+10, 1.146341e+10, 
    1.151193e+10, 1.155465e+10, 1.159146e+10, 1.162227e+10, 1.164701e+10, 
    1.166561e+10, 1.167804e+10, 1.168427e+10, 1.168427e+10, 1.167804e+10, 
    1.166561e+10, 1.164701e+10, 1.162227e+10, 1.159146e+10, 1.155465e+10, 
    1.151193e+10, 1.146341e+10, 1.14092e+10, 1.134943e+10, 1.128423e+10, 
    1.121375e+10, 1.113816e+10, 1.105763e+10, 1.097232e+10, 1.088243e+10, 
    1.078814e+10, 1.068966e+10, 1.058718e+10, 1.048091e+10, 1.037106e+10, 
    1.025783e+10, 1.014144e+10, 1.00221e+10, 9.900023e+09, 9.775411e+09, 
    9.648477e+09, 9.519426e+09, 9.388457e+09, 9.255772e+09, 9.121564e+09, 
    8.986021e+09, 8.849328e+09, 8.711665e+09, 8.573202e+09, 8.434108e+09, 
    8.294543e+09, 8.15466e+09, 8.014606e+09, 7.874522e+09, 7.734541e+09, 
    7.594789e+09, 7.455388e+09, 7.316448e+09, 7.178077e+09, 7.040374e+09, 
    6.903431e+09,
  6.878117e+09, 7.012667e+09, 7.147894e+09, 7.283705e+09, 7.420003e+09, 
    7.556683e+09, 7.693634e+09, 7.830739e+09, 7.967875e+09, 8.10491e+09, 
    8.241709e+09, 8.378128e+09, 8.514017e+09, 8.649221e+09, 8.78358e+09, 
    8.916924e+09, 9.049084e+09, 9.17988e+09, 9.309132e+09, 9.436652e+09, 
    9.562249e+09, 9.68573e+09, 9.806899e+09, 9.925557e+09, 1.00415e+10, 
    1.015454e+10, 1.026446e+10, 1.037106e+10, 1.047415e+10, 1.057352e+10, 
    1.066899e+10, 1.076036e+10, 1.084745e+10, 1.093007e+10, 1.100805e+10, 
    1.108122e+10, 1.114942e+10, 1.12125e+10, 1.127033e+10, 1.132276e+10, 
    1.136968e+10, 1.141097e+10, 1.144656e+10, 1.147634e+10, 1.150025e+10, 
    1.151823e+10, 1.153025e+10, 1.153626e+10, 1.153626e+10, 1.153025e+10, 
    1.151823e+10, 1.150025e+10, 1.147634e+10, 1.144656e+10, 1.141097e+10, 
    1.136968e+10, 1.132276e+10, 1.127033e+10, 1.12125e+10, 1.114942e+10, 
    1.108122e+10, 1.100805e+10, 1.093007e+10, 1.084745e+10, 1.076036e+10, 
    1.066899e+10, 1.057352e+10, 1.047415e+10, 1.037106e+10, 1.026446e+10, 
    1.015454e+10, 1.00415e+10, 9.925557e+09, 9.806899e+09, 9.68573e+09, 
    9.562249e+09, 9.436652e+09, 9.309132e+09, 9.17988e+09, 9.049084e+09, 
    8.916924e+09, 8.78358e+09, 8.649221e+09, 8.514017e+09, 8.378128e+09, 
    8.241709e+09, 8.10491e+09, 7.967875e+09, 7.830739e+09, 7.693634e+09, 
    7.556683e+09, 7.420003e+09, 7.283705e+09, 7.147894e+09, 7.012667e+09, 
    6.878117e+09,
  6.851641e+09, 6.98371e+09, 7.116371e+09, 7.249533e+09, 7.383099e+09, 
    7.516966e+09, 7.651027e+09, 7.785166e+09, 7.919261e+09, 8.053188e+09, 
    8.186811e+09, 8.319992e+09, 8.452588e+09, 8.584445e+09, 8.715411e+09, 
    8.845323e+09, 8.974015e+09, 9.101317e+09, 9.227054e+09, 9.351046e+09, 
    9.473112e+09, 9.593066e+09, 9.710721e+09, 9.825887e+09, 9.938373e+09, 
    1.004799e+10, 1.015454e+10, 1.025783e+10, 1.035769e+10, 1.045391e+10, 
    1.054631e+10, 1.063472e+10, 1.071896e+10, 1.079885e+10, 1.087423e+10, 
    1.094495e+10, 1.101085e+10, 1.107179e+10, 1.112763e+10, 1.117826e+10, 
    1.122356e+10, 1.126342e+10, 1.129776e+10, 1.13265e+10, 1.134958e+10, 
    1.136693e+10, 1.137852e+10, 1.138432e+10, 1.138432e+10, 1.137852e+10, 
    1.136693e+10, 1.134958e+10, 1.13265e+10, 1.129776e+10, 1.126342e+10, 
    1.122356e+10, 1.117826e+10, 1.112763e+10, 1.107179e+10, 1.101085e+10, 
    1.094495e+10, 1.087423e+10, 1.079885e+10, 1.071896e+10, 1.063472e+10, 
    1.054631e+10, 1.045391e+10, 1.035769e+10, 1.025783e+10, 1.015454e+10, 
    1.004799e+10, 9.938373e+09, 9.825887e+09, 9.710721e+09, 9.593066e+09, 
    9.473112e+09, 9.351046e+09, 9.227054e+09, 9.101317e+09, 8.974015e+09, 
    8.845323e+09, 8.715411e+09, 8.584445e+09, 8.452588e+09, 8.319992e+09, 
    8.186811e+09, 8.053188e+09, 7.919261e+09, 7.785166e+09, 7.651027e+09, 
    7.516966e+09, 7.383099e+09, 7.249533e+09, 7.116371e+09, 6.98371e+09, 
    6.851641e+09,
  6.824007e+09, 6.953512e+09, 7.083523e+09, 7.21395e+09, 7.344698e+09, 
    7.475667e+09, 7.606751e+09, 7.737838e+09, 7.868808e+09, 7.99954e+09, 
    8.129904e+09, 8.259766e+09, 8.388985e+09, 8.517416e+09, 8.64491e+09, 
    8.771312e+09, 8.896461e+09, 9.020195e+09, 9.142345e+09, 9.262742e+09, 
    9.381209e+09, 9.497571e+09, 9.61165e+09, 9.723264e+09, 9.832232e+09, 
    9.938373e+09, 1.00415e+10, 1.014144e+10, 1.023802e+10, 1.033104e+10, 
    1.042034e+10, 1.050575e+10, 1.058711e+10, 1.066424e+10, 1.0737e+10, 
    1.080523e+10, 1.08688e+10, 1.092757e+10, 1.098142e+10, 1.103023e+10, 
    1.107389e+10, 1.111231e+10, 1.11454e+10, 1.117309e+10, 1.119532e+10, 
    1.121203e+10, 1.12232e+10, 1.122879e+10, 1.122879e+10, 1.12232e+10, 
    1.121203e+10, 1.119532e+10, 1.117309e+10, 1.11454e+10, 1.111231e+10, 
    1.107389e+10, 1.103023e+10, 1.098142e+10, 1.092757e+10, 1.08688e+10, 
    1.080523e+10, 1.0737e+10, 1.066424e+10, 1.058711e+10, 1.050575e+10, 
    1.042034e+10, 1.033104e+10, 1.023802e+10, 1.014144e+10, 1.00415e+10, 
    9.938373e+09, 9.832232e+09, 9.723264e+09, 9.61165e+09, 9.497571e+09, 
    9.381209e+09, 9.262742e+09, 9.142345e+09, 9.020195e+09, 8.896461e+09, 
    8.771312e+09, 8.64491e+09, 8.517416e+09, 8.388985e+09, 8.259766e+09, 
    8.129904e+09, 7.99954e+09, 7.868808e+09, 7.737838e+09, 7.606751e+09, 
    7.475667e+09, 7.344698e+09, 7.21395e+09, 7.083523e+09, 6.953512e+09, 
    6.824007e+09,
  6.795221e+09, 6.922081e+09, 7.049361e+09, 7.176973e+09, 7.304823e+09, 
    7.432814e+09, 7.56084e+09, 7.688794e+09, 7.816561e+09, 7.94402e+09, 
    8.071048e+09, 8.197513e+09, 8.323282e+09, 8.448214e+09, 8.572165e+09, 
    8.694987e+09, 8.816526e+09, 8.936627e+09, 9.055129e+09, 9.171869e+09, 
    9.286681e+09, 9.399396e+09, 9.509846e+09, 9.61786e+09, 9.723264e+09, 
    9.825887e+09, 9.925557e+09, 1.00221e+10, 1.011536e+10, 1.020515e+10, 
    1.029132e+10, 1.037371e+10, 1.045215e+10, 1.05265e+10, 1.059662e+10, 
    1.066235e+10, 1.072358e+10, 1.078017e+10, 1.0832e+10, 1.087898e+10, 
    1.092099e+10, 1.095795e+10, 1.098979e+10, 1.101642e+10, 1.10378e+10, 
    1.105388e+10, 1.106461e+10, 1.106999e+10, 1.106999e+10, 1.106461e+10, 
    1.105388e+10, 1.10378e+10, 1.101642e+10, 1.098979e+10, 1.095795e+10, 
    1.092099e+10, 1.087898e+10, 1.0832e+10, 1.078017e+10, 1.072358e+10, 
    1.066235e+10, 1.059662e+10, 1.05265e+10, 1.045215e+10, 1.037371e+10, 
    1.029132e+10, 1.020515e+10, 1.011536e+10, 1.00221e+10, 9.925557e+09, 
    9.825887e+09, 9.723264e+09, 9.61786e+09, 9.509846e+09, 9.399396e+09, 
    9.286681e+09, 9.171869e+09, 9.055129e+09, 8.936627e+09, 8.816526e+09, 
    8.694987e+09, 8.572165e+09, 8.448214e+09, 8.323282e+09, 8.197513e+09, 
    8.071048e+09, 7.94402e+09, 7.816561e+09, 7.688794e+09, 7.56084e+09, 
    7.432814e+09, 7.304823e+09, 7.176973e+09, 7.049361e+09, 6.922081e+09, 
    6.795221e+09,
  6.76529e+09, 6.889429e+09, 7.013901e+09, 7.13862e+09, 7.263496e+09, 
    7.388432e+09, 7.513327e+09, 7.638074e+09, 7.762563e+09, 7.886679e+09, 
    8.010299e+09, 8.133301e+09, 8.255552e+09, 8.37692e+09, 8.497266e+09, 
    8.616447e+09, 8.734319e+09, 8.85073e+09, 8.96553e+09, 9.078562e+09, 
    9.18967e+09, 9.298694e+09, 9.405474e+09, 9.509846e+09, 9.61165e+09, 
    9.710721e+09, 9.806899e+09, 9.900023e+09, 9.989933e+09, 1.007647e+10, 
    1.015949e+10, 1.023883e+10, 1.031435e+10, 1.03859e+10, 1.045336e+10, 
    1.051658e+10, 1.057545e+10, 1.062985e+10, 1.067967e+10, 1.07248e+10, 
    1.076517e+10, 1.080067e+10, 1.083124e+10, 1.085682e+10, 1.087735e+10, 
    1.089278e+10, 1.090309e+10, 1.090825e+10, 1.090825e+10, 1.090309e+10, 
    1.089278e+10, 1.087735e+10, 1.085682e+10, 1.083124e+10, 1.080067e+10, 
    1.076517e+10, 1.07248e+10, 1.067967e+10, 1.062985e+10, 1.057545e+10, 
    1.051658e+10, 1.045336e+10, 1.03859e+10, 1.031435e+10, 1.023883e+10, 
    1.015949e+10, 1.007647e+10, 9.989933e+09, 9.900023e+09, 9.806899e+09, 
    9.710721e+09, 9.61165e+09, 9.509846e+09, 9.405474e+09, 9.298694e+09, 
    9.18967e+09, 9.078562e+09, 8.96553e+09, 8.85073e+09, 8.734319e+09, 
    8.616447e+09, 8.497266e+09, 8.37692e+09, 8.255552e+09, 8.133301e+09, 
    8.010299e+09, 7.886679e+09, 7.762563e+09, 7.638074e+09, 7.513327e+09, 
    7.388432e+09, 7.263496e+09, 7.13862e+09, 7.013901e+09, 6.889429e+09, 
    6.76529e+09,
  6.734221e+09, 6.855565e+09, 6.977157e+09, 7.098912e+09, 7.220742e+09, 
    7.342552e+09, 7.464245e+09, 7.585717e+09, 7.706863e+09, 7.827569e+09, 
    7.94772e+09, 8.067195e+09, 8.18587e+09, 8.303616e+09, 8.420301e+09, 
    8.53579e+09, 8.649944e+09, 8.762619e+09, 8.873673e+09, 8.982957e+09, 
    9.090322e+09, 9.195619e+09, 9.298694e+09, 9.399396e+09, 9.497571e+09, 
    9.593066e+09, 9.68573e+09, 9.775411e+09, 9.861961e+09, 9.945231e+09, 
    1.002508e+10, 1.010136e+10, 1.017395e+10, 1.02427e+10, 1.030749e+10, 
    1.03682e+10, 1.042471e+10, 1.047692e+10, 1.052472e+10, 1.056802e+10, 
    1.060673e+10, 1.064077e+10, 1.067009e+10, 1.06946e+10, 1.071428e+10, 
    1.072907e+10, 1.073895e+10, 1.07439e+10, 1.07439e+10, 1.073895e+10, 
    1.072907e+10, 1.071428e+10, 1.06946e+10, 1.067009e+10, 1.064077e+10, 
    1.060673e+10, 1.056802e+10, 1.052472e+10, 1.047692e+10, 1.042471e+10, 
    1.03682e+10, 1.030749e+10, 1.02427e+10, 1.017395e+10, 1.010136e+10, 
    1.002508e+10, 9.945231e+09, 9.861961e+09, 9.775411e+09, 9.68573e+09, 
    9.593066e+09, 9.497571e+09, 9.399396e+09, 9.298694e+09, 9.195619e+09, 
    9.090322e+09, 8.982957e+09, 8.873673e+09, 8.762619e+09, 8.649944e+09, 
    8.53579e+09, 8.420301e+09, 8.303616e+09, 8.18587e+09, 8.067195e+09, 
    7.94772e+09, 7.827569e+09, 7.706863e+09, 7.585717e+09, 7.464245e+09, 
    7.342552e+09, 7.220742e+09, 7.098912e+09, 6.977157e+09, 6.855565e+09, 
    6.734221e+09,
  6.702019e+09, 6.8205e+09, 6.939143e+09, 7.057866e+09, 7.176583e+09, 
    7.295202e+09, 7.41363e+09, 7.531766e+09, 7.649507e+09, 7.766745e+09, 
    7.883369e+09, 7.999264e+09, 8.11431e+09, 8.228386e+09, 8.341364e+09, 
    8.453116e+09, 8.563511e+09, 8.672412e+09, 8.779684e+09, 8.885187e+09, 
    8.988781e+09, 9.090322e+09, 9.18967e+09, 9.286681e+09, 9.381209e+09, 
    9.473112e+09, 9.562249e+09, 9.648477e+09, 9.731658e+09, 9.811654e+09, 
    9.88833e+09, 9.961556e+09, 1.00312e+10, 1.009715e+10, 1.015928e+10, 
    1.021748e+10, 1.027164e+10, 1.032166e+10, 1.036744e+10, 1.040891e+10, 
    1.044597e+10, 1.047856e+10, 1.050662e+10, 1.053008e+10, 1.054891e+10, 
    1.056306e+10, 1.057252e+10, 1.057725e+10, 1.057725e+10, 1.057252e+10, 
    1.056306e+10, 1.054891e+10, 1.053008e+10, 1.050662e+10, 1.047856e+10, 
    1.044597e+10, 1.040891e+10, 1.036744e+10, 1.032166e+10, 1.027164e+10, 
    1.021748e+10, 1.015928e+10, 1.009715e+10, 1.00312e+10, 9.961556e+09, 
    9.88833e+09, 9.811654e+09, 9.731658e+09, 9.648477e+09, 9.562249e+09, 
    9.473112e+09, 9.381209e+09, 9.286681e+09, 9.18967e+09, 9.090322e+09, 
    8.988781e+09, 8.885187e+09, 8.779684e+09, 8.672412e+09, 8.563511e+09, 
    8.453116e+09, 8.341364e+09, 8.228386e+09, 8.11431e+09, 7.999264e+09, 
    7.883369e+09, 7.766745e+09, 7.649507e+09, 7.531766e+09, 7.41363e+09, 
    7.295202e+09, 7.176583e+09, 7.057866e+09, 6.939143e+09, 6.8205e+09, 
    6.702019e+09,
  6.668692e+09, 6.784244e+09, 6.899874e+09, 7.015503e+09, 7.131045e+09, 
    7.246414e+09, 7.361518e+09, 7.47626e+09, 7.590542e+09, 7.704261e+09, 
    7.817309e+09, 7.929576e+09, 8.04095e+09, 8.151313e+09, 8.260545e+09, 
    8.368525e+09, 8.475127e+09, 8.580225e+09, 8.683688e+09, 8.785385e+09, 
    8.885187e+09, 8.982957e+09, 9.078562e+09, 9.171869e+09, 9.262742e+09, 
    9.351046e+09, 9.436652e+09, 9.519426e+09, 9.599237e+09, 9.67596e+09, 
    9.749469e+09, 9.819643e+09, 9.886363e+09, 9.949515e+09, 1.000899e+10, 
    1.006469e+10, 1.01165e+10, 1.016434e+10, 1.020812e+10, 1.024776e+10, 
    1.028319e+10, 1.031433e+10, 1.034114e+10, 1.036355e+10, 1.038154e+10, 
    1.039506e+10, 1.040409e+10, 1.040861e+10, 1.040861e+10, 1.040409e+10, 
    1.039506e+10, 1.038154e+10, 1.036355e+10, 1.034114e+10, 1.031433e+10, 
    1.028319e+10, 1.024776e+10, 1.020812e+10, 1.016434e+10, 1.01165e+10, 
    1.006469e+10, 1.000899e+10, 9.949515e+09, 9.886363e+09, 9.819643e+09, 
    9.749469e+09, 9.67596e+09, 9.599237e+09, 9.519426e+09, 9.436652e+09, 
    9.351046e+09, 9.262742e+09, 9.171869e+09, 9.078562e+09, 8.982957e+09, 
    8.885187e+09, 8.785385e+09, 8.683688e+09, 8.580225e+09, 8.475127e+09, 
    8.368525e+09, 8.260545e+09, 8.151313e+09, 8.04095e+09, 7.929576e+09, 
    7.817309e+09, 7.704261e+09, 7.590542e+09, 7.47626e+09, 7.361518e+09, 
    7.246414e+09, 7.131045e+09, 7.015503e+09, 6.899874e+09, 6.784244e+09, 
    6.668692e+09,
  6.634248e+09, 6.74681e+09, 6.859367e+09, 6.971842e+09, 7.084154e+09, 
    7.196217e+09, 7.307944e+09, 7.419243e+09, 7.530018e+09, 7.640172e+09, 
    7.749601e+09, 7.858201e+09, 7.965864e+09, 8.072481e+09, 8.177936e+09, 
    8.282116e+09, 8.384902e+09, 8.486173e+09, 8.585809e+09, 8.683688e+09, 
    8.779684e+09, 8.873673e+09, 8.96553e+09, 9.055129e+09, 9.142345e+09, 
    9.227054e+09, 9.309132e+09, 9.388457e+09, 9.464909e+09, 9.53837e+09, 
    9.608722e+09, 9.675857e+09, 9.739662e+09, 9.800034e+09, 9.856871e+09, 
    9.910078e+09, 9.959563e+09, 1.000524e+10, 1.004703e+10, 1.008486e+10, 
    1.011866e+10, 1.014837e+10, 1.017394e+10, 1.019532e+10, 1.021247e+10, 
    1.022536e+10, 1.023397e+10, 1.023827e+10, 1.023827e+10, 1.023397e+10, 
    1.022536e+10, 1.021247e+10, 1.019532e+10, 1.017394e+10, 1.014837e+10, 
    1.011866e+10, 1.008486e+10, 1.004703e+10, 1.000524e+10, 9.959563e+09, 
    9.910078e+09, 9.856871e+09, 9.800034e+09, 9.739662e+09, 9.675857e+09, 
    9.608722e+09, 9.53837e+09, 9.464909e+09, 9.388457e+09, 9.309132e+09, 
    9.227054e+09, 9.142345e+09, 9.055129e+09, 8.96553e+09, 8.873673e+09, 
    8.779684e+09, 8.683688e+09, 8.585809e+09, 8.486173e+09, 8.384902e+09, 
    8.282116e+09, 8.177936e+09, 8.072481e+09, 7.965864e+09, 7.858201e+09, 
    7.749601e+09, 7.640172e+09, 7.530018e+09, 7.419243e+09, 7.307944e+09, 
    7.196217e+09, 7.084154e+09, 6.971842e+09, 6.859367e+09, 6.74681e+09, 
    6.634248e+09,
  6.598693e+09, 6.708208e+09, 6.817636e+09, 6.926904e+09, 7.035934e+09, 
    7.144643e+09, 7.252946e+09, 7.360757e+09, 7.467984e+09, 7.574533e+09, 
    7.680307e+09, 7.785207e+09, 7.889131e+09, 7.991974e+09, 8.093629e+09, 
    8.193989e+09, 8.292941e+09, 8.390374e+09, 8.486173e+09, 8.580225e+09, 
    8.672412e+09, 8.762619e+09, 8.85073e+09, 8.936627e+09, 9.020195e+09, 
    9.101317e+09, 9.17988e+09, 9.255772e+09, 9.32888e+09, 9.399095e+09, 
    9.466312e+09, 9.530426e+09, 9.591338e+09, 9.64895e+09, 9.703171e+09, 
    9.753911e+09, 9.801088e+09, 9.844622e+09, 9.884442e+09, 9.920478e+09, 
    9.95267e+09, 9.980962e+09, 1.00053e+10, 1.002566e+10, 1.004198e+10, 
    1.005425e+10, 1.006244e+10, 1.006654e+10, 1.006654e+10, 1.006244e+10, 
    1.005425e+10, 1.004198e+10, 1.002566e+10, 1.00053e+10, 9.980962e+09, 
    9.95267e+09, 9.920478e+09, 9.884442e+09, 9.844622e+09, 9.801088e+09, 
    9.753911e+09, 9.703171e+09, 9.64895e+09, 9.591338e+09, 9.530426e+09, 
    9.466312e+09, 9.399095e+09, 9.32888e+09, 9.255772e+09, 9.17988e+09, 
    9.101317e+09, 9.020195e+09, 8.936627e+09, 8.85073e+09, 8.762619e+09, 
    8.672412e+09, 8.580225e+09, 8.486173e+09, 8.390374e+09, 8.292941e+09, 
    8.193989e+09, 8.093629e+09, 7.991974e+09, 7.889131e+09, 7.785207e+09, 
    7.680307e+09, 7.574533e+09, 7.467984e+09, 7.360757e+09, 7.252946e+09, 
    7.144643e+09, 7.035934e+09, 6.926904e+09, 6.817636e+09, 6.708208e+09, 
    6.598693e+09,
  6.562035e+09, 6.668449e+09, 6.774699e+09, 6.880711e+09, 6.986412e+09, 
    7.091722e+09, 7.196561e+09, 7.300845e+09, 7.404488e+09, 7.5074e+09, 
    7.60949e+09, 7.710664e+09, 7.810825e+09, 7.909876e+09, 8.007716e+09, 
    8.104243e+09, 8.199353e+09, 8.292941e+09, 8.384902e+09, 8.475127e+09, 
    8.563511e+09, 8.649944e+09, 8.734319e+09, 8.816526e+09, 8.896461e+09, 
    8.974015e+09, 9.049084e+09, 9.121564e+09, 9.191351e+09, 9.258346e+09, 
    9.322452e+09, 9.383574e+09, 9.441618e+09, 9.496498e+09, 9.548129e+09, 
    9.596429e+09, 9.641325e+09, 9.68274e+09, 9.720613e+09, 9.754878e+09, 
    9.785482e+09, 9.812372e+09, 9.835507e+09, 9.854844e+09, 9.870353e+09, 
    9.882009e+09, 9.88979e+09, 9.893683e+09, 9.893683e+09, 9.88979e+09, 
    9.882009e+09, 9.870353e+09, 9.854844e+09, 9.835507e+09, 9.812372e+09, 
    9.785482e+09, 9.754878e+09, 9.720613e+09, 9.68274e+09, 9.641325e+09, 
    9.596429e+09, 9.548129e+09, 9.496498e+09, 9.441618e+09, 9.383574e+09, 
    9.322452e+09, 9.258346e+09, 9.191351e+09, 9.121564e+09, 9.049084e+09, 
    8.974015e+09, 8.896461e+09, 8.816526e+09, 8.734319e+09, 8.649944e+09, 
    8.563511e+09, 8.475127e+09, 8.384902e+09, 8.292941e+09, 8.199353e+09, 
    8.104243e+09, 8.007716e+09, 7.909876e+09, 7.810825e+09, 7.710664e+09, 
    7.60949e+09, 7.5074e+09, 7.404488e+09, 7.300845e+09, 7.196561e+09, 
    7.091722e+09, 6.986412e+09, 6.880711e+09, 6.774699e+09, 6.668449e+09, 
    6.562035e+09,
  6.524282e+09, 6.627547e+09, 6.730571e+09, 6.833284e+09, 6.935614e+09, 
    7.037487e+09, 7.138825e+09, 7.23955e+09, 7.339579e+09, 7.438829e+09, 
    7.537212e+09, 7.634641e+09, 7.731025e+09, 7.826271e+09, 7.920287e+09, 
    8.012976e+09, 8.104243e+09, 8.193989e+09, 8.282116e+09, 8.368525e+09, 
    8.453116e+09, 8.53579e+09, 8.616447e+09, 8.694987e+09, 8.771312e+09, 
    8.845323e+09, 8.916924e+09, 8.986021e+09, 9.052518e+09, 9.116325e+09, 
    9.177352e+09, 9.235513e+09, 9.290724e+09, 9.342905e+09, 9.391978e+09, 
    9.437871e+09, 9.480515e+09, 9.519842e+09, 9.555794e+09, 9.588315e+09, 
    9.617354e+09, 9.642865e+09, 9.664807e+09, 9.683147e+09, 9.697854e+09, 
    9.708905e+09, 9.716282e+09, 9.719975e+09, 9.719975e+09, 9.716282e+09, 
    9.708905e+09, 9.697854e+09, 9.683147e+09, 9.664807e+09, 9.642865e+09, 
    9.617354e+09, 9.588315e+09, 9.555794e+09, 9.519842e+09, 9.480515e+09, 
    9.437871e+09, 9.391978e+09, 9.342905e+09, 9.290724e+09, 9.235513e+09, 
    9.177352e+09, 9.116325e+09, 9.052518e+09, 8.986021e+09, 8.916924e+09, 
    8.845323e+09, 8.771312e+09, 8.694987e+09, 8.616447e+09, 8.53579e+09, 
    8.453116e+09, 8.368525e+09, 8.282116e+09, 8.193989e+09, 8.104243e+09, 
    8.012976e+09, 7.920287e+09, 7.826271e+09, 7.731025e+09, 7.634641e+09, 
    7.537212e+09, 7.438829e+09, 7.339579e+09, 7.23955e+09, 7.138825e+09, 
    7.037487e+09, 6.935614e+09, 6.833284e+09, 6.730571e+09, 6.627547e+09, 
    6.524282e+09,
  6.485442e+09, 6.585513e+09, 6.685269e+09, 6.784643e+09, 6.883567e+09, 
    6.981969e+09, 7.079777e+09, 7.176916e+09, 7.273309e+09, 7.368877e+09, 
    7.463537e+09, 7.557208e+09, 7.649805e+09, 7.741242e+09, 7.831433e+09, 
    7.920287e+09, 8.007716e+09, 8.093629e+09, 8.177936e+09, 8.260545e+09, 
    8.341364e+09, 8.420301e+09, 8.497266e+09, 8.572165e+09, 8.64491e+09, 
    8.715411e+09, 8.78358e+09, 8.849328e+09, 8.912572e+09, 8.973229e+09, 
    9.031216e+09, 9.086456e+09, 9.138871e+09, 9.188391e+09, 9.234944e+09, 
    9.278465e+09, 9.318892e+09, 9.356163e+09, 9.390226e+09, 9.421031e+09, 
    9.448532e+09, 9.472687e+09, 9.49346e+09, 9.510819e+09, 9.524738e+09, 
    9.535196e+09, 9.542177e+09, 9.54567e+09, 9.54567e+09, 9.542177e+09, 
    9.535196e+09, 9.524738e+09, 9.510819e+09, 9.49346e+09, 9.472687e+09, 
    9.448532e+09, 9.421031e+09, 9.390226e+09, 9.356163e+09, 9.318892e+09, 
    9.278465e+09, 9.234944e+09, 9.188391e+09, 9.138871e+09, 9.086456e+09, 
    9.031216e+09, 8.973229e+09, 8.912572e+09, 8.849328e+09, 8.78358e+09, 
    8.715411e+09, 8.64491e+09, 8.572165e+09, 8.497266e+09, 8.420301e+09, 
    8.341364e+09, 8.260545e+09, 8.177936e+09, 8.093629e+09, 8.007716e+09, 
    7.920287e+09, 7.831433e+09, 7.741242e+09, 7.649805e+09, 7.557208e+09, 
    7.463537e+09, 7.368877e+09, 7.273309e+09, 7.176916e+09, 7.079777e+09, 
    6.981969e+09, 6.883567e+09, 6.784643e+09, 6.685269e+09, 6.585513e+09, 
    6.485442e+09,
  6.445522e+09, 6.54236e+09, 6.638811e+09, 6.734811e+09, 6.830297e+09, 
    6.925201e+09, 7.019455e+09, 7.112987e+09, 7.205726e+09, 7.297597e+09, 
    7.388526e+09, 7.478433e+09, 7.567242e+09, 7.654872e+09, 7.741242e+09, 
    7.826271e+09, 7.909876e+09, 7.991974e+09, 8.072481e+09, 8.151313e+09, 
    8.228386e+09, 8.303616e+09, 8.37692e+09, 8.448214e+09, 8.517416e+09, 
    8.584445e+09, 8.649221e+09, 8.711665e+09, 8.771699e+09, 8.829247e+09, 
    8.884238e+09, 8.936601e+09, 8.986266e+09, 9.033167e+09, 9.077242e+09, 
    9.118431e+09, 9.156679e+09, 9.191932e+09, 9.224142e+09, 9.253263e+09, 
    9.279254e+09, 9.302078e+09, 9.321703e+09, 9.338102e+09, 9.351248e+09, 
    9.361125e+09, 9.367718e+09, 9.371016e+09, 9.371016e+09, 9.367718e+09, 
    9.361125e+09, 9.351248e+09, 9.338102e+09, 9.321703e+09, 9.302078e+09, 
    9.279254e+09, 9.253263e+09, 9.224142e+09, 9.191932e+09, 9.156679e+09, 
    9.118431e+09, 9.077242e+09, 9.033167e+09, 8.986266e+09, 8.936601e+09, 
    8.884238e+09, 8.829247e+09, 8.771699e+09, 8.711665e+09, 8.649221e+09, 
    8.584445e+09, 8.517416e+09, 8.448214e+09, 8.37692e+09, 8.303616e+09, 
    8.228386e+09, 8.151313e+09, 8.072481e+09, 7.991974e+09, 7.909876e+09, 
    7.826271e+09, 7.741242e+09, 7.654872e+09, 7.567242e+09, 7.478433e+09, 
    7.388526e+09, 7.297597e+09, 7.205726e+09, 7.112987e+09, 7.019455e+09, 
    6.925201e+09, 6.830297e+09, 6.734811e+09, 6.638811e+09, 6.54236e+09, 
    6.445522e+09,
  6.404531e+09, 6.4981e+09, 6.591213e+09, 6.683811e+09, 6.775833e+09, 
    6.867216e+09, 6.957896e+09, 7.047806e+09, 7.136881e+09, 7.225049e+09, 
    7.312241e+09, 7.398386e+09, 7.483411e+09, 7.567242e+09, 7.649805e+09, 
    7.731025e+09, 7.810825e+09, 7.889131e+09, 7.965864e+09, 8.04095e+09, 
    8.11431e+09, 8.18587e+09, 8.255552e+09, 8.323282e+09, 8.388985e+09, 
    8.452588e+09, 8.514017e+09, 8.573202e+09, 8.630074e+09, 8.684566e+09, 
    8.736609e+09, 8.786142e+09, 8.833104e+09, 8.877434e+09, 8.919077e+09, 
    8.95798e+09, 8.994092e+09, 9.027367e+09, 9.05776e+09, 9.085231e+09, 
    9.109745e+09, 9.131267e+09, 9.14977e+09, 9.165227e+09, 9.177618e+09, 
    9.186927e+09, 9.193139e+09, 9.196247e+09, 9.196247e+09, 9.193139e+09, 
    9.186927e+09, 9.177618e+09, 9.165227e+09, 9.14977e+09, 9.131267e+09, 
    9.109745e+09, 9.085231e+09, 9.05776e+09, 9.027367e+09, 8.994092e+09, 
    8.95798e+09, 8.919077e+09, 8.877434e+09, 8.833104e+09, 8.786142e+09, 
    8.736609e+09, 8.684566e+09, 8.630074e+09, 8.573202e+09, 8.514017e+09, 
    8.452588e+09, 8.388985e+09, 8.323282e+09, 8.255552e+09, 8.18587e+09, 
    8.11431e+09, 8.04095e+09, 7.965864e+09, 7.889131e+09, 7.810825e+09, 
    7.731025e+09, 7.649805e+09, 7.567242e+09, 7.483411e+09, 7.398386e+09, 
    7.312241e+09, 7.225049e+09, 7.136881e+09, 7.047806e+09, 6.957896e+09, 
    6.867216e+09, 6.775833e+09, 6.683811e+09, 6.591213e+09, 6.4981e+09, 
    6.404531e+09,
  6.362479e+09, 6.452746e+09, 6.542493e+09, 6.631664e+09, 6.720201e+09, 
    6.808046e+09, 6.895139e+09, 6.981418e+09, 7.066822e+09, 7.151286e+09, 
    7.234745e+09, 7.317134e+09, 7.398386e+09, 7.478433e+09, 7.557208e+09, 
    7.634641e+09, 7.710664e+09, 7.785207e+09, 7.858201e+09, 7.929576e+09, 
    7.999264e+09, 8.067195e+09, 8.133301e+09, 8.197513e+09, 8.259766e+09, 
    8.319992e+09, 8.378128e+09, 8.434108e+09, 8.487873e+09, 8.539359e+09, 
    8.58851e+09, 8.635267e+09, 8.679578e+09, 8.721389e+09, 8.760649e+09, 
    8.797313e+09, 8.831335e+09, 8.862674e+09, 8.891291e+09, 8.917151e+09, 
    8.940219e+09, 8.96047e+09, 8.977876e+09, 8.992415e+09, 9.004068e+09, 
    9.012821e+09, 9.018663e+09, 9.021585e+09, 9.021585e+09, 9.018663e+09, 
    9.012821e+09, 9.004068e+09, 8.992415e+09, 8.977876e+09, 8.96047e+09, 
    8.940219e+09, 8.917151e+09, 8.891291e+09, 8.862674e+09, 8.831335e+09, 
    8.797313e+09, 8.760649e+09, 8.721389e+09, 8.679578e+09, 8.635267e+09, 
    8.58851e+09, 8.539359e+09, 8.487873e+09, 8.434108e+09, 8.378128e+09, 
    8.319992e+09, 8.259766e+09, 8.197513e+09, 8.133301e+09, 8.067195e+09, 
    7.999264e+09, 7.929576e+09, 7.858201e+09, 7.785207e+09, 7.710664e+09, 
    7.634641e+09, 7.557208e+09, 7.478433e+09, 7.398386e+09, 7.317134e+09, 
    7.234745e+09, 7.151286e+09, 7.066822e+09, 6.981418e+09, 6.895139e+09, 
    6.808046e+09, 6.720201e+09, 6.631664e+09, 6.542493e+09, 6.452746e+09, 
    6.362479e+09,
  6.319373e+09, 6.406312e+09, 6.492669e+09, 6.578392e+09, 6.663429e+09, 
    6.747724e+09, 6.831222e+09, 6.913867e+09, 6.9956e+09, 7.076365e+09, 
    7.1561e+09, 7.234745e+09, 7.312241e+09, 7.388526e+09, 7.463537e+09, 
    7.537212e+09, 7.60949e+09, 7.680307e+09, 7.749601e+09, 7.817309e+09, 
    7.883369e+09, 7.94772e+09, 8.010299e+09, 8.071048e+09, 8.129904e+09, 
    8.186811e+09, 8.241709e+09, 8.294543e+09, 8.345257e+09, 8.393798e+09, 
    8.440113e+09, 8.484152e+09, 8.525868e+09, 8.565214e+09, 8.602145e+09, 
    8.636621e+09, 8.668601e+09, 8.698051e+09, 8.724934e+09, 8.749221e+09, 
    8.770882e+09, 8.789891e+09, 8.806228e+09, 8.819871e+09, 8.830806e+09, 
    8.839017e+09, 8.844498e+09, 8.84724e+09, 8.84724e+09, 8.844498e+09, 
    8.839017e+09, 8.830806e+09, 8.819871e+09, 8.806228e+09, 8.789891e+09, 
    8.770882e+09, 8.749221e+09, 8.724934e+09, 8.698051e+09, 8.668601e+09, 
    8.636621e+09, 8.602145e+09, 8.565214e+09, 8.525868e+09, 8.484152e+09, 
    8.440113e+09, 8.393798e+09, 8.345257e+09, 8.294543e+09, 8.241709e+09, 
    8.186811e+09, 8.129904e+09, 8.071048e+09, 8.010299e+09, 7.94772e+09, 
    7.883369e+09, 7.817309e+09, 7.749601e+09, 7.680307e+09, 7.60949e+09, 
    7.537212e+09, 7.463537e+09, 7.388526e+09, 7.312241e+09, 7.234745e+09, 
    7.1561e+09, 7.076365e+09, 6.9956e+09, 6.913867e+09, 6.831222e+09, 
    6.747724e+09, 6.663429e+09, 6.578392e+09, 6.492669e+09, 6.406312e+09, 
    6.319373e+09,
  6.275223e+09, 6.35881e+09, 6.441759e+09, 6.52402e+09, 6.605544e+09, 
    6.686283e+09, 6.766183e+09, 6.845195e+09, 6.923265e+09, 7.000339e+09, 
    7.076365e+09, 7.151286e+09, 7.225049e+09, 7.297597e+09, 7.368877e+09, 
    7.438829e+09, 7.5074e+09, 7.574533e+09, 7.640172e+09, 7.704261e+09, 
    7.766745e+09, 7.827569e+09, 7.886679e+09, 7.94402e+09, 7.99954e+09, 
    8.053188e+09, 8.10491e+09, 8.15466e+09, 8.202386e+09, 8.248043e+09, 
    8.291585e+09, 8.332967e+09, 8.372148e+09, 8.409087e+09, 8.443745e+09, 
    8.476086e+09, 8.506077e+09, 8.533684e+09, 8.558878e+09, 8.581632e+09, 
    8.601922e+09, 8.619724e+09, 8.63502e+09, 8.647793e+09, 8.658028e+09, 
    8.665715e+09, 8.670843e+09, 8.673409e+09, 8.673409e+09, 8.670843e+09, 
    8.665715e+09, 8.658028e+09, 8.647793e+09, 8.63502e+09, 8.619724e+09, 
    8.601922e+09, 8.581632e+09, 8.558878e+09, 8.533684e+09, 8.506077e+09, 
    8.476086e+09, 8.443745e+09, 8.409087e+09, 8.372148e+09, 8.332967e+09, 
    8.291585e+09, 8.248043e+09, 8.202386e+09, 8.15466e+09, 8.10491e+09, 
    8.053188e+09, 7.99954e+09, 7.94402e+09, 7.886679e+09, 7.827569e+09, 
    7.766745e+09, 7.704261e+09, 7.640172e+09, 7.574533e+09, 7.5074e+09, 
    7.438829e+09, 7.368877e+09, 7.297597e+09, 7.225049e+09, 7.151286e+09, 
    7.076365e+09, 7.000339e+09, 6.923265e+09, 6.845195e+09, 6.766183e+09, 
    6.686283e+09, 6.605544e+09, 6.52402e+09, 6.441759e+09, 6.35881e+09, 
    6.275223e+09,
  6.230037e+09, 6.310255e+09, 6.38978e+09, 6.468569e+09, 6.546576e+09, 
    6.623755e+09, 6.700061e+09, 6.775447e+09, 6.849864e+09, 6.923265e+09, 
    6.9956e+09, 7.066822e+09, 7.136881e+09, 7.205726e+09, 7.273309e+09, 
    7.339579e+09, 7.404488e+09, 7.467984e+09, 7.530018e+09, 7.590542e+09, 
    7.649507e+09, 7.706863e+09, 7.762563e+09, 7.816561e+09, 7.868808e+09, 
    7.919261e+09, 7.967875e+09, 8.014606e+09, 8.059411e+09, 8.10225e+09, 
    8.143084e+09, 8.181873e+09, 8.218582e+09, 8.253174e+09, 8.285618e+09, 
    8.31588e+09, 8.343933e+09, 8.369748e+09, 8.3933e+09, 8.414565e+09, 
    8.433522e+09, 8.450151e+09, 8.464436e+09, 8.476363e+09, 8.485919e+09, 
    8.493095e+09, 8.497883e+09, 8.500278e+09, 8.500278e+09, 8.497883e+09, 
    8.493095e+09, 8.485919e+09, 8.476363e+09, 8.464436e+09, 8.450151e+09, 
    8.433522e+09, 8.414565e+09, 8.3933e+09, 8.369748e+09, 8.343933e+09, 
    8.31588e+09, 8.285618e+09, 8.253174e+09, 8.218582e+09, 8.181873e+09, 
    8.143084e+09, 8.10225e+09, 8.059411e+09, 8.014606e+09, 7.967875e+09, 
    7.919261e+09, 7.868808e+09, 7.816561e+09, 7.762563e+09, 7.706863e+09, 
    7.649507e+09, 7.590542e+09, 7.530018e+09, 7.467984e+09, 7.404488e+09, 
    7.339579e+09, 7.273309e+09, 7.205726e+09, 7.136881e+09, 7.066822e+09, 
    6.9956e+09, 6.923265e+09, 6.849864e+09, 6.775447e+09, 6.700061e+09, 
    6.623755e+09, 6.546576e+09, 6.468569e+09, 6.38978e+09, 6.310255e+09, 
    6.230037e+09,
  6.183825e+09, 6.260659e+09, 6.336752e+09, 6.412062e+09, 6.486551e+09, 
    6.560175e+09, 6.632894e+09, 6.704666e+09, 6.775447e+09, 6.845195e+09, 
    6.913867e+09, 6.981418e+09, 7.047806e+09, 7.112987e+09, 7.176916e+09, 
    7.23955e+09, 7.300845e+09, 7.360757e+09, 7.419243e+09, 7.47626e+09, 
    7.531766e+09, 7.585717e+09, 7.638074e+09, 7.688794e+09, 7.737838e+09, 
    7.785166e+09, 7.830739e+09, 7.874522e+09, 7.916475e+09, 7.956566e+09, 
    7.994759e+09, 8.031022e+09, 8.065324e+09, 8.097633e+09, 8.127923e+09, 
    8.156166e+09, 8.182336e+09, 8.20641e+09, 8.228367e+09, 8.248187e+09, 
    8.26585e+09, 8.281342e+09, 8.294647e+09, 8.305754e+09, 8.314652e+09, 
    8.321333e+09, 8.32579e+09, 8.32802e+09, 8.32802e+09, 8.32579e+09, 
    8.321333e+09, 8.314652e+09, 8.305754e+09, 8.294647e+09, 8.281342e+09, 
    8.26585e+09, 8.248187e+09, 8.228367e+09, 8.20641e+09, 8.182336e+09, 
    8.156166e+09, 8.127923e+09, 8.097633e+09, 8.065324e+09, 8.031022e+09, 
    7.994759e+09, 7.956566e+09, 7.916475e+09, 7.874522e+09, 7.830739e+09, 
    7.785166e+09, 7.737838e+09, 7.688794e+09, 7.638074e+09, 7.585717e+09, 
    7.531766e+09, 7.47626e+09, 7.419243e+09, 7.360757e+09, 7.300845e+09, 
    7.23955e+09, 7.176916e+09, 7.112987e+09, 7.047806e+09, 6.981418e+09, 
    6.913867e+09, 6.845195e+09, 6.775447e+09, 6.704666e+09, 6.632894e+09, 
    6.560175e+09, 6.486551e+09, 6.412062e+09, 6.336752e+09, 6.260659e+09, 
    6.183825e+09,
  6.136596e+09, 6.210038e+09, 6.282692e+09, 6.354524e+09, 6.425497e+09, 
    6.495574e+09, 6.564719e+09, 6.632894e+09, 6.700061e+09, 6.766183e+09, 
    6.831222e+09, 6.895139e+09, 6.957896e+09, 7.019455e+09, 7.079777e+09, 
    7.138825e+09, 7.196561e+09, 7.252946e+09, 7.307944e+09, 7.361518e+09, 
    7.41363e+09, 7.464245e+09, 7.513327e+09, 7.56084e+09, 7.606751e+09, 
    7.651027e+09, 7.693634e+09, 7.734541e+09, 7.773715e+09, 7.811129e+09, 
    7.846753e+09, 7.880559e+09, 7.912521e+09, 7.942612e+09, 7.970811e+09, 
    7.997093e+09, 8.021437e+09, 8.043825e+09, 8.064236e+09, 8.082655e+09, 
    8.099066e+09, 8.113456e+09, 8.125813e+09, 8.136126e+09, 8.144387e+09, 
    8.150589e+09, 8.154726e+09, 8.156796e+09, 8.156796e+09, 8.154726e+09, 
    8.150589e+09, 8.144387e+09, 8.136126e+09, 8.125813e+09, 8.113456e+09, 
    8.099066e+09, 8.082655e+09, 8.064236e+09, 8.043825e+09, 8.021437e+09, 
    7.997093e+09, 7.970811e+09, 7.942612e+09, 7.912521e+09, 7.880559e+09, 
    7.846753e+09, 7.811129e+09, 7.773715e+09, 7.734541e+09, 7.693634e+09, 
    7.651027e+09, 7.606751e+09, 7.56084e+09, 7.513327e+09, 7.464245e+09, 
    7.41363e+09, 7.361518e+09, 7.307944e+09, 7.252946e+09, 7.196561e+09, 
    7.138825e+09, 7.079777e+09, 7.019455e+09, 6.957896e+09, 6.895139e+09, 
    6.831222e+09, 6.766183e+09, 6.700061e+09, 6.632894e+09, 6.564719e+09, 
    6.495574e+09, 6.425497e+09, 6.354524e+09, 6.282692e+09, 6.210038e+09, 
    6.136596e+09,
  6.088361e+09, 6.158404e+09, 6.227619e+09, 6.295976e+09, 6.363442e+09, 
    6.429985e+09, 6.495574e+09, 6.560175e+09, 6.623755e+09, 6.686283e+09, 
    6.747724e+09, 6.808046e+09, 6.867216e+09, 6.925201e+09, 6.981969e+09, 
    7.037487e+09, 7.091722e+09, 7.144643e+09, 7.196217e+09, 7.246414e+09, 
    7.295202e+09, 7.342552e+09, 7.388432e+09, 7.432814e+09, 7.475667e+09, 
    7.516966e+09, 7.556683e+09, 7.594789e+09, 7.631261e+09, 7.666072e+09, 
    7.699199e+09, 7.73062e+09, 7.760311e+09, 7.788252e+09, 7.814423e+09, 
    7.838806e+09, 7.861382e+09, 7.882135e+09, 7.901051e+09, 7.918115e+09, 
    7.933316e+09, 7.946641e+09, 7.958081e+09, 7.967627e+09, 7.975273e+09, 
    7.981012e+09, 7.984841e+09, 7.986756e+09, 7.986756e+09, 7.984841e+09, 
    7.981012e+09, 7.975273e+09, 7.967627e+09, 7.958081e+09, 7.946641e+09, 
    7.933316e+09, 7.918115e+09, 7.901051e+09, 7.882135e+09, 7.861382e+09, 
    7.838806e+09, 7.814423e+09, 7.788252e+09, 7.760311e+09, 7.73062e+09, 
    7.699199e+09, 7.666072e+09, 7.631261e+09, 7.594789e+09, 7.556683e+09, 
    7.516966e+09, 7.475667e+09, 7.432814e+09, 7.388432e+09, 7.342552e+09, 
    7.295202e+09, 7.246414e+09, 7.196217e+09, 7.144643e+09, 7.091722e+09, 
    7.037487e+09, 6.981969e+09, 6.925201e+09, 6.867216e+09, 6.808046e+09, 
    6.747724e+09, 6.686283e+09, 6.623755e+09, 6.560175e+09, 6.495574e+09, 
    6.429985e+09, 6.363442e+09, 6.295976e+09, 6.227619e+09, 6.158404e+09, 
    6.088361e+09,
  6.039129e+09, 6.105772e+09, 6.171552e+09, 6.236442e+09, 6.300414e+09, 
    6.363442e+09, 6.425497e+09, 6.486551e+09, 6.546576e+09, 6.605544e+09, 
    6.663429e+09, 6.720201e+09, 6.775833e+09, 6.830297e+09, 6.883567e+09, 
    6.935614e+09, 6.986412e+09, 7.035934e+09, 7.084154e+09, 7.131045e+09, 
    7.176583e+09, 7.220742e+09, 7.263496e+09, 7.304823e+09, 7.344698e+09, 
    7.383099e+09, 7.420003e+09, 7.455388e+09, 7.489233e+09, 7.521518e+09, 
    7.552224e+09, 7.581331e+09, 7.608822e+09, 7.634681e+09, 7.65889e+09, 
    7.681435e+09, 7.702302e+09, 7.721477e+09, 7.738948e+09, 7.754704e+09, 
    7.768736e+09, 7.781033e+09, 7.791588e+09, 7.800395e+09, 7.807448e+09, 
    7.812741e+09, 7.816271e+09, 7.818037e+09, 7.818037e+09, 7.816271e+09, 
    7.812741e+09, 7.807448e+09, 7.800395e+09, 7.791588e+09, 7.781033e+09, 
    7.768736e+09, 7.754704e+09, 7.738948e+09, 7.721477e+09, 7.702302e+09, 
    7.681435e+09, 7.65889e+09, 7.634681e+09, 7.608822e+09, 7.581331e+09, 
    7.552224e+09, 7.521518e+09, 7.489233e+09, 7.455388e+09, 7.420003e+09, 
    7.383099e+09, 7.344698e+09, 7.304823e+09, 7.263496e+09, 7.220742e+09, 
    7.176583e+09, 7.131045e+09, 7.084154e+09, 7.035934e+09, 6.986412e+09, 
    6.935614e+09, 6.883567e+09, 6.830297e+09, 6.775833e+09, 6.720201e+09, 
    6.663429e+09, 6.605544e+09, 6.546576e+09, 6.486551e+09, 6.425497e+09, 
    6.363442e+09, 6.300414e+09, 6.236442e+09, 6.171552e+09, 6.105772e+09, 
    6.039129e+09,
  5.988909e+09, 6.052155e+09, 6.114508e+09, 6.175945e+09, 6.236442e+09, 
    6.295976e+09, 6.354524e+09, 6.412062e+09, 6.468569e+09, 6.52402e+09, 
    6.578392e+09, 6.631664e+09, 6.683811e+09, 6.734811e+09, 6.784643e+09, 
    6.833284e+09, 6.880711e+09, 6.926904e+09, 6.971842e+09, 7.015503e+09, 
    7.057866e+09, 7.098912e+09, 7.13862e+09, 7.176973e+09, 7.21395e+09, 
    7.249533e+09, 7.283705e+09, 7.316448e+09, 7.347746e+09, 7.377583e+09, 
    7.405943e+09, 7.432813e+09, 7.458176e+09, 7.482021e+09, 7.504335e+09, 
    7.525106e+09, 7.544322e+09, 7.561974e+09, 7.578052e+09, 7.592547e+09, 
    7.605452e+09, 7.616759e+09, 7.626462e+09, 7.634556e+09, 7.641037e+09, 
    7.645901e+09, 7.649145e+09, 7.650767e+09, 7.650767e+09, 7.649145e+09, 
    7.645901e+09, 7.641037e+09, 7.634556e+09, 7.626462e+09, 7.616759e+09, 
    7.605452e+09, 7.592547e+09, 7.578052e+09, 7.561974e+09, 7.544322e+09, 
    7.525106e+09, 7.504335e+09, 7.482021e+09, 7.458176e+09, 7.432813e+09, 
    7.405943e+09, 7.377583e+09, 7.347746e+09, 7.316448e+09, 7.283705e+09, 
    7.249533e+09, 7.21395e+09, 7.176973e+09, 7.13862e+09, 7.098912e+09, 
    7.057866e+09, 7.015503e+09, 6.971842e+09, 6.926904e+09, 6.880711e+09, 
    6.833284e+09, 6.784643e+09, 6.734811e+09, 6.683811e+09, 6.631664e+09, 
    6.578392e+09, 6.52402e+09, 6.468569e+09, 6.412062e+09, 6.354524e+09, 
    6.295976e+09, 6.236442e+09, 6.175945e+09, 6.114508e+09, 6.052155e+09, 
    5.988909e+09,
  5.937712e+09, 5.99757e+09, 6.056508e+09, 6.114508e+09, 6.171552e+09, 
    6.227619e+09, 6.282692e+09, 6.336752e+09, 6.38978e+09, 6.441759e+09, 
    6.492669e+09, 6.542493e+09, 6.591213e+09, 6.638811e+09, 6.685269e+09, 
    6.730571e+09, 6.774699e+09, 6.817636e+09, 6.859367e+09, 6.899874e+09, 
    6.939143e+09, 6.977157e+09, 7.013901e+09, 7.049361e+09, 7.083523e+09, 
    7.116371e+09, 7.147894e+09, 7.178077e+09, 7.206909e+09, 7.234377e+09, 
    7.260469e+09, 7.285175e+09, 7.308484e+09, 7.330385e+09, 7.350871e+09, 
    7.36993e+09, 7.387556e+09, 7.403741e+09, 7.418477e+09, 7.431758e+09, 
    7.443579e+09, 7.453934e+09, 7.462817e+09, 7.470226e+09, 7.476158e+09, 
    7.480609e+09, 7.483577e+09, 7.485062e+09, 7.485062e+09, 7.483577e+09, 
    7.480609e+09, 7.476158e+09, 7.470226e+09, 7.462817e+09, 7.453934e+09, 
    7.443579e+09, 7.431758e+09, 7.418477e+09, 7.403741e+09, 7.387556e+09, 
    7.36993e+09, 7.350871e+09, 7.330385e+09, 7.308484e+09, 7.285175e+09, 
    7.260469e+09, 7.234377e+09, 7.206909e+09, 7.178077e+09, 7.147894e+09, 
    7.116371e+09, 7.083523e+09, 7.049361e+09, 7.013901e+09, 6.977157e+09, 
    6.939143e+09, 6.899874e+09, 6.859367e+09, 6.817636e+09, 6.774699e+09, 
    6.730571e+09, 6.685269e+09, 6.638811e+09, 6.591213e+09, 6.542493e+09, 
    6.492669e+09, 6.441759e+09, 6.38978e+09, 6.336752e+09, 6.282692e+09, 
    6.227619e+09, 6.171552e+09, 6.114508e+09, 6.056508e+09, 5.99757e+09, 
    5.937712e+09,
  5.885548e+09, 5.942029e+09, 5.99757e+09, 6.052155e+09, 6.105772e+09, 
    6.158404e+09, 6.210038e+09, 6.260659e+09, 6.310255e+09, 6.35881e+09, 
    6.406312e+09, 6.452746e+09, 6.4981e+09, 6.54236e+09, 6.585513e+09, 
    6.627547e+09, 6.668449e+09, 6.708208e+09, 6.74681e+09, 6.784244e+09, 
    6.8205e+09, 6.855565e+09, 6.889429e+09, 6.922081e+09, 6.953512e+09, 
    6.98371e+09, 7.012667e+09, 7.040374e+09, 7.066821e+09, 7.092e+09, 
    7.115902e+09, 7.138521e+09, 7.159848e+09, 7.179877e+09, 7.198601e+09, 
    7.216014e+09, 7.23211e+09, 7.246883e+09, 7.260329e+09, 7.272444e+09, 
    7.283223e+09, 7.292662e+09, 7.30076e+09, 7.307511e+09, 7.312915e+09, 
    7.316969e+09, 7.319673e+09, 7.321026e+09, 7.321026e+09, 7.319673e+09, 
    7.316969e+09, 7.312915e+09, 7.307511e+09, 7.30076e+09, 7.292662e+09, 
    7.283223e+09, 7.272444e+09, 7.260329e+09, 7.246883e+09, 7.23211e+09, 
    7.216014e+09, 7.198601e+09, 7.179877e+09, 7.159848e+09, 7.138521e+09, 
    7.115902e+09, 7.092e+09, 7.066821e+09, 7.040374e+09, 7.012667e+09, 
    6.98371e+09, 6.953512e+09, 6.922081e+09, 6.889429e+09, 6.855565e+09, 
    6.8205e+09, 6.784244e+09, 6.74681e+09, 6.708208e+09, 6.668449e+09, 
    6.627547e+09, 6.585513e+09, 6.54236e+09, 6.4981e+09, 6.452746e+09, 
    6.406312e+09, 6.35881e+09, 6.310255e+09, 6.260659e+09, 6.210038e+09, 
    6.158404e+09, 6.105772e+09, 6.052155e+09, 5.99757e+09, 5.942029e+09, 
    5.885548e+09,
  5.832426e+09, 5.885548e+09, 5.937712e+09, 5.988909e+09, 6.039129e+09, 
    6.088361e+09, 6.136596e+09, 6.183825e+09, 6.230037e+09, 6.275223e+09, 
    6.319373e+09, 6.362479e+09, 6.404531e+09, 6.445522e+09, 6.485442e+09, 
    6.524282e+09, 6.562035e+09, 6.598693e+09, 6.634248e+09, 6.668692e+09, 
    6.702019e+09, 6.734221e+09, 6.76529e+09, 6.795221e+09, 6.824007e+09, 
    6.851641e+09, 6.878117e+09, 6.903431e+09, 6.927576e+09, 6.950547e+09, 
    6.972339e+09, 6.992947e+09, 7.012366e+09, 7.030593e+09, 7.047623e+09, 
    7.063453e+09, 7.078078e+09, 7.091497e+09, 7.103705e+09, 7.1147e+09, 
    7.124479e+09, 7.133041e+09, 7.140384e+09, 7.146505e+09, 7.151404e+09, 
    7.155078e+09, 7.157529e+09, 7.158754e+09, 7.158754e+09, 7.157529e+09, 
    7.155078e+09, 7.151404e+09, 7.146505e+09, 7.140384e+09, 7.133041e+09, 
    7.124479e+09, 7.1147e+09, 7.103705e+09, 7.091497e+09, 7.078078e+09, 
    7.063453e+09, 7.047623e+09, 7.030593e+09, 7.012366e+09, 6.992947e+09, 
    6.972339e+09, 6.950547e+09, 6.927576e+09, 6.903431e+09, 6.878117e+09, 
    6.851641e+09, 6.824007e+09, 6.795221e+09, 6.76529e+09, 6.734221e+09, 
    6.702019e+09, 6.668692e+09, 6.634248e+09, 6.598693e+09, 6.562035e+09, 
    6.524282e+09, 6.485442e+09, 6.445522e+09, 6.404531e+09, 6.362479e+09, 
    6.319373e+09, 6.275223e+09, 6.230037e+09, 6.183825e+09, 6.136596e+09, 
    6.088361e+09, 6.039129e+09, 5.988909e+09, 5.937712e+09, 5.885548e+09, 
    5.832426e+09 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01253, 0.04887, 0.10724, 0.18455, 0.27461, 0.36914, 
    0.46103, 0.54623, 0.62305, 0.69099, 0.75016, 0.8011, 0.84453, 0.88125, 
    0.9121, 0.93766, 0.95849, 0.97495, 0.98743, 0.9958, 1 ;

 pk = 1, 2.69722, 5.17136, 8.89455, 14.2479, 22.07157, 33.61283, 50.48096, 
    74.79993, 109.4006, 158.0046, 225.4411, 317.8956, 443.1935, 611.1156, 
    833.7439, 1125.834, 1505.208, 1993.158, 2614.863, 3399.784, 4382.062, 
    5600.87, 7100.731, 8931.782, 11149.97, 13817.17, 17001.21, 20775.82, 
    23967.34, 25527.65, 25671.22, 24609.3, 22640.51, 20147.13, 17477.63, 
    14859.86, 12414.93, 10201.44, 8241.503, 6534.432, 5066.179, 3815.607, 
    2758.603, 1880.646, 1169.339, 618.4799, 225, 10, 0 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.9037046, 1, 1, 0.8371245, 0.01079098, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.342301, 1, 0.9242505, 0.2324802, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1585782, 0.8988085, 0.872375, 0.8199701, 0.2036715, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04788778, 0.3358625, 0.07239318, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1174253, 0.1658257, 0.1069185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.04039344, 0.2727596, 0.3044432, 0.03935189, 0.05927679, 
    0.5426623, 0.5088302, 0.241054, 0.0411321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04967177, 0.09058292, 0.6336873, 0.9864414, 1, 0.999317, 0.9606841, 
    0.9469818, 1, 1, 1, 0.9701587, 0.6985948, 0.1660634, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04887224, 0.4892108, 0.9759328, 0.8929602, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9605891, 0.1742972, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1475878, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2927403, 
    0.1056596, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008395956, 0.8062803, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7915943, 0.001058526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003862719, 0.7844364, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4460433, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3652394, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9193342, 
    0.1419819, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2822479, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9971261, 
    0.6570057, 0.2192735, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08952717, 0.2009808, 0.4916342, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.4641593, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02373972, 
    0.2887375, 0.5454076, 0.7591597, 0.9840837, 0.9225589, 0.9569725, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2276618, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01343125, 0.2130994, 0.07166115, 
    0.1361981, 0.4062145, 0.4764926, 0.9131937, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9399245, 0.2953852, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1096427, 0.6468607, 1, 0.9679646, 
    0.8867931, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.9742239, 0.2603416, 0.000543013, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006295154, 0.4813343, 0.944672, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.811202, 0.007860967, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.3256565, 0.3595797, 0.9921021, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8934381, 0.4007365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.5127948, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8029071, 0.1827247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8530139, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6570168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0181968, 0.8725816, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7388504, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1284515, 0.9620806, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8478313, 0.01794271, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.05491119, 0.6775094, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9972597, 0.1556571, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01809847, 0.02063968, 0.5821294, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.576636, 0.0007413209, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.5811512, 0.770504, 0.5899364, 0.7125399, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9348087, 0.3177032, 0.05322447, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.7359381, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9021191, 
    0.3398403, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2397476, 0.9484219, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9444426, 0.1523203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7934542, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9452199, 
    0.4845907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.4458613, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7567984, 
    0.06867129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0058354, 0.4173073, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.4904585, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0734878, 
    0.0544353, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.3889154, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3997353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0560805, 0.6384699, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.297665, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0808603, 0.2136603, 0.223731, 0.7629656, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.1250296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1126087, 0.07242998, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.06437702, 0.4854095, 0.7614139, 0.9957509, 0.9980491, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.1323143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4987842, 0.4307159, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1129699, 0.7654874, 1, 1, 1, 1, 0.9594662, 0.2817145, 
    0.349315, 0.4800343, 0.4166909, 0.33321, 0.8587425, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5030489, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.208195, 
    0.3201258, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1805963, 0.4938805, 0.9619426, 1, 1, 0.9977201, 0.4028112, 
    0, 0, 0, 0, 0, 0.03760567, 0.4765331, 0.9889686, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6693374, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1330605, 0.07577454, 0.6408337, 1, 1, 0.8560842, 0.229482, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.7420933, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9711934, 0.8154297, 0.7031593, 0.1591314, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2664649, 0.9408039, 1, 0.9731776, 0.3734872, 0.08581278, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2477078, 0.9847024, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9874682, 0.6629098, 0.03976496, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.04098084, 0.6700594, 1, 0.9846117, 0.3915779, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002308619, 0.8402424, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9393559, 0.3334898, 0.4927699, 0.1729504, 
    0.0005183411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.05815923, 0.8921363, 0.9963881, 0.4196884, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.03001891, 0.8732678, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8185688, 0.000997816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3599489, 0.6536069, 0.2308225, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1388849, 0.9886107, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8995878, 0.6226335, 0.6108878, 0.388907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.275672, 0.4499452, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6206766, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6265669, 0.03419805, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004062632, 0.09197545, 0.07587977, 
    0.1429734, 0.07793289, 0.001982026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.09490187, 0.1736679, 0.3527791, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001625569, 0.2624141, 0.8962197, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9966809, 0.5754746, 0.03894359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2468218, 0.5043563, 0.9838024, 0.866147, 
    0.8783621, 0.9815187, 0.8271396, 0.4878259, 0.01884565, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1005597, 0.06768002, 0.1576353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.33927, 0.891219, 0.9995848, 1, 1, 0.9420939, 
    0.7670357, 0.6221464, 0.2302634, 0.2723061, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1477103, 0.6884276, 0.999054, 1, 1, 1, 0.7532653, 
    0.5085074, 0.8721771, 1, 0.3210266, 0, 0, 0, 0, 0, 0, 0, 0, 0.05677235, 
    0.0008144492, 0.04120899, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1219508, 0.1550475, 0.3309695, 0.0581816, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 2.639958e-05, 0, 0.7161255, 1, 1, 1, 1, 1, 0.7215892, 
    0.7704202, 0.9905617, 0.9987394, 0.5821542, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04867533, 0.01442351, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.04097006, 0.593925, 0.648534, 0.9974784, 1, 1, 1, 1, 
    0.999142, 0.6332727, 0.257304, 0.1315637, 0.1783369, 0.4090085, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006319822, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0159371, 0.6464633, 1, 1, 1, 1, 1, 1, 0.9379096, 0.3084929, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.05427543, 0.8169017, 1, 1, 1, 1, 1, 1, 1, 0.6480082, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0.0001631903, 0.2342296, 0.3217961, 1, 1, 1, 1, 1, 1, 1, 0.9198062, 
    0.2241177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.6364967, 0.4618171, 0.704794, 1, 1, 1, 1, 1, 1, 1, 0.4258353, 0, 0, 0, 0, 
    0, 0.01590484, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.5118697, 0.9346247, 1, 1, 1, 1, 1, 0.9876335, 0.9329823, 0.9783548, 
    0.2976481, 0, 0, 0, 0, 0.01003709, 0.4619169, 0.1022752, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.9873409, 0.253808, 0.04543634, 0.5278371, 0.002404106, 
    0, 0, 0, 0, 0.003275408, 0.6632224, 0.3422698, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.7803705, 0.005725726, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03397798, 0.01880223, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.6511014, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 0.9937965, 0.1486441, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 0.9887101, 0.3117075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.9908476, 0.4261142, 0.01644797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09772249, 0.07365502, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.7445699, 0.1342526, 0.4569494, 0.0158662, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01797347, 0.3693104, 
    0.01717718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4015935, 0.05133266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 0.9750558, 0.2528034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 0.6344764, 0.008912468, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.8986811, 0.1816702, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.2968034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.8290737, 0.01273574, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.8303954, 0.01862913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.9919094, 0.1766838, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.9953394, 0.2376448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.6380026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.6356525, 0.1226215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 orog =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7992414, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2732799, 355.3445, 661.6653, 788.604, 538.0593, 35.1188, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.84651, 302.8979, 366.1382, 
    37.41038, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39.91399, 196.7844, 215.7041, 248.1746, 36.99986, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9039114, 78.54595, 10.11436, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.704782, 26.12457, 13.85557, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005312768, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.02989985, 0.0003766294, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4189242, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1030456, 1.054963, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.143771, 12.69478, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.836948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.310095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01557077, 4.43028, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0002689204, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7.815726, 77.31487, 37.02573, 24.40091, 17.92381, 71.63206, 
    255.5557, 112.1054, 8.874227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.931261, 18.36737, 547.9603, 983.4506, 928.882, 805.4354, 755.1304, 
    606.848, 760.251, 1122.059, 1210.754, 926.5558, 393.9966, 77.59235, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18.74462, 550.8997, 873.0414, 738.3782, 1447.062, 1752.654, 1555.512, 
    1427.795, 1463.065, 1405.852, 1591.613, 1837.372, 1954.355, 1766.622, 
    1318.124, 785.6111, 74.99232, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97.7004, 1316.783, 1765.13, 1515.387, 1988.113, 2090.078, 1944.169, 
    1852.772, 1877.534, 1980.513, 2136.833, 2321.126, 2360.485, 2221.856, 
    1762.722, 1079.052, 99.97397, 6.346212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.179383, 841.1734, 1729.189, 2051.514, 2252.923, 2277.749, 2199.887, 
    2128.035, 2119.189, 2210.886, 2389.87, 2514.411, 2530.765, 2387.412, 
    2038.683, 1570.642, 1014.397, 440.8733, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.362782, 1003.385, 1800.715, 2229.933, 2275.979, 2360.229, 2311.384, 
    2315.582, 2392.034, 2497.806, 2647.774, 2647.349, 2549.216, 2306.825, 
    2075.641, 1693.824, 991.6838, 61.70815, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    118.7808, 1369.103, 1878.122, 2249.811, 2418.137, 2469.63, 2522.086, 
    2576.791, 2679.619, 2804.705, 2853.611, 2761.156, 2575.387, 2356.625, 
    2033.336, 1327.755, 445.6916, 5.287508, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3446125, 116.4755, 1433.451, 2040.093, 2321.82, 2502.561, 2570.579, 
    2649.61, 2757.851, 2852.799, 3005.241, 3050.789, 2945.686, 2746.585, 
    2492.519, 2133.578, 1679.148, 958.2936, 281.5658, 332.4458, 79.20005, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    159.5307, 500.1543, 1869.062, 2316.033, 2462.074, 2542.433, 2621.507, 
    2731.679, 2849.691, 2997.048, 3129.562, 3153.165, 3042.124, 2822.781, 
    2579.193, 2313.826, 1938.037, 1456.275, 955.3979, 723.9649, 233.088, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87.2196, 982.8452, 2074.387, 2401.657, 2479.505, 2552.033, 2644.845, 
    2764.61, 2913.177, 3071.668, 3188.252, 3187.021, 3067.563, 2877.698, 
    2677.985, 2453.64, 2217.535, 1895.206, 1415.486, 987.4891, 102.9291, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.006072, 9.248502, 51.24354, 
    117.7083, 0, 0, 0, 0, 0, 0, 1.781354, 493.788, 1756.028, 2232.431, 
    2436.472, 2528.297, 2640.581, 2788.757, 2970.408, 3126.261, 3223.229, 
    3201.013, 3098.396, 2951.579, 2787.688, 2644.104, 2469.223, 2265.754, 
    2020.998, 1603.012, 1036.609, 247.5821, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37.27396, 324.1435, 484.3052, 107.4387, 
    334.8317, 258.5734, 18.40336, 45.59911, 0, 0, 0, 0, 0, 312.953, 1500.18, 
    2183.505, 2342.897, 2491.774, 2647.206, 2829.54, 3007.807, 3145.192, 
    3213.799, 3194.5, 3103.396, 2991.563, 2858.539, 2725.452, 2602.863, 
    2442.798, 2299.817, 2079.573, 1678.872, 960.7639, 59.84979, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9005052, 143.1917, 891.4856, 1319.249, 
    1183.058, 743.5308, 625.7929, 271.4628, 29.0506, 28.26866, 0, 0, 0, 0, 0, 
    717.5844, 1521.244, 1982.313, 2315.337, 2501.919, 2714.457, 2879.019, 
    3038.052, 3144.582, 3199.439, 3176.925, 3090.616, 2991.669, 2897.744, 
    2785.427, 2687.85, 2575.268, 2434.927, 2202.157, 1748.342, 990.5164, 
    59.45817, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 138.0944, 28.26443, 859.6864, 1666.731, 1924.49, 
    1504.685, 894.1763, 626.5555, 183.7074, 1.250475, 6.993803, 0, 0, 0, 0, 
    152.5896, 1363.213, 1888.575, 2229.896, 2403.91, 2606.387, 2805.63, 
    2949.473, 3072.477, 3182.144, 3236.154, 3219.5, 3134.394, 3083.353, 
    3023.675, 2942.66, 2840.365, 2713.65, 2525.043, 2247.123, 1760.282, 
    1015.293, 69.54496, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 54.8675, 364.3715, 1548.06, 2161.363, 1988.979, 
    1423.904, 840.0815, 473.7389, 230.111, 231.5213, 70.41041, 0, 0, 0, 
    53.0154, 1249.682, 2001.559, 2304.354, 2429.361, 2548.836, 2707.271, 
    2894.569, 3029.046, 3159.696, 3279.65, 3330.228, 3323.386, 3284.032, 
    3259.254, 3244.029, 3164.147, 3039.184, 2858.268, 2653.644, 2425.572, 
    2034.225, 1328.45, 212.7939, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 138.5299, 947.9814, 1887.259, 2160.271, 1846.834, 
    1415.143, 971.5607, 604.7406, 412.5479, 333.2895, 159.8654, 26.29184, 
    1.857185, 274.4556, 1131.609, 1924.803, 2423.259, 2540.296, 2611.256, 
    2717.599, 2832.219, 2998.016, 3149.23, 3272.842, 3375.903, 3453.881, 
    3472.483, 3466.487, 3455.854, 3431.323, 3360.251, 3219.655, 3025.667, 
    2818.918, 2574.498, 2177.516, 1541.304, 418.2077, 3.786927, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.897408, 278.9847, 1150.151, 1820.023, 1906.937, 
    1710.571, 1470.08, 1188.798, 854.9822, 594.4963, 455.2799, 296.2944, 
    20.74247, 212.9633, 1377.01, 2210.266, 2531.037, 2589.832, 2729.739, 
    2779.357, 2870.47, 2960.67, 3105.383, 3254.163, 3365.769, 3484.833, 
    3561.692, 3602.843, 3610.362, 3592.779, 3537.574, 3466.485, 3340.572, 
    3139.534, 2890.738, 2605.906, 2178.262, 1557.431, 585.7548, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25.96501, 274.0147, 1064.936, 1482.375, 1656.331, 
    1647.515, 1562.002, 1335.74, 1001.996, 734.4821, 565.3111, 391.8153, 
    311.9492, 871.4916, 2073.987, 2854.189, 2770.159, 2864.382, 2882.136, 
    2935.086, 3016.186, 3112.14, 3232.739, 3376.769, 3504.886, 3614.249, 
    3695.932, 3704.89, 3713.67, 3686.838, 3614.497, 3529.63, 3396.464, 
    3164.898, 2869.117, 2545.209, 2079.768, 1444.332, 473.3306, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.198395, 148.0527, 886.8211, 1277.724, 1493.68, 
    1692.014, 1690.58, 1503.016, 1205.435, 994.3757, 848.381, 968.3361, 
    1305.293, 1773.208, 2657.443, 2950.178, 3028.504, 2998.262, 3013.121, 
    3056.479, 3144.256, 3246.656, 3377.553, 3516.235, 3644.559, 3743.524, 
    3749.271, 3708.808, 3678.306, 3622.363, 3548.655, 3468.685, 3334.021, 
    3096.724, 2813.21, 2507.742, 2064.155, 1345.841, 332.7528, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.602107, 0.03367292, 82.96276, 823.9019, 1207.387, 
    1490.124, 1792.475, 1887.241, 1801.419, 1641.348, 1457.016, 1489.465, 
    1791.969, 2173.656, 2577.651, 2800.211, 3040.854, 3063.57, 3082.433, 
    3086.433, 3130.878, 3234.532, 3374.836, 3510.101, 3641.93, 3775.546, 
    3826.162, 3739.047, 3612.842, 3507.702, 3436.104, 3394.341, 3313.844, 
    3186.941, 2981.263, 2736.921, 2428.213, 1957.258, 1192.974, 155.4329, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 87.60106, 73.32498, 112.404, 153.6019, 823.2629, 1290.737, 
    1591.929, 1899.596, 2085.203, 2131.1, 2032.692, 1952.935, 2003.027, 
    2256.183, 2444.568, 2635.164, 2807.364, 2928.302, 2931.476, 3038.824, 
    3101.363, 3169.576, 3315.562, 3484.013, 3647.621, 3791.786, 3922.948, 
    3926.845, 3723.422, 3456.011, 3269.509, 3160.537, 3127.081, 3060.512, 
    2938.832, 2773.188, 2564.738, 2217.429, 1614.816, 876.0974, 3.817307, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 174.1339, 192.5289, 595.6072, 548.1959, 902.9622, 
    1324.524, 1637.417, 1968.1, 2162.593, 2136.62, 2034.022, 1937.629, 
    2005.565, 1973.358, 2069.837, 2373.308, 2690.74, 2792.308, 2870.053, 
    3000.035, 3104.013, 3210.098, 3377.595, 3564.663, 3770.401, 3917.039, 
    4012.642, 3948.944, 3671.559, 3324.181, 3003.464, 2810.002, 2744.527, 
    2678.826, 2554.504, 2450.903, 2248.528, 1666.047, 879.4138, 217.8605, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41.24575, 171.1755, 928.2092, 911.556, 1003.465, 1333.517, 
    1742.872, 1976.593, 1971.419, 1847.775, 1596.083, 1517.469, 1510.441, 
    1449.914, 1648.969, 2160.01, 2465.792, 2611.214, 2691.124, 2869.434, 
    3045.968, 3236.557, 3398.76, 3579.36, 3797.204, 3936.64, 3975.402, 
    3863.231, 3599.677, 3223.608, 2813.848, 2505.323, 2321.725, 2250.189, 
    2064.987, 1902.286, 1638.834, 1019.027, 91.78241, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 105.7556, 967.28, 1137.105, 1125.491, 1369.858, 
    1526.296, 1610.441, 1462.915, 1195.448, 979.7076, 964.7514, 1033.812, 
    1020.986, 1503.457, 1979.614, 2248.812, 2429.502, 2603.554, 2766.973, 
    2963.375, 3182.582, 3375.808, 3529.749, 3729.817, 3856.099, 3884.153, 
    3740.839, 3498.397, 3131.312, 2677.872, 2252.273, 1934.652, 1693.907, 
    1330.782, 934.9443, 600.6172, 199.5566, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.739202, 0, 0, 0, 56.65801, 764.7597, 1177.214, 1137.807, 
    867.6033, 751.4905, 455.4625, 373.3823, 389.2663, 356.8941, 412.8959, 
    422.8545, 839.1047, 1290.905, 1814.671, 2116.265, 2387.323, 2578.228, 
    2692.938, 2810.998, 3018.81, 3251.787, 3454.09, 3636.555, 3767.025, 
    3772.435, 3602.902, 3361.617, 3049.529, 2649.456, 2152.187, 1589.401, 
    1095.306, 616.2491, 204.8285, 109.602, 22.18781, 48.89778, 9.825142, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009279916, 251.9048, 962.301, 883.4589, 677.3438, 
    361.7939, 137.7333, 20.846, 41.77541, 29.66083, 35.41616, 248.8549, 
    735.1519, 1335.172, 1731.033, 2074.124, 2359.61, 2570.465, 2604.922, 
    2667.29, 2813.544, 3063.244, 3317.592, 3564.776, 3708.774, 3713.399, 
    3546.005, 3335.875, 3064.894, 2726.397, 2302.653, 1790.918, 1349.976, 
    1108.172, 1070.336, 1060.536, 925.6852, 754.9511, 214.2521, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23.60169, 0.001468251, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 112.4058, 711.1246, 782.2984, 371.9018, 202.2023, 
    4.081332, 19.38192, 1.332851, 0.4524727, 2.236566, 63.69951, 569.4813, 
    1187.416, 1604.718, 1946.94, 2248.886, 2439.147, 2533.595, 2566.406, 
    2670.604, 2904.311, 3214.155, 3497.722, 3662.987, 3690.172, 3581.76, 
    3430.937, 3210.368, 2925.982, 2596.184, 2305.98, 2085.327, 1988.169, 
    1999.194, 2000.523, 1668.639, 1237.938, 193.779, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0277722, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.159892, 56.1418, 452.5438, 1005.819, 940.8052, 
    359.2229, 45.87414, 0.6317925, -4.440892e-16, 0.4750352, 33.37933, 
    3.9842, 295.6864, 921.4279, 1533.577, 1758.771, 2015.291, 2243.664, 
    2363.067, 2499.792, 2603.064, 2851.553, 3174.852, 3439.871, 3601.986, 
    3639.036, 3611.236, 3520.832, 3376.327, 3171.316, 2925.103, 2754.788, 
    2670.149, 2638.344, 2562.51, 2441.751, 2061.093, 1274.259, 129.2553, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 40.98916, 47.87557, 244.1692, 1334.147, 1438.746, 
    508.3959, 23.03855, -1.734723e-18, 0, 10.75564, 254.7662, 148.7082, 
    109.2365, 659.3992, 1310.688, 1593.068, 1868.237, 2051.256, 2239.637, 
    2436.269, 2622.957, 2896.737, 3180.859, 3412.578, 3564.607, 3677.027, 
    3686.917, 3618.097, 3508.476, 3355.026, 3184.518, 3051.357, 3012.698, 
    2935.528, 2832.188, 2615.409, 2041.958, 1159, 32.8907, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.57209, 3.683461, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13.15392, 21.53556, 145.4484, 166.8116, 212.421, 1456.922, 
    1442.133, 274.9966, 0, 0, 0.3660825, 97.71632, 274.119, 216.5157, 
    1.421085e-14, 355.3852, 921.0424, 1435.383, 1760.988, 2009.327, 2226.052, 
    2488.684, 2725.142, 2982.086, 3207.749, 3389.718, 3565.573, 3709.347, 
    3742.948, 3657.837, 3548.883, 3403.997, 3227.927, 3100.738, 3010.48, 
    2897.043, 2753.1, 2530.298, 1963.905, 996.7645, 20.1157, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 95.68005, 62.03844, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76.78776, 251.8225, 365.1784, 499.3779, 679.7224, 1282.687, 
    976.8096, 54.30797, 0, 0, -4.440892e-16, 3.06115, 105.1266, 7.105427e-15, 
    146.4528, 166.1453, 740.5073, 1156.732, 1667.2, 2071.25, 2311.511, 
    2561.432, 2802.865, 3051.193, 3239.81, 3403.32, 3577.332, 3697.356, 
    3695.489, 3575.418, 3467.606, 3301.877, 3080.048, 2891.024, 2773.609, 
    2640.24, 2458.685, 2296.196, 1776.581, 1080.293, 215.078, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20.15371, 42.59801, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 132.3908, 427.5094, 871.1767, 1216.166, 1215.606, 1074.381, 
    143.933, 0, 0, 0, 0, 4.440892e-16, 0.7024416, 85.66618, 422.4643, 
    753.0161, 876.0609, 1329.78, 1707.256, 2086.016, 2393.784, 2545.285, 
    2840.856, 3071.359, 3268.794, 3422.524, 3586.531, 3666.174, 3565.691, 
    3397.146, 3270.382, 3125.957, 2841.437, 2580.784, 2474.215, 2351.78, 
    2078.684, 1727.895, 1498.923, 1140.002, 539.2833, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 62.32169, 39.41545, 626.6343, 1371.758, 1347.847, 687.8185, 
    32.66976, 0, 0, 0, 0, 0, 0, -6.938894e-18, 29.09192, 611.8069, 1072.647, 
    1446.324, 1597.489, 1872.625, 2189.95, 2396.317, 2632.638, 2864.967, 
    3116.256, 3290.928, 3442.491, 3576.208, 3595.495, 3416.291, 3130.265, 
    2946.176, 2774.498, 2500.969, 2090.21, 2070.135, 2101.286, 1651.494, 
    934.1992, 472.3446, 447.5172, 68.89008, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 239.6809, 554.4179, 364.8323, 498.6555, 95.83427, 6.607563, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 132.7997, 1047.2, 1417.112, 1781.415, 2066.203, 
    2268.176, 2513.788, 2702.935, 2989.756, 3186.11, 3356.546, 3463.798, 
    3540.333, 3487.458, 3305.011, 2838.596, 2431.235, 2225.709, 1948.767, 
    1463.512, 1303.707, 1487.188, 1115.347, 344.4456, 17.17711, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.06872149, 590.6149, 255.9139, 0.4632595, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 187.6016, 678.9084, 1330.984, 2035.844, 2433.294, 
    2612.385, 2832.168, 3016.011, 3219.117, 3378.409, 3442.958, 3400.81, 
    3281.248, 3011.857, 2341.452, 1747.214, 1505.163, 1297.308, 751.0115, 
    196.1539, 377.1983, 100.9759, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 38.59026, 645.7719, 34.58854, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53.31918, 810.9399, 1739.455, 2404.192, 2757.1, 2846.992, 
    2957.257, 3148.64, 3318.68, 3306.222, 3091.919, 2659.991, 2079.938, 
    1357.805, 792.2961, 628.3082, 498.0571, 246.4902, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 235.8719, 404.9598, 19.19321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1208589, 268.1322, 1044.283, 1926.036, 2449.009, 2629.04, 
    2630.753, 3113.425, 3114.51, 2984.559, 2508.903, 1782.817, 1010.823, 
    372.2121, 24.88615, 0.03625189, 0.009416752, 86.38479, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14.21238, 250.7785, 295.3082, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 155.7787, 592.4962, 1366.038, 1963.625, 1825.582, 2069.24, 
    2485.683, 2492.135, 2126.706, 1540.313, 896.8804, 239.871, 46.3145, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.80038, 14.7334, 38.18274, 15.65409, 
    2.098015, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.28813, 129.1734, 304.9514, 
    3.314995, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 149.1334, 
    773.5136, 1044.637, 889.3293, 853.0041, 1272.865, 1052.722, 795.8773, 
    379.6655, 140.3403, 5.892643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.09859627, 30.3471, 81.51091, 108.4727, 153.5919, 
    206.7384, 204.1187, 155.7402, 96.83952, 3.76339, 0, 0, 0, 0, 0, 0, 0, 0, 
    19.27378, 11.65506, 100.7927, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26.58224, 97.38688, 141.9256, 27.09244, 26.51507, 114.4799, 
    79.36494, 31.06278, 0, 0.04206881, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 26.76524, 161.1405, 374.7367, 504.8459, 444.2382, 
    263.0925, 173.7267, 155.3289, 255.5945, 377.7833, 81.20056, 2.50277, 0, 
    0, 0, 0, 0, 0, 0, 19.48863, 0, 17.85832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 17.59249, 7.557294, 179.5778, 668.6272, 821.4158, 789.7961, 
    522.9663, 274.1659, 138.3816, 105.0803, 163.4135, 285.7044, 116.0412, 
    0.01728635, 0, 0, 0, 0, 0, 0, 0, 8.116319, 2.926316, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 13.20756, 95.12429, 260.1135, 550.1265, 864.2782, 855.9658, 
    533.712, 373.4266, 157.6363, 55.62711, 19.53305, 3.260819, 19.738, 
    47.74131, 0.02607982, 0, 0, 0, 0, 0, 0, 0, 0, 7.825083, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 4.612679, 113.7198, 483.1669, 900.5347, 984.1791, 979.368, 
    648.9869, 352.2002, 216.2779, 32.69746, 0.001431095, 0, 0, 0, 3.827783, 
    4.031102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 2.923163, 13.24115, 97.76711, 368.6615, 766.6823, 981.5728, 915.0505, 
    779.8511, 465.5477, 224.4668, 57.74731, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.630818, 0, 0, 0, 
    0, 0, 0,
  0, 26.13571, 47.18822, 329.8212, 714.1318, 817.1585, 777.6345, 720.472, 
    689.508, 412.4409, 153.8221, 13.87568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14.60614, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.904786, 0, 
    0, 0, 0, 0, 0,
  75.59756, 117.36, 464.7811, 828.5286, 914.5109, 775.4006, 524.0029, 
    525.4938, 435.8335, 205.8655, 41.74298, 0, 0, 0, 0, 0, 0.005331647, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.528418, 0, 0, 0, 0, 0, 0,
  124.0725, 609.8072, 834.5482, 960.5415, 846.6204, 569.7308, 491.7551, 
    279.8958, 218.3413, 100.8299, 12.91977, 0, 0, 0, 0, 2.74017, 34.26874, 
    4.089978, 0.006493978, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  788.1714, 924.0498, 942.0076, 910.2986, 705.7488, 565.4158, 375.6508, 
    52.00785, 10.21643, 29.34002, 0, 0, 0, 0, 0, 0.3673571, 38.30904, 
    23.26111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1149.62, 1038.71, 868.4792, 750.6149, 529.3036, 359.8947, 217.0901, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.070928, 2.819205, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1133.226, 1117.429, 1080.336, 645.8721, 348.1219, 292.5666, 127.6823, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.646089, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1091.445, 1175.159, 1047.787, 521.8422, 207.5739, 209.878, 29.33293, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3.629298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1008.184, 1060.578, 851.4131, 319.3173, 106.1258, 27.16054, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.7230543, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  712.9464, 763.3522, 556.6812, 197.0247, 47.35983, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000509836, 0, 0, 8.426788, 
    29.4048, 0.002151013, 0, 0, 0, 0.2241978, 0.5720429, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.45377, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  275.8788, 288.6921, 148.9188, 9.949349, 18.65905, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.253, 138.6072, 
    10.21046, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  162.0924, 85.03082, 25.2907, 0.1707526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  134.5873, 70.08076, 39.76377, 5.510149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.902595, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  93.36883, 48.54351, 17.077, 0.7504963, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.660882e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  42.1458, 10.08691, 0.3624226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  77.45152, 3.438473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  191.3508, 37.65026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  182.4834, 62.86003, 0.8790046, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  200.0499, 98.08273, 6.234468, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  165.0487, 101.9256, 7.986403, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  53.96191, 16.12039, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  4.127634, 1.148005, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.3091331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  6.69378, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.9037046, 1, 1, 0.8371245, 0.01079098, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.342301, 1, 0.9242505, 0.2324802, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1585782, 0.8988085, 0.872375, 0.8199701, 0.2036715, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04788778, 0.3358625, 0.07239318, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1174253, 0.1658257, 0.1069185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.04039344, 0.2727596, 0.3044432, 0.03935189, 0.05927679, 
    0.5426623, 0.5088302, 0.241054, 0.0411321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04967177, 0.09058292, 0.6336873, 0.9864414, 1, 0.999317, 0.9606841, 
    0.9469818, 1, 1, 1, 0.9701587, 0.6985948, 0.1660634, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04887224, 0.4892108, 0.9759328, 0.8929602, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9605891, 0.1742972, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1475878, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2927403, 
    0.1056596, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008395956, 0.8062803, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.7915943, 0.001058526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003862719, 0.7844364, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.4460433, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3652394, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9193342, 
    0.1419819, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2822479, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9971261, 
    0.6570057, 0.2192735, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08952717, 0.2009808, 0.4916342, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.4641593, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02373972, 
    0.2887375, 0.5454076, 0.7591597, 0.9840837, 0.9225589, 0.9569725, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.2276618, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01343125, 0.2130994, 0.07166115, 
    0.1361981, 0.4062145, 0.4764926, 0.9131937, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9399245, 0.2953852, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1096427, 0.6468607, 1, 0.9679646, 
    0.8867931, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.9742239, 0.2603416, 0.000543013, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006295154, 0.4813343, 0.944672, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.811202, 0.007860967, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.3256565, 0.3595797, 0.9921021, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8934381, 0.4007365, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.5127948, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8029071, 0.1827247, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8530139, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.6570168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0181968, 0.8725816, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.7388504, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.1284515, 0.9620806, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.8478313, 0.01794271, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.05491119, 0.6775094, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.9972597, 0.1556571, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.01809847, 0.02063968, 0.5821294, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.576636, 0.0007413209, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.5811512, 0.770504, 0.5899364, 0.7125399, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9348087, 0.3177032, 0.05322447, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.7359381, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9021191, 
    0.3398403, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2397476, 0.9484219, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9444426, 0.1523203, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.7934542, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9452199, 
    0.4845907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.4458613, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.7567984, 
    0.06867129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0058354, 0.4173073, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.4904585, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0734878, 
    0.0544353, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.3889154, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.3997353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0560805, 0.6384699, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0.297665, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0808603, 0.2136603, 0.223731, 0.7629656, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.1250296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1126087, 0.07242998, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.06437702, 0.4854095, 0.7614139, 0.9957509, 0.9980491, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0.1323143, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4987842, 0.4307159, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1129699, 0.7654874, 1, 1, 1, 1, 0.9594662, 0.2817145, 
    0.349315, 0.4800343, 0.4166909, 0.33321, 0.8587425, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.5030489, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.208195, 
    0.3201258, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1805963, 0.4938805, 0.9619426, 1, 1, 0.9977201, 0.4028112, 
    0, 0, 0, 0, 0, 0.03760567, 0.4765331, 0.9889686, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6693374, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1330605, 0.07577454, 0.6408337, 1, 1, 0.8560842, 0.229482, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.7420933, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.9711934, 0.8154297, 0.7031593, 0.1591314, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2664649, 0.9408039, 1, 0.9731776, 0.3734872, 0.08581278, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2477078, 0.9847024, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.9874682, 0.6629098, 0.03976496, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.04098084, 0.6700594, 1, 0.9846117, 0.3915779, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002308619, 0.8402424, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.9393559, 0.3334898, 0.4927699, 0.1729504, 
    0.0005183411, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.05815923, 0.8921363, 0.9963881, 0.4196884, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.03001891, 0.8732678, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.8185688, 0.000997816, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3599489, 0.6536069, 0.2308225, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1388849, 0.9886107, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.8995878, 0.6226335, 0.6108878, 0.388907, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.275672, 0.4499452, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.6206766, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.6265669, 0.03419805, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004062632, 0.09197545, 0.07587977, 
    0.1429734, 0.07793289, 0.001982026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.09490187, 0.1736679, 0.3527791, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.001625569, 0.2624141, 0.8962197, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.9966809, 0.5754746, 0.03894359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2468218, 0.5043563, 0.9838024, 0.866147, 
    0.8783621, 0.9815187, 0.8271396, 0.4878259, 0.01884565, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1005597, 0.06768002, 0.1576353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.33927, 0.891219, 0.9995848, 1, 1, 0.9420939, 
    0.7670357, 0.6221464, 0.2302634, 0.2723061, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1477103, 0.6884276, 0.999054, 1, 1, 1, 0.7532653, 
    0.5085074, 0.8721771, 1, 0.3210266, 0, 0, 0, 0, 0, 0, 0, 0, 0.05677235, 
    0.0008144492, 0.04120899, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1219508, 0.1550475, 0.3309695, 0.0581816, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 2.639958e-05, 0, 0.7161255, 1, 1, 1, 1, 1, 0.7215892, 
    0.7704202, 0.9905617, 0.9987394, 0.5821542, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04867533, 0.01442351, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.04097006, 0.593925, 0.648534, 0.9974784, 1, 1, 1, 1, 
    0.999142, 0.6332727, 0.257304, 0.1315637, 0.1783369, 0.4090085, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.006319822, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.0159371, 0.6464633, 1, 1, 1, 1, 1, 1, 0.9379096, 0.3084929, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.05427543, 0.8169017, 1, 1, 1, 1, 1, 1, 1, 0.6480082, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0.0001631903, 0.2342296, 0.3217961, 1, 1, 1, 1, 1, 1, 1, 0.9198062, 
    0.2241177, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.6364967, 0.4618171, 0.704794, 1, 1, 1, 1, 1, 1, 1, 0.4258353, 0, 0, 0, 0, 
    0, 0.01590484, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.5118697, 0.9346247, 1, 1, 1, 1, 1, 0.9876335, 0.9329823, 0.9783548, 
    0.2976481, 0, 0, 0, 0, 0.01003709, 0.4619169, 0.1022752, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.9873409, 0.253808, 0.04543634, 0.5278371, 0.002404106, 
    0, 0, 0, 0, 0.003275408, 0.6632224, 0.3422698, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.7803705, 0.005725726, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03397798, 0.01880223, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 0.6511014, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 1, 1, 1, 1, 0.9937965, 0.1486441, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 1, 0.9887101, 0.3117075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 1, 0.9908476, 0.4261142, 0.01644797, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09772249, 0.07365502, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.7445699, 0.1342526, 0.4569494, 0.0158662, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01797347, 0.3693104, 
    0.01717718, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4015935, 0.05133266, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 1, 0.9750558, 0.2528034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 1, 0.6344764, 0.008912468, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.8986811, 0.1816702, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.2968034, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1, 0.8290737, 0.01273574, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.8303954, 0.01862913, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  1, 0.9919094, 0.1766838, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.9953394, 0.2376448, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  1, 0.6380026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0.6356525, 0.1226215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7992414, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2732799, 355.3445, 661.6653, 788.604, 538.0593, 35.1188, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26.84651, 302.8979, 366.1382, 
    37.41038, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39.91399, 196.7844, 215.7041, 248.1746, 36.99986, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9039114, 78.54595, 10.11436, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.704782, 26.12457, 13.85557, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005312768, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.02989985, 0.0003766294, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4189242, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1030456, 1.054963, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.143771, 12.69478, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.836948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.310095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01557077, 4.43028, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0002689204, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7.815726, 77.31487, 37.02573, 24.40091, 17.92381, 71.63206, 
    255.5557, 112.1054, 8.874227, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.931261, 18.36737, 547.9603, 983.4506, 928.882, 805.4354, 755.1304, 
    606.848, 760.251, 1122.059, 1210.754, 926.5558, 393.9966, 77.59235, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18.74462, 550.8997, 873.0414, 738.3782, 1447.062, 1752.654, 1555.512, 
    1427.795, 1463.065, 1405.852, 1591.613, 1837.372, 1954.355, 1766.622, 
    1318.124, 785.6111, 74.99232, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97.7004, 1316.783, 1765.13, 1515.387, 1988.113, 2090.078, 1944.169, 
    1852.772, 1877.534, 1980.513, 2136.833, 2321.126, 2360.485, 2221.856, 
    1762.722, 1079.052, 99.97397, 6.346212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.179383, 841.1734, 1729.189, 2051.514, 2252.923, 2277.749, 2199.887, 
    2128.035, 2119.189, 2210.886, 2389.87, 2514.411, 2530.765, 2387.412, 
    2038.683, 1570.642, 1014.397, 440.8733, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.362782, 1003.385, 1800.715, 2229.933, 2275.979, 2360.229, 2311.384, 
    2315.582, 2392.034, 2497.806, 2647.774, 2647.349, 2549.216, 2306.825, 
    2075.641, 1693.824, 991.6838, 61.70815, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    118.7808, 1369.103, 1878.122, 2249.811, 2418.137, 2469.63, 2522.086, 
    2576.791, 2679.619, 2804.705, 2853.611, 2761.156, 2575.387, 2356.625, 
    2033.336, 1327.755, 445.6916, 5.287508, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3446125, 116.4755, 1433.451, 2040.093, 2321.82, 2502.561, 2570.579, 
    2649.61, 2757.851, 2852.799, 3005.241, 3050.789, 2945.686, 2746.585, 
    2492.519, 2133.578, 1679.148, 958.2936, 281.5658, 332.4458, 79.20005, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    159.5307, 500.1543, 1869.062, 2316.033, 2462.074, 2542.433, 2621.507, 
    2731.679, 2849.691, 2997.048, 3129.562, 3153.165, 3042.124, 2822.781, 
    2579.193, 2313.826, 1938.037, 1456.275, 955.3979, 723.9649, 233.088, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    87.2196, 982.8452, 2074.387, 2401.657, 2479.505, 2552.033, 2644.845, 
    2764.61, 2913.177, 3071.668, 3188.252, 3187.021, 3067.563, 2877.698, 
    2677.985, 2453.64, 2217.535, 1895.206, 1415.486, 987.4891, 102.9291, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.006072, 9.248502, 51.24354, 
    117.7083, 0, 0, 0, 0, 0, 0, 1.781354, 493.788, 1756.028, 2232.431, 
    2436.472, 2528.297, 2640.581, 2788.757, 2970.408, 3126.261, 3223.229, 
    3201.013, 3098.396, 2951.579, 2787.688, 2644.104, 2469.223, 2265.754, 
    2020.998, 1603.012, 1036.609, 247.5821, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37.27396, 324.1435, 484.3052, 107.4387, 
    334.8317, 258.5734, 18.40336, 45.59911, 0, 0, 0, 0, 0, 312.953, 1500.18, 
    2183.505, 2342.897, 2491.774, 2647.206, 2829.54, 3007.807, 3145.192, 
    3213.799, 3194.5, 3103.396, 2991.563, 2858.539, 2725.452, 2602.863, 
    2442.798, 2299.817, 2079.573, 1678.872, 960.7639, 59.84979, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9005052, 143.1917, 891.4856, 1319.249, 
    1183.058, 743.5308, 625.7929, 271.4628, 29.0506, 28.26866, 0, 0, 0, 0, 0, 
    717.5844, 1521.244, 1982.313, 2315.337, 2501.919, 2714.457, 2879.019, 
    3038.052, 3144.582, 3199.439, 3176.925, 3090.616, 2991.669, 2897.744, 
    2785.427, 2687.85, 2575.268, 2434.927, 2202.157, 1748.342, 990.5164, 
    59.45817, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 138.0944, 28.26443, 859.6864, 1666.731, 1924.49, 
    1504.685, 894.1763, 626.5555, 183.7074, 1.250475, 6.993803, 0, 0, 0, 0, 
    152.5896, 1363.213, 1888.575, 2229.896, 2403.91, 2606.387, 2805.63, 
    2949.473, 3072.477, 3182.144, 3236.154, 3219.5, 3134.394, 3083.353, 
    3023.675, 2942.66, 2840.365, 2713.65, 2525.043, 2247.123, 1760.282, 
    1015.293, 69.54496, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 54.8675, 364.3715, 1548.06, 2161.363, 1988.979, 
    1423.904, 840.0815, 473.7389, 230.111, 231.5213, 70.41041, 0, 0, 0, 
    53.0154, 1249.682, 2001.559, 2304.354, 2429.361, 2548.836, 2707.271, 
    2894.569, 3029.046, 3159.696, 3279.65, 3330.228, 3323.386, 3284.032, 
    3259.254, 3244.029, 3164.147, 3039.184, 2858.268, 2653.644, 2425.572, 
    2034.225, 1328.45, 212.7939, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 138.5299, 947.9814, 1887.259, 2160.271, 1846.834, 
    1415.143, 971.5607, 604.7406, 412.5479, 333.2895, 159.8654, 26.29184, 
    1.857185, 274.4556, 1131.609, 1924.803, 2423.259, 2540.296, 2611.256, 
    2717.599, 2832.219, 2998.016, 3149.23, 3272.842, 3375.903, 3453.881, 
    3472.483, 3466.487, 3455.854, 3431.323, 3360.251, 3219.655, 3025.667, 
    2818.918, 2574.498, 2177.516, 1541.304, 418.2077, 3.786927, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.897408, 278.9847, 1150.151, 1820.023, 1906.937, 
    1710.571, 1470.08, 1188.798, 854.9822, 594.4963, 455.2799, 296.2944, 
    20.74247, 212.9633, 1377.01, 2210.266, 2531.037, 2589.832, 2729.739, 
    2779.357, 2870.47, 2960.67, 3105.383, 3254.163, 3365.769, 3484.833, 
    3561.692, 3602.843, 3610.362, 3592.779, 3537.574, 3466.485, 3340.572, 
    3139.534, 2890.738, 2605.906, 2178.262, 1557.431, 585.7548, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25.96501, 274.0147, 1064.936, 1482.375, 1656.331, 
    1647.515, 1562.002, 1335.74, 1001.996, 734.4821, 565.3111, 391.8153, 
    311.9492, 871.4916, 2073.987, 2854.189, 2770.159, 2864.382, 2882.136, 
    2935.086, 3016.186, 3112.14, 3232.739, 3376.769, 3504.886, 3614.249, 
    3695.932, 3704.89, 3713.67, 3686.838, 3614.497, 3529.63, 3396.464, 
    3164.898, 2869.117, 2545.209, 2079.768, 1444.332, 473.3306, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.198395, 148.0527, 886.8211, 1277.724, 1493.68, 
    1692.014, 1690.58, 1503.016, 1205.435, 994.3757, 848.381, 968.3361, 
    1305.293, 1773.208, 2657.443, 2950.178, 3028.504, 2998.262, 3013.121, 
    3056.479, 3144.256, 3246.656, 3377.553, 3516.235, 3644.559, 3743.524, 
    3749.271, 3708.808, 3678.306, 3622.363, 3548.655, 3468.685, 3334.021, 
    3096.724, 2813.21, 2507.742, 2064.155, 1345.841, 332.7528, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.602107, 0.03367292, 82.96276, 823.9019, 1207.387, 
    1490.124, 1792.475, 1887.241, 1801.419, 1641.348, 1457.016, 1489.465, 
    1791.969, 2173.656, 2577.651, 2800.211, 3040.854, 3063.57, 3082.433, 
    3086.433, 3130.878, 3234.532, 3374.836, 3510.101, 3641.93, 3775.546, 
    3826.162, 3739.047, 3612.842, 3507.702, 3436.104, 3394.341, 3313.844, 
    3186.941, 2981.263, 2736.921, 2428.213, 1957.258, 1192.974, 155.4329, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 87.60106, 73.32498, 112.404, 153.6019, 823.2629, 1290.737, 
    1591.929, 1899.596, 2085.203, 2131.1, 2032.692, 1952.935, 2003.027, 
    2256.183, 2444.568, 2635.164, 2807.364, 2928.302, 2931.476, 3038.824, 
    3101.363, 3169.576, 3315.562, 3484.013, 3647.621, 3791.786, 3922.948, 
    3926.845, 3723.422, 3456.011, 3269.509, 3160.537, 3127.081, 3060.512, 
    2938.832, 2773.188, 2564.738, 2217.429, 1614.816, 876.0974, 3.817307, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 174.1339, 192.5289, 595.6072, 548.1959, 902.9622, 
    1324.524, 1637.417, 1968.1, 2162.593, 2136.62, 2034.022, 1937.629, 
    2005.565, 1973.358, 2069.837, 2373.308, 2690.74, 2792.308, 2870.053, 
    3000.035, 3104.013, 3210.098, 3377.595, 3564.663, 3770.401, 3917.039, 
    4012.642, 3948.944, 3671.559, 3324.181, 3003.464, 2810.002, 2744.527, 
    2678.826, 2554.504, 2450.903, 2248.528, 1666.047, 879.4138, 217.8605, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41.24575, 171.1755, 928.2092, 911.556, 1003.465, 1333.517, 
    1742.872, 1976.593, 1971.419, 1847.775, 1596.083, 1517.469, 1510.441, 
    1449.914, 1648.969, 2160.01, 2465.792, 2611.214, 2691.124, 2869.434, 
    3045.968, 3236.557, 3398.76, 3579.36, 3797.204, 3936.64, 3975.402, 
    3863.231, 3599.677, 3223.608, 2813.848, 2505.323, 2321.725, 2250.189, 
    2064.987, 1902.286, 1638.834, 1019.027, 91.78241, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 105.7556, 967.28, 1137.105, 1125.491, 1369.858, 
    1526.296, 1610.441, 1462.915, 1195.448, 979.7076, 964.7514, 1033.812, 
    1020.986, 1503.457, 1979.614, 2248.812, 2429.502, 2603.554, 2766.973, 
    2963.375, 3182.582, 3375.808, 3529.749, 3729.817, 3856.099, 3884.153, 
    3740.839, 3498.397, 3131.312, 2677.872, 2252.273, 1934.652, 1693.907, 
    1330.782, 934.9443, 600.6172, 199.5566, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.739202, 0, 0, 0, 56.65801, 764.7597, 1177.214, 1137.807, 
    867.6033, 751.4905, 455.4625, 373.3823, 389.2663, 356.8941, 412.8959, 
    422.8545, 839.1047, 1290.905, 1814.671, 2116.265, 2387.323, 2578.228, 
    2692.938, 2810.998, 3018.81, 3251.787, 3454.09, 3636.555, 3767.025, 
    3772.435, 3602.902, 3361.617, 3049.529, 2649.456, 2152.187, 1589.401, 
    1095.306, 616.2491, 204.8285, 109.602, 22.18781, 48.89778, 9.825142, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009279916, 251.9048, 962.301, 883.4589, 677.3438, 
    361.7939, 137.7333, 20.846, 41.77541, 29.66083, 35.41616, 248.8549, 
    735.1519, 1335.172, 1731.033, 2074.124, 2359.61, 2570.465, 2604.922, 
    2667.29, 2813.544, 3063.244, 3317.592, 3564.776, 3708.774, 3713.399, 
    3546.005, 3335.875, 3064.894, 2726.397, 2302.653, 1790.918, 1349.976, 
    1108.172, 1070.336, 1060.536, 925.6852, 754.9511, 214.2521, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23.60169, 0.001468251, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 112.4058, 711.1246, 782.2984, 371.9018, 202.2023, 
    4.081332, 19.38192, 1.332851, 0.4524727, 2.236566, 63.69951, 569.4813, 
    1187.416, 1604.718, 1946.94, 2248.886, 2439.147, 2533.595, 2566.406, 
    2670.604, 2904.311, 3214.155, 3497.722, 3662.987, 3690.172, 3581.76, 
    3430.937, 3210.368, 2925.982, 2596.184, 2305.98, 2085.327, 1988.169, 
    1999.194, 2000.523, 1668.639, 1237.938, 193.779, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0277722, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.159892, 56.1418, 452.5438, 1005.819, 940.8052, 
    359.2229, 45.87414, 0.6317925, -4.440892e-16, 0.4750352, 33.37933, 
    3.9842, 295.6864, 921.4279, 1533.577, 1758.771, 2015.291, 2243.664, 
    2363.067, 2499.792, 2603.064, 2851.553, 3174.852, 3439.871, 3601.986, 
    3639.036, 3611.236, 3520.832, 3376.327, 3171.316, 2925.103, 2754.788, 
    2670.149, 2638.344, 2562.51, 2441.751, 2061.093, 1274.259, 129.2553, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 40.98916, 47.87557, 244.1692, 1334.147, 1438.746, 
    508.3959, 23.03855, -1.734723e-18, 0, 10.75564, 254.7662, 148.7082, 
    109.2365, 659.3992, 1310.688, 1593.068, 1868.237, 2051.256, 2239.637, 
    2436.269, 2622.957, 2896.737, 3180.859, 3412.578, 3564.607, 3677.027, 
    3686.917, 3618.097, 3508.476, 3355.026, 3184.518, 3051.357, 3012.698, 
    2935.528, 2832.188, 2615.409, 2041.958, 1159, 32.8907, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.57209, 3.683461, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13.15392, 21.53556, 145.4484, 166.8116, 212.421, 1456.922, 
    1442.133, 274.9966, 0, 0, 0.3660825, 97.71632, 274.119, 216.5157, 
    1.421085e-14, 355.3852, 921.0424, 1435.383, 1760.988, 2009.327, 2226.052, 
    2488.684, 2725.142, 2982.086, 3207.749, 3389.718, 3565.573, 3709.347, 
    3742.948, 3657.837, 3548.883, 3403.997, 3227.927, 3100.738, 3010.48, 
    2897.043, 2753.1, 2530.298, 1963.905, 996.7645, 20.1157, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 95.68005, 62.03844, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 76.78776, 251.8225, 365.1784, 499.3779, 679.7224, 1282.687, 
    976.8096, 54.30797, 0, 0, -4.440892e-16, 3.06115, 105.1266, 7.105427e-15, 
    146.4528, 166.1453, 740.5073, 1156.732, 1667.2, 2071.25, 2311.511, 
    2561.432, 2802.865, 3051.193, 3239.81, 3403.32, 3577.332, 3697.356, 
    3695.489, 3575.418, 3467.606, 3301.877, 3080.048, 2891.024, 2773.609, 
    2640.24, 2458.685, 2296.196, 1776.581, 1080.293, 215.078, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20.15371, 42.59801, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 132.3908, 427.5094, 871.1767, 1216.166, 1215.606, 1074.381, 
    143.933, 0, 0, 0, 0, 4.440892e-16, 0.7024416, 85.66618, 422.4643, 
    753.0161, 876.0609, 1329.78, 1707.256, 2086.016, 2393.784, 2545.285, 
    2840.856, 3071.359, 3268.794, 3422.524, 3586.531, 3666.174, 3565.691, 
    3397.146, 3270.382, 3125.957, 2841.437, 2580.784, 2474.215, 2351.78, 
    2078.684, 1727.895, 1498.923, 1140.002, 539.2833, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 62.32169, 39.41545, 626.6343, 1371.758, 1347.847, 687.8185, 
    32.66976, 0, 0, 0, 0, 0, 0, -6.938894e-18, 29.09192, 611.8069, 1072.647, 
    1446.324, 1597.489, 1872.625, 2189.95, 2396.317, 2632.638, 2864.967, 
    3116.256, 3290.928, 3442.491, 3576.208, 3595.495, 3416.291, 3130.265, 
    2946.176, 2774.498, 2500.969, 2090.21, 2070.135, 2101.286, 1651.494, 
    934.1992, 472.3446, 447.5172, 68.89008, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 239.6809, 554.4179, 364.8323, 498.6555, 95.83427, 6.607563, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 132.7997, 1047.2, 1417.112, 1781.415, 2066.203, 
    2268.176, 2513.788, 2702.935, 2989.756, 3186.11, 3356.546, 3463.798, 
    3540.333, 3487.458, 3305.011, 2838.596, 2431.235, 2225.709, 1948.767, 
    1463.512, 1303.707, 1487.188, 1115.347, 344.4456, 17.17711, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.06872149, 590.6149, 255.9139, 0.4632595, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 187.6016, 678.9084, 1330.984, 2035.844, 2433.294, 
    2612.385, 2832.168, 3016.011, 3219.117, 3378.409, 3442.958, 3400.81, 
    3281.248, 3011.857, 2341.452, 1747.214, 1505.163, 1297.308, 751.0115, 
    196.1539, 377.1983, 100.9759, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 38.59026, 645.7719, 34.58854, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53.31918, 810.9399, 1739.455, 2404.192, 2757.1, 2846.992, 
    2957.257, 3148.64, 3318.68, 3306.222, 3091.919, 2659.991, 2079.938, 
    1357.805, 792.2961, 628.3082, 498.0571, 246.4902, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 235.8719, 404.9598, 19.19321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1208589, 268.1322, 1044.283, 1926.036, 2449.009, 2629.04, 
    2630.753, 3113.425, 3114.51, 2984.559, 2508.903, 1782.817, 1010.823, 
    372.2121, 24.88615, 0.03625189, 0.009416752, 86.38479, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14.21238, 250.7785, 295.3082, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 155.7787, 592.4962, 1366.038, 1963.625, 1825.582, 2069.24, 
    2485.683, 2492.135, 2126.706, 1540.313, 896.8804, 239.871, 46.3145, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.80038, 14.7334, 38.18274, 15.65409, 
    2.098015, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.28813, 129.1734, 304.9514, 
    3.314995, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 149.1334, 
    773.5136, 1044.637, 889.3293, 853.0041, 1272.865, 1052.722, 795.8773, 
    379.6655, 140.3403, 5.892643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.09859627, 30.3471, 81.51091, 108.4727, 153.5919, 
    206.7384, 204.1187, 155.7402, 96.83952, 3.76339, 0, 0, 0, 0, 0, 0, 0, 0, 
    19.27378, 11.65506, 100.7927, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 26.58224, 97.38688, 141.9256, 27.09244, 26.51507, 114.4799, 
    79.36494, 31.06278, 0, 0.04206881, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 26.76524, 161.1405, 374.7367, 504.8459, 444.2382, 
    263.0925, 173.7267, 155.3289, 255.5945, 377.7833, 81.20056, 2.50277, 0, 
    0, 0, 0, 0, 0, 0, 19.48863, 0, 17.85832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 17.59249, 7.557294, 179.5778, 668.6272, 821.4158, 789.7961, 
    522.9663, 274.1659, 138.3816, 105.0803, 163.4135, 285.7044, 116.0412, 
    0.01728635, 0, 0, 0, 0, 0, 0, 0, 8.116319, 2.926316, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 13.20756, 95.12429, 260.1135, 550.1265, 864.2782, 855.9658, 
    533.712, 373.4266, 157.6363, 55.62711, 19.53305, 3.260819, 19.738, 
    47.74131, 0.02607982, 0, 0, 0, 0, 0, 0, 0, 0, 7.825083, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 4.612679, 113.7198, 483.1669, 900.5347, 984.1791, 979.368, 
    648.9869, 352.2002, 216.2779, 32.69746, 0.001431095, 0, 0, 0, 3.827783, 
    4.031102, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 2.923163, 13.24115, 97.76711, 368.6615, 766.6823, 981.5728, 915.0505, 
    779.8511, 465.5477, 224.4668, 57.74731, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.630818, 0, 0, 0, 
    0, 0, 0,
  0, 26.13571, 47.18822, 329.8212, 714.1318, 817.1585, 777.6345, 720.472, 
    689.508, 412.4409, 153.8221, 13.87568, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 14.60614, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.904786, 0, 
    0, 0, 0, 0, 0,
  75.59756, 117.36, 464.7811, 828.5286, 914.5109, 775.4006, 524.0029, 
    525.4938, 435.8335, 205.8655, 41.74298, 0, 0, 0, 0, 0, 0.005331647, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.528418, 0, 0, 0, 0, 0, 0,
  124.0725, 609.8072, 834.5482, 960.5415, 846.6204, 569.7308, 491.7551, 
    279.8958, 218.3413, 100.8299, 12.91977, 0, 0, 0, 0, 2.74017, 34.26874, 
    4.089978, 0.006493978, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  788.1714, 924.0498, 942.0076, 910.2986, 705.7488, 565.4158, 375.6508, 
    52.00785, 10.21643, 29.34002, 0, 0, 0, 0, 0, 0.3673571, 38.30904, 
    23.26111, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  1149.62, 1038.71, 868.4792, 750.6149, 529.3036, 359.8947, 217.0901, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.070928, 2.819205, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1133.226, 1117.429, 1080.336, 645.8721, 348.1219, 292.5666, 127.6823, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.646089, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1091.445, 1175.159, 1047.787, 521.8422, 207.5739, 209.878, 29.33293, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3.629298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1008.184, 1060.578, 851.4131, 319.3173, 106.1258, 27.16054, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.7230543, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  712.9464, 763.3522, 556.6812, 197.0247, 47.35983, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000509836, 0, 0, 8.426788, 
    29.4048, 0.002151013, 0, 0, 0, 0.2241978, 0.5720429, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.45377, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  275.8788, 288.6921, 148.9188, 9.949349, 18.65905, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14.253, 138.6072, 
    10.21046, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  162.0924, 85.03082, 25.2907, 0.1707526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  134.5873, 70.08076, 39.76377, 5.510149, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.902595, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  93.36883, 48.54351, 17.077, 0.7504963, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.660882e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  42.1458, 10.08691, 0.3624226, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  77.45152, 3.438473, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  191.3508, 37.65026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  182.4834, 62.86003, 0.8790046, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  200.0499, 98.08273, 6.234468, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  165.0487, 101.9256, 7.986403, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  53.96191, 16.12039, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  4.127634, 1.148005, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0.3091331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  6.69378, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
