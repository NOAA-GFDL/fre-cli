netcdf atmos.1980-1981.aliq.11 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:23 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.11.nc reduced/atmos.1980-1981.aliq.11.nc\n",
			"Mon Aug 25 14:40:56 2025: cdo -O -s -select,month=11 merged_output.nc monthly_nc_files/all_years.11.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.477351e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004125764, 0.0001220227, 0.0002077731, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 2.133283e-07, -2.790244e-05, 0, -3.135588e-06, 0, 0, 0, 0, 0, 0, 0, 
    -5.876928e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000160211, 0, 0, 0,
  0, -6.986973e-06, -5.698249e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -1.045017e-05, -1.086787e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.0003880856, -2.663957e-05, 0.0007909854, 
    0.0004360115, 0.00018059, 0.0003995473, 0, 1.328684e-05, 0, 0, 
    -6.018905e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.983225e-05, -4.000842e-07, -1.793312e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.955553e-05, 0, 0, 0,
  0, 0, -3.943291e-06, -7.270707e-05, 0.0001046347, -1.887175e-05, 0, 0, 0, 
    0, 0, 0, 0, -9.900304e-05, -6.882213e-06, 0.001967175, 0, 0, 0, 0, 0, 0, 
    0, 0, -2.144113e-05, 0.001086961, 0, 0, 0,
  0, 0.000504988, -5.930079e-06, 0, -5.309697e-06, 0, 0, 0, 2.919231e-06, 0, 
    0, 0, 0, -9.836776e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003591845, 
    -1.828804e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.001081229, -8.113584e-05, 0.002275015, 0.001246437, 
    0.0005141768, 0.001243126, 0.001150693, 6.944773e-06, 0, 0.0008218914, 
    -2.285294e-05, 0, -2.792115e-05, -4.122836e-05, 0, 0, -3.063232e-06, 0, 
    -4.269799e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.32758e-06, -2.327206e-06, -9.723382e-07, 
    -4.626169e-05, 7.441124e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0.0003200208, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.230005e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, -3.13166e-05, 0, 0, 0,
  0, 0, 0.0002745432, -2.203883e-05, 0.0003511936, 2.503707e-05, 0.001311897, 
    -2.064802e-05, 0, 0, 0, 0, 0, 0.000231019, 0.001728961, 0.002582901, 0, 
    0, 0, 0, 0, 0, 0, -4.004056e-06, -4.758954e-05, 0.002813295, 0, 0, 0,
  0, 0.001181712, -1.004493e-05, 0, -3.604913e-05, 0.000606424, 0, 0, 
    -2.339874e-05, -2.804195e-05, 0, 0, 0, 5.125105e-05, 0, -6.117293e-07, 0, 
    0, 0, 0, 0, 0, 0, 0.0003907428, -3.444554e-05, 0, 0.0001556521, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.004014635, -0.0001695841, 0.004724398, 0.003190717, 
    0.001470751, 0.00298365, 0.003462777, 0.0002495023, -3.686141e-06, 
    0.003140341, 0.0006952575, 0.0005981278, -9.317166e-05, 0.00251773, 0, 0, 
    -3.227113e-05, 0, 0.0002360819, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.994822e-05, 0.002150742, -1.077876e-06, 
    -0.0001188753, 0.002713965, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004455626, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.593581e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -4.873743e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0004671463, -1.036831e-05, -1.516479e-05, 0, 0,
  0, 0, 0.001516126, 0, -7.130448e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.697364e-05, -1.494886e-05, 0, 0, 0, 0, 0, 0, 0, -9.631022e-05, 
    0.0004869055, 0, 0,
  0, -1.745142e-05, 0.001038432, 0.001337317, 0.001297986, 0.002931188, 
    0.002551123, 0.0001133972, -7.745618e-06, 0, 0, -2.274146e-05, 0, 
    0.005131501, 0.004419999, 0.003362385, 0.0006224072, 0, 0, 0, 0, 0, 0, 
    7.114512e-05, -8.374075e-05, 0.00420707, 0, 0, 0,
  0, 0.002462932, 0.0003772919, 0, -7.624932e-05, 0.0009660443, 0, 0, 
    0.0001171861, -7.488056e-05, -1.490287e-05, -1.209894e-05, -1.202274e-06, 
    0.000469847, 0, 1.333847e-05, -1.073856e-05, 0, 0, 0, 0, 0, 0, 
    0.0003904286, -2.753084e-05, 0, 0.001243333, 0, 0,
  0, 0, 0, 0, 0, -3.187805e-06, 0, 0.009049562, -6.999614e-05, 0.01009295, 
    0.005153945, 0.002634415, 0.007595866, 0.006279867, 0.0006324413, 
    -9.453547e-06, 0.005347097, 0.002350325, 0.00223577, 0.0006247329, 
    0.01095329, -5.388135e-06, -4.139106e-05, -6.464512e-05, -1.586336e-05, 
    0.0003055907, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.000109378, -4.658612e-05, 0.008589149, 
    -4.704762e-05, 0.0003007344, 0.007755606, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004946164, 0.00641626, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -9.094725e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -2.424584e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.236681e-05, -6.354287e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.432863e-05, 0, 0, 0, 0, 0, 0, 0, 0, -6.691657e-07, 0, 0, 0, 
    0, 0.0002888344, 0, 0, 0, 0, 0, 0.0009273991, -7.410922e-07, 0, 0, 0,
  0, 0, 0, 4.112464e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.868107e-06, 0, 0, 
    -1.57437e-05, 0, -9.838264e-06, -4.80627e-06, 0, 0, 0, 0, 0.001048995, 
    0.000450581, 0.0001563275, 0, 0,
  0, 0, 0.002395728, 0.0002975923, -1.556965e-05, 0.0007390097, 0, 0, 0, 0, 
    0, 0, 0, 5.41995e-05, -5.594662e-06, 0.0006552096, 0.002381678, 
    0.0001136452, -1.75048e-05, 0, 0, 0, 0, 0, 7.353174e-05, -5.697366e-05, 
    0.00180935, 0, 0,
  0, -4.899598e-05, 0.001370668, 0.002465692, 0.002120931, 0.005038876, 
    0.004965415, 0.0005635393, -3.49211e-05, 0, 0, -4.316232e-05, 
    -3.389539e-05, 0.009337727, 0.007292184, 0.005425583, 0.003323818, 0, 0, 
    0, 0, 0, 0, 1.07275e-05, 0.0004004702, 0.00507328, 0, 0, 0,
  -2.537373e-06, 0.004184441, 0.002876065, 0, 0.0003202703, 0.001005957, 
    -4.030988e-06, 0, 0.006087746, -0.0001145157, -0.0001111752, -2.654e-05, 
    -8.906187e-06, 0.001187145, -2.451168e-06, 3.908518e-05, -4.767404e-05, 
    0, 0, 0, 0, 0, 0, 0.0003939636, 2.854815e-05, 0.0002439318, 0.002958971, 
    0, 0,
  0, 0, 0, 0, -7.936641e-07, -1.303779e-05, -3.121918e-05, 0.01572987, 
    0.003476398, 0.02050146, 0.009261896, 0.004906115, 0.01221337, 
    0.01492883, 0.002460585, 0.0003969151, 0.009339701, 0.01051425, 
    0.004352438, 0.001330144, 0.02153202, -0.0001012431, -8.180452e-05, 
    -7.80923e-05, -5.228081e-05, 0.001505001, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0001261044, -8.113834e-05, 0.01803552, 
    -0.0001068998, 0.001254336, 0.01648497, 0, 0, 0, 0, 0, 0, 0.0002863174, 
    0.0001088715, 0.002517245, 0.0074139, -8.802403e-06, 0.0005233938, 0, 0, 0,
  0, 0, 0, 0, -5.063834e-05, 0, 0, 0, 0, 0, 0, 0, -2.676287e-05, 
    -7.756474e-06, 0.0006201902, -1.253525e-05, 0, 0, 0, 0, 0, 0, 
    0.0005696531, -1.358377e-06, 0, 0.001006961, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000240067, 0, -5.244455e-06, 
    0.000445804, 0.001218446, 0, 0, 0, 0, 0, 0, 0.0004225352, -3.55253e-05, 
    1.444347e-05, -1.553482e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000195677, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004048589, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, -1.230647e-05, 2.678423e-05, -6.930444e-06, 0, 0, 0, 0, 0, 0, 0, 
    -1.762436e-05, 0, 0, 0, 0, 0.001752747, 0, 0, 0, 0, 0, 0.002355175, 
    0.001462034, -4.057874e-05, 0, 0,
  0, 0, -2.029617e-06, 0.0008505313, 1.876858e-05, 0, 0, 0, 0, 0, 0, 
    0.0003081867, 0, -9.772799e-05, 0, 0, 0.002829224, 0.0006820983, 
    0.0005129733, -5.276488e-05, -5.570498e-07, 0, 0, 0, 0.002678894, 
    0.002348858, 0.0007018151, 0, 0,
  0, 0, 0.00337042, 0.0007442307, -5.391715e-05, 0.002767946, 0, 0, 0, 0, 0, 
    0, 0, 0.001219061, -2.96172e-05, 0.001205075, 0.005141148, 0.0001423465, 
    0.0001319875, 0, 0, 0, 0, -4.643726e-08, 0.0006427958, 0.001612782, 
    0.003450837, 0, 0,
  0, -0.0001148498, 0.001649596, 0.004193448, 0.004115804, 0.006825165, 
    0.008434437, 0.00208797, 0.0003598997, 0, 0, -7.829331e-05, 
    -0.0001611206, 0.01580672, 0.01123743, 0.008486304, 0.006748339, 0, 0, 0, 
    0, 0, 0, 5.117965e-05, 0.001244955, 0.005998129, 0.001967682, 0, 0,
  -6.013729e-05, 0.007008546, 0.005524156, 0, 0.001235794, 0.002282878, 
    -4.030988e-06, -4.903346e-06, 0.01378163, 0.0008898253, 3.68383e-05, 
    -6.815032e-05, 0.00181714, 0.0057132, -1.227016e-05, 9.899977e-06, 
    -0.0001418853, 0, -1.075792e-05, 0, 0, 0, 0, 0.004226848, 6.428984e-05, 
    0.001179283, 0.004931308, 0, 0,
  0, 0, 0, 0, 6.828045e-06, 1.97129e-05, -6.002247e-05, 0.02390185, 
    0.01136036, 0.03285182, 0.01894946, 0.01272062, 0.02140753, 0.03140511, 
    0.005500703, 0.001732347, 0.01706045, 0.01998507, 0.005827788, 
    0.003369878, 0.03651967, -0.0002122247, -0.0003096875, 0.0002178839, 
    0.0001429274, 0.003509085, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 1.509204e-05, 0.001132872, 4.170081e-05, 0.03098722, 
    0.0002493937, 0.003244847, 0.03039163, -2.428139e-05, 0, -1.687678e-05, 
    -1.287775e-05, -3.127331e-06, 0, 0.0004791944, 0.001762783, 0.003850843, 
    0.009204227, 4.817305e-06, 0.003157841, 0, 0, 0,
  0, 0, 0, 0, -4.631731e-05, 0, 0, 0, 0, 0, 0, 0, 0.002266586, 0.001059432, 
    0.002869412, 6.681136e-05, 0, 0, 0, 0, 0, 9.005817e-06, 0.002103495, 
    0.000997716, 0.0006184727, 0.00300972, 0, 0, 0,
  0, 0, 0, 0, -1.146806e-05, 0, 0, 0, 0, 0, 0, 0, -1.468191e-05, 0.001661214, 
    -1.519745e-05, 0.001141524, 0.00123827, 0.004389889, 0, 0, 0, 0, 0, 
    -2.026092e-06, 0.002081159, 0.0003608517, 0.001924255, -3.766322e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004400677, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.867018e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0.001791267, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, -1.460918e-05, -8.916952e-06, 0, 0,
  -2.092594e-07, 0, 0, 0.001273299, 0.001806439, 0.0005535411, 0, 0, 0, 0, 0, 
    -8.333863e-08, -8.22365e-06, 0.001624995, 4.874559e-05, 0, 0, 0, 
    0.002432482, -8.03036e-05, 0, 0, 0, 0, 0.00544023, 0.008811524, 
    0.001728278, 0, -5.385761e-06,
  0, 0, 3.840539e-05, 0.006784768, 0.002208099, -4.63254e-05, 0, 0, 0, 0, 0, 
    0.002262071, -7.946885e-06, 0.002259508, 0, -1.658218e-06, 0.008478372, 
    0.005647837, 0.007308967, -9.317845e-05, 0.0002938031, 0, 0, 0, 
    0.006925656, 0.008600023, 0.002097765, -1.674487e-05, 0,
  0, 0.0001156039, 0.007814094, 0.001363918, -9.113066e-05, 0.00506007, 
    -5.537489e-05, 0.0007398846, 0, 0, -2.879259e-06, -1.780021e-08, 0, 
    0.003087872, -0.0001542438, 0.00406194, 0.008980745, 0.003929342, 
    0.002310989, 0, 0, 0, 0, -8.398717e-07, 0.003048202, 0.004547142, 
    0.006808838, 0, 0,
  0, 0.0004797601, 0.002500763, 0.008541073, 0.01601351, 0.01715452, 
    0.01522249, 0.006905605, 0.002163098, -4.267688e-06, -6.321066e-10, 
    0.0001522749, 0.001032133, 0.02578574, 0.01774425, 0.01598591, 0.0153484, 
    0, 0, 0, 0, 0, 0, 0.001445064, 0.005986538, 0.009137388, 0.004499671, 0, 0,
  3.915761e-05, 0.01334399, 0.01537121, -8.266292e-06, 0.002357649, 
    0.004956239, -1.35187e-05, -2.851793e-05, 0.02718825, 0.003093038, 
    0.0008371481, -0.0002412922, 0.003006778, 0.01948612, 0.000671806, 
    0.002603787, 0.0002543737, -9.813846e-07, 1.024341e-05, 0, 0, 0, 
    -1.22592e-08, 0.008446775, 0.001649352, 0.002887106, 0.01138494, 
    -6.230671e-06, 0,
  0, 0, 3.511051e-05, 0, -1.65319e-05, 0.0004816196, -0.0001790848, 
    0.02941906, 0.01941605, 0.04953501, 0.03624672, 0.02620699, 0.03951008, 
    0.05189727, 0.01154376, 0.005007359, 0.03054061, 0.03435552, 0.00987619, 
    0.008707414, 0.06507914, -0.0003283766, 0.000549556, 0.002230686, 
    0.0005491596, 0.008366155, 0.0002883508, 0, 0,
  0, 0, 0, 0, 0, -1.130842e-06, 0, 0.0013457, 0.002560136, 0.002257941, 
    0.04506641, 0.003498377, 0.009025826, 0.0393202, -2.709675e-05, 0, 
    0.0001524563, -1.929008e-05, -1.250932e-05, 0, 0.001724557, 0.0036091, 
    0.0063367, 0.01688083, 6.97625e-06, 0.005076066, 0, 0, 0,
  0, 0, 0, 0.001308808, 0.0004996121, 0, 0, 0, -7.224586e-08, 0, 
    -3.748968e-06, -4.375389e-05, 0.003657336, 0.002831189, 0.005915017, 
    0.001579794, 0, 0, 0, 0, 0, 0.002020941, 0.003847953, 0.002987432, 
    0.002044396, 0.007391315, -1.710713e-05, 0, 0,
  0, 0, 0, 0, 0.0001329038, 0, 0, 0, 0, 0, 0, 1.510949e-09, 0.001033053, 
    0.004280454, 0.0002793568, 0.006431458, 0.003264181, 0.006399704, 
    -2.917744e-08, -1.556995e-05, 0, 0, 0.0001751746, 0.002654744, 
    0.007430259, 0.001667044, 0.002833065, -9.27119e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002278431, 0, 0, 0, -1.506004e-05, 
    -3.476864e-05, 0, 0, 0, 0, 0, 0.0007914159, -4.968683e-05, 0.00156927, 
    -3.640386e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.227345e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -6.717799e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.806564e-06, 
    0, 0, 0, 0, 0, 0, 0.0008954047, 0,
  -9.376837e-06, -1.519174e-06, 0, 0, -4.343024e-05, 0.0002473389, 
    0.0001049113, -4.475553e-06, 0, 0, 0, 0, 0, -1.120965e-05, 0.002155864, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001893331, -1.120957e-05, -1.653441e-06, 
    -3.245294e-06,
  0.0004266569, -1.308905e-05, 0, 0.006165482, 0.009724301, 0.006353055, 
    0.001134011, -8.74227e-06, 0, 0, -2.391447e-06, -5.479804e-05, 
    0.0004617036, 0.006641957, 0.0004421158, -4.515589e-06, -5.862138e-07, 
    0.001888093, 0.00530354, 0.001645858, 2.355691e-05, 0.001284021, 0, 0, 
    0.009638148, 0.019984, 0.007044812, -2.912896e-06, 0.000774572,
  -9.189308e-07, 0, 0.0008541866, 0.02056008, 0.005890124, 0.001588945, 
    1.67356e-05, 0, 6.453297e-05, 4.595551e-06, 5.776785e-06, 0.003577319, 
    1.678231e-05, 0.008221057, -3.8677e-05, -3.226438e-05, 0.01545244, 
    0.01479235, 0.02829047, -0.0002639732, 0.0005146668, 0, 0, 0, 0.01879479, 
    0.0178772, 0.008599302, 0.0007851913, 0,
  0, 0.000312858, 0.01090161, 0.004181319, -0.0001041513, 0.009074887, 
    0.000833623, 0.001366976, 0, 4.937311e-07, -2.676405e-05, -4.704075e-06, 
    7.153638e-08, 0.008525055, 0.0002205179, 0.009501483, 0.01869337, 
    0.01354873, 0.007515265, -2.222219e-06, -4.777598e-07, 0, 0, 
    -3.599975e-05, 0.008738667, 0.0150323, 0.01497688, 2.351363e-05, 0,
  0, 0.002801489, 0.008570719, 0.02338148, 0.03205356, 0.03945876, 
    0.03173136, 0.01458305, 0.005192414, 2.569064e-05, 0.000469512, 
    0.002620277, 0.01036754, 0.06312788, 0.03556569, 0.03232877, 0.02613014, 
    -1.31683e-10, 0, 0, 0, 0, 0, 0.01694212, 0.04637478, 0.01972925, 
    0.006380854, -1.254545e-09, 0,
  0.005823598, 0.02399264, 0.04217618, 0.0001568015, 0.0160207, 0.01604182, 
    0.00153513, 0.0001676067, 0.05150342, 0.01215326, 0.01184472, 
    0.004194974, 0.01585532, 0.05079409, 0.001719136, 0.005161857, 
    0.001403498, -3.393686e-05, 0.0007087258, 0.00134436, -7.782212e-05, 
    3.754681e-09, 6.147573e-06, 0.02970159, 0.02050443, 0.004996873, 
    0.0180375, -6.699934e-06, 9.248982e-10,
  0, 3.47295e-07, 0.0001016657, -7.080019e-09, 0.001888586, 0.0007055108, 
    0.0002465713, 0.03882707, 0.02972602, 0.06876324, 0.05462411, 0.04841963, 
    0.08212633, 0.09009221, 0.02759699, 0.01334896, 0.04983095, 0.05514219, 
    0.02022299, 0.02032844, 0.09334358, 0.002431408, 0.01948021, 0.009101802, 
    0.004758341, 0.01471261, 0.002339773, -8.017597e-07, 2.057134e-07,
  0, 0, 0, 5.294922e-08, 0, -3.102897e-05, -3.721132e-05, 0.009097881, 
    0.007232971, 0.006475901, 0.06411575, 0.01226395, 0.01581149, 0.04823498, 
    0.001326722, 0.000315781, 0.0006528943, 0.002560876, 0.000526401, 
    -3.065649e-05, 0.006040166, 0.008894907, 0.008487659, 0.02229089, 
    0.0008429189, 0.01010909, 0.0004196698, 0.0002941838, -5.044771e-05,
  0, 0, 0, 0.004127591, 0.002673443, 1.209943e-05, 0, 0, -1.543469e-05, 
    1.711948e-05, -5.368473e-07, -3.554701e-06, 0.005888891, 0.01060233, 
    0.01179099, 0.007612505, 0.0007496625, 2.273771e-05, 5.934473e-06, 0, 
    -1.633201e-05, 0.01132295, 0.01076492, 0.004829364, 0.006303975, 
    0.0168708, -6.777008e-05, -3.117685e-05, -1.921976e-05,
  0, 0, 0, 2.902174e-05, 0.0003289914, 0, 0, 0, 0, 0, 0, 2.781635e-05, 
    0.003079541, 0.0121718, 0.006313776, 0.01485773, 0.008326847, 0.01145746, 
    0.001009202, 0.0001647281, 0, 0, 0.0001685926, 0.007995575, 0.01816829, 
    0.00510408, 0.007207152, 0.000125759, 5.507865e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.34044e-05, 0.004040684, 0.001057412, 
    1.00606e-05, 0, 0.0004521555, 0.001604904, -1.061772e-05, -7.740157e-06, 
    0, 0, 0, 0.00629694, 0.0001299825, 0.00368468, 1.561761e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.491515e-07, 0, 0, 0, 0, 
    -3.054579e-06, 0, 0, 0, 0, 0.0005397886, 0.002802128, 0.001219945, 
    -6.423506e-06, 1.586813e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.753837e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.484081e-07, 0, 0, 0, 0, 
    0.0005765828, 0, -9.840624e-06, 0, 0, 0, 0, 0.001340917, -6.238783e-06,
  0.001870104, 7.203154e-05, -3.290702e-06, -3.31265e-05, 0.00162106, 
    0.001221374, 0.002772423, 0.002028716, -1.337344e-07, -1.981924e-05, 
    -4.564636e-06, -2.775392e-06, -3.635882e-06, 0.001340023, 0.00319997, 
    0.0002824032, 5.682399e-05, 0, -7.819501e-06, -9.365313e-05, 
    -4.35774e-06, 0, 0.000671284, -3.15568e-09, -2.636131e-06, 0.002862602, 
    0.002739625, 0.002809773, 0.0008646392,
  0.001429032, 0.000102478, 2.772842e-05, 0.01707794, 0.02383697, 0.01508781, 
    0.004973792, 0.0007759312, -8.492404e-06, -3.014176e-05, 4.600523e-06, 
    0.000295558, 0.00168904, 0.01972902, 0.004745156, 0.002264338, 
    -3.356483e-05, 0.005931552, 0.01534554, 0.008658933, 0.00333451, 
    0.00592449, -3.536375e-05, -2.993494e-05, 0.01665925, 0.03513266, 
    0.02173118, 0.0007431306, 0.006121492,
  -1.189296e-05, 0.0002192449, 0.002872763, 0.0414615, 0.01467746, 
    0.009509637, 0.0001194786, 0.002385502, 0.001486001, 5.167018e-05, 
    -1.706263e-05, 0.005922901, 0.0003396698, 0.01176016, 0.00183743, 
    0.006268308, 0.02211409, 0.02507001, 0.06015055, 0.00286248, 0.003029915, 
    0, -2.706853e-10, 8.05257e-08, 0.02869587, 0.02921458, 0.02263099, 
    0.00272287, 1.161e-05,
  3.106197e-08, 0.001641297, 0.03529473, 0.01140322, 0.00174866, 0.01291739, 
    0.005395774, 0.002887632, 9.864594e-07, 7.749152e-05, 0.0009513408, 
    -2.417132e-05, 4.671795e-05, 0.01927387, 0.006532091, 0.01905655, 
    0.03459336, 0.03586431, 0.01859245, 0.0004090248, 0.0003544353, 
    8.384545e-06, 0, 0.01288344, 0.07631589, 0.02929925, 0.03055245, 
    0.00019083, -3.583044e-06,
  -5.529226e-06, 0.09186114, 0.03466508, 0.04250204, 0.05385505, 0.06201155, 
    0.06721924, 0.05534011, 0.01158171, 0.0003757526, 0.002979167, 0.0211115, 
    0.06934631, 0.161765, 0.1059415, 0.1090891, 0.04240549, -1.341265e-06, 
    0.0002072314, -1.782906e-08, -5.862504e-09, 6.761217e-08, -6.904949e-05, 
    0.1076551, 0.213328, 0.07795016, 0.02655236, 0.001361231, 8.07779e-05,
  0.008612702, 0.0577831, 0.12307, 0.0009568684, 0.0255247, 0.02093209, 
    0.01305523, 0.008604567, 0.1054726, 0.0619157, 0.07835902, 0.05563957, 
    0.1059951, 0.1079287, 0.01945571, 0.0236427, 0.001987901, -0.0001127556, 
    0.003025463, 0.004765781, 0.001016075, 6.399085e-05, 0.0001658584, 
    0.1291701, 0.175283, 0.01158867, 0.03673806, 2.942205e-05, 1.875157e-07,
  -5.372574e-09, -5.491655e-05, 0.0004629133, -7.539822e-07, 0.006347195, 
    0.009132134, 0.004638183, 0.05467713, 0.04497922, 0.1667812, 0.1661281, 
    0.1676078, 0.2157898, 0.2021717, 0.1170395, 0.03534597, 0.07099693, 
    0.08665186, 0.03058977, 0.05201672, 0.1219542, 0.02060618, 0.03005149, 
    0.03373512, 0.03497289, 0.03260374, 0.004089429, 0.0002956849, 
    0.0003566587,
  -7.39631e-07, 0, -1.46933e-06, 9.282389e-06, 2.889062e-05, 0.000351817, 
    0.0009815437, 0.01839018, 0.009298611, 0.01439816, 0.106541, 0.07885869, 
    0.03915907, 0.06664185, 0.03020617, 0.005049553, 0.004644516, 0.01576014, 
    0.008859063, 0.002912953, 0.01355165, 0.02936731, 0.0187575, 0.02796439, 
    0.006551004, 0.01852587, 0.001680761, 0.005082182, -8.787538e-05,
  0, -6.322604e-07, -5.00217e-08, 0.008277742, 0.007865738, 0.002743364, 
    -6.306096e-05, 0, 0.0007412895, 0.004344632, 0.0001357116, 0.002266832, 
    0.02025117, 0.02410409, 0.02339877, 0.01372054, 0.008501014, 0.003262882, 
    0.004444534, 0.0002540641, -0.0001337736, 0.02232242, 0.03051133, 
    0.01135324, 0.01621264, 0.02871061, 0.0005048388, -9.047472e-05, 
    -0.0001109052,
  4.796169e-06, 0.0003794217, -5.652495e-08, 0.001574605, 0.000648381, 0, 0, 
    0, 0, 0, 0, 0.00780883, 0.01394524, 0.02793373, 0.01508139, 0.03493081, 
    0.02221755, 0.02099367, 0.01224594, 0.0006376221, 0, -2.095592e-05, 
    0.0005473698, 0.0176232, 0.03730283, 0.0172809, 0.02442297, 0.001503066, 
    0.0001233189,
  -1.082729e-05, 0, 0.0002470764, 0.0006041992, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002464385, 0.006640268, 0.004397736, 0.002497448, 0.0004901875, 
    0.005085078, 0.009478696, -8.69784e-06, 0.001219827, 0, 0, 0.000852299, 
    0.01169315, 0.003797567, 0.01260717, 0.00274749, 0.001986391,
  0.0005360738, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.313986e-06, 0, 0, 0, 
    -6.180413e-06, 0.000135254, 0.0004098339, 0, 0, 0, 0.003148558, 
    0.008748157, 0.003229071, 0.001241525, 0.004982785,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.848825e-05, -6.672883e-05, 0, 0, 0, 0,
  7.774938e-05, 0, -3.68421e-06, -1.657245e-06, 0, 0, -1.737325e-06, 
    -6.677705e-06, -1.9686e-06, -3.914308e-07, 0, 0, 0, 0, 0, 0.0004858565, 
    0, -3.126253e-06, 0, 0, 0.001783053, 0, -1.638676e-05, -1.392195e-06, 0, 
    0, -7.266574e-06, 0.002403107, -3.551537e-05,
  0.005850736, 0.003423715, 0.0001822289, 0.0003392209, 0.004854121, 
    0.003870693, 0.00836759, 0.005511285, 2.742366e-05, 0.001387555, 
    -1.830474e-05, 8.920466e-06, -1.831692e-05, 0.002368475, 0.00421702, 
    0.005156858, 0.000401561, 0.001515724, 0.0005577743, 0.001174763, 
    0.0004759053, -2.707226e-05, 0.002278935, 0.001522562, 0.0002064662, 
    0.007192633, 0.01013719, 0.009518711, 0.006289697,
  0.008268749, 0.0008966038, 0.0002622285, 0.03226857, 0.06714312, 
    0.05143894, 0.02924045, 0.007153574, 0.0001637064, -7.077748e-05, 
    0.0007337838, 0.001127666, 0.004874628, 0.03084311, 0.01510314, 
    0.005590278, 0.002157229, 0.01253969, 0.02886207, 0.02598572, 0.01265319, 
    0.01727667, 0.001064384, -1.428517e-05, 0.03037473, 0.05707961, 
    0.04275248, 0.01962424, 0.015647,
  0.002681593, 0.002355951, 0.006466704, 0.1433279, 0.06734421, 0.04849006, 
    0.02640064, 0.006672438, 0.03134306, 0.02538116, 0.006535854, 0.01169394, 
    0.00515204, 0.01917878, 0.0162537, 0.0129148, 0.03778843, 0.06656969, 
    0.1167455, 0.0471389, 0.01839841, 0.001598186, 0.0001672845, 
    0.0002481407, 0.05853652, 0.1005306, 0.07231951, 0.03152121, 0.02450979,
  0.0003645776, 0.0176429, 0.1768847, 0.0704347, 0.03368696, 0.0435376, 
    0.02474886, 0.0199338, 0.00451386, 0.02639955, 0.04583666, -0.0001282873, 
    0.002812146, 0.0489085, 0.04209861, 0.06925294, 0.1530264, 0.2386809, 
    0.1808845, 0.05477968, 0.01647234, 0.001332526, 6.947743e-07, 0.04326195, 
    0.1111211, 0.1391943, 0.1392419, 0.06754752, 0.02091517,
  0.0009054022, 0.1245454, 0.2610784, 0.1191739, 0.1078303, 0.1017586, 
    0.1148677, 0.0836003, 0.03789772, 0.003734842, 0.01691537, 0.03383449, 
    0.0711937, 0.1886719, 0.1504807, 0.1623733, 0.07882285, 0.001833682, 
    0.0002976781, -5.867156e-06, 3.647012e-07, 3.238324e-07, 0.00348753, 
    0.3402942, 0.3202892, 0.3356413, 0.1004744, 0.08185863, 0.0003199135,
  0.01669252, 0.2692906, 0.4566098, 0.02206318, 0.04008881, 0.06269286, 
    0.04042087, 0.03092877, 0.2922764, 0.2706323, 0.1706168, 0.1224854, 
    0.132892, 0.1063985, 0.01439682, 0.009618878, 0.002844718, 0.002157439, 
    0.003711884, 0.008426813, 0.001546641, 0.0002242207, 0.02222048, 
    0.4309114, 0.3368606, 0.03523077, 0.07614416, 0.02788356, 4.90003e-06,
  0.006130631, 0.004947115, 0.02634149, 0.002395461, 0.03572199, 0.05166136, 
    0.03846115, 0.09539565, 0.06918015, 0.2202617, 0.1522616, 0.1601987, 
    0.2123958, 0.1943319, 0.1002788, 0.09665941, 0.1237242, 0.1657835, 
    0.06313323, 0.1180845, 0.1744907, 0.05872836, 0.1001465, 0.08530103, 
    0.06812713, 0.08050897, 0.1206243, 0.08145486, 0.01412642,
  0.01951166, 0.0004676849, 0.0006798537, 0.01109952, 0.01880601, 0.03467222, 
    0.03275534, 0.04425561, 0.0242551, 0.01634385, 0.09452296, 0.06692325, 
    0.033625, 0.08021447, 0.04733059, 0.06001183, 0.05141599, 0.0591553, 
    0.07143383, 0.04767345, 0.07441491, 0.08870067, 0.08883129, 0.114691, 
    0.07006398, 0.06764384, 0.01877814, 0.0960047, 0.02130785,
  -2.427447e-06, 0.0002418652, 1.914122e-06, 0.01544305, 0.01228855, 
    0.004876236, 0.0003104609, -8.315987e-06, 0.002137498, 0.04659089, 
    0.003513803, 0.01166195, 0.04631121, 0.06087858, 0.08214646, 0.05354175, 
    0.04460357, 0.04201986, 0.01365706, 0.005755298, 0.003275501, 0.05309641, 
    0.07046347, 0.04850187, 0.08656543, 0.07778828, 0.009471305, 
    0.0003706813, -0.0003709699,
  0.001512787, 0.003328419, -4.219866e-05, 0.004112873, 0.002129923, 
    -4.587998e-06, 0, 0, 0, 0, 1.119034e-05, 0.02152935, 0.02944605, 
    0.0589192, 0.03834763, 0.07641485, 0.04208951, 0.04626788, 0.03596453, 
    0.002171558, 0, 7.24686e-05, 0.001901953, 0.03984678, 0.06284419, 
    0.03547197, 0.05962686, 0.01069877, 0.002173895,
  0.003993542, -1.825285e-06, 0.002224272, 0.001657272, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0003754157, 0.00891171, 0.009236748, 0.0108931, 0.004110973, 
    0.01461412, 0.02056944, 0.0031999, 0.001896106, -1.079927e-06, 
    -4.487157e-05, 0.00442268, 0.02185853, 0.01301647, 0.02177291, 
    0.01010776, 0.01268248,
  0.002336992, 3.921537e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.280434e-07, 
    -4.009228e-08, 0.0002564965, 0, 0, 0.0005504567, 0.0006131678, 
    0.001662909, -3.461296e-05, 0, 0.0002004893, 0.005719494, 0.02018415, 
    0.008282932, 0.007141235, 0.009370733,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.289291e-06, -8.135546e-05, 0.001121583, 0, 0, 0, 0,
  0.004323658, 4.428888e-05, 3.232504e-05, -2.178076e-05, 4.132732e-05, 
    -9.363222e-06, 0.0007702473, 0.00107331, 0.0001437442, 0.001115978, 
    -6.975107e-07, -3.416607e-06, 0, -1.533264e-06, -5.550362e-05, 
    0.0009322833, 0.002110993, 0.0002940015, 0.001209341, -1.526902e-05, 
    0.003043873, -3.281679e-05, 0.001373399, -1.756922e-06, 0, -5.220901e-06, 
    5.010485e-05, 0.003933067, 0.003243603,
  0.01866329, 0.009574756, 0.005296913, 0.002198876, 0.009856623, 0.01233428, 
    0.02196034, 0.01673999, 0.01560965, 0.01019894, 0.002913075, 
    0.0002650004, 0.0009114753, 0.007419819, 0.006746712, 0.01056954, 
    0.006030148, 0.006444597, 0.003159205, 0.006323603, 0.00628358, 
    0.0007744142, 0.01066543, 0.002931429, 0.00115823, 0.01562122, 
    0.03309087, 0.03619874, 0.02357404,
  0.02911193, 0.01386902, 0.03373174, 0.08368558, 0.1214687, 0.1045574, 
    0.08353534, 0.04876347, 0.03682984, 0.03070724, 0.04722717, 0.02804486, 
    0.0238337, 0.04577794, 0.03500151, 0.04430639, 0.0152923, 0.02428302, 
    0.06833236, 0.08957884, 0.07384492, 0.0516989, 0.02514726, 0.001447518, 
    0.0493973, 0.1226274, 0.09131406, 0.08505304, 0.06310116,
  0.03600439, 0.02424569, 0.04395102, 0.136213, 0.09569928, 0.09064974, 
    0.0540342, 0.07064834, 0.0756878, 0.06446154, 0.07183097, 0.05005646, 
    0.03292862, 0.04271739, 0.05222209, 0.05702757, 0.08687977, 0.1150577, 
    0.2640084, 0.1707786, 0.1167045, 0.08101587, 0.01657776, 0.01174249, 
    0.07009224, 0.09498921, 0.1410589, 0.1153227, 0.09141812,
  0.001718368, 0.01523433, 0.1861189, 0.05629854, 0.02429085, 0.03766741, 
    0.01237266, 0.01729128, 0.0004373865, 0.02467059, 0.04368369, 
    0.006664284, 0.00534285, 0.06076168, 0.06293868, 0.07710292, 0.1376641, 
    0.2472186, 0.1627, 0.04766618, 0.01981492, 0.0007347836, -3.09481e-09, 
    0.03536627, 0.08279555, 0.1404427, 0.1487319, 0.1005408, 0.01561309,
  0.001335003, 0.08886485, 0.215555, 0.1004742, 0.08698297, 0.07882649, 
    0.08544269, 0.06717196, 0.03106551, 0.002750672, 0.007966849, 0.02206551, 
    0.04549529, 0.1481836, 0.1292337, 0.1271386, 0.05967498, 0.001604571, 
    5.856988e-06, 3.475659e-07, 2.276218e-07, 3.380337e-07, 0.001024167, 
    0.2861719, 0.2666436, 0.2991808, 0.08376405, 0.07357494, 1.863314e-05,
  0.01375583, 0.2318592, 0.3660809, 0.01650458, 0.02438396, 0.03710333, 
    0.02234462, 0.01778085, 0.2353033, 0.2054302, 0.1157924, 0.08024544, 
    0.0885497, 0.08336826, 0.01264605, 0.007953389, 0.00198109, 8.042745e-05, 
    0.0008478715, 0.001223566, 0.0006320686, -2.096644e-05, 0.02247588, 
    0.3346014, 0.263034, 0.0338629, 0.05980513, 0.01358747, 3.678295e-06,
  0.002455857, 0.0005336969, 0.01874893, 0.02353276, 0.02138866, 0.03907742, 
    0.02571, 0.0724494, 0.05944321, 0.175995, 0.1217256, 0.1243992, 0.190098, 
    0.1633898, 0.07230247, 0.07644325, 0.1121649, 0.1152576, 0.05221809, 
    0.092457, 0.1481532, 0.0290055, 0.07076686, 0.05798611, 0.05989051, 
    0.06319042, 0.08231745, 0.06262605, 0.01408022,
  0.08512726, 0.009070973, 0.000675978, 0.004706529, 0.02750808, 0.02709579, 
    0.04995384, 0.03704383, 0.01975745, 0.0129817, 0.08411232, 0.05042183, 
    0.02354682, 0.07043462, 0.04587401, 0.04932322, 0.04253352, 0.04543225, 
    0.0562745, 0.03676433, 0.05088791, 0.08519536, 0.06887121, 0.08649376, 
    0.04781628, 0.07569986, 0.09777185, 0.1474153, 0.1727757,
  0.02535914, 0.0202705, 0.03800346, 0.03598235, 0.0232956, 0.02108714, 
    0.05263074, -3.419473e-05, 0.00753232, 0.06185337, 0.01990391, 
    0.03290044, 0.05469389, 0.08062288, 0.1294056, 0.1428831, 0.1237893, 
    0.1070965, 0.09944978, 0.0567051, 0.01644244, 0.1013956, 0.1439269, 
    0.09679499, 0.1826383, 0.1851705, 0.09239489, 0.0241339, 0.02330917,
  0.003479245, 0.006150597, 0.0008416314, 0.009299591, 0.009100011, 
    0.0001107115, -1.187424e-05, -1.555139e-06, 8.04328e-07, -2.161159e-07, 
    0.002465931, 0.02745469, 0.04599246, 0.08467075, 0.07313183, 0.1210745, 
    0.1140546, 0.131863, 0.1104438, 0.01057257, -2.151307e-05, 0.0007398553, 
    0.005257881, 0.06545369, 0.09818587, 0.09258753, 0.157358, 0.04731273, 
    0.01379776,
  0.01323406, 0.003020325, 0.007685808, 0.00415311, -5.391745e-05, 
    -2.148215e-07, 0, -1.535965e-06, 0, 0, 0, 0, 0.003357035, 0.01495015, 
    0.02507281, 0.02993501, 0.02371807, 0.05404851, 0.06871254, 0.01476528, 
    0.005390243, 0.001763754, 0.002374004, 0.00924604, 0.04148187, 
    0.03806143, 0.04501008, 0.03438656, 0.04542281,
  0.005005496, 0.0005574824, 0.0009217056, 0, 3.500127e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, -2.090292e-06, 0.0006309851, 0.001423815, -7.351533e-05, 
    0.0003718202, 0.002985972, 0.00250323, 0.002809457, 7.935715e-05, 0, 
    0.003409148, 0.0115016, 0.04288189, 0.01999593, 0.01779556, 0.01618227,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00089126, 8.600475e-05, -7.904715e-06, -8.17131e-09, -3.757263e-06, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.542892e-06, -2.173826e-06, 0, 0, 0, 0, 0, 0, 0, 
    -4.536137e-06, 0.001308146, 0.0003695053, -1.476006e-10, 3.655213e-05, 0, 
    -1.813499e-06, 0.001558798, 0.001789474, 0, 2.247219e-05, 0, 0,
  0.006730796, 0.005623158, 0.005536207, 0.0002781991, 0.001217616, 
    0.002705671, 0.003868626, 0.01197441, 0.02286302, 0.01673102, 
    0.002386898, 0.002677328, 0.0111947, 0.01249324, 0.008523032, 
    0.006012322, 0.01124381, 0.00578472, 0.008892598, 0.009131613, 
    0.009361469, 0.002232511, 0.002050182, 0.001571547, 1.266434e-05, 
    4.620589e-05, 0.001993229, 0.00602303, 0.008600348,
  0.04620545, 0.04128275, 0.03327928, 0.04602429, 0.06341377, 0.05875139, 
    0.0714674, 0.05826521, 0.08190377, 0.06572101, 0.06425655, 0.06817999, 
    0.05933998, 0.07985987, 0.04387908, 0.06557287, 0.04599547, 0.03117976, 
    0.03759149, 0.05597157, 0.05108989, 0.02912082, 0.03615739, 0.008350213, 
    0.02167969, 0.07674511, 0.1142311, 0.09826483, 0.06652153,
  0.07439257, 0.0497214, 0.05930179, 0.1104417, 0.1443626, 0.1310305, 
    0.1361314, 0.1420245, 0.1205711, 0.1140781, 0.1328675, 0.1136567, 
    0.05573123, 0.1009218, 0.08396223, 0.1068905, 0.08845118, 0.05727898, 
    0.1226318, 0.142769, 0.1426564, 0.1458943, 0.09761554, 0.03184137, 
    0.1246186, 0.1430257, 0.114492, 0.1052331, 0.1148917,
  0.02381962, 0.01243066, 0.06285694, 0.1144529, 0.09611157, 0.06951585, 
    0.03853815, 0.0659316, 0.06471783, 0.0488488, 0.05637091, 0.04658405, 
    0.04049382, 0.03702824, 0.08042774, 0.0692528, 0.1273624, 0.1346516, 
    0.253438, 0.1403772, 0.1318969, 0.08291419, 0.01413617, 0.006535026, 
    0.08398435, 0.09177719, 0.1360299, 0.101166, 0.06817748,
  -1.228719e-05, 0.01258868, 0.1649726, 0.04131132, 0.02293674, 0.03748773, 
    0.01003221, 0.02210975, 2.294604e-05, 0.02647284, 0.04459649, 
    0.004061989, 0.008784286, 0.0887693, 0.06174023, 0.06772789, 0.1266452, 
    0.1981762, 0.1392216, 0.03088216, 0.02063495, 0.0006991612, 
    -4.062333e-07, 0.02471787, 0.06113998, 0.1416629, 0.1281629, 0.07805118, 
    0.006120154,
  0.0007936645, 0.07542179, 0.1727957, 0.1013594, 0.07209504, 0.07116, 
    0.07903653, 0.05449554, 0.03316116, 0.002892724, 0.00560563, 0.02154315, 
    0.03375205, 0.1338224, 0.1132014, 0.1073469, 0.05757844, 0.0004380648, 
    1.054885e-05, 7.23601e-08, 4.847153e-08, 2.045701e-07, 0.000181969, 
    0.2438991, 0.2390662, 0.2759053, 0.0747713, 0.06174341, 1.879484e-06,
  0.01474955, 0.2063476, 0.3038127, 0.01440834, 0.02523189, 0.02883674, 
    0.01849515, 0.01539785, 0.1939711, 0.1568831, 0.08613864, 0.06149901, 
    0.07892331, 0.06929485, 0.01506844, 0.008318854, 0.001426905, 
    -7.780681e-05, 0.0006879823, -2.640412e-06, -5.98198e-05, -8.373585e-07, 
    0.01861553, 0.2844633, 0.2109969, 0.04558557, 0.06406429, 0.008304144, 
    0.0002075144,
  0.002105332, 6.692422e-05, 0.01560312, 0.01260073, 0.01167153, 0.0328498, 
    0.02270769, 0.0720266, 0.06094532, 0.1455143, 0.1120291, 0.1097546, 
    0.1747485, 0.1487615, 0.06283244, 0.0601497, 0.1035641, 0.09964973, 
    0.04968445, 0.07936727, 0.1354339, 0.02702763, 0.05083906, 0.05109573, 
    0.05366888, 0.06009852, 0.05732686, 0.0499764, 0.01458584,
  0.05364916, 0.001361, 0.0001494031, 0.002574291, 0.0248299, 0.02902856, 
    0.06101193, 0.02614922, 0.02013878, 0.01048636, 0.08589826, 0.04136305, 
    0.02005114, 0.06590462, 0.04284042, 0.04077645, 0.03862853, 0.0376606, 
    0.0447152, 0.02318401, 0.03264096, 0.06707084, 0.05302337, 0.0701858, 
    0.03768824, 0.06024185, 0.08004734, 0.12686, 0.1546164,
  0.04314461, 0.0497068, 0.06966733, 0.08431684, 0.06188111, 0.06068353, 
    0.1217701, 0.0002179447, 0.01462248, 0.07701133, 0.0292088, 0.06498156, 
    0.06962933, 0.08961189, 0.1175681, 0.1224283, 0.1124724, 0.1031534, 
    0.1264763, 0.06912179, 0.05991147, 0.1201274, 0.1332818, 0.09053686, 
    0.1306556, 0.1541783, 0.08308326, 0.04208959, 0.05582166,
  0.05225482, 0.05257349, 0.05129667, 0.02198057, 0.05253711, 0.02952287, 
    0.0003959156, 0.002409299, -7.532732e-06, -1.772e-05, 0.0107915, 
    0.05761612, 0.06546935, 0.1376093, 0.1357724, 0.1799701, 0.1857081, 
    0.2317852, 0.157483, 0.06054252, 0.001336231, 0.01808904, 0.06985656, 
    0.113563, 0.1409421, 0.1695137, 0.2454858, 0.1354875, 0.06331599,
  0.06238222, 0.01300095, 0.02189268, 0.007654227, 0.006249675, 0.008503584, 
    0.001217256, -1.661983e-05, 0, 0, 0, 0, 0.006065893, 0.02077, 0.02885664, 
    0.03255422, 0.07050289, 0.1387755, 0.2320507, 0.03885054, 0.02146028, 
    0.0167961, 0.01212828, 0.02166778, 0.07509752, 0.06577599, 0.09922135, 
    0.09300522, 0.09900287,
  0.02480132, 0.004415603, 0.001164927, 8.262299e-05, 0.0003065091, 
    0.002509165, 0, 2.936391e-05, 0, 0, 0, 0, 0, -1.197631e-05, 0.003854297, 
    0.004517985, 0.0006441524, 0.004622472, 0.01167678, 0.005010599, 
    0.009091211, 0.004616185, -0.0001179985, 0.009602845, 0.02567757, 
    0.07191366, 0.05887948, 0.03653934, 0.03062997,
  0, 0, 0, 0, 0, 0, 0.0001032337, 0, 0, 0, 0, 0, 0, 0, 0, -2.179655e-06, 
    1.326529e-06, 0, 0, 0, 0, 0, -0.0001293449, 0.001826222, 0.003212135, 
    0.0001367857, -3.203206e-07, 0.0001395964, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -9.383631e-05, -0.0003574492, 0.006573272, -1.793836e-05, -3.23454e-06, 0, 
    0.0001711008, -8.64538e-05, -4.08748e-05, -3.110437e-09, 0, 0, 
    -2.307641e-08, 0.0002986565, 0.0001125254, -0.0002576837, 0.0009200297, 
    0.002166267, 0.002479538, -9.367411e-05, -1.664959e-05, -0.0001223418, 
    0.004942814, 0.008216976, 0.01192338, 0.005599496, 0.005399605, 
    0.001274595, 0.001152828,
  0.02924184, 0.02752674, 0.02527961, 0.02550967, 0.02697039, 0.02502702, 
    0.01864884, 0.04229356, 0.04208269, 0.04554883, 0.02903594, 0.02878458, 
    0.04788225, 0.07325352, 0.08765981, 0.07574622, 0.08918431, 0.06130882, 
    0.04772865, 0.02913767, 0.04708989, 0.06629222, 0.06625812, 0.05119907, 
    0.03496699, 0.03427059, 0.03586194, 0.04199721, 0.03798424,
  0.08646432, 0.09264232, 0.1056883, 0.1188716, 0.1123324, 0.1143162, 
    0.129828, 0.1121319, 0.1401569, 0.1331551, 0.1361327, 0.1458421, 
    0.1425792, 0.1513073, 0.118538, 0.1354912, 0.1010395, 0.1333719, 
    0.1203994, 0.1350347, 0.1094715, 0.1062741, 0.09527084, 0.04107023, 
    0.0811657, 0.1525387, 0.1801987, 0.1486209, 0.1002489,
  0.08452888, 0.05776927, 0.04758894, 0.09423382, 0.1203698, 0.1238654, 
    0.1323138, 0.1347821, 0.1259404, 0.1185863, 0.1148547, 0.1123425, 
    0.07957716, 0.116987, 0.09358689, 0.1286974, 0.115511, 0.0699231, 
    0.1238497, 0.1536349, 0.1568928, 0.1679804, 0.1187953, 0.07492702, 
    0.1235433, 0.1435161, 0.1188634, 0.1055063, 0.1256327,
  0.00994582, 0.001645591, 0.0469065, 0.1046796, 0.09447464, 0.05837772, 
    0.02438834, 0.05210418, 0.0566497, 0.03287755, 0.04182941, 0.04295228, 
    0.03067838, 0.03732047, 0.06963276, 0.05803972, 0.1027341, 0.124947, 
    0.2295168, 0.102254, 0.1065262, 0.07180555, 0.01449678, 0.00364772, 
    0.08206514, 0.0795826, 0.1297304, 0.08948526, 0.06364141,
  3.72932e-06, 0.01129575, 0.1627377, 0.04869338, 0.02113356, 0.03835375, 
    0.006890747, 0.02582197, 1.395866e-06, 0.01387336, 0.03789767, 
    0.002595276, 0.005353938, 0.08756939, 0.0614007, 0.0721555, 0.1154436, 
    0.1619031, 0.1185644, 0.0111854, 0.02662361, -7.789366e-06, 1.873376e-08, 
    0.01179453, 0.04560072, 0.1387453, 0.1156377, 0.05158479, 0.002971977,
  0.0001282773, 0.07490018, 0.1395414, 0.09551379, 0.05485306, 0.07275226, 
    0.06899038, 0.03631104, 0.03439962, 0.002563408, 0.003116153, 0.02228602, 
    0.02767527, 0.1113458, 0.1052525, 0.08824479, 0.05927089, 0.0005683133, 
    5.944859e-07, -6.486733e-09, -2.622388e-10, 3.807368e-08, 0.0004655429, 
    0.1899613, 0.1972997, 0.2247991, 0.07402225, 0.03521182, 3.000469e-07,
  0.01682616, 0.1698632, 0.2433956, 0.01303105, 0.03375376, 0.02293002, 
    0.01191366, 0.01221387, 0.1462121, 0.1186225, 0.0554667, 0.05185941, 
    0.06092201, 0.05592472, 0.01721211, 0.009339161, 0.001449246, 
    -3.517851e-05, 0.0007535774, -9.680332e-06, -0.0001334267, 4.686313e-07, 
    0.003543971, 0.2289992, 0.1470666, 0.05469146, 0.06979531, 0.005027188, 
    8.887775e-05,
  0.00121081, 3.797642e-05, 0.008139093, 0.006434542, 0.01495069, 0.02562455, 
    0.02001998, 0.06845886, 0.0641676, 0.1228192, 0.09839039, 0.08990489, 
    0.1509343, 0.1284305, 0.05068798, 0.04784522, 0.09979761, 0.08500366, 
    0.04183964, 0.0735689, 0.1293435, 0.02033864, 0.03538869, 0.04278957, 
    0.04690861, 0.05798684, 0.04445736, 0.04078216, 0.01595677,
  0.03326327, 0.0001113732, -1.820928e-05, 0.0009975748, 0.01926273, 
    0.01884906, 0.04145526, 0.02490884, 0.02222062, 0.00754996, 0.08789325, 
    0.03391941, 0.01752164, 0.05978522, 0.03590782, 0.02758464, 0.03671543, 
    0.03242492, 0.03127674, 0.02108859, 0.03266746, 0.06709743, 0.04286053, 
    0.06930817, 0.03233004, 0.05598691, 0.05981025, 0.1111041, 0.1190797,
  0.02505356, 0.05091789, 0.06512126, 0.08037065, 0.08622074, 0.07819302, 
    0.1186291, 0.001656524, 0.02304972, 0.08140512, 0.02170105, 0.09236998, 
    0.06486763, 0.08832879, 0.1025626, 0.09435432, 0.09016092, 0.09413861, 
    0.1145744, 0.0443302, 0.07970149, 0.09322658, 0.1038811, 0.08428752, 
    0.08845023, 0.1335185, 0.06140196, 0.03182587, 0.06229464,
  0.08735673, 0.09628388, 0.09060521, 0.08373247, 0.1129509, 0.1046367, 
    0.001777874, 0.03916929, 0.01627049, 0.01350591, 0.0638249, 0.1222457, 
    0.1265855, 0.1808057, 0.1699775, 0.1776874, 0.1934777, 0.2245338, 
    0.1531259, 0.1041855, 0.02271996, 0.05553947, 0.1365926, 0.1597587, 
    0.1903811, 0.1654305, 0.2481361, 0.1297371, 0.07554312,
  0.1206761, 0.09949517, 0.09988848, 0.1230849, 0.1581367, 0.0916553, 
    0.02405109, 1.882949e-05, 4.617086e-05, -1.063368e-05, 0.00492805, 
    0.0008213573, 0.01871905, 0.03569172, 0.04783634, 0.06086384, 0.1243104, 
    0.1926059, 0.2940583, 0.1159107, 0.05378872, 0.08355155, 0.04570718, 
    0.04704064, 0.1283789, 0.1268277, 0.1315635, 0.1294582, 0.1536777,
  0.05610788, 0.0218037, 0.009798932, 0.006276542, 0.01883693, 0.02070157, 
    0.008483552, 0.004920431, 6.553611e-05, 0, 0, 0, 0, 0.004696334, 
    0.009568031, 0.04903629, 0.01280389, 0.02162475, 0.02171522, 0.03204099, 
    0.02188736, 0.01242358, 0.003892209, 0.02242209, 0.06993061, 0.1055763, 
    0.107209, 0.09734689, 0.06509297,
  0.0001149343, -2.87178e-05, -1.229018e-06, 0, 0, 0, 0.001891331, 0, 0, 0, 
    0, 0, 0, 0, 0.01357863, 0.01982018, 0.007462295, 0.01705507, 0.002632413, 
    1.257175e-05, 0, -0.0003728429, 0.007525565, 0.01001718, 0.02564717, 
    0.003031628, -4.127464e-05, 0.01815604, -7.30651e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.959096e-06, 0.0009348413, 
    3.10926e-05, 0.001231868, 0.0002477365, -5.997825e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.87945e-06, -7.317223e-06, 0, 0,
  0.005751668, 0.01518849, 0.02387616, 0.01128999, -8.012862e-05, 
    -0.0002944376, 0.01187537, -7.656013e-05, 1.34644e-05, -4.369467e-05, 
    -2.637391e-07, -1.628614e-06, -0.0004394332, 0.009480952, 0.01589115, 
    0.03353389, 0.03791384, 0.05352143, 0.03716537, 0.03319791, 0.01177542, 
    0.003277327, 0.005974563, 0.01719539, 0.03649902, 0.04231725, 0.02766541, 
    0.02727389, 0.01402461,
  0.1165242, 0.1108455, 0.08469354, 0.1063737, 0.08407799, 0.08320387, 
    0.1035521, 0.08161844, 0.05682613, 0.09445177, 0.07357452, 0.0766435, 
    0.1061814, 0.1173767, 0.1571461, 0.1683315, 0.1588286, 0.163747, 
    0.1298552, 0.1474037, 0.1332016, 0.1501288, 0.1484682, 0.1358075, 
    0.141944, 0.1091501, 0.1142832, 0.1379728, 0.1299315,
  0.1054464, 0.1157709, 0.1333842, 0.1506523, 0.1356395, 0.1373715, 
    0.1685969, 0.1556921, 0.1635618, 0.1455714, 0.1544676, 0.1625986, 
    0.1694517, 0.1574846, 0.1405326, 0.1423869, 0.1179332, 0.1338274, 
    0.1384078, 0.1376169, 0.1348504, 0.123424, 0.1372324, 0.09514605, 
    0.104647, 0.1804408, 0.1633464, 0.1582476, 0.1282346,
  0.086463, 0.06580286, 0.0382042, 0.07392919, 0.1018031, 0.1092956, 
    0.1265467, 0.1188011, 0.1100671, 0.1173772, 0.1054625, 0.1004598, 
    0.06789791, 0.1257686, 0.08992228, 0.1077208, 0.1065479, 0.0720797, 
    0.1013715, 0.1430942, 0.1541176, 0.1781763, 0.110985, 0.0748595, 
    0.108284, 0.1436329, 0.1139419, 0.1131487, 0.1117989,
  0.002565917, 0.0003619793, 0.04152016, 0.1088011, 0.08353122, 0.04636892, 
    0.0286462, 0.04089058, 0.0477153, 0.02916226, 0.03953221, 0.04118568, 
    0.02729923, 0.04086234, 0.06790195, 0.04740553, 0.08268084, 0.1118351, 
    0.2004611, 0.09457734, 0.1040866, 0.0500325, 0.007740181, 0.0007144416, 
    0.0750734, 0.06705532, 0.1261978, 0.07909962, 0.02508235,
  3.746608e-06, 0.009179822, 0.151379, 0.05681428, 0.01972697, 0.03576671, 
    0.006133542, 0.01751745, 8.616602e-06, 0.003498277, 0.02614942, 
    0.001726906, 0.006528839, 0.09084105, 0.06006797, 0.07559531, 0.09513154, 
    0.1244647, 0.1039259, 0.005964803, 0.02170477, -5.911329e-06, 
    5.590764e-10, 0.004703218, 0.03073182, 0.141795, 0.1085188, 0.03607824, 
    0.0009603607,
  1.707993e-06, 0.06553348, 0.1097081, 0.0825126, 0.04474168, 0.07405686, 
    0.05906592, 0.03262555, 0.03456741, 0.002145821, 0.004648527, 0.01879906, 
    0.02255243, 0.08923833, 0.07417299, 0.08087328, 0.0501715, 0.0005982183, 
    6.104978e-07, 8.695913e-09, 0, 1.238622e-08, 0.0002259414, 0.1439074, 
    0.1645877, 0.1698783, 0.06650344, 0.009620016, 1.001179e-07,
  0.02224491, 0.1519801, 0.1937068, 0.01095982, 0.03279326, 0.01964488, 
    0.0100841, 0.01129298, 0.1095131, 0.09472568, 0.03308971, 0.04519108, 
    0.04497294, 0.04215919, 0.01906782, 0.01059646, 0.002793204, 0.003308823, 
    0.00022342, -9.989699e-06, -8.494107e-05, 1.489526e-06, 5.434499e-05, 
    0.1801843, 0.08590004, 0.06227073, 0.09079789, 0.009732557, 2.807433e-05,
  0.0004433483, 0.0001505047, 0.00350009, 0.006312367, 0.02034928, 
    0.02231968, 0.02184943, 0.06522186, 0.06450751, 0.1095602, 0.08193129, 
    0.07798524, 0.1259838, 0.1056804, 0.04396483, 0.04169603, 0.09367813, 
    0.071638, 0.03412757, 0.07609001, 0.124288, 0.01558533, 0.02951878, 
    0.03533697, 0.03528952, 0.06126964, 0.03801123, 0.03134886, 0.01333,
  0.0242261, 0.001675555, -1.944574e-05, 0.001004688, 0.01657374, 
    0.009474767, 0.03165223, 0.02198501, 0.02142873, 0.005020373, 0.07984079, 
    0.02362755, 0.01473287, 0.05703947, 0.02415413, 0.01249084, 0.03302362, 
    0.0234539, 0.01107731, 0.01600386, 0.03451169, 0.07120015, 0.03996624, 
    0.06637433, 0.02588721, 0.05440355, 0.05222113, 0.09272445, 0.08520679,
  0.02229323, 0.05039587, 0.05154354, 0.06696251, 0.09155141, 0.07430695, 
    0.09636925, 0.005900121, 0.05030565, 0.08011844, 0.02441519, 0.06854594, 
    0.05765438, 0.07138523, 0.08292394, 0.07560733, 0.07821256, 0.0835323, 
    0.07128288, 0.02618403, 0.05812213, 0.0686718, 0.08839549, 0.07002026, 
    0.06945449, 0.1206325, 0.05800886, 0.02287997, 0.06281211,
  0.09117442, 0.1133145, 0.1080443, 0.1535659, 0.1127459, 0.1166675, 
    0.01414459, 0.08161412, 0.03494475, 0.03775942, 0.1006661, 0.1433741, 
    0.164611, 0.1918628, 0.1787752, 0.1782484, 0.1935903, 0.2240326, 
    0.173953, 0.1136313, 0.0521313, 0.06152857, 0.1348049, 0.1486089, 
    0.1909221, 0.1477965, 0.2475068, 0.1095042, 0.08149792,
  0.1565029, 0.1517659, 0.1929142, 0.2346244, 0.2550775, 0.2342272, 0.118673, 
    0.001335243, 0.001162123, 0.01170248, 0.01909021, 0.00977614, 0.04642483, 
    0.08266658, 0.08129261, 0.1065742, 0.1526156, 0.2415608, 0.3139652, 
    0.1869698, 0.08345392, 0.1218375, 0.101969, 0.1041711, 0.1633007, 
    0.1566652, 0.1419258, 0.1402584, 0.1704851,
  0.1270227, 0.07754839, 0.05092103, 0.05761259, 0.1053805, 0.1549946, 
    0.1467356, 0.1366443, 0.04464674, 0.007972877, 0, 0, -0.0001190042, 
    0.02148967, 0.05970616, 0.09626434, 0.04892527, 0.03685983, 0.08434178, 
    0.1023436, 0.07995357, 0.05612794, 0.0355899, 0.06846409, 0.1075048, 
    0.1357776, 0.1800479, 0.1267681, 0.1110311,
  0.008209018, 0.01262766, 0.002179352, 0.001221765, 0.01584655, 0.02553314, 
    0.01814563, 0.001224499, 0.0003684458, 0, 0, -2.539555e-07, 0, 
    0.001055255, 0.03022695, 0.03823163, 0.04613848, 0.05376984, 0.02808453, 
    0.005960463, 0.005407878, 0.01063698, 0.01899705, 0.01623815, 0.04050541, 
    0.01195484, 2.63985e-05, 0.06371678, 0.02038763,
  0.003238543, -9.528439e-05, -2.117331e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001022395, 0.01499154, 0.01478353, 0.01612712, 0.01396193, 0.01026834, 
    0.0001475316, 0, -1.146161e-05, -0.0001221365, -0.0009056836, 
    0.0005349577, -5.528332e-09, 0, -0.000796065, 0.005233258,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.748793e-06, 2.038361e-05, 
    0.0002058607, 0.01085147, 0.004399417, 0.0001274045, 0, 0, 0, 
    -1.037644e-09, 0.01947315, 0.000611551, -0.001961021, -0.000909151, 0, 0,
  0.04853756, 0.08043733, 0.07876286, 0.05427569, -5.797434e-05, 
    0.0003117399, 0.04942842, 0.0005236921, -0.0001951304, -0.0002692542, 
    -1.169568e-05, 6.76595e-05, -0.0003276217, 0.04072656, 0.06203247, 
    0.07734136, 0.104215, 0.1084731, 0.08993328, 0.06696313, 0.05781535, 
    0.05224116, 0.05818302, 0.08087726, 0.0979417, 0.09775563, 0.1280728, 
    0.09022263, 0.0615911,
  0.1667505, 0.1639833, 0.1279036, 0.1490812, 0.1488742, 0.1657121, 
    0.1928576, 0.1362531, 0.1043116, 0.1428018, 0.1294584, 0.1113759, 
    0.1522246, 0.1595186, 0.2084812, 0.2005723, 0.1996161, 0.2112043, 
    0.17117, 0.1732978, 0.1728345, 0.2000476, 0.2158971, 0.206004, 0.2002503, 
    0.1530243, 0.1474845, 0.1631516, 0.1849196,
  0.1101887, 0.1258857, 0.1387772, 0.1762967, 0.1581924, 0.1464453, 
    0.1810664, 0.1635021, 0.1712957, 0.155663, 0.1653804, 0.1605304, 
    0.1692732, 0.1538917, 0.1515645, 0.139641, 0.1175273, 0.1342617, 
    0.123164, 0.1385354, 0.1487771, 0.1314854, 0.1459646, 0.1185153, 
    0.1099461, 0.1665899, 0.1741754, 0.1457619, 0.1301303,
  0.07671525, 0.06592557, 0.0321533, 0.05988038, 0.08708067, 0.0975402, 
    0.1271512, 0.1175699, 0.10368, 0.1094136, 0.09652308, 0.08765675, 
    0.05677473, 0.1278166, 0.08877425, 0.1030719, 0.09426104, 0.07226849, 
    0.08390341, 0.1345913, 0.1599103, 0.1733562, 0.1053959, 0.06819014, 
    0.09494548, 0.1431805, 0.1087864, 0.1064006, 0.1039787,
  0.0006292469, 0.0005401847, 0.03910111, 0.122443, 0.06848919, 0.04968737, 
    0.02196578, 0.02923373, 0.04021038, 0.01904262, 0.04919689, 0.04448604, 
    0.02667228, 0.04282701, 0.06669975, 0.04326544, 0.06027986, 0.09955651, 
    0.181393, 0.07941121, 0.09057128, 0.03849836, 0.002565647, -1.383712e-05, 
    0.06413308, 0.06269728, 0.1001763, 0.06983395, 0.01444293,
  2.109758e-06, 0.007423257, 0.1283258, 0.04823362, 0.01450665, 0.03765076, 
    0.009295742, 0.01351549, 0.0001303874, 0.0004925135, 0.01519564, 
    0.001632235, 0.004960496, 0.09843336, 0.06099887, 0.07158735, 0.08932003, 
    0.09517418, 0.08436679, 0.006907851, 0.01506194, -1.127239e-07, 
    7.184325e-09, 0.004617732, 0.02166519, 0.1356074, 0.09771577, 0.02943282, 
    -1.847629e-07,
  0.0002153181, 0.05656422, 0.08711511, 0.07802814, 0.05020377, 0.08264928, 
    0.05854937, 0.0297831, 0.0323871, 0.002312667, 0.003026163, 0.01159562, 
    0.02140576, 0.07078607, 0.05889288, 0.07613009, 0.0478336, 0.0006515106, 
    8.302576e-08, 1.068641e-09, 0, 2.582874e-11, 0.0008158213, 0.100059, 
    0.1377007, 0.1248485, 0.05264313, 0.0008321554, 2.805338e-08,
  0.03152668, 0.1431855, 0.1471152, 0.01923396, 0.03136242, 0.01920548, 
    0.009859901, 0.009787703, 0.07794251, 0.09478605, 0.02048691, 0.03551411, 
    0.03413316, 0.04132929, 0.01861296, 0.01111837, 0.006025591, 0.00121013, 
    2.190762e-05, 1.01352e-05, 0.0004348482, 2.935472e-06, 0.003225998, 
    0.1460071, 0.05527434, 0.06224734, 0.1105554, 0.00703904, 9.493794e-05,
  0.001288649, 7.503951e-05, 0.00258385, 0.006373304, 0.009421581, 
    0.01898669, 0.02078438, 0.06099843, 0.07020593, 0.1045581, 0.07268355, 
    0.07465722, 0.1118967, 0.08826531, 0.04076339, 0.03257319, 0.08267264, 
    0.07339957, 0.03424155, 0.0886704, 0.1275156, 0.0134093, 0.02371236, 
    0.02825447, 0.02754023, 0.06657091, 0.0296744, 0.02245377, 0.009196938,
  0.0080402, 0.0005231482, -4.353811e-07, 0.001397678, 0.01637711, 
    0.007140429, 0.01198341, 0.01545098, 0.01967959, 0.002854428, 0.06808481, 
    0.01924595, 0.01499082, 0.05016102, 0.01760769, 0.00548102, 0.03926544, 
    0.01925128, 0.01211614, 0.01721095, 0.0370358, 0.07854241, 0.03091267, 
    0.07140195, 0.02302459, 0.05283403, 0.03875323, 0.06989354, 0.06030294,
  0.02119791, 0.0478126, 0.03622758, 0.05414822, 0.08432062, 0.07302884, 
    0.07846342, 0.01032359, 0.08671407, 0.07534856, 0.02425986, 0.05158048, 
    0.05707491, 0.06411953, 0.07635078, 0.06589734, 0.06709254, 0.07136934, 
    0.04139881, 0.01743368, 0.03745034, 0.05369144, 0.07874587, 0.06111129, 
    0.06710238, 0.108373, 0.05261441, 0.01719653, 0.06539655,
  0.09419671, 0.1080737, 0.09665758, 0.1816823, 0.0894064, 0.1004981, 
    0.03603882, 0.1106731, 0.05054259, 0.04890358, 0.1073606, 0.1302779, 
    0.1715101, 0.1805927, 0.1873045, 0.1701923, 0.2051015, 0.2098568, 
    0.1623982, 0.1321116, 0.083094, 0.05610518, 0.115252, 0.1359704, 
    0.1694147, 0.1334501, 0.2096821, 0.1118025, 0.08388988,
  0.1771584, 0.1974091, 0.2522769, 0.248976, 0.2384904, 0.2150415, 0.1340403, 
    0.01200757, 0.0191536, 0.04524916, 0.07344393, 0.03316189, 0.1313644, 
    0.126481, 0.1220148, 0.1403852, 0.1626247, 0.2377288, 0.3091289, 
    0.211547, 0.1099327, 0.1512677, 0.169461, 0.1872277, 0.1731774, 
    0.1596227, 0.1272967, 0.1490348, 0.1741031,
  0.1656615, 0.1465389, 0.2009412, 0.1821191, 0.2005423, 0.2495012, 
    0.2314709, 0.2499047, 0.1872692, 0.05589769, 0.01533126, 0.0009982859, 
    0.001840775, 0.05599608, 0.09502146, 0.1685439, 0.09355653, 0.08071534, 
    0.1452204, 0.1373355, 0.1239965, 0.1147061, 0.08248824, 0.1629993, 
    0.1836938, 0.2090473, 0.2042158, 0.1870418, 0.1692249,
  0.04585986, 0.03907195, 0.0312032, 0.1288394, 0.1368725, 0.1165633, 
    0.1154594, 0.07383046, 0.0335367, 0.0423228, 0.02144098, 0.01200114, 
    0.03101267, 0.07983855, 0.1193638, 0.09960631, 0.08626562, 0.07640942, 
    0.0708776, 0.05994992, 0.0406714, 0.0411416, 0.06626825, 0.03889108, 
    0.1119501, 0.03558722, 0.000280291, 0.08413956, 0.05216199,
  0.02666161, 0.01859129, 0.01377738, 0.01518791, 0.01600685, 0.01343262, 
    0.01081929, -4.631803e-05, 0, 0, 9.30843e-05, 0.01033771, 0.0129538, 
    0.01925164, 0.02510132, 0.02913775, 0.03374222, 0.02701987, 0.02384098, 
    0.01462898, 0.006611825, 0.0001621037, 0.005234743, 0.004389932, 
    0.007792829, 0.0002354103, -0.0008819308, 0.0002600187, 0.04009675,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.676701e-06, 0.0003262333, 0.01447836, 
    0.01892986, 0.01890995, 0.01660418, 0.006232093, 0.0001152946, 0, 0, 
    0.002752311, 0.05186916, 0.05074182, 0.02239884, 0.03522383, 
    -0.001302465, 6.967922e-08,
  0.0980105, 0.1421855, 0.1529444, 0.1130454, 0.001804433, 0.005456191, 
    0.09568183, 0.001622665, 0.002346084, -0.001225256, 0.000186284, 
    0.0002214295, 0.02141748, 0.1346278, 0.150993, 0.1708618, 0.1654254, 
    0.1481416, 0.1306322, 0.1178428, 0.1239332, 0.1281092, 0.13243, 
    0.1924775, 0.2011997, 0.1880925, 0.1824205, 0.1263863, 0.09053326,
  0.211491, 0.1888041, 0.1808104, 0.2129109, 0.2181577, 0.2231427, 0.2565684, 
    0.2129017, 0.1493649, 0.165736, 0.1663481, 0.1646372, 0.2149052, 
    0.188883, 0.2694206, 0.232355, 0.2012929, 0.21708, 0.188033, 0.198369, 
    0.2007746, 0.2416052, 0.2396626, 0.2343365, 0.2408635, 0.1842063, 
    0.1703759, 0.1691827, 0.2149684,
  0.1139891, 0.1232165, 0.1396981, 0.1753881, 0.1577898, 0.1458017, 
    0.1666028, 0.1673351, 0.1695318, 0.1532511, 0.1609513, 0.1549428, 
    0.173357, 0.1543704, 0.1499867, 0.1304288, 0.1094274, 0.1313863, 
    0.1204909, 0.1363087, 0.1595048, 0.1363706, 0.1495768, 0.1394114, 
    0.09900756, 0.1514699, 0.169986, 0.1387331, 0.1262385,
  0.0781137, 0.05841386, 0.02594788, 0.05510327, 0.08490181, 0.0932108, 
    0.1237314, 0.1167568, 0.1081551, 0.09573409, 0.08393132, 0.08982472, 
    0.04945679, 0.1248825, 0.08634189, 0.1030262, 0.09371042, 0.07642575, 
    0.06961298, 0.120448, 0.1618629, 0.1696717, 0.1190249, 0.0600672, 
    0.09119998, 0.1465444, 0.100118, 0.1044415, 0.09279656,
  5.234222e-05, 0.003517938, 0.03142425, 0.111842, 0.05816511, 0.03562889, 
    0.01429961, 0.02502544, 0.04301002, 0.0159379, 0.06202834, 0.0512009, 
    0.02527591, 0.04611921, 0.06695417, 0.04056536, 0.04978961, 0.09193741, 
    0.1481529, 0.06185187, 0.08801221, 0.02196725, 0.002739605, 
    -2.101977e-06, 0.06347512, 0.05516348, 0.09269412, 0.06328265, 0.01007004,
  1.91669e-06, 0.005186181, 0.1046364, 0.03932052, 0.01302574, 0.03858023, 
    0.01588354, 0.01395418, 2.66084e-06, 0.0004915746, 0.01441428, 
    0.001320886, 0.006323976, 0.09614037, 0.0535131, 0.06829375, 0.07500455, 
    0.08397849, 0.07167584, 0.009655913, 0.003249475, 1.044983e-07, 
    2.484974e-08, 0.002370774, 0.0166341, 0.1408847, 0.0937258, 0.03877098, 
    4.664711e-06,
  0.0005768651, 0.04669406, 0.0730744, 0.07534844, 0.04987957, 0.08980145, 
    0.06977452, 0.02908642, 0.02726462, 0.003156889, 0.005619033, 
    0.009558154, 0.02637414, 0.06419446, 0.06096699, 0.0647095, 0.04429869, 
    0.002072824, 7.641717e-06, 0, 0, 1.883774e-09, 0.0009629886, 0.07351088, 
    0.129693, 0.1092005, 0.03437359, -5.73023e-06, 3.755893e-08,
  0.05223534, 0.1491754, 0.1241723, 0.017162, 0.03429664, 0.02602954, 
    0.01427741, 0.008584268, 0.06398235, 0.09174184, 0.01896764, 0.0262201, 
    0.02929541, 0.03514442, 0.01700146, 0.0101528, 0.0007962101, 
    0.0009622908, 1.81746e-05, 0.001378414, 0.0004954368, 0.0001535798, 
    0.001509075, 0.1217079, 0.04374569, 0.0698006, 0.1243628, 0.004963616, 
    6.528186e-05,
  0.0008036529, 6.497547e-05, 0.001926019, 0.006603331, 0.01282089, 
    0.01741518, 0.008775543, 0.06265132, 0.0707987, 0.1025196, 0.06145487, 
    0.06976695, 0.09849501, 0.0767014, 0.0438805, 0.03167696, 0.06447658, 
    0.0750639, 0.03454112, 0.108244, 0.1402753, 0.02196193, 0.01953726, 
    0.02618617, 0.02361081, 0.06801355, 0.02761779, 0.009148736, 0.008984573,
  0.004163309, 2.351362e-05, 2.1743e-06, 0.0008650538, 0.01441138, 
    0.007331558, 0.006337184, 0.01271408, 0.02296886, 0.002618507, 
    0.06453174, 0.01888788, 0.01668187, 0.05122289, 0.01482025, 0.004970506, 
    0.03080795, 0.01433474, 0.02130983, 0.01405564, 0.03681136, 0.08692578, 
    0.02314149, 0.07119133, 0.01689788, 0.05274165, 0.04250816, 0.05261043, 
    0.06840857,
  0.02341837, 0.04002797, 0.03057884, 0.04507129, 0.07037421, 0.06305057, 
    0.06435026, 0.03487466, 0.1329668, 0.07489525, 0.0232396, 0.04328914, 
    0.05405967, 0.05726771, 0.06708927, 0.06568822, 0.05301786, 0.06900853, 
    0.03202783, 0.02012161, 0.02041987, 0.03994331, 0.07344541, 0.06323721, 
    0.06588121, 0.1019352, 0.04100042, 0.01572887, 0.06350878,
  0.09180625, 0.09488969, 0.0925327, 0.1865195, 0.06604843, 0.07591896, 
    0.07530431, 0.1152992, 0.05200056, 0.0509984, 0.112892, 0.1316065, 
    0.1738496, 0.1714127, 0.198016, 0.167981, 0.2179105, 0.2100524, 
    0.1433576, 0.125993, 0.09190764, 0.05984075, 0.107288, 0.1281386, 
    0.1689524, 0.1219001, 0.2062974, 0.1011311, 0.09074342,
  0.1961412, 0.1841259, 0.2609278, 0.2481301, 0.2163512, 0.1954002, 
    0.1340308, 0.06159968, 0.04203114, 0.08662967, 0.1441855, 0.09281789, 
    0.1777078, 0.1626363, 0.1382035, 0.1628063, 0.1805479, 0.2315098, 
    0.2905514, 0.2326434, 0.1315126, 0.1799358, 0.2252111, 0.2396878, 
    0.1950279, 0.1600669, 0.1218773, 0.1628931, 0.1862803,
  0.1776851, 0.2075153, 0.2695413, 0.2627434, 0.2647898, 0.2918684, 
    0.2581893, 0.273882, 0.2550638, 0.1272447, 0.04881462, 0.02119768, 
    0.04770485, 0.1164765, 0.1829237, 0.2139999, 0.1417481, 0.1412006, 
    0.1930249, 0.1870469, 0.1624131, 0.185262, 0.1678145, 0.2340677, 
    0.2648062, 0.26185, 0.2704061, 0.2425385, 0.2156523,
  0.05162469, 0.09867361, 0.1470255, 0.2200781, 0.2296351, 0.2049212, 
    0.1620403, 0.1374021, 0.09319857, 0.1024615, 0.05091599, 0.05909659, 
    0.1091937, 0.146595, 0.198756, 0.1137924, 0.09757401, 0.1253617, 
    0.1386551, 0.1403199, 0.09218408, 0.09775504, 0.1089349, 0.08554551, 
    0.1587668, 0.05514494, 0.01231987, 0.1246277, 0.08332344,
  0.08064879, 0.05916972, 0.04963804, 0.05889451, 0.05947641, 0.04486977, 
    0.0221377, 0.0007078745, -0.001194193, 0.01938718, 0.03142609, 
    0.04542109, 0.06050589, 0.06725408, 0.03965984, 0.03364341, 0.03484869, 
    0.04744199, 0.05448268, 0.06153758, 0.04118346, 0.02108778, 0.01039227, 
    0.004404223, 0.01279119, 0.002983671, -0.002491468, 0.03370275, 0.1155765,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -8.590152e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005929175, 0.03591404, 
    0.0494383, 0.05177244, 0.06388514, 0.04896549, 0.01563518, 0.008946348, 
    0.002072666, -4.844051e-05, 0.01804049, 0.1880745, 0.1529724, 0.08128556, 
    0.08537956, 0.02883077, 1.43448e-05,
  0.1875481, 0.1984502, 0.1997339, 0.1519067, 0.02128236, 0.02670459, 
    0.1529766, 0.009711899, 0.006248387, 0.004000575, 0.005622691, 
    0.006111812, 0.0532533, 0.2064821, 0.1899277, 0.2039168, 0.182911, 
    0.1719239, 0.2199649, 0.171575, 0.2224883, 0.252441, 0.2398038, 
    0.2993666, 0.2781792, 0.2086292, 0.226654, 0.1867065, 0.1600757,
  0.2340153, 0.2017802, 0.1765856, 0.2402429, 0.2442092, 0.2536099, 
    0.2973092, 0.2360272, 0.175926, 0.1941257, 0.2032894, 0.2126814, 
    0.249355, 0.2209922, 0.2801557, 0.2526897, 0.2123877, 0.2137147, 
    0.1897327, 0.226004, 0.2072722, 0.2568453, 0.2380937, 0.2584431, 
    0.2307312, 0.183231, 0.1699403, 0.1821921, 0.2538507,
  0.115565, 0.1179968, 0.1380177, 0.1796971, 0.1566296, 0.1408704, 0.1616175, 
    0.1728373, 0.1633599, 0.1468356, 0.1511819, 0.1558692, 0.1729063, 
    0.1493548, 0.1486906, 0.1226684, 0.1067828, 0.1302662, 0.1256068, 
    0.143545, 0.1514876, 0.125352, 0.1583317, 0.1412672, 0.09684061, 
    0.1465015, 0.1605565, 0.1311144, 0.123246,
  0.08441348, 0.05686557, 0.02378753, 0.05047548, 0.09186981, 0.08998981, 
    0.1230003, 0.09562621, 0.09635539, 0.08103105, 0.07665347, 0.08783331, 
    0.04873742, 0.1271491, 0.09036671, 0.1017221, 0.09094034, 0.07298295, 
    0.06275813, 0.1100855, 0.1572739, 0.1588599, 0.1239182, 0.04900148, 
    0.09309641, 0.1378632, 0.08947827, 0.1092009, 0.09200095,
  4.877505e-05, 0.001429179, 0.02820712, 0.1076791, 0.05449361, 0.03591114, 
    0.007483065, 0.01940483, 0.02960109, 0.008147486, 0.07775191, 0.05813384, 
    0.02357071, 0.04548762, 0.0578748, 0.02947804, 0.03939104, 0.0861617, 
    0.1378943, 0.05337985, 0.09157842, 0.02357014, 0.005917205, 0.0008490626, 
    0.05986755, 0.05228699, 0.09204154, 0.06631285, 0.006624277,
  1.823358e-06, 0.004236327, 0.08986273, 0.03960621, 0.01796996, 0.03894547, 
    0.01721365, 0.01421193, 8.331526e-08, 0.0001196524, 0.02089607, 
    0.003097081, 0.007216498, 0.07010598, 0.04645897, 0.06479886, 0.06151644, 
    0.06336671, 0.05895057, 0.008772705, 0.0001354676, 5.033856e-09, 
    1.337076e-08, 0.002364264, 0.01749839, 0.1326379, 0.08293925, 0.03408218, 
    -6.302628e-06,
  0.001704512, 0.04905779, 0.07380345, 0.07680818, 0.05117262, 0.0941897, 
    0.08054117, 0.02678863, 0.02608422, 0.004144448, 0.008727764, 0.01021875, 
    0.02499823, 0.05878359, 0.05471246, 0.06109506, 0.03913236, 0.002922536, 
    3.807569e-05, -2.125948e-11, 4.259611e-11, 2.382299e-09, 0.0005721248, 
    0.05365063, 0.1183255, 0.1074889, 0.01509384, 2.802591e-07, -7.884688e-06,
  0.1092439, 0.163668, 0.1076264, 0.01706254, 0.03315039, 0.03376211, 
    0.01980675, 0.006362174, 0.05829344, 0.09049898, 0.02262656, 0.01527481, 
    0.0269765, 0.0290811, 0.01539955, 0.01594021, 0.003384946, 0.0002654956, 
    0.003371733, -5.252984e-06, 0.0004153322, 2.803964e-05, 0.004164078, 
    0.1108562, 0.04018514, 0.06247885, 0.1237588, 0.003715359, 0.007264388,
  0.006024324, 8.84446e-05, 0.001512947, 0.01443643, 0.01364485, 0.01520569, 
    0.005530829, 0.05649232, 0.070421, 0.1042926, 0.05319184, 0.06366997, 
    0.09055461, 0.07605737, 0.04102109, 0.0390834, 0.04377449, 0.07771732, 
    0.03958476, 0.1239448, 0.1351506, 0.03426594, 0.01917676, 0.02094979, 
    0.02124524, 0.05937445, 0.02591484, 0.003200335, 0.01366574,
  0.0003838775, 1.191182e-06, 1.153013e-06, 0.0007431262, 0.01265123, 
    0.007575963, 0.004319211, 0.009108985, 0.03428584, 0.001921316, 
    0.06571499, 0.02294811, 0.01726172, 0.05286649, 0.01372377, 0.005434519, 
    0.02520016, 0.009806865, 0.01339873, 0.01145362, 0.03435091, 0.09471116, 
    0.02104012, 0.06837764, 0.01480915, 0.04965593, 0.04555527, 0.04684991, 
    0.04925799,
  0.02558794, 0.01757269, 0.01997587, 0.03383757, 0.06365445, 0.04805643, 
    0.0532507, 0.04338313, 0.1743131, 0.0810198, 0.01673921, 0.04669721, 
    0.05054907, 0.05232542, 0.06052223, 0.0524587, 0.0443932, 0.0519725, 
    0.02694418, 0.01505637, 0.01104202, 0.03949266, 0.06292652, 0.06575996, 
    0.06161363, 0.09534572, 0.03122273, 0.01355106, 0.06966974,
  0.09543311, 0.09207049, 0.08414863, 0.1706583, 0.05190158, 0.05495013, 
    0.1039799, 0.1100914, 0.04143182, 0.04944444, 0.1146512, 0.1382308, 
    0.1795101, 0.1766912, 0.2031434, 0.1634365, 0.2209328, 0.1936783, 
    0.1202522, 0.1185027, 0.08405129, 0.0613409, 0.1111836, 0.114833, 
    0.1765917, 0.1126533, 0.1781124, 0.09921374, 0.07237881,
  0.2039062, 0.1805261, 0.2407703, 0.2433293, 0.1936447, 0.1654158, 
    0.1194346, 0.09404424, 0.0906374, 0.1327491, 0.1655118, 0.1450704, 
    0.1886775, 0.1976608, 0.15966, 0.1796992, 0.1934183, 0.2184211, 0.271636, 
    0.2424151, 0.1504084, 0.2050463, 0.2390112, 0.2765002, 0.2142874, 
    0.1569382, 0.120282, 0.1706239, 0.1891098,
  0.173043, 0.2705677, 0.2734131, 0.2900325, 0.3068188, 0.2986419, 0.2513616, 
    0.2906403, 0.3078206, 0.1681694, 0.09641573, 0.1114156, 0.07537651, 
    0.1349882, 0.209273, 0.2395411, 0.1849443, 0.1890387, 0.2412153, 
    0.230446, 0.1825493, 0.2853748, 0.2490155, 0.2818372, 0.3159594, 
    0.3480048, 0.2827724, 0.2496573, 0.2376367,
  0.1041814, 0.1428072, 0.2043031, 0.291929, 0.3297573, 0.3147901, 0.2540807, 
    0.2583689, 0.1855399, 0.1729362, 0.1086161, 0.1537534, 0.1769346, 
    0.2161653, 0.2748762, 0.1454436, 0.1267495, 0.1540541, 0.2102806, 
    0.208183, 0.1194871, 0.1545536, 0.2529286, 0.1581912, 0.1965741, 
    0.07291602, 0.04471258, 0.1450415, 0.1114838,
  0.1697828, 0.1422437, 0.1105826, 0.1209888, 0.1257514, 0.1220715, 
    0.0948497, 0.04396021, 0.05170697, 0.07153527, 0.06766798, 0.07331432, 
    0.09281716, 0.1239673, 0.129872, 0.08809659, 0.05559462, 0.09405929, 
    0.1202043, 0.1040047, 0.09016181, 0.110446, 0.08138746, 0.01039764, 
    0.03149229, 0.007113433, 0.01589416, 0.07693754, 0.1646079,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.692992e-05, -2.692992e-05, -2.692992e-05, -2.692992e-05, 
    -2.692992e-05, -2.692992e-05, -2.692992e-05, 0,
  0.0002840183, 0.0001694444, -5.375794e-11, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.367746e-06, 0.0003935203, 0.07625142, 0.06616335, 0.08683121, 0.129998, 
    0.133035, 0.07424547, 0.04290663, 0.02092523, 0.004345085, 0.05002764, 
    0.2303437, 0.1755193, 0.1176577, 0.1711196, 0.07922576, 0.002679704,
  0.2055646, 0.2378625, 0.212854, 0.2162931, 0.08044438, 0.0944239, 
    0.1712665, 0.04919759, 0.02765334, 0.0488019, 0.01423507, 0.0362935, 
    0.08774523, 0.2497547, 0.2222295, 0.2047706, 0.2050294, 0.2233108, 
    0.2624264, 0.2108062, 0.2495466, 0.295354, 0.2912482, 0.3923836, 
    0.2873334, 0.2012167, 0.2220204, 0.1960614, 0.1870659,
  0.2367342, 0.2206618, 0.2108482, 0.2295694, 0.2339822, 0.2562712, 
    0.3168112, 0.2371275, 0.1955307, 0.2135096, 0.2228265, 0.2431158, 
    0.2547272, 0.2248255, 0.2780697, 0.2386349, 0.227347, 0.2179718, 
    0.1849712, 0.2448221, 0.2217408, 0.2621289, 0.2377157, 0.2449886, 
    0.2261185, 0.1695428, 0.1679733, 0.174197, 0.2467821,
  0.1046312, 0.113768, 0.1453332, 0.1801066, 0.1528934, 0.1391231, 0.1642343, 
    0.1767504, 0.1664697, 0.1564489, 0.146306, 0.1620583, 0.1795811, 
    0.1768555, 0.150228, 0.1190087, 0.1038688, 0.1280714, 0.1313298, 
    0.1299786, 0.1432838, 0.1284157, 0.167076, 0.1329304, 0.07955064, 
    0.1428603, 0.1612036, 0.1368964, 0.1197478,
  0.08830158, 0.0649703, 0.02439448, 0.05544651, 0.09385598, 0.08930982, 
    0.1175552, 0.08854973, 0.09738181, 0.05433835, 0.07299344, 0.08554928, 
    0.05861606, 0.1407232, 0.09228197, 0.103055, 0.08609626, 0.07721899, 
    0.05641548, 0.1041497, 0.1497303, 0.1317092, 0.1149754, 0.03809346, 
    0.1006414, 0.1261975, 0.0847282, 0.1119737, 0.10761,
  0.0004209535, 0.0002544036, 0.03823235, 0.09904736, 0.04647794, 0.0272947, 
    0.008367981, 0.01597009, 0.02342441, 0.005545649, 0.07159986, 0.03570876, 
    0.02264869, 0.04031108, 0.04972955, 0.0312592, 0.03607901, 0.07145254, 
    0.125181, 0.0456178, 0.08407255, 0.02300143, 0.009235642, 0.0004244549, 
    0.05388198, 0.04961352, 0.09106107, 0.07379244, 0.004530262,
  1.678607e-06, 0.004774285, 0.0984567, 0.03604349, 0.02272113, 0.03819665, 
    0.01166393, 0.01256283, 4.325052e-09, -1.115625e-05, 0.05696496, 
    0.01104434, 0.007675905, 0.06195544, 0.06606792, 0.06291747, 0.0471454, 
    0.05098335, 0.05636904, 0.003672727, 3.336013e-06, 7.46857e-09, 
    9.105301e-09, 0.002108096, 0.02322438, 0.1435475, 0.09377542, 0.01785224, 
    1.622757e-06,
  0.005276978, 0.0623537, 0.07085455, 0.07432369, 0.05368318, 0.08973929, 
    0.08068289, 0.02502943, 0.01527845, 0.00392343, 0.01457673, 0.009622228, 
    0.0259521, 0.05999446, 0.05894912, 0.06368668, 0.03948161, 0.003999253, 
    0.0001920502, 1.790118e-09, 7.585336e-10, 5.274345e-08, 0.000376962, 
    0.05434822, 0.1299484, 0.1176734, 0.01687028, 6.751865e-07, 0.008125525,
  0.2082038, 0.1748517, 0.1022863, 0.01956778, 0.03188084, 0.0314437, 
    0.02250203, 0.004459708, 0.07527671, 0.1005137, 0.03423334, 0.01931623, 
    0.02554827, 0.02699719, 0.01572557, 0.0121889, 0.005114235, 0.0002173865, 
    0.008080094, -5.0914e-06, 0.002213202, 1.345119e-06, 0.01348544, 
    0.1188418, 0.04790507, 0.044344, 0.1298701, 0.003942067, 0.02844969,
  0.01333327, 7.223369e-05, 0.001334813, 0.01843352, 0.01794706, 0.01885995, 
    0.006688739, 0.05726716, 0.07459473, 0.1139146, 0.06904327, 0.06418222, 
    0.09569322, 0.08368462, 0.05224972, 0.047079, 0.03828567, 0.08381557, 
    0.0495429, 0.1348759, 0.1518271, 0.03678221, 0.02164203, 0.0205458, 
    0.02213125, 0.04643244, 0.02395802, 0.002828317, 0.01046963,
  -7.194564e-05, -5.648261e-06, 1.337074e-06, 0.001057704, 0.008146429, 
    0.008343922, 0.004765542, 0.005648397, 0.04039225, 0.005215916, 
    0.07183192, 0.02958954, 0.01847943, 0.05354238, 0.01043725, 0.006697562, 
    0.02374875, 0.01124724, 0.005034247, 0.009343765, 0.02518179, 0.1032925, 
    0.01845632, 0.06332427, 0.01646401, 0.04824605, 0.03473343, 0.03592321, 
    0.03936296,
  0.02332738, 0.009750949, 0.01099945, 0.01872199, 0.06481645, 0.03919132, 
    0.04598548, 0.07565621, 0.1942622, 0.07631613, 0.01190699, 0.05220994, 
    0.0492828, 0.05230813, 0.04960912, 0.05009262, 0.04321712, 0.04655096, 
    0.02640019, 0.008071218, 0.007563103, 0.03795202, 0.06074636, 0.06361365, 
    0.05341973, 0.09593064, 0.03001555, 0.01822572, 0.07700507,
  0.09121467, 0.09118876, 0.08529633, 0.1627522, 0.04292722, 0.04231431, 
    0.1050925, 0.09696607, 0.03306963, 0.04545536, 0.116032, 0.1318076, 
    0.1802899, 0.1767063, 0.1927006, 0.155705, 0.2132043, 0.1873418, 
    0.1107796, 0.1054269, 0.06932481, 0.05721749, 0.1146559, 0.1196808, 
    0.173704, 0.1004086, 0.1752761, 0.09308466, 0.07676835,
  0.2198985, 0.1753549, 0.2230934, 0.2225709, 0.1797685, 0.1488721, 
    0.1148392, 0.1173524, 0.1189839, 0.1456798, 0.1716898, 0.1740475, 
    0.1795854, 0.1967764, 0.1554418, 0.1804476, 0.1961583, 0.2217141, 
    0.2639519, 0.254499, 0.1696588, 0.2215405, 0.2457674, 0.2923148, 
    0.2082384, 0.1670199, 0.1177134, 0.1715064, 0.1762102,
  0.1803826, 0.271341, 0.2711074, 0.3027206, 0.3163419, 0.2992042, 0.2441638, 
    0.3074036, 0.3500124, 0.2174452, 0.1679826, 0.1440685, 0.1011588, 
    0.1525172, 0.2033159, 0.2413723, 0.2011143, 0.2100691, 0.2602617, 
    0.2648557, 0.2009814, 0.3173772, 0.3273096, 0.3250865, 0.3361083, 
    0.3915604, 0.2643067, 0.2351609, 0.2364427,
  0.1298622, 0.1548654, 0.2075242, 0.3196908, 0.3834276, 0.3455192, 
    0.3011637, 0.3234182, 0.3031794, 0.2485874, 0.154812, 0.1755879, 
    0.2216284, 0.2628376, 0.3390569, 0.2223152, 0.1780229, 0.1738813, 
    0.2460339, 0.2195927, 0.1226806, 0.2052597, 0.2568268, 0.1961205, 
    0.179688, 0.1185681, 0.07618991, 0.1476556, 0.1149835,
  0.1870828, 0.2146778, 0.1701331, 0.1463053, 0.1537665, 0.1928985, 
    0.1433089, 0.08269006, 0.09414194, 0.1076907, 0.1010374, 0.1240466, 
    0.1650174, 0.1823662, 0.200528, 0.1445879, 0.1307336, 0.1171283, 
    0.1534547, 0.1680712, 0.1502632, 0.1586871, 0.1285231, 0.03559443, 
    0.06846153, 0.01014424, 0.02706062, 0.08960765, 0.1715747,
  0.002885053, 0.002619625, 0.002354198, 0.00208877, 0.001823342, 
    0.001557915, 0.001292487, 0.0008760469, 0.0008197398, 0.0007634327, 
    0.0007071256, 0.0006508185, 0.0005945113, 0.0005382043, -0.00024381, 
    -5.376531e-05, 0.0001362794, 0.0003263241, 0.0005163688, 0.0007064135, 
    0.0008964582, 0.002520886, 0.002652576, 0.002784267, 0.002915957, 
    0.003047647, 0.003179337, 0.003311027, 0.003097395,
  -0.002324194, 0.001531891, 0.0007328395, -1.683752e-06, 0, -5.788262e-06, 
    0, 0, 0, 0, -3.578059e-06, 7.331951e-05, 0.004252374, 0.1058109, 
    0.06541005, 0.08129141, 0.1328717, 0.176687, 0.1345307, 0.09458347, 
    0.06056878, 0.02484219, 0.144198, 0.230754, 0.1573068, 0.1064929, 
    0.1607907, 0.1894016, 0.0252807,
  0.1905488, 0.2471258, 0.2027548, 0.2468309, 0.1558058, 0.1566019, 
    0.1814251, 0.1023225, 0.04582926, 0.14348, 0.09710219, 0.08173276, 
    0.1246515, 0.2556099, 0.2345387, 0.2153937, 0.2152047, 0.2398185, 
    0.277662, 0.2269595, 0.2438404, 0.3064911, 0.3043824, 0.422257, 
    0.2827285, 0.1901317, 0.2220711, 0.2030534, 0.186741,
  0.2371058, 0.2253668, 0.2289917, 0.2352894, 0.2318948, 0.2682635, 
    0.3323267, 0.2411255, 0.2033693, 0.22958, 0.2168754, 0.2483692, 
    0.2446355, 0.2264692, 0.2787554, 0.2475851, 0.2406096, 0.2013719, 
    0.1887215, 0.2406135, 0.2269343, 0.2556782, 0.2380814, 0.2464458, 
    0.1993614, 0.1632414, 0.1591125, 0.1694952, 0.2360171,
  0.110833, 0.1204557, 0.1547028, 0.1876168, 0.1487322, 0.1479037, 0.163685, 
    0.1644474, 0.1668608, 0.1566105, 0.1428886, 0.1715124, 0.1927267, 
    0.1771801, 0.1449852, 0.111089, 0.1151463, 0.1266202, 0.1291037, 
    0.1305059, 0.1413246, 0.125178, 0.1628086, 0.1241078, 0.07904857, 
    0.1532331, 0.1400371, 0.1519569, 0.1332791,
  0.09206128, 0.06712885, 0.02146118, 0.05799432, 0.09489758, 0.08569199, 
    0.1110669, 0.08311941, 0.09353764, 0.04501423, 0.07531783, 0.06768522, 
    0.06365652, 0.1322894, 0.09309123, 0.1049419, 0.07057522, 0.0898684, 
    0.05031873, 0.1029105, 0.1211534, 0.1335371, 0.1252935, 0.02858375, 
    0.103882, 0.1283343, 0.0866963, 0.1168444, 0.1097502,
  0.001224765, 0.0001028462, 0.05873117, 0.09974083, 0.03166361, 0.02823341, 
    0.009282244, 0.01619428, 0.01476508, 0.005131125, 0.03716904, 0.01855426, 
    0.03160301, 0.03740488, 0.04005653, 0.03221699, 0.04238838, 0.0763675, 
    0.1312371, 0.04292168, 0.07445112, 0.02554462, 0.01015137, -4.694132e-05, 
    0.05996108, 0.04879193, 0.09084252, 0.08033352, 0.001500061,
  4.36794e-06, 0.01600476, 0.1400148, 0.0316352, 0.02907545, 0.05067873, 
    0.008177261, 0.01474649, 4.467397e-05, 0.0008108775, 0.08431073, 
    0.03395782, 0.01283778, 0.061189, 0.06541557, 0.06513424, 0.04672239, 
    0.05302951, 0.05528062, 0.002623634, 5.315061e-07, 4.536543e-08, 
    1.435209e-07, 0.002783174, 0.02656938, 0.156989, 0.09408523, 0.006978, 
    3.843643e-06,
  0.004223532, 0.08427061, 0.09180127, 0.0706193, 0.05876324, 0.09992725, 
    0.09867584, 0.03081293, 0.01184658, 0.003548962, 0.01635025, 0.0209706, 
    0.03206562, 0.07171483, 0.07369705, 0.06841834, 0.03760386, 0.004077883, 
    0.0001071387, 6.925339e-08, 9.577743e-09, 6.490258e-07, 0.001567128, 
    0.0766166, 0.1689139, 0.1360181, 0.008692073, 8.094884e-07, 0.001607817,
  0.2802067, 0.2148476, 0.1303757, 0.02464329, 0.03182069, 0.03069465, 
    0.02211709, 0.006083699, 0.08942796, 0.1167762, 0.05087303, 0.03713244, 
    0.03622275, 0.03252498, 0.01479714, 0.008053401, 0.00795936, 0.006553705, 
    0.0004834027, -3.162877e-05, 0.0002424251, 3.64809e-06, 0.01938197, 
    0.1432992, 0.07622464, 0.04296758, 0.1287136, 0.005235371, 0.06468923,
  0.00188061, 0.0001817679, 0.001997674, 0.01002324, 0.02691363, 0.02677632, 
    0.0100888, 0.06323911, 0.08482549, 0.1324552, 0.08041596, 0.07482778, 
    0.1168971, 0.1066772, 0.0658758, 0.05607652, 0.04125369, 0.09243862, 
    0.06691752, 0.1465536, 0.1659978, 0.04754174, 0.03387879, 0.02329228, 
    0.02401959, 0.0458192, 0.027795, 0.003119356, 0.008864064,
  -3.420188e-05, -1.257521e-05, 1.113043e-06, 0.001785044, 0.005564552, 
    0.008157904, 0.006833513, 0.002876801, 0.03710456, 0.02830407, 0.1005104, 
    0.03610219, 0.02154106, 0.05873462, 0.01093787, 0.009680416, 0.02010977, 
    0.01496156, 0.001462751, 0.009922701, 0.02457039, 0.1144137, 0.0188049, 
    0.05823655, 0.02170818, 0.05294941, 0.02884353, 0.03402076, 0.02203144,
  0.01441254, 0.006701487, 0.007218291, 0.0141482, 0.06635482, 0.03604285, 
    0.05108953, 0.1173858, 0.1927428, 0.07317561, 0.008115753, 0.06549642, 
    0.05385473, 0.05675677, 0.05483614, 0.0475874, 0.04851522, 0.05364995, 
    0.01890086, 0.01564426, 0.006057156, 0.04094068, 0.05732754, 0.06709385, 
    0.04654789, 0.09183685, 0.03487024, 0.01972506, 0.08965068,
  0.07916066, 0.09473635, 0.07361132, 0.1584839, 0.03895423, 0.03123734, 
    0.1005439, 0.07843955, 0.02952321, 0.04277372, 0.1147, 0.1259345, 
    0.1607567, 0.1731625, 0.1742207, 0.1524554, 0.220189, 0.1860274, 
    0.103577, 0.09149146, 0.05984899, 0.04389966, 0.1234108, 0.1128742, 
    0.1620239, 0.1017878, 0.1622892, 0.09069382, 0.06152441,
  0.2068222, 0.1575663, 0.2215476, 0.2169447, 0.1552372, 0.1314707, 
    0.09534341, 0.1355995, 0.1458296, 0.1570231, 0.1600834, 0.1643343, 
    0.1818401, 0.2027394, 0.1642517, 0.1794305, 0.1919194, 0.2258376, 
    0.2469589, 0.2602942, 0.1926492, 0.2015845, 0.2446013, 0.2987086, 
    0.2231994, 0.1592818, 0.1151367, 0.1793253, 0.1923358,
  0.1909515, 0.3047611, 0.2530697, 0.3051168, 0.3159758, 0.293637, 0.2524164, 
    0.3177318, 0.3823228, 0.2452784, 0.2159699, 0.1556039, 0.1244938, 
    0.1660849, 0.1895965, 0.2239614, 0.2137852, 0.2226015, 0.2815177, 
    0.2665291, 0.1937252, 0.3373871, 0.3744329, 0.3630269, 0.3461699, 
    0.4131269, 0.2518958, 0.2461878, 0.2504829,
  0.1121256, 0.1771327, 0.2269591, 0.3608768, 0.4478396, 0.3571166, 
    0.3046891, 0.3231044, 0.3256846, 0.2651265, 0.1957594, 0.2169766, 
    0.2390336, 0.2840692, 0.3284528, 0.2208894, 0.1792703, 0.1744313, 
    0.2433798, 0.2178645, 0.1456661, 0.2460564, 0.2933492, 0.2264217, 
    0.1754796, 0.1818506, 0.1179665, 0.1483514, 0.1474629,
  0.1742069, 0.1962118, 0.1815938, 0.1305444, 0.1340927, 0.1871103, 
    0.1515477, 0.1093857, 0.1375845, 0.1511987, 0.136527, 0.1654423, 
    0.2171585, 0.1927538, 0.2253554, 0.1723696, 0.196308, 0.2175285, 
    0.2133014, 0.2027478, 0.1915573, 0.1942255, 0.141678, 0.04562453, 
    0.09008254, 0.02214474, 0.03504823, 0.08630635, 0.1817326,
  0.007322111, 0.006927454, 0.006532797, 0.00613814, 0.005743483, 
    0.005348826, 0.00495417, 0.005313458, 0.005212031, 0.005110605, 
    0.005009178, 0.004907752, 0.004806325, 0.004704899, 0.002888232, 
    0.003330464, 0.003772696, 0.004214928, 0.00465716, 0.005099392, 
    0.005541624, 0.009325228, 0.00937908, 0.009432931, 0.009486782, 
    0.009540634, 0.009594485, 0.009648337, 0.007637836,
  0.02336146, 0.005978274, 0.01053564, 0.004766244, 0.0008449229, 
    -0.0002347623, -0.0005948729, -0.0001344659, 2.61303e-05, 0.0006933106, 
    -8.849106e-05, 0.00406252, 0.03451995, 0.1081036, 0.06174272, 0.07465912, 
    0.1352689, 0.1677174, 0.1579991, 0.1444231, 0.157028, 0.1260784, 
    0.2587851, 0.2171391, 0.1501777, 0.100787, 0.157203, 0.1875056, 0.06212506,
  0.1865405, 0.2554677, 0.1919626, 0.2592681, 0.2037094, 0.2007933, 
    0.1920654, 0.1641484, 0.111858, 0.2430481, 0.188261, 0.09730603, 
    0.1565888, 0.2503891, 0.2296237, 0.2130667, 0.2167582, 0.2362731, 
    0.301425, 0.2501584, 0.2497837, 0.3176529, 0.290812, 0.4440589, 
    0.2813691, 0.1800092, 0.2339039, 0.2192735, 0.1941324,
  0.2305031, 0.2281256, 0.2423362, 0.2558612, 0.2759827, 0.2647026, 
    0.3224841, 0.2613696, 0.2162578, 0.2285466, 0.2275875, 0.2605889, 
    0.2701299, 0.2239537, 0.2793351, 0.2440286, 0.2147742, 0.2138352, 
    0.1851469, 0.2376238, 0.2518257, 0.2313792, 0.2342299, 0.2517933, 
    0.2001797, 0.1654684, 0.1574922, 0.1735389, 0.2344005,
  0.1103941, 0.123662, 0.1673875, 0.1901257, 0.1440035, 0.128943, 0.1522542, 
    0.174867, 0.1901004, 0.1714308, 0.159894, 0.187805, 0.2271641, 0.1777006, 
    0.1396042, 0.116093, 0.1095287, 0.1240246, 0.1122864, 0.1249749, 
    0.1444195, 0.1283491, 0.1655445, 0.1231955, 0.08984049, 0.1671203, 
    0.1468389, 0.1335192, 0.1176844,
  0.08973247, 0.05868992, 0.02014764, 0.06452554, 0.097756, 0.08784559, 
    0.1094636, 0.09220681, 0.08699928, 0.04225488, 0.06694306, 0.05796009, 
    0.07185662, 0.1218414, 0.107518, 0.106691, 0.05898852, 0.08837067, 
    0.05060884, 0.1027434, 0.11353, 0.1118359, 0.1121484, 0.0236663, 
    0.102952, 0.1397102, 0.09352349, 0.1169317, 0.1098581,
  0.002824869, 0.0001683448, 0.06712471, 0.1104942, 0.02762699, 0.02922278, 
    0.01452301, 0.01676223, 0.0142771, 0.004916705, 0.02509518, 0.003344054, 
    0.03403559, 0.04093469, 0.04078071, 0.03903424, 0.03911531, 0.08529468, 
    0.1454722, 0.05199272, 0.07894967, 0.01853037, 0.007683172, -3.69389e-06, 
    0.08088519, 0.05212085, 0.1141617, 0.06815182, 0.0009800587,
  5.541808e-06, 0.01525081, 0.1653091, 0.02898707, 0.03803107, 0.05818427, 
    0.006803414, 0.008853077, 0.0008721639, 0.0009906131, 0.07272491, 
    0.04912021, 0.01517871, 0.06284485, 0.06089798, 0.06534756, 0.04935631, 
    0.05949376, 0.06600227, 0.003769685, 3.429621e-07, 7.619035e-08, 
    8.665819e-08, 0.001683775, 0.0405938, 0.1731813, 0.08457069, 0.00174852, 
    -5.504452e-06,
  0.004921835, 0.1068982, 0.1310802, 0.07946768, 0.06411432, 0.1101298, 
    0.1110504, 0.03826396, 0.01059306, 0.00352943, 0.01504376, 0.02719197, 
    0.03614491, 0.08103455, 0.07972544, 0.08496657, 0.0357262, 0.003649971, 
    5.94666e-05, -9.209475e-08, 2.807742e-08, -2.098392e-07, 0.002345267, 
    0.09865755, 0.205394, 0.1865643, 0.004728941, 9.31058e-07, 0.0001313535,
  0.2671608, 0.2751245, 0.1753916, 0.04075804, 0.03150344, 0.0342648, 
    0.02219674, 0.008189941, 0.1189811, 0.1537748, 0.06164587, 0.04705754, 
    0.04237511, 0.03254625, 0.01539768, 0.01249127, 0.008078271, 0.007132858, 
    -0.0001576559, 7.282825e-05, 0.001336913, -3.716935e-05, 0.02979395, 
    0.1799299, 0.1118783, 0.03806837, 0.1386961, 0.008092377, 0.04377146,
  0.001041601, 0.000336234, 0.0046369, 0.0224417, 0.04179011, 0.03409225, 
    0.02403619, 0.06732822, 0.09934875, 0.1410007, 0.09307204, 0.08273233, 
    0.1323989, 0.1226619, 0.08048572, 0.0543841, 0.04998768, 0.09084006, 
    0.07122972, 0.1650292, 0.174518, 0.0550652, 0.0474027, 0.03158256, 
    0.02445451, 0.0469595, 0.03272852, 0.006822421, 0.006219794,
  4.751597e-05, 2.765049e-06, 1.007832e-05, 0.003905902, 0.004615545, 
    0.00940311, 0.01205263, 0.008937966, 0.03533316, 0.04266633, 0.1273855, 
    0.03845599, 0.02383651, 0.0550036, 0.01346116, 0.01686851, 0.02976581, 
    0.01635317, 0.006574128, 0.0009806638, 0.02785259, 0.1214207, 0.02272037, 
    0.06299707, 0.02680032, 0.05896537, 0.02848875, 0.04433793, 0.01433031,
  0.004149776, 0.01077318, 0.005575472, 0.0129373, 0.0677869, 0.03524071, 
    0.04484299, 0.1412072, 0.194596, 0.08255643, 0.008958893, 0.06853294, 
    0.06673245, 0.06311911, 0.06471291, 0.04966187, 0.04842175, 0.05834341, 
    0.01171374, 0.008032587, 0.009648377, 0.04357485, 0.05710577, 0.07194076, 
    0.04467675, 0.1023464, 0.04051423, 0.02939925, 0.0763125,
  0.06939357, 0.09335375, 0.06807353, 0.1610613, 0.04244152, 0.03575572, 
    0.0952739, 0.05782559, 0.02422073, 0.03667034, 0.1175482, 0.1247894, 
    0.1473429, 0.1641627, 0.1593094, 0.1581206, 0.2146916, 0.1889087, 
    0.09460601, 0.0895196, 0.05511387, 0.042637, 0.1132459, 0.1146779, 
    0.1619924, 0.08829971, 0.1522468, 0.08032797, 0.06506778,
  0.1874171, 0.1549069, 0.2263485, 0.2044991, 0.1403567, 0.1197125, 
    0.0968706, 0.1471881, 0.1390423, 0.165564, 0.1522061, 0.1548227, 
    0.183648, 0.2102676, 0.1717244, 0.1723515, 0.1917174, 0.225627, 
    0.2345659, 0.2485944, 0.1841684, 0.2049409, 0.2447073, 0.2980488, 
    0.232362, 0.1724255, 0.1206136, 0.1851818, 0.1810119,
  0.1971665, 0.327818, 0.2769821, 0.3830854, 0.3380004, 0.2918318, 0.2482514, 
    0.3246671, 0.3966099, 0.2533024, 0.2349029, 0.1555422, 0.1269166, 
    0.1534959, 0.1790123, 0.2252796, 0.2180917, 0.2281114, 0.3009245, 
    0.2778659, 0.2069927, 0.322467, 0.3853447, 0.3856639, 0.354912, 
    0.4184095, 0.2621672, 0.2589384, 0.2419483,
  0.1280542, 0.1578591, 0.2115757, 0.382691, 0.4560579, 0.3578841, 0.3028149, 
    0.3232182, 0.3307639, 0.257386, 0.204571, 0.2343195, 0.2268827, 
    0.2872438, 0.322522, 0.2078355, 0.1627408, 0.1612131, 0.2503685, 
    0.1969363, 0.144133, 0.2576705, 0.2845371, 0.2421059, 0.163462, 
    0.2084021, 0.1467084, 0.1377235, 0.1406325,
  0.1537154, 0.1697122, 0.1557723, 0.1382406, 0.133397, 0.1703218, 0.1534203, 
    0.1208509, 0.1492067, 0.1903021, 0.1907213, 0.1788977, 0.2249602, 
    0.2153211, 0.2325531, 0.1916, 0.2212905, 0.2337112, 0.2459568, 0.2192178, 
    0.2232899, 0.2103813, 0.1572664, 0.07720304, 0.1085559, 0.02072829, 
    0.04537354, 0.07548632, 0.1949901,
  0.01425812, 0.01320771, 0.01215729, 0.01110687, 0.01005646, 0.009006043, 
    0.007955628, 0.009788658, 0.009936175, 0.01008369, 0.01023121, 
    0.01037873, 0.01052624, 0.01067376, 0.01021756, 0.0112874, 0.01235724, 
    0.01342709, 0.01449693, 0.01556677, 0.01663661, 0.01336876, 0.01320182, 
    0.01303487, 0.01286793, 0.01270099, 0.01253404, 0.0123671, 0.01509846,
  0.06188417, 0.01565153, 0.02441133, 0.01598232, 0.01456384, 0.002306861, 
    0.00727271, 0.007746764, 0.00638034, 0.001226452, 0.006391138, 
    0.03585936, 0.05319009, 0.1044492, 0.04696066, 0.0565262, 0.1328971, 
    0.1586233, 0.1490631, 0.1363515, 0.2053941, 0.2768015, 0.2642936, 
    0.206998, 0.141009, 0.1014612, 0.1481119, 0.1767442, 0.1027448,
  0.2043784, 0.2509941, 0.2008637, 0.2915278, 0.2721847, 0.2259323, 
    0.1999387, 0.2092979, 0.1713624, 0.28777, 0.2295878, 0.1378275, 
    0.1744162, 0.2543255, 0.2414157, 0.2155364, 0.2342812, 0.2617915, 
    0.3141792, 0.2482602, 0.2591714, 0.3179757, 0.2728736, 0.4664163, 
    0.2826868, 0.1774618, 0.2270527, 0.2545297, 0.2158805,
  0.2386769, 0.2397561, 0.2763134, 0.2922809, 0.3197921, 0.293768, 0.3206071, 
    0.2634886, 0.2380907, 0.2594303, 0.2341715, 0.2739614, 0.25222, 
    0.2311871, 0.2685627, 0.2545687, 0.2406786, 0.2202266, 0.1975711, 
    0.2512464, 0.268945, 0.2509108, 0.23973, 0.2430051, 0.1777327, 0.1573424, 
    0.1534116, 0.1855683, 0.233762,
  0.1189711, 0.1248336, 0.1710685, 0.2063262, 0.1446193, 0.146989, 0.1583991, 
    0.1628579, 0.1893506, 0.1601802, 0.1726089, 0.2054661, 0.2027709, 
    0.1750241, 0.1248809, 0.1107018, 0.1080682, 0.1243232, 0.1178416, 
    0.114784, 0.1354193, 0.1313325, 0.16735, 0.1296941, 0.09545238, 
    0.1581589, 0.1273161, 0.1281138, 0.1147822,
  0.0953341, 0.07303992, 0.02981503, 0.08322011, 0.1037719, 0.09386881, 
    0.1091522, 0.0946725, 0.08715899, 0.04666709, 0.05542243, 0.05090979, 
    0.06534991, 0.1146018, 0.114649, 0.1033738, 0.06387873, 0.0930387, 
    0.05629076, 0.1151022, 0.1189891, 0.1021607, 0.112235, 0.02397688, 
    0.09544673, 0.1359548, 0.09982519, 0.1110632, 0.1210615,
  0.004556129, 0.0003505309, 0.07575444, 0.1252696, 0.02018074, 0.03901201, 
    0.01922366, 0.01921064, 0.02399039, 0.006057371, 0.00975379, 
    0.0005699329, 0.03937704, 0.05223703, 0.0482556, 0.05073956, 0.04350342, 
    0.08554278, 0.1524924, 0.06068683, 0.09302722, 0.01304701, 0.004602644, 
    1.817135e-07, 0.08618622, 0.06435813, 0.1339155, 0.06925465, 0.0002695777,
  3.155395e-06, 0.0116974, 0.1455683, 0.02796321, 0.03434025, 0.05931411, 
    0.003083094, 0.00360272, 1.025155e-05, 0.0004062563, 0.02685141, 
    0.0249429, 0.01413621, 0.06442252, 0.05497053, 0.07188682, 0.0555091, 
    0.06389751, 0.0810595, 0.004111668, 3.637008e-07, 9.91458e-08, 
    7.492838e-08, 0.0002019277, 0.05081452, 0.1954566, 0.08950351, 
    0.000850612, 8.283685e-06,
  0.0005995234, 0.08169958, 0.1526772, 0.08093527, 0.06579033, 0.109457, 
    0.09236656, 0.04059791, 0.009673716, 0.006260299, 0.01617567, 0.01486373, 
    0.02998118, 0.06491557, 0.07200438, 0.08247974, 0.03741978, 0.006098222, 
    0.001148465, -6.423121e-06, 3.076229e-08, 0.0001550147, 0.001078946, 
    0.1093949, 0.1923609, 0.2163144, 0.004685567, 7.214686e-07, 1.731467e-05,
  0.2675889, 0.3435622, 0.1977095, 0.06300828, 0.03336355, 0.03293307, 
    0.02226806, 0.01029305, 0.1394484, 0.1753238, 0.05848357, 0.03907013, 
    0.03260277, 0.02851976, 0.01345647, 0.01170874, 0.007080168, 0.001656575, 
    -2.390992e-05, 8.958632e-05, 0.005723943, 0.004564405, 0.04826963, 
    0.1829917, 0.1306726, 0.03558418, 0.1211302, 0.01199532, 0.04228017,
  0.001132079, 0.0002966001, 0.012114, 0.03396202, 0.04970107, 0.03056083, 
    0.04070232, 0.06018342, 0.09696936, 0.115833, 0.08722378, 0.06746715, 
    0.1071241, 0.1041794, 0.0836326, 0.05313058, 0.05793642, 0.08651963, 
    0.08157534, 0.1463909, 0.1689645, 0.05466016, 0.06119481, 0.03733957, 
    0.02765457, 0.04394571, 0.04540979, 0.007315657, 0.002948768,
  1.365815e-05, 2.215208e-06, 0.0008378291, 0.006999122, 0.006631635, 
    0.01119734, 0.0169024, 0.01504372, 0.03787484, 0.05545564, 0.1226022, 
    0.03277775, 0.0235985, 0.05367514, 0.01111882, 0.01922192, 0.03596081, 
    0.01915958, 0.01244205, 0.001454592, 0.03501572, 0.1256629, 0.02280088, 
    0.06936095, 0.02895344, 0.06450339, 0.03403791, 0.04381436, 0.008972902,
  0.001526403, 0.006482777, 0.008536622, 0.01237903, 0.07102579, 0.03975531, 
    0.03808717, 0.1507647, 0.2020648, 0.08640133, 0.01162596, 0.06782098, 
    0.07267934, 0.07674806, 0.09263727, 0.05836612, 0.05024759, 0.06070599, 
    0.007283966, 0.003054092, 0.01594638, 0.04284003, 0.06272257, 0.0738705, 
    0.05031963, 0.1047498, 0.04956651, 0.03554404, 0.05849287,
  0.06035344, 0.09405962, 0.07309344, 0.1664874, 0.04714069, 0.02668888, 
    0.1024715, 0.04509798, 0.02025533, 0.02596737, 0.1173045, 0.1249537, 
    0.1364561, 0.1494763, 0.1562073, 0.1597094, 0.2077914, 0.1898875, 
    0.09751031, 0.08340681, 0.05860171, 0.03241324, 0.09814586, 0.1144793, 
    0.1650618, 0.09467924, 0.1454367, 0.08232458, 0.07735714,
  0.1914532, 0.1537893, 0.217001, 0.1977736, 0.1393358, 0.1368262, 
    0.09893954, 0.1494134, 0.1297619, 0.1633927, 0.1483187, 0.1480744, 
    0.181506, 0.2239707, 0.1873735, 0.1715415, 0.1788577, 0.2262725, 
    0.2291384, 0.2470914, 0.1727179, 0.2022545, 0.2657636, 0.2996261, 
    0.2458217, 0.1728897, 0.1341486, 0.1897123, 0.1825707,
  0.2362361, 0.3539295, 0.2779524, 0.3477868, 0.3159381, 0.3141899, 
    0.2548248, 0.3332152, 0.3946577, 0.2716873, 0.2473106, 0.1583805, 
    0.1362718, 0.1431139, 0.1950999, 0.2189522, 0.2160636, 0.2832207, 
    0.2826726, 0.2652679, 0.2209675, 0.3850779, 0.377148, 0.3565398, 
    0.3329299, 0.4103604, 0.2616633, 0.2685609, 0.2529227,
  0.1522557, 0.1913525, 0.2624469, 0.3921525, 0.4748372, 0.3704835, 
    0.2799014, 0.3375497, 0.3454133, 0.2684556, 0.1948842, 0.251917, 
    0.2200966, 0.275808, 0.3278463, 0.1972633, 0.1527596, 0.1688464, 
    0.2434198, 0.2124877, 0.1349741, 0.2716718, 0.2625651, 0.2587477, 
    0.1333505, 0.2233119, 0.1868646, 0.1507607, 0.161476,
  0.1331151, 0.1534023, 0.1452876, 0.1375772, 0.1531833, 0.1523893, 0.146366, 
    0.1263786, 0.1427404, 0.1803611, 0.1806371, 0.2077905, 0.2508851, 
    0.2132121, 0.2401879, 0.2059677, 0.1794342, 0.2110357, 0.237997, 
    0.2574214, 0.2322577, 0.2212157, 0.1572391, 0.09386614, 0.1141505, 
    0.04804079, 0.05319955, 0.08612634, 0.1894526,
  0.07344697, 0.06918188, 0.0649168, 0.06065173, 0.05638665, 0.05212156, 
    0.04785649, 0.04129569, 0.0397647, 0.03823371, 0.03670273, 0.03517174, 
    0.03364075, 0.03210976, 0.02876972, 0.03402761, 0.0392855, 0.04454338, 
    0.04980127, 0.05505915, 0.06031704, 0.06802224, 0.06856042, 0.0690986, 
    0.06963678, 0.07017496, 0.07071315, 0.07125133, 0.07685903,
  0.0899163, 0.03632374, 0.04382326, 0.04420722, 0.04468509, 0.01898697, 
    0.01510913, 0.008048198, 0.01071481, 0.007094273, 0.03918767, 0.05620306, 
    0.0712432, 0.1016021, 0.03767214, 0.0551956, 0.1187024, 0.1479517, 
    0.1311637, 0.1273638, 0.2085519, 0.3523703, 0.2697138, 0.2047571, 
    0.1374466, 0.1037304, 0.1450793, 0.1734396, 0.1057221,
  0.2184602, 0.24404, 0.2062081, 0.3049279, 0.3312264, 0.2347499, 0.2197476, 
    0.2312132, 0.2357684, 0.290293, 0.2512952, 0.1497397, 0.1842512, 
    0.2857274, 0.2475052, 0.2373887, 0.2699772, 0.2994015, 0.3251245, 
    0.2545491, 0.2933009, 0.3423433, 0.3072043, 0.5010046, 0.2664154, 
    0.1836529, 0.2694853, 0.2787637, 0.2276444,
  0.2555249, 0.2537009, 0.2782408, 0.370664, 0.3038462, 0.3163301, 0.3181458, 
    0.3149907, 0.2827842, 0.2952219, 0.2786371, 0.3076859, 0.2692172, 
    0.2349207, 0.2758809, 0.2405386, 0.2288206, 0.2319221, 0.1938246, 
    0.2500085, 0.2848307, 0.270498, 0.2482198, 0.2465957, 0.1876756, 
    0.1599204, 0.1713114, 0.196659, 0.2512545,
  0.1180698, 0.1413112, 0.1940432, 0.2162924, 0.1546345, 0.1488308, 
    0.1627846, 0.1746656, 0.2085562, 0.1863053, 0.1850709, 0.2036997, 
    0.1804556, 0.1570416, 0.120953, 0.1338857, 0.1214955, 0.1232147, 
    0.1299515, 0.1282256, 0.1307943, 0.1392017, 0.176745, 0.1401028, 
    0.1155953, 0.1517658, 0.1291166, 0.1424788, 0.1165159,
  0.1048341, 0.07833754, 0.04569275, 0.09898202, 0.1183131, 0.09768546, 
    0.1207487, 0.08936333, 0.08820737, 0.0666766, 0.03936584, 0.03125505, 
    0.06194516, 0.1246022, 0.1048117, 0.1169106, 0.07378103, 0.09561763, 
    0.05949479, 0.1198346, 0.1287807, 0.1044192, 0.1091446, 0.02856543, 
    0.08739059, 0.1491068, 0.09689503, 0.1202371, 0.1254285,
  0.00648796, 0.0003689197, 0.0690489, 0.1140133, 0.02206568, 0.03648817, 
    0.01590413, 0.02212278, 0.03625552, 0.004842889, 0.003771264, 
    0.0004019806, 0.03698774, 0.06803737, 0.05985714, 0.05718267, 0.05870554, 
    0.08963279, 0.1677834, 0.06475972, 0.09604447, 0.01517077, 0.005935817, 
    6.926331e-08, 0.05594431, 0.06901146, 0.1265415, 0.07994723, 0.001885065,
  1.073778e-06, 0.005143603, 0.1026357, 0.01795146, 0.02954878, 0.05260685, 
    0.001471951, 0.001165907, 3.207462e-06, 4.859887e-05, 0.006140009, 
    0.00757697, 0.01543886, 0.05146286, 0.05566632, 0.06729618, 0.06153587, 
    0.0644976, 0.08105338, 0.02458335, 1.848118e-07, -1.667497e-08, 
    6.178077e-08, 1.163338e-05, 0.06161567, 0.2167974, 0.08342868, 
    0.000575297, 5.521588e-06,
  0.001191668, 0.0513798, 0.1237694, 0.07204277, 0.06547635, 0.1037961, 
    0.08476841, 0.0408245, 0.007980966, 0.004019182, 0.01635042, 0.01141876, 
    0.02772117, 0.05216487, 0.06862312, 0.07185945, 0.03792703, 0.01094248, 
    0.001997837, 0.0001551599, 4.459541e-08, 6.670633e-06, 5.927458e-05, 
    0.07121202, 0.1383645, 0.1713665, 0.006855043, 5.329952e-07, -1.034263e-05,
  0.2163882, 0.3297725, 0.1303165, 0.07939755, 0.02925891, 0.03427452, 
    0.0244296, 0.009222353, 0.1299781, 0.1672397, 0.05311176, 0.03524418, 
    0.02706227, 0.02487124, 0.01110899, 0.009641225, 0.003162499, 
    4.066225e-05, -5.458369e-05, 0.0003325984, 0.003086802, 0.01115824, 
    0.03431364, 0.131767, 0.1374397, 0.02907066, 0.1180695, 0.01873767, 
    0.04589473,
  0.0009991002, 0.001181276, 0.02016929, 0.09267809, 0.05571458, 0.02811223, 
    0.04760529, 0.05527952, 0.08621274, 0.09804694, 0.08607041, 0.05372189, 
    0.08691454, 0.09098163, 0.08701853, 0.05562394, 0.05696399, 0.0765609, 
    0.09266306, 0.142687, 0.1728896, 0.04726136, 0.06816921, 0.04002901, 
    0.027515, 0.03572503, 0.03631141, 0.004899938, 0.001608747,
  1.253491e-05, 1.235052e-06, 0.006887572, 0.008058645, 0.01503496, 
    0.01311428, 0.0233373, 0.0160878, 0.04105883, 0.05854372, 0.0987187, 
    0.03448842, 0.02293092, 0.05704406, 0.0120265, 0.02256064, 0.03586114, 
    0.01653348, 0.01446237, 0.0009925128, 0.02417062, 0.1383726, 0.02296503, 
    0.06187383, 0.02950921, 0.06825215, 0.03002318, 0.03922638, 0.002410906,
  0.004293157, 0.006748767, 0.01087363, 0.01624635, 0.07518859, 0.03038095, 
    0.04040858, 0.1560026, 0.2148342, 0.0892565, 0.01682321, 0.0751469, 
    0.08182068, 0.09614614, 0.1161608, 0.06812122, 0.05453943, 0.06300718, 
    0.01137461, 0.001519778, 0.02333415, 0.04648926, 0.07146558, 0.06261966, 
    0.05303133, 0.1050313, 0.06296267, 0.04237056, 0.0467552,
  0.0536028, 0.09559225, 0.07986241, 0.1827668, 0.04403914, 0.02150433, 
    0.1136131, 0.03893907, 0.01737033, 0.01844118, 0.1124132, 0.1208896, 
    0.1357797, 0.1387348, 0.1577038, 0.1593204, 0.2145799, 0.18018, 
    0.1027767, 0.07958082, 0.06332619, 0.02593215, 0.09384668, 0.1211128, 
    0.1712866, 0.1142328, 0.1567122, 0.09260401, 0.0857779,
  0.1847561, 0.1740725, 0.2292714, 0.1893628, 0.1225097, 0.11405, 0.08695699, 
    0.1467623, 0.1224866, 0.1595836, 0.1414052, 0.1424279, 0.1946113, 
    0.2339005, 0.2043871, 0.1814151, 0.1751653, 0.2210352, 0.2332723, 
    0.248831, 0.1866632, 0.2183256, 0.2565913, 0.3396717, 0.2302547, 
    0.1781948, 0.147821, 0.2028898, 0.1769333,
  0.2415053, 0.3742223, 0.2982789, 0.3389317, 0.3266498, 0.3076041, 
    0.2875252, 0.3610525, 0.4249462, 0.315578, 0.2487395, 0.1373828, 
    0.1569582, 0.1414574, 0.2017016, 0.2016615, 0.2260741, 0.3017383, 
    0.2723483, 0.2829193, 0.287771, 0.373936, 0.4332891, 0.3592166, 
    0.3312369, 0.4220353, 0.2439416, 0.2629757, 0.2622889,
  0.1826778, 0.2335222, 0.2905671, 0.4031871, 0.4967479, 0.3819862, 
    0.3174996, 0.3871245, 0.3605674, 0.2809078, 0.2125897, 0.2335236, 
    0.2199075, 0.2720736, 0.3164207, 0.1875143, 0.1859771, 0.1993184, 
    0.245533, 0.210286, 0.1576477, 0.3368509, 0.3003209, 0.2948783, 
    0.1371561, 0.242794, 0.2214266, 0.1591924, 0.1675802,
  0.141227, 0.1805038, 0.1698615, 0.1435761, 0.1604853, 0.1310373, 0.1422818, 
    0.1323057, 0.1393893, 0.1748295, 0.185531, 0.2022, 0.2436388, 0.2027859, 
    0.2527569, 0.2195389, 0.1814171, 0.2042712, 0.2806088, 0.2663722, 
    0.2274656, 0.2322027, 0.1630364, 0.09681869, 0.1134975, 0.06212626, 
    0.04945113, 0.09087642, 0.1869232,
  0.1503744, 0.1446773, 0.1389803, 0.1332833, 0.1275862, 0.1218892, 
    0.1161922, 0.1060858, 0.1038447, 0.1016037, 0.09936265, 0.09712161, 
    0.09488057, 0.09263954, 0.08411256, 0.09251054, 0.1009085, 0.1093065, 
    0.1177045, 0.1261024, 0.1345004, 0.1507321, 0.1502722, 0.1498123, 
    0.1493524, 0.1488925, 0.1484326, 0.1479727, 0.154932,
  0.1050879, 0.07286543, 0.03549129, 0.06734918, 0.05725231, 0.05134323, 
    0.03522866, 0.02771749, 0.02795805, 0.03481917, 0.07211442, 0.06617235, 
    0.1010357, 0.1030376, 0.03328482, 0.03864888, 0.09808222, 0.1266696, 
    0.1324222, 0.1145249, 0.1944697, 0.3696703, 0.2826009, 0.234821, 
    0.1726926, 0.1105949, 0.1387273, 0.1727581, 0.1105165,
  0.2258997, 0.2533511, 0.2123982, 0.3226923, 0.3338705, 0.2495776, 
    0.2309247, 0.2210667, 0.2329495, 0.2863722, 0.2646553, 0.1686507, 
    0.2234965, 0.2907363, 0.2318562, 0.2356678, 0.2545527, 0.2760234, 
    0.3266187, 0.2568368, 0.343115, 0.3468433, 0.3486873, 0.5266832, 
    0.2387199, 0.1849178, 0.2493133, 0.3038087, 0.2394398,
  0.2615631, 0.2666524, 0.2516302, 0.3798787, 0.3084808, 0.3136398, 
    0.3599353, 0.3165663, 0.2591256, 0.2952539, 0.3019491, 0.2818414, 
    0.3033569, 0.2580569, 0.2826456, 0.262404, 0.2440099, 0.2497925, 
    0.2446262, 0.2790461, 0.2971659, 0.2794648, 0.2520587, 0.2629267, 
    0.1917812, 0.1683598, 0.183272, 0.2112227, 0.2539073,
  0.1339726, 0.1661509, 0.2052364, 0.2357881, 0.1574592, 0.1593441, 
    0.1766397, 0.1811971, 0.2145704, 0.2072526, 0.1907127, 0.2083259, 
    0.1722107, 0.1736918, 0.115485, 0.1225193, 0.1372138, 0.1566078, 
    0.1396636, 0.1311533, 0.1543519, 0.1487226, 0.1789451, 0.1486402, 
    0.1254402, 0.1465532, 0.1326861, 0.135307, 0.1373902,
  0.1178624, 0.08392341, 0.06068147, 0.1185086, 0.125696, 0.1067591, 0.13218, 
    0.09290245, 0.1003632, 0.06865776, 0.05543786, 0.02928152, 0.06481448, 
    0.1355146, 0.115868, 0.1120835, 0.08844705, 0.09930056, 0.07360761, 
    0.1336358, 0.1513853, 0.1232667, 0.1183333, 0.03084614, 0.08675813, 
    0.1575268, 0.100262, 0.1309424, 0.1357622,
  0.005673377, 0.0006523214, 0.05905588, 0.08482274, 0.0263191, 0.03323307, 
    0.02427896, 0.03175382, 0.0429743, 0.001907409, 0.001496649, 
    0.0009885365, 0.02885534, 0.07729732, 0.07668238, 0.06094614, 0.08619066, 
    0.09287883, 0.1597158, 0.07212679, 0.1020813, 0.02187135, 0.0195666, 
    1.405641e-07, 0.03362204, 0.06973576, 0.1118798, 0.07426371, 0.006194589,
  8.833943e-07, 0.00228351, 0.04573521, 0.01283327, 0.03027991, 0.05338135, 
    0.003707152, 0.006665844, 1.314166e-06, -4.396176e-07, 0.001824522, 
    0.001147862, 0.01289201, 0.04801792, 0.05871302, 0.05701145, 0.05970449, 
    0.06325878, 0.08081719, 0.04970079, 0.0008278809, -2.216414e-06, 
    7.206591e-08, -4.522441e-06, 0.0655624, 0.2109419, 0.08648808, 
    0.0008526891, 6.496072e-06,
  0.0031055, 0.03893925, 0.07808512, 0.0698873, 0.06541058, 0.09822825, 
    0.08491465, 0.04685856, 0.009417949, 0.003961715, 0.01139471, 0.00701731, 
    0.02842302, 0.04548808, 0.06330107, 0.06494309, 0.04082676, 0.02098357, 
    0.007570747, 0.001609353, 4.271608e-08, 7.099632e-07, 1.446481e-05, 
    0.0556039, 0.1244957, 0.147375, 0.008599504, 5.396675e-07, 1.598104e-07,
  0.1630753, 0.2807042, 0.1028103, 0.09397557, 0.02588502, 0.03549983, 
    0.02463053, 0.01186141, 0.1384714, 0.1756814, 0.04757431, 0.02774705, 
    0.02430872, 0.02312187, 0.009929959, 0.01022789, 0.003376444, 
    0.0001965457, 1.095801e-05, 5.669473e-05, 0.008743202, 0.01791624, 
    0.03123722, 0.1181643, 0.1610354, 0.02109213, 0.116485, 0.03101583, 
    0.04676546,
  0.0007986804, 0.001009002, 0.01631821, 0.1067083, 0.05610301, 0.02643004, 
    0.05102389, 0.06059658, 0.08759294, 0.08976375, 0.08412528, 0.04811238, 
    0.07849506, 0.08717808, 0.08169923, 0.05297638, 0.05565579, 0.07936568, 
    0.09626838, 0.1478332, 0.1676945, 0.04598076, 0.07662033, 0.04375483, 
    0.02947956, 0.03084994, 0.02764317, 0.001821183, 0.0006844596,
  1.152778e-05, 5.292468e-07, 0.0004255701, 0.008678375, 0.01673569, 
    0.01088739, 0.02637148, 0.01367113, 0.03681277, 0.04507606, 0.08550707, 
    0.042909, 0.02828706, 0.05926856, 0.01697679, 0.02692085, 0.04201915, 
    0.01351151, 0.01382744, 0.0008645485, 0.01623126, 0.1568111, 0.02428219, 
    0.06327158, 0.03714496, 0.0731342, 0.02421741, 0.02096852, -3.881471e-06,
  0.0008816366, 0.01033902, 0.01653278, 0.02165501, 0.0831739, 0.02669797, 
    0.03689786, 0.1513565, 0.2058364, 0.08356483, 0.01356441, 0.07760242, 
    0.0796504, 0.106272, 0.1229664, 0.07430132, 0.06409217, 0.06505676, 
    0.02833389, 0.002184371, 0.02663861, 0.05664169, 0.08504072, 0.05596696, 
    0.04875576, 0.1033279, 0.06106827, 0.0446028, 0.03500447,
  0.05134596, 0.1034828, 0.09155126, 0.1748538, 0.05057107, 0.01757751, 
    0.1168916, 0.03683108, 0.01403254, 0.01552696, 0.1108538, 0.1298784, 
    0.1462153, 0.1308274, 0.1666054, 0.1631458, 0.2130767, 0.1838006, 
    0.1098813, 0.08904499, 0.06230026, 0.02074532, 0.09814352, 0.1384204, 
    0.1834251, 0.1380423, 0.1626463, 0.1100219, 0.09360961,
  0.1943451, 0.1892082, 0.2484818, 0.1951946, 0.1621811, 0.1108809, 
    0.08475346, 0.1549174, 0.1163681, 0.1594102, 0.1378902, 0.1473307, 
    0.2303406, 0.2577822, 0.2209471, 0.1834799, 0.1890506, 0.2235293, 
    0.2307827, 0.2548966, 0.1646554, 0.1611456, 0.2563293, 0.3784133, 
    0.2206504, 0.1847004, 0.1615095, 0.2278551, 0.1828538,
  0.2603572, 0.3781346, 0.3941262, 0.3448562, 0.3528547, 0.3338577, 
    0.3057905, 0.3693998, 0.3801386, 0.3190647, 0.2780027, 0.1254395, 
    0.1847344, 0.1495769, 0.1838821, 0.2099105, 0.2210224, 0.3274524, 
    0.2783191, 0.2720454, 0.2324461, 0.3636374, 0.431587, 0.3459413, 0.35663, 
    0.4196708, 0.2556445, 0.27448, 0.2652684,
  0.2465099, 0.2928877, 0.3301105, 0.4132509, 0.5056924, 0.3912581, 0.308674, 
    0.4349634, 0.3869816, 0.2829874, 0.2181608, 0.2329938, 0.208421, 
    0.2558562, 0.3068062, 0.1747868, 0.2167766, 0.2173107, 0.2018369, 
    0.2059936, 0.152936, 0.3113091, 0.2401131, 0.2916761, 0.1482022, 
    0.285069, 0.2262097, 0.1613401, 0.1978528,
  0.1594323, 0.2114829, 0.1897825, 0.1578303, 0.1558019, 0.127169, 0.139966, 
    0.1402428, 0.1400628, 0.1648784, 0.2005018, 0.1935176, 0.2223028, 
    0.2134673, 0.2413486, 0.2314761, 0.206813, 0.2246376, 0.2868668, 
    0.3191476, 0.2381062, 0.2515149, 0.1808176, 0.08950044, 0.1140569, 
    0.09417479, 0.06608734, 0.09496796, 0.1989291,
  0.1790929, 0.1753616, 0.1716303, 0.167899, 0.1641676, 0.1604363, 0.156705, 
    0.1671094, 0.1653738, 0.1636382, 0.1619027, 0.1601671, 0.1584316, 
    0.156696, 0.1514136, 0.1590555, 0.1666974, 0.1743393, 0.1819813, 
    0.1896232, 0.1972651, 0.1968967, 0.1947216, 0.1925466, 0.1903715, 
    0.1881965, 0.1860214, 0.1838463, 0.1820779,
  0.1221126, 0.09743369, 0.05938799, 0.07570966, 0.06545101, 0.07217167, 
    0.06268746, 0.04623236, 0.04186805, 0.09859364, 0.09995405, 0.09194535, 
    0.1390046, 0.1199317, 0.04865463, 0.04060958, 0.07924919, 0.1073494, 
    0.1305343, 0.1021543, 0.2036595, 0.3766513, 0.3063813, 0.2304379, 
    0.2037442, 0.1546147, 0.1337231, 0.1609323, 0.1270361,
  0.2109683, 0.2307574, 0.1952257, 0.3077726, 0.3251687, 0.2710517, 
    0.2153344, 0.2102386, 0.2303762, 0.3030411, 0.2599767, 0.1714215, 
    0.2304468, 0.2459564, 0.2001697, 0.2411971, 0.2656338, 0.2572934, 
    0.3165833, 0.2485014, 0.2719538, 0.3465114, 0.3010481, 0.5284239, 
    0.1993705, 0.1889303, 0.2932811, 0.3447155, 0.2502925,
  0.2456813, 0.2809061, 0.2868896, 0.3499693, 0.3598433, 0.3238817, 
    0.3852033, 0.2847362, 0.2586153, 0.3161206, 0.3202784, 0.3076343, 
    0.3024808, 0.2747262, 0.293489, 0.2717988, 0.278417, 0.2749936, 
    0.2552153, 0.2924692, 0.3152948, 0.2824412, 0.2781944, 0.2879701, 
    0.1996099, 0.1705767, 0.1780314, 0.1839063, 0.2464192,
  0.1415462, 0.1854379, 0.2262974, 0.2482835, 0.1723267, 0.1446359, 
    0.1666138, 0.2002005, 0.2405212, 0.2261375, 0.2252087, 0.2122006, 
    0.1761793, 0.1823748, 0.1139489, 0.135952, 0.1607629, 0.1669649, 
    0.1606033, 0.1518806, 0.1684452, 0.1879205, 0.2164277, 0.1580801, 
    0.1125582, 0.1577708, 0.1397686, 0.1457667, 0.1397065,
  0.1258848, 0.09839451, 0.08853806, 0.1422153, 0.1417886, 0.1153111, 
    0.1483103, 0.1103133, 0.114878, 0.06337652, 0.05699682, 0.03811447, 
    0.07024599, 0.1506732, 0.1405341, 0.1128184, 0.1205023, 0.1081935, 
    0.08358912, 0.1371504, 0.1529044, 0.1349344, 0.1385957, 0.03977152, 
    0.07185369, 0.1516818, 0.1058528, 0.1412598, 0.1598478,
  0.006098142, 0.001166914, 0.03717886, 0.05365229, 0.03298236, 0.03438231, 
    0.02838344, 0.03235115, 0.04813316, 0.001246152, 0.0002182126, 
    0.002024114, 0.02545135, 0.06925599, 0.0854586, 0.06454931, 0.08777692, 
    0.0895862, 0.1459291, 0.06720591, 0.1006684, 0.03315975, 0.01607107, 
    4.639052e-07, 0.02994547, 0.05800751, 0.1009941, 0.07338312, 0.0168955,
  4.032958e-07, 0.0009612183, 0.0259275, 0.01066154, 0.03248772, 0.0597648, 
    0.01122968, 0.01230733, -1.90184e-05, 2.042564e-07, 0.000858454, 
    0.0001669677, 0.01373111, 0.05560688, 0.06147425, 0.05453169, 0.06023789, 
    0.06424491, 0.07692115, 0.06488175, 0.005276927, -7.943154e-07, 
    3.025112e-08, -3.70365e-06, 0.05705946, 0.2010315, 0.08838098, 
    0.004168362, 0.0002867298,
  0.002499519, 0.03534898, 0.06374114, 0.07688276, 0.07177636, 0.08995953, 
    0.08978737, 0.05805724, 0.0145194, 0.003979632, 0.004765767, 0.006122324, 
    0.03145882, 0.04186386, 0.05839778, 0.05922838, 0.04342145, 0.03687575, 
    0.02179366, 0.003890443, -2.668066e-06, 1.506163e-07, 6.149889e-06, 
    0.04731396, 0.1085974, 0.1041965, 0.01099587, 2.264877e-06, 3.250601e-07,
  0.1203085, 0.2364849, 0.09187099, 0.1235299, 0.02466208, 0.03454073, 
    0.02673801, 0.01306334, 0.1440623, 0.1793579, 0.03749559, 0.02588094, 
    0.02276085, 0.02255129, 0.0107391, 0.01239888, 0.003625988, 0.0002086828, 
    0.001358753, 0.0007930789, 0.01530156, 0.02291108, 0.02322911, 0.1024238, 
    0.1504255, 0.01617987, 0.1216685, 0.05244591, 0.06355805,
  0.0002641383, 0.0004436584, 0.002788684, 0.0987938, 0.06476428, 0.0301856, 
    0.05859999, 0.06734973, 0.09821154, 0.08515906, 0.08946031, 0.04601561, 
    0.07325079, 0.08490536, 0.07890174, 0.05571139, 0.05595212, 0.08335053, 
    0.1001565, 0.1593167, 0.1626243, 0.04876014, 0.09726955, 0.04963215, 
    0.03198096, 0.03143021, 0.02546689, 0.0006695124, 0.0004016203,
  7.659358e-06, 2.970179e-07, 0.009136692, 0.009756216, 0.01673446, 
    0.01152488, 0.03811278, 0.01794533, 0.03701875, 0.05103267, 0.07579726, 
    0.0492432, 0.0345416, 0.06167987, 0.02429821, 0.02625365, 0.04526891, 
    0.01830606, 0.01686517, 0.01010303, 0.01646293, 0.1754987, 0.03134583, 
    0.06274433, 0.04526871, 0.07338981, 0.02794465, 0.008845931, 5.75487e-06,
  0.001152488, 0.01493908, 0.01872139, 0.02651297, 0.08489749, 0.02502692, 
    0.0186385, 0.1299517, 0.1717869, 0.08230965, 0.02571047, 0.07978472, 
    0.07959947, 0.108648, 0.1308661, 0.08563913, 0.07633006, 0.07412897, 
    0.03392789, 0.003192931, 0.01985479, 0.05015626, 0.0956829, 0.05442453, 
    0.05716732, 0.1095164, 0.06273174, 0.05125163, 0.02499378,
  0.04714888, 0.1125487, 0.1015446, 0.1638516, 0.04954229, 0.02298243, 
    0.1178486, 0.02740441, 0.008532003, 0.0176595, 0.1123177, 0.1454147, 
    0.1613938, 0.1457291, 0.1893739, 0.1684315, 0.2302972, 0.1996434, 
    0.1173996, 0.1020596, 0.06159943, 0.01700403, 0.09939419, 0.1372306, 
    0.1922906, 0.1366282, 0.1750665, 0.1208816, 0.1088234,
  0.2093494, 0.2080143, 0.2692688, 0.2109187, 0.169264, 0.1177016, 
    0.08502899, 0.1700003, 0.1030602, 0.1623928, 0.1434749, 0.1562068, 
    0.2528274, 0.2925608, 0.2270187, 0.2045057, 0.2125346, 0.242315, 
    0.2333415, 0.2707043, 0.1348155, 0.1634312, 0.2796496, 0.3769462, 
    0.2275102, 0.2040635, 0.1767035, 0.250926, 0.1952603,
  0.2539347, 0.378974, 0.3521209, 0.4035739, 0.3544089, 0.3036631, 0.2818704, 
    0.365018, 0.370219, 0.3663478, 0.3264821, 0.1197845, 0.1921697, 
    0.1306239, 0.2000935, 0.2577794, 0.2007684, 0.3234712, 0.266864, 
    0.2514971, 0.2147964, 0.3370214, 0.4207419, 0.3377286, 0.3588181, 
    0.4117206, 0.2880067, 0.2762226, 0.2692261,
  0.2679441, 0.2780165, 0.3033708, 0.4102083, 0.5147189, 0.3722929, 
    0.3274135, 0.4531306, 0.3816045, 0.2788796, 0.2293718, 0.2176625, 
    0.1951192, 0.2458549, 0.2926185, 0.1730569, 0.1951254, 0.2287476, 
    0.2015612, 0.1905108, 0.1434638, 0.2465175, 0.2200464, 0.264966, 
    0.1616607, 0.3246517, 0.2245678, 0.1829068, 0.2061174,
  0.1958522, 0.1999094, 0.1848658, 0.1448812, 0.148247, 0.1402744, 0.1324417, 
    0.1378879, 0.1542718, 0.1922881, 0.2134315, 0.230848, 0.2329534, 
    0.1861328, 0.2217217, 0.1897443, 0.1874892, 0.2149992, 0.2347701, 
    0.2723571, 0.2271817, 0.2337769, 0.1692068, 0.1071295, 0.1282315, 
    0.1094766, 0.069879, 0.1102076, 0.2113817,
  0.2035707, 0.2016974, 0.1998241, 0.1979507, 0.1960773, 0.194204, 0.1923307, 
    0.2001759, 0.1989935, 0.197811, 0.1966285, 0.1954461, 0.1942636, 
    0.1930811, 0.1921096, 0.1991467, 0.2061839, 0.213221, 0.2202581, 
    0.2272953, 0.2343324, 0.2194073, 0.215426, 0.2114447, 0.2074634, 
    0.203482, 0.1995007, 0.1955194, 0.2050694,
  0.1253891, 0.1195525, 0.08599807, 0.07734853, 0.07055968, 0.09122869, 
    0.07390572, 0.05360465, 0.08006046, 0.127666, 0.1099074, 0.107674, 
    0.14666, 0.1017025, 0.03891945, 0.03900864, 0.08117791, 0.08899741, 
    0.1310972, 0.09778561, 0.2084182, 0.3781064, 0.3235139, 0.2039858, 
    0.1746408, 0.1625134, 0.0958057, 0.1473797, 0.1280805,
  0.2215768, 0.2517751, 0.2219599, 0.2952597, 0.3347203, 0.3040879, 
    0.2252911, 0.204673, 0.2398595, 0.3099995, 0.2572181, 0.1655934, 
    0.2236224, 0.2276334, 0.1937425, 0.2117264, 0.2458667, 0.2318806, 
    0.2882767, 0.2566805, 0.2695795, 0.3524703, 0.3108101, 0.5115632, 
    0.1697624, 0.1822456, 0.3059429, 0.3248594, 0.2916984,
  0.2669996, 0.2775259, 0.3029056, 0.3240711, 0.3714353, 0.3657446, 0.348285, 
    0.2925108, 0.2567778, 0.2940599, 0.3232856, 0.2961457, 0.268317, 
    0.2640162, 0.2989709, 0.2743815, 0.27551, 0.2636248, 0.2609663, 
    0.2910362, 0.3155966, 0.280281, 0.2711148, 0.2855647, 0.1967634, 
    0.193103, 0.2116046, 0.1958116, 0.2334155,
  0.1602936, 0.203152, 0.2293076, 0.2478069, 0.1766748, 0.152115, 0.1784491, 
    0.2215909, 0.2728786, 0.245277, 0.2572014, 0.2199951, 0.1946819, 
    0.1838444, 0.1092055, 0.1393383, 0.1685937, 0.1772242, 0.1751657, 
    0.1793773, 0.1923165, 0.2265498, 0.2201251, 0.1640275, 0.08518057, 
    0.1545928, 0.1537578, 0.1480919, 0.1531966,
  0.1235546, 0.1141837, 0.1202844, 0.1554081, 0.1416726, 0.1482087, 
    0.1722622, 0.1402878, 0.1345165, 0.05877278, 0.05467007, 0.04941733, 
    0.07051519, 0.1583361, 0.1594962, 0.1244304, 0.1303965, 0.1278053, 
    0.1135027, 0.1259913, 0.1499711, 0.1472675, 0.1508646, 0.04760048, 
    0.05478986, 0.1513446, 0.1172535, 0.1498986, 0.1526375,
  0.0130457, 0.003064678, 0.02838852, 0.04204328, 0.05511867, 0.04641896, 
    0.0365291, 0.04003824, 0.05161182, 0.003319571, 8.075163e-05, 
    0.002006636, 0.01790133, 0.06787995, 0.08494588, 0.05555907, 0.09164865, 
    0.08668237, 0.1396078, 0.07979068, 0.1001918, 0.05763081, 0.01406479, 
    3.759523e-07, 0.02448701, 0.05107963, 0.09685767, 0.08032583, 0.03736449,
  -9.209087e-06, 0.000206031, 0.02127932, 0.007442337, 0.03738736, 
    0.06746447, 0.01693991, 0.02654238, 0.0007666473, 1.472846e-07, 
    0.0004197787, 4.304926e-05, 0.01174647, 0.04538439, 0.06439938, 
    0.05187561, 0.05759839, 0.06370784, 0.06999466, 0.08155654, 0.0382406, 
    0.001964636, 1.886431e-07, 5.825529e-06, 0.05548763, 0.1870147, 
    0.08205655, 0.02804965, 0.002088572,
  0.000398487, 0.03074501, 0.05994788, 0.08564685, 0.07889234, 0.08546872, 
    0.08488442, 0.06852684, 0.01682414, 0.003806665, 0.003886535, 0.00583102, 
    0.03437715, 0.03442208, 0.05216673, 0.04768311, 0.04159311, 0.0341044, 
    0.03448393, 0.02746648, 0.0002605787, 3.723766e-07, 3.222979e-06, 
    0.04226515, 0.09755638, 0.0758674, 0.02654965, 4.792369e-05, 1.224402e-06,
  0.1057492, 0.2135864, 0.08738635, 0.1608171, 0.02736049, 0.04113936, 
    0.02683783, 0.01382225, 0.1467578, 0.1853557, 0.02993983, 0.0182536, 
    0.0200861, 0.02171558, 0.01200641, 0.01515726, 0.003479171, 0.001414454, 
    0.002083234, 0.01141698, 0.01699999, 0.01645727, 0.0184916, 0.08944695, 
    0.1205673, 0.01280483, 0.1206128, 0.08187983, 0.07271546,
  9.653719e-05, 2.269107e-05, 0.001448676, 0.0815176, 0.07618531, 0.02901174, 
    0.06733272, 0.06676725, 0.08781622, 0.07847334, 0.08654365, 0.03863845, 
    0.06384124, 0.07521167, 0.0754162, 0.05304452, 0.05788893, 0.08112351, 
    0.1080691, 0.1584072, 0.1550541, 0.04555002, 0.1153391, 0.05175314, 
    0.03134751, 0.03310476, 0.025564, 0.0008095592, 3.811172e-05,
  2.895659e-06, 1.282836e-07, 0.00594318, 0.01115656, 0.01160587, 0.01695546, 
    0.03200628, 0.01803069, 0.06356916, 0.06310654, 0.07301329, 0.05323578, 
    0.04496387, 0.06362255, 0.03531912, 0.03601143, 0.06566414, 0.02633351, 
    0.01916496, 0.02220159, 0.0152525, 0.2034987, 0.04099793, 0.06453586, 
    0.04425735, 0.06131129, 0.0286818, 0.006019951, 5.586847e-06,
  0.002135214, 0.03114298, 0.01830227, 0.02673479, 0.07885026, 0.02964038, 
    0.006491075, 0.09574091, 0.1482903, 0.06268592, 0.05793121, 0.09217186, 
    0.09385031, 0.1040533, 0.1357856, 0.09558395, 0.09864336, 0.08211885, 
    0.02454466, 0.003646243, 0.01274295, 0.03624957, 0.0847214, 0.06370737, 
    0.07070336, 0.101766, 0.05531099, 0.06498785, 0.016351,
  0.04132219, 0.1182709, 0.1111521, 0.1669166, 0.04073868, 0.0316114, 
    0.1120381, 0.01866965, 0.006107855, 0.02866863, 0.1138037, 0.1814692, 
    0.1827244, 0.1849176, 0.2163555, 0.1785533, 0.240407, 0.2055299, 
    0.1270504, 0.101676, 0.05391242, 0.01738456, 0.09968854, 0.1285334, 
    0.2105417, 0.1274076, 0.1708199, 0.1412431, 0.1215669,
  0.2186475, 0.2095887, 0.2587531, 0.2317871, 0.1682817, 0.1122124, 
    0.09395553, 0.1834478, 0.09249068, 0.1658612, 0.1542101, 0.1741525, 
    0.2816445, 0.3371624, 0.2544574, 0.233373, 0.2142722, 0.2550266, 
    0.2439281, 0.2955583, 0.1278247, 0.1716863, 0.2786876, 0.3538327, 
    0.2389748, 0.21304, 0.1910847, 0.2603682, 0.2101368,
  0.2581384, 0.3629743, 0.3360915, 0.4136834, 0.2876674, 0.2940258, 
    0.2460276, 0.3272542, 0.3791858, 0.395067, 0.3508818, 0.1290204, 
    0.202369, 0.1608943, 0.2352951, 0.2746785, 0.2204379, 0.3273968, 
    0.2583217, 0.2496006, 0.2469373, 0.3394361, 0.4462295, 0.3679068, 
    0.3715501, 0.374837, 0.2949178, 0.2907816, 0.290673,
  0.25565, 0.2909756, 0.3245703, 0.3980098, 0.4710447, 0.378824, 0.3044856, 
    0.417021, 0.3636497, 0.3260459, 0.2515257, 0.2172989, 0.1841635, 
    0.2840027, 0.2833393, 0.161548, 0.1859445, 0.2424168, 0.1758755, 
    0.2410106, 0.1842354, 0.2278683, 0.2555838, 0.2376566, 0.1511215, 
    0.3439026, 0.2433864, 0.2021924, 0.2359022,
  0.2280626, 0.1889092, 0.1894425, 0.1472175, 0.1414365, 0.1602477, 
    0.1338449, 0.1431052, 0.1777455, 0.2047913, 0.2022339, 0.2128564, 
    0.2200877, 0.1848896, 0.1923966, 0.1773659, 0.1729397, 0.1920487, 
    0.2549151, 0.318606, 0.2548181, 0.1942986, 0.1278995, 0.1204305, 
    0.1440974, 0.1315666, 0.05740439, 0.1355885, 0.2520228,
  0.2238133, 0.2214547, 0.219096, 0.2167373, 0.2143787, 0.21202, 0.2096614, 
    0.2073528, 0.207474, 0.2075952, 0.2077164, 0.2078376, 0.2079588, 0.20808, 
    0.2166639, 0.2224937, 0.2283235, 0.2341533, 0.2399831, 0.2458129, 
    0.2516427, 0.2409128, 0.2373204, 0.2337281, 0.2301357, 0.2265434, 
    0.222951, 0.2193587, 0.2257002,
  0.1333709, 0.1305471, 0.1141588, 0.1181752, 0.09293275, 0.1299541, 
    0.1187031, 0.06781124, 0.1210369, 0.1468144, 0.1214715, 0.1114799, 
    0.1616359, 0.1034686, 0.09741025, 0.0895419, 0.08382792, 0.07547863, 
    0.1110464, 0.09054604, 0.2335229, 0.3974927, 0.3596885, 0.1853035, 
    0.1851183, 0.1415076, 0.1249541, 0.1277325, 0.1340293,
  0.2244355, 0.2587568, 0.2169385, 0.2514784, 0.3260345, 0.3279405, 0.220403, 
    0.195232, 0.2466473, 0.3114589, 0.2592307, 0.147082, 0.2020969, 
    0.2282642, 0.2434711, 0.2070744, 0.2509333, 0.2429199, 0.2689621, 
    0.2643933, 0.3038192, 0.3613084, 0.3305972, 0.5230316, 0.1545229, 
    0.2292667, 0.3369372, 0.3079701, 0.2866993,
  0.2884834, 0.2978873, 0.3383538, 0.3709821, 0.3605033, 0.3335303, 
    0.4155833, 0.3066777, 0.3254668, 0.3384503, 0.3345253, 0.2765126, 
    0.2944898, 0.3004647, 0.3001776, 0.2827783, 0.2872086, 0.3009153, 
    0.2844909, 0.3392196, 0.3310217, 0.3078655, 0.2836134, 0.2998613, 
    0.1837623, 0.2001219, 0.2290324, 0.2587638, 0.2814821,
  0.1884062, 0.2404705, 0.2434906, 0.2597373, 0.2070293, 0.1852742, 
    0.2200087, 0.2846922, 0.2880332, 0.2492697, 0.3096795, 0.2547567, 
    0.2370892, 0.1837846, 0.1075456, 0.1679381, 0.1967161, 0.2103568, 
    0.2048643, 0.205601, 0.2140447, 0.2412803, 0.2480243, 0.1795498, 
    0.06823877, 0.1588655, 0.1653158, 0.1632603, 0.1766625,
  0.1686746, 0.171858, 0.150771, 0.1767045, 0.1677284, 0.1999654, 0.201247, 
    0.1802696, 0.1657283, 0.09264391, 0.0697352, 0.06728371, 0.07641992, 
    0.1602392, 0.1845093, 0.1349427, 0.1737617, 0.1557153, 0.1461386, 
    0.1347469, 0.190116, 0.1778048, 0.1812003, 0.05449729, 0.05376971, 
    0.1773717, 0.1296467, 0.1729798, 0.1522813,
  0.04246613, 0.01577681, 0.0283097, 0.06031064, 0.07562077, 0.06319474, 
    0.04267409, 0.06273974, 0.06037851, 0.007126577, 6.283639e-05, 
    0.0002546838, 0.02901243, 0.07060329, 0.09751809, 0.06696501, 0.09920292, 
    0.09939441, 0.1426386, 0.09209457, 0.1052107, 0.08699502, 0.02165511, 
    5.52736e-07, 0.01420525, 0.06041297, 0.1076123, 0.09762671, 0.06415592,
  0.0007452663, 2.962294e-05, 0.01796935, 0.006250432, 0.04314692, 
    0.06087417, 0.03317231, 0.04315197, 0.004492331, 1.042157e-07, 
    0.0001269696, 7.169901e-06, 0.0151905, 0.0363111, 0.06872642, 0.05477259, 
    0.03916213, 0.0604139, 0.05891946, 0.08933808, 0.07099885, 0.02125319, 
    2.358307e-06, 2.944847e-05, 0.06967053, 0.186589, 0.07771935, 0.09676678, 
    0.02523579,
  2.881132e-05, 0.02103969, 0.05724724, 0.09066702, 0.07343444, 0.0823618, 
    0.07562857, 0.07187938, 0.02082175, 0.005686848, 0.004242225, 
    0.006437711, 0.04048181, 0.03265007, 0.04590043, 0.04106176, 0.03619647, 
    0.0309606, 0.03250588, 0.0462229, 0.009565827, 0.0001433218, 
    2.544196e-06, 0.03918894, 0.08820307, 0.06326339, 0.04657881, 
    0.003459402, 3.949067e-05,
  0.09945771, 0.193679, 0.08297411, 0.1841419, 0.02758832, 0.04034486, 
    0.0249977, 0.01374366, 0.1458742, 0.1993016, 0.02799934, 0.01610134, 
    0.02014701, 0.02107863, 0.01340059, 0.01768039, 0.005916457, 0.002519531, 
    0.001822531, 0.00592088, 0.01047239, 0.006888435, 0.01911976, 0.07555471, 
    0.09015752, 0.01443821, 0.1125752, 0.08019369, 0.07635547,
  3.449933e-05, 4.619618e-06, 0.0002709697, 0.06505211, 0.08712347, 
    0.0284121, 0.07258362, 0.05862703, 0.07984932, 0.07192125, 0.07476741, 
    0.03289685, 0.05317308, 0.06300264, 0.06586585, 0.049346, 0.06730004, 
    0.07691996, 0.114105, 0.1412975, 0.1402393, 0.04103466, 0.1089726, 
    0.05992409, 0.03092317, 0.03309274, 0.02400513, 0.0007630747, 0.0001119051,
  9.940652e-07, 3.853068e-08, 3.795898e-05, 0.02153982, 0.007263305, 
    0.04177663, 0.03032082, 0.01725429, 0.08965321, 0.07292084, 0.1025761, 
    0.06359418, 0.052538, 0.06823575, 0.04456959, 0.06563775, 0.06766276, 
    0.03745454, 0.03365363, 0.01679279, 0.01621708, 0.2306145, 0.05678774, 
    0.06949525, 0.04101631, 0.04537663, 0.02887512, 0.001644114, 2.711024e-06,
  8.681523e-05, 0.03338492, 0.03171931, 0.03319481, 0.07919046, 0.02753014, 
    0.002930928, 0.06621791, 0.146506, 0.03816584, 0.1297542, 0.1434929, 
    0.1237965, 0.1231456, 0.164548, 0.1401537, 0.1277882, 0.09005949, 
    0.04444206, 0.003694917, 0.01038991, 0.04431523, 0.08081906, 0.07292423, 
    0.08932448, 0.0944725, 0.05025944, 0.07850185, 0.01341804,
  0.03290758, 0.1299018, 0.1213482, 0.1628089, 0.03712923, 0.01336829, 
    0.1100203, 0.0145965, 0.002938477, 0.02712836, 0.1139955, 0.2224682, 
    0.234434, 0.2196881, 0.2571262, 0.2011329, 0.2681734, 0.2339235, 
    0.1337115, 0.1048746, 0.04832037, 0.02281262, 0.109921, 0.1457106, 
    0.2472322, 0.155183, 0.1923213, 0.1730043, 0.1377635,
  0.2276818, 0.2315944, 0.279707, 0.2686772, 0.1552095, 0.09696927, 
    0.08980056, 0.1934029, 0.08790653, 0.1812108, 0.1855106, 0.191121, 
    0.3294788, 0.3653165, 0.289069, 0.2720705, 0.2750994, 0.3069095, 
    0.2932566, 0.3173888, 0.1444619, 0.2128839, 0.3070847, 0.3652742, 
    0.270674, 0.2501588, 0.2256767, 0.2917376, 0.2153114,
  0.2572375, 0.3709412, 0.3425975, 0.4094372, 0.2970487, 0.2533973, 
    0.2788366, 0.3910496, 0.4139235, 0.4366287, 0.3940266, 0.1538266, 
    0.1886588, 0.2126945, 0.3152542, 0.3026349, 0.2441783, 0.3327451, 
    0.2700201, 0.2833082, 0.2864574, 0.3338152, 0.4726422, 0.3422585, 
    0.4267765, 0.3375165, 0.2974004, 0.2977858, 0.29541,
  0.2386622, 0.2640558, 0.3406761, 0.4120677, 0.4648764, 0.3773323, 
    0.3164041, 0.411883, 0.3620265, 0.3428182, 0.2706226, 0.2295374, 
    0.2120275, 0.3114319, 0.2967823, 0.1648524, 0.2270819, 0.2830985, 
    0.1614985, 0.284118, 0.2336984, 0.2309681, 0.2170042, 0.2319386, 
    0.1466516, 0.3430409, 0.2257205, 0.2169704, 0.286734,
  0.228348, 0.1963353, 0.1823034, 0.1707732, 0.1370191, 0.1539414, 0.1204397, 
    0.1388953, 0.1839736, 0.2146413, 0.2413753, 0.2123234, 0.2437037, 
    0.195654, 0.2090714, 0.1957101, 0.2265965, 0.2262706, 0.281152, 
    0.3293548, 0.217446, 0.2212054, 0.1103237, 0.1555264, 0.1730231, 
    0.1683882, 0.06162887, 0.1602474, 0.2943027,
  0.239329, 0.2373471, 0.2353651, 0.2333831, 0.2314012, 0.2294192, 0.2274373, 
    0.2369586, 0.2376538, 0.238349, 0.2390442, 0.2397394, 0.2404347, 
    0.2411299, 0.2423108, 0.2480323, 0.2537538, 0.2594754, 0.2651969, 
    0.2709184, 0.2766399, 0.2614665, 0.2570317, 0.2525969, 0.2481622, 
    0.2437274, 0.2392926, 0.2348579, 0.2409146,
  0.1420546, 0.14006, 0.1425999, 0.1357504, 0.1191852, 0.1709619, 0.1600291, 
    0.09672549, 0.1396873, 0.1539332, 0.1178827, 0.1149914, 0.1799656, 
    0.08417568, 0.1253543, 0.1858236, 0.1336689, 0.1063605, 0.09029976, 
    0.08762123, 0.2581331, 0.4035068, 0.4118643, 0.269693, 0.1884749, 
    0.1597546, 0.1215621, 0.1046852, 0.1410816,
  0.2669128, 0.2496384, 0.2246366, 0.2139201, 0.307771, 0.3385029, 0.1863074, 
    0.2038464, 0.2512836, 0.3139808, 0.2544441, 0.1337214, 0.1932678, 
    0.2245486, 0.269699, 0.2717497, 0.2910791, 0.2491829, 0.3150767, 
    0.2672046, 0.3012953, 0.3648446, 0.3332968, 0.5440735, 0.1461944, 
    0.2308441, 0.4052878, 0.3725891, 0.3095086,
  0.3632731, 0.3489857, 0.3732746, 0.4127621, 0.4290323, 0.3768985, 
    0.4713707, 0.3630701, 0.4081026, 0.3526006, 0.3504045, 0.360032, 
    0.3812475, 0.3702627, 0.3233463, 0.3249543, 0.3281333, 0.3366174, 
    0.2870841, 0.3611589, 0.3353969, 0.3322993, 0.3023583, 0.3160929, 
    0.2110581, 0.243952, 0.2701821, 0.2688804, 0.319309,
  0.2558888, 0.307722, 0.3065382, 0.3167059, 0.2673039, 0.2310321, 0.2967828, 
    0.36349, 0.3333681, 0.3285401, 0.3287694, 0.2808248, 0.26422, 0.2388674, 
    0.1407155, 0.2154533, 0.2852352, 0.2207897, 0.229701, 0.2649859, 
    0.2693786, 0.292094, 0.2872443, 0.1720475, 0.05690904, 0.1656123, 
    0.1901855, 0.176249, 0.2412922,
  0.2441754, 0.2262786, 0.196641, 0.2112844, 0.2299103, 0.2080821, 0.235448, 
    0.2203477, 0.2234447, 0.1618069, 0.1008234, 0.12048, 0.08890584, 
    0.1786966, 0.1994644, 0.1651745, 0.2344362, 0.2094948, 0.190321, 
    0.177686, 0.2595281, 0.2437323, 0.2472025, 0.06205673, 0.04422725, 
    0.2132273, 0.1658924, 0.2128046, 0.2249217,
  0.07625458, 0.03959407, 0.02800539, 0.08020316, 0.1306413, 0.1445141, 
    0.1017328, 0.1120331, 0.09328949, 0.01854679, -2.356899e-05, 
    6.737045e-05, 0.03438899, 0.09115652, 0.1079087, 0.07806389, 0.1139408, 
    0.1195467, 0.1484417, 0.131463, 0.1271748, 0.1272926, 0.07435949, 
    1.316519e-06, 0.008985294, 0.06980111, 0.1161852, 0.1255962, 0.121873,
  0.04311868, -3.581615e-05, 0.01299539, 0.00881446, 0.04173779, 0.06229334, 
    0.05820099, 0.0591699, 0.01303076, 6.684371e-08, 5.653533e-05, 
    -5.969613e-07, 0.0187127, 0.03923241, 0.06481299, 0.05079937, 0.0445303, 
    0.06157039, 0.0522519, 0.07659046, 0.1582944, 0.1282123, 0.0005108092, 
    5.548797e-05, 0.06955485, 0.2106875, 0.06875579, 0.1463787, 0.2335135,
  0.0004797834, 0.01881657, 0.04779168, 0.0991068, 0.0643099, 0.07874869, 
    0.06468161, 0.06096171, 0.02872273, 0.007685019, 0.006191002, 0.00888612, 
    0.04180893, 0.03239259, 0.04081399, 0.04455924, 0.03491188, 0.03196611, 
    0.03165832, 0.04274526, 0.07421142, 0.005272981, 9.894566e-05, 
    0.03591655, 0.07675716, 0.04732145, 0.05855179, 0.03943397, 0.00544444,
  0.09457765, 0.17734, 0.07744807, 0.1890703, 0.02775865, 0.03742376, 
    0.02554791, 0.01624438, 0.156196, 0.209557, 0.02883969, 0.0179598, 
    0.02452528, 0.02153521, 0.01666107, 0.02160366, 0.009609513, 0.005069519, 
    0.008773934, 0.003649584, 0.01157437, 0.00219409, 0.01341348, 0.06836397, 
    0.06776686, 0.02156887, 0.09553462, 0.07584652, 0.08782781,
  2.238336e-05, 1.694263e-06, 8.136805e-05, 0.04009297, 0.08195712, 
    0.02717401, 0.05979763, 0.05407238, 0.09092861, 0.07219446, 0.06697185, 
    0.03201315, 0.04456744, 0.05431491, 0.05734454, 0.0446042, 0.06939091, 
    0.07509778, 0.1148184, 0.1217328, 0.1268632, 0.0430627, 0.106268, 
    0.06561101, 0.03428226, 0.03531685, 0.03119769, 0.000821342, 3.726432e-05,
  3.430933e-07, 1.170476e-08, 4.388902e-06, 0.03476328, 0.001833473, 
    0.05905111, 0.02985791, 0.02774943, 0.1057233, 0.1208579, 0.147971, 
    0.0890801, 0.0596393, 0.06700068, 0.06222942, 0.0668842, 0.07920171, 
    0.06169474, 0.06818993, 0.04028083, 0.01863958, 0.2508729, 0.07143422, 
    0.0729294, 0.0405279, 0.04345256, 0.04277287, 0.01423549, 1.349995e-06,
  3.771202e-06, 0.02579622, 0.0318124, 0.03225253, 0.07975871, 0.02308237, 
    0.0008095844, 0.04364927, 0.1450246, 0.02735632, 0.219537, 0.1837606, 
    0.1673584, 0.1509399, 0.1776224, 0.1629378, 0.145101, 0.108564, 
    0.1074337, 0.02010662, 0.0111556, 0.05180506, 0.0929049, 0.1469662, 
    0.1115531, 0.1027995, 0.05346248, 0.1153909, 0.01879235,
  0.01993836, 0.1044442, 0.125401, 0.1611856, 0.0435745, 0.03150413, 
    0.09213162, 0.008432483, 0.001163157, 0.02454871, 0.1115491, 0.3363654, 
    0.2884754, 0.2559219, 0.2438109, 0.2105706, 0.2998545, 0.2363659, 
    0.1722144, 0.1148754, 0.04287231, 0.03841573, 0.1519012, 0.1671735, 
    0.2803207, 0.1851719, 0.220598, 0.2016869, 0.1683214,
  0.2341251, 0.2716939, 0.3201029, 0.2898895, 0.1506219, 0.1158648, 
    0.1158436, 0.2033772, 0.0903413, 0.2224131, 0.1789956, 0.1928126, 
    0.3873037, 0.3951775, 0.2632058, 0.2971169, 0.289906, 0.3525972, 
    0.3489125, 0.3279201, 0.1466914, 0.2542809, 0.3453099, 0.3993383, 
    0.2878348, 0.2898281, 0.2712459, 0.2946925, 0.2201028,
  0.250798, 0.3791338, 0.3691275, 0.4505312, 0.3622067, 0.2628447, 0.3286009, 
    0.4251547, 0.4475321, 0.470128, 0.4365506, 0.1902875, 0.1870849, 
    0.2346433, 0.4268, 0.3482447, 0.2758645, 0.3397869, 0.300455, 0.3160192, 
    0.3251058, 0.3597458, 0.5508322, 0.3751493, 0.435422, 0.3089865, 
    0.3126963, 0.3319702, 0.2928538,
  0.2449176, 0.2510963, 0.3364673, 0.4215121, 0.4795879, 0.393682, 0.3423777, 
    0.4290525, 0.3912379, 0.3879298, 0.313065, 0.2531811, 0.2135776, 
    0.3362046, 0.3306037, 0.1736404, 0.25468, 0.3127859, 0.1631223, 
    0.3283723, 0.2651052, 0.2407029, 0.2552967, 0.2819379, 0.1795436, 
    0.338003, 0.2342989, 0.2631522, 0.3331926,
  0.2090392, 0.2178873, 0.2115133, 0.1514233, 0.1349937, 0.178034, 0.160007, 
    0.1561715, 0.1933076, 0.2431146, 0.2800376, 0.22973, 0.2363276, 
    0.2535316, 0.2705754, 0.2523108, 0.2664974, 0.2951995, 0.3419784, 
    0.2941284, 0.2205505, 0.2109893, 0.1336039, 0.1511078, 0.1974143, 
    0.2013996, 0.06524002, 0.1916288, 0.2903086,
  0.2555861, 0.2545555, 0.2535249, 0.2524943, 0.2514637, 0.2504331, 
    0.2494026, 0.2584325, 0.2594099, 0.2603872, 0.2613645, 0.2623418, 
    0.2633191, 0.2642965, 0.2869905, 0.2929273, 0.2988641, 0.3048009, 
    0.3107377, 0.3166746, 0.3226114, 0.289979, 0.2840955, 0.278212, 
    0.2723284, 0.2664448, 0.2605613, 0.2546777, 0.2564105,
  0.1483276, 0.1527277, 0.1534702, 0.154526, 0.1447712, 0.2019109, 0.1906839, 
    0.1206931, 0.1530938, 0.1739904, 0.1401478, 0.1279005, 0.1856014, 
    0.04990642, 0.1175656, 0.1459466, 0.1299887, 0.09132442, 0.06578198, 
    0.07468365, 0.2814082, 0.4104736, 0.4162142, 0.2404297, 0.2147155, 
    0.1926508, 0.1179351, 0.09124774, 0.1363916,
  0.2589787, 0.2325573, 0.2061357, 0.1710739, 0.2748051, 0.3464334, 
    0.1524111, 0.2136372, 0.2714017, 0.3147526, 0.2463516, 0.1237627, 
    0.1916958, 0.2041444, 0.2668033, 0.2930086, 0.3302949, 0.3115808, 
    0.3818634, 0.2854013, 0.3464882, 0.3978971, 0.3595379, 0.5872952, 
    0.1363161, 0.258645, 0.4132046, 0.4051434, 0.3519582,
  0.4537735, 0.4014385, 0.3973296, 0.4148617, 0.4973191, 0.4384506, 
    0.4402761, 0.4185801, 0.4027483, 0.3663853, 0.3495806, 0.3999393, 
    0.350756, 0.3520525, 0.3284367, 0.3757995, 0.3795357, 0.4005717, 
    0.3292909, 0.3547746, 0.3631938, 0.3491749, 0.3020909, 0.3176906, 
    0.2538289, 0.2755944, 0.3460038, 0.3138597, 0.3583883,
  0.3485909, 0.342851, 0.3664609, 0.3154913, 0.2900119, 0.2944045, 0.3444951, 
    0.3859888, 0.3589789, 0.3539317, 0.3021089, 0.2742324, 0.2504224, 
    0.3038512, 0.2025051, 0.2399459, 0.3123575, 0.2535269, 0.2507197, 
    0.2935563, 0.3359863, 0.3500246, 0.3163974, 0.1687073, 0.04771744, 
    0.1980124, 0.2440161, 0.2827936, 0.2925746,
  0.2947438, 0.2768446, 0.1809198, 0.2166716, 0.2627077, 0.2843489, 
    0.3166902, 0.3036895, 0.277412, 0.2298325, 0.1717499, 0.1272142, 
    0.09375501, 0.190746, 0.2312936, 0.2411195, 0.2592141, 0.2878914, 
    0.245225, 0.2874795, 0.3038668, 0.3135437, 0.2902526, 0.06954566, 
    0.04615383, 0.2488407, 0.1984582, 0.2555913, 0.311877,
  0.1757177, 0.08395839, 0.02795581, 0.1172951, 0.1294031, 0.1632147, 
    0.1814405, 0.1643774, 0.1818996, 0.03304117, -4.629871e-05, 2.225408e-05, 
    0.0165229, 0.1351541, 0.1507828, 0.112239, 0.1333541, 0.1903853, 
    0.1930863, 0.2015772, 0.1814312, 0.1528646, 0.2317695, 1.155291e-05, 
    0.008345695, 0.1233186, 0.142194, 0.1889223, 0.1854544,
  0.2950794, -0.0001473831, 0.01053463, 0.02601278, 0.05840949, 0.0692879, 
    0.07747933, 0.09072073, 0.08619319, 6.433789e-08, 2.37885e-05, 
    -4.176798e-07, 0.05423319, 0.07955071, 0.09571683, 0.08578045, 
    0.09827154, 0.08032203, 0.05637282, 0.09444162, 0.1584871, 0.3346539, 
    0.0640644, 0.0002459509, 0.0505346, 0.2214957, 0.08104566, 0.1879604, 
    0.3688,
  0.01861384, 0.03224168, 0.03389265, 0.09714969, 0.07000016, 0.08370389, 
    0.06958547, 0.07260762, 0.07378994, 0.01605261, 0.01072101, 0.01758106, 
    0.0574026, 0.03729181, 0.06541657, 0.06606956, 0.04688528, 0.0535213, 
    0.04791938, 0.06392852, 0.1613377, 0.09390497, 0.002341653, 0.03210286, 
    0.05800506, 0.03493337, 0.09629948, 0.1122173, 0.06049018,
  0.09041273, 0.1524259, 0.06701379, 0.1807032, 0.04008716, 0.03994445, 
    0.04033341, 0.02184631, 0.1489252, 0.1961398, 0.04577067, 0.02799922, 
    0.06308182, 0.04377358, 0.05395909, 0.06055844, 0.04003928, 0.02247524, 
    0.01733125, 0.02960266, 0.01235764, 0.007168008, 0.004856981, 0.05080514, 
    0.04397913, 0.02996205, 0.08463062, 0.07383652, 0.08548345,
  1.092905e-05, 1.523094e-06, 3.626687e-05, 0.0203367, 0.06951597, 0.1045484, 
    0.02926866, 0.07911131, 0.1457908, 0.09175659, 0.07283668, 0.05256142, 
    0.04492103, 0.05857106, 0.07669199, 0.05100794, 0.07521287, 0.09368189, 
    0.1118841, 0.1059627, 0.1178101, 0.04469085, 0.1014236, 0.06182288, 
    0.05955236, 0.09854353, 0.1216725, 0.001798032, 1.397835e-05,
  1.246423e-07, 2.729424e-09, 2.309594e-06, 0.02509971, 0.0009501975, 
    0.07969929, 0.02411656, 0.05420681, 0.1146855, 0.1801873, 0.1464418, 
    0.1438272, 0.07211789, 0.07980169, 0.06625366, 0.08377551, 0.08937014, 
    0.06456003, 0.142572, 0.1045682, 0.02409354, 0.2661179, 0.1077928, 
    0.07770828, 0.04821181, 0.05766678, 0.08820586, 0.01108535, 5.359365e-07,
  8.151076e-07, 0.03400949, 0.02209491, 0.03381331, 0.08144026, 0.02378817, 
    -7.575587e-05, 0.02315857, 0.1222198, 0.01992422, 0.2005877, 0.1413065, 
    0.140586, 0.1485424, 0.2140912, 0.1447124, 0.1793489, 0.1122214, 
    0.2472471, 0.0146088, 0.007305047, 0.06256001, 0.1130622, 0.13539, 
    0.1333074, 0.1126753, 0.06201182, 0.1365447, 0.01808797,
  0.01982678, 0.08939575, 0.1283237, 0.1679213, 0.06243688, 0.01783495, 
    0.08827665, 0.004480189, 0.000108617, 0.01961162, 0.141877, 0.2667225, 
    0.2729447, 0.215384, 0.2219003, 0.231225, 0.2946608, 0.2565677, 
    0.2384122, 0.1234343, 0.04092497, 0.05159362, 0.2248542, 0.1909631, 
    0.2586214, 0.2013246, 0.2227835, 0.2118362, 0.2018569,
  0.2579227, 0.3365558, 0.3235754, 0.2927501, 0.2107083, 0.168492, 0.1605732, 
    0.2122847, 0.08931753, 0.2681733, 0.1711145, 0.2603642, 0.3826545, 
    0.3562526, 0.2755704, 0.2946747, 0.2974877, 0.3167866, 0.3292615, 
    0.3508017, 0.1525109, 0.2981173, 0.3766816, 0.4853352, 0.2828184, 
    0.3039678, 0.2377103, 0.256183, 0.2311307,
  0.2176311, 0.4014354, 0.4188666, 0.4859053, 0.4352627, 0.3880696, 0.406852, 
    0.4638715, 0.4686898, 0.5392333, 0.4253376, 0.2190629, 0.1892756, 
    0.2271551, 0.5618337, 0.3350616, 0.2982074, 0.3356218, 0.3809577, 
    0.3108757, 0.3694112, 0.3861167, 0.4418094, 0.3910343, 0.3971488, 
    0.2658352, 0.2937129, 0.313256, 0.2499054,
  0.1543817, 0.2155097, 0.3515524, 0.3732017, 0.4664147, 0.4428531, 
    0.3530079, 0.488266, 0.420897, 0.4292747, 0.3375111, 0.2927842, 
    0.2390649, 0.38463, 0.4014439, 0.1796041, 0.2302444, 0.328659, 0.2285898, 
    0.3862022, 0.2757618, 0.2656366, 0.2926763, 0.2933571, 0.2285835, 
    0.3396333, 0.2344702, 0.2527991, 0.3333332,
  0.1875418, 0.244575, 0.2348374, 0.1545659, 0.1816456, 0.2307126, 0.21444, 
    0.1881851, 0.2115879, 0.2923194, 0.305425, 0.3050584, 0.2398508, 
    0.316566, 0.324333, 0.3351627, 0.3366123, 0.3417244, 0.3758692, 
    0.3075934, 0.2682475, 0.2415713, 0.1727305, 0.1787405, 0.2181844, 
    0.2383672, 0.08674347, 0.2153921, 0.2689934,
  0.2717947, 0.2725414, 0.2732881, 0.2740348, 0.2747815, 0.2755282, 
    0.2762749, 0.305345, 0.3053209, 0.3052967, 0.3052726, 0.3052485, 
    0.3052243, 0.3052002, 0.3180347, 0.324004, 0.3299733, 0.3359426, 
    0.3419118, 0.3478811, 0.3538504, 0.326802, 0.3201101, 0.3134183, 
    0.3067265, 0.3000346, 0.2933428, 0.2866509, 0.2711973,
  0.1452533, 0.165338, 0.161042, 0.1827312, 0.1776144, 0.2222392, 0.2255479, 
    0.1403827, 0.176667, 0.1884447, 0.1560501, 0.14537, 0.1827753, 
    0.03535711, 0.06847298, 0.09477926, 0.1221133, 0.1121086, 0.07308704, 
    0.06317015, 0.3066368, 0.415369, 0.4074395, 0.211781, 0.2088638, 
    0.2164157, 0.09698066, 0.07056835, 0.1199541,
  0.2634178, 0.1944943, 0.1939727, 0.1390525, 0.2377153, 0.3376287, 
    0.1165015, 0.2069017, 0.2695739, 0.3042062, 0.2190462, 0.1125686, 
    0.1879209, 0.1968572, 0.2708598, 0.3183513, 0.3230451, 0.3265204, 
    0.3856073, 0.3092871, 0.3460089, 0.3707318, 0.3813966, 0.625611, 
    0.1253774, 0.267511, 0.3653692, 0.4029356, 0.3336867,
  0.4262312, 0.427579, 0.4416826, 0.4335853, 0.4874514, 0.4318558, 0.4157208, 
    0.4270779, 0.3960753, 0.3487039, 0.3715327, 0.3764656, 0.3723081, 
    0.3628812, 0.3264664, 0.4258352, 0.4003096, 0.4560711, 0.3726132, 
    0.35123, 0.3431343, 0.3157094, 0.3217043, 0.3751312, 0.3115177, 
    0.3207079, 0.3600594, 0.3857129, 0.4261492,
  0.3766162, 0.3819997, 0.3766557, 0.3438373, 0.3541398, 0.356944, 0.3641928, 
    0.3406167, 0.3376014, 0.3561605, 0.28256, 0.2846094, 0.2326862, 
    0.3282008, 0.253662, 0.2801214, 0.3385642, 0.3335781, 0.3029856, 
    0.332026, 0.3374655, 0.3572372, 0.3768672, 0.161649, 0.0452536, 
    0.2368429, 0.3322086, 0.2853587, 0.2887604,
  0.334559, 0.2478075, 0.1487706, 0.228037, 0.2240088, 0.2250173, 0.261554, 
    0.3099748, 0.3189767, 0.2867377, 0.2645592, 0.1268204, 0.08798378, 
    0.2291653, 0.2521032, 0.3302211, 0.3003286, 0.2762186, 0.2617583, 
    0.3441603, 0.3222268, 0.2716473, 0.2820058, 0.09390645, 0.0431686, 
    0.2621168, 0.2816171, 0.2919783, 0.3284986,
  0.305263, 0.1256661, 0.02609495, 0.1109717, 0.1728958, 0.1551387, 
    0.1618575, 0.1949617, 0.2680718, 0.05761439, -0.0001167873, 1.555366e-05, 
    0.008268477, 0.1293722, 0.1683227, 0.1891696, 0.1348024, 0.1666881, 
    0.2343985, 0.2302783, 0.2126983, 0.1472253, 0.3727272, 0.0003655844, 
    0.009703092, 0.08450009, 0.1436939, 0.153264, 0.2002802,
  0.4969989, 0.0004364823, 0.01577485, 0.05749838, 0.1122046, 0.08695699, 
    0.1089246, 0.127298, 0.1720647, -0.0002100067, 2.91346e-05, 
    -1.668198e-07, 0.0868867, 0.0832396, 0.1330172, 0.1289599, 0.1215946, 
    0.09978811, 0.07646804, 0.08601819, 0.1127896, 0.3022588, 0.5390134, 
    0.002296705, 0.03840179, 0.2179868, 0.07643994, 0.1073332, 0.3580676,
  0.2077406, 0.08528998, 0.02188079, 0.1092288, 0.08763985, 0.08798113, 
    0.09171669, 0.09055022, 0.1752008, 0.1079784, 0.02601875, 0.05962949, 
    0.07857421, 0.05662123, 0.07801347, 0.06982384, 0.06756043, 0.1027945, 
    0.06940576, 0.06944403, 0.1636652, 0.4493634, 0.06057849, 0.01671673, 
    0.03738484, 0.02528174, 0.1171293, 0.1123451, 0.3641221,
  0.08316782, 0.1340823, 0.04811959, 0.1631368, 0.1028314, 0.1286889, 
    0.1523164, 0.07286991, 0.1268467, 0.158124, 0.06439148, 0.0768632, 
    0.125347, 0.1092559, 0.1137504, 0.09763669, 0.1070082, 0.0825514, 
    0.09316161, 0.09407014, 0.08954723, 0.03253271, 0.030401, 0.03168904, 
    0.02192791, 0.04777563, 0.0916808, 0.07883698, 0.08759815,
  5.550519e-06, 4.381632e-07, 1.923238e-05, 0.01054741, 0.08813789, 
    0.1237979, 0.01664331, 0.07605141, 0.1454956, 0.1052671, 0.06608652, 
    0.05413438, 0.06976059, 0.07641778, 0.05793978, 0.06655926, 0.08517581, 
    0.1273629, 0.1465297, 0.1066322, 0.1297657, 0.05737163, 0.1239748, 
    0.07106899, 0.06720354, 0.06771831, 0.1033944, 0.04627041, 6.109165e-06,
  7.555845e-08, 1.114135e-09, 1.546296e-06, 0.01754727, 0.0007365327, 
    0.04102313, 0.01399574, 0.0654261, 0.07705428, 0.1459792, 0.107751, 
    0.1205994, 0.1025875, 0.1042669, 0.09388101, 0.07852598, 0.127531, 
    0.06830113, 0.2577125, 0.201506, 0.08641992, 0.2826662, 0.06550974, 
    0.06202397, 0.06327632, 0.05600743, 0.09294339, 0.02037046, 2.108724e-07,
  4.506663e-07, 0.03296422, 0.02011725, 0.04468564, 0.07173922, 0.01431438, 
    -0.0006114971, 0.01247459, 0.1175761, 0.01110725, 0.1195975, 0.1163561, 
    0.1115205, 0.1259946, 0.1724238, 0.1262844, 0.1277412, 0.08514234, 
    0.257349, 0.02801942, 0.009512072, 0.07731552, 0.1232832, 0.08648592, 
    0.1299269, 0.154115, 0.0596114, 0.09265067, 0.02039927,
  0.01920703, 0.08901705, 0.138199, 0.1767105, 0.04832996, 0.006417659, 
    0.1031557, 0.00225899, -2.758244e-05, 0.01814498, 0.1602054, 0.1498076, 
    0.1824123, 0.1639236, 0.2040138, 0.2161696, 0.2631667, 0.2816327, 
    0.2497451, 0.1369111, 0.04038428, 0.08101256, 0.2742911, 0.1820166, 
    0.1930951, 0.2256906, 0.2243284, 0.2347203, 0.1624216,
  0.2494873, 0.3675204, 0.3283206, 0.3603257, 0.2788665, 0.172125, 0.157277, 
    0.224098, 0.09380025, 0.285055, 0.1409019, 0.2786848, 0.2488323, 
    0.2738851, 0.2558877, 0.2619633, 0.2918463, 0.3166224, 0.3183215, 
    0.3847302, 0.1843942, 0.288227, 0.3458494, 0.6007056, 0.3090201, 
    0.2841627, 0.2309001, 0.2354532, 0.2048011,
  0.1796895, 0.4006446, 0.5174059, 0.5519655, 0.5128806, 0.4070134, 
    0.4932067, 0.5449857, 0.506794, 0.5785071, 0.4695985, 0.2389331, 
    0.1704763, 0.2141708, 0.5915806, 0.328777, 0.3166496, 0.3345931, 
    0.3976114, 0.3074965, 0.4343424, 0.3806475, 0.3470943, 0.3836264, 
    0.3022864, 0.2161327, 0.2493479, 0.2494179, 0.2063465,
  0.09969594, 0.1412963, 0.3214893, 0.2816359, 0.4022149, 0.4896767, 
    0.3954591, 0.5258345, 0.4255263, 0.4497444, 0.3738609, 0.3233213, 
    0.2794482, 0.4636551, 0.443724, 0.2398617, 0.2627275, 0.3537797, 
    0.2994702, 0.4373058, 0.3154141, 0.2880799, 0.3030289, 0.3359986, 
    0.2672453, 0.3472645, 0.2401596, 0.2160129, 0.215721,
  0.2379825, 0.3323638, 0.2670512, 0.2018834, 0.2115869, 0.2784097, 
    0.2228546, 0.2308422, 0.245696, 0.3856189, 0.3801385, 0.3656298, 
    0.3281156, 0.372396, 0.3705637, 0.3641911, 0.3778813, 0.3699495, 
    0.3887011, 0.3436427, 0.3328676, 0.2562347, 0.2050826, 0.172625, 
    0.2266066, 0.2852515, 0.1336786, 0.2427998, 0.2993919,
  0.324219, 0.3280234, 0.3318278, 0.3356322, 0.3394367, 0.343241, 0.3470455, 
    0.3534856, 0.350188, 0.3468903, 0.3435926, 0.3402949, 0.3369972, 
    0.3336995, 0.3597578, 0.3649035, 0.3700493, 0.375195, 0.3803408, 
    0.3854865, 0.3906322, 0.3472135, 0.3415611, 0.3359086, 0.3302562, 
    0.3246037, 0.3189512, 0.3132988, 0.3211754,
  0.13681, 0.1613663, 0.1621262, 0.2115435, 0.2246166, 0.2555985, 0.2455645, 
    0.1563981, 0.2328153, 0.221071, 0.1826443, 0.1577478, 0.1946003, 
    0.03175826, 0.08822198, 0.1858066, 0.1974794, 0.1437773, 0.1127325, 
    0.07057802, 0.2953242, 0.4345082, 0.3898675, 0.204633, 0.1692941, 
    0.203742, 0.07489089, 0.05350364, 0.1303888,
  0.2408373, 0.1542477, 0.1884048, 0.1141745, 0.1994561, 0.3162435, 
    0.08514784, 0.1761139, 0.2342883, 0.2718489, 0.1866477, 0.1021119, 
    0.1433859, 0.1796593, 0.2774795, 0.3174732, 0.3212596, 0.2994502, 
    0.3794591, 0.3436052, 0.3364416, 0.3628315, 0.3552611, 0.588432, 
    0.1067989, 0.2584006, 0.3813363, 0.4150633, 0.3275207,
  0.3902704, 0.3903287, 0.43825, 0.4226742, 0.4483536, 0.4300404, 0.3947438, 
    0.3922324, 0.4067192, 0.3315844, 0.3525906, 0.3452513, 0.3838398, 
    0.3424743, 0.3483146, 0.4551737, 0.4375555, 0.4907698, 0.4135453, 
    0.3156957, 0.3102016, 0.281412, 0.3027812, 0.4004228, 0.3311321, 
    0.3780533, 0.3451804, 0.4245256, 0.4659406,
  0.4198641, 0.4160924, 0.3940642, 0.3448561, 0.3229021, 0.3244484, 
    0.3518659, 0.3152728, 0.321587, 0.3393381, 0.2569997, 0.2665001, 
    0.1891934, 0.2720788, 0.2275499, 0.2882319, 0.3117341, 0.3753062, 
    0.4296498, 0.3473934, 0.3521393, 0.3796524, 0.3800239, 0.1449524, 
    0.04458649, 0.2529066, 0.4019382, 0.3050748, 0.3292364,
  0.2932105, 0.2006488, 0.1071414, 0.1835425, 0.1823227, 0.1675732, 
    0.2138715, 0.2638925, 0.3219383, 0.2364612, 0.2353631, 0.09095658, 
    0.06661545, 0.1865368, 0.2631968, 0.335656, 0.2803742, 0.2204775, 
    0.2437311, 0.2568864, 0.317607, 0.2614664, 0.2493114, 0.1162177, 
    0.03944264, 0.2101173, 0.2807801, 0.3119616, 0.3099133,
  0.1350721, 0.09132721, 0.02220302, 0.09763901, 0.1738845, 0.1086577, 
    0.1067756, 0.1454227, 0.2530937, 0.05065287, 0.000427093, 4.268659e-06, 
    0.003436753, 0.1327978, 0.1479882, 0.09276138, 0.07900098, 0.1044041, 
    0.1891274, 0.1452988, 0.1596958, 0.0720531, 0.2708278, 0.01488765, 
    0.01059277, 0.09121475, 0.1404447, 0.09717697, 0.09201614,
  0.3220425, 0.0002242259, 0.01961921, 0.06820722, 0.05734254, 0.05551627, 
    0.06682557, 0.09393483, 0.2128471, -0.0002208253, 1.71598e-05, 
    -1.836299e-06, 0.1221342, 0.05913406, 0.06961246, 0.07854325, 0.03947151, 
    0.1149916, 0.05935568, 0.03515685, 0.03319805, 0.09718205, 0.4693117, 
    0.08117595, 0.02377072, 0.1984209, 0.05060884, 0.02229742, 0.1509639,
  0.4626772, 0.1902121, 0.01094582, 0.1450606, 0.09947857, 0.0700352, 
    0.05683452, 0.03993985, 0.07783733, 0.1010363, 0.02258482, 0.05739067, 
    0.06767593, 0.03472755, 0.03837065, 0.03111825, 0.02796127, 0.0387302, 
    0.01546875, 0.01665368, 0.05644376, 0.3072394, 0.5943828, 0.006933151, 
    0.02460599, 0.01840549, 0.03104955, 0.04462606, 0.2222117,
  0.07776591, 0.1144004, 0.03118586, 0.1517969, 0.1180393, 0.1112497, 
    0.1120134, 0.2135277, 0.1054499, 0.1104412, 0.01874498, 0.06264222, 
    0.01894139, 0.02177333, 0.04033624, 0.04122005, 0.04913493, 0.07810267, 
    0.09878865, 0.1426553, 0.3393423, 0.3346532, 0.1481166, 0.0233673, 
    0.008261534, 0.04942112, 0.08752511, 0.08022408, 0.1207334,
  1.950637e-06, -4.142082e-09, 9.735064e-06, 0.01125985, 0.0970113, 
    0.06034735, 0.01355237, 0.03338131, 0.04736379, 0.05286074, 0.05113502, 
    0.03533297, 0.03716992, 0.03908189, 0.02710688, 0.0362901, 0.05870728, 
    0.07694916, 0.1172985, 0.09368353, 0.09873566, 0.08868504, 0.2247567, 
    0.06527165, 0.02250472, 0.01918607, 0.03430801, 0.04888843, 2.942747e-06,
  7.360912e-08, 6.981394e-10, 1.20068e-06, 0.007067774, 0.0003133018, 
    0.02040922, 0.01564607, 0.01851678, 0.04829933, 0.06960943, 0.05347146, 
    0.04582214, 0.05703133, 0.04623232, 0.03422769, 0.0229781, 0.0548273, 
    0.08015253, 0.1430936, 0.1594442, 0.05840527, 0.2182238, 0.01738892, 
    0.0316189, 0.04645529, 0.01716662, 0.01992296, 0.002643096, 1.16562e-07,
  6.75665e-08, 0.02568294, 0.01228477, 0.04333727, 0.06362577, 0.0132266, 
    -0.0006036562, 0.00589807, 0.113011, 0.007814202, 0.07264737, 0.09378463, 
    0.09386124, 0.1023491, 0.1267731, 0.0911914, 0.09004023, 0.05489598, 
    0.1877104, 0.03378706, 0.009934333, 0.0857006, 0.1274381, 0.0429308, 
    0.06661127, 0.1119528, 0.01959277, 0.03046995, 0.01761992,
  0.02305113, 0.05824098, 0.1231786, 0.1737356, 0.02475782, 0.003659421, 
    0.1169445, 0.003009497, -1.20926e-05, 0.0192989, 0.1791299, 0.09363885, 
    0.1162634, 0.1174563, 0.1691694, 0.175017, 0.2167922, 0.2522653, 
    0.2358883, 0.1511419, 0.02781802, 0.09748006, 0.2462876, 0.1372351, 
    0.1517309, 0.2260572, 0.2033107, 0.1765931, 0.1260463,
  0.2112165, 0.3933132, 0.3411216, 0.4107705, 0.2804218, 0.1901093, 
    0.1388439, 0.2238252, 0.09271412, 0.2915779, 0.09926501, 0.2967155, 
    0.1686383, 0.2120351, 0.215703, 0.2180686, 0.2621417, 0.293456, 
    0.2796748, 0.4127911, 0.1993686, 0.2529868, 0.293521, 0.6462932, 
    0.2920792, 0.2459198, 0.2029935, 0.2260961, 0.1813075,
  0.1329616, 0.4299504, 0.5171055, 0.6383076, 0.6532993, 0.4017554, 
    0.5578228, 0.6169946, 0.5861584, 0.5697139, 0.5217924, 0.3008116, 
    0.1661393, 0.2376092, 0.4510593, 0.2954489, 0.3427874, 0.317987, 
    0.3976959, 0.3432662, 0.4939589, 0.344613, 0.2259989, 0.3624124, 
    0.2397998, 0.1689821, 0.2014378, 0.1951892, 0.1672619,
  0.07080146, 0.0832444, 0.3013935, 0.1670475, 0.3203522, 0.4490204, 
    0.4834222, 0.5258505, 0.4312336, 0.4843254, 0.4180414, 0.3297105, 
    0.3215103, 0.5309957, 0.4702041, 0.3197352, 0.2867166, 0.3533911, 
    0.3224592, 0.4585681, 0.3902468, 0.3642855, 0.3160722, 0.3427316, 
    0.2086343, 0.3497536, 0.2530023, 0.1869931, 0.1403993,
  0.2096654, 0.328943, 0.2955874, 0.2093382, 0.2273926, 0.2947989, 0.2960318, 
    0.2739733, 0.3134287, 0.4828175, 0.4291776, 0.4230373, 0.4001644, 
    0.4525986, 0.4584713, 0.4474224, 0.4301004, 0.4393487, 0.4110544, 
    0.3961423, 0.3724934, 0.2548871, 0.2236664, 0.1777133, 0.2216, 0.3037745, 
    0.1606732, 0.2668588, 0.3060291,
  0.4185333, 0.4224356, 0.426338, 0.4302404, 0.4341427, 0.4380451, 0.4419475, 
    0.4230013, 0.4185313, 0.4140612, 0.4095911, 0.4051211, 0.400651, 
    0.3961809, 0.4230217, 0.4264905, 0.4299593, 0.4334281, 0.436897, 
    0.4403658, 0.4438346, 0.4026106, 0.3997095, 0.3968084, 0.3939072, 
    0.3910061, 0.388105, 0.3852039, 0.4154114,
  0.1372469, 0.1588346, 0.158629, 0.2225762, 0.2597044, 0.2802697, 0.2610403, 
    0.1712912, 0.2670675, 0.265698, 0.2054272, 0.1499897, 0.2022686, 
    0.01984158, 0.1582877, 0.2317424, 0.2146435, 0.1554654, 0.1240886, 
    0.0807133, 0.2681056, 0.4195309, 0.3759897, 0.1790414, 0.1371235, 
    0.2093574, 0.05890474, 0.05453779, 0.1260133,
  0.1906236, 0.1233503, 0.1493092, 0.09093477, 0.1539881, 0.275511, 
    0.05314644, 0.1224843, 0.1807573, 0.2106897, 0.144671, 0.08358192, 
    0.1057382, 0.1557718, 0.265484, 0.3081834, 0.3281364, 0.2799031, 
    0.3795832, 0.3138399, 0.3090777, 0.3207008, 0.3426454, 0.5177409, 
    0.08025832, 0.2645079, 0.3753167, 0.3935991, 0.2981372,
  0.3595257, 0.3558837, 0.4061903, 0.4044865, 0.3946289, 0.3985135, 
    0.4036667, 0.3693419, 0.3920508, 0.3010931, 0.3118106, 0.3160638, 
    0.3714951, 0.3120672, 0.3403919, 0.4383765, 0.4652746, 0.501894, 
    0.4116476, 0.2954242, 0.2809243, 0.260139, 0.2715088, 0.3468906, 
    0.3213955, 0.3973771, 0.370426, 0.4562252, 0.4736512,
  0.3867968, 0.3831501, 0.3698082, 0.2970343, 0.2843792, 0.2875192, 
    0.3215438, 0.2868368, 0.298547, 0.3158859, 0.2229395, 0.2412432, 
    0.1484305, 0.2382875, 0.1896306, 0.276081, 0.3047036, 0.3409731, 
    0.3746552, 0.3520201, 0.3169776, 0.367248, 0.3133972, 0.1268147, 
    0.05778328, 0.275639, 0.4016468, 0.2986247, 0.3636566,
  0.2394294, 0.1336295, 0.0579517, 0.1566894, 0.1667114, 0.1576246, 0.178351, 
    0.2187012, 0.2717865, 0.1842065, 0.1462279, 0.0478861, 0.03193475, 
    0.152855, 0.262801, 0.2736815, 0.2570417, 0.1693089, 0.1928675, 
    0.2128742, 0.2790471, 0.2306062, 0.1888868, 0.1231487, 0.03735661, 
    0.1775163, 0.2427674, 0.2649728, 0.2683787,
  0.04391322, 0.06237398, 0.01700803, 0.1163593, 0.1541368, 0.06308955, 
    0.06277269, 0.08101733, 0.1453497, 0.02069051, 0.0003266745, 
    1.139016e-06, 0.002967487, 0.1333555, 0.1115971, 0.06777922, 0.04052275, 
    0.07415831, 0.1500748, 0.0920549, 0.09423581, 0.03019825, 0.1136053, 
    0.01997658, 0.009906535, 0.07784204, 0.1386099, 0.05594629, 0.02971793,
  0.1175482, 0.01098084, 0.01510576, 0.02425648, 0.01723649, 0.02353222, 
    0.03146401, 0.04315383, 0.1065841, -6.45354e-05, 5.293763e-06, 
    -1.631488e-06, 0.04913376, 0.02169309, 0.02541512, 0.03213794, 
    0.01523364, 0.05663795, 0.02936649, 0.01485994, 0.007490172, 0.02959387, 
    0.1847726, 0.1280925, 0.01575791, 0.1901272, 0.03013852, 0.0042852, 
    0.04596245,
  0.2346841, 0.1513935, 0.006317044, 0.2073942, 0.01916326, 0.03268696, 
    0.01994071, 0.007529764, 0.02261355, 0.02445601, 0.009481657, 0.01416814, 
    0.02616166, 0.007946373, 0.01545851, 0.009575434, 0.003604243, 
    0.005775275, 0.002473716, 0.003327263, 0.01498541, 0.1036777, 0.3674768, 
    0.003302305, 0.02120696, 0.01598153, 0.0003675183, 0.006983151, 0.09079036,
  0.09772269, 0.09605893, 0.02091307, 0.1427632, 0.02270734, 0.02159748, 
    0.01776973, 0.02782912, 0.092953, 0.06868076, 0.006936054, 0.006778213, 
    0.004122015, 0.007809972, 0.009487783, 0.009038188, 0.008543111, 
    0.01895905, 0.02751739, 0.05272263, 0.1685515, 0.4566821, 0.371122, 
    0.0112006, 0.005300403, 0.01570294, 0.04875451, 0.04006114, 0.1395953,
  2.594871e-06, 1.997558e-07, 5.36607e-06, 0.009731774, 0.08068638, 
    0.01213988, 0.005091743, 0.01357558, 0.01492105, 0.0363284, 0.02841695, 
    0.008547232, 0.0171663, 0.02147254, 0.01015217, 0.0106475, 0.02068833, 
    0.03851645, 0.07245426, 0.06806287, 0.06351096, 0.03302155, 0.2902772, 
    0.05626535, 0.006534118, 0.007764717, 0.009899606, 0.008431777, 
    1.63118e-06,
  7.24087e-08, 5.81675e-10, 1.033262e-06, 0.003183236, 0.0001114739, 
    0.005656744, 0.01072003, 0.004744483, 0.03813071, 0.02627994, 0.02467034, 
    0.01604014, 0.0150619, 0.0174995, 0.0101006, 0.006128273, 0.02806844, 
    0.03660034, 0.07447971, 0.07071552, 0.0205585, 0.1592461, 0.004069503, 
    0.0137659, 0.008497464, 0.005169821, 0.005356461, 0.0006619347, 
    8.917793e-08,
  -8.229693e-07, 0.02051751, 0.003812296, 0.03494602, 0.06067374, 0.02115892, 
    -0.0008125041, 0.002881024, 0.09932169, 0.008309661, 0.02576685, 
    0.05757134, 0.06446853, 0.06611059, 0.09783405, 0.04949273, 0.05094416, 
    0.04347486, 0.1368289, 0.03822805, 0.01056042, 0.07248557, 0.1108748, 
    0.02298355, 0.03326028, 0.05571561, 0.005159322, 0.009734631, 0.01845611,
  0.01053741, 0.02794671, 0.09203419, 0.1686543, 0.0230407, 0.003028035, 
    0.1200021, 0.002758815, -6.017894e-05, 0.01632152, 0.1846837, 0.06217858, 
    0.0851402, 0.08783132, 0.1295974, 0.1363488, 0.1874251, 0.2080777, 
    0.2000668, 0.1551818, 0.01921594, 0.08816709, 0.1969711, 0.1088679, 
    0.1141068, 0.1823022, 0.1733943, 0.1157738, 0.08736133,
  0.1728036, 0.3859516, 0.3428082, 0.399709, 0.2227258, 0.1770248, 0.1244475, 
    0.213529, 0.06954607, 0.2349689, 0.08334339, 0.3132099, 0.1154684, 
    0.165421, 0.1725181, 0.196358, 0.2208081, 0.2547735, 0.2420215, 0.436371, 
    0.1891591, 0.2157442, 0.2807769, 0.6583039, 0.2455899, 0.2011055, 
    0.1839205, 0.2090253, 0.1616104,
  0.09947853, 0.448545, 0.4768468, 0.7435763, 0.741574, 0.4225194, 0.624428, 
    0.6231753, 0.5951318, 0.5645487, 0.5841337, 0.3717058, 0.1654373, 
    0.2110913, 0.3438739, 0.2485341, 0.3624369, 0.2854815, 0.3823273, 
    0.3888307, 0.5799905, 0.2677122, 0.1490767, 0.3401825, 0.1865957, 
    0.1293044, 0.170075, 0.1408043, 0.1239327,
  0.04634804, 0.05798686, 0.2888946, 0.09575844, 0.2207632, 0.3830765, 
    0.5669655, 0.5085838, 0.4090387, 0.5107404, 0.4443821, 0.3397895, 
    0.3631199, 0.5666655, 0.4843789, 0.3422138, 0.3352966, 0.3585384, 
    0.3663541, 0.4537441, 0.4073184, 0.4569283, 0.328097, 0.3785667, 
    0.1375355, 0.3532361, 0.2647754, 0.1592688, 0.0947166,
  0.2510653, 0.3569729, 0.3074085, 0.2597833, 0.2650741, 0.3311239, 
    0.3597882, 0.366847, 0.4360824, 0.5325093, 0.4976272, 0.4732625, 
    0.4778178, 0.5520097, 0.5500571, 0.5245506, 0.4978805, 0.4945617, 
    0.5136874, 0.4745664, 0.4388962, 0.2459257, 0.2596678, 0.2219398, 
    0.207021, 0.3204734, 0.1712158, 0.2890783, 0.3381322,
  0.4728012, 0.4780032, 0.4832052, 0.4884072, 0.4936092, 0.4988112, 
    0.5040131, 0.4757563, 0.4749997, 0.474243, 0.4734863, 0.4727296, 
    0.4719729, 0.4712163, 0.5265635, 0.5253418, 0.5241201, 0.5228984, 
    0.5216768, 0.5204551, 0.5192333, 0.4710826, 0.4678589, 0.4646353, 
    0.4614117, 0.4581881, 0.4549644, 0.4517408, 0.4686397,
  0.1314775, 0.1593983, 0.1564441, 0.2154764, 0.275385, 0.266441, 0.2585962, 
    0.1935101, 0.2766041, 0.2625926, 0.1936657, 0.1157099, 0.1649372, 
    0.01141609, 0.1619837, 0.2193021, 0.2077176, 0.1828271, 0.1315722, 
    0.0798504, 0.2292084, 0.3693984, 0.3362695, 0.1402015, 0.09972738, 
    0.1724856, 0.03851631, 0.05386204, 0.109033,
  0.1511755, 0.0954344, 0.1122164, 0.06949177, 0.1123262, 0.2264163, 
    0.03049101, 0.08042295, 0.1314653, 0.153151, 0.09558824, 0.06654779, 
    0.07386259, 0.1330793, 0.2469386, 0.3050272, 0.2816948, 0.2554294, 
    0.3482269, 0.266862, 0.271423, 0.2688706, 0.3065366, 0.4632766, 
    0.06871553, 0.2773214, 0.3415342, 0.3243722, 0.2545642,
  0.3187073, 0.2982773, 0.3554196, 0.3366057, 0.3386951, 0.3481885, 
    0.3616816, 0.3113535, 0.3465413, 0.2708977, 0.2694057, 0.2860059, 
    0.3368415, 0.2744795, 0.2983572, 0.3990361, 0.4329516, 0.4663318, 
    0.3618819, 0.2619646, 0.2558691, 0.2251366, 0.2331605, 0.2987692, 
    0.2986957, 0.3941269, 0.4127926, 0.4349309, 0.4114288,
  0.3322351, 0.3233, 0.3264546, 0.2602137, 0.2509888, 0.2434648, 0.2800724, 
    0.2363045, 0.266951, 0.2931914, 0.1830222, 0.2040642, 0.1096065, 
    0.1909137, 0.1844908, 0.2397341, 0.2592758, 0.2633056, 0.2782416, 
    0.2733158, 0.2649313, 0.3262105, 0.2568156, 0.106597, 0.06042581, 
    0.2889875, 0.3792188, 0.3082118, 0.3746575,
  0.1796949, 0.07320932, 0.03042648, 0.1320275, 0.1406696, 0.1216532, 
    0.1367967, 0.1803293, 0.2072512, 0.1206384, 0.07832678, 0.02313768, 
    0.01916019, 0.1296902, 0.2460643, 0.2304836, 0.2206589, 0.1483394, 
    0.1701194, 0.1683224, 0.2499358, 0.1938492, 0.1585507, 0.1186623, 
    0.02956564, 0.1522263, 0.1977788, 0.2256386, 0.1996528,
  0.01941978, 0.02976836, 0.01358381, 0.1244643, 0.1040676, 0.03137477, 
    0.03485804, 0.03670444, 0.08109322, 0.03810358, 0.0002008834, 
    4.305163e-07, 0.004407463, 0.08840479, 0.06028533, 0.04150108, 
    0.02680266, 0.05215368, 0.1309431, 0.06664395, 0.05257227, 0.009729415, 
    0.05001158, 0.03153189, 0.006312639, 0.05462547, 0.09719466, 0.0346169, 
    0.01192389,
  0.04691183, 0.0180827, 0.007627151, 0.009410284, 0.001563959, 0.006962951, 
    0.01298913, 0.02267532, 0.05351869, -3.093027e-05, 3.579017e-07, 
    -7.57285e-07, 0.01434682, 0.009113488, 0.01125701, 0.0160168, 
    0.004739564, 0.02268632, 0.01292444, 0.00726535, 0.002543868, 0.01169586, 
    0.07634412, 0.05506194, 0.01086224, 0.1797644, 0.01538055, 0.001550242, 
    0.01547762,
  0.09514502, 0.04741861, 0.00443323, 0.2048938, 0.004792563, 0.01103716, 
    0.006524479, 0.001465111, 0.006134677, 0.006651592, 0.003219318, 
    0.005008878, 0.008715402, 0.0009942537, 0.00650399, 0.004885026, 
    0.0002860251, 0.001541896, 0.0009887643, 0.001424565, 0.006136095, 
    0.04145357, 0.1451349, 0.00361447, 0.01853043, 0.01539084, -0.00114988, 
    0.002072396, 0.03033341,
  0.02541262, 0.09830632, 0.02024764, 0.1223903, 0.005894662, 0.00712167, 
    0.004380603, 0.00811534, 0.08540668, 0.04656333, 0.001554862, 
    0.001700581, 0.001524266, 0.002879813, 0.003829277, 0.003375941, 
    0.00250542, 0.005265919, 0.007539192, 0.01364483, 0.04749381, 0.173889, 
    0.1538545, 0.008243097, 0.002011667, 0.002260355, 0.03595278, 
    0.005094931, 0.03500715,
  3.797409e-06, 5.381309e-08, 2.929778e-06, 0.006380895, 0.06099021, 
    0.003998886, 4.80318e-05, 0.005346365, 0.004928521, 0.01651298, 
    0.01259451, 0.002087681, 0.005519562, 0.009617891, 0.002951708, 
    0.001898731, 0.0103863, 0.01340724, 0.03441713, 0.02631645, 0.03538103, 
    0.007368444, 0.2475607, 0.04735191, 0.00256262, 0.003373775, 0.003550984, 
    0.003216243, -2.904061e-07,
  7.077649e-08, 5.460696e-10, 7.71513e-07, 0.001648693, 0.001088678, 
    0.002382508, 0.006379708, 0.002250252, 0.03082664, 0.00992288, 
    0.00758609, 0.006375299, 0.005069952, 0.006969799, 0.002096395, 
    0.001898331, 0.01070483, 0.01524024, 0.02862085, 0.024631, 0.008846958, 
    0.1214185, 0.001318835, 0.004047867, 0.002494585, 0.002056587, 
    0.002398478, 0.000314725, 8.375931e-08,
  -9.605486e-06, 0.0133498, 0.000620669, 0.02876841, 0.04829914, 0.01224917, 
    -0.0006242328, 0.001732323, 0.08618842, 0.01382811, 0.01201436, 
    0.0390824, 0.04021747, 0.03568156, 0.06757765, 0.02515874, 0.02445091, 
    0.02519356, 0.08802484, 0.03073389, 0.009327454, 0.05755906, 0.09391906, 
    0.01515361, 0.01761533, 0.03409051, 0.001712264, 0.004056687, 0.01371526,
  0.006431371, 0.010781, 0.05974988, 0.1628997, 0.009187873, 0.00221106, 
    0.1142817, 0.002711162, -9.766503e-05, 0.01179225, 0.1788734, 0.0433266, 
    0.06625713, 0.06709628, 0.1008985, 0.1086843, 0.1645018, 0.1691948, 
    0.138702, 0.1524014, 0.01226471, 0.08243895, 0.1615598, 0.08531892, 
    0.08214545, 0.1412054, 0.1371778, 0.0727766, 0.05346575,
  0.1239123, 0.3663799, 0.3350332, 0.3552235, 0.2428618, 0.1565547, 
    0.09784718, 0.2005953, 0.04976258, 0.1761954, 0.07201168, 0.3130987, 
    0.08623414, 0.1242792, 0.1286694, 0.1741815, 0.1838508, 0.2204017, 
    0.2198602, 0.4507513, 0.1673839, 0.1726738, 0.237184, 0.6407361, 
    0.1935394, 0.1768035, 0.1624317, 0.1944204, 0.128141,
  0.0718731, 0.4657638, 0.4487099, 0.7506394, 0.7184306, 0.4147989, 
    0.6357707, 0.6023139, 0.5907739, 0.5229979, 0.5668116, 0.4167489, 
    0.1586768, 0.2058563, 0.2694861, 0.2183293, 0.3726593, 0.2432219, 
    0.3423087, 0.4025289, 0.6381185, 0.2109792, 0.102132, 0.2989233, 
    0.1399663, 0.1077591, 0.1366133, 0.09695613, 0.094327,
  0.03076933, 0.03130636, 0.2863602, 0.05823173, 0.1586937, 0.3013152, 
    0.591264, 0.4263384, 0.394702, 0.5039443, 0.4731661, 0.3633453, 
    0.4364098, 0.5822929, 0.5032033, 0.3798396, 0.3628014, 0.3753816, 
    0.3910547, 0.4419123, 0.4591851, 0.5356132, 0.3695683, 0.4507759, 
    0.1017509, 0.3347616, 0.2708104, 0.1308839, 0.06798519,
  0.3630989, 0.3724338, 0.3710351, 0.3215636, 0.2681529, 0.4237081, 
    0.4656607, 0.4849907, 0.5068181, 0.5997059, 0.5618758, 0.5455566, 
    0.585636, 0.6031506, 0.6141537, 0.5801357, 0.5603579, 0.6182033, 
    0.6415449, 0.5456219, 0.4577947, 0.2594198, 0.3019566, 0.2830925, 
    0.2194297, 0.3297224, 0.1772329, 0.3089396, 0.4685544,
  0.497998, 0.5033593, 0.5087206, 0.514082, 0.5194433, 0.5248047, 0.530166, 
    0.4774241, 0.4796249, 0.4818257, 0.4840265, 0.4862273, 0.4884281, 
    0.4906288, 0.5726797, 0.5690777, 0.5654758, 0.5618739, 0.5582719, 
    0.55467, 0.5510681, 0.5271969, 0.5232367, 0.5192765, 0.5153164, 
    0.5113562, 0.507396, 0.5034358, 0.4937089,
  0.1160916, 0.1603948, 0.139739, 0.1881765, 0.2746814, 0.2333064, 0.2401636, 
    0.2137266, 0.2253875, 0.1935889, 0.1392443, 0.06839187, 0.1077424, 
    0.008062276, 0.1753322, 0.2447745, 0.2067068, 0.181825, 0.1074582, 
    0.08866853, 0.1823287, 0.3277254, 0.2827378, 0.09751922, 0.08238621, 
    0.1571723, 0.03042769, 0.04736832, 0.08606156,
  0.1295578, 0.07486141, 0.09063414, 0.05509307, 0.08350955, 0.1758304, 
    0.02023106, 0.0534263, 0.09896072, 0.1088382, 0.06761094, 0.05644394, 
    0.05240599, 0.1067578, 0.2347237, 0.2688226, 0.235522, 0.2264496, 
    0.3080786, 0.223385, 0.2499135, 0.2254739, 0.2536944, 0.4079362, 
    0.05661563, 0.262285, 0.2794711, 0.2558309, 0.2248368,
  0.2709503, 0.2411103, 0.2923763, 0.2541568, 0.2728575, 0.2646172, 
    0.2653158, 0.2411091, 0.2824731, 0.2118265, 0.2236976, 0.2400469, 
    0.2854168, 0.2319359, 0.2469653, 0.3460455, 0.379226, 0.3889914, 
    0.2986658, 0.2298722, 0.2103819, 0.1769957, 0.1802711, 0.2410833, 
    0.2567124, 0.3772908, 0.3924155, 0.3626497, 0.3200628,
  0.289814, 0.2589266, 0.2567511, 0.2089163, 0.1963558, 0.1832408, 0.2287201, 
    0.1827798, 0.2228819, 0.2407383, 0.1415934, 0.1566172, 0.06859353, 
    0.1386149, 0.1847934, 0.1980609, 0.193292, 0.1890594, 0.2124214, 
    0.1912047, 0.1858292, 0.2577405, 0.1967266, 0.0874209, 0.0762568, 
    0.263353, 0.3471775, 0.2921776, 0.3407736,
  0.1270251, 0.03823682, 0.01791021, 0.1050802, 0.1013291, 0.08481129, 
    0.1006537, 0.1305438, 0.1471823, 0.07579188, 0.04587265, 0.01162468, 
    0.01285137, 0.1109745, 0.2121764, 0.1777033, 0.181322, 0.137398, 
    0.139616, 0.1429775, 0.2249282, 0.1576115, 0.1232495, 0.1089384, 
    0.02903205, 0.1288741, 0.1418459, 0.1820955, 0.161164,
  0.0116925, 0.01532187, 0.01118148, 0.08563209, 0.06299801, 0.01474288, 
    0.01842308, 0.0165661, 0.0476144, 0.02458079, 0.0001014291, 2.284248e-07, 
    0.00261577, 0.03938878, 0.02954572, 0.02420225, 0.01636787, 0.03169239, 
    0.09178156, 0.04515507, 0.03327049, 0.003922731, 0.02612503, 0.02905371, 
    0.004117684, 0.02532467, 0.05865912, 0.01785108, 0.006312794,
  0.02363524, 0.01380037, 0.004378391, 0.004321266, -0.000624681, 
    0.002583642, 0.003214176, 0.006657987, 0.027047, 5.894635e-07, 
    7.05268e-08, -9.100106e-07, 0.005680332, 0.003072805, 0.006045103, 
    0.007036512, 0.001903671, 0.009343482, 0.006332651, 0.004648557, 
    0.001224115, 0.006317159, 0.03905512, 0.02675376, 0.007287828, 0.1568716, 
    0.006680343, 0.0008282227, 0.006801853,
  0.0500368, 0.0179688, 0.003830299, 0.1561228, 0.001697528, 0.003873056, 
    0.002380214, 0.0005182119, 0.003010063, 0.003586221, 0.001047205, 
    0.003045795, 0.002537046, 0.000140726, 0.003804479, 0.002215924, 
    0.0001067749, 0.0008087237, 0.000558304, 0.0008068132, 0.003396334, 
    0.02201657, 0.07450512, 0.004917853, 0.01575379, 0.01367199, 
    -0.0003010041, 0.001009534, 0.01498666,
  0.008360609, 0.09621482, 0.01843491, 0.1061082, 0.002782359, 0.003429403, 
    0.001879877, 0.004070279, 0.07177394, 0.04530556, 0.0006894107, 
    0.0007862798, 0.0007503451, 0.001112005, 0.002199043, 0.001591602, 
    0.001302822, 0.002537566, 0.00346534, 0.005424437, 0.01793411, 
    0.07513951, 0.07737607, 0.00931987, 0.001435575, 0.0008091682, 
    0.02177049, 0.001100217, 0.01980142,
  1.855318e-06, -1.544611e-08, 4.561613e-06, 0.005775675, 0.03836076, 
    0.002005085, -0.001802243, 0.001789807, 0.001799744, 0.006346509, 
    0.006374603, 0.0008097357, 0.00197649, 0.003883623, 0.0008739592, 
    0.0005056769, 0.005676622, 0.00494883, 0.01679416, 0.01092443, 
    0.01488391, 0.002188323, 0.1830228, 0.04341898, 0.001028253, 0.001497005, 
    0.001782639, 0.001777972, -1.257617e-07,
  6.91173e-08, 5.192801e-10, 7.300492e-07, 0.001085633, 0.001174185, 
    0.00138015, 0.006617589, 0.0013752, 0.02386976, 0.00477703, 0.002461549, 
    0.002530379, 0.0020077, 0.002420881, 0.0008722055, 0.001067404, 
    0.003856921, 0.00402747, 0.01271253, 0.01329875, 0.004742999, 0.09252967, 
    0.0007068021, 0.001079663, 0.001200116, 0.0009405754, 0.001405152, 
    0.0001744638, 8.508466e-08,
  -2.036251e-05, 0.007964378, 0.000359473, 0.02012524, 0.03603794, 
    0.007632369, -0.0002450175, 0.002644254, 0.07485884, 0.01347266, 
    0.007551852, 0.02530421, 0.02405668, 0.01847254, 0.04046249, 0.01110278, 
    0.01138975, 0.0131236, 0.05110299, 0.01935591, 0.006905825, 0.0494271, 
    0.08087251, 0.009327589, 0.00661805, 0.01953825, 0.0007667181, 
    0.002316839, 0.01265235,
  0.004223479, 0.005256818, 0.03763117, 0.1556615, 0.004720157, 0.001376377, 
    0.1108735, 0.002085557, -7.692131e-05, 0.009060068, 0.1686259, 
    0.03051757, 0.05264252, 0.04974107, 0.07253599, 0.0867293, 0.1347559, 
    0.1291167, 0.08533141, 0.1426032, 0.008451954, 0.07286, 0.1353815, 
    0.06662696, 0.0554872, 0.1014017, 0.09899842, 0.03975692, 0.03565782,
  0.08221506, 0.3142985, 0.2802994, 0.329764, 0.2241002, 0.1285573, 
    0.07394465, 0.1774255, 0.04065299, 0.1374882, 0.06265287, 0.2899019, 
    0.066879, 0.09105687, 0.09517646, 0.1409601, 0.1404112, 0.1782518, 
    0.1728792, 0.4427927, 0.146594, 0.1305532, 0.1831242, 0.5865133, 
    0.1527867, 0.1531647, 0.1342336, 0.1540992, 0.1004338,
  0.04382824, 0.4700314, 0.4011231, 0.6990813, 0.6595023, 0.392139, 
    0.5719131, 0.5525229, 0.5503753, 0.4595854, 0.5216129, 0.4161644, 
    0.158111, 0.2051183, 0.2244335, 0.1798553, 0.3902822, 0.1954021, 
    0.2886707, 0.3702029, 0.6363555, 0.1866642, 0.06638395, 0.306102, 
    0.1056149, 0.09068683, 0.1034576, 0.06594443, 0.06633411,
  0.02103392, 0.01613363, 0.2687264, 0.03718391, 0.1167903, 0.2392325, 
    0.541451, 0.3413485, 0.3653045, 0.5091451, 0.5423501, 0.3700652, 
    0.5034652, 0.5463356, 0.4669801, 0.400044, 0.3106207, 0.3272262, 
    0.3826253, 0.3734012, 0.454654, 0.5889454, 0.3443958, 0.518733, 
    0.07908887, 0.2997838, 0.2907923, 0.09941731, 0.05179185,
  0.4393222, 0.3506702, 0.4360263, 0.3628901, 0.3216701, 0.4917417, 
    0.5611203, 0.5937763, 0.6271101, 0.7040415, 0.6689957, 0.6101357, 
    0.6327984, 0.63267, 0.6301774, 0.5988358, 0.5932439, 0.6709117, 
    0.6576765, 0.6125524, 0.5493035, 0.2691739, 0.3619036, 0.3873887, 
    0.1883363, 0.3199491, 0.1702724, 0.3176221, 0.4881335,
  0.4430829, 0.4487509, 0.4544188, 0.4600868, 0.4657547, 0.4714227, 
    0.4770906, 0.396861, 0.3988021, 0.4007432, 0.4026843, 0.4046254, 
    0.4065664, 0.4085075, 0.5301265, 0.5266436, 0.5231607, 0.5196778, 
    0.5161948, 0.5127119, 0.509229, 0.4824051, 0.478279, 0.4741529, 
    0.4700268, 0.4659007, 0.4617745, 0.4576485, 0.4385486,
  0.101826, 0.1439929, 0.1119697, 0.1653754, 0.2494695, 0.1983509, 0.1970417, 
    0.2052764, 0.1638479, 0.1332218, 0.08094867, 0.0384996, 0.07621513, 
    0.006957516, 0.1895764, 0.2393041, 0.170358, 0.1695509, 0.08090194, 
    0.1021466, 0.1369285, 0.2958013, 0.2360031, 0.06961065, 0.0663705, 
    0.1429054, 0.01927013, 0.03937092, 0.07698083,
  0.1015999, 0.06153607, 0.07941607, 0.04494298, 0.06222683, 0.1381198, 
    0.01583753, 0.04060267, 0.0745022, 0.07660588, 0.05394554, 0.04891646, 
    0.03898134, 0.08985268, 0.2153571, 0.2257122, 0.1927871, 0.1857137, 
    0.2410624, 0.182337, 0.2003926, 0.1798826, 0.1980385, 0.3377196, 
    0.05350696, 0.2135036, 0.2136506, 0.1864333, 0.1883027,
  0.201085, 0.1813124, 0.2163672, 0.1799963, 0.1959352, 0.1911732, 0.1870813, 
    0.1802312, 0.2152888, 0.1561689, 0.1694023, 0.1881038, 0.224631, 
    0.1872844, 0.1894724, 0.2738055, 0.3101558, 0.3042896, 0.2389219, 
    0.1870707, 0.1616442, 0.1253515, 0.1249305, 0.1689231, 0.2121511, 
    0.315845, 0.3240837, 0.2805636, 0.2364336,
  0.242658, 0.1980882, 0.1981247, 0.1548137, 0.1421007, 0.140299, 0.173748, 
    0.1302165, 0.1662552, 0.1839443, 0.09642871, 0.1022666, 0.03947319, 
    0.09603523, 0.1502072, 0.140566, 0.1269284, 0.1307707, 0.1594695, 
    0.1280203, 0.1185264, 0.187198, 0.1298299, 0.07078291, 0.07029422, 
    0.2181133, 0.2949406, 0.2478126, 0.2888435,
  0.07871428, 0.01991796, 0.01098375, 0.07347678, 0.06629943, 0.05739396, 
    0.0666339, 0.08555938, 0.0874446, 0.04372929, 0.02864455, 0.007572779, 
    0.009741532, 0.09051913, 0.1818718, 0.1137681, 0.1315617, 0.1145738, 
    0.1046877, 0.1139392, 0.1837014, 0.1201622, 0.0776979, 0.09962012, 
    0.03204358, 0.09859123, 0.08633927, 0.1284358, 0.1168005,
  0.008254549, 0.009403221, 0.00770419, 0.0413691, 0.03264261, 0.005797906, 
    0.00816124, 0.00846573, 0.02873018, 0.01851217, 4.137451e-05, 
    1.597126e-07, 0.001110833, 0.02012508, 0.01558005, 0.01563124, 
    0.009125462, 0.01779351, 0.05649976, 0.02962131, 0.02016232, 0.002161146, 
    0.01614719, 0.02271833, 0.00277142, 0.01148334, 0.02883654, 0.008277448, 
    0.004253666,
  0.01473306, 0.0154939, 0.002589943, 0.002579376, -0.0005296163, 
    0.001377283, 0.001459808, 0.00345797, 0.01648161, -1.078606e-05, 
    6.048209e-08, -2.074575e-06, 0.003259691, 0.001270863, 0.002803814, 
    0.00320437, 0.001015211, 0.004040473, 0.002147768, 0.002716596, 
    0.0007311186, 0.004086112, 0.0244422, 0.01720112, 0.004996931, 0.1278744, 
    0.002471962, 0.0005327863, 0.003862043,
  0.03172177, 0.007940128, 0.003267694, 0.1184676, 0.000930434, 0.001544101, 
    0.001043867, 0.0002718134, 0.001903942, 0.002470208, 0.0004910598, 
    0.001604122, 0.001030239, 5.697389e-05, 0.002033499, 0.0009279515, 
    8.97896e-05, 0.0005298767, 0.0003708745, 0.0005387745, 0.002236464, 
    0.01422757, 0.04669661, 0.00573915, 0.01174278, 0.01164715, 1.989025e-05, 
    0.0006154048, 0.009368462,
  0.00314744, 0.08163403, 0.01681733, 0.0857996, 0.001696584, 0.001690061, 
    0.001148187, 0.002545833, 0.06635105, 0.04679295, 0.000329613, 
    0.0004676743, 0.0004717202, 0.0005040453, 0.001310259, 0.0009056866, 
    0.0008372525, 0.001599922, 0.002128864, 0.003049766, 0.009745616, 
    0.04345511, 0.04700631, 0.01018107, 0.001662428, 0.0004280557, 
    0.01021286, 0.0003715214, 0.008075885,
  -1.457499e-06, -7.162545e-08, 1.989962e-06, 0.006348442, 0.02480428, 
    0.001273397, -0.001604997, 0.000618833, 0.0006460929, 0.002399225, 
    0.002673828, 0.0003438883, 0.0008453474, 0.001532458, 0.0003281665, 
    0.0002236584, 0.00280885, 0.001894018, 0.007156114, 0.004810559, 
    0.005626324, 0.001123672, 0.1328864, 0.03995766, 0.0004707109, 
    0.0006801609, 0.0009787192, 0.00115769, -1.684745e-06,
  6.692903e-08, 5.184945e-10, 6.617364e-07, 0.0006612057, 0.0004080639, 
    0.0009414227, 0.008386141, 0.0009459711, 0.01589887, 0.002778958, 
    0.001067907, 0.001186762, 0.0009903363, 0.0009365326, 0.0005401157, 
    0.000709738, 0.001952089, 0.001997711, 0.007331511, 0.008706152, 
    0.002745559, 0.06910418, 0.0004724799, -0.000511999, 0.0007764131, 
    0.0005260165, 0.0009497963, 0.0001039922, 8.640252e-08,
  -2.152781e-05, 0.00419959, 0.0003940932, 0.013962, 0.02619129, 0.005262296, 
    -0.000311892, 0.005795497, 0.06546497, 0.008410334, 0.005553265, 
    0.01362155, 0.01069703, 0.007372614, 0.01980745, 0.005056524, 
    0.005537238, 0.005036261, 0.02645985, 0.01352049, 0.005093704, 
    0.04382014, 0.06863463, 0.002913032, 0.002793587, 0.009148898, 
    0.0004481591, 0.001647921, 0.009495756,
  0.002639164, 0.002816394, 0.02353665, 0.1475321, 0.002780987, 0.0009080691, 
    0.0958918, 0.001681811, -5.306085e-05, 0.007112225, 0.15069, 0.02171031, 
    0.0381404, 0.03373998, 0.04841466, 0.0620947, 0.1005084, 0.09217023, 
    0.04830782, 0.1313961, 0.007200575, 0.06424019, 0.1133307, 0.05200073, 
    0.03251592, 0.06055434, 0.06075696, 0.02077774, 0.02304115,
  0.05339234, 0.2651169, 0.2239722, 0.2706402, 0.1878789, 0.1133853, 
    0.05692376, 0.1519516, 0.04181627, 0.1129399, 0.05523517, 0.2612612, 
    0.05214309, 0.06686999, 0.07032323, 0.1015138, 0.09977903, 0.1285615, 
    0.1155393, 0.421704, 0.1231912, 0.1011669, 0.1357051, 0.5117139, 
    0.1246288, 0.1317385, 0.09981802, 0.1037342, 0.06861314,
  0.02718949, 0.457891, 0.365116, 0.6236914, 0.6008805, 0.3543847, 0.4990134, 
    0.4690487, 0.4682212, 0.3914538, 0.4343789, 0.4206508, 0.1949978, 
    0.2019947, 0.189083, 0.1345875, 0.4055439, 0.1553971, 0.2388115, 
    0.3400533, 0.6088684, 0.1541229, 0.04754928, 0.3290451, 0.08196582, 
    0.07580986, 0.07295647, 0.04413488, 0.04421793,
  0.01480522, 0.009960163, 0.2767528, 0.02605717, 0.089212, 0.1970373, 
    0.4771407, 0.315137, 0.3414963, 0.4816577, 0.5624021, 0.3358577, 
    0.5152822, 0.422928, 0.3680782, 0.3445399, 0.281718, 0.2489359, 
    0.3667606, 0.2822976, 0.373427, 0.6158463, 0.325007, 0.5600848, 
    0.0639448, 0.2722617, 0.3441135, 0.07824224, 0.03975538,
  0.4517927, 0.3337802, 0.4583157, 0.3675917, 0.3889325, 0.4727884, 0.530009, 
    0.5802624, 0.5844434, 0.638317, 0.6825696, 0.6103629, 0.6053241, 
    0.5801957, 0.5149739, 0.604404, 0.5271579, 0.5832021, 0.5869421, 
    0.6140814, 0.5667929, 0.289083, 0.4133685, 0.476545, 0.1710498, 
    0.2874725, 0.1611949, 0.3148034, 0.488014,
  0.3267463, 0.3320991, 0.3374518, 0.3428046, 0.3481573, 0.3535101, 
    0.3588629, 0.2699016, 0.2703467, 0.2707918, 0.271237, 0.2716821, 
    0.2721272, 0.2725723, 0.3923752, 0.3893393, 0.3863033, 0.3832674, 
    0.3802314, 0.3771955, 0.3741595, 0.3456641, 0.3429022, 0.3401403, 
    0.3373784, 0.3346164, 0.3318545, 0.3290926, 0.3224641,
  0.09289858, 0.1107737, 0.08461954, 0.1341361, 0.2259889, 0.1666136, 
    0.1464667, 0.1603117, 0.1165281, 0.09011409, 0.05323497, 0.02384339, 
    0.059299, 0.006267394, 0.2130611, 0.2166228, 0.1517762, 0.1574819, 
    0.06861477, 0.1070621, 0.1127784, 0.2591559, 0.2004867, 0.05973397, 
    0.07564279, 0.1341403, 0.0165168, 0.03292689, 0.06983186,
  0.09782998, 0.05708093, 0.08123255, 0.03815696, 0.05005676, 0.1176008, 
    0.01297798, 0.03245836, 0.06349927, 0.05772665, 0.04569394, 0.04314125, 
    0.02932986, 0.08027677, 0.1912234, 0.1911618, 0.1555992, 0.158951, 
    0.1894218, 0.1535534, 0.1600155, 0.1377943, 0.1580679, 0.2798682, 
    0.04528492, 0.1692641, 0.1737939, 0.1478796, 0.152223,
  0.1558049, 0.1431212, 0.1726855, 0.1415726, 0.1514051, 0.1513226, 
    0.1453948, 0.1383332, 0.167602, 0.1254711, 0.135024, 0.152535, 0.1795191, 
    0.1533611, 0.1493503, 0.2226376, 0.2578741, 0.2587174, 0.196838, 
    0.1501468, 0.1293347, 0.09556971, 0.09133202, 0.1246993, 0.1719754, 
    0.2556982, 0.2672958, 0.2271697, 0.1882932,
  0.2010263, 0.1591206, 0.1619504, 0.1206241, 0.110925, 0.1185591, 0.1370286, 
    0.09793782, 0.1247392, 0.1377706, 0.06769183, 0.07013743, 0.0256964, 
    0.06688079, 0.1110358, 0.09906079, 0.08849438, 0.09110638, 0.1159967, 
    0.08552285, 0.08197542, 0.1382953, 0.09096881, 0.06124815, 0.05254197, 
    0.1728332, 0.2462565, 0.1982692, 0.2435232,
  0.05110062, 0.0126188, 0.007222492, 0.04699025, 0.04166483, 0.03928961, 
    0.04119269, 0.05782698, 0.05673226, 0.02629369, 0.01784415, 0.005646722, 
    0.007153627, 0.06410861, 0.158769, 0.07463998, 0.09937507, 0.07586361, 
    0.07333795, 0.08843581, 0.1340857, 0.08513101, 0.05145727, 0.08586006, 
    0.03233106, 0.07154633, 0.0541901, 0.09038574, 0.07810672,
  0.006467939, 0.007003997, 0.005504995, 0.02327459, 0.01870161, 0.003363397, 
    0.005028669, 0.005329644, 0.02078997, 0.01478062, 2.136755e-05, 
    1.297678e-07, 0.0003346484, 0.01209051, 0.008078102, 0.009233426, 
    0.00528266, 0.009814324, 0.03486189, 0.01774752, 0.01093144, 0.001592751, 
    0.01175736, 0.01839419, 0.002061668, 0.006068175, 0.01533671, 
    0.005982344, 0.003342455,
  0.01063609, 0.01112723, 0.001379103, 0.001776004, -0.0003482445, 
    0.0008657841, 0.001008224, 0.00245538, 0.01189252, -9.134505e-06, 
    5.671721e-08, -3.581142e-07, 0.002300418, 0.0008481344, 0.001408321, 
    0.001784823, 0.0006472393, 0.002124772, 0.001094627, 0.001319888, 
    0.000510855, 0.003014085, 0.01757746, 0.01286579, 0.003560274, 0.103741, 
    0.001051456, 0.0003925471, 0.002617727,
  0.02322131, 0.003849097, 0.004594302, 0.09780961, 0.0006414519, 
    0.0006897631, 0.0005520022, 0.0001916907, 0.001383889, 0.001867747, 
    0.0003281969, 0.0009019896, 0.0006608571, 6.400645e-05, 0.001011563, 
    0.0005055865, 7.360586e-05, 0.0003946197, 0.0002776115, 0.0004047954, 
    0.001666991, 0.01048993, 0.03395925, 0.007043209, 0.009298319, 
    0.008837679, 8.822513e-05, 0.0004402957, 0.006804631,
  0.001500672, 0.06866327, 0.01057082, 0.07391927, 0.001178867, 0.00107916, 
    0.0008266635, 0.001823549, 0.0647929, 0.04971654, 0.0002112881, 
    0.0003285696, 0.0003386479, 0.0003342531, 0.0009261904, 0.0006104876, 
    0.0006150987, 0.001158186, 0.001524685, 0.002070874, 0.006506108, 
    0.03030114, 0.03340336, 0.007560001, 0.001832211, 0.0002875083, 
    0.004616642, 0.0001710191, 0.003260805,
  -5.517477e-07, -4.386212e-06, 3.856365e-07, 0.00808073, 0.01972603, 
    0.0009471941, -0.001179634, 0.0003066116, 0.000417819, 0.001092138, 
    0.001261271, 0.000213091, 0.0004570788, 0.0008326569, 0.0001739323, 
    0.0001470792, 0.001382095, 0.00101467, 0.003340347, 0.002141296, 
    0.002342385, 0.0007629268, 0.108043, 0.0339522, 0.0002613578, 
    0.0003498618, 0.0006565818, 0.000856644, -1.96715e-05,
  6.57652e-08, 5.224004e-10, 5.865289e-07, 0.0003548741, 0.0001743516, 
    0.0007080235, 0.01143969, 0.0007120605, 0.01211387, 0.001900871, 
    0.0006317209, 0.0007517769, 0.0006183943, 0.000491723, 0.0003940858, 
    0.0005380915, 0.001145025, 0.001330815, 0.005202752, 0.006607377, 
    0.001804581, 0.05805766, 0.0003661409, -0.0008229914, 0.0005746273, 
    0.0003469382, 0.0007187987, 7.730927e-05, 8.613618e-08,
  -1.738336e-05, 0.002941823, 0.000140606, 0.0109887, 0.01959418, 
    0.003279551, -0.0005700538, 0.00802175, 0.0637563, 0.006559485, 
    0.004504795, 0.008378942, 0.005307969, 0.003788156, 0.009933714, 
    0.002817241, 0.003428006, 0.002361976, 0.01495559, 0.0095545, 
    0.003953839, 0.04244613, 0.05853294, 0.001728811, 0.001661216, 
    0.004347248, 0.0003269863, 0.001285063, 0.007825724,
  0.003161102, 0.001724087, 0.0151755, 0.1399078, 0.00198894, 0.0006185912, 
    0.0896225, 0.001106509, -3.764679e-05, 0.005476831, 0.1349499, 
    0.01701086, 0.02706648, 0.02245446, 0.03015603, 0.04223944, 0.0762623, 
    0.05817756, 0.03054588, 0.1201276, 0.00598062, 0.05959278, 0.09605341, 
    0.0419849, 0.01998363, 0.03471812, 0.03204566, 0.01194073, 0.01639067,
  0.03765715, 0.2330911, 0.1919481, 0.2332043, 0.1619966, 0.1053675, 
    0.04848146, 0.1444564, 0.05876261, 0.09666084, 0.04915077, 0.2526759, 
    0.04151466, 0.0542644, 0.05375337, 0.07339732, 0.07269929, 0.09092508, 
    0.07938245, 0.4090649, 0.1077519, 0.07929856, 0.1135115, 0.4493163, 
    0.1051538, 0.1156333, 0.07630456, 0.06967232, 0.04585207,
  0.01923336, 0.4211115, 0.3373781, 0.5534322, 0.5594519, 0.3229771, 
    0.4484888, 0.4138703, 0.4009202, 0.3281425, 0.3580634, 0.4400614, 
    0.2402441, 0.2149396, 0.1614948, 0.1071612, 0.4072553, 0.1409278, 
    0.2118764, 0.3135859, 0.5528608, 0.1487389, 0.03788003, 0.3562213, 
    0.07008402, 0.06522356, 0.0560292, 0.03210769, 0.03224776,
  0.01090936, 0.007284683, 0.3108526, 0.02016526, 0.07262985, 0.1604826, 
    0.4286838, 0.3266652, 0.3397353, 0.4405437, 0.5614969, 0.3067504, 
    0.4558522, 0.3237023, 0.2832919, 0.2893984, 0.2613961, 0.1998911, 
    0.3032959, 0.2168774, 0.2716924, 0.5368749, 0.3395811, 0.5762204, 
    0.05269269, 0.2514658, 0.4323809, 0.06279044, 0.03185373,
  0.4692232, 0.3206043, 0.4468362, 0.3400627, 0.3615684, 0.3973252, 
    0.4221947, 0.4497923, 0.445039, 0.4750656, 0.4767813, 0.4055793, 
    0.4103283, 0.4191252, 0.3617086, 0.4255057, 0.3869942, 0.4368163, 
    0.409879, 0.4082022, 0.4049399, 0.2866455, 0.4302759, 0.5677292, 
    0.172438, 0.2493077, 0.1726852, 0.2994722, 0.4173578,
  0.2128464, 0.2166433, 0.2204402, 0.2242371, 0.2280341, 0.231831, 0.2356279, 
    0.1905023, 0.1917098, 0.1929172, 0.1941246, 0.195332, 0.1965394, 
    0.1977468, 0.269731, 0.2673698, 0.2650087, 0.2626476, 0.2602865, 
    0.2579254, 0.2555643, 0.2666344, 0.2639912, 0.261348, 0.2587048, 
    0.2560616, 0.2534183, 0.2507751, 0.2098089,
  0.1059392, 0.098052, 0.07207775, 0.1158308, 0.2018186, 0.1363353, 
    0.1285619, 0.148889, 0.09238175, 0.06969389, 0.04245215, 0.01828593, 
    0.04485846, 0.006338859, 0.2452876, 0.2028243, 0.1600949, 0.1663072, 
    0.06411521, 0.1242283, 0.1065908, 0.230909, 0.1760156, 0.06063301, 
    0.09760183, 0.1287406, 0.02616319, 0.03084959, 0.06375111,
  0.09623244, 0.06948148, 0.09898067, 0.03389095, 0.04784286, 0.1090773, 
    0.01315206, 0.02839141, 0.05703623, 0.05043416, 0.04088669, 0.04600859, 
    0.02638295, 0.07895287, 0.1904521, 0.1762841, 0.1362111, 0.143992, 
    0.1653968, 0.1318158, 0.1428789, 0.1196256, 0.1397957, 0.2474619, 
    0.0406546, 0.1493214, 0.1544347, 0.1283379, 0.1312932,
  0.1354037, 0.1271286, 0.1503784, 0.1237795, 0.1274111, 0.127808, 0.1214, 
    0.1185276, 0.1421438, 0.1081359, 0.1168556, 0.1313314, 0.1486866, 
    0.1308643, 0.1258542, 0.189161, 0.2206748, 0.2266012, 0.1715305, 
    0.1270573, 0.1098007, 0.08044538, 0.07498217, 0.1020963, 0.1414479, 
    0.2188921, 0.2378331, 0.1999324, 0.1644843,
  0.1733651, 0.1371002, 0.1366097, 0.101286, 0.09423018, 0.1028511, 
    0.1119725, 0.08066477, 0.1028163, 0.1129244, 0.05285172, 0.05308734, 
    0.01831069, 0.05206622, 0.08861314, 0.07582651, 0.06520816, 0.06820816, 
    0.09004339, 0.06349969, 0.06399766, 0.107537, 0.07246664, 0.06362177, 
    0.03955242, 0.1369798, 0.2066992, 0.166852, 0.2090986,
  0.03861114, 0.009632777, 0.005137896, 0.03226783, 0.02946714, 0.02795812, 
    0.02786563, 0.0434531, 0.03873888, 0.01882562, 0.01296247, 0.004759937, 
    0.005386699, 0.04696928, 0.1681221, 0.05272094, 0.07106449, 0.05220189, 
    0.05488588, 0.06565872, 0.1001252, 0.06211542, 0.03840757, 0.07994176, 
    0.02857873, 0.05079721, 0.03734374, 0.066329, 0.05655873,
  0.005538297, 0.00586962, 0.01131314, 0.01653307, 0.01168829, 0.002562179, 
    0.003755617, 0.004066954, 0.01483235, 0.01260061, 1.425624e-05, 
    1.148355e-07, 0.002521505, 0.008748466, 0.004657389, 0.005925518, 
    0.003378997, 0.006322883, 0.02236955, 0.01175646, 0.006395269, 
    0.001317491, 0.009749288, 0.01631559, 0.00192511, 0.003816386, 
    0.009671128, 0.003899244, 0.002832134,
  0.008741877, 0.008359486, 0.0007993355, 0.001376387, -0.0004064832, 
    0.0006828627, 0.0007848406, 0.00199019, 0.009679427, -7.876517e-06, 
    5.615131e-08, -5.708372e-08, 0.001845332, 0.0006896133, 0.0009552443, 
    0.001276761, 0.0005046434, 0.001510598, 0.0007582092, 0.0008143811, 
    0.0004120863, 0.00251334, 0.01439591, 0.01052919, 0.009628769, 0.1291037, 
    0.0006985702, 0.0003273332, 0.002095021,
  0.01904218, 0.002114741, 0.02004927, 0.1238829, 0.0005113414, 0.0004379365, 
    0.0003905334, 0.0001597187, 0.001138571, 0.001254088, 0.0002609915, 
    0.0006156124, 0.0004512301, 6.208084e-05, 0.0006568859, 0.0003529773, 
    6.226885e-05, 0.0003259355, 0.0002309822, 0.000339006, 0.00139351, 
    0.008686573, 0.02772191, 0.03596154, 0.01805111, 0.008119066, 
    9.943819e-05, 0.0003623904, 0.005592855,
  0.001022696, 0.08684957, 0.01150708, 0.07531323, 0.0009410483, 
    0.0008213097, 0.0006660273, 0.001475196, 0.08981119, 0.07721926, 
    0.0001691216, 0.000261455, 0.0002651406, 0.0002622716, 0.0007396424, 
    0.0004960612, 0.0005072248, 0.0009455368, 0.001229489, 0.001637449, 
    0.005057454, 0.02404746, 0.02684259, 0.04153452, 0.02402439, 
    0.0002247461, 0.002694749, 0.0001160263, 0.001845682,
  -2.410425e-05, -5.508396e-05, -1.273903e-07, 0.01608139, 0.01564826, 
    0.0007890009, -0.001390425, 0.0002112366, -1.722125e-05, 0.0007478521, 
    0.0007817182, 0.0001657003, 0.0003172448, 0.0005992158, 0.0001325344, 
    0.0001169358, 0.0009093729, 0.0007455309, 0.001994915, 0.001255874, 
    0.00145098, 0.0006078333, 0.1450295, 0.03265353, 0.0002020041, 
    0.0002589185, 0.0005029125, 0.000705555, -7.741697e-05,
  6.588785e-08, 5.320347e-10, -6.415276e-08, 0.0002313409, 0.0001004993, 
    0.0005853871, 0.01441962, 0.0005309301, 0.01178075, 0.001218289, 
    0.0005110453, 0.0006008575, 0.000476714, 0.0003544715, 0.0003246191, 
    0.0004517519, 0.0008422998, 0.001058181, 0.004232391, 0.005521099, 
    0.001422959, 0.05468452, 0.0003141421, -0.001235785, 0.0004693196, 
    0.0002682684, 0.0006053424, 6.515585e-05, 8.716507e-08,
  -1.372968e-05, 0.002426057, 0.0003179469, 0.01065719, 0.01844934, 
    0.003681997, 0.001011968, 0.01333662, 0.06927608, 0.007384009, 
    0.003966616, 0.006117264, 0.003529662, 0.002649438, 0.00554911, 
    0.001942201, 0.002637912, 0.001534325, 0.009625781, 0.007128765, 
    0.00310734, 0.04629205, 0.06696758, 0.001452999, 0.001267589, 
    0.002837266, 0.0002713388, 0.001077671, 0.008099026,
  0.004167296, 0.0008581337, 0.01108109, 0.1407932, 0.001591367, 
    0.0005186662, 0.08480191, 0.0008360443, -3.660032e-05, 0.004634986, 
    0.1435605, 0.01489458, 0.02192362, 0.01720355, 0.02213513, 0.03113817, 
    0.05938305, 0.04086477, 0.02200485, 0.1155081, 0.004752863, 0.05833346, 
    0.100845, 0.03483283, 0.01443648, 0.02383563, 0.0178536, 0.008512933, 
    0.01386396,
  0.02846352, 0.2379571, 0.1904137, 0.23588, 0.1539291, 0.1053922, 
    0.04611517, 0.2072437, 0.09526714, 0.09599952, 0.06787542, 0.2795959, 
    0.03618741, 0.04866844, 0.0450992, 0.05880224, 0.05701677, 0.071022, 
    0.05945177, 0.43291, 0.1044548, 0.0733799, 0.1293594, 0.4458643, 
    0.1010341, 0.09907073, 0.06220895, 0.05346479, 0.03310538,
  0.01538502, 0.4321544, 0.3287627, 0.5314441, 0.5544928, 0.3601449, 
    0.4520952, 0.4284737, 0.3834875, 0.3126374, 0.3381446, 0.5193986, 
    0.3367136, 0.2580802, 0.1462401, 0.09281883, 0.4321353, 0.1412139, 
    0.2445926, 0.3349971, 0.538146, 0.1663112, 0.03339414, 0.4069262, 
    0.06286101, 0.05977746, 0.04747989, 0.02661993, 0.02689107,
  0.009026401, 0.006125784, 0.3631184, 0.01658184, 0.06379717, 0.1397499, 
    0.4025908, 0.349808, 0.3791965, 0.4404498, 0.6178308, 0.3441011, 
    0.4495798, 0.2649727, 0.2449035, 0.2639917, 0.2966475, 0.1783079, 
    0.2638293, 0.183855, 0.2226241, 0.4777764, 0.3315459, 0.5681455, 
    0.04696926, 0.2274182, 0.5162534, 0.05673754, 0.02740966,
  0.4800027, 0.31591, 0.4003987, 0.2675982, 0.3107324, 0.323075, 0.3235577, 
    0.3423087, 0.33815, 0.3409396, 0.3264423, 0.2863331, 0.2934329, 
    0.3184902, 0.260287, 0.3240471, 0.2955882, 0.3298383, 0.3152619, 
    0.3071314, 0.3036175, 0.2989596, 0.4720376, 0.6256486, 0.173578, 
    0.2263957, 0.1944792, 0.3079453, 0.3605 ;

 average_DT = 730 ;

 average_T1 = 320 ;

 average_T2 = 1050 ;

 climatology_bounds =
  320, 1050 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
