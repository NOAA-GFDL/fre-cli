netcdf \00010101.river_month.tile1.rv_o_h2o {
dimensions:
	time = UNLIMITED ; // (12 currently)
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float rv_o_h2o(time, grid_yt, grid_xt) ;
		rv_o_h2o:_FillValue = -1.e+08f ;
		rv_o_h2o:missing_value = -1.e+08f ;
		rv_o_h2o:units = "kg/m2/s" ;
		rv_o_h2o:long_name = "river outflow, h2o mass" ;
		rv_o_h2o:cell_methods = "time: mean" ;
		rv_o_h2o:time_avg_info = "average_T1,average_T2,average_DT" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "areacellr: 00010101.river_static_cmip.nc land_area: 00010101.river_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Sep  5 12:38:46 2025: ncatted -O -a coordinates,,d,, /work/cew/scratch/workflow-test/river_month//split-netcdf//00010101.river_month.tile1.rv_o_h2o.nc\nFri Sep  5 12:38:28 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 /work/cew/scratch//00010101.river_month.tile1.nc -O /work/cew/scratch/workflow-test/river_month//ncks_out//00010101.river_month.tile1.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365 ;

 rv_o_h2o =
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.783949e-12, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.754725e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  5.370085e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  8.173346e-08, 6.418787e-13, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.141853e-08, 3.706681e-07, 2.288766e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.55106e-08, 1.047896e-07, 1.18621e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  3.458532e-06, 1.852095e-06, 1.069637e-05, 1.142035e-11, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  2.319162e-06, 2.64238e-06, 7.163104e-07, 5.245058e-06, 2.825562e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.453269e-12, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.43408e-08, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  5.179931e-08, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.366156e-06, 1.778598e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  5.885338e-08, 3.200078e-07, 6.965727e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.517018e-08, 4.57346e-07, 4.334787e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  3.46297e-06, 1.661024e-06, 9.343751e-06, 9.460297e-12, 0, 0, _, _, _, _, _, 
    _, _, _, _,
  1.700426e-06, 1.932523e-06, 3.435822e-07, 4.441563e-06, 5.817318e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.173501e-12, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.692413e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  3.34457e-08, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.527236e-08, 7.696157e-09, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.246274e-09, 3.458272e-07, 2.424648e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.159908e-09, 1.12311e-08, 8.695477e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.930972e-06, 1.839331e-06, 9.74838e-06, 7.929491e-12, 0, 0, _, _, _, _, _, 
    _, _, _, _,
  1.871002e-06, 2.437646e-06, 9.614423e-07, 4.835775e-06, 4.858274e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.926663e-12, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.350512e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  3.988207e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.67404e-07, 1.50401e-09, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.115685e-07, 4.065391e-07, 1.591828e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  8.011843e-08, 1.521109e-07, 1.210448e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  4.154814e-06, 1.869857e-06, 1.159446e-05, 4.058029e-08, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  2.144441e-06, 2.980537e-06, 1.350278e-06, 4.7859e-06, 8.845695e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.026505e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.632753e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  3.256443e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.841992e-08, 5.396015e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.841604e-08, 3.584104e-07, 1.044741e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.01403e-09, 8.954152e-08, 8.094626e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.763084e-06, 1.780599e-06, 9.088204e-06, 8.32863e-08, 0, 0, _, _, _, _, _, 
    _, _, _, _,
  1.664419e-06, 2.136979e-06, 6.021688e-07, 4.00265e-06, 9.128241e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9.614267e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.218107e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  1.622921e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.19915e-08, 2.519898e-10, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.239342e-08, 3.44725e-07, 6.766038e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.545081e-10, 1.041748e-07, 8.21075e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.708135e-06, 1.781257e-06, 8.726299e-06, 1.285764e-07, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  1.551048e-06, 2.080922e-06, 6.336949e-07, 3.797761e-06, 9.355174e-07, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.852475e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.580138e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  6.055403e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  8.716285e-08, 2.272584e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.882848e-08, 4.290145e-07, 1.862803e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.674542e-08, 2.995227e-07, 1.091762e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.869512e-06, 1.837604e-06, 9.349597e-06, 5.134834e-08, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  1.687709e-06, 2.375356e-06, 7.590771e-07, 3.743873e-06, 1.018836e-06, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.095259e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.963832e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  1.621293e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.675391e-08, 1.721222e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.268218e-08, 4.572776e-07, 2.772999e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  8.107595e-08, 1.656344e-06, 1.600403e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.765611e-06, 1.880544e-06, 1.059338e-05, 2.771205e-07, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  1.48227e-06, 2.182951e-06, 7.748583e-07, 3.688564e-06, 1.051489e-06, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.174346e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.164013e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  3.133352e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.43002e-07, 5.891942e-09, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.248717e-08, 4.69442e-07, 1.027973e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.680072e-09, 7.870566e-07, 1.875703e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.897054e-06, 1.883745e-06, 1.08927e-05, 4.610299e-07, 0, 0, _, _, _, _, _, 
    _, _, _, _,
  1.669194e-06, 2.538543e-06, 1.194217e-06, 3.890069e-06, 1.807028e-06, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.721434e-08, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.064937e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  6.363212e-07, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.289753e-07, 5.0667e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.019959e-09, 4.363419e-07, 7.853914e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.736772e-10, 1.900696e-07, 1.292923e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.703483e-06, 1.794684e-06, 8.022034e-06, 2.409837e-07, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  1.235817e-06, 1.856054e-06, 5.498907e-07, 3.000923e-06, 1.190648e-06, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.272583e-09, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.965654e-07, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  6.276038e-09, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.071777e-07, 7.580739e-09, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  8.926763e-10, 4.787742e-07, 1.098006e-06, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.067065e-10, 2.155925e-07, 1.313095e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.759327e-06, 1.844869e-06, 8.094425e-06, 1.954345e-07, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  1.204259e-06, 1.885949e-06, 6.692941e-07, 3.164022e-06, 1.472084e-06, 0, 0, 
    _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.103318e-09, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.467109e-08, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  1.192214e-09, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.654616e-07, 1.46936e-09, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.365767e-10, 4.750335e-07, 2.507245e-07, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.486241e-11, 2.445026e-08, 1.107022e-06, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  2.938859e-06, 1.955711e-06, 8.338474e-06, 7.487669e-08, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  2.16795e-06, 2.650416e-06, 9.170484e-07, 3.098445e-06, 4.559905e-07, 0, 0, 
    _, _, _, _, _, _, _, _ ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 349.5 ;
}
