netcdf atmos.1980-1981.alb_sfc.09 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:21 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.09.nc reduced/atmos.1980-1981.alb_sfc.09.nc\n",
			"Mon Aug 25 14:40:08 2025: cdo -O -s -select,month=9 merged_output.nc monthly_nc_files/all_years.9.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  20.66323, 20.66323, 20.66323, 20.66323, 20.66323, 20.66323, 20.66323, 
    20.58856, 20.58856, 20.58856, 20.58856, 20.58856, 20.58856, 20.58856, 
    20.42933, 20.42933, 20.42933, 20.42933, 20.42933, 20.42933, 20.42933, 
    20.50862, 20.50862, 20.50862, 20.50862, 20.50862, 20.50862, 20.50862, 
    20.66323,
  33.02045, 32.92193, 32.90263, 32.77621, 32.72767, 32.66845, 32.67631, 
    32.75317, 32.767, 32.90293, 33.0189, 33.04833, 33.10769, 33.17324, 
    33.20422, 33.50983, 33.3208, 33.29965, 33.11493, 33.10618, 33.10583, 
    33.1887, 33.19465, 33.51388, 33.49552, 33.51531, 33.67562, 33.36684, 
    33.15046,
  41.52293, 41.56403, 43.09171, 40.14873, 36.54132, 36.48971, 39.89568, 
    36.53849, 36.59326, 36.70491, 36.67489, 36.64999, 36.98787, 42.9565, 
    43.18962, 42.5639, 42.39352, 42.70868, 42.23248, 42.04861, 41.74931, 
    40.74972, 40.7514, 38.72163, 42.57952, 43.20123, 43.29587, 43.36191, 
    43.28548,
  43.47955, 43.76934, 8.859238, 4.225399, 7.922081, 16.25109, 42.78152, 
    25.71103, 20.68662, 4.543509, 4.446462, 4.362767, 4.021481, 4.105857, 
    4.296268, 4.016517, 3.859648, 3.656593, 4.020806, 4.266135, 4.194271, 
    4.23074, 4.13394, 4.034355, 14.59998, 29.85413, 38.79991, 40.99497, 
    42.7914,
  3.821842, 3.864328, 3.901444, 3.807488, 3.908346, 3.907754, 3.877761, 
    4.045282, 4.073135, 4.069674, 4.01515, 3.977728, 3.95337, 3.968427, 
    3.900409, 3.924134, 3.833704, 3.729463, 3.886237, 3.800952, 3.881865, 
    3.961741, 3.800235, 8.401329, 4.224381, 3.80261, 3.698251, 3.578206, 
    3.723454,
  3.702379, 3.745209, 3.78032, 3.594174, 3.612713, 3.710622, 3.736301, 
    3.883488, 3.752656, 3.95553, 3.802466, 3.977048, 4.063, 3.807789, 
    13.84426, 3.726971, 3.955099, 3.754842, 3.629945, 3.779317, 3.845484, 
    3.894812, 3.833145, 10.97887, 4.332592, 3.895722, 3.646708, 3.734929, 
    3.590675,
  3.665452, 3.735859, 12.73534, 3.612913, 3.733438, 3.65388, 3.774567, 
    3.835169, 3.747289, 4.112978, 9.480423, 14.10804, 11.43204, 3.790099, 
    3.693535, 3.621714, 3.723859, 3.597898, 3.343357, 3.472167, 3.754168, 
    3.656986, 3.566717, 4.528167, 8.841412, 3.518774, 3.568186, 3.53184, 
    3.608103,
  3.277508, 9.679306, 10.09781, 3.733357, 3.746872, 3.756079, 3.624061, 
    3.636028, 3.657395, 3.829741, 11.92314, 11.70178, 3.708552, 3.591596, 
    3.556084, 3.456469, 3.582799, 3.688466, 3.756582, 3.830585, 3.564949, 
    3.267758, 3.276315, 3.593744, 8.917823, 9.045326, 3.799617, 3.687589, 
    3.493907,
  3.080974, 6.082598, 9.040388, 9.105547, 3.624725, 3.591949, 3.273056, 
    3.299476, 3.43743, 3.508, 4.743412, 3.44821, 4.20923, 3.245314, 3.289592, 
    3.342466, 3.563619, 3.773612, 3.63663, 3.732333, 3.568008, 3.268701, 
    3.325814, 8.741015, 8.591301, 12.00813, 3.721806, 3.416591, 3.239951,
  3.206051, 8.170681, 8.205413, 9.928078, 3.454987, 3.238625, 3.109753, 
    3.076408, 8.55699, 8.239193, 3.310597, 3.374115, 3.356166, 3.472544, 
    3.505334, 3.541268, 3.566093, 3.742085, 3.510695, 3.540003, 3.386259, 
    3.177172, 3.173014, 8.476091, 8.579597, 3.423398, 3.421369, 3.29805, 
    3.153507,
  9.535032, 9.799501, 9.728287, 9.36434, 14.6009, 3.267204, 4.962337, 
    3.078237, 3.189939, 3.132822, 4.000747, 3.12495, 3.265537, 3.202188, 
    3.1882, 3.260356, 3.29556, 3.437104, 3.387794, 3.226074, 3.151515, 
    3.137635, 8.591904, 7.332052, 3.44105, 3.187157, 3.096544, 3.113197, 
    8.472248,
  17.83367, 20.17626, 21.8405, 3.385727, 22.44984, 3.130757, 10.18964, 
    3.093315, 8.628801, 3.357168, 3.321045, 3.28263, 3.385703, 3.486458, 
    3.463739, 3.683282, 3.624532, 3.724292, 3.4833, 3.447575, 3.190724, 
    6.067308, 3.413317, 4.006247, 3.41606, 3.268721, 3.151448, 3.152757, 
    22.91566,
  23.02053, 19.35734, 20.09576, 18.86843, 12.61588, 14.50615, 11.85608, 
    9.933898, 7.166511, 9.940439, 3.492388, 3.567873, 3.723592, 3.67032, 
    3.713316, 3.739949, 3.678763, 3.854204, 3.528728, 3.762489, 11.9292, 
    11.91544, 8.771135, 3.527946, 3.579979, 3.555734, 3.688622, 3.621299, 
    10.57927,
  6.188347, 3.862209, 6.195559, 9.967353, 1.976844, 14.72065, 8.719292, 
    14.62524, 12.64574, 10.90428, 7.285124, 3.795602, 3.614068, 3.563422, 
    3.606153, 3.49991, 3.585889, 3.625772, 3.588534, 11.79068, 10.68945, 
    12.86331, 12.10933, 4.350485, 3.749884, 3.693425, 3.74259, 3.756849, 
    5.166119,
  5.84121, 11.06509, 12.22004, 12.81276, 12.31121, 11.25619, 7.534362, 11.58, 
    8.168203, 6.882803, 6.816991, 6.200529, 3.828244, 3.858465, 3.944414, 
    3.956304, 3.752263, 3.916388, 3.910429, 8.463642, 9.951468, 9.316036, 
    6.373158, 6.19451, 5.002342, 3.825631, 3.726788, 3.921892, 4.083949,
  4.397814, 6.446847, 7.501013, 6.190328, 6.828495, 6.785339, 6.719504, 
    6.742296, 6.769308, 7.307252, 6.732722, 10.84201, 10.56142, 6.234003, 
    4.327715, 4.277146, 9.019155, 12.71124, 10.06658, 6.999386, 6.013795, 
    10.58687, 3.787417, 9.969274, 3.85788, 7.626759, 4.252257, 4.232515, 
    4.361547,
  4.105151, 4.61524, 6.938627, 4.119861, 4.101231, 4.920473, 11.18737, 
    11.72035, 12.52407, 12.09229, 10.7132, 9.338655, 11.93761, 4.911802, 
    17.50594, 4.236989, 9.246899, 12.01605, 7.611715, 6.906734, 17.70159, 
    11.29195, 15.12267, 27.89269, 4.47335, 42.39854, 43.15886, 8.870539, 
    4.261112,
  24.1229, 5.420525, 11.20607, 12.05765, 15.08401, 26.26855, 39.43262, 
    33.89502, 33.60452, 44.37672, 44.32983, 45.43599, 45.86336, 45.93732, 
    46.56146, 46.49811, 45.70898, 44.7709, 44.80893, 45.70079, 46.80277, 
    43.02631, 39.87453, 44.5517, 45.94991, 47.21799, 47.65586, 43.87235, 
    31.49117 ;

 average_DT = 730 ;

 average_T1 = 259 ;

 average_T2 = 989 ;

 climatology_bounds =
  259, 989 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
