netcdf atmos.1980-1981.alb_sfc.07 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float alb_sfc(time, lat, lon) ;
		alb_sfc:long_name = "Surface Albedo for  Flux" ;
		alb_sfc:units = "percent" ;
		alb_sfc:_FillValue = 1.e+20f ;
		alb_sfc:missing_value = 1.e+20f ;
		alb_sfc:cell_measures = "area: area" ;
		alb_sfc:interp_method = "conserve_order1" ;
		alb_sfc:cell_methods = "time: mean within months time: mean over years" ;
		alb_sfc:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:19 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.alb_sfc.07.nc reduced/atmos.1980-1981.alb_sfc.07.nc\n",
			"Mon Aug 25 14:40:06 2025: cdo -O -s -select,month=7 merged_output.nc monthly_nc_files/all_years.7.nc\n",
			"Mon Aug 25 14:40:01 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.alb_sfc.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.alb_sfc.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 alb_sfc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  3.893769, 3.957814, 3.984975, 3.75982, 3.360525, 3.367844, 3.736684, 
    3.297889, 3.443738, 3.492855, 3.329947, 3.218516, 3.29508, 4.035928, 
    4.120365, 4.198918, 4.370879, 4.013604, 2.189337, 3.905518, 4.230511, 
    4.157845, 4.062459, 3.720376, 4.363034, 4.448526, 4.215519, 4.233375, 
    4.171025,
  24.64448, 22.11505, 2.51651, 2.951343, 3.030559, 2.898912, 20.71697, 
    5.303041, 3.136072, 3.257371, 3.138627, 2.844691, 2.779058, 2.813788, 
    2.812222, 2.758431, 2.618274, 2.668301, 2.966527, 3.180755, 3.1746, 
    3.102262, 3.143943, 2.846476, 8.250247, 18.641, 24.69358, 24.64685, 
    25.08932,
  3.268646, 2.981042, 3.065086, 3.028602, 3.125591, 3.443169, 3.532747, 
    3.919787, 3.737343, 3.653876, 3.659802, 3.674549, 3.512769, 3.715965, 
    3.473058, 3.661293, 3.808983, 3.550088, 3.699895, 3.526358, 3.728127, 
    3.6411, 3.661794, 8.168527, 3.782351, 3.668315, 3.236194, 3.464187, 
    3.285471,
  3.55271, 3.888999, 3.984056, 3.939133, 3.819123, 3.836473, 4.023032, 
    3.836723, 3.995898, 3.917907, 4.141827, 4.046985, 4.351769, 4.122092, 
    11.4769, 4.095002, 3.914773, 3.926031, 3.737213, 3.699249, 3.557942, 
    3.506707, 3.626276, 9.389973, 4.265119, 3.791682, 3.961382, 3.592037, 
    3.760844,
  3.959295, 4.213758, 11.47938, 4.210011, 4.002475, 3.981825, 3.941133, 
    3.739111, 4.02416, 4.331559, 8.734747, 12.73454, 10.68067, 4.278761, 
    3.978963, 3.989288, 3.855234, 3.847867, 3.771066, 3.74169, 3.884342, 
    4.131775, 3.661839, 4.346064, 8.539532, 3.901964, 3.965643, 4.070668, 
    3.964937,
  3.388689, 9.420258, 9.72988, 3.827368, 4.084201, 4.100616, 3.720517, 
    3.919013, 3.55412, 4.232073, 11.52419, 11.77317, 3.942879, 3.730154, 
    3.665559, 3.610971, 3.920919, 3.740543, 4.034106, 3.817398, 3.923012, 
    3.404066, 3.238661, 3.849156, 8.793956, 8.850889, 3.829705, 3.669417, 
    3.426335,
  3.305635, 6.248497, 9.306512, 9.117855, 3.70272, 3.668977, 3.440277, 
    3.461504, 3.443296, 3.784505, 4.709443, 3.667914, 4.126745, 3.30078, 
    3.450619, 3.548276, 3.922378, 3.766535, 4.031528, 3.77492, 3.833939, 
    3.464999, 3.38008, 8.891066, 8.849451, 9.147311, 3.8194, 4.0281, 3.538044,
  3.191148, 8.637932, 8.512736, 10.1732, 3.523946, 3.251534, 3.168823, 
    3.19142, 8.69614, 8.449436, 3.318681, 3.301401, 3.535558, 3.42249, 
    3.432887, 3.579743, 3.675519, 3.806186, 3.6483, 3.719849, 3.653842, 
    3.515404, 3.409293, 8.467526, 8.642493, 3.565739, 3.553222, 3.453924, 
    3.407778,
  9.730167, 10.20761, 9.975561, 9.387707, 15.01674, 3.196598, 5.018166, 
    3.02397, 3.528544, 3.170757, 4.24186, 3.248659, 3.294413, 3.367255, 
    3.358724, 3.442703, 3.419716, 3.574326, 3.308482, 3.405231, 3.24552, 
    3.228845, 8.924456, 7.61975, 3.333212, 3.17745, 3.197472, 3.131694, 
    8.701424,
  19.19147, 21.59842, 23.48695, 3.345978, 23.91034, 3.093387, 10.24592, 
    3.263543, 8.846461, 3.334408, 3.416669, 3.341785, 3.470773, 3.539012, 
    3.550277, 3.815123, 3.75862, 3.819625, 3.503144, 3.437288, 3.352797, 
    6.697916, 3.430224, 4.072087, 3.491013, 3.404324, 3.418198, 3.204288, 
    24.67139,
  25.35246, 21.54479, 22.6327, 20.61969, 13.57708, 15.85847, 12.56262, 
    10.13175, 7.459718, 10.74393, 3.628049, 3.820002, 3.511331, 3.692544, 
    4.053599, 3.853418, 4.006166, 3.86092, 3.735098, 3.926968, 11.83777, 
    12.11118, 9.513004, 3.643644, 3.668504, 4.00719, 3.983634, 3.701885, 
    11.6777,
  8.25515, 4.137305, 6.753142, 11.156, 2.289236, 16.81276, 9.487543, 
    16.89839, 14.45383, 11.5083, 7.843853, 3.918589, 3.720922, 3.728784, 
    3.666089, 3.656257, 3.793622, 3.83622, 3.968376, 13.4553, 12.53626, 
    14.69349, 13.74583, 4.671746, 3.860129, 3.937924, 3.959774, 3.993908, 
    5.541318,
  6.644896, 13.56631, 15.12451, 15.84409, 14.99307, 13.53935, 9.132669, 
    11.84106, 8.346721, 7.887961, 7.744296, 7.315935, 4.119781, 4.168202, 
    4.007197, 4.035099, 4.001596, 4.05704, 4.163233, 10.35844, 11.73738, 
    10.88496, 7.751626, 7.443059, 5.695897, 4.219515, 4.335897, 4.17465, 
    4.544651,
  5.131839, 8.645904, 10.08397, 8.46305, 8.950133, 8.822401, 8.814001, 
    8.79633, 9.012403, 8.947889, 8.740297, 13.21627, 13.25886, 8.051533, 
    5.020106, 4.985484, 11.46976, 16.4708, 12.78504, 8.829653, 7.975107, 
    13.85026, 5.802172, 13.22037, 5.470679, 10.218, 5.02393, 5.002809, 
    4.825701,
  6.135005, 6.560645, 11.448, 7.154935, 6.887377, 48.50443, 19.64494, 
    17.77319, 18.71438, 18.31274, 13.54437, 12.59713, 18.28409, 34.90093, 
    54.33942, 14.93266, 26.75996, 24.5584, 19.83979, 25.44018, 28.28759, 
    45.12157, 33.73246, 41.93322, 9.736616, 66.60789, 71.50674, 15.79074, 
    6.44587,
  60.07027, 46.72136, 48.63533, 52.91319, 32.72775, 52.54621, 59.66739, 
    36.3352, 59.72209, 60.16356, 60.22125, 60.18361, 60.19011, 60.20282, 
    60.20239, 60.22253, 60.26421, 60.3139, 60.42854, 60.50266, 60.30748, 
    51.33521, 52.29346, 60.01953, 70.46642, 65.95874, 72.70717, 60.40523, 
    52.16167 ;

 average_DT = 730 ;

 average_T1 = 197.5 ;

 average_T2 = 927.5 ;

 climatology_bounds =
  197.5, 927.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 time = 0 ;
}
