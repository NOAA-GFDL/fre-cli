netcdf atmos.1980-1981.aliq.08 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:21 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.08.nc reduced/atmos.1980-1981.aliq.08.nc\n",
			"Mon Aug 25 14:40:48 2025: cdo -O -s -select,month=8 merged_output.nc monthly_nc_files/all_years.8.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.652274e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 3.698578e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.888449e-05, 0.0001594647, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0006555094, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -6.381267e-05, 0, 0, 0, 0.0001368089, 0.001304981, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -9.947018e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.001862315, 0, 0, 0, 1.371525e-05, 0, 0, 0.0001185111, 
    2.628516e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.071078e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -7.065535e-05, 0.0002230425, 0, 
    0.0007496308, 8.359431e-05, 0.0001433148, -7.280933e-06, -1.713477e-06, 
    0, 0, -1.727013e-05, 0.0021883, 0, 0, 0, 0, -1.581091e-06, -1.109009e-05,
  0, 0, 0, 0, 0, 0, -0.0001160855, 0, 0, -1.111657e-05, 0.0004641321, 
    0.002217565, -4.180533e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001427431, -2.149742e-05, 0, 0.0001580095, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.882883e-06, -5.00201e-05, 0, 0, 0, 0, 0, 0, 
    0.0002438873, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.002763859, 0, 0, -1.826303e-05, 0.001748657, 0, 
    1.143265e-05, 0.00266966, 0.0002294348, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.421495e-05, 0, 0, 0, 0, 0,
  0, 0, 9.090858e-05, 0, 0, 0, 0, 0, 0, 0, 0, 8.51205e-05, 0.001399778, 
    -5.589213e-05, 0.001066934, 0.00105064, 0.00037559, 0.0005513346, 
    -3.302932e-05, 0.0003754325, 0.0001677334, -3.775347e-05, 0.003831376, 
    3.149447e-05, -1.589167e-07, -1.095613e-05, 0.0002218378, 0.001635568, 
    0.002286826,
  0, 0, 0, 0, 0, -6.830212e-06, 0.0008857743, -1.890416e-07, 0.0004508504, 
    -8.542529e-05, 0.0007656344, 0.006052435, 4.194541e-05, -6.373176e-06, 0, 
    0, 0, 0, 0, 0, 0, 0.000117662, 0, -6.440996e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.0001988255, -0.0001168095, 0.0005414542, 0.0005260508, 
    0.0003642856, -3.656668e-06, 0.0002443249, 0.00129681, -2.190415e-06, 0, 
    0, 0, 0, 0, 0, 0, 9.645633e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.691587e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -8.009506e-05, 0.001028444, -6.734044e-06, 0, 0, 
    -9.900752e-08, 0, -1.157864e-05, 0.0002160664, -2.767234e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.003784267, 0, -2.788607e-06, -2.78047e-05, 0.005014447, 0, 
    2.248378e-05, 0.01282601, 0.0008931575, -1.229324e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.478048e-05, 0, 0, 0, 0, 0,
  -3.958909e-06, -6.136224e-06, 0.001903058, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004368455, 0.003366099, 0.001408234, 0.002003203, 0.002425299, 
    0.001585906, 0.002789217, 0.002582291, 0.001212471, 0.001148689, 
    0.001868543, 0.006151642, 5.018943e-05, -2.890508e-05, -0.0001095118, 
    0.001403147, 0.003716098, 0.00490715,
  0, 0, 0, -7.306974e-07, 0.0001196093, -3.812737e-05, 0.005016319, 
    -9.979087e-06, 0.00135808, 0.000158372, 0.0019754, 0.01164891, 
    0.0002815752, 0.0005721791, 0, 0, 0, 0, 0, 0, 7.01372e-05, 0.0002035778, 
    -1.167734e-05, -3.972592e-05, -9.263425e-08, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.00114281, 0.0002064498, 0.001837465, 0.001837983, 
    0.006199575, -3.249494e-05, 0.0008497524, 0.002315718, 0.0003426731, 0, 
    0, 0, 0, 0, 0, 0, 0.0007839616, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -3.536437e-06, 0, 3.231224e-05, -1.692309e-05, 
    -2.262667e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001566377, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.655974e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -7.608459e-08, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001047727, 0.002648997, 0.0002588793, 0, 0, 
    -9.900752e-08, -1.546134e-05, -4.682324e-05, 0.0003076358, -6.718512e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.006708466, 0, 3.106242e-05, 5.711806e-05, 0.009787591, 
    -2.141242e-05, 0.0007285324, 0.02567421, 0.00271529, -1.651118e-05, 
    -6.72263e-07, 0, 0, 0, 0, 0, 0, 0, 8.402942e-05, 0, 0, 0, 0, 0,
  0.0006684466, 0.001192118, 0.002371184, -1.866009e-06, 0, 0, 0, 
    5.859594e-05, 0, 0, -1.219612e-05, 0.001355455, 0.01191959, 0.004600439, 
    0.003666542, 0.005678718, 0.00391179, 0.007596191, 0.00646003, 
    0.005285614, 0.003609085, 0.003459329, 0.009093767, 0.001732937, 
    -4.523187e-05, -0.0001208922, 0.003059768, 0.006117956, 0.009857683,
  0, 0, 0, 0.0001152542, 0.0001724668, -5.145518e-05, 0.009775581, 
    -8.947824e-05, 0.002806188, 0.001351488, 0.006295675, 0.02046358, 
    0.001313394, 0.003424622, 0, 0, 0, 0, 0, 0, 0.0001703547, 0.001346229, 
    -1.766079e-05, 8.664321e-05, -6.625921e-06, 0, 0, 0, 0,
  0, 0, 0, 0, -7.046049e-09, -4.408154e-06, 0.001911226, 0.002720857, 
    0.003754077, 0.006296472, 0.01764978, 0.0008837918, 0.003074033, 
    0.005840648, 0.0005625472, 0, 0, 0, 0, 0, 0, -2.09257e-05, 0.001294535, 
    -3.086862e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 8.058516e-05, 0.001425135, 0.001265546, 
    1.321747e-05, -8.498667e-06, 0.0006503032, -1.597088e-05, 0, 0, 0, 0, 0, 
    -1.771611e-05, 0.0002599237, -1.486839e-05, 0.002366461, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.902531e-05, -1.19945e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -8.464258e-07, 0.0001090241, 0.0002514766, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.496168e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.071441e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.073639e-05, 0, 0, 0, 
    0, 0, 0, 0, -3.335398e-07, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.399504e-05, 
    -8.270905e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007389698, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -2.088978e-07, 3.832809e-05, 0.004735212, 0.008479377, 
    0.003399666, 0, 0, -6.481371e-05, -3.775122e-05, 0.0008025585, 
    0.0005057703, -1.881835e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -3.131014e-06, -1.054526e-06, 0, 0, 0.01142298, -2.285931e-05, 
    5.382284e-06, 6.738835e-05, 0.01707942, 7.854251e-06, 0.003767076, 
    0.03843018, 0.004770827, 0.0006018092, -5.779141e-06, 0, 0, 0, 0, 0, 0, 
    0, 0.0001135397, 0, 0, 0, 0, 0,
  0.002762041, 0.004124341, 0.005536465, 0.0002618307, 0, -6.750832e-06, 0, 
    0.0005169587, 4.491413e-06, -2.039735e-05, 6.041489e-06, 0.004753659, 
    0.02738479, 0.009953546, 0.005975806, 0.01240098, 0.0105553, 0.01458251, 
    0.01137685, 0.0130945, 0.006938923, 0.008747404, 0.01352682, 0.003919263, 
    -0.0001077136, -6.941861e-05, 0.0052484, 0.009191696, 0.02019214,
  0, 0, 0, 0.001135092, 0.002279564, 0.0006129806, 0.03179893, 0.0006195262, 
    0.005057697, 0.003208674, 0.02002673, 0.02851292, 0.006711654, 
    0.009147577, 4.673247e-05, 0, 0, 0, -7.343365e-09, 0, 0.0002209925, 
    0.007072779, -2.199997e-05, 0.0003941419, -2.14223e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 1.31418e-06, -1.560566e-05, 0.005563319, 0.004427244, 
    0.008517604, 0.01061075, 0.03676164, 0.002325779, 0.006509417, 
    0.008518226, 0.002990078, 0, 0, 0, 0, 0, 0, 0.0008382808, 0.002567373, 
    0.0001226171, -2.286075e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.001088121, 0.001891633, 0.007431107, 0.009892809, 
    0.002411412, 0.0007348278, 0.002399178, 0.000580915, 8.533599e-05, 0, 0, 
    0, 0, 4.648743e-05, 0.002612285, -2.613276e-05, 0.00431772, 0, 
    4.246275e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.369888e-05, 9.366283e-05, -0.0002366067, 
    0.0005163724, 0, -6.37436e-05, -4.667415e-05, 0, 0, 0, 0, 0, 
    -2.200469e-06, 0.001504201, 0.003049321, 0.003054612, -5.669046e-05, 
    0.0008787694, -4.362439e-06, -2.272088e-05, 0.0006228622,
  0, -3.322391e-05, -2.178938e-06, 0, 0, -1.030849e-05, 0, 0, 0, 
    -9.392525e-06, -2.456041e-06, -2.624874e-05, 0, 0, 0, 0.0001008359, 0, 0, 
    0, 0, 0, 0, 4.363852e-06, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -1.23238e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6.235456e-05, 0, 0, 0, 0, 0.0005731456, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.470881e-05, 
    0.0002858571, -3.571398e-06, 8.261855e-06, 2.286437e-05, 0, 0, 0, 
    -1.111716e-05, -3.39816e-05, -2.797232e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.626424e-05, 0.004425106, 
    0.0001638143, -3.265628e-05, 0.0005103695, 0, 0, 0, 0, 0.0005539014, 
    0.003002672, -5.469334e-09, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.70365e-07, 2.233482e-06, 
    0.005169475, 4.872838e-06, 0, 0, 0, 0, -2.348807e-07, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -4.123702e-06, 2.925888e-05, 0.01015358, 0.01688106, 
    0.004624524, 0, -1.303517e-08, 0.002231017, -5.54587e-05, 0.002809848, 
    0.002199383, -5.25028e-05, 0, 0, 0, 0, 0, 0, 0, 0, -6.845168e-09, 0, 0, 
    0, 0,
  0, 3.090392e-06, 7.613453e-06, 0, 0, 0.01817716, -0.0001954051, 
    0.0003447773, 0.00117044, 0.02688071, 0.0003311815, 0.007994307, 
    0.05626146, 0.01112283, 0.001448184, 5.112011e-06, 0, 0, 0, 0, 0, 
    -1.398686e-05, -3.045147e-08, 0.0002696418, -1.129939e-05, 0, 0, 0, 
    -4.57721e-06,
  0.005316976, 0.006558179, 0.009243253, 0.001564346, 0, 2.993204e-05, 
    0.0002056806, 0.001592153, 0.0001097654, 5.802079e-05, 0.0005886358, 
    0.009020722, 0.04907306, 0.01819211, 0.007787392, 0.02389486, 0.0241975, 
    0.02728859, 0.01761148, 0.02263271, 0.0177323, 0.02285476, 0.0261957, 
    0.006150529, 3.345702e-05, 0.001084166, 0.009224971, 0.02054889, 
    0.02990026,
  0, -1.05201e-09, -3.237701e-11, 0.006498009, 0.005357284, 0.008577231, 
    0.07459214, 0.003724085, 0.008712511, 0.01240261, 0.04405206, 0.04545785, 
    0.01642704, 0.02378056, 0.0004343051, 0, 0, 0, -2.386482e-05, 
    0.001817647, 0.004079864, 0.01576178, 0.000388629, 0.0006961696, 
    4.099405e-05, 0, 0, 0, 0,
  0, 0, 0, -3.195532e-11, 0.0004527931, 0.0006886117, 0.0166792, 0.006873737, 
    0.01447955, 0.02139492, 0.04734825, 0.006675069, 0.01884214, 0.01515663, 
    0.0149416, 7.317549e-05, 0, 0, 0, -2.936954e-05, -1.742067e-05, 
    0.001245233, 0.008145795, 0.003476419, 4.159046e-05, 0, 0, 0, 0,
  0, 0, 0, -6.716633e-11, 0, 0, -8.391756e-11, -1.233796e-07, 0.001766689, 
    0.003681768, 0.01374557, 0.01843089, 0.009815693, 0.007159052, 
    0.01039547, 0.002192586, 5.171548e-05, -3.044061e-06, -1.064797e-08, 0, 
    -5.160754e-06, 0.002100657, 0.005786197, -2.342719e-05, 0.007949532, 
    -1.818906e-05, 0.001957511, 0.0008040982, 0,
  0.0003490846, -9.333189e-06, 4.090191e-05, 0.0002033341, 0.000587024, 
    -1.630881e-05, 0, 0, 0.0001419959, 0.006052287, 0.006878374, 0.005411881, 
    0.0002848773, 0.00701471, 0.001565491, -5.730688e-06, 0.0001823577, 0, 0, 
    0, 0.0002630574, 0.003335344, 0.01201767, 0.007720803, 0.003579561, 
    0.001441541, 0.0002949419, -7.223551e-05, 0.00213902,
  2.770971e-05, -6.315604e-05, 0.001507682, 0, -1.159903e-06, -8.415601e-05, 
    -2.774331e-05, 0, -2.376825e-06, 0.0007409721, -0.0001138236, 
    0.005404236, -2.575551e-05, 0.0001702073, -2.2592e-05, 0.001504658, 
    -7.879928e-05, 0, 0, 0, 3.611562e-05, 2.247022e-05, 9.101594e-05, 
    -2.926281e-06, -1.051976e-05, -6.323211e-06, 2.320957e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.482301e-05, 1.465882e-08, 0, 2.953862e-10, 
    0, 0, 0, 0, 0, 0, -1.795511e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.492364e-10, 6.185945e-08, 
    2.07216e-07, -2.082601e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.002202114, 7.8426e-05, -1.51862e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0001493546, 0, 0, 0, -1.594291e-05, 0, 0.0001332498, 0, 0, 0, 
    0.0001299666, 0.00130506, 0,
  -3.10651e-05, 0, -2.786025e-06, 0.0002764458, 3.542402e-06, -9.17352e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, -1.884289e-05, 0.0003110505, -2.455704e-05, 
    0.0009661144, 0.002370244, 6.493995e-05, 0.0004945006, 0.003810009, 
    -1.470632e-07, 0, 0.0006874473, 0.003703195, 0.001131029, 0.0006008146, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -1.181826e-10, 0, 0, 0, 0, 0, 1.822753e-07, 
    0.003991412, 0.0155568, 0.008769193, 0.00275519, 0.003727196, 0, 0, 0, 0, 
    0.002466679, 0.01277015, -5.19435e-06, 0, 0,
  0, 0, 0, 0, 0, 0, -1.680057e-06, 0, 0, 0, 0, 0, 0, -3.202214e-06, 
    0.0001667409, 0.006160459, 0.01041931, 0.001645401, -8.836311e-09, 0, 0, 
    -3.874255e-06, -4.366079e-08, -9.066865e-10, 0, -5.170263e-06, 0, 0, 0,
  1.340317e-07, -1.140284e-09, 0, 0, -6.546262e-06, 1.842047e-05, 0.02322339, 
    0.03685343, 0.006638482, 3.640238e-05, 2.006838e-05, 0.008701769, 
    0.0006249663, 0.007592229, 0.004799304, 4.203234e-05, 3.054033e-09, 0, 0, 
    6.531881e-08, -3.512598e-10, -1.105024e-09, 1.039461e-08, -1.958375e-06, 
    -1.3429e-05, 2.868846e-07, 0, -6.778028e-10, 0,
  -1.865688e-08, 0.0008765397, 0.0002534478, 0, -3.268145e-10, 0.03307074, 
    0.002557522, 0.005939513, 0.008698484, 0.04451287, 0.005346856, 
    0.01975377, 0.0856054, 0.02715562, 0.002880072, 0.0002107636, 0, 
    -6.504555e-08, -5.071641e-08, -1.228198e-07, 0.0001754882, 0.0002083672, 
    -1.069797e-05, 0.006134507, 2.748059e-05, -1.497158e-05, -4.550253e-06, 
    0, 4.248029e-06,
  0.01277557, 0.0122525, 0.01445961, 0.007042388, 2.694049e-05, 
    -4.402898e-05, 0.001476819, 0.01547335, 0.002802554, 0.003031387, 
    0.001818358, 0.02099684, 0.09414043, 0.03306141, 0.02279331, 0.04647544, 
    0.04984127, 0.04256277, 0.03095949, 0.03765305, 0.04350568, 0.05390585, 
    0.06083368, 0.01446653, 0.00134447, 0.005930008, 0.01539984, 0.04152716, 
    0.04576828,
  -4.208983e-08, -9.124881e-07, -1.914603e-05, 0.01733253, 0.0217604, 
    0.05097523, 0.1220534, 0.05602919, 0.03902819, 0.07471213, 0.08012308, 
    0.07729402, 0.05064628, 0.05580765, 0.00479422, 6.369738e-05, 
    -1.69049e-09, 0, 0.0009199069, 0.003542409, 0.008567515, 0.03971674, 
    0.002339451, 0.002138612, 0.002126416, -5.828964e-10, 0, 5.767264e-07, 0,
  0, 0, 0, -1.116934e-06, 0.001302398, 0.002297872, 0.1007302, 0.01132421, 
    0.02522387, 0.05868024, 0.08608991, 0.02072765, 0.0534368, 0.03137793, 
    0.03101185, 0.003236482, -2.261718e-05, 0, 0, -4.839166e-05, 
    8.089066e-05, 0.005679377, 0.02430134, 0.008483564, 0.0002206952, 
    0.0007234249, 0, 0, 0,
  0, -3.543101e-06, 0.0005040363, 1.577367e-07, 5.598963e-06, 4.863743e-05, 
    -1.1201e-07, -2.534519e-05, 0.005362091, 0.007845447, 0.03273614, 
    0.03503481, 0.01817677, 0.01853233, 0.02700548, 0.005413725, 0.00311692, 
    0.0005267612, -2.632943e-05, 0, -4.325579e-05, 0.006139485, 0.008809648, 
    0.003661814, 0.01358603, 0.001843586, 0.006492358, 0.004733223, 0,
  0.002333681, -2.636293e-05, 0.002531859, 0.001207433, 0.002545994, 
    -2.365797e-05, 0, 0.0002079033, 0.007727662, 0.01661526, 0.01811774, 
    0.01673686, 0.007164346, 0.02902251, 0.005392442, 7.906639e-06, 
    0.004139422, 3.972252e-05, 0.001625706, -1.31472e-05, 0.001249713, 
    0.006790605, 0.02359813, 0.01473549, 0.01597552, 0.008682293, 
    0.005647712, 0.0005761366, 0.005407164,
  0.0004894946, 0.002503067, 0.004085143, -5.391599e-07, 0.0007259414, 
    0.0006274637, 9.742715e-06, 0.0002473875, 0.0003775614, 0.003136158, 
    0.0001863731, 0.02319202, 0.004897221, 0.002385754, 0.001875607, 
    0.004878907, 0.00357787, 0, 0, 0, 0.001100155, 0.0001981158, 0.002452759, 
    -1.646629e-05, 0.002854259, 0.001764519, 0.0007021066, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001077516, 0, 0, 0, -2.424341e-05, -4.318081e-05, 
    -5.832257e-05, -5.374396e-05, 0, 0, 0, 0, 0, -4.331338e-05, 0.0004408853, 
    -8.642678e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.918994e-11, -8.278917e-10, 
    1.189969e-07, 1.279739e-07, 0, 0, 1.226717e-09, -7.196587e-11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.0005656705, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0.0004555797, 0.0001877487, 0, -2.639765e-05, 0.004763741, 6.911719e-05, 
    1.584527e-05, -1.299354e-05, -5.677521e-07, 0, 0, 0, 0, 0, -4.640924e-06, 
    0, 0.001824928, 0, 0, 0, 0.001289187, -3.029093e-07, 0.0004703579, 
    -4.439526e-06, 0.0002792577, 0, 0.0002444582, 0.00198192, 0,
  0.0003768936, 0, -5.428823e-06, 0.006821977, 0.003336985, 0.005765096, 
    3.379334e-05, 0, 0, 1.69326e-10, 0, 0, 0, -3.449401e-06, -6.245911e-05, 
    0.003783349, 0.0001153133, 0.004972429, 0.006096335, 0.007984142, 
    0.005571235, 0.005652494, 0.00110588, 0, 0.00156864, 0.008485315, 
    0.005783051, 0.005664723, -4.362572e-05,
  0, 0.0003104046, 0, -1.139444e-10, 0.003547589, -1.134131e-05, 
    1.633021e-07, -8.534208e-10, -5.923754e-07, 1.596002e-07, -1.05825e-09, 
    0, -1.060051e-11, -7.29808e-09, 0.001379196, 0.01616247, 0.03336878, 
    0.02905606, 0.01460876, 0.006351864, 0.0004116173, 1.312052e-05, 0, 
    0.0002657648, 0.005563246, 0.02094823, 0.0001226805, 2.51297e-07, 
    -7.346669e-06,
  1.74581e-07, -1.685414e-08, 0, 2.535165e-09, 5.434324e-08, 3.22945e-07, 
    1.283075e-05, 3.993889e-07, -1.198076e-06, 3.962987e-07, 1.809811e-05, 
    1.368827e-07, -2.630312e-05, 0.0009441528, 0.001713102, 0.02053577, 
    0.01905261, 0.006937662, 2.041673e-05, 4.180219e-05, 0, -3.573865e-07, 
    2.340094e-05, 7.038201e-06, 6.855096e-05, 5.962599e-05, 1.262698e-07, 
    -1.588097e-08, 0,
  2.098014e-05, 0.0003854625, -4.591507e-06, -5.093695e-09, -8.236768e-06, 
    0.00244367, 0.04128925, 0.05928023, 0.01834019, 0.005823236, 0.005033182, 
    0.05732573, 0.01105254, 0.02905831, 0.02488582, 0.001916725, 
    1.226833e-06, -8.195827e-09, 2.69764e-08, 0.0002609071, 0.0002768322, 
    -6.831045e-07, -5.476414e-06, 6.208775e-05, 0.0006169862, -2.682262e-05, 
    5.481169e-06, 2.078972e-05, 4.766888e-06,
  9.518231e-05, 0.008159673, 0.004565825, -1.984837e-06, 2.317528e-07, 
    0.05302193, 0.01058816, 0.03234924, 0.05871098, 0.08808316, 0.1150698, 
    0.1502549, 0.1991307, 0.08514975, 0.049671, 0.004589343, 0.0003699562, 
    -3.808604e-06, 4.325615e-05, 0.00043171, 0.0004550161, 0.002503481, 
    0.003072579, 0.0249102, 0.0009828383, -6.065518e-06, 0.0002352304, 
    0.006893455, 0.002258027,
  0.06598078, 0.03694388, 0.04396147, 0.01946142, 0.0004590529, 0.0106791, 
    0.1454325, 0.4618304, 0.3426508, 0.1950972, 0.2592062, 0.2313686, 
    0.3006229, 0.1511305, 0.1604839, 0.1589874, 0.1036902, 0.08231296, 
    0.0752764, 0.08555038, 0.1245874, 0.1917668, 0.1361217, 0.05184621, 
    0.01543313, 0.01389976, 0.02613293, 0.08271962, 0.07631144,
  4.846373e-07, 0.0001277046, 0.01010928, 0.07560734, 0.1124781, 0.1724168, 
    0.320585, 0.2110961, 0.3313785, 0.2507125, 0.2916431, 0.2404893, 
    0.2989798, 0.216263, 0.05000447, 0.0005848515, -3.274516e-05, 
    -8.418855e-08, 0.006768824, 0.008440555, 0.07762978, 0.1478839, 
    0.05980444, 0.01798822, 0.009789786, -1.271153e-06, 3.592071e-05, 
    0.0004068327, -1.510706e-07,
  2.773436e-06, 0, -5.146841e-08, 0.0006791416, 0.009483863, 0.01396749, 
    0.1100026, 0.0257672, 0.04294714, 0.1777575, 0.1683473, 0.1386429, 
    0.1660375, 0.0915371, 0.08941906, 0.006809768, 0.0001578665, 
    0.0002720541, 0.0001276835, 0.0001139737, 0.001870238, 0.03851826, 
    0.09350432, 0.02373222, 0.002659808, 0.001183441, -6.122121e-08, 
    -3.558845e-08, -7.71339e-09,
  1.093763e-05, -1.896166e-05, 0.00199194, 2.774903e-06, 0.0005214174, 
    0.001422112, 5.841794e-07, 0.001479976, 0.03004301, 0.03081188, 
    0.1130766, 0.1474964, 0.07239791, 0.06685227, 0.08163976, 0.0201274, 
    0.01833012, 0.002224269, -3.206957e-05, -1.402981e-07, 0.0006994058, 
    0.0117981, 0.01752839, 0.01301281, 0.03421038, 0.002154568, 0.01156598, 
    0.008190843, 5.078454e-07,
  0.006211947, 0.0006841468, 0.01655798, 0.003746848, 0.004697828, 
    0.002201982, 0.000176012, 0.0007548335, 0.02212741, 0.03821238, 
    0.04708483, 0.04134085, 0.03411504, 0.06373682, 0.03669009, 0.008841012, 
    0.01422039, 0.006547656, 0.004883289, 0.000127712, 0.002308398, 
    0.02013862, 0.0391358, 0.02925295, 0.02554647, 0.02497625, 0.01457969, 
    0.008460695, 0.01202771,
  0.006054656, 0.004702494, 0.009936098, 0.0009006578, 0.001722643, 
    0.002492123, 0.004320945, 0.0003160174, 0.00184827, 0.01182956, 
    0.008278655, 0.04015507, 0.009313982, 0.004708658, 0.007543526, 
    0.009520301, 0.007033297, 9.322585e-05, 0, -8.515458e-07, 0.003439033, 
    0.002229544, 0.0163239, 0.001302054, 0.01435731, 0.007402523, 
    0.006909199, 0.0007658936, 0.0001939165,
  0, 0, 0, 0, 0, -1.094601e-05, 0.004225889, 0.002841741, 0, 0.0009326469, 
    0.001950751, 0.0001159953, 0.0004141722, 0.0003907925, 0, -6.992776e-06, 
    -2.472969e-06, 0, -3.589849e-06, 4.620526e-05, 0.004236362, 
    -5.951908e-06, 0, 0, 0, 0, 0, 0, 0.0004162709,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.326676e-10, 2.226536e-08, 0.000181536, 
    -0.0001764729, -9.55098e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -8.420706e-06, 0, 0, 0.001693768, 0, 0, 0, 0, 0, 0, 2.789592e-05, 
    -3.165372e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.002712206, 0.001129945, -7.451581e-06, 0.0003893364, 0.01148579, 
    0.001431185, 0.001931534, -1.460029e-05, 0.0009913873, 2.414665e-06, 
    -2.707957e-06, 0.00077718, -3.200269e-05, -2.61329e-06, 0.001378254, 
    1.089259e-05, 0.00432927, 0.001006635, -8.566334e-06, -6.101843e-05, 
    0.004283405, 0.0003348638, 0.003182712, 0.0002177054, 0.001255461, 
    -1.027765e-05, 0.001256113, 0.00351583, -8.164742e-06,
  0.0005630614, -2.764095e-08, -2.434606e-05, 0.01572609, 0.008443064, 
    0.01319254, 0.003282448, -2.830821e-06, 4.904968e-08, 2.252088e-08, 
    3.178329e-10, -5.509075e-06, 1.773563e-05, 0.001347907, 0.003189229, 
    0.00703638, 0.00293695, 0.01675795, 0.0207289, 0.03057392, 0.03909796, 
    0.01759838, 0.003291425, 0.002771625, 0.003042832, 0.0142772, 0.01646636, 
    0.01956756, 0.003958018,
  7.44692e-06, 0.0005218916, 0, -1.778398e-06, 0.007973797, 0.0006862427, 
    3.149367e-05, -1.670386e-06, -1.683502e-05, 6.316648e-05, 1.267282e-05, 
    -7.759111e-07, 2.505127e-07, 1.587272e-06, 0.004465358, 0.03217318, 
    0.06492706, 0.07374177, 0.04431751, 0.009379529, 0.002979277, 
    0.002322022, -6.01353e-06, 0.0007123533, 0.009948333, 0.02953854, 
    0.007268595, 0.0006278863, 1.573987e-05,
  1.661711e-05, 0.000212372, 1.978263e-07, -3.398883e-09, 7.886993e-07, 
    -1.416685e-08, -2.030164e-05, -1.400008e-05, 9.963701e-06, 3.916788e-07, 
    1.431997e-05, 2.546047e-07, -0.0001388141, 0.002239035, 0.006500952, 
    0.04365885, 0.05626742, 0.02651628, 0.0018339, 3.935676e-05, 
    3.444724e-05, 0.0001335448, -1.453463e-05, 0.009500069, 0.005637588, 
    -1.211261e-05, 0.003610167, 6.72395e-05, 5.067517e-05,
  0.00236097, 0.002275012, 8.393795e-06, -5.066837e-05, 0.005432102, 
    0.03026713, 0.0688182, 0.1178294, 0.04352283, 0.01472755, 0.009058164, 
    0.06228906, 0.01849445, 0.03990769, 0.02635373, 0.02080719, 0.0005359931, 
    0.0001959555, 8.442902e-07, 0.005596729, 0.0008627641, 0.0004906374, 
    0.008970116, 0.01829791, 0.0249613, 0.02158594, 0.01101055, 0.003196789, 
    3.72441e-05,
  0.0452944, 0.3164829, 0.2783229, 0.0001393469, 0.00272487, 0.1704731, 
    0.207268, 0.2670916, 0.3811911, 0.3135194, 0.2681372, 0.1908341, 
    0.2074602, 0.07590513, 0.04594443, 0.005009956, 0.0006988413, 
    7.382863e-05, 3.200745e-05, 0.02500135, 0.05077571, 0.02252074, 
    0.08651562, 0.1836336, 0.03473162, 0.008349389, 0.02967981, 0.07182424, 
    0.0277875,
  0.3221187, 0.3885759, 0.3561699, 0.03622339, 0.01253652, 0.04549533, 
    0.2053465, 0.3843206, 0.2273778, 0.115434, 0.1927173, 0.1764074, 
    0.2553051, 0.1286731, 0.1521401, 0.1668375, 0.1199418, 0.1383794, 
    0.1168609, 0.1485026, 0.1959517, 0.2471237, 0.3389073, 0.1463476, 
    0.08076721, 0.09981749, 0.1275427, 0.2174919, 0.3073595,
  1.1583e-05, 0.003329137, 0.0108685, 0.0700502, 0.125145, 0.1427362, 
    0.2892318, 0.1576418, 0.3072074, 0.1788841, 0.2233354, 0.2049548, 
    0.2596296, 0.2925079, 0.2238364, 0.08916185, 0.00655014, 9.954599e-06, 
    0.007216158, 0.009334078, 0.06100628, 0.1990014, 0.1135986, 0.07829981, 
    0.08096841, 0.02297807, 0.00412745, 0.002511142, 0.0001961537,
  2.615849e-06, 0, -4.531548e-08, 0.001099439, 0.007146536, 0.01155082, 
    0.08803722, 0.05452286, 0.07912733, 0.139117, 0.1460431, 0.1080638, 
    0.1580833, 0.1598466, 0.2077342, 0.03384293, 0.05854866, 0.01390014, 
    0.004657701, 0.01205184, 0.06072743, 0.1486767, 0.2823825, 0.166934, 
    0.08680016, 0.07666851, 0.01225434, -1.456493e-06, -6.214254e-05,
  0.008830891, 0.001691513, 0.003270466, 0.0001191317, 0.001243848, 
    0.00322327, 0.0001762415, 0.03503127, 0.08901387, 0.09114146, 0.1920254, 
    0.1937277, 0.1028744, 0.1773977, 0.2365913, 0.1523257, 0.1208158, 
    0.06567401, 0.02639172, 0.0004217575, 0.005128711, 0.05718173, 
    0.07466104, 0.1114476, 0.1953021, 0.05769841, 0.07025644, 0.03479917, 
    0.00657717,
  0.009390041, 0.009536467, 0.03569212, 0.005971317, 0.009664728, 0.01082414, 
    0.0004716778, 0.00146082, 0.03713211, 0.07475747, 0.1291916, 0.1665657, 
    0.143874, 0.1966877, 0.1217894, 0.1102406, 0.06401471, 0.04317709, 
    0.03061233, 0.00159922, 0.008848267, 0.03832221, 0.07117417, 0.0503284, 
    0.04594411, 0.06355673, 0.05185675, 0.03533827, 0.02506768,
  0.01457277, 0.007677603, 0.01504141, 0.005159033, 0.002384, 0.01226086, 
    0.01129371, 0.0003070573, 0.007168634, 0.03086893, 0.0411261, 0.06447995, 
    0.02187307, 0.02354042, 0.0311069, 0.02650683, 0.00974884, 0.005249634, 
    0.0002341661, 0.0001983382, 0.009384025, 0.01041172, 0.03175559, 
    0.004487108, 0.02670798, 0.01431426, 0.01821644, 0.005351439, 0.003699068,
  -2.687331e-05, -6.351037e-06, 0.0006898812, -0.000138528, 0.0004517646, 
    0.004462833, 0.007171158, 0.006622877, -3.816764e-05, 0.003091329, 
    0.004320919, 0.00120875, 0.0004641954, 0.001437472, -9.49263e-05, 
    -9.829282e-06, 6.468501e-05, -1.602355e-05, 6.569504e-05, 0.001121861, 
    0.009190267, 0.003853785, 0.0004704317, -3.755081e-05, 0, 0, 
    -1.433997e-06, -1.189336e-05, 0.002205608,
  0, 0, 0, 0, 0, 0, 0, -6.896069e-05, -2.082604e-05, -3.010855e-05, 
    6.188806e-10, 5.986385e-07, 4.240272e-07, 0.0006931183, 0.001922521, 
    -1.439707e-09, -2.286105e-07, -1.09286e-05, 2.488431e-06, -1.884308e-06, 
    0.002295281, -3.920203e-05, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, -3.230685e-05, -1.383309e-06, -5.213577e-06, 0.00280636, -8.563659e-06, 
    -6.751319e-06, 0, 0.000332462, 0.0003793885, -2.964663e-05, 0.0006109062, 
    0.0009812926, 3.086727e-05, -5.175315e-07, 0, -1.046639e-05, 
    0.0002709469, 0, 0, 0.0001447232, 0, -7.355875e-06, -9.601407e-06, 
    -1.871133e-06, 0, 0, 0, 0,
  0.006322276, 0.002580796, 0.002873675, 0.003097221, 0.02399402, 
    0.005168067, 0.008003555, 0.00315195, 0.002006737, 0.0005406251, 
    -3.256138e-05, 0.001896219, -1.269097e-05, 0.002090941, 0.007083653, 
    3.289618e-05, 0.005931011, 0.002123202, -4.414761e-05, -0.0002956858, 
    0.008660389, 0.003983012, 0.01376923, 0.004857301, 0.001786437, 
    0.0009809432, 0.007523373, 0.009212805, 0.0003016463,
  0.003869709, 4.259756e-05, 0.0002479689, 0.0328057, 0.01529577, 0.0197725, 
    0.01392584, -3.479305e-05, -1.430076e-05, 2.903941e-06, 2.508805e-05, 
    0.0007639765, 0.002368708, 0.002898096, 0.01291371, 0.0177924, 
    0.008317208, 0.04088214, 0.05403607, 0.05470736, 0.07912399, 0.04391599, 
    0.01660583, 0.01295648, 0.01127934, 0.03216702, 0.04830842, 0.03553817, 
    0.01417781,
  0.004710885, 0.009266108, 2.069765e-05, 0.000789058, 0.01041289, 
    0.007614116, 0.003445706, 0.0002528643, 2.455431e-07, 0.003354046, 
    0.003086531, -8.24497e-06, 0.0001940544, 0.001223404, 0.006209401, 
    0.0461714, 0.1124049, 0.1285862, 0.08775778, 0.04209484, 0.03774262, 
    0.02279662, 0.003100947, 0.003006484, 0.01773069, 0.06394287, 0.03457184, 
    0.01936495, 0.005517287,
  4.488651e-06, 2.345703e-05, 4.204554e-06, -1.964994e-09, 2.382838e-05, 
    -1.42895e-07, -5.050209e-07, 1.697912e-05, 2.600887e-06, 5.469087e-07, 
    1.382497e-06, 4.080913e-07, -2.831714e-05, 0.002307257, 0.01848835, 
    0.04653544, 0.04539193, 0.01828902, 0.008629918, 7.497591e-05, 
    8.400842e-06, 1.608425e-05, 3.737581e-06, 0.005223048, 0.009313015, 
    0.01100838, 0.000533175, 7.802336e-05, 3.25538e-06,
  2.799465e-05, 5.510981e-05, 2.915907e-05, -8.132278e-06, 0.0009399969, 
    0.01266184, 0.06263213, 0.09749921, 0.03066149, 0.00628097, 0.006723185, 
    0.04449525, 0.010404, 0.03397819, 0.01846985, 0.01512789, 0.000122433, 
    0.0002286764, 7.035338e-08, 9.253283e-05, 5.869499e-05, 4.003496e-05, 
    0.002839154, 0.002569166, 0.01913483, 0.01381496, 0.00362737, 
    0.0001405914, 1.191917e-06,
  0.035159, 0.230138, 0.1781139, 0.00068793, 0.000788091, 0.1158897, 
    0.1252041, 0.1983612, 0.3195668, 0.278708, 0.1747161, 0.1529769, 
    0.196378, 0.06668016, 0.02851142, 0.002776749, 2.759664e-05, 
    9.015785e-06, 8.582312e-06, 0.003397201, 0.007361929, 0.008349586, 
    0.05625449, 0.132427, 0.01761998, 0.003928115, 0.016472, 0.05172434, 
    0.009451735,
  0.2792962, 0.3423209, 0.287104, 0.1387457, 0.005508089, 0.02386414, 
    0.1061606, 0.2685746, 0.1466844, 0.05350457, 0.09902298, 0.1237507, 
    0.217887, 0.09946521, 0.1164654, 0.1200015, 0.08657797, 0.106542, 
    0.09092167, 0.11265, 0.1717732, 0.2118585, 0.2792098, 0.09932128, 
    0.04887329, 0.06396553, 0.08988178, 0.1814685, 0.2643825,
  2.462531e-05, 0.001319328, 0.006624364, 0.06842388, 0.136937, 0.1184931, 
    0.2519423, 0.1251337, 0.2896037, 0.1407357, 0.2081391, 0.1906319, 
    0.2166159, 0.2236515, 0.1804298, 0.06231515, 0.0003522068, 3.133932e-06, 
    0.005110295, 0.007056527, 0.05056387, 0.1493757, 0.07073043, 0.04817275, 
    0.04441967, 0.01371457, 0.005066233, 0.0004988679, 0.0005672821,
  -6.97673e-07, 0, -3.756452e-09, 0.001029293, 0.006108555, 0.008580186, 
    0.08013318, 0.1344844, 0.1405296, 0.1082559, 0.1347449, 0.07915264, 
    0.1393668, 0.13523, 0.2073886, 0.03912587, 0.1147837, 0.01638518, 
    0.00117263, 0.007353137, 0.09935943, 0.09402677, 0.2048795, 0.1267984, 
    0.06059685, 0.06616677, 0.01656548, 1.573009e-05, 0.0002508429,
  0.05178108, 0.01154552, 0.007144047, 0.001839666, 0.003439747, 0.01123352, 
    0.001370768, 0.06715987, 0.1433772, 0.1362136, 0.1931441, 0.1862669, 
    0.08925804, 0.16142, 0.2283756, 0.2243189, 0.1657127, 0.1325061, 
    0.03848755, 0.003138364, 0.07444727, 0.07952601, 0.1071802, 0.09084626, 
    0.1885842, 0.07806124, 0.1098563, 0.07040242, 0.03725098,
  0.101574, 0.05128865, 0.08048761, 0.02852373, 0.03974029, 0.06735196, 
    0.04591278, 0.002148806, 0.05873299, 0.1499436, 0.1947362, 0.2234562, 
    0.1841494, 0.2305043, 0.1892176, 0.1304612, 0.1052991, 0.1060847, 
    0.1076528, 0.003339, 0.0609658, 0.1198836, 0.1120425, 0.1181081, 
    0.1137447, 0.1466599, 0.1554154, 0.1432207, 0.1349097,
  0.06964059, 0.01478752, 0.02768141, 0.01330302, 0.007101772, 0.04801981, 
    0.05125879, 0.01718432, 0.02792574, 0.09604473, 0.1450396, 0.1327936, 
    0.03831466, 0.07319729, 0.1241182, 0.1133467, 0.05594474, 0.0406388, 
    0.002621555, 0.02437618, 0.02276101, 0.05527509, 0.08483236, 0.03986254, 
    0.06131712, 0.03776854, 0.04118401, 0.04265657, 0.02858161,
  -0.0001634556, 4.31047e-05, 0.0009130876, 0.003020674, 0.004687418, 
    0.007678588, 0.01671776, 0.01292518, 0.01197355, 0.02598942, 0.03890168, 
    0.02799665, 0.03753575, 0.03613788, 0.01608394, 0.01188474, 0.009522131, 
    0.01112043, 0.01632416, 0.01256894, 0.02646793, 0.01744252, 0.01096734, 
    0.002436377, -3.512061e-05, -1.168391e-05, -2.823416e-05, 0.006677787, 
    0.005592848,
  -1.959337e-08, 0, -2.900557e-07, 8.840285e-05, -2.885335e-05, 0, 0, 
    -0.0002370214, -1.364637e-05, -1.027766e-05, 1.068577e-06, -3.402474e-06, 
    -2.560736e-05, 0.001117005, 0.002497558, -4.013871e-05, 0.001174868, 
    0.0006346415, 0.001479977, -2.393295e-05, 0.003755467, 0.001558985, 
    1.276259e-05, -8.974877e-08, -1.008615e-05, -9.577627e-07, 0, 
    -2.095102e-07, 6.720733e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.418303e-07, -1.078852e-05, 
    9.02117e-05, -3.27673e-05, 0, -2.202278e-05, 0, -2.604834e-05, 0, 
    -7.028292e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0.001156266, -6.961943e-06, 0.000662536, 0.004169847, 0.002241714, 
    0.001156526, 3.529595e-05, 0.0008273991, 0.001841684, 0.0009520049, 
    0.001048582, 0.002235732, 0.004331763, 0.001037385, 0.0002729122, 
    -6.146642e-05, 0.001579301, -3.441007e-06, 0.001851998, 0.002412209, 
    2.943336e-05, -4.291614e-05, 0.0005503928, 0.000461732, 0.0002778833, 
    -1.234428e-05, -3.793192e-06, 0,
  0.0130715, 0.004434277, 0.01321332, 0.007203941, 0.0452522, 0.02089349, 
    0.01506826, 0.007343008, 0.00577862, 0.002890648, 0.003952476, 
    0.00598581, 0.002007527, 0.01254284, 0.02398045, 0.002456536, 0.01061285, 
    0.01391733, 0.003066401, 0.002839266, 0.01772504, 0.0148841, 0.03196844, 
    0.02061572, 0.008320872, 0.01740195, 0.02316232, 0.02803778, 0.006299078,
  0.04123166, 0.02333361, 0.02786135, 0.08190709, 0.03387602, 0.04087812, 
    0.04733483, 0.02245989, 0.01137606, 0.005621682, 0.00748426, 0.009540852, 
    0.01402137, 0.01021642, 0.03278091, 0.04815955, 0.03447497, 0.07775754, 
    0.0981722, 0.1105267, 0.1363364, 0.1118396, 0.08449072, 0.04014604, 
    0.06310029, 0.1232337, 0.1427727, 0.1149192, 0.08217497,
  0.003994868, 0.005281176, 0.003946054, 0.01033315, 0.02836339, 0.01408681, 
    0.007828907, 0.005382475, 0.003338203, 0.005684927, 0.004687242, 
    0.005313322, 0.005746773, 0.000934243, 0.01047796, 0.05717872, 0.1499194, 
    0.1773992, 0.1172583, 0.07176957, 0.04880901, 0.03205168, 0.01708764, 
    0.006685887, 0.0233367, 0.07014292, 0.04839526, 0.02485495, 0.01021948,
  1.271038e-06, 4.050452e-06, 1.387691e-06, -1.097574e-09, 0.0001462917, 
    8.796277e-08, 1.807177e-06, 0.0008981993, 0.0005506595, 1.238404e-06, 
    2.896278e-06, 2.867104e-07, 4.386971e-07, 0.002900621, 0.02972186, 
    0.04441554, 0.03491854, 0.01136549, 0.004572003, 9.541732e-06, 
    2.894596e-07, 3.028313e-06, 3.095399e-06, 2.82438e-05, 0.009346818, 
    0.02193682, 0.0002449796, 0.0001234818, -6.071978e-05,
  7.074743e-06, 1.300023e-05, 2.361551e-06, 5.518425e-06, 3.446726e-06, 
    0.005017398, 0.05481938, 0.09075947, 0.02952164, 0.005533168, 0.00450416, 
    0.04333169, 0.01166204, 0.03378916, 0.01935983, 0.01491252, 0.0005864305, 
    7.02456e-05, -2.127922e-09, 2.839192e-06, 1.196931e-05, 1.815334e-06, 
    0.0001715337, 0.0008260711, 0.01610083, 0.005073, 5.266569e-05, 
    2.907128e-06, 2.054612e-07,
  0.01226185, 0.1519312, 0.09863899, 0.00158203, 0.0002615104, 0.09186308, 
    0.0802534, 0.1467668, 0.2815251, 0.2449568, 0.1251622, 0.1437092, 
    0.202633, 0.06999275, 0.02913286, 0.002745885, 2.465879e-05, 
    5.560768e-06, 8.535509e-06, 5.504869e-05, 0.00108258, 0.00309824, 
    0.03882883, 0.09839867, 0.01491211, 0.002012888, 0.002554901, 0.03333763, 
    0.006899679,
  0.2640393, 0.3318661, 0.2500642, 0.1146201, 0.001118846, 0.009400243, 
    0.06766233, 0.1513292, 0.1110391, 0.0327752, 0.05647565, 0.1066988, 
    0.2033277, 0.09629364, 0.1061284, 0.1003727, 0.07890686, 0.09706409, 
    0.07801673, 0.1067566, 0.1606602, 0.1880076, 0.2552895, 0.08471385, 
    0.04844905, 0.05469438, 0.08176528, 0.1665078, 0.2611929,
  2.094012e-05, 0.00114483, 0.007536661, 0.06641623, 0.1233649, 0.1226132, 
    0.2279295, 0.091777, 0.2711612, 0.1042204, 0.1837283, 0.1765975, 
    0.1808342, 0.1832999, 0.1569229, 0.04976888, 0.000272047, 2.002456e-06, 
    0.005920666, 0.005651874, 0.04697603, 0.1227909, 0.0548703, 0.03552673, 
    0.03432402, 0.007630925, 0.004861695, 0.0003082642, 0.002051316,
  -1.659785e-08, 0, -2.162279e-08, 0.001041129, 0.005584022, 0.008710471, 
    0.07187001, 0.1932836, 0.1420941, 0.08495407, 0.1280567, 0.05451049, 
    0.1320398, 0.1196709, 0.179706, 0.02708191, 0.07411777, 0.006050439, 
    0.0001030575, 0.01022759, 0.0723343, 0.06106587, 0.1778834, 0.1181752, 
    0.05550461, 0.05238127, 0.009798413, 3.663285e-06, -1.016026e-05,
  0.04917599, 0.01432708, 0.01278742, 0.01186951, 0.004580276, 0.01153666, 
    0.009283788, 0.09243415, 0.167446, 0.1585075, 0.1743858, 0.1682487, 
    0.08464341, 0.1529548, 0.2073649, 0.2043886, 0.1477943, 0.1200627, 
    0.03753597, 0.0036328, 0.09166248, 0.06189446, 0.08705463, 0.06902176, 
    0.1520445, 0.0679186, 0.09246371, 0.05950671, 0.03105394,
  0.1581659, 0.1485366, 0.1755555, 0.1191603, 0.0975391, 0.1192283, 
    0.07200482, 0.02466057, 0.1214942, 0.2139429, 0.1847848, 0.1820257, 
    0.1614748, 0.2045141, 0.1630146, 0.1282702, 0.1034935, 0.1285091, 
    0.1334814, 0.04634234, 0.08959398, 0.1146422, 0.119058, 0.1343956, 
    0.1318298, 0.1720404, 0.1777551, 0.1803966, 0.1934233,
  0.1910457, 0.1444605, 0.1238013, 0.07303328, 0.08537178, 0.1435922, 
    0.1469965, 0.09431568, 0.1007916, 0.1566227, 0.1837655, 0.1812296, 
    0.07227978, 0.1569427, 0.1572055, 0.1445143, 0.1093876, 0.1289233, 
    0.04979781, 0.0989067, 0.1060703, 0.1458894, 0.1361976, 0.08954518, 
    0.1548018, 0.1108386, 0.1159911, 0.09448527, 0.09198714,
  0.0523092, 0.04088208, 0.02090039, 0.02066852, 0.03474085, 0.04470788, 
    0.06311258, 0.0782124, 0.070738, 0.0861817, 0.135334, 0.1000123, 
    0.1321457, 0.1176318, 0.131289, 0.07543126, 0.07655257, 0.04430371, 
    0.0301475, 0.08028389, 0.09286984, 0.1171586, 0.06146247, 0.01627709, 
    0.06627928, 3.120982e-05, 0.0006580051, 0.09962541, 0.08625436,
  0.01318395, 0.01731147, 0.02575401, 0.0296526, 0.02126958, 0.02744657, 
    0.01519262, 0.01692263, 0.01976075, 0.01751183, 0.0130963, 0.004891935, 
    -0.0007244991, 0.0101839, 0.008196753, 0.009362426, 0.01161831, 
    0.02201113, 0.0138253, 0.02719108, 0.06978572, 0.07861553, 0.03554647, 
    -0.0001950899, -0.001048622, -0.0001084304, -0.0005087229, 0.001784202, 
    0.01382067,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001576696, -7.60969e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.418303e-07, -1.078852e-05, 
    0.000857948, 0.0005736649, 0, -0.000128098, 0.001762262, 0.0003706609, 
    0.0004230943, -1.364229e-05, 0.0003435969, -0.0001569057, 0, 0, 
    6.326837e-05, 0, 0,
  0.004397072, 0.002481357, 4.893167e-05, 0.001046587, 0.005912405, 
    0.006111207, 0.008751845, 0.002203167, 0.002246658, 0.002508991, 
    0.00512232, 0.005516317, 0.004952817, 0.01018579, 0.01324214, 0.02084274, 
    0.01308754, 0.005004968, 0.007325562, 0.01490483, 0.01689057, 0.01288763, 
    0.004953873, 0.004521598, 0.008926987, 0.007148708, 0.0004136061, 
    0.003000357, 0.003781075,
  0.05950706, 0.02677288, 0.0348588, 0.03716942, 0.1055752, 0.0801734, 
    0.0608962, 0.03330999, 0.03291526, 0.02530312, 0.02666495, 0.01420421, 
    0.01176949, 0.02883108, 0.0602821, 0.03441405, 0.04178201, 0.03391395, 
    0.03972496, 0.01636881, 0.04381773, 0.05076911, 0.07838196, 0.05266299, 
    0.05879704, 0.07543761, 0.06389499, 0.06776139, 0.05490833,
  0.1524615, 0.09782425, 0.07175577, 0.1441789, 0.05962276, 0.07475932, 
    0.08423696, 0.05244317, 0.03697307, 0.02228534, 0.02945368, 0.04161005, 
    0.03595209, 0.03719822, 0.06430028, 0.1098301, 0.05011661, 0.1088674, 
    0.1388673, 0.1612168, 0.1812414, 0.1681363, 0.1478288, 0.06942293, 
    0.1382792, 0.1546752, 0.1738597, 0.1490236, 0.1714213,
  0.0005321497, 0.00339365, 0.01105452, 0.006757443, 0.02833639, 0.01653553, 
    0.007810113, 0.004567026, 0.003593447, 0.01168141, 0.008375325, 
    0.004883604, 0.01135535, 0.001590142, 0.01445773, 0.05798753, 0.1620449, 
    0.1693907, 0.1079301, 0.06834288, 0.04351912, 0.02648742, 0.007597956, 
    0.005090264, 0.0263343, 0.06892507, 0.05725866, 0.02662087, 0.004917054,
  2.872438e-07, 6.369384e-07, 2.435251e-07, -6.04469e-11, 0.0002367875, 
    -8.042961e-07, -3.845637e-06, 0.003140393, 0.005363508, 5.874623e-06, 
    3.625292e-05, 9.928528e-06, -1.09678e-06, 0.007179117, 0.04243454, 
    0.04039788, 0.03398066, 0.01046814, 0.004379372, 9.595974e-07, 
    6.365386e-09, 3.751872e-07, 9.159891e-07, 4.200922e-06, 0.006651593, 
    0.01050667, 0.001339691, 0.00389436, 7.182921e-05,
  3.593274e-06, 3.877416e-06, 1.74016e-06, 6.286783e-06, -7.987993e-05, 
    0.004078362, 0.06663999, 0.0965941, 0.02327019, 0.00492268, 0.003389982, 
    0.04509651, 0.02083188, 0.03650397, 0.01905468, 0.01467388, 0.0002614992, 
    2.279163e-05, 6.024515e-10, 8.685974e-07, 1.529329e-06, 3.040942e-07, 
    5.314599e-07, 0.001095464, 0.01288164, 0.001660995, 3.745704e-06, 
    2.488256e-07, 1.589121e-07,
  0.001840724, 0.09168343, 0.05728814, 0.00081777, 0.000553575, 0.07322556, 
    0.05320028, 0.09703535, 0.2277318, 0.2150259, 0.08547147, 0.1361219, 
    0.2065966, 0.0701696, 0.02838513, 0.002558089, 9.214054e-05, 
    -2.581544e-07, 8.654417e-06, 9.662195e-06, 6.119166e-05, 0.003850649, 
    0.02968196, 0.06020966, 0.01024523, 0.001501934, 0.0006800005, 
    0.006025835, 0.01136085,
  0.2360838, 0.2906965, 0.1934219, 0.1142433, 0.001925179, 0.004794751, 
    0.05466418, 0.07812817, 0.09368196, 0.02618493, 0.03812883, 0.08735938, 
    0.1830045, 0.08364324, 0.08533937, 0.08413455, 0.06651117, 0.08697597, 
    0.06699505, 0.1064623, 0.1482295, 0.1603829, 0.2054297, 0.06244352, 
    0.03975703, 0.0452202, 0.07097897, 0.1520425, 0.2565956,
  9.699936e-05, 0.002336568, 0.007082445, 0.0667285, 0.1085222, 0.1179429, 
    0.2216298, 0.06189752, 0.2599495, 0.07776125, 0.155841, 0.1510594, 
    0.1392831, 0.1519876, 0.1277823, 0.04648051, 0.003760101, 1.438761e-06, 
    0.006537815, 0.01089749, 0.0426277, 0.09808116, 0.03500693, 0.02210443, 
    0.0230446, 0.005748101, 0.001799981, 0.0002059871, 0.001774105,
  8.088935e-08, 2.611094e-10, -1.993298e-09, 0.002081407, 0.003395203, 
    0.01098161, 0.06905915, 0.1807156, 0.1461024, 0.06901272, 0.1143851, 
    0.0450839, 0.1226298, 0.1055337, 0.1699678, 0.02957489, 0.0514866, 
    0.002976731, 7.156515e-05, 0.01304876, 0.05510745, 0.04124178, 0.1426828, 
    0.103708, 0.04453804, 0.03881684, 0.003511709, 3.655822e-07, -3.188077e-05,
  0.03957182, 0.01559626, 0.01113146, 0.01054487, 0.006315151, 0.01364279, 
    0.01786758, 0.1084201, 0.1729277, 0.1441258, 0.1672202, 0.1448766, 
    0.09145708, 0.1531587, 0.1879729, 0.1960841, 0.1281107, 0.1049774, 
    0.03892092, 0.002935334, 0.06847073, 0.06189171, 0.07071337, 0.05681035, 
    0.1290107, 0.05826005, 0.08167831, 0.05204985, 0.01910802,
  0.1540627, 0.1464957, 0.1706902, 0.1047384, 0.08503784, 0.1174405, 
    0.07312879, 0.05979828, 0.1698706, 0.2076505, 0.1546543, 0.1525947, 
    0.1430204, 0.1846706, 0.139421, 0.1226891, 0.1084064, 0.1321692, 
    0.1336779, 0.06370793, 0.08301391, 0.1040314, 0.1041915, 0.1280814, 
    0.1100312, 0.14755, 0.1520697, 0.1737489, 0.1718022,
  0.1922713, 0.1500699, 0.1588079, 0.1373883, 0.1266594, 0.1608177, 
    0.2375687, 0.1454352, 0.1411185, 0.2057131, 0.2072295, 0.1811547, 
    0.09245512, 0.1502505, 0.1485576, 0.1713879, 0.1124042, 0.1895134, 
    0.1892698, 0.1657672, 0.1215142, 0.149033, 0.1406846, 0.1159427, 0.20767, 
    0.2225232, 0.1407548, 0.1522172, 0.1779751,
  0.1339814, 0.1409914, 0.09225906, 0.1102489, 0.1474472, 0.1322815, 
    0.1577147, 0.1971391, 0.1626604, 0.1433608, 0.1577159, 0.1401641, 
    0.1753901, 0.1994918, 0.206114, 0.1269061, 0.1235646, 0.1455526, 
    0.1565108, 0.2191488, 0.1624746, 0.1440634, 0.08907082, 0.04062026, 
    0.1333281, 0.006719582, 0.0009840353, 0.1988278, 0.1702804,
  0.1000201, 0.1129673, 0.1037187, 0.1242274, 0.1314671, 0.08813009, 
    0.06946573, 0.06707112, 0.06559625, 0.0663556, 0.1043048, 0.0789195, 
    0.04540099, 0.05624126, 0.06082413, 0.05044373, 0.08919737, 0.1499788, 
    0.1835629, 0.1593088, 0.1509408, 0.1641224, 0.1133984, 0.06118749, 
    0.04156967, 0.002403719, -0.001637875, 0.02265244, 0.07269236,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.966308e-06, 3.954257e-05, 0, 0, 
    -7.339196e-05, 0.001717396, -2.002164e-05, 0, 0, 0.0008743581, 
    0.0001498518, 0, 0, 0, 0, 0,
  -6.673887e-06, -0.0001225499, 0.004407434, 0.0004522294, -2.115342e-05, 0, 
    0, 0, 0, 0, 0, 0.0001613803, -7.284074e-05, 3.860724e-05, 0.001269291, 
    0.00258993, 0.005204106, 0.001823067, 0.006399679, 0.007666904, 
    0.005383106, 0.002408713, 0.01007253, 0.0003931228, 0.00106949, 
    0.0001381222, 0.001306928, -1.174056e-05, -4.409662e-05,
  0.03730453, 0.02439343, 0.0141285, 0.02081248, 0.02589918, 0.03269396, 
    0.0395546, 0.03702952, 0.022902, 0.01191818, 0.02831407, 0.02429654, 
    0.02785787, 0.04671717, 0.05687057, 0.06590237, 0.05290428, 0.05956057, 
    0.02802053, 0.03506, 0.02813819, 0.0184613, 0.01435566, 0.02214114, 
    0.03643076, 0.03844408, 0.02516863, 0.02484151, 0.03475471,
  0.1135175, 0.1039222, 0.1806905, 0.175638, 0.2053185, 0.18462, 0.1243829, 
    0.09359236, 0.1017689, 0.09204422, 0.09069327, 0.1050437, 0.08519804, 
    0.09716427, 0.179031, 0.1405004, 0.09999307, 0.08308052, 0.08569191, 
    0.05479094, 0.09322095, 0.1032615, 0.1312664, 0.09911008, 0.120668, 
    0.1677305, 0.1180037, 0.1122983, 0.100388,
  0.1995132, 0.1111455, 0.07899766, 0.1491158, 0.05922842, 0.07969112, 
    0.09390283, 0.06727895, 0.05455614, 0.04779306, 0.05949089, 0.09038791, 
    0.05363257, 0.09072089, 0.1044237, 0.162975, 0.07786053, 0.1335919, 
    0.1508779, 0.19253, 0.1946718, 0.1894838, 0.1607608, 0.1052423, 
    0.1216304, 0.1305505, 0.1526317, 0.1516858, 0.1952522,
  0.0004839799, 0.001874781, 0.008901311, 0.003506332, 0.03002507, 
    0.02123724, 0.007999197, 0.004113511, 0.002010274, 0.01349831, 
    0.009695618, 0.003311531, 0.01164391, 0.001808749, 0.02167146, 
    0.06268921, 0.1735193, 0.1635948, 0.09927793, 0.0627775, 0.03338136, 
    0.01292633, 0.002717373, 0.004314615, 0.03067938, 0.07480909, 0.06240898, 
    0.02549133, 0.004551909,
  1.197804e-08, 1.089291e-07, 9.325765e-08, -1.927389e-07, 0.0002107932, 
    -3.035203e-05, 1.019446e-06, 0.01621594, 0.001213025, 0.0001541064, 
    0.001975695, 0.000612586, 2.556244e-06, 0.01524087, 0.04310435, 
    0.04091518, 0.03889235, 0.005887719, 0.00260725, 1.992901e-06, 
    -2.989411e-10, -3.021378e-06, 8.694986e-08, 6.983544e-07, 0.006054608, 
    0.004115786, 0.0006782926, 4.747631e-05, 6.446838e-07,
  1.123191e-06, 9.363872e-07, 2.515738e-07, 1.014711e-05, 0.001669859, 
    0.004433533, 0.06989144, 0.09691687, 0.02024787, 0.005512836, 
    0.002216994, 0.03592025, 0.03135474, 0.03545864, 0.01400515, 0.01441945, 
    0.0002965351, 3.780077e-06, 0, 2.348591e-07, 3.489621e-07, 1.452779e-07, 
    2.179388e-06, 0.001441022, 0.01046283, 0.0006457567, 1.317624e-06, 
    8.304392e-08, 1.104044e-07,
  0.001826897, 0.0566534, 0.04254729, 0.004235878, 0.000798521, 0.06496943, 
    0.03183007, 0.05099664, 0.1569415, 0.1965748, 0.05852715, 0.1210538, 
    0.200898, 0.06131519, 0.0264604, 0.002190944, 0.000116988, -3.927756e-06, 
    7.564087e-06, -2.495424e-06, 1.178253e-07, 0.001305913, 0.02306548, 
    0.03417137, 0.008455141, 0.001044386, 3.270166e-05, 0.0001208501, 
    0.00924681,
  0.2072501, 0.2396829, 0.1618402, 0.1161329, 0.003889784, 0.004142862, 
    0.04038938, 0.03234537, 0.08258659, 0.01709256, 0.02519947, 0.06412474, 
    0.1565215, 0.06568605, 0.06598361, 0.08138928, 0.05956625, 0.08822994, 
    0.0712591, 0.1203566, 0.1298195, 0.1321453, 0.172688, 0.04961558, 
    0.03491511, 0.03562474, 0.05543274, 0.1491918, 0.2505225,
  8.945199e-05, 0.001809278, 0.006561426, 0.07004596, 0.1293937, 0.1520816, 
    0.1911254, 0.04072695, 0.2520305, 0.05605187, 0.135566, 0.128417, 
    0.0907849, 0.1161371, 0.08383543, 0.03775586, 0.001062183, 2.724497e-06, 
    0.006146527, 0.007078793, 0.0417238, 0.07481125, 0.02253665, 0.01268432, 
    0.01572401, 0.003705358, 0.0001210233, 0.0002368999, 0.002025678,
  2.158603e-08, -1.535431e-08, 0, 0.00971524, 0.004154043, 0.009884096, 
    0.06189115, 0.1644423, 0.1500758, 0.05216826, 0.1046344, 0.03633882, 
    0.1128507, 0.09072129, 0.1514511, 0.03356532, 0.039154, 0.002033681, 
    2.760226e-05, 0.02264766, 0.04241696, 0.02601857, 0.1074481, 0.07893337, 
    0.03133788, 0.02555263, 0.0008830196, 2.974591e-08, 3.183113e-05,
  0.03286557, 0.01681911, 0.01153743, 0.007358694, 0.01028563, 0.01915797, 
    0.04151408, 0.116304, 0.1746328, 0.1261799, 0.1673331, 0.1282537, 
    0.08537918, 0.1412837, 0.1970244, 0.1807003, 0.1181693, 0.09739088, 
    0.02932803, 0.006367447, 0.05691256, 0.05787464, 0.05405805, 0.04787304, 
    0.1062047, 0.05543013, 0.06886721, 0.04889517, 0.01734955,
  0.1521194, 0.1248456, 0.1552279, 0.0889981, 0.07586198, 0.1039651, 
    0.06594214, 0.06666718, 0.1806097, 0.1900881, 0.1325269, 0.1337435, 
    0.1246719, 0.1765092, 0.1273054, 0.1201296, 0.1048403, 0.1270175, 
    0.1274852, 0.05527834, 0.0680953, 0.09752911, 0.09455576, 0.1082319, 
    0.0971908, 0.1271075, 0.1536356, 0.1613493, 0.1482605,
  0.172043, 0.172043, 0.1466335, 0.1390983, 0.1303402, 0.163679, 0.2648624, 
    0.1649648, 0.1543428, 0.207602, 0.1900213, 0.1661946, 0.08335441, 
    0.1424417, 0.1371984, 0.1726816, 0.1758032, 0.2269469, 0.259591, 
    0.1550859, 0.130114, 0.1334073, 0.1332576, 0.1199985, 0.2102975, 
    0.2330159, 0.1508589, 0.1658643, 0.197136,
  0.141077, 0.1862262, 0.1885049, 0.1648149, 0.1950458, 0.1859673, 0.1846538, 
    0.2458209, 0.1983463, 0.1505373, 0.1826362, 0.1725349, 0.1661942, 
    0.2007515, 0.2290333, 0.1267684, 0.1838113, 0.1838324, 0.1737166, 
    0.254885, 0.215932, 0.1480664, 0.104182, 0.1086551, 0.15404, 0.05842837, 
    0.01224808, 0.2328941, 0.1752226,
  0.1848632, 0.2111472, 0.1812902, 0.1812853, 0.1702554, 0.1616198, 
    0.1348932, 0.1181523, 0.1173907, 0.1044145, 0.1221604, 0.1076428, 
    0.07246952, 0.1081081, 0.09844883, 0.1257842, 0.1780595, 0.2288978, 
    0.251231, 0.2267116, 0.1910788, 0.2179543, 0.1538327, 0.1121891, 
    0.09243228, 0.04779949, 0.03540738, 0.0825566, 0.1619688,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000241079, -8.225258e-05, 
    -7.147421e-05, 0, -5.846091e-05, 0.007907982, 0.0009808567, 
    -1.056048e-05, -5.368418e-06, 0.001298506, 0.003088747, -2.42743e-06, 0, 
    0, 0, 0,
  0.0006935099, 0.005641871, 0.0333344, 0.02015736, -7.492094e-05, 0, 
    0.0001199993, -3.441839e-06, 0, -1.985709e-05, -5.590743e-06, 
    0.0005505074, 0.0002099358, 0.02525862, 0.03212954, 0.02493228, 
    0.01923627, 0.0154977, 0.03651228, 0.03900137, 0.02245735, 0.0154778, 
    0.02471514, 0.00865043, 0.009683324, 0.01909878, 0.006430042, 
    0.001269524, 0.002377439,
  0.08322182, 0.08488113, 0.06543375, 0.06474315, 0.09171076, 0.1028912, 
    0.100209, 0.07978834, 0.06444497, 0.05084615, 0.06219498, 0.07851839, 
    0.128476, 0.1979357, 0.2009043, 0.2095363, 0.1783347, 0.1669684, 
    0.1006968, 0.08350999, 0.05983102, 0.05025724, 0.03892341, 0.05626486, 
    0.09669132, 0.1324554, 0.06252246, 0.09081084, 0.08057266,
  0.15278, 0.1443976, 0.2537076, 0.2374156, 0.2340118, 0.2075754, 0.1431083, 
    0.1362666, 0.1475112, 0.1232471, 0.1814065, 0.1890502, 0.1936894, 
    0.195493, 0.218317, 0.1556401, 0.1569853, 0.1529238, 0.1668876, 
    0.1060612, 0.1790283, 0.1757694, 0.1887678, 0.1588551, 0.1613915, 
    0.2057517, 0.1854583, 0.1594757, 0.1451712,
  0.1743276, 0.0920532, 0.08588684, 0.1455601, 0.06083515, 0.08217168, 
    0.09889111, 0.07089061, 0.06498033, 0.06603402, 0.0829026, 0.1175414, 
    0.08207548, 0.1133173, 0.1355205, 0.1619, 0.08250678, 0.1412102, 
    0.1392532, 0.1785981, 0.1896339, 0.1884828, 0.1702619, 0.1234316, 
    0.1060375, 0.107033, 0.1203934, 0.1480169, 0.1770896,
  -4.986567e-05, 0.0009116894, 0.004869009, 0.002038191, 0.03175587, 
    0.03625277, 0.008148258, 0.002862742, 1.588913e-05, 0.005429874, 
    0.01233415, 0.00327328, 0.01345033, 0.00580183, 0.02677979, 0.07520736, 
    0.1613813, 0.1651825, 0.1039333, 0.0619956, 0.0263527, 0.003790127, 
    0.0001789319, 0.002165949, 0.0333504, 0.08090113, 0.06974165, 0.02774673, 
    0.006027493,
  -6.261225e-10, 3.993313e-08, 6.520748e-08, 2.867226e-05, 7.747365e-05, 
    0.001296084, 4.157843e-08, 0.03073773, 3.570953e-05, 0.001123024, 
    0.001911957, 0.002226903, 0.0001616763, 0.01583736, 0.03791283, 
    0.05405007, 0.03373837, 0.002259352, 0.002387121, 1.809478e-06, 
    1.849325e-08, -2.759965e-06, 1.216526e-08, 2.403386e-07, 0.009355535, 
    0.00485927, 4.379654e-05, 1.150709e-06, 2.696032e-08,
  2.048146e-07, 1.08803e-06, 3.157747e-10, 1.214344e-05, 0.002920916, 
    0.004688977, 0.07867543, 0.09226315, 0.01983917, 0.009336563, 
    0.002298783, 0.02441747, 0.0393643, 0.04225665, 0.01127102, 0.01909573, 
    0.0003251958, -2.599396e-05, 0, 3.428823e-08, 1.12143e-08, 1.024773e-09, 
    2.315435e-06, 0.001276107, 0.008051983, 0.0007245177, 4.061342e-07, 
    8.550411e-08, 7.283629e-08,
  0.01316639, 0.04268994, 0.03321741, 0.006033272, 0.001302828, 0.05406058, 
    0.02001602, 0.02557763, 0.09553546, 0.2009788, 0.04414327, 0.1212886, 
    0.2052043, 0.0560339, 0.02108529, 0.002458443, 0.0001289025, 
    -3.224352e-06, 0.0001269463, -1.019326e-05, 7.101554e-06, 0.009448137, 
    0.02586926, 0.02168685, 0.009426582, 0.001344554, 0.0002919585, 
    5.698885e-05, 0.003674733,
  0.1840595, 0.2031878, 0.1485004, 0.1202163, 0.007003898, 0.004112548, 
    0.03791111, 0.01500661, 0.0687246, 0.0117378, 0.01965877, 0.04728489, 
    0.134816, 0.05210716, 0.0562978, 0.07887921, 0.05739061, 0.09645845, 
    0.08220027, 0.1350087, 0.137949, 0.109966, 0.1582262, 0.04251929, 
    0.0295231, 0.03025753, 0.05179677, 0.1605715, 0.256225,
  9.273747e-05, 0.002165618, 0.01155929, 0.09057176, 0.1203349, 0.1326197, 
    0.1954015, 0.03031765, 0.2260349, 0.04496884, 0.1270187, 0.1145179, 
    0.06851824, 0.09244154, 0.04990084, 0.02911603, 9.397319e-05, 
    4.615664e-06, 0.00323839, 0.008912949, 0.04267913, 0.06656167, 
    0.01496562, 0.009662999, 0.01147816, 0.002396337, 5.808919e-05, 
    0.0001541703, 0.003602583,
  0.0001234696, -4.685878e-05, 0, 0.01787416, 0.003208356, 0.007316052, 
    0.05294061, 0.1652808, 0.1600591, 0.05363588, 0.09262305, 0.03824962, 
    0.1081327, 0.082932, 0.1214477, 0.02743408, 0.0345043, 0.003532154, 
    3.499819e-05, 0.0114637, 0.03325596, 0.01697704, 0.07970203, 0.05431052, 
    0.01869736, 0.01436344, 0.0001966142, 1.361496e-07, 0.0006834124,
  0.02468794, 0.01625352, 0.01187448, 0.006731449, 0.0193198, 0.0174642, 
    0.06090338, 0.1106877, 0.1574264, 0.1102186, 0.1649397, 0.1164531, 
    0.07998785, 0.1563982, 0.1872091, 0.1687163, 0.1169955, 0.09437397, 
    0.02538936, 0.01028885, 0.04466805, 0.06688221, 0.04330962, 0.04014271, 
    0.08410516, 0.05005316, 0.05367751, 0.0439583, 0.01273175,
  0.1498426, 0.1163637, 0.1396686, 0.07697837, 0.07054394, 0.09559458, 
    0.06346636, 0.05600827, 0.1906483, 0.1765099, 0.12436, 0.1160643, 
    0.1255338, 0.1577819, 0.11612, 0.1116671, 0.1020301, 0.1238575, 
    0.1355711, 0.04581798, 0.05510353, 0.102685, 0.09616188, 0.1046396, 
    0.09568387, 0.1251278, 0.1492266, 0.149738, 0.1314144,
  0.1546498, 0.1486998, 0.1336683, 0.1297923, 0.1146059, 0.1619601, 
    0.2451216, 0.1474513, 0.1334703, 0.1837231, 0.1632635, 0.1501383, 
    0.0827097, 0.1375731, 0.1391762, 0.1751207, 0.1940423, 0.2412053, 
    0.2990135, 0.1469831, 0.1189622, 0.1304087, 0.132872, 0.1174116, 
    0.202176, 0.2437797, 0.1504546, 0.1660884, 0.2064854,
  0.1348678, 0.1755184, 0.1925392, 0.1474751, 0.1828814, 0.1761285, 
    0.1852649, 0.2366972, 0.1821662, 0.1430173, 0.1714447, 0.1719122, 
    0.1522477, 0.2000677, 0.2321351, 0.1281385, 0.1839551, 0.1868618, 
    0.1634911, 0.2442329, 0.2306648, 0.1627996, 0.09810311, 0.1466127, 
    0.1738383, 0.1587804, 0.05396006, 0.2166273, 0.1623545,
  0.1869071, 0.2080676, 0.1770074, 0.1791587, 0.1651532, 0.1552964, 
    0.1251012, 0.1210527, 0.120816, 0.1176012, 0.1396204, 0.1187774, 
    0.1034502, 0.138827, 0.1403006, 0.1687705, 0.2003849, 0.2284802, 
    0.2617823, 0.2354646, 0.1871902, 0.2320631, 0.1766787, 0.1156275, 
    0.1408938, 0.06191466, 0.06577811, 0.1120813, 0.1691887,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007731061, 0.01338651, 
    0.008684147, 0.004297201, 0.002602088, 0.01111273, 0.003268472, 
    0.0007665544, -2.615899e-05, 0.001838654, 0.02220652, 0.02118701, 
    -0.003541231, 9.893411e-06, -0.0002151148, 0,
  0.05021225, 0.0550763, 0.052539, 0.04061257, -0.000335602, -0.0002388426, 
    0.004359111, 0, -4.595448e-05, 0.0001950811, 0.0005033527, 0.001499741, 
    0.02090226, 0.1336062, 0.1425794, 0.1336455, 0.1366726, 0.1095579, 
    0.09383069, 0.1171554, 0.08715177, 0.07877129, 0.09365399, 0.04142141, 
    0.08689101, 0.06255849, 0.03834151, 0.02102597, 0.06124967,
  0.1147387, 0.1182392, 0.1122863, 0.130729, 0.1895229, 0.1712148, 0.1451919, 
    0.1376263, 0.1033475, 0.1200802, 0.1504373, 0.2085688, 0.2402225, 
    0.2852687, 0.2504256, 0.2377324, 0.2480738, 0.2475546, 0.1771793, 
    0.1466745, 0.1288253, 0.1172814, 0.1370063, 0.1596035, 0.227361, 
    0.1903334, 0.1348178, 0.1587149, 0.1382966,
  0.1551456, 0.1442269, 0.25781, 0.2258376, 0.2137802, 0.186726, 0.1514861, 
    0.1607412, 0.1764894, 0.1757013, 0.2190571, 0.2244581, 0.2100366, 
    0.1805952, 0.2179791, 0.1492258, 0.1517813, 0.149255, 0.16989, 0.1317765, 
    0.209851, 0.2073869, 0.2298404, 0.1941708, 0.1740211, 0.1968115, 
    0.1876254, 0.1641379, 0.1651996,
  0.1588641, 0.09104899, 0.07653234, 0.1364143, 0.06353043, 0.08317183, 
    0.09525099, 0.07965324, 0.07066463, 0.06002236, 0.07642032, 0.1075875, 
    0.07410953, 0.1117008, 0.1190291, 0.1510099, 0.07794132, 0.1385261, 
    0.1294943, 0.1601982, 0.1917494, 0.193245, 0.1795193, 0.1360287, 
    0.1060045, 0.0889996, 0.1062014, 0.1371247, 0.1578319,
  0.0005913929, 0.0003370011, 0.001812955, 0.002218735, 0.03073161, 
    0.05581735, 0.009197685, 0.0003748735, 4.52069e-05, 0.002171547, 
    0.006058118, 0.005517698, 0.01395685, 0.01088133, 0.03583868, 0.08008806, 
    0.1492108, 0.1790181, 0.1045433, 0.04873534, 0.02235759, 0.002670203, 
    0.0001008675, 0.002556924, 0.03449322, 0.084025, 0.06677817, 0.02589174, 
    0.009260315,
  4.37308e-09, 6.959036e-09, 2.995941e-07, 7.631932e-05, 8.441681e-06, 
    0.005626902, 1.496908e-06, 0.03498174, 0.001486786, 0.005749656, 
    0.009487594, 0.001620526, 0.0001835533, 0.01618088, 0.03924833, 
    0.06930504, 0.0320015, 0.003327806, 0.007260816, 2.351283e-06, 
    -2.287801e-08, -1.678319e-07, 5.207531e-09, 7.563622e-08, 0.006704257, 
    0.01101395, -3.095401e-05, 1.531503e-08, 2.222152e-08,
  3.64222e-07, 4.057732e-06, 3.101417e-08, 0.0006592069, 0.008271739, 
    0.005429678, 0.06059083, 0.08470938, 0.01777893, 0.01411417, 0.003680319, 
    0.0143118, 0.05367226, 0.04793102, 0.01525747, 0.01759917, 0.0006316271, 
    -2.134646e-05, 0, 6.216936e-09, 6.600431e-09, 1.048598e-08, 2.343053e-06, 
    0.001086316, 0.006266785, 0.0004453812, 3.243106e-08, 1.70872e-08, 
    1.219518e-08,
  0.01092428, 0.04052401, 0.02923265, 0.009041323, 0.006346802, 0.0550125, 
    0.01398224, 0.01870218, 0.0692654, 0.1925696, 0.03576284, 0.1192533, 
    0.2108419, 0.0566257, 0.01756205, 0.004940697, 0.000302098, 
    -8.626417e-06, 0.001555073, -4.960192e-05, 3.980388e-05, 0.007305774, 
    0.0286069, 0.01955466, 0.01044277, 0.003056797, 0.002221874, 0.001095634, 
    0.000776499,
  0.1749815, 0.1871258, 0.1521124, 0.1391586, 0.01540181, 0.004865299, 
    0.04644587, 0.008639463, 0.05965684, 0.01066776, 0.01571393, 0.03362929, 
    0.129463, 0.04598467, 0.04876446, 0.07108648, 0.06534213, 0.1017226, 
    0.1305537, 0.1375924, 0.1352243, 0.1035269, 0.1445063, 0.03814443, 
    0.02617433, 0.02880177, 0.05174116, 0.1740532, 0.266167,
  0.000211128, 0.002684746, 0.02470078, 0.08183411, 0.1161471, 0.1543122, 
    0.2203223, 0.03085215, 0.21568, 0.04331451, 0.1292064, 0.114146, 
    0.05905861, 0.08261477, 0.03220915, 0.02609418, 0.004756679, 
    2.261205e-06, 0.001650633, 0.01132028, 0.03530974, 0.0613891, 0.01249482, 
    0.008934841, 0.00884846, 0.001681244, 0.002684696, 0.0002005909, 
    0.004535872,
  0.003225423, 0.001691168, -2.810547e-10, 0.02877959, 0.004517831, 
    0.004854872, 0.04838199, 0.1715096, 0.1669413, 0.04444511, 0.08711824, 
    0.04460576, 0.1043926, 0.07339537, 0.1106241, 0.02493965, 0.02931155, 
    0.01074789, -6.699593e-05, 0.01897048, 0.02360308, 0.01180102, 
    0.06286358, 0.03927306, 0.01399034, 0.008235549, 0.0002456353, 
    2.993203e-08, 0.002164525,
  0.02025859, 0.01550618, 0.0126927, 0.006858883, 0.03938475, 0.01336241, 
    0.05881206, 0.0892249, 0.1333262, 0.1111076, 0.1637847, 0.09370887, 
    0.06881047, 0.1123843, 0.1834033, 0.1590047, 0.1151773, 0.07651407, 
    0.01615107, 0.002027672, 0.05730879, 0.06470396, 0.03418169, 0.03357507, 
    0.07318301, 0.0423445, 0.04952621, 0.04332079, 0.008389717,
  0.1306699, 0.1092205, 0.1298568, 0.06969014, 0.06691546, 0.08985101, 
    0.05503215, 0.05690051, 0.1687686, 0.166198, 0.1100991, 0.1034059, 
    0.1050704, 0.1443976, 0.1153161, 0.08631642, 0.103977, 0.1186882, 
    0.1315617, 0.03753505, 0.04924467, 0.1111946, 0.08969695, 0.0915705, 
    0.0970736, 0.1239729, 0.1464899, 0.1387997, 0.1352522,
  0.1414118, 0.1278757, 0.1247686, 0.1237577, 0.1052731, 0.1580046, 
    0.2246147, 0.1309609, 0.1131377, 0.1600998, 0.1491907, 0.1380307, 
    0.08435227, 0.1384292, 0.1395059, 0.1726562, 0.1903696, 0.2343692, 
    0.2950946, 0.14989, 0.1135994, 0.1242252, 0.1359866, 0.1173919, 
    0.1959642, 0.2591948, 0.1560102, 0.1701794, 0.1867932,
  0.1382399, 0.1690697, 0.1927018, 0.1462004, 0.1825997, 0.1550044, 
    0.1762928, 0.2205947, 0.1624331, 0.1415813, 0.1720714, 0.1713213, 
    0.1497796, 0.2052795, 0.2285289, 0.1202922, 0.1819881, 0.1838577, 
    0.1542374, 0.2281739, 0.224223, 0.1672805, 0.1315577, 0.1404307, 
    0.1791784, 0.2179377, 0.1206905, 0.2173372, 0.1656968,
  0.1855395, 0.2033163, 0.1616935, 0.15448, 0.1537594, 0.1567847, 0.1228403, 
    0.1195725, 0.1173799, 0.1258966, 0.1469205, 0.1152472, 0.1176658, 
    0.1668169, 0.1819571, 0.1934912, 0.2040324, 0.2227869, 0.2563138, 
    0.2250512, 0.1814315, 0.2344024, 0.1910055, 0.1173474, 0.1550665, 
    0.07308903, 0.08842936, 0.1037818, 0.1523278,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -2.017528e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04213101, 0.07063045, 
    0.05622707, 0.04257831, 0.02994414, 0.0243081, 0.01439363, 0.001991927, 
    -8.963331e-05, 0.01094984, 0.1257322, 0.09377091, 0.02954368, 0.02063587, 
    0.0004303431, 0.0002734868,
  0.1053381, 0.1134131, 0.1069114, 0.04725285, -0.0002012994, -0.0004974518, 
    0.03580968, -0.0001472423, -0.0004665057, 0.001758565, 0.001672964, 
    0.004016793, 0.09682083, 0.2082567, 0.2221335, 0.2038148, 0.2028071, 
    0.1638275, 0.1502256, 0.1583739, 0.1364465, 0.1667528, 0.2235748, 
    0.1481673, 0.1845248, 0.1404655, 0.1365447, 0.114873, 0.1339999,
  0.1793348, 0.1783254, 0.1652301, 0.1978565, 0.2297184, 0.2214676, 
    0.1781671, 0.1889763, 0.1498896, 0.1882421, 0.2613105, 0.2770959, 
    0.2998163, 0.2895541, 0.2446551, 0.2232195, 0.2423694, 0.2343588, 
    0.178212, 0.1751217, 0.1764053, 0.1964361, 0.2446479, 0.2234763, 
    0.2792574, 0.255091, 0.2012429, 0.2184366, 0.2144937,
  0.1633435, 0.1547429, 0.2579213, 0.2294974, 0.2082466, 0.1759976, 
    0.1505632, 0.1758828, 0.1824671, 0.1972685, 0.2361997, 0.2251767, 
    0.2020642, 0.1629822, 0.2099282, 0.1506517, 0.1354641, 0.1441787, 
    0.1589072, 0.1361306, 0.2062519, 0.1891936, 0.2271658, 0.2177388, 
    0.1742902, 0.1944742, 0.1863993, 0.1672759, 0.1704397,
  0.1492942, 0.09283094, 0.07514809, 0.1351123, 0.06372879, 0.07644233, 
    0.1026425, 0.08318526, 0.06846985, 0.05810459, 0.07330035, 0.09743859, 
    0.07278991, 0.1019269, 0.1212275, 0.1426785, 0.0811711, 0.14022, 
    0.1202253, 0.1421054, 0.1901189, 0.1939722, 0.1749163, 0.1432651, 
    0.09928774, 0.08722779, 0.1005351, 0.1307786, 0.1382465,
  0.001382306, 0.0001154104, 0.005717108, 0.003503778, 0.02865396, 
    0.06007437, 0.007009478, -3.194659e-05, -2.628289e-05, 3.207892e-05, 
    0.0005901514, 0.01460734, 0.01771547, 0.01872858, 0.04276089, 0.08084251, 
    0.143728, 0.1899195, 0.1114443, 0.04883462, 0.02106916, 0.004466976, 
    7.117448e-05, 0.002726926, 0.03790952, 0.08613872, 0.06575933, 
    0.02472559, 0.01004387,
  2.281224e-08, 2.13104e-09, 2.271127e-07, 0.0001502309, 0.003895031, 
    0.007506207, -0.0002500105, 0.03108766, 0.0005477347, 0.007858762, 
    0.008008232, 0.0007194437, 4.804803e-05, 0.01862095, 0.05094281, 
    0.05925274, 0.03246717, 0.0003786823, 0.01319966, 3.294731e-06, 
    -2.676318e-07, 8.073674e-08, -5.95572e-11, 8.485399e-08, 0.004961497, 
    0.0171573, -0.0001091837, 1.817717e-09, 4.344367e-09,
  2.162909e-07, 2.473842e-05, 2.118391e-07, 0.0004387459, 0.01175133, 
    0.005946027, 0.05529086, 0.07790691, 0.02449867, 0.01943847, 0.002320073, 
    0.007613678, 0.06294125, 0.06035259, 0.01649104, 0.02192128, 0.001684236, 
    -4.963205e-05, -1.14164e-09, 2.330488e-09, 4.669034e-09, 6.245436e-08, 
    1.7705e-06, 0.001653672, 0.003685238, 0.0001652206, 3.271005e-10, 
    5.455668e-10, -2.03298e-10,
  0.01398394, 0.04975912, 0.03729644, 0.01876737, 0.01566244, 0.05107614, 
    0.01329495, 0.01529424, 0.06179528, 0.1888862, 0.03392649, 0.1197558, 
    0.2198789, 0.05837142, 0.01632616, 0.006646587, 0.001652411, 0.002131911, 
    0.002423591, 0.003647022, 0.0008547023, 0.001072459, 0.02729088, 
    0.01529999, 0.01315693, 0.008341128, 0.001557316, 0.004889564, 
    -6.114355e-05,
  0.1747165, 0.1807835, 0.148943, 0.1527444, 0.03244532, 0.007050105, 
    0.05080806, 0.007178905, 0.05722733, 0.011702, 0.01619371, 0.02667511, 
    0.1164682, 0.04008108, 0.04764795, 0.07806462, 0.06898433, 0.1100373, 
    0.1661948, 0.1654412, 0.1319687, 0.1146532, 0.1443455, 0.04130213, 
    0.02150945, 0.02904032, 0.05373242, 0.1793693, 0.2776839,
  0.001990864, 0.004481226, 0.02410092, 0.08016405, 0.09894562, 0.1310862, 
    0.2259894, 0.0364336, 0.2120701, 0.04337447, 0.1335675, 0.1195401, 
    0.05867016, 0.07129869, 0.02301857, 0.02147665, 0.002962241, 4.0684e-08, 
    0.006476287, 0.005949138, 0.03808877, 0.05531044, 0.01060468, 0.00814732, 
    0.006794967, 0.001409288, 0.001691767, 0.0006147701, 0.01140164,
  0.01685947, 0.001280454, -1.448917e-07, 0.04553905, 0.009994527, 
    0.00247478, 0.04934701, 0.1830907, 0.1821613, 0.04880621, 0.0814394, 
    0.0498398, 0.1116496, 0.06746907, 0.09894496, 0.02063514, 0.03487571, 
    0.00711883, 0.0005305754, 0.03504621, 0.01897096, 0.0141745, 0.05158876, 
    0.0288368, 0.01460815, 0.00459647, 0.0002628738, 8.000133e-10, 0.01946048,
  0.01641931, 0.01173723, 0.01380859, 0.007702702, 0.04047226, 0.007671059, 
    0.06840955, 0.06904881, 0.107717, 0.09814617, 0.1649618, 0.08268301, 
    0.06764201, 0.09776157, 0.1712258, 0.1428903, 0.1313545, 0.08093775, 
    0.01504821, 0.000375023, 0.0938707, 0.0689232, 0.03072752, 0.03141423, 
    0.06822208, 0.04196703, 0.04522986, 0.03183959, 0.006727709,
  0.1073646, 0.1039185, 0.1199495, 0.06420036, 0.06215216, 0.08884131, 
    0.044226, 0.05921057, 0.1587709, 0.1615224, 0.1013399, 0.09421334, 
    0.08736741, 0.1354868, 0.1135317, 0.09513295, 0.1103718, 0.1219937, 
    0.1253774, 0.02613583, 0.0522359, 0.1126927, 0.09683628, 0.09419154, 
    0.09695652, 0.1136437, 0.1426658, 0.1367961, 0.1259941,
  0.1471642, 0.1216641, 0.1207297, 0.1184354, 0.1005374, 0.1464598, 
    0.2063327, 0.1287247, 0.09986596, 0.133434, 0.1386027, 0.1311715, 
    0.08807075, 0.1496149, 0.1479226, 0.156358, 0.1891117, 0.219703, 
    0.3055292, 0.1422646, 0.1129208, 0.1241872, 0.1320133, 0.1493571, 
    0.1958974, 0.2677065, 0.1453621, 0.1830994, 0.2003821,
  0.1437893, 0.2018522, 0.2294597, 0.1567132, 0.1837903, 0.1467796, 
    0.1863656, 0.2293967, 0.1550056, 0.1467101, 0.1632291, 0.177751, 
    0.1755475, 0.2155163, 0.2339996, 0.1083749, 0.1803563, 0.1945074, 
    0.142634, 0.2193149, 0.216089, 0.1686124, 0.1312127, 0.1478495, 
    0.1675906, 0.2517973, 0.1637491, 0.2290867, 0.1630221,
  0.1811654, 0.1981502, 0.1520574, 0.1534996, 0.1416072, 0.1611995, 
    0.1204685, 0.1291588, 0.1109919, 0.126213, 0.1564315, 0.1248944, 
    0.1549763, 0.2329193, 0.2407206, 0.2369151, 0.2272313, 0.2270982, 
    0.2639585, 0.2209778, 0.1841839, 0.2337332, 0.1852232, 0.108792, 
    0.1640323, 0.09360406, 0.09992145, 0.09188247, 0.135106,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -0.0001257764, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004517217, 0.1086498, 
    0.1072079, 0.09273887, 0.08352949, 0.06924812, 0.06404485, 0.03062756, 
    0.005394268, 0.00125113, 0.03626431, 0.182825, 0.1542586, 0.1057045, 
    0.1103754, 0.01370537, 0.00189458,
  0.2031802, 0.2316645, 0.1711847, 0.09722656, 0.002577776, 0.001549833, 
    0.09245005, -0.001832861, -2.624889e-05, 0.001807084, 0.004325802, 
    0.003306349, 0.1820036, 0.2738171, 0.2445834, 0.2413737, 0.2383773, 
    0.1788616, 0.1828687, 0.2086688, 0.2167278, 0.2323079, 0.2781018, 
    0.2657782, 0.2575648, 0.1946231, 0.1933631, 0.1650236, 0.1798484,
  0.2211596, 0.218961, 0.2321694, 0.2582201, 0.256182, 0.2411847, 0.2175817, 
    0.2353474, 0.1904013, 0.2512496, 0.3306121, 0.3244293, 0.3015909, 
    0.2728876, 0.235787, 0.2195393, 0.2326967, 0.226458, 0.1832281, 0.175146, 
    0.1857893, 0.2182111, 0.2608189, 0.2263175, 0.276595, 0.2509561, 
    0.1943963, 0.2403843, 0.2475021,
  0.1802362, 0.1737904, 0.2346375, 0.2188384, 0.197476, 0.1712528, 0.1510186, 
    0.1911223, 0.1854836, 0.2159254, 0.2416951, 0.2188376, 0.1951494, 
    0.1442456, 0.2087345, 0.1513617, 0.1317654, 0.1411975, 0.1659551, 
    0.1257192, 0.1938662, 0.1801527, 0.220755, 0.2188346, 0.1687631, 
    0.1830019, 0.1660109, 0.1604792, 0.1699503,
  0.1448865, 0.09663476, 0.06934366, 0.1273188, 0.06663312, 0.0743724, 
    0.1016809, 0.07516351, 0.07200097, 0.05445617, 0.06700163, 0.09147621, 
    0.07636442, 0.10639, 0.133574, 0.1572805, 0.08741543, 0.1359938, 
    0.1122785, 0.1398877, 0.1689675, 0.188785, 0.1680558, 0.1414384, 
    0.09320986, 0.0924842, 0.08836073, 0.1359858, 0.1471939,
  0.001702424, 2.012316e-05, 0.01495917, 0.005561565, 0.02971068, 0.06561732, 
    0.008756144, 0.001151776, -3.982409e-05, -0.0001021327, 0.0007875012, 
    0.02709485, 0.02652593, 0.02787217, 0.04357263, 0.08441633, 0.1470649, 
    0.1922679, 0.1164087, 0.04484056, 0.02961615, 0.00762317, 0.0001516015, 
    0.005608802, 0.05149681, 0.09034198, 0.0673257, 0.02090664, 0.01115674,
  4.162951e-08, 8.600706e-09, -4.0377e-07, 0.0001735085, 0.009837197, 
    0.007886432, 0.0007439344, 0.02138048, 0.001399572, 0.00647301, 
    0.02047836, 4.896148e-05, 0.0004886089, 0.02435666, 0.05689189, 
    0.06398429, 0.03662556, 0.0006374072, 0.01943646, 2.077098e-05, 
    -1.878182e-07, -4.361272e-08, 5.296978e-09, 3.389553e-07, 0.007905769, 
    0.02098276, -0.0002191425, 1.120525e-08, 1.355728e-08,
  3.033022e-07, 9.42456e-05, 2.097125e-06, 0.006869293, 0.01785046, 
    0.008015627, 0.06109859, 0.07667316, 0.02482, 0.01753883, 0.005581157, 
    0.00825001, 0.07529622, 0.07322858, 0.02061396, 0.02914236, 0.001805941, 
    -8.141891e-06, 1.85101e-09, 1.198015e-08, 5.089535e-09, 5.754672e-08, 
    2.873876e-06, 0.00208112, 0.003651671, 0.0001250035, 2.9516e-08, 
    1.208173e-08, 1.392324e-08,
  0.01947268, 0.04339114, 0.06508327, 0.02495971, 0.006045854, 0.05274954, 
    0.01313281, 0.01369936, 0.05753834, 0.2022882, 0.03454974, 0.1251957, 
    0.2383159, 0.05832884, 0.0191114, 0.007920328, 0.003704686, 0.007760673, 
    0.005354194, 0.01201015, 0.007099148, 0.001643389, 0.03390561, 
    0.01797016, 0.01888286, 0.01212409, 0.0119262, 0.002908961, 0.006773296,
  0.1846144, 0.1800579, 0.1576782, 0.1823379, 0.05312619, 0.0199765, 
    0.05284068, 0.008012432, 0.07083973, 0.0210645, 0.01740324, 0.02748021, 
    0.118421, 0.0440019, 0.05472521, 0.09116992, 0.0839862, 0.1193563, 
    0.2103016, 0.1951492, 0.1353537, 0.1147389, 0.1598243, 0.04839382, 
    0.01996891, 0.03203645, 0.06699826, 0.181808, 0.3012512,
  0.004099428, 0.005091693, 0.01622521, 0.08748959, 0.08094093, 0.1254732, 
    0.2534974, 0.0517181, 0.2326313, 0.05324218, 0.1607006, 0.1352211, 
    0.06316326, 0.06956112, 0.02092409, 0.02120578, 1.367683e-05, 
    4.405055e-05, 0.008697726, 0.009931361, 0.0482645, 0.05614086, 
    0.01207422, 0.01013556, 0.006820585, 0.001028983, 0.001281371, 
    0.002907308, 0.006980738,
  0.001224844, 0.005637135, -6.416167e-07, 0.04271426, 0.01674706, 
    0.00137076, 0.05803761, 0.1872096, 0.2087263, 0.06312443, 0.08363244, 
    0.061535, 0.1192339, 0.07168479, 0.120782, 0.01828424, 0.0259017, 
    0.006180637, 3.945314e-05, 0.02791149, 0.03279557, 0.01609467, 
    0.04776909, 0.02405648, 0.01520838, 0.002749479, 0.0003961182, 
    -1.20992e-07, 0.03566992,
  0.01220332, 0.007362043, 0.01552633, 0.01018897, 0.02692039, 0.002958818, 
    0.07971587, 0.05268851, 0.07954331, 0.09103697, 0.1595804, 0.07894136, 
    0.07256915, 0.08625949, 0.1569948, 0.1443965, 0.1035148, 0.06867857, 
    0.01192179, 0.000548267, 0.1197422, 0.06836003, 0.03566033, 0.03480516, 
    0.06518182, 0.03774937, 0.04487419, 0.03033904, 0.005370024,
  0.08563171, 0.1239477, 0.1140896, 0.06374932, 0.05888937, 0.08109657, 
    0.04148189, 0.06830735, 0.1455603, 0.1644301, 0.09565538, 0.07886486, 
    0.09724222, 0.130113, 0.1102984, 0.0788384, 0.1113896, 0.1083157, 
    0.1141023, 0.0246329, 0.05400144, 0.1057857, 0.09875892, 0.08645203, 
    0.09410863, 0.1152163, 0.1336917, 0.1292785, 0.1058865,
  0.1212818, 0.1074452, 0.1192974, 0.1240425, 0.1048738, 0.1442725, 
    0.2040153, 0.1487281, 0.09466438, 0.1148985, 0.1240142, 0.1353878, 
    0.09380854, 0.1651442, 0.1379107, 0.1500677, 0.1738292, 0.2274405, 
    0.3217822, 0.1324556, 0.1047846, 0.1292263, 0.1406508, 0.1410019, 
    0.201347, 0.2778498, 0.1696656, 0.2222129, 0.1683411,
  0.1254159, 0.195494, 0.2209167, 0.1600183, 0.2079584, 0.1384717, 0.1805935, 
    0.2322534, 0.1640864, 0.146784, 0.1511181, 0.1839926, 0.1978512, 
    0.2007845, 0.2369222, 0.1170643, 0.1776736, 0.1842692, 0.1490612, 
    0.2092996, 0.2051111, 0.1620983, 0.1428656, 0.1445107, 0.148239, 
    0.2729352, 0.1781134, 0.2302188, 0.1492838,
  0.1671271, 0.2166768, 0.1376323, 0.1467904, 0.1701745, 0.1708598, 
    0.1176916, 0.1283042, 0.1373, 0.1378494, 0.1748573, 0.1460142, 0.1777801, 
    0.2755288, 0.2944945, 0.2798797, 0.2551792, 0.2663839, 0.2931084, 
    0.2619691, 0.2205386, 0.2815065, 0.1736454, 0.101667, 0.1655765, 
    0.1162014, 0.1093948, 0.1021612, 0.1398428,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.000119819, -0.000119819, 
    -0.000119819, -0.000119819, -0.000119819, -0.000119819, -0.000119819, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0.001432168, -2.705993e-05, 0.0003082, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.063804e-05, 0.007702447, 0.1504241, 0.1344234, 0.1169741, 0.129958, 
    0.1186536, 0.09147026, 0.1139159, 0.04437303, 0.01615797, 0.08950764, 
    0.2242964, 0.1910312, 0.147202, 0.1640046, 0.08248062, 0.002724848,
  0.2637108, 0.2826845, 0.2161895, 0.1406557, 0.01198417, 0.007019589, 
    0.1249942, 0.001670685, 0.004058809, 0.01119353, 0.02151635, 0.05650794, 
    0.2632719, 0.2836009, 0.2646526, 0.2608331, 0.2506551, 0.1957589, 
    0.2059395, 0.2538617, 0.2735141, 0.3143199, 0.3337592, 0.317602, 
    0.2709558, 0.1887186, 0.1812619, 0.1830089, 0.1934853,
  0.2461308, 0.2596047, 0.2543988, 0.2702027, 0.2651345, 0.2464351, 
    0.2475315, 0.2499532, 0.2077745, 0.2688213, 0.3235128, 0.3074528, 
    0.2927234, 0.2712122, 0.2317598, 0.2107771, 0.2346859, 0.2144991, 
    0.1777704, 0.1901567, 0.1858625, 0.2020637, 0.2590124, 0.2243054, 
    0.2700321, 0.2379054, 0.2023407, 0.2410903, 0.2675593,
  0.1785128, 0.1696368, 0.214416, 0.216348, 0.1982447, 0.1615736, 0.1574667, 
    0.196635, 0.1920063, 0.2117638, 0.2259206, 0.2233434, 0.1866588, 
    0.1433238, 0.2018536, 0.1665163, 0.1311617, 0.139031, 0.1866503, 
    0.133385, 0.188526, 0.1653378, 0.2066097, 0.2066219, 0.1568877, 
    0.1746032, 0.1559781, 0.1592469, 0.1644374,
  0.1430475, 0.09540077, 0.06649323, 0.1244373, 0.06940241, 0.08260268, 
    0.102694, 0.07836305, 0.07114801, 0.05757517, 0.07428968, 0.09784701, 
    0.0844284, 0.1058867, 0.1380404, 0.1537925, 0.08901294, 0.1366801, 
    0.1162434, 0.1374009, 0.1716876, 0.1772769, 0.1636041, 0.1408488, 
    0.08500292, 0.07881276, 0.08184886, 0.1297294, 0.1406274,
  0.002499806, 0.0001773154, 0.02631313, 0.01155114, 0.03744414, 0.07231945, 
    0.007478782, 0.002590176, 1.882225e-05, 0.003830166, 0.006121602, 
    0.02789108, 0.03708138, 0.03195125, 0.06224415, 0.0851364, 0.1506923, 
    0.2046826, 0.1096741, 0.04613596, 0.03987043, 0.01500802, 0.0006842988, 
    0.006468352, 0.06539203, 0.09720513, 0.06554748, 0.02303611, 0.01531723,
  3.454319e-07, 3.230625e-07, 3.451102e-05, 0.001221915, 0.01770556, 
    0.0123839, -8.540865e-06, 0.007390562, 0.0008487931, 0.01201774, 
    0.02805673, 8.345971e-06, 0.0004680299, 0.03151048, 0.05335859, 
    0.07736488, 0.04093335, 0.001136183, 0.02532293, 5.742053e-06, 
    -6.556048e-06, -5.198299e-07, 1.018398e-08, 5.276485e-07, 0.01134064, 
    0.0222264, 0.0005120079, 1.04371e-07, 1.773235e-07,
  7.440393e-07, 0.001047601, 4.598685e-05, 0.00826089, 0.02197077, 
    0.01398375, 0.06094752, 0.07515317, 0.02999331, 0.02078914, 0.01117022, 
    0.01372331, 0.08337466, 0.08141919, 0.02802206, 0.03631026, 0.006747419, 
    0.0002608543, 8.280374e-08, 4.85113e-08, 9.469534e-08, 3.421813e-07, 
    6.426038e-06, 0.003064502, 0.002143672, 0.0003137541, 2.05539e-07, 
    4.707977e-08, 8.071012e-08,
  0.01480123, 0.04683298, 0.1072246, 0.02730804, 0.003384016, 0.05869784, 
    0.01549627, 0.02146294, 0.06936999, 0.2359006, 0.0512295, 0.1393389, 
    0.2444044, 0.0682646, 0.01970994, 0.008791054, 0.006850306, 0.00717902, 
    0.005499185, 0.001638916, 0.002106533, 0.002729712, 0.03762534, 
    0.02164041, 0.01929737, 0.01998265, 0.03197892, 0.0008667685, 0.003780143,
  0.1955028, 0.2170011, 0.1908893, 0.2288238, 0.07629935, 0.01876771, 
    0.06179894, 0.02232127, 0.1106605, 0.03792136, 0.02928182, 0.04146037, 
    0.1320128, 0.05476244, 0.07326745, 0.1173888, 0.1034542, 0.1640401, 
    0.2479843, 0.2493366, 0.1466182, 0.1424244, 0.173184, 0.06979431, 
    0.02618366, 0.04526479, 0.08928239, 0.2295163, 0.3424764,
  0.04351998, 0.001621477, 0.01118186, 0.07650658, 0.07129518, 0.1365053, 
    0.2926199, 0.08618437, 0.2761814, 0.06993853, 0.1960968, 0.1582573, 
    0.07768381, 0.08522069, 0.02827338, 0.02302743, 0.0007098907, 
    0.002289562, 0.008572373, 0.02136357, 0.06530615, 0.06687745, 0.01622205, 
    0.01541341, 0.009441413, 0.00424507, 0.001455861, 0.003372011, 0.007498301,
  -5.939843e-05, 0.02504417, 1.300116e-08, 0.02075204, 0.01309443, 
    0.002745501, 0.06886841, 0.1994928, 0.2423205, 0.07829189, 0.09839524, 
    0.082581, 0.1341045, 0.08618227, 0.1292116, 0.01654745, 0.01818563, 
    0.002326184, 7.423123e-06, 0.008904609, 0.05463159, 0.02161559, 
    0.0545052, 0.0248002, 0.01970871, 0.003074316, 0.0004762974, 
    6.601437e-08, 0.02443255,
  0.008278504, 0.003941812, 0.01509133, 0.01573133, 0.01602175, 0.004209322, 
    0.09196918, 0.04802906, 0.06200205, 0.08869766, 0.1542714, 0.07239682, 
    0.07980339, 0.08864483, 0.1611441, 0.142134, 0.09706894, 0.06075965, 
    0.01526216, 0.0003233713, 0.08016565, 0.06416856, 0.03892307, 0.043556, 
    0.06760534, 0.03805014, 0.04626396, 0.02801132, 0.002823486,
  0.07846696, 0.1144142, 0.1088125, 0.07068671, 0.05707708, 0.07481691, 
    0.04158618, 0.07225315, 0.1422469, 0.1783777, 0.0953957, 0.08466858, 
    0.1027089, 0.134178, 0.09995791, 0.07728184, 0.1199423, 0.1108023, 
    0.1164097, 0.0232478, 0.06302794, 0.08828569, 0.1004237, 0.09817559, 
    0.101238, 0.1121195, 0.1342607, 0.1222202, 0.1025241,
  0.1283089, 0.1016779, 0.1140129, 0.09915952, 0.106292, 0.1567039, 
    0.1979052, 0.1575243, 0.1033244, 0.1182607, 0.1143475, 0.1405487, 
    0.1073353, 0.1820939, 0.1209442, 0.1499827, 0.1665778, 0.2163366, 
    0.3482395, 0.1258748, 0.109181, 0.1329779, 0.1594385, 0.1634033, 
    0.2017645, 0.2837901, 0.1530271, 0.1974073, 0.1766476,
  0.1256154, 0.1582389, 0.2318584, 0.118973, 0.225358, 0.1761993, 0.1989144, 
    0.269015, 0.161435, 0.1619556, 0.1659048, 0.1962756, 0.1758363, 
    0.2046104, 0.2246379, 0.1187821, 0.200622, 0.1958671, 0.1643728, 
    0.2491591, 0.2232006, 0.1952411, 0.1496052, 0.1508588, 0.1253295, 
    0.2802583, 0.1801061, 0.2049312, 0.1479538,
  0.1586336, 0.190086, 0.1348083, 0.1433127, 0.1468464, 0.1671288, 0.131861, 
    0.1319885, 0.1495553, 0.1653879, 0.1856681, 0.169757, 0.2369166, 
    0.3354105, 0.3815629, 0.3425662, 0.3067321, 0.2829304, 0.3177267, 
    0.2765037, 0.2060386, 0.2789348, 0.1901415, 0.1158914, 0.1753236, 
    0.1352266, 0.136446, 0.1040077, 0.1210045,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.412013e-05, -9.412013e-05, 
    -9.412013e-05, -9.412013e-05, -9.412013e-05, -9.412013e-05, 
    -9.412013e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0.004290987, 0.002368123, 0.004686478, 0.001724849, -1.391719e-05, 
    -1.851805e-07, 0, 0, 0, 0, -0.0001562552, 0.009775683, 0.02144496, 
    0.1804214, 0.1326332, 0.1275388, 0.1485269, 0.1660641, 0.1362134, 
    0.161138, 0.1137933, 0.09660627, 0.1574296, 0.2207689, 0.1854029, 
    0.1670909, 0.1750757, 0.1821157, 0.008999678,
  0.2795089, 0.288817, 0.236144, 0.1646553, 0.01879881, 0.01730827, 
    0.1349159, 0.03059185, 0.02414412, 0.06713082, 0.08631521, 0.1753085, 
    0.3029793, 0.2856231, 0.2618202, 0.2783862, 0.2453365, 0.206691, 
    0.2243961, 0.2624839, 0.2791789, 0.3196456, 0.339069, 0.313426, 
    0.2612345, 0.1850101, 0.1676401, 0.1825988, 0.204479,
  0.2485441, 0.2499255, 0.235145, 0.2709728, 0.2577828, 0.24452, 0.2351639, 
    0.2500021, 0.2075492, 0.2881811, 0.3225003, 0.2804002, 0.282609, 0.2696, 
    0.2356355, 0.2012013, 0.2226895, 0.2240458, 0.1781266, 0.2130741, 
    0.1996705, 0.2047367, 0.2733554, 0.2132744, 0.271041, 0.2264097, 
    0.1970313, 0.234843, 0.258427,
  0.182498, 0.1676066, 0.1934129, 0.2072576, 0.2082188, 0.1755225, 0.1583095, 
    0.2043311, 0.183529, 0.1995665, 0.2338238, 0.2275817, 0.1994134, 
    0.1563174, 0.1903206, 0.1711158, 0.1313707, 0.1379809, 0.1717869, 
    0.1331289, 0.1835724, 0.171048, 0.1928423, 0.1982575, 0.1494761, 
    0.1619445, 0.1498832, 0.1581923, 0.1569327,
  0.1289099, 0.09700911, 0.07240465, 0.1167084, 0.0692991, 0.08736119, 
    0.1067088, 0.0818945, 0.07364552, 0.06856903, 0.08296504, 0.1060587, 
    0.084181, 0.1035557, 0.1332105, 0.1375354, 0.08820772, 0.1439006, 
    0.1157215, 0.1358076, 0.1615672, 0.1592062, 0.1474747, 0.1411676, 
    0.0792862, 0.07236398, 0.07647645, 0.137268, 0.1493885,
  0.002560718, 0.0005055397, 0.06335402, 0.02025506, 0.03997242, 0.09087363, 
    0.008768192, 0.003266694, 0.0007252641, 0.01564026, 0.02188497, 
    0.0420101, 0.05082886, 0.03572232, 0.07099259, 0.09273627, 0.1536719, 
    0.1885455, 0.1000037, 0.05021403, 0.05245274, 0.02438383, 0.001044705, 
    0.00635739, 0.08415819, 0.1036693, 0.06682017, 0.03363844, 0.01855315,
  3.654035e-07, 5.810731e-05, 0.005447558, 0.001054389, 0.03513524, 
    0.01447365, 0.00586543, 0.0003201757, 0.0004656803, 0.01256813, 
    0.03447808, 0.0001930568, 0.0001456687, 0.03342322, 0.05084752, 
    0.09080116, 0.04513259, 0.001259927, 0.03826167, 5.586318e-05, 
    -4.195696e-05, -1.0859e-06, 9.416825e-09, 3.75281e-07, 0.02167253, 
    0.02517822, 0.00195982, 4.905071e-07, 1.474992e-07,
  9.850221e-07, 0.003080966, 0.002193437, 0.007217445, 0.02403687, 
    0.02060898, 0.0688405, 0.08385134, 0.041575, 0.01985059, 0.01332765, 
    0.01192637, 0.09803598, 0.09838862, 0.03886183, 0.03998074, 0.01049022, 
    0.0004639876, 2.592123e-05, 5.767081e-08, 1.668676e-07, 4.000392e-07, 
    8.931822e-06, 0.006406605, 0.007192138, 0.002670142, 1.421634e-07, 
    5.375934e-08, 9.803217e-08,
  0.01299996, 0.06009491, 0.16583, 0.02394782, 0.008255994, 0.06975938, 
    0.01826236, 0.03258629, 0.1016832, 0.2794727, 0.06193518, 0.1574121, 
    0.2491253, 0.08086672, 0.02058836, 0.009923194, 0.007396218, 0.006970818, 
    0.002930071, 0.0002631826, 0.00376612, 0.0004818079, 0.03626016, 
    0.0409531, 0.03082512, 0.0231259, 0.0310387, 0.006199307, 0.008613787,
  0.2406838, 0.2733089, 0.2310183, 0.2884386, 0.09275851, 0.01489078, 
    0.06948706, 0.04543288, 0.1384932, 0.0423165, 0.04319202, 0.05498068, 
    0.1476266, 0.07025156, 0.09157614, 0.1388611, 0.119026, 0.19481, 
    0.2708402, 0.3096859, 0.1489395, 0.1612529, 0.190612, 0.09620094, 
    0.03008625, 0.0554587, 0.1073927, 0.2459897, 0.3717998,
  0.03985071, 0.003950653, 0.003325718, 0.05459358, 0.05551116, 0.09488763, 
    0.3527172, 0.09167092, 0.3251171, 0.0718313, 0.1855976, 0.154335, 
    0.0795275, 0.09773942, 0.03801687, 0.02536439, 0.0005519209, 
    0.0003377263, 0.003354297, 0.01707701, 0.08741681, 0.0787824, 0.01705742, 
    0.01713958, 0.01001394, 0.002258351, 0.0003432906, 0.001150873, 
    0.003173099,
  -7.533595e-06, 0.01166807, 6.643732e-08, 0.007867665, 0.0069121, 
    0.003334154, 0.06481465, 0.2126047, 0.254592, 0.07413451, 0.1019146, 
    0.08352838, 0.1479224, 0.09598957, 0.1423242, 0.0147761, 0.01702608, 
    0.006748377, 0.002636867, 0.0005786379, 0.06412412, 0.02632139, 
    0.06168728, 0.03324244, 0.02196646, 0.004659191, 0.001224905, 
    7.046222e-08, 0.008249029,
  0.002705822, 0.003322588, 0.01521322, 0.01740187, 0.01274539, 0.005980926, 
    0.08357296, 0.04617368, 0.04837178, 0.1030746, 0.1563657, 0.07651076, 
    0.08693583, 0.09570169, 0.1703772, 0.1466621, 0.09244613, 0.05988947, 
    0.01348231, 0.0007068783, 0.03646126, 0.04599079, 0.04782759, 0.0583777, 
    0.08346428, 0.04251884, 0.05720551, 0.02896078, 0.001398678,
  0.07450821, 0.1196858, 0.1106664, 0.06927945, 0.0641958, 0.07624325, 
    0.05213274, 0.07563224, 0.1423036, 0.1712036, 0.1059567, 0.09667802, 
    0.1051336, 0.1479607, 0.09282735, 0.07778105, 0.1267826, 0.1206018, 
    0.127864, 0.02036634, 0.06424787, 0.06886458, 0.1047829, 0.1028361, 
    0.116286, 0.1249334, 0.1323982, 0.1303323, 0.1086602,
  0.1141948, 0.09873645, 0.09702997, 0.09026487, 0.1042155, 0.1755177, 
    0.2090963, 0.1420788, 0.09974311, 0.1262685, 0.1190829, 0.1596941, 
    0.1191548, 0.200533, 0.1395959, 0.1529507, 0.1556488, 0.2290355, 
    0.3586532, 0.1232286, 0.1096326, 0.1414801, 0.1759533, 0.1737324, 
    0.2123061, 0.3002777, 0.168945, 0.1780683, 0.1648053,
  0.1119294, 0.1462303, 0.2215967, 0.1505647, 0.2464816, 0.1692576, 
    0.2119983, 0.2636816, 0.2353574, 0.171328, 0.1764003, 0.2057619, 
    0.1894393, 0.2046767, 0.2319608, 0.1232414, 0.2052181, 0.2036738, 
    0.1599811, 0.2553811, 0.2229293, 0.1925884, 0.1299167, 0.1389899, 
    0.1039455, 0.3159978, 0.18626, 0.2081478, 0.1320595,
  0.166194, 0.2168273, 0.1422911, 0.1245811, 0.1583177, 0.1659445, 0.1685059, 
    0.1656138, 0.1893815, 0.1897963, 0.2283669, 0.2310403, 0.2553645, 
    0.3795694, 0.4062472, 0.3342283, 0.3144949, 0.309669, 0.3350005, 
    0.269315, 0.2031358, 0.2715428, 0.1873, 0.1202152, 0.1586801, 0.1719657, 
    0.1520615, 0.115589, 0.1366315,
  0.000182111, 5.738459e-05, -6.734183e-05, -0.0001920682, -0.0003167946, 
    -0.0004415211, -0.0005662475, -5.834131e-05, -4.202552e-05, 
    -2.570974e-05, -9.393963e-06, 6.921817e-06, 2.32376e-05, 3.955338e-05, 
    -0.001355608, -0.001089019, -0.0008224298, -0.0005558408, -0.0002892518, 
    -2.266276e-05, 0.0002439263, -0.0003395235, -0.0004977019, -0.0006558803, 
    -0.0008140586, -0.000972237, -0.001130415, -0.001288594, 0.0002818921,
  0.003284797, 0.01100269, 0.01899751, 0.006940732, -0.0003074774, 
    1.087629e-06, 5.243484e-07, 0, 0, 0, 0.001776835, 0.01941988, 0.02524109, 
    0.184343, 0.1237057, 0.1273303, 0.1688494, 0.1908592, 0.199616, 
    0.2244426, 0.1974209, 0.1525175, 0.1892286, 0.2314003, 0.1693403, 
    0.157817, 0.1598497, 0.2179061, 0.04431425,
  0.2863667, 0.3014667, 0.2451231, 0.1765083, 0.0377835, 0.06135879, 
    0.1411218, 0.08127666, 0.06326856, 0.1313403, 0.1472262, 0.2144334, 
    0.3122729, 0.3010107, 0.2954096, 0.2985184, 0.2671543, 0.2399984, 
    0.222927, 0.2930628, 0.2702885, 0.3254847, 0.3450959, 0.3390974, 
    0.2699162, 0.1725005, 0.1688231, 0.1952198, 0.2161847,
  0.255215, 0.2420032, 0.2427889, 0.2781036, 0.249804, 0.232968, 0.2441875, 
    0.2722185, 0.217964, 0.2971063, 0.3205201, 0.2721882, 0.2899323, 
    0.2665756, 0.2496893, 0.2036349, 0.2217399, 0.2291892, 0.1943781, 
    0.2246362, 0.2072932, 0.2215744, 0.2657824, 0.2230555, 0.2748967, 
    0.2229982, 0.1884302, 0.2227974, 0.2711249,
  0.1851512, 0.1703193, 0.1961112, 0.203182, 0.1966321, 0.1792425, 0.1662891, 
    0.2129569, 0.1833143, 0.219782, 0.2573839, 0.2379892, 0.2054046, 
    0.1629053, 0.1909917, 0.1714942, 0.1321641, 0.14123, 0.1674877, 
    0.1519078, 0.1866257, 0.1627726, 0.1825131, 0.1961409, 0.1383952, 
    0.1566162, 0.1501936, 0.1621874, 0.1559506,
  0.1296898, 0.105888, 0.08189966, 0.1102449, 0.0735205, 0.08074791, 
    0.1020886, 0.08757411, 0.07470806, 0.07733472, 0.09036027, 0.114036, 
    0.08724442, 0.1077373, 0.1334287, 0.1405633, 0.09450488, 0.1455713, 
    0.1090122, 0.1299126, 0.1528466, 0.1578246, 0.1410401, 0.1417737, 
    0.07975309, 0.06316248, 0.07275395, 0.1377925, 0.157585,
  0.004601878, 0.000589977, 0.07832053, 0.01944556, 0.04586257, 0.09553104, 
    0.01325219, 0.003886679, 0.001744397, 0.01233613, 0.03197676, 0.0365024, 
    0.06617747, 0.04166566, 0.07232878, 0.1067397, 0.156663, 0.1768704, 
    0.1010758, 0.06141502, 0.05528783, 0.03340982, 0.001543704, 0.006241491, 
    0.1077034, 0.1102117, 0.06905178, 0.03681581, 0.02478483,
  1.292277e-07, 4.278101e-07, 0.001382427, 0.001728142, 0.04186055, 
    0.01503816, 0.01107796, 0.0003195036, -0.0001444537, 0.005635826, 
    0.04483251, 0.004310696, 0.006478033, 0.03448287, 0.04247952, 0.09034363, 
    0.05321991, 0.002848893, 0.04525315, 0.001890046, -5.860454e-05, 
    -2.934187e-06, 4.821916e-09, 1.885033e-07, 0.01918838, 0.02977908, 
    0.003279108, 4.000556e-07, 1.217621e-07,
  3.202828e-06, 0.0001914767, 0.01372272, 0.003081465, 0.02491687, 
    0.02009643, 0.08295007, 0.07728033, 0.04230469, 0.01820003, 0.01299609, 
    0.009047434, 0.1029976, 0.09799781, 0.04215297, 0.04463343, 0.01276343, 
    0.001116662, 6.798233e-05, 5.263732e-08, 1.901706e-07, 3.515109e-07, 
    9.450911e-06, 0.01031939, 0.03864225, 0.01465617, 4.449029e-05, 
    1.12859e-07, 1.184655e-07,
  0.01611808, 0.07724151, 0.1961927, 0.02615405, 0.002154165, 0.06627867, 
    0.0199587, 0.03068416, 0.112402, 0.3092461, 0.04228026, 0.1154389, 
    0.2250525, 0.07108335, 0.02184937, 0.01009425, 0.01075435, 0.00754645, 
    0.006817858, 0.008687308, 0.00529151, 0.001918023, 0.03038216, 
    0.06925013, 0.03829855, 0.01794765, 0.01404936, 0.004940504, 0.01210055,
  0.2394052, 0.293245, 0.2429482, 0.343123, 0.06890754, 0.02604982, 
    0.06871305, 0.04248447, 0.07851478, 0.03881913, 0.02840648, 0.03336334, 
    0.1102652, 0.0574396, 0.07754917, 0.1349284, 0.1304186, 0.2155696, 
    0.2702782, 0.3126528, 0.1206359, 0.1378793, 0.20188, 0.1023654, 
    0.02726708, 0.052898, 0.09626888, 0.207321, 0.4058967,
  0.01176956, 0.006593659, 0.0001621235, 0.02570896, 0.02958916, 0.0494, 
    0.2632438, 0.08383863, 0.3463473, 0.06193088, 0.1366524, 0.1080511, 
    0.05269634, 0.06983999, 0.02758992, 0.02375884, 0.0004413842, 
    1.628242e-05, 0.001694034, 0.01027398, 0.06570157, 0.08215272, 
    0.01392843, 0.01346398, 0.009434487, 0.001441759, 0.0001101184, 
    0.000642499, 0.002449466,
  1.963389e-06, 0.002826883, 2.335874e-09, 0.002102937, 0.003064672, 
    0.002217408, 0.06147126, 0.2621414, 0.2754975, 0.05517595, 0.08550353, 
    0.06818816, 0.1244442, 0.07923819, 0.1265001, 0.01405681, 0.01437411, 
    0.003751249, 0.000660888, 2.093051e-05, 0.06496003, 0.02400238, 
    0.05438264, 0.03139867, 0.01510597, 0.005709673, 0.0009849726, 
    2.749427e-08, 0.0006383012,
  0.001178912, 0.002544553, 0.01888896, 0.01735152, 0.007292284, 0.006315029, 
    0.06211246, 0.03408854, 0.03461265, 0.1092181, 0.1629999, 0.0708975, 
    0.09470046, 0.095654, 0.1877438, 0.1768152, 0.1022599, 0.08064934, 
    0.01717986, 0.0003275722, 0.01591512, 0.02885297, 0.04840326, 0.06304812, 
    0.08880998, 0.04852942, 0.06688988, 0.03046153, 0.001838227,
  0.07538739, 0.1215297, 0.1246316, 0.1041379, 0.0723317, 0.06863252, 
    0.06491945, 0.07586718, 0.1391141, 0.1648224, 0.123193, 0.1046481, 
    0.1192887, 0.1693084, 0.1000118, 0.0843861, 0.1533228, 0.1208444, 
    0.1366584, 0.03005344, 0.07175022, 0.05252929, 0.1003771, 0.1205479, 
    0.13044, 0.1428787, 0.1370102, 0.140417, 0.1492134,
  0.1152198, 0.1124532, 0.1014565, 0.1028843, 0.1034385, 0.1918447, 
    0.2010732, 0.143495, 0.10841, 0.1361742, 0.1255169, 0.1788028, 0.1326873, 
    0.2241562, 0.1419431, 0.1576427, 0.1529028, 0.2841389, 0.3825078, 
    0.130877, 0.1139527, 0.1656739, 0.2068803, 0.1747736, 0.241389, 
    0.3107474, 0.1831504, 0.1705887, 0.1594215,
  0.1054731, 0.1601275, 0.247499, 0.1340658, 0.1875923, 0.15754, 0.1926488, 
    0.2765388, 0.2016657, 0.1887318, 0.1894424, 0.2261221, 0.235072, 
    0.2351851, 0.2532644, 0.1591415, 0.2053126, 0.1890362, 0.164446, 
    0.2549669, 0.2263802, 0.1885388, 0.1331899, 0.1781238, 0.09903312, 
    0.3455822, 0.2115977, 0.189222, 0.144325,
  0.1673836, 0.1818065, 0.1417841, 0.1080287, 0.1288981, 0.1842226, 
    0.1544239, 0.1653518, 0.179671, 0.2313954, 0.262557, 0.2571791, 
    0.2861346, 0.3907936, 0.376195, 0.3311194, 0.2970233, 0.2677022, 
    0.2979096, 0.2673986, 0.1954494, 0.2812456, 0.2152195, 0.1432404, 
    0.1702601, 0.1785052, 0.1587521, 0.1232458, 0.1367531,
  0.01049956, 0.009294025, 0.008088488, 0.006882951, 0.005677413, 
    0.004471876, 0.003266339, 0.002917122, 0.002986768, 0.003056414, 
    0.00312606, 0.003195706, 0.003265352, 0.003334997, 0.003971966, 
    0.005796439, 0.007620911, 0.009445383, 0.01126985, 0.01309433, 0.0149188, 
    0.01441591, 0.01372733, 0.01303875, 0.01235017, 0.01166159, 0.010973, 
    0.01028442, 0.01146399,
  0.0255123, 0.01688533, 0.03235952, 0.02635251, 0.001984937, 0.0001793288, 
    0.0004559533, 0, 0, 2.644692e-05, 0.01263774, 0.02359732, 0.03632148, 
    0.1695189, 0.1033699, 0.1527133, 0.2025202, 0.2111405, 0.2397762, 
    0.2716205, 0.2549937, 0.2376015, 0.204483, 0.2222475, 0.1611048, 
    0.148723, 0.1633382, 0.2101464, 0.1145331,
  0.2815211, 0.2995844, 0.2586238, 0.1808058, 0.07475406, 0.1295093, 
    0.1567261, 0.1227877, 0.1114131, 0.2134741, 0.1989004, 0.2607631, 
    0.3208975, 0.323123, 0.3124122, 0.3383759, 0.3069243, 0.2813966, 
    0.2728807, 0.3073403, 0.299405, 0.3296066, 0.3774669, 0.3717095, 
    0.2888017, 0.1799799, 0.1922368, 0.1844457, 0.2303885,
  0.2856798, 0.2717665, 0.2705649, 0.2985785, 0.2713451, 0.2381196, 
    0.2595766, 0.3061353, 0.2733315, 0.3011773, 0.3446295, 0.2700801, 
    0.2833477, 0.2762191, 0.2631944, 0.2267554, 0.2497664, 0.2638114, 
    0.2310475, 0.2377085, 0.2377518, 0.2643341, 0.2778674, 0.2292559, 
    0.26539, 0.207544, 0.1973063, 0.2329238, 0.2811573,
  0.2106279, 0.1818934, 0.2055678, 0.2017642, 0.1907794, 0.1918203, 
    0.1824192, 0.2393124, 0.2062801, 0.2270218, 0.2631418, 0.2585993, 
    0.2193488, 0.1850132, 0.2013767, 0.1794008, 0.128175, 0.1805307, 
    0.2007732, 0.1891491, 0.2114766, 0.1807358, 0.1909882, 0.1926897, 
    0.1395264, 0.1504488, 0.1546168, 0.1812195, 0.1576159,
  0.1442801, 0.1396, 0.09096283, 0.1019145, 0.08697487, 0.09121075, 
    0.1055647, 0.08803916, 0.08150388, 0.09892523, 0.09761767, 0.1173335, 
    0.08991807, 0.107279, 0.1321241, 0.1442601, 0.09826152, 0.148151, 
    0.1070655, 0.1275987, 0.1539259, 0.1729089, 0.1366518, 0.1423202, 
    0.06486746, 0.05782909, 0.08043844, 0.1418798, 0.1722348,
  0.008650023, 0.0008056573, 0.06524801, 0.02054632, 0.05961661, 0.09934851, 
    0.01683722, 0.008503936, 0.004398989, 0.01464093, 0.02583018, 0.02278686, 
    0.06717025, 0.04694042, 0.07690876, 0.1217656, 0.1654578, 0.165859, 
    0.1026615, 0.07336269, 0.07612298, 0.03969339, 0.003368238, 0.006942962, 
    0.1138294, 0.1083705, 0.07374383, 0.04571381, 0.02837907,
  6.404964e-08, -3.053447e-05, 0.004672214, 0.005788706, 0.046028, 
    0.02392998, 0.01089418, 0.003873874, 0.0004443362, 0.001347973, 
    0.03104804, 0.01901524, 0.01887939, 0.04497794, 0.07068501, 0.08329859, 
    0.0793848, 0.01011815, 0.04347354, 0.01483651, 5.51265e-05, 
    -4.229241e-05, 5.078352e-09, 2.166496e-07, 0.02093341, 0.03162182, 
    0.008408044, 5.539397e-07, 5.377716e-06,
  -1.365756e-07, -0.0001588801, 0.02030521, 0.02293919, 0.0232849, 
    0.02287006, 0.06616452, 0.07432042, 0.03930524, 0.00842139, 0.01352147, 
    0.00621099, 0.1097335, 0.1010405, 0.03934618, 0.04892887, 0.01662683, 
    0.002098992, 0.0006501405, 5.595437e-08, 2.006295e-07, 2.645656e-07, 
    4.615101e-06, 0.01162704, 0.08095138, 0.02351161, 0.00428109, 
    8.656381e-06, 1.107257e-07,
  0.004493368, 0.07010422, 0.1624592, 0.01903192, 0.0008527923, 0.05920408, 
    0.01721203, 0.03168208, 0.08135357, 0.256988, 0.03625347, 0.08181822, 
    0.2009371, 0.06358667, 0.02319655, 0.009042194, 0.007287886, 0.003313535, 
    0.01007249, 0.006199365, 0.0004034067, 0.00335116, 0.02957108, 
    0.07357574, 0.03565717, 0.01482448, 0.006562209, 0.006462593, 0.004471392,
  0.1263199, 0.1840599, 0.1571842, 0.4318432, 0.06389265, 0.02074272, 
    0.07447585, 0.04101556, 0.04883612, 0.03374293, 0.02123011, 0.02162897, 
    0.08649167, 0.04820417, 0.06870357, 0.1287809, 0.1349871, 0.211185, 
    0.2578774, 0.3062762, 0.09995414, 0.1252917, 0.1814935, 0.09867181, 
    0.02727873, 0.04869575, 0.09319907, 0.1737577, 0.326041,
  0.002000682, 0.004119924, -4.040329e-05, 0.0253371, 0.02000618, 0.03190625, 
    0.2155994, 0.08645177, 0.3180504, 0.05861184, 0.1176017, 0.08077753, 
    0.04106595, 0.05183487, 0.02083181, 0.01626855, 0.0001370146, 
    2.705877e-07, 0.001527017, 0.006951686, 0.04950698, 0.08518146, 
    0.01202502, 0.01004512, 0.00844148, 0.001436549, 3.571378e-05, 
    3.188304e-05, 0.001232439,
  1.612472e-06, 0.00359091, 3.612096e-09, 0.0001226229, 0.0006830083, 
    0.001420564, 0.05562945, 0.288632, 0.313272, 0.05315586, 0.07548106, 
    0.06659111, 0.09079199, 0.0552576, 0.09139889, 0.008714902, 0.01472982, 
    0.004131927, 0.0005242582, 1.060405e-05, 0.05723914, 0.0255268, 
    0.0435177, 0.01728048, 0.0121375, 0.00556306, 0.0003905578, 2.648681e-08, 
    7.322981e-05,
  0.001182699, 0.001060159, 0.0153199, 0.02286128, 0.001863325, 0.00696028, 
    0.04926241, 0.02338575, 0.03140975, 0.1156187, 0.1501187, 0.05647583, 
    0.09466064, 0.09775116, 0.1437529, 0.177164, 0.1377364, 0.08417383, 
    0.02242629, 0.0006691227, 0.007961622, 0.009780828, 0.04329468, 
    0.05028049, 0.06621732, 0.04984078, 0.05855848, 0.02950535, 0.001757066,
  0.07774408, 0.139962, 0.1226269, 0.1189926, 0.08194098, 0.05829685, 
    0.06128838, 0.08034751, 0.1528186, 0.1727746, 0.1302413, 0.1111464, 
    0.1010015, 0.1768609, 0.1070151, 0.08890394, 0.1562054, 0.1227696, 
    0.1400901, 0.0396104, 0.07009761, 0.03665855, 0.09412032, 0.1337305, 
    0.1395502, 0.1484336, 0.1511747, 0.1454566, 0.1449844,
  0.1647994, 0.1153445, 0.123339, 0.136894, 0.1170873, 0.2000433, 0.2338237, 
    0.1887121, 0.14501, 0.1531345, 0.1309361, 0.2017163, 0.1554479, 
    0.2636567, 0.1605184, 0.1709638, 0.1741545, 0.3237437, 0.3823294, 
    0.1550874, 0.1156252, 0.1663786, 0.2134936, 0.1808018, 0.2264411, 
    0.3022307, 0.1655857, 0.1730015, 0.164239,
  0.1295479, 0.1656489, 0.2373712, 0.1422945, 0.202538, 0.1385976, 0.2064632, 
    0.279312, 0.1882651, 0.1721207, 0.1830747, 0.2016811, 0.2189706, 
    0.221236, 0.2397209, 0.1745942, 0.2090692, 0.2251229, 0.1493266, 
    0.2817842, 0.2154387, 0.2254427, 0.1560198, 0.1569499, 0.1147044, 
    0.353999, 0.2638599, 0.1999247, 0.1677081,
  0.1441895, 0.1710203, 0.1168803, 0.1334689, 0.1457797, 0.1549993, 
    0.1477778, 0.176005, 0.1770626, 0.2032643, 0.2011701, 0.2671624, 
    0.2954974, 0.3968126, 0.4418556, 0.3309909, 0.3384444, 0.3143404, 
    0.2840416, 0.2301687, 0.1952165, 0.2632824, 0.2261112, 0.1860295, 
    0.1431247, 0.1674738, 0.1543838, 0.1006506, 0.1472713,
  0.02556998, 0.02315734, 0.02074469, 0.01833204, 0.01591939, 0.01350674, 
    0.0110941, 0.0168636, 0.01790016, 0.01893672, 0.01997328, 0.02100984, 
    0.0220464, 0.02308296, 0.01137329, 0.01633821, 0.02130313, 0.02626805, 
    0.03123297, 0.03619789, 0.04116281, 0.05038941, 0.04680058, 0.04321174, 
    0.03962291, 0.03603408, 0.03244524, 0.02885641, 0.0275001,
  0.0802985, 0.01740697, 0.03626468, 0.03751057, 0.004856537, 0.0001722798, 
    0.001266265, -8.176555e-06, 7.298369e-06, 0.004073134, 0.02002039, 
    0.02822093, 0.06312357, 0.142352, 0.08155864, 0.1336103, 0.1992683, 
    0.252601, 0.2657968, 0.2861849, 0.3243453, 0.282614, 0.2041509, 
    0.2329211, 0.1611364, 0.1487048, 0.1634543, 0.2090993, 0.1734794,
  0.2727232, 0.2982784, 0.2852666, 0.1907119, 0.1261796, 0.1816559, 
    0.1809727, 0.1621439, 0.1723537, 0.2860861, 0.2612287, 0.3129315, 
    0.3202933, 0.3233656, 0.3429512, 0.3520136, 0.3064204, 0.2814838, 
    0.3032541, 0.3430521, 0.3220706, 0.3454812, 0.3790498, 0.392499, 
    0.3196752, 0.2075011, 0.2003281, 0.2089862, 0.2443898,
  0.3261234, 0.2618606, 0.2836617, 0.3046922, 0.2947882, 0.261041, 0.2756747, 
    0.3111714, 0.3387805, 0.3297292, 0.3687856, 0.2884389, 0.3284159, 
    0.3290027, 0.3230034, 0.2586037, 0.2756251, 0.2880241, 0.2673445, 
    0.2635815, 0.2705818, 0.2825775, 0.2864379, 0.2486787, 0.2876085, 
    0.2366117, 0.243348, 0.2678872, 0.3222784,
  0.2308928, 0.2211735, 0.2190078, 0.2215567, 0.218217, 0.2081609, 0.2193085, 
    0.2710865, 0.2322029, 0.2513657, 0.2840327, 0.2882121, 0.2320457, 
    0.201414, 0.1867123, 0.1887394, 0.1341982, 0.1933126, 0.1987399, 
    0.2037619, 0.2428294, 0.2116951, 0.2235119, 0.196823, 0.1281886, 
    0.1525075, 0.1709136, 0.2063317, 0.1957797,
  0.1697842, 0.1626366, 0.1000547, 0.1045903, 0.1172511, 0.1028555, 0.123133, 
    0.09717597, 0.09474325, 0.1151184, 0.1043041, 0.1381082, 0.09725207, 
    0.1111741, 0.1395816, 0.1695216, 0.119121, 0.1583451, 0.1148615, 
    0.1354766, 0.1706907, 0.1890844, 0.1437327, 0.1459599, 0.05535702, 
    0.05853292, 0.103403, 0.1609362, 0.1911647,
  0.01640274, 0.001866142, 0.05034737, 0.01831393, 0.06106427, 0.107828, 
    0.02708725, 0.02006623, 0.01081175, 0.01808253, 0.02063349, 0.01801867, 
    0.07359459, 0.05339945, 0.08806591, 0.1373229, 0.1733511, 0.1644083, 
    0.1192193, 0.09129753, 0.08636049, 0.06194039, 0.006934678, 0.007151055, 
    0.1038359, 0.1027074, 0.08024926, 0.05222484, 0.03587674,
  1.049162e-07, -1.71391e-06, 0.01917097, 0.008127267, 0.05339291, 
    0.02439664, 0.020568, 0.02803637, 0.0120636, 0.004246467, 0.008024592, 
    0.01806008, 0.03751709, 0.04034144, 0.08252049, 0.07058443, 0.09755801, 
    0.03357466, 0.04615295, 0.02529178, 0.002508439, -1.321616e-05, 
    2.918e-08, 2.182294e-06, 0.02409809, 0.03670012, 0.01856932, 
    0.0006023785, 0.001165951,
  6.660483e-08, -3.710783e-05, 0.01238327, 0.08639188, 0.02359243, 
    0.02734729, 0.05249236, 0.07500679, 0.03508935, 0.005678817, 0.01638719, 
    0.006325763, 0.1313436, 0.101535, 0.04300902, 0.05508143, 0.02213436, 
    0.003755019, 0.0008558011, 1.919166e-06, 3.332579e-07, 2.014556e-07, 
    1.217156e-06, 0.01228203, 0.02880247, 0.01562112, 0.02058558, 
    0.0006334089, 9.749882e-08,
  0.0001654378, 0.06808186, 0.08506334, 0.01863873, 0.001173031, 0.052439, 
    0.01447349, 0.0311616, 0.07426641, 0.2283484, 0.03787497, 0.05532386, 
    0.1704139, 0.05994414, 0.02813311, 0.01542914, 0.008790421, 0.001390441, 
    0.004189143, 0.004274736, 0.0001995525, 0.005175074, 0.02618981, 
    0.06724098, 0.02781253, 0.01033377, 0.007803247, 0.0006774931, 0.001608388,
  0.09886888, 0.1284863, 0.1191226, 0.4723929, 0.04359157, 0.01103975, 
    0.08029088, 0.0456798, 0.03498502, 0.02507783, 0.01822526, 0.01860629, 
    0.07859319, 0.0433813, 0.06687364, 0.1263891, 0.1471596, 0.2009807, 
    0.2445957, 0.297267, 0.08416504, 0.114077, 0.1711186, 0.09317122, 
    0.02646836, 0.04900494, 0.09837055, 0.1638716, 0.2718105,
  0.0003008637, 0.0003370371, -2.06923e-07, 0.02858698, 0.007583395, 
    0.02569655, 0.1989967, 0.09386867, 0.3202042, 0.0604853, 0.1080252, 
    0.07254282, 0.03791845, 0.04771216, 0.02204967, 0.02032233, 0.0004045347, 
    3.666955e-07, 0.001982133, 0.00605138, 0.0410893, 0.09011661, 0.01171761, 
    0.009570215, 0.01136161, 0.002226966, 9.716698e-07, 4.646283e-06, 
    0.0004215399,
  1.3499e-06, 0.00180738, 9.175613e-09, 6.504702e-06, 0.0002622826, 
    0.0005643038, 0.05048349, 0.2969512, 0.3462024, 0.0560775, 0.07371332, 
    0.07271366, 0.07209155, 0.04805303, 0.06731369, 0.01091903, 0.01608636, 
    0.0007381325, 0.0001589215, 4.022981e-06, 0.02891766, 0.03541063, 
    0.03939769, 0.01352059, 0.01216112, 0.007284381, 0.0008887108, 
    1.745965e-08, 1.6129e-05,
  0.00246374, 0.0009418063, 0.01248107, 0.01916359, 8.080463e-05, 
    0.004244258, 0.03329267, 0.0129923, 0.02478825, 0.1169382, 0.1384984, 
    0.05584922, 0.1014363, 0.09602924, 0.1258044, 0.1369983, 0.1234663, 
    0.08808148, 0.03139601, 0.0008671691, 0.006587659, 0.005425749, 
    0.04337988, 0.04401608, 0.05499806, 0.04332002, 0.0636986, 0.0296255, 
    0.002592298,
  0.09961596, 0.1592868, 0.1296623, 0.131368, 0.07668278, 0.06151181, 
    0.06901971, 0.09310266, 0.1706933, 0.1794516, 0.1211337, 0.1028783, 
    0.1061809, 0.1744528, 0.08604957, 0.08628311, 0.1619134, 0.1464075, 
    0.1534401, 0.0471772, 0.06881041, 0.02094171, 0.08543187, 0.1443628, 
    0.1551258, 0.1558984, 0.1558725, 0.150036, 0.1455826,
  0.1717662, 0.1366128, 0.1449653, 0.1683802, 0.1578448, 0.2264752, 
    0.2509565, 0.1913864, 0.1642893, 0.1857359, 0.1464463, 0.2090548, 
    0.1762664, 0.2835298, 0.18986, 0.1836396, 0.2246864, 0.3665108, 
    0.4195385, 0.1796799, 0.1267462, 0.1719019, 0.2118322, 0.1857427, 
    0.2096211, 0.3080604, 0.2057972, 0.1965715, 0.1840516,
  0.1610441, 0.1771224, 0.2283501, 0.161915, 0.2094339, 0.1778939, 0.2441766, 
    0.3388645, 0.2397941, 0.1775098, 0.1858019, 0.2119326, 0.2296592, 
    0.2138783, 0.2560461, 0.1997969, 0.244972, 0.2375884, 0.1763768, 
    0.2751207, 0.2338473, 0.2540666, 0.1481214, 0.1294161, 0.104319, 
    0.3580457, 0.2664903, 0.1884871, 0.1710313,
  0.1852717, 0.1947237, 0.1719781, 0.1347354, 0.1744099, 0.1880524, 
    0.1929489, 0.21945, 0.2454694, 0.2308334, 0.2656361, 0.3147386, 
    0.3285867, 0.414647, 0.4436367, 0.3561719, 0.3299253, 0.3083932, 
    0.285094, 0.262971, 0.200884, 0.2627749, 0.2100025, 0.172468, 0.1442469, 
    0.1403233, 0.1659648, 0.09658352, 0.1895043,
  0.05945751, 0.0549075, 0.0503575, 0.04580749, 0.04125749, 0.03670748, 
    0.03215747, 0.04486239, 0.04911573, 0.05336908, 0.05762242, 0.06187576, 
    0.0661291, 0.07038245, 0.07863493, 0.08522812, 0.09182131, 0.0984145, 
    0.1050077, 0.1116009, 0.1181941, 0.1058566, 0.09956011, 0.09326358, 
    0.08696705, 0.08067054, 0.07437401, 0.06807747, 0.06309751,
  0.1082973, 0.0364138, 0.03499579, 0.04170767, 0.007916664, -1.824995e-05, 
    0.001437563, -0.0003817521, 0.004767635, 0.03493117, 0.02499589, 
    0.05596177, 0.07497671, 0.1255053, 0.06591526, 0.1240305, 0.201945, 
    0.2529929, 0.2853217, 0.2685547, 0.3572011, 0.3297281, 0.2174374, 
    0.2257028, 0.1630997, 0.1462065, 0.1674491, 0.2233861, 0.2003068,
  0.2876478, 0.2874336, 0.2622258, 0.1820165, 0.1816348, 0.1981728, 
    0.2026762, 0.2291735, 0.2432619, 0.3330643, 0.3064332, 0.3328233, 
    0.2987209, 0.3115174, 0.3081638, 0.3101585, 0.2560865, 0.2493863, 
    0.2268204, 0.3091294, 0.3386146, 0.3414702, 0.3394756, 0.3877358, 
    0.3256918, 0.2069539, 0.1843248, 0.1878603, 0.2479301,
  0.3125258, 0.2535641, 0.2981955, 0.3070229, 0.3311458, 0.2851949, 
    0.2721558, 0.3027816, 0.3214694, 0.3244887, 0.3678629, 0.2901603, 
    0.3174437, 0.3340561, 0.3050082, 0.2453851, 0.2781205, 0.3321854, 
    0.2969352, 0.2567709, 0.3225695, 0.2876098, 0.271564, 0.2575864, 
    0.2754026, 0.246017, 0.2401937, 0.2538866, 0.306747,
  0.2667947, 0.2356569, 0.2315031, 0.2412938, 0.2292133, 0.2341082, 
    0.2446665, 0.2873893, 0.240029, 0.2595531, 0.2880739, 0.2833286, 
    0.2539673, 0.2056593, 0.19582, 0.2157979, 0.1460569, 0.1971917, 
    0.1979447, 0.223096, 0.2417342, 0.2158824, 0.2270304, 0.2023904, 
    0.1224943, 0.1623801, 0.1829201, 0.2196199, 0.2092153,
  0.1890996, 0.1863807, 0.1161111, 0.1286403, 0.1289774, 0.1211568, 
    0.1387777, 0.1186032, 0.1344012, 0.1403949, 0.1191038, 0.1513983, 
    0.1020892, 0.1124272, 0.1594748, 0.2113444, 0.132349, 0.180964, 
    0.1359696, 0.1494172, 0.2063134, 0.201399, 0.1581466, 0.1533999, 
    0.05428683, 0.0743133, 0.1256131, 0.1679565, 0.2249695,
  0.02949759, 0.005348749, 0.03611617, 0.02154759, 0.06161088, 0.1129122, 
    0.03174271, 0.02530684, 0.02109161, 0.03070112, 0.01290875, 0.01008758, 
    0.08678497, 0.05937052, 0.100736, 0.1550348, 0.1717208, 0.1515383, 
    0.1220397, 0.1087193, 0.09527276, 0.08556225, 0.009712134, 0.00953728, 
    0.07434151, 0.09705902, 0.07744661, 0.06598216, 0.04660317,
  -1.262064e-07, -8.566249e-08, 0.01238788, 0.01282558, 0.05724036, 
    0.02816103, 0.03152996, 0.02787854, 0.02652465, 0.003965938, 
    0.0004391203, 0.04122256, 0.05005368, 0.04651099, 0.07311814, 0.05705569, 
    0.1084709, 0.04024034, 0.06002959, 0.03709189, 0.01253697, 6.953889e-05, 
    1.748964e-07, 3.280946e-05, 0.007745604, 0.03850462, 0.04439625, 
    0.01138799, 0.003857554,
  9.61806e-08, -1.568862e-06, 0.002264882, 0.1492903, 0.0269921, 0.03300187, 
    0.04129282, 0.0875061, 0.03579777, 0.006602746, 0.02307998, 0.009623263, 
    0.1498285, 0.1011864, 0.04794647, 0.05947815, 0.02624297, 0.01127155, 
    0.003793469, 0.0003920642, 5.260175e-07, 1.139233e-07, 5.914793e-07, 
    0.01215331, 0.004244795, 0.00417907, 0.03862443, 0.001709347, 2.486212e-07,
  7.491485e-05, 0.07461943, 0.04292882, 0.02848988, 0.005018668, 0.04846538, 
    0.01397022, 0.03037957, 0.07455466, 0.2182076, 0.04130382, 0.04079146, 
    0.1547001, 0.04965463, 0.03001103, 0.02759621, 0.01697975, 0.002327684, 
    0.0009090651, 0.001581382, 0.00204515, 0.004838389, 0.02148405, 
    0.05804076, 0.02328718, 0.00782521, 0.009678027, 0.001338032, 0.0009789325,
  0.07788152, 0.1049974, 0.1024008, 0.4163425, 0.02692372, 0.004007488, 
    0.08466206, 0.04155277, 0.03007062, 0.02072285, 0.01709059, 0.01889994, 
    0.0738952, 0.04068474, 0.06223296, 0.1191727, 0.1470941, 0.1876336, 
    0.2400925, 0.2726775, 0.0774091, 0.1087733, 0.1846412, 0.08880946, 
    0.02660021, 0.0480692, 0.1003078, 0.1644937, 0.238926,
  8.066892e-05, 0.0002717715, 5.96805e-07, 0.02732901, 0.004012973, 
    0.02084116, 0.1959909, 0.1049185, 0.3249007, 0.05794513, 0.09521067, 
    0.07015865, 0.03592404, 0.04357007, 0.02316956, 0.02341311, 0.003153674, 
    9.488429e-05, 0.003913245, 0.006310264, 0.03383143, 0.09555199, 
    0.01291435, 0.009615823, 0.01755058, 0.009453846, 4.220166e-05, 
    9.61996e-07, 0.0001280623,
  1.058387e-06, 0.0002082132, -5.266297e-08, 3.171942e-06, 0.0001493302, 
    0.0001311773, 0.04227293, 0.3498871, 0.3333969, 0.07374803, 0.07444434, 
    0.07908574, 0.06243478, 0.04542927, 0.05472568, 0.01397235, 0.02698737, 
    0.00387691, 5.679197e-06, 1.690828e-06, 0.01045121, 0.03024791, 
    0.03764787, 0.01330606, 0.01585212, 0.00893662, 0.004781605, 7.95782e-06, 
    6.919089e-06,
  0.0008407101, 0.001273573, 0.01176026, 0.02254164, -8.26617e-05, 
    0.001437295, 0.02191898, 0.00854042, 0.01557769, 0.0845677, 0.1386721, 
    0.06747804, 0.1069275, 0.1008624, 0.1227081, 0.1312846, 0.09328575, 
    0.09709291, 0.03690745, 0.0003563283, 0.004586771, 0.00221844, 
    0.04026654, 0.04245137, 0.05160492, 0.0430155, 0.06784196, 0.03687846, 
    0.002974671,
  0.08533173, 0.1633386, 0.1317267, 0.1373168, 0.051215, 0.04297192, 
    0.0692932, 0.1062059, 0.185069, 0.1748963, 0.1198179, 0.1028047, 
    0.08860161, 0.1664584, 0.09901646, 0.08603394, 0.1599207, 0.1610832, 
    0.1522594, 0.05838493, 0.05079183, 0.01302274, 0.07946116, 0.1533383, 
    0.1513999, 0.1691396, 0.1648149, 0.1437097, 0.139753,
  0.2119986, 0.1443343, 0.1650003, 0.1707379, 0.2109482, 0.2279111, 
    0.2470818, 0.219467, 0.1972529, 0.2028725, 0.1916401, 0.2346355, 
    0.1821915, 0.3120671, 0.1961055, 0.1971977, 0.2695612, 0.3805837, 
    0.421375, 0.1926377, 0.1194013, 0.1525276, 0.1981439, 0.2106447, 
    0.194413, 0.3199657, 0.2415541, 0.260345, 0.2187373,
  0.1827663, 0.2251358, 0.2807099, 0.2010277, 0.2949719, 0.2313189, 
    0.2717414, 0.3469739, 0.2488335, 0.2145604, 0.1967597, 0.2496395, 
    0.2540253, 0.2339182, 0.2885185, 0.19343, 0.2807124, 0.278903, 0.1891432, 
    0.2817384, 0.2457553, 0.2883233, 0.1851606, 0.1210961, 0.1003735, 
    0.3524046, 0.2195067, 0.2035908, 0.1908558,
  0.2355807, 0.2781647, 0.2042975, 0.1509754, 0.1846857, 0.2231409, 
    0.1776723, 0.2399291, 0.2520137, 0.2767064, 0.2975579, 0.312551, 
    0.3118348, 0.4184254, 0.4344749, 0.3712133, 0.3724818, 0.293507, 
    0.2898781, 0.3094504, 0.2222753, 0.2980783, 0.2152475, 0.1741691, 
    0.1253993, 0.1131678, 0.1351884, 0.1059546, 0.2270324,
  0.1256261, 0.1216478, 0.1176696, 0.1136913, 0.109713, 0.1057348, 0.1017565, 
    0.1409045, 0.14797, 0.1550356, 0.1621012, 0.1691668, 0.1762323, 
    0.1832979, 0.1758728, 0.181172, 0.1864712, 0.1917704, 0.1970696, 
    0.2023688, 0.2076679, 0.171023, 0.1626365, 0.15425, 0.1458635, 0.137477, 
    0.1290905, 0.120704, 0.1288087,
  0.1421196, 0.06351845, 0.04902601, 0.0430668, 0.01317557, 0.0005345093, 
    0.002190765, 0.000933696, 0.02818434, 0.0451278, 0.05152698, 0.07108556, 
    0.1065315, 0.1201444, 0.06448396, 0.1426252, 0.21129, 0.2472753, 
    0.2772937, 0.2491974, 0.3891217, 0.3650215, 0.2491609, 0.2313867, 
    0.1600896, 0.1671644, 0.1660443, 0.2230172, 0.1968658,
  0.2953975, 0.270042, 0.270124, 0.1827255, 0.2167381, 0.2012747, 0.2303717, 
    0.2862406, 0.2832031, 0.3608797, 0.330931, 0.3515056, 0.2735779, 
    0.3135764, 0.2846418, 0.2752023, 0.2043976, 0.2144364, 0.2063964, 
    0.3155912, 0.3387686, 0.3320279, 0.3133805, 0.3769986, 0.3276798, 
    0.1565883, 0.1640352, 0.2227143, 0.2538493,
  0.2853655, 0.2429676, 0.2787455, 0.3153621, 0.3443164, 0.2999154, 0.310984, 
    0.3263115, 0.3056692, 0.314492, 0.36659, 0.2812824, 0.2929227, 0.2805863, 
    0.2514696, 0.2229431, 0.2547567, 0.2746145, 0.2877499, 0.3142245, 
    0.3352374, 0.2770908, 0.271954, 0.2384121, 0.2665987, 0.2130107, 
    0.2155249, 0.2414899, 0.2982904,
  0.301283, 0.2438219, 0.2473167, 0.2607035, 0.252139, 0.2643954, 0.2536744, 
    0.311301, 0.2580292, 0.2663379, 0.2970171, 0.27639, 0.2793156, 0.2192615, 
    0.2164783, 0.2294417, 0.163075, 0.2419994, 0.2239028, 0.2343919, 
    0.2464177, 0.2171501, 0.22231, 0.2069294, 0.1112096, 0.1819452, 
    0.1969992, 0.2236732, 0.2382453,
  0.2181656, 0.2182254, 0.1382362, 0.1683518, 0.1449711, 0.1424478, 
    0.1501858, 0.1419507, 0.1636261, 0.1725902, 0.1418851, 0.1628354, 
    0.1047585, 0.1172412, 0.1818372, 0.2193599, 0.1509404, 0.1910958, 
    0.1479639, 0.1558053, 0.2288966, 0.2094521, 0.179015, 0.1644151, 
    0.05466849, 0.09938277, 0.1469254, 0.1927508, 0.2612926,
  0.05191363, 0.01809441, 0.02807988, 0.02922344, 0.06326907, 0.09574109, 
    0.05214522, 0.03167664, 0.04106049, 0.05575731, 0.006426411, 0.005757933, 
    0.07911386, 0.07178675, 0.0967896, 0.1612256, 0.1742653, 0.1504013, 
    0.1251725, 0.1196719, 0.1134182, 0.09261759, 0.01540209, 0.007697331, 
    0.056964, 0.09257741, 0.07806095, 0.07192615, 0.07282402,
  4.786691e-06, 1.869432e-08, 0.001227075, 0.02166271, 0.06693177, 
    0.02723284, 0.03873321, 0.03471445, 0.0325876, 0.001064963, 2.016335e-05, 
    0.008130251, 0.06340864, 0.05322415, 0.07336409, 0.04961874, 0.1219036, 
    0.05077622, 0.06743004, 0.05069233, 0.05212463, 0.001741341, 
    4.668561e-06, 0.0001619355, 0.001451671, 0.06784467, 0.06349643, 
    0.0438687, 0.0168,
  2.044166e-07, 1.755626e-07, 9.695695e-05, 0.1165615, 0.03056344, 
    0.03623931, 0.04728088, 0.09068707, 0.0559388, 0.0152722, 0.03047398, 
    0.02320525, 0.1575432, 0.09618521, 0.05107567, 0.05135513, 0.02483817, 
    0.01309453, 0.009666514, 0.004485783, 6.192441e-05, 5.602566e-07, 
    4.648639e-07, 0.01302926, 0.001401644, 0.0005320398, 0.04328895, 
    0.004791189, 3.468084e-05,
  0.0002305494, 0.09648401, 0.02212874, 0.03484106, 0.01801419, 0.04412003, 
    0.01292685, 0.02965723, 0.07379501, 0.2128091, 0.04273701, 0.03224024, 
    0.1288218, 0.03888128, 0.02650763, 0.02895493, 0.02491822, 0.00741011, 
    0.002908688, 0.002643959, 0.002662481, 0.007205375, 0.01875812, 
    0.05685525, 0.02237626, 0.007373439, 0.01330156, 0.002502181, 0.0001431375,
  0.07317652, 0.08901853, 0.09045186, 0.3472079, 0.007218047, 0.002472345, 
    0.07306282, 0.03504261, 0.02342644, 0.01826051, 0.01923318, 0.01936016, 
    0.06310575, 0.03658079, 0.05394492, 0.1072706, 0.1325822, 0.1784974, 
    0.233734, 0.2511351, 0.08605248, 0.1014411, 0.2007373, 0.08789398, 
    0.02419586, 0.04551658, 0.09308653, 0.1707922, 0.2092912,
  2.659454e-05, 6.207072e-05, 1.129775e-07, 0.02165842, 0.00267705, 
    0.01090292, 0.1931182, 0.1112388, 0.3188812, 0.05406904, 0.0797319, 
    0.06509835, 0.03151423, 0.0378995, 0.02208287, 0.02569966, 0.01117016, 
    0.001902066, 0.008686117, 0.00930262, 0.027264, 0.09206793, 0.01221951, 
    0.009374876, 0.02625589, 0.02517777, 0.002560855, 4.370882e-07, 
    4.282675e-05,
  8.719803e-07, 4.607833e-05, 3.617968e-05, 1.487355e-06, 0.000121822, 
    2.977341e-05, 0.03029615, 0.3408734, 0.331015, 0.0879743, 0.07314051, 
    0.08113679, 0.06007879, 0.04386773, 0.04769772, 0.022337, 0.03956969, 
    0.01261096, 5.341354e-06, 8.095266e-07, 0.004765661, 0.02971116, 
    0.03715113, 0.0125668, 0.01879982, 0.02059608, 0.01873013, 0.00133994, 
    3.268954e-06,
  0.001642838, 0.002190598, 0.01142499, 0.03613704, -4.438447e-05, 
    0.001697159, 0.01288318, 0.00435488, 0.009756068, 0.07319385, 0.1483434, 
    0.08147541, 0.1189657, 0.1058932, 0.1316023, 0.141883, 0.08687162, 
    0.09609444, 0.03630246, 3.878967e-05, 0.002229511, 0.001414312, 
    0.03178985, 0.04193284, 0.05810305, 0.04916281, 0.07700397, 0.05598414, 
    0.006645898,
  0.07984822, 0.1514819, 0.1319928, 0.105004, 0.02541615, 0.04229169, 
    0.04306549, 0.08928191, 0.1848589, 0.1569304, 0.1112436, 0.1077871, 
    0.077402, 0.1745444, 0.1190111, 0.1024984, 0.1545108, 0.1755756, 
    0.1645063, 0.06159416, 0.0315584, 0.01048589, 0.0791071, 0.1542995, 
    0.1599342, 0.1630902, 0.1722165, 0.1538191, 0.138982,
  0.2092164, 0.1494836, 0.1775643, 0.1672886, 0.2000472, 0.2227818, 
    0.2440605, 0.234219, 0.1859344, 0.1850307, 0.1705417, 0.2305582, 
    0.1760834, 0.3355392, 0.1924837, 0.2113322, 0.3083969, 0.3763534, 
    0.4213714, 0.1758358, 0.1280324, 0.1413827, 0.1839236, 0.2365516, 
    0.1931058, 0.3205505, 0.265469, 0.2524941, 0.2243832,
  0.2107897, 0.1967881, 0.3608612, 0.2086264, 0.3340489, 0.2031154, 
    0.2516864, 0.3376598, 0.2688157, 0.2041464, 0.2379756, 0.2435385, 
    0.2284558, 0.1984804, 0.2681358, 0.1677097, 0.2658857, 0.2885812, 
    0.1935559, 0.2873335, 0.2706609, 0.2808392, 0.2224903, 0.1496446, 
    0.1020186, 0.3625186, 0.2405749, 0.2030257, 0.2092135,
  0.2360002, 0.3003553, 0.2524471, 0.1524708, 0.1743976, 0.246767, 0.2288733, 
    0.2126713, 0.192497, 0.2531263, 0.2438702, 0.3227958, 0.3196487, 
    0.3815818, 0.3857933, 0.3682842, 0.35917, 0.2844356, 0.274519, 0.292989, 
    0.2316652, 0.3254811, 0.2354714, 0.1937694, 0.1097975, 0.1140399, 
    0.118269, 0.1450588, 0.249254,
  0.152943, 0.1496197, 0.1462963, 0.142973, 0.1396497, 0.1363264, 0.133003, 
    0.1583239, 0.1679548, 0.1775858, 0.1872168, 0.1968478, 0.2064788, 
    0.2161098, 0.2378643, 0.2415025, 0.2451406, 0.2487788, 0.2524169, 
    0.2560551, 0.2596932, 0.2012059, 0.1912601, 0.1813143, 0.1713685, 
    0.1614227, 0.1514769, 0.1415311, 0.1556017,
  0.1527207, 0.09464213, 0.05208113, 0.0452634, 0.02575453, 0.01769404, 
    0.01700715, 0.01542488, 0.04285257, 0.04675931, 0.07758487, 0.08016931, 
    0.1178656, 0.1157755, 0.06854306, 0.1537098, 0.1928808, 0.2400818, 
    0.2654023, 0.2399223, 0.425823, 0.3894928, 0.280385, 0.231698, 0.1625708, 
    0.1729839, 0.1755211, 0.2167507, 0.1939783,
  0.2905613, 0.2510581, 0.2673617, 0.1776049, 0.2303346, 0.2138076, 
    0.2428627, 0.3194268, 0.3066346, 0.3640121, 0.3389944, 0.3551199, 
    0.2617633, 0.3097214, 0.2899489, 0.2621443, 0.2093066, 0.2131544, 
    0.2298516, 0.3491078, 0.3652123, 0.3348519, 0.2990302, 0.3747735, 
    0.3169369, 0.1615355, 0.1638801, 0.2515129, 0.3010085,
  0.2965737, 0.2471085, 0.3186267, 0.3974752, 0.385933, 0.3231025, 0.3110446, 
    0.3534855, 0.3334281, 0.3566, 0.3620899, 0.3118284, 0.3000337, 0.28628, 
    0.2863498, 0.2658051, 0.2659724, 0.2813898, 0.3213447, 0.3650562, 
    0.3434534, 0.302251, 0.2774275, 0.2365222, 0.280987, 0.2160561, 
    0.2616314, 0.2383033, 0.3290757,
  0.3287098, 0.2833036, 0.2742428, 0.2817942, 0.2961099, 0.291688, 0.2847304, 
    0.3454604, 0.2728748, 0.2821719, 0.3145461, 0.2867877, 0.2752433, 
    0.2389618, 0.2256655, 0.2414571, 0.2206642, 0.2771237, 0.2529835, 
    0.2696219, 0.2655166, 0.2363849, 0.2302565, 0.2187773, 0.1149275, 
    0.2072879, 0.2244296, 0.303095, 0.2880803,
  0.2564633, 0.2562994, 0.1931343, 0.2414418, 0.1986909, 0.224695, 0.1802679, 
    0.159418, 0.2025534, 0.2001058, 0.1847505, 0.1893535, 0.1145981, 
    0.1382263, 0.1983957, 0.2377707, 0.1813493, 0.2038387, 0.1788455, 
    0.1809374, 0.245158, 0.2327574, 0.1953464, 0.1813128, 0.05533149, 
    0.1469101, 0.217147, 0.2764102, 0.308619,
  0.1137693, 0.03408568, 0.02074648, 0.04664692, 0.07432877, 0.09467636, 
    0.08135015, 0.06896316, 0.08825164, 0.1024982, 0.005533015, 0.0002910214, 
    0.05406506, 0.1320633, 0.1141117, 0.166245, 0.1734867, 0.1635869, 
    0.1640251, 0.1284252, 0.138532, 0.1275163, 0.04713168, 0.008763922, 
    0.05726344, 0.1006261, 0.1063329, 0.1098268, 0.09211513,
  0.03303909, -1.65626e-07, 3.364481e-05, 0.02111483, 0.07120219, 0.03378589, 
    0.06801215, 0.1092402, 0.1543132, 0.0130524, -6.197032e-06, 0.0009762351, 
    0.06050926, 0.07851557, 0.08775806, 0.04444882, 0.1135954, 0.05600727, 
    0.06469214, 0.06956698, 0.08966838, 0.07023493, 0.005882432, 
    0.0002064037, 0.000837252, 0.02735725, 0.05356086, 0.1155308, 0.05868324,
  2.517384e-06, 4.027862e-06, 2.200668e-05, 0.05642125, 0.03139924, 
    0.04439459, 0.06030216, 0.08957319, 0.06546818, 0.02876041, 0.03098062, 
    0.03292921, 0.1814447, 0.0897608, 0.05197205, 0.04312446, 0.0247582, 
    0.01510902, 0.01614155, 0.01915412, 0.002134508, 5.983998e-05, 
    2.86912e-07, 0.01544396, 0.0008400059, 8.901765e-05, 0.03958204, 
    0.02735963, 0.001005533,
  0.0010345, 0.1185948, 0.01610952, 0.02788824, 0.03034917, 0.04501187, 
    0.01245228, 0.02681119, 0.06780019, 0.1991163, 0.04161617, 0.02433409, 
    0.1052497, 0.03211139, 0.02384125, 0.02392829, 0.02878283, 0.01733452, 
    0.01446288, 0.01233986, 0.002006226, 0.006213626, 0.01437419, 0.05957277, 
    0.02449924, 0.007407051, 0.01641485, 0.01206318, 0.001172237,
  0.0872069, 0.07887784, 0.08150515, 0.2938668, 0.0007944938, 0.005627946, 
    0.05732104, 0.03073451, 0.01716366, 0.01753076, 0.04997048, 0.02007268, 
    0.05161481, 0.03098948, 0.04350742, 0.09123309, 0.1131391, 0.1669789, 
    0.2024537, 0.224151, 0.08503924, 0.08811273, 0.2033967, 0.08888878, 
    0.02246073, 0.04052128, 0.08044761, 0.1539272, 0.1844035,
  4.650168e-06, 8.677749e-06, 3.076092e-08, 0.0152731, 0.002083613, 
    0.004600297, 0.1960874, 0.1051322, 0.3054398, 0.04848351, 0.06463826, 
    0.05528091, 0.0278286, 0.03267151, 0.0233755, 0.03233991, 0.02424105, 
    0.01006538, 0.01076418, 0.01763829, 0.02342649, 0.09034157, 0.0130099, 
    0.01064379, 0.03365947, 0.03809637, 0.008871318, 2.547797e-07, 
    1.185694e-05,
  7.423145e-07, 1.261446e-05, 2.332792e-05, 6.389678e-07, 4.411678e-05, 
    3.558192e-06, 0.02122292, 0.3013015, 0.3316602, 0.09190004, 0.07062506, 
    0.07572643, 0.05799134, 0.04017866, 0.03971829, 0.0283716, 0.04642327, 
    0.05365874, 0.0005399601, 2.959614e-07, 0.001817926, 0.0295364, 
    0.03575943, 0.0133343, 0.01894267, 0.0270912, 0.04054206, 0.005303744, 
    1.913861e-06,
  0.003112558, 0.005173332, 0.006027049, 0.06589851, -4.266014e-05, 
    0.000487147, 0.008283583, 0.001657922, 0.009542472, 0.07149561, 
    0.1635723, 0.09813508, 0.1342382, 0.120806, 0.1552825, 0.1584484, 
    0.1143106, 0.1302448, 0.05936393, -5.867008e-05, 0.0006399213, 
    0.000701444, 0.02656485, 0.04255658, 0.06454237, 0.0534223, 0.105016, 
    0.09542488, 0.009550005,
  0.1078561, 0.1646518, 0.1413558, 0.08236526, 0.02311282, 0.03031895, 
    0.0377388, 0.09068161, 0.182729, 0.1331331, 0.1120705, 0.1062437, 
    0.09220413, 0.2029076, 0.1285803, 0.1011818, 0.1834499, 0.2036318, 
    0.2166711, 0.07694621, 0.02146376, 0.01007505, 0.08935578, 0.1637045, 
    0.1580605, 0.1774957, 0.222637, 0.1831804, 0.1404129,
  0.1994071, 0.1767402, 0.1796045, 0.1896458, 0.2086428, 0.2125438, 
    0.2376374, 0.2265862, 0.1879893, 0.197364, 0.1799529, 0.2575133, 
    0.1972584, 0.3596313, 0.2123076, 0.2649409, 0.3425776, 0.3948286, 
    0.429356, 0.1642882, 0.1472562, 0.1518315, 0.1664531, 0.2613516, 
    0.2043654, 0.2971806, 0.3025268, 0.3053415, 0.2488932,
  0.2354089, 0.2331908, 0.3765048, 0.271093, 0.2999812, 0.1868026, 0.259935, 
    0.366222, 0.2899125, 0.2116394, 0.2486876, 0.2833977, 0.2489613, 
    0.2447427, 0.3005517, 0.1809802, 0.2980247, 0.2676569, 0.2091969, 
    0.2747377, 0.276577, 0.2944849, 0.2312935, 0.1420487, 0.1107279, 
    0.3823275, 0.2527185, 0.2037971, 0.2234828,
  0.2895382, 0.3072222, 0.2749277, 0.2277993, 0.2075745, 0.2908115, 
    0.2654389, 0.231244, 0.2159815, 0.2576781, 0.2290449, 0.402571, 
    0.3625677, 0.4298698, 0.4194004, 0.3771191, 0.3531646, 0.3014767, 
    0.2983172, 0.2799985, 0.2355762, 0.3302328, 0.2744096, 0.2250082, 
    0.1178628, 0.1426869, 0.1395537, 0.1522393, 0.2962198,
  0.1899526, 0.1873677, 0.1847828, 0.1821979, 0.179613, 0.1770281, 0.1744432, 
    0.1919765, 0.201686, 0.2113955, 0.221105, 0.2308145, 0.240524, 0.2502335, 
    0.2666636, 0.2693407, 0.2720178, 0.274695, 0.2773722, 0.2800493, 
    0.2827265, 0.2378759, 0.2280742, 0.2182725, 0.2084707, 0.198669, 
    0.1888673, 0.1790655, 0.1920206,
  0.1569602, 0.1078829, 0.05281364, 0.05192288, 0.03439905, 0.03999233, 
    0.04988926, 0.03335383, 0.06427953, 0.06820808, 0.08874188, 0.08913197, 
    0.1377326, 0.1049217, 0.0693945, 0.1572587, 0.1962253, 0.2310944, 
    0.2572458, 0.2173293, 0.4479937, 0.4032569, 0.3011772, 0.2401865, 
    0.180791, 0.1633871, 0.1835751, 0.2025393, 0.1939783,
  0.3029061, 0.2373115, 0.2682916, 0.1707682, 0.2383013, 0.213745, 0.2093377, 
    0.3393687, 0.3274879, 0.370876, 0.3451579, 0.3264824, 0.2651005, 
    0.311424, 0.3147324, 0.296504, 0.2614462, 0.2203209, 0.301706, 0.3762456, 
    0.3741979, 0.3174778, 0.3077059, 0.3780556, 0.2997546, 0.1791723, 
    0.1583299, 0.254848, 0.3131693,
  0.3412758, 0.3096282, 0.4297695, 0.4337969, 0.4272294, 0.3619059, 
    0.3047236, 0.3952638, 0.4013363, 0.3801046, 0.3596377, 0.3188355, 
    0.3699219, 0.3247963, 0.3415694, 0.3353299, 0.3271018, 0.34224, 
    0.3780218, 0.4241183, 0.2798667, 0.2545786, 0.2855609, 0.2337034, 
    0.2821063, 0.2294168, 0.272158, 0.3114022, 0.3824177,
  0.2887788, 0.2729639, 0.2680832, 0.2997177, 0.3067728, 0.3094921, 
    0.3110962, 0.328021, 0.2714347, 0.2822576, 0.2989916, 0.3022928, 
    0.2851608, 0.2666204, 0.2619964, 0.2832764, 0.3039348, 0.3216913, 
    0.287895, 0.3344885, 0.3011178, 0.2347053, 0.2493364, 0.2359174, 
    0.1239293, 0.2283555, 0.3060608, 0.331529, 0.2921777,
  0.3086409, 0.2569554, 0.190732, 0.2260425, 0.2540014, 0.241504, 0.2271295, 
    0.2155558, 0.212773, 0.1728872, 0.1656942, 0.1597973, 0.09673724, 
    0.1794768, 0.2230669, 0.2418321, 0.2305166, 0.234347, 0.2063721, 
    0.230737, 0.2558904, 0.272781, 0.2226094, 0.1995806, 0.05453774, 
    0.1992523, 0.2673558, 0.2786237, 0.2999548,
  0.1740204, 0.07254665, 0.01479414, 0.08609332, 0.08995843, 0.1085243, 
    0.08683833, 0.207144, 0.138767, 0.1604497, 0.002815901, -3.331551e-06, 
    0.03855339, 0.1231633, 0.1393739, 0.1802298, 0.2067103, 0.183101, 
    0.1620492, 0.1601244, 0.1597311, 0.2029083, 0.1178238, 0.01188981, 
    0.06224542, 0.1318129, 0.1738191, 0.1558064, 0.1362112,
  0.1112285, -4.505083e-05, -5.564128e-06, 0.04491006, 0.06768808, 
    0.04842804, 0.09132448, 0.1943038, 0.1905859, 0.01408214, -7.286753e-07, 
    0.0001970936, 0.09454612, 0.1650014, 0.119432, 0.06018924, 0.09715501, 
    0.05240599, 0.07445341, 0.1148132, 0.1826122, 0.2100437, 0.06139717, 
    -0.0002354923, 0.0003692391, 0.01347256, 0.05784892, 0.149049, 0.3075446,
  0.0005806152, 3.152341e-05, -6.194962e-05, 0.02315601, 0.0343884, 
    0.0436174, 0.06048495, 0.08284467, 0.06590781, 0.03775499, 0.02899516, 
    0.03496211, 0.1975997, 0.0907837, 0.05314307, 0.04315203, 0.03001574, 
    0.02094535, 0.02293567, 0.03493945, 0.03924045, 0.02774503, -3.06966e-05, 
    0.01682333, 0.0004066905, 1.355609e-05, 0.06074934, 0.05836374, 0.012702,
  0.01657931, 0.1432717, 0.01431577, 0.0221799, 0.03607405, 0.04621439, 
    0.01470192, 0.02735418, 0.05969723, 0.1848267, 0.04031911, 0.02291823, 
    0.0830005, 0.02884844, 0.02388715, 0.02170989, 0.02221913, 0.01390182, 
    0.01569293, 0.0266706, 0.002729244, 0.003726445, 0.00961569, 0.07418942, 
    0.02728114, 0.01070086, 0.02334784, 0.03941124, 0.01145014,
  0.09578885, 0.07391109, 0.06578179, 0.2581411, -0.0002825177, 0.01453263, 
    0.04476388, 0.02831282, 0.01416667, 0.01968243, 0.03006064, 0.02541865, 
    0.04191285, 0.02810173, 0.03793932, 0.07496982, 0.09163009, 0.1453756, 
    0.1663155, 0.1909581, 0.08051753, 0.07786597, 0.2002907, 0.08639215, 
    0.02282445, 0.03949865, 0.06918398, 0.1396694, 0.1712856,
  4.15175e-07, 2.843489e-07, 1.847878e-08, 0.009530176, 0.001964525, 
    0.002770931, 0.1899313, 0.09877482, 0.2750086, 0.04380603, 0.05127507, 
    0.0466177, 0.02727031, 0.03328653, 0.02686998, 0.03800036, 0.08110986, 
    0.06339717, 0.008810965, 0.03361773, 0.02302993, 0.08894931, 0.01594476, 
    0.01379018, 0.04260841, 0.0608657, 0.04015383, -4.054072e-06, 2.057653e-06,
  6.508374e-07, 2.055679e-06, 0.0006037169, 2.766508e-07, 4.100029e-05, 
    -2.908273e-06, 0.01265834, 0.2702884, 0.3358538, 0.08276458, 0.07608593, 
    0.07444204, 0.05266699, 0.04292382, 0.0410955, 0.03524087, 0.06238349, 
    0.1067408, 0.02022118, 9.341013e-08, 0.0009522729, 0.02757317, 
    0.03835234, 0.01808702, 0.02792068, 0.03675805, 0.07975268, 0.01580754, 
    1.259442e-06,
  0.009581791, 0.0027034, 0.003105912, 0.1107652, -2.613731e-05, 
    -2.018434e-05, 0.006685938, 0.0003283119, 0.008903999, 0.06574731, 
    0.1690379, 0.1001934, 0.1480493, 0.1394801, 0.1843291, 0.1841853, 
    0.1676559, 0.1777987, 0.09638909, -5.055311e-05, 9.200423e-05, 
    0.0003739324, 0.02751509, 0.04033534, 0.07450847, 0.08694349, 0.1129936, 
    0.1242835, 0.01105732,
  0.112299, 0.190487, 0.1370647, 0.09106954, 0.02390279, 0.02413236, 
    0.03246383, 0.1026489, 0.1941065, 0.1355529, 0.1129058, 0.1157028, 
    0.09821771, 0.2305151, 0.1402792, 0.1272035, 0.203051, 0.219066, 
    0.2504075, 0.06477454, 0.01859461, 0.009187241, 0.08991572, 0.177423, 
    0.1509558, 0.2179061, 0.2733911, 0.2106836, 0.1748956,
  0.2137519, 0.1764893, 0.1785874, 0.1733294, 0.1820325, 0.1811825, 
    0.2296608, 0.1962077, 0.1716991, 0.1909421, 0.173551, 0.2875588, 
    0.2145545, 0.3810868, 0.2325017, 0.2909702, 0.3673537, 0.38495, 
    0.4352747, 0.1526715, 0.1329581, 0.163538, 0.1718808, 0.3051781, 
    0.2207298, 0.2639981, 0.4192891, 0.3521692, 0.299054,
  0.2857021, 0.3037386, 0.4506967, 0.3050439, 0.2940736, 0.2154288, 
    0.3323328, 0.3782418, 0.2898396, 0.28022, 0.3028001, 0.3302668, 
    0.3241633, 0.2823047, 0.3214154, 0.2487529, 0.3139177, 0.2697491, 
    0.1793792, 0.2797889, 0.2749824, 0.3254883, 0.2515785, 0.1531082, 
    0.0998048, 0.3672439, 0.253576, 0.2039093, 0.2500364,
  0.3105076, 0.346968, 0.2430729, 0.2401669, 0.2523497, 0.3073258, 0.2630881, 
    0.2874887, 0.2700584, 0.3126327, 0.3840786, 0.4377915, 0.4318588, 
    0.4801807, 0.4550918, 0.4091584, 0.375773, 0.3349604, 0.3259818, 
    0.3231165, 0.3107404, 0.3478263, 0.2975527, 0.2601093, 0.1396259, 
    0.1648715, 0.1271707, 0.1818313, 0.2969216,
  0.1991061, 0.1983532, 0.1976003, 0.1968474, 0.1960945, 0.1953416, 
    0.1945887, 0.2239542, 0.2336641, 0.2433741, 0.2530841, 0.262794, 
    0.272504, 0.2822139, 0.2851718, 0.2861609, 0.2871501, 0.2881393, 
    0.2891285, 0.2901176, 0.2911068, 0.2544462, 0.2444999, 0.2345537, 
    0.2246074, 0.2146612, 0.204715, 0.1947687, 0.1997084,
  0.1576476, 0.1074659, 0.05795636, 0.05845407, 0.05215759, 0.06615621, 
    0.06911514, 0.07434314, 0.06866469, 0.0733102, 0.09753773, 0.1088839, 
    0.1499306, 0.0766804, 0.06597398, 0.156928, 0.2190626, 0.2178586, 
    0.2421428, 0.2068596, 0.4674426, 0.419568, 0.3221657, 0.2309765, 
    0.1740732, 0.1522599, 0.1722528, 0.1997607, 0.1965015,
  0.2996612, 0.2409067, 0.2564923, 0.1544662, 0.2559356, 0.2186112, 
    0.1668589, 0.3403562, 0.3440505, 0.3819926, 0.3499166, 0.2983322, 
    0.2623817, 0.289352, 0.3255294, 0.3593954, 0.3217748, 0.2633821, 
    0.3886095, 0.3709301, 0.369012, 0.3517618, 0.3426937, 0.396212, 
    0.3099843, 0.2126214, 0.1953673, 0.2330502, 0.3162095,
  0.4131509, 0.3627578, 0.498586, 0.4185869, 0.4345143, 0.4073091, 0.3212414, 
    0.4556385, 0.4392178, 0.3600021, 0.3767527, 0.3294674, 0.4026071, 
    0.3848885, 0.3545767, 0.3537332, 0.3710203, 0.4465573, 0.4401799, 
    0.3411218, 0.247345, 0.2318951, 0.2640088, 0.2550713, 0.3064122, 
    0.2721351, 0.3135291, 0.3574107, 0.3910123,
  0.2526216, 0.2547881, 0.2575623, 0.287118, 0.3094225, 0.315598, 0.3273201, 
    0.3063595, 0.2574091, 0.2453367, 0.2646328, 0.3024985, 0.2572414, 
    0.2693334, 0.3278797, 0.2928821, 0.3367904, 0.3268797, 0.3220652, 
    0.3010012, 0.2795544, 0.2689037, 0.2748484, 0.2712371, 0.1328676, 
    0.232017, 0.3577023, 0.318407, 0.275385,
  0.2738447, 0.2150237, 0.148812, 0.2100846, 0.2412428, 0.2274626, 0.2383854, 
    0.232245, 0.209547, 0.155022, 0.1374018, 0.112799, 0.05705197, 0.1739185, 
    0.2693129, 0.2210358, 0.2140559, 0.2748511, 0.1770338, 0.2116469, 
    0.2128354, 0.2526311, 0.1871004, 0.2465779, 0.0504848, 0.1986426, 
    0.2414085, 0.232453, 0.2892796,
  0.2217519, 0.1135038, 0.01385244, 0.08913622, 0.1347531, 0.1176823, 
    0.2297498, 0.2824008, 0.2223048, 0.08452755, 0.000516855, 0.0001230569, 
    0.02610132, 0.08241273, 0.09927857, 0.1661836, 0.1779445, 0.1582051, 
    0.1347065, 0.1281375, 0.1417698, 0.1929584, 0.1528258, 0.01474168, 
    0.06146839, 0.1554477, 0.1966635, 0.1649617, 0.1775623,
  0.3410548, 6.317579e-05, -1.117754e-05, 0.04258352, 0.08157608, 0.05769902, 
    0.09918136, 0.1791151, 0.1934784, 0.01104189, 6.755972e-08, 8.499315e-05, 
    0.1223669, 0.1935135, 0.1579461, 0.09269296, 0.0952128, 0.06059655, 
    0.09070858, 0.1770616, 0.1986082, 0.3506227, 0.2048269, 0.002649155, 
    0.001285323, 0.00859383, 0.1090108, 0.1456336, 0.4364308,
  0.009413899, 0.002207555, -3.212476e-05, 0.01140102, 0.04489569, 
    0.05406378, 0.07041138, 0.08638974, 0.08009906, 0.1017341, 0.03183287, 
    0.06051769, 0.1997356, 0.101694, 0.06246497, 0.05919272, 0.0741632, 
    0.04936597, 0.04248001, 0.07821223, 0.1500415, 0.1371476, 0.004165297, 
    0.01302885, 0.0001744716, 2.373434e-06, 0.09892999, 0.07393971, 0.1667618,
  0.09207815, 0.2084053, 0.00971311, 0.02492078, 0.04227126, 0.04770476, 
    0.03175187, 0.03100415, 0.05115535, 0.1681058, 0.04644229, 0.02428378, 
    0.07360646, 0.03144474, 0.03256711, 0.02397717, 0.0168094, 0.01128684, 
    0.01211038, 0.03309389, 0.0221776, 0.001063183, 0.006886984, 0.06163747, 
    0.01880555, 0.02117748, 0.04370133, 0.07185347, 0.0579765,
  0.09697109, 0.07284051, 0.04628703, 0.2306457, -0.0003081537, 0.01786416, 
    0.03268467, 0.03226572, 0.01096133, 0.0250987, 0.01606097, 0.03257107, 
    0.04034591, 0.0374622, 0.03691821, 0.06741057, 0.08246689, 0.1259005, 
    0.1412247, 0.1508555, 0.07747274, 0.06998694, 0.1964766, 0.08251752, 
    0.02765742, 0.04280357, 0.06513463, 0.12142, 0.1553516,
  -3.707493e-08, -5.587047e-07, 1.448486e-08, 0.007852237, 0.001493588, 
    0.01497252, 0.1544293, 0.09001338, 0.2442507, 0.02964103, 0.04546671, 
    0.05266266, 0.03262933, 0.03725972, 0.03385711, 0.04962977, 0.1661037, 
    0.1627054, 0.05379915, 0.05178964, 0.02568865, 0.09413431, 0.02362599, 
    0.01683288, 0.04973772, 0.08919307, 0.07471915, 0.0004674544, 1.148287e-06,
  5.951679e-07, -5.200836e-06, 0.001704989, 1.470606e-07, 2.908045e-06, 
    -8.411772e-07, 0.006848652, 0.2795717, 0.3156701, 0.0619711, 0.09386224, 
    0.07734716, 0.05999032, 0.04859208, 0.04696973, 0.0422609, 0.07433274, 
    0.1431473, 0.07491945, 3.925053e-07, 0.0003486575, 0.02507807, 
    0.03454625, 0.02798837, 0.04215893, 0.0500133, 0.1050221, 0.08841512, 
    -9.835087e-07,
  0.01201436, 0.001844438, 0.001183589, 0.1594197, -2.28387e-05, 
    -4.963285e-05, 0.007837069, 3.83954e-05, 0.006884815, 0.05670559, 
    0.1601313, 0.1077282, 0.2002113, 0.1881473, 0.2226704, 0.1920237, 
    0.2246989, 0.2210554, 0.2143407, -3.703311e-05, 3.058297e-05, 
    0.000194172, 0.02335582, 0.03373738, 0.08552548, 0.1137771, 0.1516398, 
    0.2164135, 0.03102622,
  0.1076411, 0.169641, 0.1526027, 0.07840261, 0.0238925, 0.01640251, 
    0.01935109, 0.1097716, 0.1820383, 0.1367345, 0.1077236, 0.1086101, 
    0.1031637, 0.2617254, 0.1698212, 0.2426486, 0.3268856, 0.3140993, 
    0.2604611, 0.04736131, 0.01535769, 0.005911615, 0.09413606, 0.1675245, 
    0.1337811, 0.2514448, 0.3170404, 0.2812094, 0.2213042,
  0.2334076, 0.1396278, 0.153327, 0.1438, 0.1498201, 0.1779167, 0.2051295, 
    0.1840839, 0.140257, 0.1915995, 0.1611605, 0.2995068, 0.2119129, 
    0.4014055, 0.2621193, 0.3331346, 0.376782, 0.3625398, 0.426807, 
    0.1429588, 0.1187448, 0.1709815, 0.2174753, 0.3084306, 0.278357, 
    0.2311458, 0.4941074, 0.4125528, 0.2825263,
  0.397141, 0.3465287, 0.466997, 0.3227862, 0.3659382, 0.2565033, 0.3772144, 
    0.3835009, 0.259518, 0.3117512, 0.3268085, 0.3380785, 0.3682985, 
    0.3201727, 0.2989171, 0.334248, 0.3393744, 0.2891558, 0.2338821, 
    0.3057783, 0.2991486, 0.3778118, 0.2849053, 0.1772203, 0.1054591, 
    0.3437062, 0.242954, 0.2065044, 0.3281763,
  0.3237242, 0.4066604, 0.3053725, 0.293391, 0.3351859, 0.3490773, 0.322468, 
    0.3731727, 0.3887001, 0.4049703, 0.4896611, 0.5205384, 0.5289316, 
    0.5289187, 0.4924778, 0.4585075, 0.4601367, 0.3816351, 0.4123089, 
    0.4154891, 0.3824637, 0.3549902, 0.3066249, 0.2858559, 0.1851812, 
    0.1536447, 0.1321899, 0.2120527, 0.2807019,
  0.2091736, 0.208894, 0.2086144, 0.2083348, 0.2080552, 0.2077757, 0.2074961, 
    0.2240416, 0.2341419, 0.2442421, 0.2543423, 0.2644426, 0.2745428, 
    0.2846431, 0.2956977, 0.2947975, 0.2938974, 0.2929972, 0.2920971, 
    0.291197, 0.2902968, 0.2582927, 0.2493722, 0.2404517, 0.2315312, 
    0.2226107, 0.2136902, 0.2047697, 0.2093973,
  0.1618874, 0.1090603, 0.05651961, 0.06026833, 0.0636774, 0.08707343, 
    0.09816337, 0.09338923, 0.07007517, 0.07873838, 0.1082794, 0.1314171, 
    0.1602998, 0.05110544, 0.06606212, 0.1408305, 0.225884, 0.2102787, 
    0.2213265, 0.1957614, 0.5073708, 0.4736948, 0.3310791, 0.212315, 
    0.166934, 0.1538488, 0.1692411, 0.1977163, 0.2043113,
  0.2820315, 0.2378459, 0.2329247, 0.1222488, 0.2511088, 0.2262381, 
    0.1062004, 0.3316643, 0.358105, 0.3805946, 0.3515905, 0.2739066, 
    0.2384735, 0.2580105, 0.345715, 0.3829608, 0.3663706, 0.2830783, 
    0.4330493, 0.3464611, 0.3787657, 0.3789707, 0.3742802, 0.4049429, 
    0.3153681, 0.2565651, 0.2620004, 0.2349479, 0.3207108,
  0.4323368, 0.3928556, 0.4745009, 0.3213065, 0.3862137, 0.4904205, 
    0.3435079, 0.5029229, 0.4138335, 0.2818644, 0.3407069, 0.3443335, 
    0.4345902, 0.443665, 0.3922786, 0.3840848, 0.4526327, 0.4526865, 
    0.416523, 0.2488489, 0.1890785, 0.1891697, 0.2573067, 0.2824336, 
    0.3341327, 0.3167043, 0.3488611, 0.3905819, 0.4318472,
  0.2510794, 0.2318687, 0.2318352, 0.2866542, 0.3166893, 0.3301099, 
    0.3278245, 0.2771202, 0.2492286, 0.2259815, 0.2269313, 0.2802824, 
    0.2324371, 0.2236218, 0.3084008, 0.2532744, 0.2755182, 0.309993, 
    0.2639033, 0.2363283, 0.2428115, 0.2617071, 0.2546158, 0.2956407, 
    0.1248156, 0.2518755, 0.340615, 0.2945434, 0.2632126,
  0.2322126, 0.1533191, 0.09346724, 0.2013154, 0.2016672, 0.1874196, 
    0.1954746, 0.1746463, 0.18671, 0.1138841, 0.1292186, 0.07121451, 
    0.02791234, 0.1265986, 0.30493, 0.1680502, 0.1679108, 0.252331, 
    0.1397285, 0.1769011, 0.193417, 0.2177718, 0.1907856, 0.2804459, 
    0.04659494, 0.1349757, 0.1946579, 0.2146417, 0.2951404,
  0.1912685, 0.1431254, 0.01180636, 0.06443037, 0.1218986, 0.1335569, 
    0.1821686, 0.1713515, 0.1631595, 0.02096593, 0.0001459844, 2.597173e-05, 
    0.02165212, 0.04128136, 0.08075073, 0.1550503, 0.1360074, 0.145716, 
    0.1198, 0.1061547, 0.1262396, 0.1889889, 0.1504802, 0.01660118, 
    0.06610553, 0.1232535, 0.1389407, 0.1561337, 0.1707386,
  0.5374123, 0.001769205, -4.044621e-06, 0.03703816, 0.1023097, 0.03966533, 
    0.04837288, 0.07968503, 0.114919, 0.003226602, 4.972393e-08, 
    2.346831e-05, 0.07106645, 0.117001, 0.1335157, 0.105088, 0.1168713, 
    0.1059555, 0.09844309, 0.0952521, 0.0942148, 0.29667, 0.5056099, 
    0.003265492, 0.003756697, 0.009976627, 0.05134933, 0.07604508, 0.2218918,
  0.2746548, 0.03566857, -3.835941e-05, 0.008523071, 0.04696511, 0.06229679, 
    0.09666941, 0.08119697, 0.06738575, 0.08303865, 0.04247662, 0.05516884, 
    0.196657, 0.1204175, 0.06370354, 0.04276307, 0.0419166, 0.02727188, 
    0.02128848, 0.03859203, 0.1280451, 0.4051092, 0.0198745, 0.00601674, 
    6.967372e-05, 6.287823e-07, 0.07484508, 0.06582874, 0.3636883,
  0.2338684, 0.2193418, 0.004605583, 0.03224361, 0.04653992, 0.1140367, 
    0.1307141, 0.1094809, 0.03345881, 0.1452479, 0.07683796, 0.03223957, 
    0.08886627, 0.04188322, 0.03005494, 0.02578627, 0.01962053, 0.01512683, 
    0.01582535, 0.02306848, 0.08674014, 0.01871646, 0.007896574, 0.03245784, 
    0.007184988, 0.07631834, 0.07512207, 0.1415998, 0.1588155,
  0.09067526, 0.0613519, 0.03101332, 0.2017881, -0.0001897905, 0.01676788, 
    0.02824886, 0.04775298, 0.008298095, 0.05399939, 0.01207799, 0.1285708, 
    0.05269372, 0.04662566, 0.04264132, 0.06039934, 0.07867329, 0.1152499, 
    0.1312169, 0.1293674, 0.09855981, 0.07010714, 0.1816063, 0.07290231, 
    0.05061885, 0.05880333, 0.07921447, 0.1199768, 0.1382853,
  -8.546189e-08, -1.24074e-07, 1.261174e-08, 0.004802225, 0.0006577535, 
    0.03999544, 0.107058, 0.07863366, 0.2061425, 0.02397209, 0.05533557, 
    0.05507722, 0.03577747, 0.062877, 0.033466, 0.05230777, 0.09605761, 
    0.2147657, 0.3322473, 0.07380684, 0.02939105, 0.1068415, 0.04648231, 
    0.0281534, 0.05526184, 0.1143267, 0.1880825, 0.01761853, -6.297797e-07,
  5.594758e-07, -6.387368e-05, 0.003222199, 1.038654e-07, 4.963362e-07, 
    -1.494217e-06, 0.003041422, 0.312393, 0.2951374, 0.0419567, 0.1220118, 
    0.07317943, 0.1020161, 0.07220348, 0.0728936, 0.05904776, 0.07117409, 
    0.1676579, 0.3112669, 0.0001067898, 0.0001654961, 0.02142627, 0.02700313, 
    0.1352411, 0.06002488, 0.1057018, 0.1149965, 0.2312286, -0.0002343321,
  0.01311635, 0.001176094, 0.0005799185, 0.2046418, -2.887742e-05, 
    -2.441882e-05, 0.005602067, -1.943778e-06, 0.005286977, 0.05174428, 
    0.1425164, 0.1253805, 0.2418812, 0.2332432, 0.2406446, 0.2101749, 
    0.3330408, 0.2130729, 0.3927395, -6.382962e-05, 1.227444e-05, 
    5.297148e-05, 0.01457181, 0.0519803, 0.1170178, 0.2145322, 0.210497, 
    0.2468047, 0.06200017,
  0.09937686, 0.1617816, 0.1076731, 0.06696214, 0.02283245, 0.01748182, 
    0.01430916, 0.1069465, 0.1655945, 0.1333094, 0.08946264, 0.103044, 
    0.1207325, 0.3060211, 0.3103791, 0.3762242, 0.4568107, 0.4188234, 
    0.3067262, 0.04364425, 0.01857129, 0.01001491, 0.1035716, 0.1588707, 
    0.1280776, 0.2849938, 0.3557727, 0.2802421, 0.2277983,
  0.2430542, 0.1325741, 0.1208607, 0.1114096, 0.1353126, 0.1391178, 
    0.1809971, 0.1451627, 0.1205403, 0.1869726, 0.1426652, 0.2882776, 
    0.1985548, 0.3912716, 0.249538, 0.4294795, 0.3754453, 0.3374236, 
    0.3923548, 0.112514, 0.08511962, 0.1766738, 0.2660013, 0.2968083, 
    0.3517157, 0.1971574, 0.4985859, 0.3747204, 0.2931918,
  0.5562117, 0.3986478, 0.484482, 0.3892382, 0.4652857, 0.3640357, 0.4403176, 
    0.4212415, 0.252663, 0.3251545, 0.3494796, 0.3945775, 0.3671934, 
    0.3700663, 0.3381753, 0.4767874, 0.3884636, 0.3619849, 0.2971946, 
    0.3609542, 0.395963, 0.4685188, 0.3343872, 0.2468047, 0.1866558, 
    0.3204626, 0.2554264, 0.217085, 0.4785624,
  0.4111169, 0.4803041, 0.4852755, 0.4883272, 0.5130004, 0.4459836, 
    0.4193791, 0.5064046, 0.5467199, 0.5477792, 0.5277939, 0.5560545, 
    0.5625955, 0.6000968, 0.6174493, 0.5916239, 0.6381575, 0.538167, 
    0.5256637, 0.5245125, 0.5165728, 0.4210191, 0.3462832, 0.3260294, 
    0.2158521, 0.1749265, 0.13989, 0.2546629, 0.3510175,
  0.207143, 0.2068332, 0.2065234, 0.2062136, 0.2059038, 0.205594, 0.2052842, 
    0.2074384, 0.2178737, 0.2283089, 0.2387441, 0.2491794, 0.2596146, 
    0.2700499, 0.2831745, 0.2802994, 0.2774243, 0.2745492, 0.271674, 
    0.2687989, 0.2659238, 0.2377022, 0.2304519, 0.2232016, 0.2159513, 
    0.2087009, 0.2014506, 0.1942003, 0.2073908,
  0.1862756, 0.1030397, 0.05583272, 0.05967657, 0.07056529, 0.09719772, 
    0.121256, 0.106005, 0.06181004, 0.07774016, 0.1164767, 0.1441994, 
    0.1790445, 0.03406688, 0.07092611, 0.142527, 0.2328318, 0.2193845, 
    0.2062255, 0.1784787, 0.515889, 0.4921881, 0.3307137, 0.2052948, 
    0.1538553, 0.1624093, 0.2042334, 0.1971259, 0.2203535,
  0.264904, 0.2147519, 0.2172283, 0.0823358, 0.2257798, 0.2264192, 
    0.05564352, 0.3257957, 0.3773424, 0.377439, 0.3327971, 0.2650169, 
    0.1980883, 0.2193075, 0.3567296, 0.4048292, 0.3977709, 0.3067371, 
    0.4393747, 0.3453757, 0.4057195, 0.3672602, 0.3890045, 0.3935187, 
    0.3201977, 0.3121429, 0.2920645, 0.2629534, 0.3144774,
  0.4484037, 0.4037579, 0.3929296, 0.2589816, 0.3192397, 0.4945121, 
    0.3216933, 0.5144178, 0.3527269, 0.2085126, 0.2897164, 0.2988308, 
    0.4292028, 0.4931619, 0.412551, 0.4048827, 0.5043832, 0.465446, 
    0.3874624, 0.1867708, 0.1461052, 0.1533938, 0.220691, 0.248274, 
    0.3352388, 0.3507115, 0.3945411, 0.4459842, 0.4913782,
  0.2142965, 0.2183163, 0.229172, 0.2773091, 0.3208411, 0.347277, 0.3317437, 
    0.2639901, 0.2327452, 0.2106003, 0.1970219, 0.2601098, 0.2317804, 
    0.1988752, 0.2340489, 0.2113852, 0.1877836, 0.2680691, 0.2230952, 
    0.2107468, 0.2076551, 0.2370277, 0.2308778, 0.2884638, 0.1367304, 
    0.2589515, 0.2935582, 0.2718047, 0.2313978,
  0.2035644, 0.1056508, 0.06557432, 0.1814452, 0.1892353, 0.1605596, 
    0.1657607, 0.1475503, 0.1514201, 0.06061844, 0.09173754, 0.04293007, 
    0.01160307, 0.0834083, 0.3120416, 0.1503934, 0.1393291, 0.198219, 
    0.1268885, 0.1374338, 0.1830187, 0.2074525, 0.1610337, 0.2932617, 
    0.04380498, 0.1127736, 0.168781, 0.1800227, 0.2729133,
  0.09832899, 0.08601874, 0.009200648, 0.02878515, 0.136488, 0.1019062, 
    0.08017451, 0.07477328, 0.0525089, 0.006975585, 6.859885e-05, 
    -2.797997e-05, 0.01998768, 0.01920374, 0.05665489, 0.1321895, 0.1056323, 
    0.1224538, 0.105954, 0.09145936, 0.1351287, 0.1140938, 0.126851, 
    0.0183282, 0.07229541, 0.1506883, 0.08904053, 0.09001066, 0.1054914,
  0.2522176, 0.003409756, -1.572395e-05, 0.01999306, 0.06867724, 0.01349289, 
    0.01284003, 0.02333356, 0.03644852, 0.002728769, 3.472178e-08, 
    1.885745e-06, 0.03569786, 0.06885891, 0.09797125, 0.1022942, 0.1513575, 
    0.0807905, 0.03847271, 0.03204595, 0.03077559, 0.1237144, 0.2820821, 
    0.003134224, 0.004521598, 0.01194219, 0.02078928, 0.02336811, 0.06473136,
  0.5039541, 0.1506057, -1.029076e-05, 0.01281697, 0.03219111, 0.02702689, 
    0.04103711, 0.05025928, 0.02559096, 0.03568451, 0.03357328, 0.02396274, 
    0.1567573, 0.06939735, 0.02361144, 0.0164862, 0.009870885, 0.005563888, 
    0.0050304, 0.008272119, 0.03946282, 0.2429364, 0.2076157, 0.002619147, 
    3.731795e-05, 2.58365e-07, 0.01285515, 0.01345453, 0.1431471,
  0.312913, 0.1556361, 0.001726113, 0.03176103, 0.04447263, 0.05261573, 
    0.05227298, 0.04572451, 0.03827111, 0.1143334, 0.05331938, 0.04268888, 
    0.06758443, 0.02422835, 0.01346263, 0.009935398, 0.01527791, 0.01133151, 
    0.0145005, 0.02218244, 0.1366945, 0.2583562, 0.04245355, 0.01189204, 
    0.001977619, 0.03583482, 0.02035305, 0.04951117, 0.2698535,
  0.06012012, 0.04642194, 0.01971, 0.1907272, -0.0001082698, 0.01348265, 
    0.03409253, 0.01956175, 0.001028115, 0.01917222, 0.004998902, 0.09769397, 
    0.0412921, 0.09182949, 0.04102174, 0.0526692, 0.07186791, 0.1028374, 
    0.1298007, 0.1403821, 0.1080289, 0.1177636, 0.1926982, 0.06065141, 
    0.01983413, 0.03892398, 0.08278601, 0.1090741, 0.1109455,
  -5.960369e-08, -3.365299e-08, 1.189107e-08, 0.004433276, 0.0002140434, 
    0.06671515, 0.1013705, 0.05280508, 0.1796659, 0.03262333, 0.04532748, 
    0.03645936, 0.01668749, 0.02973239, 0.01151337, 0.01188374, 0.02368032, 
    0.08568136, 0.304768, 0.2224062, 0.06806926, 0.1263138, 0.005242413, 
    0.004056365, 0.01809124, 0.04785673, 0.233187, 0.09024144, -1.604514e-05,
  5.361871e-07, 2.705163e-05, 0.001542608, 4.459048e-08, 3.368445e-07, 
    -4.258673e-07, -0.001697235, 0.3357794, 0.2874787, 0.02978891, 0.1076444, 
    0.08721188, 0.09880796, 0.06116767, 0.09806907, 0.1056275, 0.05386281, 
    0.09425129, 0.4266005, 0.01902384, 7.525743e-05, 0.02287835, 0.01843067, 
    0.06436655, 0.07048076, 0.1123997, 0.1016431, 0.1827758, -0.0003959013,
  0.006549942, 0.0006161877, 0.0001757947, 0.2560772, -4.473471e-05, 
    -3.89459e-06, 0.004462989, -1.135313e-05, 0.004214288, 0.04631897, 
    0.1276112, 0.1612655, 0.3352703, 0.2418141, 0.2769194, 0.2915716, 
    0.3538287, 0.215553, 0.3716429, -0.0001174328, 5.986997e-06, 
    0.0004852809, 0.004662449, 0.06821486, 0.1569563, 0.1909449, 0.1794304, 
    0.1991469, 0.1384758,
  0.1051902, 0.1184919, 0.07883526, 0.05306896, 0.01537156, 0.01499789, 
    0.01001002, 0.09782913, 0.1682309, 0.1317969, 0.07746052, 0.08196771, 
    0.2025552, 0.39669, 0.4303733, 0.4917608, 0.5294113, 0.4731506, 
    0.3219636, 0.04795092, 0.01468243, 0.0126467, 0.0933971, 0.1386153, 
    0.1273385, 0.3420596, 0.3276708, 0.2920473, 0.2451766,
  0.2298088, 0.1304914, 0.1015955, 0.09129215, 0.09921908, 0.109164, 
    0.1693178, 0.1098363, 0.1014762, 0.1664546, 0.1274427, 0.2867154, 
    0.226566, 0.3998848, 0.2897562, 0.4581524, 0.3574969, 0.3093665, 
    0.3714093, 0.09891699, 0.06662678, 0.1751063, 0.2575351, 0.3025481, 
    0.4854323, 0.1766708, 0.4870675, 0.3738873, 0.313845,
  0.5433918, 0.3469954, 0.4661449, 0.3537002, 0.4858413, 0.4065409, 
    0.4397103, 0.4266456, 0.2071058, 0.2878451, 0.3346261, 0.4107318, 
    0.3802437, 0.4370974, 0.4398923, 0.5133104, 0.4763544, 0.3540227, 
    0.3584016, 0.4084597, 0.4617409, 0.5510408, 0.2911499, 0.2970371, 
    0.2404545, 0.3456584, 0.2540343, 0.2651285, 0.6320376,
  0.5350568, 0.5462912, 0.583434, 0.6306361, 0.7154861, 0.7085605, 0.6234736, 
    0.6336843, 0.668659, 0.6855506, 0.6648164, 0.6967342, 0.7127877, 0.77553, 
    0.7463763, 0.7107611, 0.7459949, 0.7263942, 0.739219, 0.7059318, 
    0.6419591, 0.4886131, 0.3306689, 0.3819023, 0.2690057, 0.1516638, 
    0.1588723, 0.3200572, 0.4936145,
  0.1669144, 0.1655347, 0.1641551, 0.1627755, 0.1613958, 0.1600162, 
    0.1586365, 0.1545202, 0.1658204, 0.1771206, 0.1884208, 0.199721, 
    0.2110212, 0.2223215, 0.23868, 0.2346987, 0.2307174, 0.2267361, 
    0.2227548, 0.2187735, 0.2147922, 0.2076001, 0.2016608, 0.1957216, 
    0.1897823, 0.183843, 0.1779037, 0.1719645, 0.1680181,
  0.1991926, 0.0970774, 0.0454226, 0.05824613, 0.0529388, 0.08872264, 
    0.1090032, 0.09137765, 0.04704492, 0.06162827, 0.07925261, 0.1265291, 
    0.2189377, 0.02708572, 0.08458205, 0.1842511, 0.2722981, 0.2520279, 
    0.206919, 0.175493, 0.5223945, 0.5038951, 0.3078599, 0.1912199, 
    0.1784481, 0.1687813, 0.2289607, 0.1958279, 0.2394687,
  0.2305105, 0.1828674, 0.1863339, 0.04681944, 0.1741521, 0.2033857, 
    0.02047978, 0.3144798, 0.3766074, 0.3573065, 0.3003877, 0.2672936, 
    0.1644924, 0.1845272, 0.3603202, 0.4365223, 0.4272286, 0.3434893, 
    0.4378909, 0.3845212, 0.4295046, 0.3751874, 0.3755464, 0.3761266, 
    0.3296522, 0.3514135, 0.3226835, 0.311754, 0.3252171,
  0.4943676, 0.3960618, 0.2989381, 0.2064256, 0.2597201, 0.4170705, 
    0.3431499, 0.4755096, 0.2905428, 0.1499679, 0.2378894, 0.2613809, 
    0.4051644, 0.4702935, 0.4138586, 0.4034925, 0.4943705, 0.489814, 
    0.3299667, 0.1441745, 0.1154434, 0.1191301, 0.1849764, 0.203407, 
    0.3041644, 0.3785102, 0.4332933, 0.5012028, 0.5461061,
  0.1761573, 0.1865018, 0.2308011, 0.2798733, 0.3227066, 0.3605853, 0.320984, 
    0.2478131, 0.2061831, 0.1842037, 0.1564199, 0.2008395, 0.1793117, 
    0.2021437, 0.2000187, 0.1844603, 0.138794, 0.2197994, 0.1791806, 
    0.1807193, 0.1689699, 0.2124443, 0.1930838, 0.2446973, 0.1291866, 
    0.2264082, 0.2453089, 0.2272768, 0.1928605,
  0.1760166, 0.06959321, 0.04623891, 0.1508964, 0.1614457, 0.1467375, 
    0.1383494, 0.0962349, 0.09835112, 0.02904006, 0.05185703, 0.02473672, 
    0.004605642, 0.05300856, 0.2672032, 0.1154549, 0.1062998, 0.1630611, 
    0.1012459, 0.1140966, 0.1709507, 0.1905353, 0.1340365, 0.3007688, 
    0.03179723, 0.08991691, 0.1482324, 0.1506343, 0.2352729,
  0.03463565, 0.03595685, 0.006449138, 0.01582138, 0.1101142, 0.07350634, 
    0.04759935, 0.02552551, 0.02133149, 0.003333496, 2.12786e-05, 
    -0.0001073186, 0.01748753, 0.01046128, 0.03749342, 0.1078682, 0.08374945, 
    0.1246924, 0.09670299, 0.08745724, 0.09157165, 0.06723551, 0.07261077, 
    0.01350496, 0.07650156, 0.1238182, 0.05645115, 0.04326378, 0.04361221,
  0.09513114, 0.005976744, -2.025925e-05, 0.005015734, 0.01979122, 
    0.001659923, 0.004078669, 0.006093587, 0.01120488, 0.0006921653, 
    2.613447e-08, 3.61142e-07, 0.02284807, 0.04377423, 0.07359485, 
    0.08562791, 0.07575336, 0.01865779, 0.01680895, 0.009650003, 0.006193769, 
    0.04292725, 0.1342255, 0.01165822, 0.005434519, 0.01885638, 0.01233881, 
    0.007209619, 0.01919918,
  0.2590993, 0.3098691, 4.91705e-05, 0.02142654, 0.009536176, 0.008369246, 
    0.01610618, 0.02961151, 0.007402054, 0.006151918, 0.02118039, 
    0.004678019, 0.1101277, 0.03584207, 0.00464044, 0.006171862, 0.001249489, 
    0.0005272103, 0.0003561537, 0.0008949746, 0.007482853, 0.08717378, 
    0.1804987, 0.0006542196, 1.300534e-05, 1.191026e-07, -0.001493781, 
    0.00294799, 0.04886281,
  0.1289674, 0.110636, 0.0009867409, 0.0178003, 0.03240852, 0.02072146, 
    0.007281112, 0.01414266, 0.04087321, 0.08183506, 0.02425658, 0.01721786, 
    0.06047924, 0.008737119, 0.002883142, 0.0007036852, 0.003976001, 
    0.003108814, 0.009521088, 0.01656285, 0.07744258, 0.5304207, 0.2444113, 
    0.005280348, 0.0006058508, 0.004563337, 0.00272804, 0.008485198, 0.1132785,
  0.03906582, 0.04248971, 0.01430732, 0.1886144, -6.370498e-05, 0.005368257, 
    0.04683884, 0.00379746, -0.002371148, 0.003259589, 0.002221803, 
    0.02054998, 0.02547322, 0.01964935, 0.01433815, 0.03847037, 0.04782251, 
    0.07804655, 0.08646709, 0.1119182, 0.03554077, 0.05847956, 0.2406133, 
    0.04261932, 0.004545247, 0.01273086, 0.04554122, 0.08492585, 0.09558736,
  -9.96512e-09, 4.81516e-09, 1.14976e-08, 0.002510455, 8.524963e-05, 
    0.05886921, 0.08592348, 0.02209664, 0.1839767, 0.01896423, 0.02183542, 
    0.01519503, 0.003263887, 0.009918935, 0.001462392, 0.001364686, 
    0.004763601, 0.02705298, 0.1637002, 0.4344103, 0.1618768, 0.1092177, 
    0.0003987164, -0.002026169, 0.004025101, 0.01099188, 0.1004976, 
    0.1539869, -1.03969e-05,
  5.203702e-07, 0.0002713088, 0.000812506, -1.136533e-08, 2.81785e-07, 
    -5.767441e-08, -0.00355887, 0.3340833, 0.2805199, 0.02129581, 0.09162666, 
    0.07131649, 0.03996122, 0.01782351, 0.04986637, 0.02088593, 0.01115497, 
    0.03491942, 0.214542, 0.1567736, 2.661165e-05, 0.01761556, 0.01027823, 
    0.01752452, 0.01453722, 0.01983468, 0.03461636, 0.08391668, -0.0005705435,
  0.003050188, 0.0001742054, 6.245795e-05, 0.3081045, -4.92762e-05, 
    -1.015964e-06, 0.003947251, -1.294329e-06, 0.004690778, 0.04286044, 
    0.1277919, 0.148297, 0.4532106, 0.2970029, 0.3191837, 0.4102241, 
    0.3247307, 0.1637403, 0.259106, -0.0003894191, 7.519461e-06, 0.004987303, 
    0.002324592, 0.09717961, 0.1484194, 0.1627858, 0.1114118, 0.1597309, 
    0.1561547,
  0.1044305, 0.09342738, 0.06531081, 0.04053234, 0.007493069, 0.01016303, 
    0.006888575, 0.1039094, 0.1556702, 0.1216527, 0.06948416, 0.07215596, 
    0.3588257, 0.5157757, 0.6273919, 0.6159155, 0.5480469, 0.4487462, 
    0.2837011, 0.05272901, 0.01220903, 0.01279852, 0.09481978, 0.115649, 
    0.1289568, 0.3284652, 0.2873695, 0.2349217, 0.2280821,
  0.2901502, 0.1321411, 0.07571644, 0.08025665, 0.08069553, 0.09103963, 
    0.1510299, 0.0867013, 0.09150901, 0.1592285, 0.1184823, 0.3095692, 
    0.28396, 0.4414086, 0.3428342, 0.4713368, 0.3349817, 0.2902671, 
    0.3735905, 0.08828752, 0.05533379, 0.167563, 0.2449286, 0.2943377, 
    0.5260648, 0.1513526, 0.4382091, 0.333516, 0.3217179,
  0.4472594, 0.2828199, 0.4153054, 0.2687734, 0.4436165, 0.3672518, 
    0.4410955, 0.3964803, 0.1964535, 0.2125514, 0.3010393, 0.3774226, 
    0.3354677, 0.4123048, 0.4265427, 0.4416233, 0.3992445, 0.3008749, 
    0.3441085, 0.3718268, 0.4890906, 0.5432671, 0.2541272, 0.312498, 
    0.4157834, 0.3353632, 0.2281658, 0.302162, 0.5921011,
  0.591798, 0.5839053, 0.5063107, 0.5870223, 0.6761688, 0.697695, 0.7078768, 
    0.6916217, 0.6742439, 0.7194835, 0.6645335, 0.6874467, 0.6964201, 
    0.7273362, 0.7183566, 0.6975753, 0.6965051, 0.7206515, 0.7216002, 
    0.7870595, 0.6740987, 0.5147398, 0.3279789, 0.4646683, 0.3043392, 
    0.1348951, 0.1348283, 0.3331747, 0.515381,
  0.1108561, 0.1108225, 0.1107889, 0.1107552, 0.1107216, 0.110688, 0.1106543, 
    0.1070303, 0.1174268, 0.1278234, 0.13822, 0.1486165, 0.1590131, 
    0.1694097, 0.1690061, 0.1649284, 0.1608507, 0.156773, 0.1526953, 
    0.1486176, 0.1445399, 0.160963, 0.1546778, 0.1483925, 0.1421073, 
    0.135822, 0.1295368, 0.1232515, 0.110883,
  0.2001731, 0.08619949, 0.03696572, 0.05555185, 0.04262707, 0.05743385, 
    0.06677265, 0.0702839, 0.02496833, 0.02817556, 0.04919433, 0.07062161, 
    0.2037442, 0.02233272, 0.1169102, 0.2660596, 0.3203005, 0.3006509, 
    0.201814, 0.203692, 0.5261437, 0.525142, 0.2879987, 0.1836868, 0.2016221, 
    0.2061512, 0.2645864, 0.1787346, 0.2480647,
  0.2051509, 0.1502924, 0.1688177, 0.0281817, 0.1172871, 0.1819094, 
    0.01063641, 0.2848088, 0.3596938, 0.3245889, 0.2735517, 0.2816853, 
    0.1299092, 0.1435241, 0.3719954, 0.4766556, 0.474081, 0.3803201, 
    0.4545414, 0.4328478, 0.4501063, 0.3820135, 0.3727767, 0.355658, 
    0.3445197, 0.3989501, 0.3601801, 0.3816648, 0.3534484,
  0.5370909, 0.4145588, 0.2324531, 0.1568231, 0.2070349, 0.3226931, 
    0.3632751, 0.4465924, 0.226783, 0.1073227, 0.1832193, 0.2249113, 
    0.3659411, 0.4104044, 0.3736618, 0.3936768, 0.4551526, 0.4720212, 
    0.2675048, 0.1089348, 0.09404141, 0.09602602, 0.1537403, 0.1648415, 
    0.2655877, 0.3800154, 0.4316569, 0.5020281, 0.5896512,
  0.1449762, 0.1606137, 0.2150428, 0.2619401, 0.2976743, 0.3253092, 
    0.2852269, 0.2130336, 0.1737953, 0.1520294, 0.115317, 0.1485725, 
    0.1230281, 0.1793226, 0.1567338, 0.1427659, 0.1000281, 0.1823132, 
    0.134454, 0.1373871, 0.1333703, 0.1641914, 0.1421238, 0.2046518, 
    0.09999808, 0.173749, 0.2138569, 0.1915953, 0.1619387,
  0.1411225, 0.04178696, 0.03677573, 0.1127921, 0.1363007, 0.1268879, 
    0.09592238, 0.06424588, 0.07200988, 0.01375942, 0.02900485, 0.01331056, 
    0.002159294, 0.0366481, 0.2131605, 0.08361167, 0.07615757, 0.138101, 
    0.09077215, 0.09424339, 0.1438189, 0.1640669, 0.09881143, 0.2947732, 
    0.02183261, 0.06750114, 0.1184103, 0.107638, 0.1823513,
  0.01214832, 0.0150017, 0.00443182, 0.006086688, 0.07067484, 0.052097, 
    0.02853084, 0.01384006, 0.011824, 0.00206011, 2.835882e-06, 
    -0.0002933553, 0.01312194, 0.006383696, 0.02982102, 0.08249943, 
    0.06690896, 0.1163052, 0.07319288, 0.05581648, 0.05529361, 0.03553473, 
    0.02811733, 0.01098688, 0.07445069, 0.05986066, 0.0296629, 0.02241041, 
    0.01774392,
  0.04169708, 0.01075361, -1.948935e-05, 0.001983957, 0.003914719, 
    0.0003065284, 0.001537727, 0.002281036, 0.004863406, 0.0002788338, 
    2.135289e-08, 1.963628e-07, 0.01615147, 0.03425354, 0.03815935, 
    0.04887173, 0.03634981, 0.005147505, 0.009719891, 0.004412102, 
    0.001741316, 0.01721314, 0.05995807, 0.01288041, 0.003073993, 0.02961954, 
    0.006842197, 0.0028356, 0.0078338,
  0.1212505, 0.1952366, 0.0001104036, 0.02857387, 0.002672064, 0.0024093, 
    0.004725422, 0.0163767, 0.00117777, -0.0009413175, 0.0122797, 
    0.0006308502, 0.0640623, 0.01267816, 0.001054895, 0.006375195, 
    0.0003509989, 0.0001242454, 0.0001394464, 0.000333349, 0.002717976, 
    0.03244642, 0.07448809, 0.0001226006, 4.893382e-06, 7.511177e-08, 
    -0.001312052, 0.001213023, 0.0186867,
  0.04454651, 0.09051886, 0.0005419547, 0.008142446, 0.005711059, 0.00827287, 
    0.001946304, 0.00354776, 0.04574762, 0.06651839, 0.002862484, 
    0.006373552, 0.04003768, 0.003770401, 0.000343708, 3.155721e-05, 
    0.0001263484, 5.304129e-05, 0.0004881379, 0.003818483, 0.0144868, 
    0.2312188, 0.2026387, 0.002015373, 0.0002039254, 0.001224082, 
    0.0005560183, 0.00339611, 0.03353184,
  0.02678169, 0.04017637, 0.009759446, 0.1945756, -3.300063e-05, 
    0.0005057282, 0.05770637, 0.0004867785, -0.003164062, 0.000815886, 
    0.0002891995, 0.005679496, 0.01416815, 0.005983322, 0.002284219, 
    0.0209386, 0.02338506, 0.0537837, 0.05063797, 0.05832805, 0.01131648, 
    0.02290619, 0.2773644, 0.02914439, 0.001256619, 0.003305316, 0.01235251, 
    0.03886537, 0.08144711,
  2.442337e-08, 2.533291e-08, 1.13603e-08, 0.001446091, 2.672951e-05, 
    0.02123261, 0.05198882, 0.002016398, 0.1940384, 0.006150673, 0.006100004, 
    0.005349951, 0.0001745424, 0.004531909, 6.592815e-05, 0.0003706453, 
    0.001648657, 0.008835535, 0.06321931, 0.2376148, 0.04466475, 0.08664532, 
    7.632259e-05, -0.002027027, 0.001027764, 0.002904051, 0.03381321, 
    0.1167053, -2.030391e-06,
  5.089064e-07, 0.0004580657, 0.0006762762, -5.966712e-07, 2.498797e-07, 
    -4.635154e-09, -0.004733284, 0.3118465, 0.2711846, 0.01373539, 0.0551916, 
    0.01994952, 0.01409339, 0.006896717, 0.01666839, 0.006044888, 
    0.002298692, 0.02109169, 0.08545594, 0.1846174, 8.203348e-06, 0.01190136, 
    0.0069914, 0.005316982, 0.003683511, 0.005759561, 0.009423682, 
    0.03351781, -1.672006e-05,
  0.001474074, -4.292053e-05, 1.401801e-05, 0.3203008, -5.505776e-05, 
    -5.264411e-07, 0.004188512, 2.245212e-07, 0.00746179, 0.03390321, 
    0.1279756, 0.1457424, 0.4245593, 0.2990147, 0.3335899, 0.4019518, 
    0.2544823, 0.1053634, 0.1794586, -0.001135851, 6.178871e-06, 0.01040541, 
    0.003673866, 0.1123053, 0.1239834, 0.1303913, 0.07139236, 0.1148444, 
    0.1251278,
  0.08334419, 0.07818894, 0.05457431, 0.03342886, 0.00287068, 0.006457123, 
    0.004502982, 0.09674264, 0.138164, 0.1165442, 0.06095225, 0.06893196, 
    0.4352669, 0.5965083, 0.6810902, 0.6477528, 0.5001624, 0.3574971, 
    0.2327323, 0.05171599, 0.01013074, 0.009675153, 0.08608216, 0.09784344, 
    0.1361002, 0.3258177, 0.237131, 0.1822489, 0.2260424,
  0.2604471, 0.1224637, 0.05595485, 0.06730153, 0.06928779, 0.079948, 
    0.1326649, 0.07164101, 0.0835905, 0.1493247, 0.1099102, 0.3061092, 
    0.2972289, 0.4319865, 0.3734585, 0.4291049, 0.3167311, 0.2710792, 
    0.3456862, 0.07961445, 0.04812994, 0.1567191, 0.2244279, 0.2834865, 
    0.5024458, 0.1434412, 0.3792056, 0.258159, 0.3453201,
  0.391259, 0.2309887, 0.3814916, 0.2402653, 0.3601021, 0.4007002, 0.3709585, 
    0.3526497, 0.1778167, 0.1737784, 0.2564422, 0.3364365, 0.3094171, 
    0.3819727, 0.3365835, 0.3588484, 0.3148456, 0.267729, 0.2989588, 
    0.313668, 0.487098, 0.4995624, 0.2386864, 0.2786156, 0.5056359, 
    0.3014525, 0.1984165, 0.2745702, 0.5177732,
  0.6246467, 0.5164756, 0.4076349, 0.4828942, 0.5608009, 0.6050645, 
    0.6360205, 0.5908799, 0.5880532, 0.64588, 0.5887482, 0.6556622, 
    0.6242166, 0.6435945, 0.6541213, 0.6375631, 0.61834, 0.6285819, 
    0.6409562, 0.750156, 0.6335875, 0.4642454, 0.4013447, 0.4964092, 
    0.2610937, 0.1310098, 0.098842, 0.3140017, 0.5093465,
  0.04760742, 0.04655469, 0.04550196, 0.04444923, 0.0433965, 0.04234376, 
    0.04129103, 0.06029951, 0.06972641, 0.07915331, 0.08858021, 0.09800711, 
    0.107434, 0.1168609, 0.1187813, 0.1168691, 0.1149569, 0.1130447, 
    0.1111325, 0.1092203, 0.107308, 0.1219414, 0.1154794, 0.1090175, 
    0.1025555, 0.09609354, 0.08963158, 0.08316962, 0.04844961,
  0.1727674, 0.07179354, 0.02256852, 0.03738889, 0.03738884, 0.02765396, 
    0.03114915, 0.03678808, 0.001867832, 0.002353607, 0.009859001, 
    0.04470035, 0.1815989, 0.01690336, 0.1558236, 0.3736518, 0.3446867, 
    0.3270884, 0.1748076, 0.2268572, 0.5442013, 0.5579773, 0.2455844, 
    0.1553337, 0.2285811, 0.2775171, 0.2697144, 0.1634174, 0.2338951,
  0.1923821, 0.1189573, 0.1598729, 0.01915316, 0.08005162, 0.1573056, 
    0.004417872, 0.223493, 0.3271778, 0.2691083, 0.2333134, 0.2884416, 
    0.101392, 0.105182, 0.4040505, 0.4939105, 0.4487351, 0.3730195, 
    0.4052809, 0.4183916, 0.4460081, 0.3812687, 0.3692002, 0.3144384, 
    0.3297305, 0.4137067, 0.3970802, 0.4206944, 0.3520628,
  0.5222409, 0.3925931, 0.1746949, 0.1102031, 0.1508899, 0.2438462, 
    0.3431291, 0.3875423, 0.1744316, 0.07084264, 0.1374541, 0.185793, 
    0.315751, 0.3391786, 0.3009919, 0.3163339, 0.3808302, 0.4123475, 
    0.2069501, 0.07932541, 0.07713483, 0.07764249, 0.1185792, 0.1300843, 
    0.2388712, 0.3374511, 0.3948419, 0.4522554, 0.5346105,
  0.1161774, 0.1321357, 0.1772323, 0.2242741, 0.2552856, 0.2609293, 
    0.2369116, 0.1623514, 0.1367585, 0.113188, 0.07993889, 0.09884556, 
    0.07787803, 0.126448, 0.1266492, 0.1046122, 0.07124122, 0.1420455, 
    0.09345412, 0.09541808, 0.1002352, 0.1165615, 0.09741271, 0.1719645, 
    0.07692222, 0.1333703, 0.1748984, 0.1465915, 0.1278862,
  0.1014465, 0.02482891, 0.02993742, 0.08181251, 0.0957312, 0.08743261, 
    0.05909777, 0.0405345, 0.05217354, 0.006367447, 0.01237616, 0.006674326, 
    0.0009506276, 0.02420766, 0.1586221, 0.06293705, 0.05627995, 0.1087013, 
    0.07518202, 0.06897295, 0.1163011, 0.1289276, 0.06312979, 0.2699706, 
    0.01600433, 0.050381, 0.07650701, 0.07042093, 0.1306399,
  0.006889455, 0.008828293, 0.002678578, 0.002368881, 0.039346, 0.03204978, 
    0.01549373, 0.008380516, 0.007988815, 0.001469209, 2.193448e-06, 
    -0.0003891652, 0.008738504, 0.003804246, 0.02045051, 0.05725972, 
    0.05141278, 0.08444662, 0.04849761, 0.03015346, 0.03044897, 0.0212718, 
    0.01483087, 0.006149057, 0.06658089, 0.03192717, 0.01570995, 0.01295401, 
    0.009794901,
  0.02325844, 0.01124713, -1.462708e-05, 0.001173011, 9.206642e-05, 
    0.0001390124, 0.0004692086, 0.001164375, 0.00271148, 0.0001651129, 
    1.846606e-08, -6.596956e-09, 0.009645741, 0.01314745, 0.01640299, 
    0.02096741, 0.01242397, 0.002176554, 0.005123854, 0.002107302, 
    0.0008522343, 0.008760316, 0.03221013, 0.00827591, 0.001083293, 
    0.0409596, 0.003734084, 0.001455753, 0.004245515,
  0.06521168, 0.08915354, 4.542888e-05, 0.02923284, 0.0007522634, 
    0.001003952, 0.001413006, 0.00705268, 0.0002459979, -0.001613076, 
    0.009255962, 0.0002298133, 0.03216607, 0.004518795, 0.0003038624, 
    0.004729239, 0.0002018295, 6.991842e-05, 7.425897e-05, 0.0001876591, 
    0.001415148, 0.01584946, 0.03916603, 0.0003769783, 1.360823e-06, 
    1.084072e-07, -0.001174543, 0.000666945, 0.00975095,
  0.02281524, 0.0833884, 0.0005366516, 0.003318435, 0.0008313, 0.003533709, 
    0.00102124, 0.001409927, 0.04100575, 0.06460222, 0.0005554993, 
    0.003872393, 0.02115658, 0.001860874, 7.956514e-05, 9.945596e-06, 
    3.025291e-05, 1.198986e-05, 4.405449e-05, 0.0003612236, 0.004131515, 
    0.1014186, 0.1006355, 0.0007915612, 0.0001009864, 0.0006113234, 
    0.0002997129, 0.001919175, 0.016041,
  0.02196761, 0.03915966, 0.00402688, 0.1842604, -1.534118e-05, 5.021522e-05, 
    0.04814869, 0.0001533575, -0.00186998, 0.0004220909, 2.060795e-05, 
    0.002717409, 0.006633426, 0.0026012, 0.0003262922, 0.009076477, 
    0.01005793, 0.03747315, 0.02421242, 0.02451092, 0.004564741, 0.01020115, 
    0.2337965, 0.02640729, 0.0005776642, 0.001785747, 0.003460095, 
    0.01563095, 0.06253918,
  3.985416e-08, 2.040045e-08, 1.134925e-08, 0.0006299394, 7.068177e-06, 
    0.003857469, 0.02023599, -0.0002365188, 0.1888149, 0.001271667, 
    0.002020305, 0.002075056, 1.571756e-05, 0.002014899, 2.652108e-05, 
    0.0001810172, 0.0008515861, 0.00430989, 0.0259752, 0.1267964, 0.0140252, 
    0.07179363, 3.151746e-05, -0.001509553, 0.0003270385, 0.001335463, 
    0.0145475, 0.06570319, -4.920616e-07,
  5.004248e-07, 0.0003180925, 0.0006973757, -8.021668e-07, 2.298456e-07, 
    -9.108995e-10, -0.004120102, 0.2862983, 0.2511468, 0.008715521, 
    0.02893687, 0.006798012, 0.004378402, 0.003075954, 0.008379636, 
    0.002973981, 0.001127942, 0.01080406, 0.04090425, 0.1295625, 1.93018e-06, 
    0.00880964, 0.004918857, 0.002741985, 0.001717923, 0.002834075, 
    0.00471219, 0.01493827, 8.651429e-05,
  0.0009745386, -8.706575e-05, -1.119181e-05, 0.3085289, -4.688802e-05, 
    -6.649836e-08, 0.003817281, 3.814663e-07, 0.004960208, 0.02514672, 
    0.1171751, 0.1605994, 0.358756, 0.2412845, 0.2859637, 0.2855253, 
    0.1547755, 0.05200263, 0.1202179, -0.001643494, 4.493314e-06, 0.01204064, 
    0.00266272, 0.1217853, 0.07350508, 0.07642931, 0.03886394, 0.0762932, 
    0.1249058,
  0.06320435, 0.06617695, 0.03850018, 0.02463079, 0.001108009, 0.003253283, 
    0.002366473, 0.08678694, 0.1177255, 0.1122372, 0.05257526, 0.06753496, 
    0.4751717, 0.5921718, 0.6232122, 0.6164401, 0.4463802, 0.2877155, 
    0.1843013, 0.04752526, 0.008183794, 0.005685589, 0.07926781, 0.08370094, 
    0.1325304, 0.3352394, 0.1901177, 0.141954, 0.199104,
  0.2475792, 0.1089282, 0.03792636, 0.05228264, 0.05648272, 0.07101478, 
    0.1119483, 0.05624742, 0.07714245, 0.1415606, 0.09645551, 0.2869577, 
    0.2879306, 0.383833, 0.3694348, 0.3648262, 0.2905518, 0.2461495, 0.29151, 
    0.07088336, 0.03775242, 0.1448444, 0.210186, 0.2680022, 0.4357271, 
    0.1436172, 0.3224477, 0.2072603, 0.3006037,
  0.3596987, 0.1817611, 0.3297832, 0.1988922, 0.2932502, 0.3752196, 
    0.3068594, 0.2963172, 0.1574427, 0.1483972, 0.2235761, 0.2995836, 
    0.2763288, 0.350825, 0.27524, 0.305734, 0.2691799, 0.2555608, 0.2675925, 
    0.2669117, 0.4722132, 0.4677132, 0.2200537, 0.2440968, 0.4686035, 
    0.2594724, 0.1790685, 0.2636447, 0.4660295,
  0.596349, 0.4463083, 0.3339185, 0.4119416, 0.4503836, 0.5090347, 0.5625702, 
    0.5072039, 0.5034599, 0.5481517, 0.5016363, 0.5489542, 0.5239334, 
    0.551071, 0.5554806, 0.5527325, 0.5365319, 0.5571777, 0.5707395, 
    0.6594322, 0.5761338, 0.3618714, 0.3781179, 0.4568744, 0.2135441, 
    0.1094791, 0.07747231, 0.2722478, 0.4976467,
  0.02233258, 0.02051677, 0.01870096, 0.01688515, 0.01506934, 0.01325352, 
    0.01143771, 0.0191949, 0.02499907, 0.03080324, 0.0366074, 0.04241157, 
    0.04821574, 0.05401991, 0.06361858, 0.06506033, 0.06650209, 0.06794384, 
    0.0693856, 0.07082735, 0.07226911, 0.07162088, 0.06619077, 0.06076066, 
    0.05533055, 0.04990044, 0.04447033, 0.03904022, 0.02378523,
  0.1480693, 0.04568762, 0.01709957, 0.04831766, 0.03025722, 0.01055329, 
    0.02078542, 0.01458847, 0.007215346, 0.005496575, 0.008780966, 
    0.02007752, 0.1110888, 0.009563995, 0.2305155, 0.3819325, 0.2799461, 
    0.3649918, 0.1677531, 0.2792771, 0.5395105, 0.5764391, 0.2248647, 
    0.1407673, 0.240117, 0.3548111, 0.2548494, 0.1424595, 0.2113792,
  0.1783888, 0.08854515, 0.1532504, 0.0148938, 0.06425972, 0.1325956, 
    0.00328832, 0.1622808, 0.2872117, 0.2065715, 0.1964354, 0.2695674, 
    0.0817939, 0.08860675, 0.410705, 0.4663979, 0.4131526, 0.3482423, 
    0.368228, 0.3927431, 0.4071431, 0.3701551, 0.3688717, 0.2672574, 
    0.2996674, 0.4256954, 0.4190639, 0.3871403, 0.307302,
  0.4318958, 0.3352944, 0.1347542, 0.07579962, 0.1107277, 0.1878924, 
    0.313291, 0.3287998, 0.1378261, 0.04762282, 0.1019997, 0.1439084, 
    0.2595972, 0.265954, 0.220642, 0.2335718, 0.2968971, 0.3410436, 
    0.1604489, 0.06058076, 0.06192136, 0.06031259, 0.09267785, 0.09842294, 
    0.2004822, 0.278003, 0.3525651, 0.3889139, 0.4461229,
  0.09094816, 0.1034199, 0.1345074, 0.1783549, 0.2148701, 0.205249, 
    0.1904524, 0.1213698, 0.1048776, 0.08161899, 0.05307452, 0.06217147, 
    0.04568473, 0.0769539, 0.09650169, 0.07513168, 0.05041445, 0.09430967, 
    0.06484608, 0.06421529, 0.0708008, 0.07840903, 0.06277777, 0.1442638, 
    0.05326406, 0.08954606, 0.131019, 0.1105415, 0.09597863,
  0.06820571, 0.01402236, 0.02167108, 0.04990026, 0.05409269, 0.05057151, 
    0.03474997, 0.02449002, 0.03312075, 0.003352981, 0.006205287, 
    0.003797146, 0.0005526387, 0.01480574, 0.1177424, 0.04193908, 0.03588378, 
    0.07874103, 0.05647686, 0.04422852, 0.08677211, 0.09042913, 0.03772621, 
    0.238676, 0.01071967, 0.03420477, 0.04785584, 0.0459485, 0.08752099,
  0.004790072, 0.006148955, 0.001399764, 0.001280245, 0.02017893, 0.01569152, 
    0.008974365, 0.00567178, 0.006025127, 0.001138247, 4.044637e-07, 
    -0.0002410008, 0.005374178, 0.002258714, 0.01192018, 0.03717443, 
    0.03196427, 0.05212223, 0.02863397, 0.01442373, 0.01465204, 0.01214921, 
    0.009952216, 0.004040518, 0.05610979, 0.01463362, 0.008491733, 
    0.00668037, 0.006686809,
  0.01537587, 0.009907913, -1.050003e-05, 0.0008160658, -0.0006577286, 
    8.516066e-05, 0.0002140369, 0.0007279392, 0.001771523, 0.0001149517, 
    1.827072e-08, -2.606411e-06, 0.004336197, 0.00612031, 0.006757148, 
    0.007123712, 0.005289691, 0.001394005, 0.002570185, 0.0009682403, 
    0.000525643, 0.005417133, 0.02145027, 0.006518778, 0.0005426791, 
    0.0373898, 0.001979597, 0.0008957664, 0.002737005,
  0.04210608, 0.04134148, 1.454383e-05, 0.02684899, 0.0004062379, 
    0.0003124615, 0.000650019, 0.00264273, 0.0001191258, -0.0008169132, 
    0.006174917, 0.0001421049, 0.01295679, 0.001608441, 0.000133176, 
    0.00262072, 0.0001362155, 4.714409e-05, 4.806202e-05, 0.0001255922, 
    0.0008975922, 0.009673972, 0.02481888, 0.0002115724, 5.341762e-07, 
    4.781765e-08, -0.0006920893, 0.0004342462, 0.006220461,
  0.01469991, 0.06955329, 0.0003869005, 0.001474899, 0.0003655872, 
    0.001663592, 0.0006587066, 0.0008115473, 0.03072764, 0.06353644, 
    0.0002845676, 0.002113604, 0.009220053, 0.0008981776, 4.053415e-05, 
    5.409167e-06, 1.49552e-05, 5.293353e-06, 1.953268e-05, 0.00013362, 
    0.002173421, 0.05685586, 0.06709454, 0.00114111, -8.113075e-05, 
    0.0003842089, 0.0001958824, 0.001278318, 0.01002846,
  0.01244764, 0.02807987, 0.001519681, 0.1610917, -6.692819e-06, 
    2.276837e-05, 0.0285456, 9.491923e-05, -0.000752208, 0.0002618911, 
    -6.815163e-06, 0.001678492, 0.002734937, 0.001242516, 9.310543e-05, 
    0.003574374, 0.00406771, 0.01853339, 0.01070436, 0.01019011, 0.002066627, 
    0.004555497, 0.1888525, 0.02854284, 0.0002119369, 0.0009054839, 
    0.001135064, 0.006406242, 0.04043174,
  4.476358e-08, 2.709732e-08, 1.135962e-08, 0.0003394521, 9.829594e-07, 
    0.001515086, 0.004708712, -0.0002184821, 0.1564614, 0.0002430988, 
    0.0008436621, 0.0008208753, 9.906635e-06, 0.0008838734, 1.421893e-05, 
    0.0001086524, 0.000540034, 0.002400148, 0.01446381, 0.07526652, 
    0.007130017, 0.05957913, 1.645945e-05, -0.001097008, 0.0001536733, 
    0.0008229515, 0.008458695, 0.03499697, -1.441466e-07,
  4.939545e-07, 0.0001106947, 0.0002644013, -1.376532e-06, 2.171758e-07, 
    -7.866158e-10, -0.005076933, 0.2616943, 0.2242774, 0.004379349, 
    0.0115218, 0.003067207, 0.001793504, 0.001029425, 0.004112164, 
    0.001952443, 0.0007306485, 0.004496328, 0.02473536, 0.1040661, 
    -3.810722e-07, 0.005755594, 0.002737481, 0.001761346, 0.001100941, 
    0.001778165, 0.002990703, 0.00886978, -1.249624e-05,
  0.0006544128, -0.0001092192, -2.95807e-05, 0.2802989, -4.496014e-05, 
    -1.167107e-07, 0.0033732, 4.246133e-07, 0.002534661, 0.01803937, 
    0.1064821, 0.1413164, 0.2824419, 0.1814073, 0.203346, 0.181789, 
    0.07858604, 0.02431177, 0.08151628, -0.00203121, 3.465607e-06, 
    0.01024788, 0.003837867, 0.1075414, 0.03649178, 0.03812686, 0.01753441, 
    0.04045137, 0.1070073,
  0.03970408, 0.05220726, 0.02491669, 0.01531539, 0.0005565647, 0.001534623, 
    0.001280787, 0.08022177, 0.09993746, 0.1047753, 0.04732522, 0.05823641, 
    0.4459142, 0.5474033, 0.5383565, 0.5446771, 0.3950942, 0.2173713, 
    0.1303583, 0.04431482, 0.006026482, 0.003213061, 0.07271868, 0.06933652, 
    0.1167085, 0.3139957, 0.1392563, 0.09803744, 0.1329639,
  0.2058872, 0.0931377, 0.02547104, 0.0350301, 0.04516237, 0.05805804, 
    0.0923619, 0.04063128, 0.07174947, 0.1266462, 0.0806064, 0.2520703, 
    0.2703268, 0.3177288, 0.308477, 0.2954728, 0.2557121, 0.2089472, 
    0.2228081, 0.05963737, 0.02897917, 0.1361559, 0.183841, 0.2407137, 
    0.3589989, 0.1367209, 0.2268885, 0.1506495, 0.2449455,
  0.2946722, 0.1414284, 0.2791001, 0.1517745, 0.2350268, 0.3253927, 
    0.2499975, 0.2502376, 0.1357107, 0.1250174, 0.1878335, 0.2579297, 
    0.2398905, 0.3375527, 0.2284513, 0.2699962, 0.2241022, 0.2364122, 
    0.2404696, 0.240822, 0.4066046, 0.4376578, 0.1968383, 0.2155943, 
    0.4256227, 0.2201231, 0.1755695, 0.2455922, 0.4193097,
  0.5632377, 0.3899843, 0.2813371, 0.3531522, 0.3572773, 0.4201474, 
    0.4731287, 0.418901, 0.416862, 0.4408188, 0.4010752, 0.3990768, 
    0.3686198, 0.3870756, 0.3995532, 0.4039741, 0.4200966, 0.4540919, 
    0.480267, 0.5389861, 0.5011486, 0.2864101, 0.3314529, 0.4193898, 
    0.1794348, 0.08303151, 0.06034918, 0.2359916, 0.4575048,
  0.01063811, 0.01023984, 0.009841574, 0.009443304, 0.009045033, 0.008646763, 
    0.008248492, 0.0150442, 0.01870375, 0.02236331, 0.02602287, 0.02968242, 
    0.03334198, 0.03700154, 0.04372801, 0.04408812, 0.04444823, 0.04480834, 
    0.04516844, 0.04552855, 0.04588866, 0.03377788, 0.03015648, 0.02653509, 
    0.02291369, 0.0192923, 0.01567091, 0.01204951, 0.01095673,
  0.0685776, 0.03365948, 0.03529307, 0.05073692, 0.02655786, 0.01763459, 
    0.01757267, 0.003371959, 0.007660978, 0.006642671, 0.004338789, 
    0.01525102, 0.07803261, 0.007341032, 0.3144997, 0.2942623, 0.2507063, 
    0.3845112, 0.1531827, 0.3419797, 0.5467981, 0.6085024, 0.2151739, 
    0.1334001, 0.2269424, 0.343783, 0.2616015, 0.1074552, 0.1776232,
  0.1453911, 0.07336332, 0.1370049, 0.01104783, 0.04420181, 0.1079429, 
    0.002627889, 0.1289995, 0.2330031, 0.1692759, 0.1771321, 0.2491104, 
    0.07017951, 0.07345012, 0.3887235, 0.4313931, 0.3838905, 0.3104842, 
    0.3478841, 0.355608, 0.3616235, 0.3497702, 0.3571143, 0.2383453, 
    0.2726984, 0.4083802, 0.39193, 0.3261866, 0.2499074,
  0.3533099, 0.2766253, 0.1132541, 0.05854423, 0.0844055, 0.1570902, 
    0.2835306, 0.288835, 0.1156092, 0.03581133, 0.07974664, 0.1189092, 
    0.212593, 0.2148911, 0.1690115, 0.179772, 0.2484957, 0.2865223, 
    0.1303881, 0.04829337, 0.05089535, 0.05113892, 0.0762977, 0.07937568, 
    0.1689465, 0.2411704, 0.3156719, 0.3382116, 0.3750574,
  0.07333597, 0.08459486, 0.1059794, 0.1512566, 0.1911708, 0.1708034, 
    0.1607268, 0.09578641, 0.08560072, 0.06229798, 0.0391801, 0.04356523, 
    0.02860809, 0.05143378, 0.06711903, 0.05041549, 0.03602552, 0.06664554, 
    0.04906506, 0.04674245, 0.05311488, 0.05665337, 0.0447449, 0.1304765, 
    0.03964802, 0.06347362, 0.1006362, 0.08865274, 0.07632779,
  0.04577911, 0.009352478, 0.0152076, 0.0313923, 0.03220801, 0.03146588, 
    0.0212157, 0.0148584, 0.02196472, 0.002156547, 0.004091572, 0.002528024, 
    0.0004177501, 0.009000385, 0.091985, 0.02783842, 0.02261043, 0.05509806, 
    0.0414027, 0.02837147, 0.0660589, 0.06184588, 0.02358034, 0.2139087, 
    0.007604538, 0.02302649, 0.03126341, 0.03042362, 0.06061475,
  0.003731713, 0.004818494, 0.0008029871, 0.000902163, 0.01223994, 
    0.008676732, 0.005961423, 0.004295428, 0.00492104, 0.000939401, 
    2.884373e-07, -7.864712e-05, 0.004110755, 0.001473021, 0.007486301, 
    0.02199852, 0.0187063, 0.02756929, 0.01662592, 0.008378856, 0.007991253, 
    0.007397974, 0.007655285, 0.003335358, 0.04538146, 0.008098693, 
    0.004558168, 0.004356289, 0.00518816,
  0.01150695, 0.007959883, -8.25471e-06, 0.0006204033, -0.0005525891, 
    6.165601e-05, 0.0001327883, 0.0005258259, 0.001312634, 8.922053e-05, 
    1.724239e-08, -4.106908e-06, 0.002120709, 0.003621121, 0.003514047, 
    0.003469129, 0.002937497, 0.001040403, 0.001445651, 0.0006247612, 
    0.0003766025, 0.003875189, 0.01617117, 0.00576583, 0.0003280504, 
    0.03114097, 0.001030611, 0.0006362464, 0.002008819,
  0.0309848, 0.0241627, 4.890734e-06, 0.02153921, 0.0002822174, 0.0001447032, 
    0.0004192307, 0.001017084, 7.993425e-05, -0.000332007, 0.003754832, 
    0.000102664, 0.005962491, 0.0007728665, 7.992303e-05, 0.001232784, 
    0.0001033251, 3.5883e-05, 3.558178e-05, 9.520812e-05, 0.0006585199, 
    0.006885611, 0.01814669, 0.0006856791, 5.640245e-07, 4.488229e-08, 
    -0.0004054447, 0.0003220615, 0.004556818,
  0.01090349, 0.06518649, 0.0002380143, 0.0007529648, 0.0002359652, 
    0.0008920989, 0.0004869803, 0.0005730282, 0.02772353, 0.06506225, 
    0.0001919628, 0.0009889537, 0.004430759, 0.0004579794, 2.797481e-05, 
    3.862719e-06, 9.801238e-06, 3.297057e-06, 1.190633e-05, 7.989553e-05, 
    0.001452946, 0.0388375, 0.05082269, 0.00363343, 0.0006532529, 
    0.0002795486, 0.0001459969, 0.0009594553, 0.007246311,
  0.007753349, 0.01664046, 0.0007137058, 0.1310963, -3.236243e-06, 
    1.484884e-05, 0.01627569, 6.949668e-05, -0.0003991756, 0.0001894608, 
    -6.233267e-07, 0.001204009, 0.001246091, 0.0006907419, 6.094882e-05, 
    0.00158324, 0.001720001, 0.007857597, 0.004838623, 0.004381154, 
    0.001050776, 0.002084349, 0.1541378, 0.03110302, 9.573216e-05, 
    0.0004506756, 0.0004790449, 0.002762234, 0.02273968,
  4.284535e-08, 2.689331e-08, 1.139205e-08, 0.0002149907, 1.172872e-07, 
    0.0009012822, 0.001869724, -0.0001155095, 0.1154297, 5.821451e-05, 
    0.0004404864, 0.0004081273, 1.050734e-05, 0.0004870563, 1.002983e-05, 
    7.658733e-05, 0.0003816066, 0.001698704, 0.009886676, 0.05052954, 
    0.00481644, 0.05057077, 1.035816e-05, -0.0009541545, 9.892012e-05, 
    0.0005898039, 0.0058473, 0.02066166, -6.155729e-08,
  4.889725e-07, 5.536988e-05, 0.0001720456, -1.048933e-06, 2.078233e-07, 
    -7.539471e-10, -0.005199101, 0.241577, 0.1995535, 0.002260728, 
    0.00575295, 0.001960081, 0.001020856, 0.0005754032, 0.002607882, 
    0.001447491, 0.0005357093, 0.002469018, 0.01694575, 0.08805149, 
    -1.222886e-06, 0.004727012, 0.005469231, 0.001291215, 0.0008076284, 
    0.001283641, 0.002176966, 0.006295117, -6.958714e-05,
  0.0006173056, -0.0001285845, -3.019939e-05, 0.2502548, -4.610783e-05, 
    -8.999824e-08, 0.002858645, 4.312876e-07, 0.001465371, 0.01250329, 
    0.09625222, 0.1133448, 0.2049797, 0.1348378, 0.1466893, 0.1157125, 
    0.03921383, 0.01215059, 0.05860432, -0.002245025, 3.289813e-06, 
    0.008310097, 0.005423734, 0.08918819, 0.02250625, 0.02159073, 
    0.009597061, 0.02333977, 0.08616692,
  0.02654123, 0.04450247, 0.01943418, 0.01032454, 0.0003395059, 0.000876096, 
    0.0008461814, 0.07554197, 0.08854379, 0.09684871, 0.049932, 0.04816052, 
    0.3915281, 0.4777235, 0.4379341, 0.4248265, 0.3142969, 0.1554169, 
    0.08879808, 0.04249121, 0.004914404, 0.002017687, 0.06429003, 0.06490158, 
    0.09900307, 0.2663591, 0.09929916, 0.06652847, 0.09004097,
  0.1627425, 0.08153629, 0.01899467, 0.02705412, 0.03826711, 0.04896627, 
    0.07953948, 0.03140325, 0.07758224, 0.112053, 0.07258362, 0.2252671, 
    0.2556394, 0.2497867, 0.2333108, 0.2073646, 0.2201166, 0.1818326, 
    0.1682755, 0.05070405, 0.02191707, 0.1311401, 0.1528277, 0.2136314, 
    0.2866347, 0.1277377, 0.1554152, 0.1030515, 0.2037206,
  0.2129025, 0.1075959, 0.235601, 0.1094204, 0.1966494, 0.2830842, 0.2099369, 
    0.2118447, 0.1164313, 0.1021969, 0.160058, 0.2253194, 0.2096263, 
    0.3083578, 0.2007518, 0.2285159, 0.1912158, 0.2158466, 0.2278038, 
    0.2387851, 0.3379616, 0.4201937, 0.1715996, 0.1947775, 0.3689676, 
    0.1930539, 0.1767898, 0.2210677, 0.3552095,
  0.5280558, 0.3523086, 0.2367244, 0.2961058, 0.2954976, 0.3518423, 
    0.4013979, 0.3690097, 0.3487965, 0.3521875, 0.3236125, 0.3128492, 
    0.2833363, 0.2878568, 0.2973697, 0.3094811, 0.33084, 0.3671616, 
    0.3906819, 0.4565267, 0.4326625, 0.2401776, 0.2942113, 0.3832873, 
    0.1561508, 0.0714043, 0.04744088, 0.2110931, 0.4094348,
  0.00733426, 0.006980754, 0.006627249, 0.006273742, 0.005920236, 
    0.005566731, 0.005213225, 0.007330619, 0.00993062, 0.01253062, 
    0.01513062, 0.01773063, 0.02033063, 0.02293063, 0.03112542, 0.03186237, 
    0.03259933, 0.03333628, 0.03407323, 0.03481019, 0.03554714, 0.02623771, 
    0.02325426, 0.02027082, 0.01728737, 0.01430392, 0.01132047, 0.008337021, 
    0.007617065,
  0.04083214, 0.02809243, 0.04436368, 0.02329945, 0.01594151, 0.009243914, 
    0.01597996, 0.003213633, 0.01182834, 0.006126458, 0.001271446, 0.0124461, 
    0.0585412, 0.006344193, 0.3528533, 0.1841285, 0.2079494, 0.452164, 
    0.1911647, 0.3777639, 0.5421022, 0.6307691, 0.2228208, 0.1303445, 
    0.230073, 0.3218163, 0.2558647, 0.1090071, 0.1207478,
  0.1306965, 0.07188068, 0.1188306, 0.009585799, 0.02044882, 0.09728295, 
    0.002623167, 0.1223703, 0.2163673, 0.1513413, 0.1691989, 0.2450452, 
    0.06482954, 0.0672929, 0.366879, 0.4114579, 0.3575917, 0.2971813, 
    0.3220024, 0.3360547, 0.3372186, 0.3380627, 0.3320657, 0.2123919, 
    0.2632543, 0.3845601, 0.3527799, 0.2967206, 0.2225017,
  0.3177933, 0.2501245, 0.1021746, 0.05076647, 0.07235745, 0.1427594, 
    0.2592134, 0.272935, 0.1051217, 0.03064362, 0.06781013, 0.105301, 
    0.1824608, 0.1860515, 0.1415824, 0.1503357, 0.2170407, 0.2497145, 
    0.1122721, 0.04169594, 0.04379959, 0.04541976, 0.06685487, 0.06955259, 
    0.1570196, 0.2266011, 0.2987587, 0.3108796, 0.3428846,
  0.06342666, 0.07143039, 0.09005723, 0.1294486, 0.1667792, 0.1509098, 
    0.1396167, 0.08230847, 0.07580099, 0.05321345, 0.03306633, 0.0351643, 
    0.02182458, 0.03818284, 0.04868643, 0.03727719, 0.02762631, 0.05030934, 
    0.03538148, 0.03647152, 0.04428399, 0.04647929, 0.03683378, 0.1530848, 
    0.03268237, 0.05114862, 0.08556705, 0.07649036, 0.06741507,
  0.0341128, 0.007685425, 0.01015493, 0.02272481, 0.02236016, 0.02239148, 
    0.01582749, 0.0108664, 0.01649771, 0.001733895, 0.003229324, 0.002019839, 
    0.0003633391, 0.006311744, 0.08518238, 0.01940206, 0.01593945, 0.0403452, 
    0.03166955, 0.02106948, 0.0519184, 0.04548675, 0.01756234, 0.2108804, 
    0.005532339, 0.01639341, 0.0232323, 0.02292107, 0.04473496,
  0.003188174, 0.004122047, 0.0005144541, 0.0007409157, 0.007369223, 
    0.005523153, 0.004462652, 0.003655186, 0.004315845, 0.000809208, 
    1.258496e-07, -9.76333e-05, 0.005297273, 0.001125479, 0.005336177, 
    0.01360928, 0.01065912, 0.01533302, 0.01022094, 0.00573923, 0.005201821, 
    0.005524285, 0.006434494, 0.002958949, 0.04571974, 0.005096637, 
    0.00313037, 0.003355903, 0.004410833,
  0.00963827, 0.006650776, -7.982179e-06, 0.0005391793, -0.0005848292, 
    5.198288e-05, 0.0001062058, 0.0004409543, 0.001107481, 7.699768e-05, 
    1.657208e-08, -2.190772e-06, 0.001392965, 0.00255253, 0.002342586, 
    0.002312632, 0.002085455, 0.0008501743, 0.001018928, 0.0004838544, 
    0.000309117, 0.00316278, 0.01362213, 0.005260725, 0.0002263398, 
    0.03342439, 0.0006814856, 0.0005207935, 0.001668339,
  0.02550407, 0.01688468, 4.191618e-06, 0.01852055, 0.0002254384, 
    0.0001018941, 0.0003470407, 0.0005639876, 6.474375e-05, -0.0002660174, 
    0.002652348, 8.610411e-05, 0.003757665, 0.0005416843, 6.047767e-05, 
    0.0007233766, 8.989252e-05, 3.078873e-05, 3.050447e-05, 8.170409e-05, 
    0.0005515274, 0.005627622, 0.01490692, 0.007873468, 1.724817e-07, 
    5.246056e-08, -0.0003410441, 0.000271001, 0.003781035,
  0.009002563, 0.1162284, 0.002735275, 0.0004734837, 0.000181924, 
    0.0006295225, 0.0003698037, 0.0004566998, 0.0433401, 0.09966969, 
    0.0001534557, 0.0005996805, 0.002889614, 0.0002958033, 2.299863e-05, 
    3.337385e-06, 8.112683e-06, 2.750699e-06, 9.719267e-06, 6.046926e-05, 
    0.001142446, 0.0304582, 0.04232103, 0.02427844, 0.02283988, 0.0002321277, 
    0.0001234936, 0.0008039342, 0.005861878,
  0.03080849, 0.02327426, 0.0007905925, 0.121053, -1.984797e-06, 
    1.189854e-05, 0.01803022, 5.153758e-05, -0.00167738, 0.0001572678, 
    4.397933e-06, 0.0009691581, 0.0008190579, 0.0005016073, 4.957918e-05, 
    0.0009925682, 0.001022861, 0.004408264, 0.002905616, 0.002772106, 
    0.0006821995, 0.001304265, 0.219196, 0.04076367, 6.381297e-05, 
    0.0003042124, 0.0003415616, 0.001709793, 0.03477518,
  4.160193e-08, 2.005184e-08, 1.142904e-08, 0.0001605946, 9.556524e-08, 
    0.0006873425, 0.0008050824, -0.0001025014, 0.1575837, -0.0006746521, 
    0.0002964733, 0.0002752763, 9.827736e-06, 0.0003529307, 8.465096e-06, 
    6.306209e-05, 0.0003171204, 0.001397796, 0.007874586, 0.03938219, 
    0.003632108, 0.04740674, 7.926034e-06, -0.001659756, 7.871227e-05, 
    0.0004851335, 0.004687282, 0.01486338, -3.01279e-08,
  4.847988e-07, 3.539187e-05, 0.0004422448, -6.713344e-07, 2.021698e-07, 
    -7.257921e-10, -0.004510285, 0.2446772, 0.1994692, 0.001990137, 
    0.003853472, 0.001512153, 0.0007817104, 0.0004001881, 0.00179398, 
    0.001183862, 0.0004400248, 0.001792075, 0.01350661, 0.07814658, 
    -9.985422e-07, 0.02137164, 0.02772192, 0.00106101, 0.0006601933, 
    0.001037422, 0.00176395, 0.005123041, -8.428771e-05,
  0.001112848, -0.0001732839, -0.0001301233, 0.2436902, -5.538172e-05, 
    -7.576935e-08, 0.002550413, 4.262413e-07, 0.001081182, 0.010491, 
    0.1193115, 0.07976884, 0.1467321, 0.09696397, 0.1037274, 0.07463956, 
    0.02668655, 0.008264212, 0.03518128, -0.002599062, 3.319455e-06, 
    0.007292361, 0.02591634, 0.06937908, 0.01682618, 0.01427273, 0.006765373, 
    0.01480151, 0.06922957,
  0.01917736, 0.05749384, 0.02835356, 0.008037627, 0.0002481722, 
    0.0005933649, 0.0006980827, 0.08226229, 0.09701198, 0.1080374, 0.1245143, 
    0.06758796, 0.3254743, 0.3958012, 0.3521636, 0.3357032, 0.2334779, 
    0.1090198, 0.06411739, 0.04473411, 0.0052162, 0.001582531, 0.07232386, 
    0.1125914, 0.09274045, 0.218442, 0.07388806, 0.04995539, 0.06652792,
  0.1391927, 0.09507097, 0.02612723, 0.02735914, 0.05276757, 0.06453703, 
    0.08984864, 0.0575504, 0.1143762, 0.1299084, 0.09512288, 0.2496852, 
    0.2554263, 0.2232517, 0.1801733, 0.1602486, 0.2182452, 0.169549, 
    0.1609172, 0.0521794, 0.02081237, 0.1531261, 0.1198337, 0.2162994, 
    0.2330699, 0.1054228, 0.1191895, 0.07672474, 0.1736444,
  0.1668833, 0.08255437, 0.2183824, 0.0822276, 0.1623233, 0.2565547, 
    0.2062953, 0.2099515, 0.1178034, 0.09763403, 0.1622089, 0.22463, 
    0.2044906, 0.2764481, 0.1864671, 0.1848502, 0.1762059, 0.1920287, 
    0.2185059, 0.2354876, 0.2908173, 0.41356, 0.1638961, 0.186509, 0.3268174, 
    0.1750456, 0.2002557, 0.1989796, 0.2896272,
  0.4538513, 0.308951, 0.2091895, 0.2389524, 0.2498452, 0.3027318, 0.3535951, 
    0.3326328, 0.3092522, 0.3018671, 0.2708823, 0.2606898, 0.2343166, 
    0.2342298, 0.2461066, 0.2598691, 0.2803805, 0.3140673, 0.3307661, 
    0.4064739, 0.3877879, 0.2114448, 0.2693477, 0.3628927, 0.1424319, 
    0.06723358, 0.04278444, 0.198616, 0.3550046 ;

 average_DT = 730 ;

 average_T1 = 228.5 ;

 average_T2 = 958.5 ;

 climatology_bounds =
  228.5, 958.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
