netcdf atmos.1980-1981.aliq.12 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:23 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.12.nc reduced/atmos.1980-1981.aliq.12.nc\n",
			"Mon Aug 25 14:40:59 2025: cdo -O -s -select,month=12 merged_output.nc monthly_nc_files/all_years.12.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.017685e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -5.691084e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002279972, -1.968573e-05, 0, 
    -4.900259e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 9.004445e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.930638e-05, 0, 0, 0, 0,
  0, 0, 0, 0, -3.627932e-05, 0.0002584162, 0, -9.854371e-06, 0, 0, 0, 
    -1.466907e-05, 0, 0, 7.115689e-05, -8.710068e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.940235e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.745156e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004475706, -5.772568e-05, 0, 
    -5.220146e-06, -2.648391e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.15545e-06, -3.027788e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 3.597157e-05, 0, -1.701017e-05, 0, 0, 0, 0, 0, 0, -4.029116e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.21061e-05, 0.0001114764, 0, 0, 0,
  0, 0, 0, 0, 0.0001567389, 0.001291634, -7.125455e-05, 0.001003805, 0, 0, 0, 
    0.0001812679, 0, -3.29269e-05, 2.331869e-05, -1.167314e-05, 0, 0, 0, 0, 
    0, 0, 0, -8.740531e-06, 0.0008449883, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 5.119384e-06, 0, 0, -2.122534e-06, 
    -9.614941e-06, -9.520201e-07, 0, 0, 0, 0, 0, 0, 0, 0, 2.722227e-05, 
    0.0004292151, 2.071871e-05, 0.0002197014, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0001590287, 0, 0.0006294117, -0.0001431906, 
    -4.796604e-06, -7.439354e-05, -7.946302e-05, 0, 0, -3.479822e-06, 
    -7.842289e-06, 0, 0.0005203128, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001131924, -1.561369e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.793836e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -3.556745e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -3.903052e-06, 0, 0,
  0, 0, 1.019555e-05, 0, -7.082415e-05, 0, 0, 0, 0, 0, 0, -4.029116e-06, 0, 
    0, -1.269778e-06, 0, -3.479244e-06, 0, 0, 0, 0, 0, 0, 0, -8.216253e-05, 
    0.00192304, 0, 0, 0,
  0, 0, -1.215e-05, 0, 0.0003200324, 0.005519748, -0.0002126032, 0.001680847, 
    0, 0, 2.486364e-06, 0.0007018389, -1.98194e-05, 0.0001611629, 
    0.0003155575, 0.0006349063, 0, -8.12719e-06, 0, 0, 0, 0, 0, 
    -2.246194e-05, 0.002468074, 0, 0, 0, 0,
  0, 0, 0, 0, -3.409582e-07, -8.458317e-06, 0.0009191822, 9.771567e-05, 
    -1.461653e-05, 0.001290417, 4.673511e-06, 0, 1.771616e-05, 0.0008052397, 
    -7.625119e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006478633, 0.00136389, 
    0.0001146547, 0.001346277, 0, 0,
  0, 0, 0, 0, 0, -7.301156e-06, 0, 0, 0.002150281, 0.0006027027, 0.00192108, 
    0.001566686, 0.0004320119, -6.20561e-05, -0.0002071653, -3.17315e-05, 0, 
    0.0003593857, -4.399881e-05, -5.095437e-05, 0.001842941, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00116883, 0.0002128293, 0, 0, 0, 0, 0, 0, 
    0, 0, -4.008055e-05, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -6.072227e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, -1.330456e-10, 0, 0, 0,
  0, 0, 0, -4.669686e-05, 0, 3.983078e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002094171, 0, 8.869178e-05, 0, 0, 0, 0, 0, 0, 0, 0.0001130429, 
    0.0001202487, 0, 0,
  0, 0.0002762708, 0.0002715797, 0, -0.0001827082, 0, 0, 0, 0, 0, 
    -9.260352e-06, -4.029116e-06, 0, 0, -1.480779e-06, -3.798981e-06, 
    -2.091411e-05, 0, 0, 0, 0, 0, 0, 0, 0.0001380299, 0.004108055, 0, 0, 0,
  0, 0, 0.001363308, 0, 0.0005661197, 0.009941622, 0.0008865789, 0.00535397, 
    0, 0, 4.935203e-06, 0.003011122, -8.113884e-05, 0.0008088634, 
    0.0005109975, 0.00114446, 0.0001554077, -9.292138e-08, 0, 0, 0, 0, 0, 
    -5.103356e-05, 0.006141276, -2.003123e-06, 0, 0, 0,
  0, 0, -7.726129e-11, 0, -3.382712e-06, -1.322627e-05, 0.001231522, 
    0.0002605251, -5.115688e-05, 0.00307654, 1.869404e-05, -2.708329e-06, 
    -3.981342e-06, 0.003894791, 0.0002539794, 0, -5.049582e-06, 0, 0, 0, 0, 
    0, 0.0004456897, 0.002451656, 0.002779541, 0.0003003302, 0.002733629, 0, 0,
  0, 0, 0, 0, 0, -1.388393e-05, 0, -2.332907e-06, 0.003467432, 0.002149973, 
    0.003542678, 0.005299153, 0.002660238, 0.0008221365, -0.0003717663, 
    -0.0001434582, -7.14959e-05, 0.00137893, -9.968647e-05, 0.0007499311, 
    0.008849273, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002476494, 0.0003105662, 0, 0, 0, 0, 0, 0, 
    0.0004385968, 0, -7.79507e-05, 0, -2.442638e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -3.020341e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.88842e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.000868176, 0, 0, 1.917823e-05, 0, 0, 0, 0, -2.622015e-05, 
    -2.145826e-05, 0.0002347803, 0, 0, 0, 0, 0, -5.713448e-06, 0, 0, 0, 0, 
    6.040756e-05, -4.374959e-06, 9.852936e-05, 0, 0,
  0, 0, 0, -8.655633e-05, 0, 0.002009238, 0, 0, 0, 0, 0, -4.953867e-06, 
    -1.246051e-05, 0, 0, 0.0009473325, 0.0002566448, 0.003464454, 
    -1.238787e-05, 0, 0, 0, 0, 0, -6.63525e-08, 0.001150432, 0.002317872, 0, 0,
  0, 0.0003869241, 0.0007023637, 0, 0.0003602413, 1.187522e-05, 0, 0, 0, 0, 
    -2.31509e-05, -1.972333e-05, -1.397779e-05, 0, -1.099189e-05, 
    -3.216981e-05, -4.1677e-05, 0.0005755675, 0, 0, 0, 0, 0, 0, 0.0005449491, 
    0.005590935, 0, 0, 0,
  0, 0, 0.001272023, -3.123963e-05, 0.005367992, 0.01991529, 0.005016883, 
    0.009628177, 0, 0, 2.515165e-06, 0.007575216, -1.224489e-05, 0.002894268, 
    0.001453926, 0.004558312, 0.001017923, 0.0001510163, 0, 0, 0, 0, 0, 
    0.0003328049, 0.007577901, 0.000208994, 0, 0, 0,
  0, 0, -4.245728e-07, 0, -1.399284e-05, -8.784946e-06, 0.003185188, 
    0.0007295914, -7.943852e-05, 0.007255838, 0.0004982528, -4.286457e-05, 
    0.0001253646, 0.006463114, 0.000504034, 0, -2.998677e-05, -1.383031e-05, 
    0, 0, 0, 0, 0.00191228, 0.00466488, 0.00332498, 0.001626086, 0.0061153, 
    0, 0,
  0, 0, 0, 0, 0, -2.515201e-05, 0, -2.612549e-05, 0.00561646, 0.007321109, 
    0.008227731, 0.009698111, 0.007255747, 0.001963311, -0.0004944741, 
    -0.0001121842, 0.0006180631, 0.002775188, 0.001162166, 0.00254247, 
    0.02429472, 0, 0, 0, 0, -8.264202e-06, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004256283, 0.001249199, 0, 0, 0, 0, 
    -3.277293e-06, 0, 0.001230435, -9.976776e-07, 0.0005914559, 0, 
    -3.506594e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, -6.040682e-06, 0, 0, 0, 0, 0, 0, 1.923571e-05, 0, 0, 0, 0, 0, 
    -2.455672e-07, 0, 0, 0, 0, 0, 0, 0, -1.670039e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.001334547, 0, 0, 0, 0, 0, 0, 0, 0.001748101, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -4.908235e-06, -2.613733e-06, 0, 0, 0,
  0, 0, 5.551909e-05, 0.002772148, 0.0008430912, 1.506348e-06, 0.0004017961, 
    0, 0, 0, -4.779234e-05, 0.000164054, -7.597198e-05, 0.001635151, 
    -2.52116e-06, -1.340148e-05, 0, 0, 0.0007401066, -8.589362e-05, 0, 0, 0, 
    0, 0.00131347, 0.0008806604, 0.003117369, 0.0001696669, 0,
  0, 0, 0, 0.001162468, -1.742042e-06, 0.006466532, -2.011328e-05, 0, 0, 0, 
    0.0001085376, 0.0001988559, 7.55939e-05, 0.001071674, -4.283777e-07, 
    0.004492879, 0.0007548435, 0.007229215, 0.0005391391, 0, -4.353191e-06, 
    0, 0, 0, -2.126933e-05, 0.004667848, 0.006953672, 0, 0,
  0, 0.001174161, 0.001774616, 7.363917e-05, 0.001369552, 2.852408e-05, 
    -5.359485e-05, 0, 0, 0, 1.844018e-05, 3.822849e-05, -4.921162e-05, 0, 
    0.0004467412, 0.0009982232, 0.0002818756, 0.001993093, 0, 0, 0, 0, 0, 0, 
    0.001333836, 0.01025808, -1.626091e-05, 0, 0,
  0, -5.688536e-05, 0.00158552, 9.451846e-05, 0.01282771, 0.03155096, 
    0.0109334, 0.01814008, -7.848477e-06, -2.88364e-05, 5.431191e-08, 
    0.009813515, -8.620472e-05, 0.007490262, 0.006071514, 0.009006287, 
    0.002203851, 0.000427748, 0, 0, 0, 0, 0, 0.001427744, 0.01128869, 
    0.0009966416, -8.553231e-06, 0, 0,
  0, -1.124787e-06, 1.268981e-06, 0, -1.94979e-05, 0.0001301181, 0.005944446, 
    0.0008170521, -8.186264e-05, 0.01660684, 0.002296361, -0.0001743557, 
    0.001645383, 0.008585982, 0.001015463, -7.014029e-07, 0.0003189554, 
    1.280311e-05, 0, 0, 0, 0, 0.004193635, 0.006240788, 0.003887203, 
    0.002795121, 0.0100577, 0, 0,
  0, 0, 0, 0, -1.020033e-05, 0.001178012, 0, -0.0001356743, 0.01019479, 
    0.01163536, 0.01857657, 0.01751699, 0.01376103, 0.007730367, 0.001015725, 
    0.001355276, 0.002592047, 0.005921593, 0.005750212, 0.005870024, 
    0.04441396, 0, 1.795688e-05, -9.876458e-07, 0, -2.952158e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01655432, 0.002498665, 0, 0, 0, 0, 
    -3.781983e-05, 4.628642e-05, 0.003255776, 1.979706e-05, 0.002658939, 0, 
    0.000197004, 0, 0.001559653, 0, 0, 0, 0,
  0, 0, 0, 0, 6.17065e-05, 1.943625e-05, 0, 0, 0, 0, -2.725538e-09, 
    0.0001009811, 8.769913e-05, 0, -1.01364e-05, -2.139528e-05, 3.830948e-05, 
    8.971494e-05, 0, 0, 0, 0, 0, 0, 0, -2.060635e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.519398e-06, 0, 0.0005006049, 0, 
    0, 0, 0, 0, 0, 0, 0, -1.64639e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0006330149, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.26096e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.004936228, 0, 0, 0, 0, 0, 0, 0, 0.003492933, 0, 
    -1.108918e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.439916e-05, 0.0006529766, 
    -1.330983e-05, 0, 0,
  0, 0, 0.001819958, 0.006916337, 0.005035556, 0.0007589535, 0.0005377234, 0, 
    0, 0, 0.0008770577, 0.005374419, 0.0008492257, 0.009971553, 0.0001108644, 
    -3.573729e-05, -9.598997e-06, -7.097804e-06, 0.001650749, 0.0003857785, 
    1.939061e-05, -4.083854e-05, 0, 0, 0.004303087, 0.002360615, 0.006218667, 
    0.00128986, -3.57103e-06,
  0, 0, 0.0001042252, 0.008012928, -1.278119e-05, 0.01526895, 0.0003222484, 
    0, 0, 0, 0.002913956, 0.004338033, 0.0004487916, 0.00179887, 0.001707407, 
    0.01152971, 0.003890698, 0.01257799, 0.001954856, 0.0001129725, 
    -8.01869e-05, 0, 0, 0, 0.0009312046, 0.01030969, 0.01522215, 0, 
    0.001358928,
  0, 0.00275486, 0.005589302, 0.0001598085, 0.009725421, 0.0003969175, 
    -0.000127241, -3.625146e-05, 0, 0, 0.0003580764, 0.001062025, 
    0.001111676, -4.680744e-06, 0.00326779, 0.003033396, 0.001885414, 
    0.004685682, -4.106138e-06, 0, 0, 0, 0, -4.965875e-05, 0.004894787, 
    0.01515878, 0.0004808209, 0, 0,
  0, 0.000315061, 0.002363361, 0.0009816698, 0.02904657, 0.04929632, 
    0.02500018, 0.0305419, 6.422686e-05, -9.366201e-05, -6.829454e-06, 
    0.01696309, 0.002196284, 0.02057437, 0.01900556, 0.01514627, 0.006072058, 
    0.001493353, 0, 0, 0, 0, 0, 0.005197863, 0.01525152, 0.005264149, 
    7.239306e-05, 0, 0,
  0, 0.0003440462, 8.856977e-05, 0, 2.315755e-05, 0.00198976, 0.01811874, 
    0.004082712, 0.0002759924, 0.02932095, 0.005160963, 0.0006194514, 
    0.01039532, 0.01563858, 0.005305634, -2.115906e-06, 0.003930181, 
    0.0002391789, 0, -1.051866e-07, 0, 0, 0.008452528, 0.01343854, 
    0.005397201, 0.006898136, 0.01358325, -8.863488e-06, -3.864124e-06,
  0, 0, 0, 0, -4.834733e-05, 0.003404496, 0, 0.0005515544, 0.01537213, 
    0.01935133, 0.03234244, 0.02925576, 0.02314004, 0.016198, 0.007634101, 
    0.007091613, 0.006648027, 0.01070416, 0.02012781, 0.01835752, 0.07026235, 
    -1.809314e-05, 6.286937e-05, 1.740213e-05, -4.96756e-06, 0.0008061249, 
    -2.009439e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -5.393255e-05, 0.03366809, 0.003639346, 
    -9.667299e-06, -1.216049e-06, 0, -7.531497e-06, 0.001554895, 0.003166331, 
    0.007329543, 0.0004634726, 0.005040338, 0, 0.0008580978, 0, 0.009179786, 
    -2.595753e-05, 0, 0, 0,
  0, 0, 0, 0, 9.384136e-05, 0.0002958461, 0, 0, 0, -1.998962e-06, 
    5.229912e-07, 0.001919215, 0.002603594, 4.034823e-05, 0.000718596, 
    0.003148637, 0.002610768, 0.002246368, -1.020843e-05, -5.6275e-06, 0, 0, 
    0, 0, -3.748686e-05, -2.547164e-05, -2.1045e-05, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.622943e-05, 1.008051e-05, -1.324502e-05, 
    0.001559349, 0.001192375, 0.001831397, 0, 0, 0, 0, 0, 0.0003561321, 
    9.061439e-05, 0.001227798, 0.0004427558, 0.0002189899, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.208248e-07, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.002315547, 0, 1.152643e-05, 3.41755e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0006598555, 0, -1.102687e-07, 
    0.0003771278, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -9.147374e-06, 0.0001552117, 0, 0, 0.009134897, 0.0004571671, 0, 
    0.0007720534, 0, 0, 0, -1.564602e-06, 0.008141765, 0, -4.135179e-05, 
    -1.606031e-05, 0, 0, -1.142178e-05, -8.013115e-06, 0, 0, 0.000263271, 0, 
    -1.382353e-05, 0.001751291, 0.0005020029, -1.338715e-06, 0,
  -8.553295e-06, 0, 0.003904719, 0.01301585, 0.009344733, 0.002372699, 
    0.004640733, -4.852638e-06, -6.524123e-06, -4.622034e-06, 0.00312757, 
    0.01565763, 0.004556616, 0.02132373, 0.003403265, 0.001751684, 
    0.0008484413, 0.00111275, 0.004226472, 0.006166362, 0.0006487322, 
    0.002817199, -3.040841e-06, 0, 0.008601004, 0.01109593, 0.02092604, 
    0.004555974, 4.284708e-05,
  0, -6.056581e-09, 0.001777771, 0.01673104, 0.002825969, 0.03245518, 
    0.004174107, -1.463521e-05, 0, 6.505504e-05, 0.004031953, 0.01527101, 
    0.001502756, 0.00401224, 0.006509021, 0.02410458, 0.01374277, 0.02735744, 
    0.009744771, 0.0005442171, -0.0001797125, 0, 0, 2.524201e-07, 
    0.005788569, 0.01438539, 0.02585757, -1.0939e-05, 0.001961659,
  0, 0.006226792, 0.01380421, 0.0006860313, 0.01479731, 0.005964266, 
    0.001602034, 0.0002036034, -2.883469e-06, 0, 0.01278906, 0.008892126, 
    0.01301894, 7.597417e-05, 0.01190098, 0.0132699, 0.006139921, 0.01117923, 
    -9.676643e-06, -1.57459e-09, 0, 0, 0, 0.0006737126, 0.03315821, 
    0.0258349, 0.004923562, 0, -2.046209e-10,
  0, 0.005680981, 0.007923299, 0.003840078, 0.05335159, 0.06150495, 
    0.05377366, 0.04910532, 0.0009396473, -5.512245e-05, 0.0001910698, 
    0.03640256, 0.00967068, 0.04528738, 0.04795385, 0.02819178, 0.01026662, 
    0.003586433, -4.620831e-11, -1.90256e-08, 0, 0, -2.577101e-07, 
    0.02879843, 0.03879239, 0.01611618, 3.092066e-05, -3.699468e-10, 0,
  0.0004353736, 0.001284211, 0.003319572, -1.468435e-05, 0.001460542, 
    0.007339335, 0.04613065, 0.01501593, 0.007670288, 0.04823717, 
    0.009848313, 0.007346013, 0.03909918, 0.03433497, 0.006482441, 
    -1.264126e-05, 0.004680316, 0.0005683959, -5.013048e-06, -5.071443e-06, 
    0, 8.028862e-07, 0.0113626, 0.03465694, 0.009050895, 0.01853202, 
    0.02060479, -3.487458e-05, 4.664329e-05,
  0, 0, 0, 1.923899e-05, 0.0006512421, 0.00648889, 0, 0.004342723, 
    0.02110626, 0.03097169, 0.04896105, 0.05221894, 0.03478921, 0.03806211, 
    0.01815388, 0.02047104, 0.01392005, 0.01528773, 0.04306782, 0.03719369, 
    0.09347989, -0.0001036291, 0.0001572923, 1.836611e-05, -3.740851e-05, 
    0.001925545, -1.737645e-05, -8.37505e-10, 0,
  0, 0, -7.832245e-08, 0, -3.119595e-09, 0, 0.0001884913, 2.916494e-06, 0, 
    -2.386203e-05, 0.04693428, 0.004610772, -0.0001187895, -8.388909e-06, 
    0.001153284, 0.001388012, 0.01110695, 0.01475332, 0.01682766, 0.0010424, 
    0.009567702, 0.0007340294, 0.003368528, 0, 0.01341104, -4.878531e-05, 0, 
    0, -8.103657e-06,
  0, 0, 0, 0, 0.0007059738, 0.000751043, -5.898804e-07, 0, 0, 3.893142e-05, 
    0.002150419, 0.005400893, 0.006441818, 0.001917786, 0.00857034, 
    0.01442433, 0.01134507, 0.009739741, 0.00618441, 0.002417067, 
    -1.644687e-05, 0.003164823, 0.0002201146, -2.142925e-05, 0.001808052, 
    0.001202003, 3.727996e-05, 0, 0,
  0, 0, 0, 0, -8.559221e-07, 0, 0, 0, 0, 0, 0, 0.0007098406, 0.000375716, 
    0.0005009408, 0.004554025, 0.007635498, 0.005615995, 2.57805e-05, 0, 
    8.805842e-05, 0, 0, 0.001896941, 0.001471705, 0.006332266, 0.003958655, 
    0.001081008, 5.875745e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001096257, 0, 0, 0, 0, 0, 
    0, -5.644052e-06, -3.832281e-06, 0.004642262, 0.002231209, 0.0008746614, 
    0.0004928517,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, -3.095979e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001040912, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -7.61623e-08, 0, 0, 0, 0, 0, 0, 0, 0.002667575, 0.001555475, 
    -1.626401e-05, 0.001945851, 0, 0, 0, 0, 3.552723e-05, 0, 0, 0, 0, 0, 0, 0,
  0.00044908, 0.002793838, 0.001284136, 2.502181e-05, 0.01739308, 0.00465097, 
    -5.204735e-06, 0.001542685, -8.581799e-05, 0, -1.325217e-05, 
    0.0006549025, 0.013077, -5.529304e-05, 0.003837309, -2.39777e-05, 
    7.980711e-05, 0, 0.0002851292, 0.001632331, 0.0001753652, -5.186496e-06, 
    0.001516226, 0.0002626792, 0.0001925533, 0.003003007, 0.004469072, 
    0.0001262591, 0.0008143859,
  0.0007269791, -1.715666e-05, 0.005937039, 0.02499973, 0.02200554, 
    0.007801463, 0.0109894, 0.001885631, -4.426834e-05, -1.478791e-05, 
    0.006281158, 0.02690348, 0.008969171, 0.03025697, 0.01020026, 
    0.009649873, 0.003805246, 0.005862678, 0.01402298, 0.01268504, 
    0.008359982, 0.005899531, 4.984421e-05, 0, 0.01965218, 0.02661351, 
    0.04198319, 0.01267819, 0.0006719327,
  3.757092e-07, 7.716352e-05, 0.01077675, 0.03934458, 0.01873725, 0.05887251, 
    0.01825687, 0.001111503, 8.814872e-05, 0.002078374, 0.009074738, 
    0.03707587, 0.00584785, 0.007950808, 0.01247351, 0.04559854, 0.03609259, 
    0.0533358, 0.02678644, 0.004626143, 0.001295656, 0, 1.942205e-05, 
    8.132483e-05, 0.02151838, 0.03021784, 0.04592113, 0.000801223, 0.003610817,
  -5.563351e-07, 0.03121738, 0.06151444, 0.009888788, 0.04422234, 0.06633157, 
    0.02045942, 0.003975923, 0.0001180376, 2.178921e-06, 0.06420951, 
    0.03342054, 0.06130262, 0.02942393, 0.09410045, 0.07287641, 0.02548623, 
    0.02811608, 0.002392049, -1.006173e-06, -1.223477e-05, -8.879189e-07, 
    -2.246704e-06, 0.04305236, 0.1755139, 0.04165592, 0.01503892, 
    -2.410031e-05, 0.0001178215,
  -2.147971e-05, 0.07317939, 0.04500684, 0.01632123, 0.117003, 0.117224, 
    0.108391, 0.09814735, 0.02577212, 0.01252221, 0.01015515, 0.1305941, 
    0.06427479, 0.1503929, 0.1555048, 0.09795181, 0.01314366, 0.005744706, 
    -1.443974e-05, 2.787722e-06, 0, 0, 0.0005268293, 0.1408476, 0.2010786, 
    0.04102941, 0.002733186, 0.0002720039, -2.637969e-09,
  0.002282541, 0.007443378, 0.01623324, 0.001149472, 0.01312654, 0.0274434, 
    0.07940214, 0.08644648, 0.05382692, 0.1092857, 0.06227028, 0.06521257, 
    0.1660092, 0.09051032, 0.02433662, 0.005602207, 0.004780137, 0.005261126, 
    -3.337929e-05, 0.006118667, -7.927603e-06, 1.401737e-05, 0.0146547, 
    0.1281487, 0.07803307, 0.03781416, 0.03432581, -2.540689e-05, 4.208219e-05,
  1.882274e-06, -8.503695e-07, -6.676137e-07, 0.0003342972, 0.003006797, 
    0.01232534, -7.668961e-06, 0.01819559, 0.02394476, 0.06909317, 0.1375636, 
    0.1055089, 0.09942845, 0.08131997, 0.05417862, 0.04836167, 0.01967276, 
    0.02224161, 0.06845459, 0.05320622, 0.1141674, -1.237527e-05, 
    0.0004996634, 0.0004721688, 0.0001248606, 0.005909649, -0.0001634264, 
    0.0002470269, 1.406831e-05,
  3.039876e-05, 0, 0.0001831695, 3.881345e-07, -3.495051e-06, -4.329463e-10, 
    0.001924778, 0.0003158938, 4.410515e-05, 0.001998509, 0.06972208, 
    0.01936704, 0.01689616, 0.002380681, 0.001943368, 0.01240435, 0.03206206, 
    0.03420398, 0.03747378, 0.01395765, 0.02117474, 0.006904008, 0.005780834, 
    5.851658e-06, 0.01894397, -5.666608e-05, 4.774227e-05, -2.776004e-06, 
    -6.435207e-05,
  0, 0, 0, -3.641831e-06, 0.001348356, 0.0028432, -1.367173e-05, 0, 0, 
    0.01037489, 0.01617661, 0.01652486, 0.01413141, 0.006118326, 0.01886042, 
    0.02446441, 0.02548779, 0.01839428, 0.01696978, 0.009788115, 
    -8.310264e-06, 0.01141993, 0.003457264, 9.717388e-05, 0.007845796, 
    0.003003357, 0.001040798, -1.974795e-12, 0,
  0, 0, 1.804146e-06, -2.048992e-05, 0.0001113411, 0, -6.802669e-06, 0, 0, 0, 
    -1.277094e-07, 0.003440913, 0.00438217, 0.005306876, 0.01146282, 
    0.0252818, 0.01759732, 0.004609216, -5.722319e-06, 0.0002002229, 0, 
    0.0003780427, 0.005315168, 0.01800632, 0.02666198, 0.01732016, 
    0.01024331, 0.001029453, 0,
  -1.304894e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.221159e-05, 
    -2.802373e-05, 0.0001218802, 0.003025181, -1.392973e-05, -1.58417e-05, 0, 
    0, 0, 0, 0.0001964526, 0.001414222, 0.0141819, 0.01185801, 0.003846261, 
    0.002075044,
  0, 9.325429e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003028993, 
    0, 0, 0, 0, 0, 0, 0, 0.0001094737, 0.001152001, 0.0007387777, 6.156986e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.361554e-05, 0.001771405, 0, 
    -2.684002e-10, -4.557146e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0002073535, -7.690728e-06, -3.742173e-06, 0, 0, -9.59561e-07, 
    0, 4.19531e-06, -1.139078e-05, 0.002929395, 0.002856505, 0.0009275535, 
    0.004817314, 0.0001067222, -9.757451e-06, 0, 0, 0.0002695724, 0, 
    0.0003979912, 1.974216e-05, 0.0005467314, 0.001055224, 0.0002221097, 0,
  0.004099922, 0.006057248, 0.005600041, 0.001994872, 0.03430948, 0.01436026, 
    0.004269898, 0.007945146, 0.0008679376, 0.0001940851, -0.0001366168, 
    0.001719827, 0.01571343, 0.0004349313, 0.01133968, 0.0002054959, 
    0.003350679, 0.0001652273, 0.004201058, 0.005388035, 0.0008997653, 
    0.002200237, 0.00917747, 0.002938162, 0.001579837, 0.007150091, 
    0.01824013, 0.008758312, 0.00445468,
  0.01199155, 0.001773483, 0.01042747, 0.04751623, 0.0560362, 0.02865591, 
    0.02530126, 0.00904835, 0.0164507, 0.002149568, 0.01612397, 0.03681342, 
    0.02186311, 0.04291143, 0.01792888, 0.01713411, 0.00980323, 0.01721198, 
    0.02794787, 0.03083508, 0.02076199, 0.01259652, 4.760943e-05, 
    -6.023994e-06, 0.0309439, 0.0512557, 0.09127749, 0.02731516, 0.01678073,
  0.0002320421, 0.0008968791, 0.06338898, 0.1339725, 0.1033679, 0.1456502, 
    0.0821071, 0.04803991, 0.02622129, 0.02250795, 0.02905993, 0.1042604, 
    0.03554155, 0.02889526, 0.04756685, 0.1184319, 0.1066952, 0.1402168, 
    0.1834412, 0.05227648, 0.008726358, 0.000703097, 0.006773489, 0.0102608, 
    0.07532863, 0.1287526, 0.1352978, 0.0476623, 0.01711244,
  8.667949e-05, 0.09615234, 0.3206681, 0.0430757, 0.05506137, 0.09577124, 
    0.07982256, 0.01157042, 0.007041134, 8.806113e-06, 0.1355013, 0.1181109, 
    0.09016392, 0.05301901, 0.1721251, 0.2040331, 0.1524749, 0.2623653, 
    0.09513992, 0.009447211, 0.00289267, 0.0001969157, 0.001578579, 
    0.07099828, 0.1789457, 0.2400285, 0.1377496, 0.01830189, 0.002736095,
  0.002432154, 0.1870869, 0.3406356, 0.1292912, 0.1657239, 0.1610283, 
    0.1908166, 0.1538012, 0.04994366, 0.0280952, 0.02444264, 0.1363011, 
    0.08061011, 0.1757912, 0.1685094, 0.1109914, 0.04440508, 0.03701898, 
    0.003645262, 2.864212e-05, 0.0001428586, 2.843301e-06, 0.0111547, 
    0.2998097, 0.327267, 0.2464106, 0.1089992, 0.0410485, -4.414534e-06,
  0.01274833, 0.1237901, 0.153423, 0.07573787, 0.0848083, 0.0941211, 
    0.145289, 0.1327013, 0.2520628, 0.3747506, 0.1199519, 0.08020475, 
    0.1700685, 0.0933442, 0.04274876, 0.006104245, 0.01671857, 0.01704242, 
    0.0008907442, 0.01188458, 4.865084e-06, 0.0004231746, 0.01869356, 
    0.3577825, 0.2872974, 0.1077524, 0.1893839, 0.01072657, 0.0004321571,
  0.001100827, 0.004799495, 0.0001425862, 0.0006301937, 0.02573141, 
    0.04264165, -8.055902e-05, 0.0267512, 0.04558485, 0.1088052, 0.1442583, 
    0.1140295, 0.08519712, 0.06693593, 0.0672783, 0.07628161, 0.05553281, 
    0.1283563, 0.1286273, 0.147063, 0.2245922, 0.05980797, 0.01518381, 
    0.007531014, 0.02533415, 0.03022839, 0.0162554, 0.1003397, 0.001126567,
  9.334052e-05, 0.0001516216, 0.001719581, 0.002088678, -1.35665e-05, 
    1.09349e-06, 0.003476922, 0.0003955585, 0.004394499, 0.01424508, 
    0.07078872, 0.04857857, 0.01340934, 0.004544938, 0.02442974, 0.03755367, 
    0.1065539, 0.1073581, 0.1372845, 0.1082259, 0.1400848, 0.0460446, 
    0.02369965, 0.007394114, 0.04002463, 0.008120893, 0.003777252, 
    0.02988423, 0.003954103,
  -1.023226e-06, -2.051867e-06, -7.692981e-09, -2.355531e-05, 0.001431639, 
    0.01464051, 3.658076e-05, -6.248487e-08, 0, 0.02213205, 0.04119711, 
    0.06032718, 0.03935346, 0.009674238, 0.07056859, 0.08865999, 0.04545335, 
    0.04199706, 0.03736141, 0.03925315, 0.00622252, 0.04465249, 0.01722799, 
    0.03678282, 0.02708719, 0.008824631, 0.004361256, 3.716786e-05, 
    -2.784013e-05,
  1.625504e-05, 0, -1.799938e-06, 0.0004499054, 0.0009711965, 0.0003132423, 
    0.000783999, 0, 0, 0, -2.812855e-07, 0.01122038, 0.007651605, 0.01305732, 
    0.03105997, 0.05982205, 0.05282706, 0.025557, 0.008061831, 0.0007462895, 
    0, 0.002784893, 0.01607034, 0.04724664, 0.05865712, 0.04304473, 
    0.02959405, 0.007688425, -1.12739e-05,
  0.001755299, 0.000314038, 0, 0, 0, -3.638567e-08, 0, 0, 0, 0, 0, 0, 
    -3.060588e-05, 0.002915426, 0.00105311, 0.001640489, 0.01191898, 
    0.00211437, 0.001074011, -3.573105e-06, -4.316776e-07, 0, -5.833459e-05, 
    0.0003330119, 0.007637164, 0.03276474, 0.03321756, 0.02021605, 0.00606279,
  0.0002938969, 9.814647e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.021407e-05, 
    0, 0, 0.0005143805, 0.001653911, -1.420893e-05, 0, 0.000425225, 0, 0, 0, 
    0, 0.004267422, 0.006423465, 0.002235062, 0.001870128,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.331034e-06, 0, 0, 0, 0, 0, 0.0002649977, 0.0001008414, 
    0.003752243, 2.008997e-05, 5.652541e-06, -2.921585e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0.001533877, 0, 0, 0, 0.001700824, 0.002587442, 0.006992721, 0.0003579513, 
    -2.293326e-05, -1.339616e-05, -7.016132e-06, 0.002973138, -7.626584e-05, 
    0.01234594, 0.01814359, 0.01164874, 0.0100104, 0.004461279, 6.853276e-05, 
    -1.536062e-05, 3.877116e-05, 0.001000077, -1.452116e-05, 0.0006709825, 
    0.00268844, 0.004589137, 0.002481242, 0.000647251, 0.0002143954,
  0.01228904, 0.01226167, 0.0118936, 0.01187972, 0.06631086, 0.06469032, 
    0.02668108, 0.02964105, 0.02113956, 0.009897323, 0.01635586, 0.009077445, 
    0.02630075, 0.02662264, 0.03167569, 0.02954836, 0.01501596, 0.006530331, 
    0.01646603, 0.01101279, 0.009382539, 0.007459274, 0.02066341, 
    0.008599217, 0.008763856, 0.02853274, 0.03636807, 0.03954658, 0.01998288,
  0.08094704, 0.05248946, 0.03529153, 0.07732838, 0.09609957, 0.08565959, 
    0.09793057, 0.05994122, 0.05228132, 0.0448746, 0.07547912, 0.0883126, 
    0.06431854, 0.09540299, 0.0518599, 0.09153026, 0.07344463, 0.06601679, 
    0.102009, 0.1557347, 0.1273327, 0.07293119, 0.01642236, 0.00275019, 
    0.06769382, 0.1325762, 0.1725408, 0.1155264, 0.09338017,
  0.001210947, 0.0002554712, 0.07701518, 0.1267821, 0.1013976, 0.1453212, 
    0.09567514, 0.06580239, 0.03673596, 0.04613933, 0.09183107, 0.1710085, 
    0.1317342, 0.1347892, 0.146135, 0.1862425, 0.151544, 0.1944431, 0.33215, 
    0.189876, 0.08462887, 0.03551735, 0.01839191, 0.005095339, 0.09078471, 
    0.1484268, 0.1779139, 0.07943676, 0.01622418,
  7.31759e-05, 0.06531214, 0.2748097, 0.03055377, 0.04633952, 0.07820351, 
    0.07305901, 0.009371927, 0.003578066, 1.934755e-05, 0.1198037, 
    0.09517669, 0.06400955, 0.04052104, 0.1495709, 0.1734661, 0.1158906, 
    0.2220777, 0.07394711, 0.01855928, 0.01410486, 0.0002920715, 0.002539712, 
    0.06747708, 0.1469034, 0.2805196, 0.1067153, 0.009007718, 0.0001643401,
  0.0008498275, 0.147083, 0.2954655, 0.09301288, 0.134568, 0.1289955, 
    0.1532151, 0.1305699, 0.03254378, 0.02493603, 0.01513156, 0.1181412, 
    0.06524473, 0.1329082, 0.1254723, 0.0714886, 0.02660413, 0.0171743, 
    0.0001708975, 1.146194e-05, 1.524575e-05, 8.675796e-08, 0.001530804, 
    0.2706405, 0.278742, 0.216446, 0.09386764, 0.007310184, -4.911913e-06,
  0.004857638, 0.08856444, 0.08945584, 0.0377373, 0.05405152, 0.07470541, 
    0.1174289, 0.09783771, 0.1902265, 0.3300709, 0.09103127, 0.06221564, 
    0.1265739, 0.07694001, 0.02808064, 0.005508166, 0.01322427, 0.01196902, 
    0.0003011975, 0.003642717, 1.156195e-06, 0.001220708, 0.02037599, 
    0.2719882, 0.1963976, 0.08830607, 0.1357717, 0.002284392, 0.0002064323,
  3.393248e-05, 0.001989534, 0.000518956, 0.008682909, 0.02223213, 0.0245305, 
    -6.248691e-05, 0.02075456, 0.03560098, 0.08378235, 0.120197, 0.09672385, 
    0.06332886, 0.05617486, 0.05977318, 0.06036992, 0.04376611, 0.1113722, 
    0.09911905, 0.1148575, 0.1864633, 0.03296317, 0.005396113, 0.001780825, 
    0.01662426, 0.0255033, 0.03097716, 0.1009716, 0.04611934,
  0.09399657, 0.01303249, 0.0003429574, 0.001807153, 4.004827e-05, 
    0.001186177, 0.002623143, 0.001065291, 0.007118654, 0.01775291, 
    0.06449007, 0.03933818, 0.004933944, 0.004862866, 0.02379349, 0.0387246, 
    0.09632346, 0.1129017, 0.1539957, 0.1394462, 0.1164714, 0.03652053, 
    0.01470518, 0.004711299, 0.03594388, 0.04327382, 0.03600515, 0.09260939, 
    0.1408816,
  0.00673929, -0.0001310354, 0.006676686, 0.001252273, 0.003831072, 
    0.03898488, 0.01518882, -6.747054e-05, -3.047404e-06, 0.0332986, 
    0.06533293, 0.08497062, 0.04847801, 0.01954788, 0.1049765, 0.1708482, 
    0.1101379, 0.08730322, 0.08542923, 0.1028142, 0.03019065, 0.1305962, 
    0.1117491, 0.091683, 0.1300195, 0.1143499, 0.04685047, 0.0216635, 
    0.004732528,
  0.001364428, 0.0006050003, 0.0008536904, 0.002304361, 0.005978041, 
    0.002134873, 0.0009644593, 0, 0, 0, 8.728589e-05, 0.02238532, 0.01705174, 
    0.0304431, 0.07374054, 0.0979587, 0.09645486, 0.08969504, 0.0350453, 
    0.003667716, 0.0006045279, 0.01149563, 0.04779489, 0.1008153, 0.1106077, 
    0.1025207, 0.09174962, 0.02905143, 0.001162592,
  0.006018111, 0.004293935, -2.601655e-05, -2.375451e-06, 0, -1.015208e-05, 
    -7.175354e-07, 0, 0, 0, 0, 0, 0.0001246594, 0.005764627, 0.01148477, 
    0.008616449, 0.02916675, 0.01344917, 0.01465775, 0.001821817, 
    0.0001338759, -3.447459e-12, -0.0001421471, 0.002090506, 0.01690245, 
    0.0521127, 0.06749926, 0.05017008, 0.01569223,
  0.003332161, 0.001144043, -3.575514e-05, -1.798589e-08, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.444683e-05, 0.001010449, 0.001872302, 0.003777059, 
    0.008319822, 0.004555371, -1.2221e-05, 0.001905204, -1.064693e-05, 0, 0, 
    -4.468784e-06, 0.006571374, 0.01595473, 0.01447761, 0.01068334,
  0, 9.830676e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.908135e-06, 0, 0, 0, 0, 0, 0, 0, 0, -1.491554e-05, -1.922079e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0001585295, 0.001705572, -2.008108e-06, 0, 0, 0, 0, 
    0.001030536, 0.00149596, 0.007718335, 0.006141066, 0.003840259, 
    0.003006722, 0.000580955, -7.728425e-06, 0, 0, 0, 0, 0.0008433021, 0, 
    3.124887e-06, 0, 0,
  0.003249152, -4.322218e-05, -5.226993e-08, 0.0006294579, 0.005952267, 
    0.0150941, 0.02693466, 0.01438488, 0.009839699, 0.0001431344, 
    8.181398e-05, 0.003793129, 0.006683839, 0.02054188, 0.03484105, 
    0.03901917, 0.03366996, 0.02330522, 0.01321421, 0.005042277, 0.003561708, 
    0.003633197, 0.001759039, 0.003427912, 0.01324605, 0.01354882, 
    0.006689708, 0.009968141, 0.0011217,
  0.09441214, 0.08499011, 0.08732392, 0.1116035, 0.1358424, 0.1382987, 
    0.1234132, 0.1370002, 0.1113225, 0.0766037, 0.06256828, 0.06524196, 
    0.08042089, 0.09781979, 0.1130995, 0.1253358, 0.1027653, 0.1006143, 
    0.1214797, 0.08587722, 0.07754637, 0.08376843, 0.1060525, 0.03136829, 
    0.06894179, 0.101297, 0.115819, 0.09775884, 0.09434479,
  0.0889487, 0.0612468, 0.04119765, 0.07604495, 0.1141921, 0.1056167, 
    0.1249773, 0.119105, 0.09064112, 0.05861411, 0.09382781, 0.09794639, 
    0.09911284, 0.164533, 0.1203188, 0.1384868, 0.140053, 0.09750725, 
    0.1281919, 0.1846234, 0.1565619, 0.145013, 0.05804865, 0.02814997, 
    0.09517903, 0.1320372, 0.2103981, 0.1602062, 0.1077235,
  0.001209015, 0.0002163271, 0.08724865, 0.1078684, 0.09181623, 0.126393, 
    0.1198648, 0.05874289, 0.02623381, 0.03816741, 0.08073105, 0.1549683, 
    0.1215841, 0.1013959, 0.1236135, 0.1852403, 0.1282697, 0.1900554, 
    0.3021314, 0.1908453, 0.07045761, 0.02273654, 0.001725141, 0.003148134, 
    0.07437745, 0.1212101, 0.1515842, 0.05716291, 0.01150621,
  2.06085e-05, 0.05358591, 0.2416939, 0.03001096, 0.04074831, 0.07007165, 
    0.07019222, 0.01404687, 0.00200382, 1.08083e-05, 0.1102274, 0.08052513, 
    0.03719134, 0.03786657, 0.1342578, 0.1511196, 0.08710817, 0.1980606, 
    0.05996967, 0.01654792, 0.008826058, -5.087898e-05, 0.003964427, 
    0.05831819, 0.1244215, 0.2397877, 0.06720006, 0.002280907, 0.0007079446,
  7.493541e-05, 0.1069008, 0.2580048, 0.08093041, 0.1240705, 0.1223362, 
    0.1374221, 0.1236239, 0.02929731, 0.02375539, 0.01403654, 0.09907939, 
    0.06564142, 0.107276, 0.110696, 0.0588518, 0.02239922, 0.01496372, 
    0.0006096208, 2.303351e-06, 1.006609e-06, 3.375533e-07, 0.001523423, 
    0.2507301, 0.2737127, 0.1965042, 0.06954556, 0.0006105628, 1.033116e-06,
  0.003663315, 0.0675619, 0.05136579, 0.01868917, 0.03958707, 0.07054409, 
    0.1099879, 0.08178394, 0.1390136, 0.2941713, 0.06920112, 0.04559314, 
    0.1130576, 0.08047704, 0.02425517, 0.005072239, 0.009088845, 0.003976794, 
    0.0001125681, 0.0002276935, 8.125261e-07, 0.0006416682, 0.02230584, 
    0.1971652, 0.1634554, 0.0846806, 0.1103541, 0.001373033, 0.001120768,
  3.272628e-06, 0.0004065773, 0.0003314922, 0.007913874, 0.02579575, 
    0.02042854, -1.663899e-05, 0.01909087, 0.03779749, 0.07307176, 0.1038681, 
    0.08695962, 0.05964611, 0.05173737, 0.05460225, 0.0563326, 0.04357557, 
    0.09846543, 0.0833324, 0.1099088, 0.1701361, 0.02221022, 0.004312826, 
    0.002091554, 0.01073173, 0.02825366, 0.04705575, 0.08757125, 0.0269845,
  0.07314491, 0.005840543, 9.785912e-05, 0.0002336286, 9.125811e-06, 
    0.0005546053, 0.006637566, 0.002582058, 0.005570912, 0.02692036, 
    0.06470188, 0.03223753, 0.001487448, 0.01128933, 0.016397, 0.0321326, 
    0.08833857, 0.113728, 0.1618011, 0.09507106, 0.0976783, 0.02617204, 
    0.01124265, 0.00358273, 0.03598091, 0.03798118, 0.03954676, 0.07660889, 
    0.1595318,
  0.0499844, 0.01826786, 0.02080192, 0.0007377184, 0.01116019, 0.07391233, 
    0.06181901, -7.930532e-05, -3.279675e-06, 0.04233503, 0.07559653, 
    0.08734803, 0.05698003, 0.03396734, 0.1352806, 0.196289, 0.1077509, 
    0.1215032, 0.1159465, 0.1093301, 0.08982585, 0.1566608, 0.1324271, 
    0.07844312, 0.1241451, 0.1211772, 0.0959475, 0.04744056, 0.02384125,
  0.01991605, 0.003913933, 0.009485632, 0.007479368, 0.02936044, 0.01164457, 
    0.001953613, 0, -5.944968e-07, -5.16762e-10, 0.0008023161, 0.03716182, 
    0.0358858, 0.06964804, 0.118566, 0.1593886, 0.1847032, 0.1548615, 
    0.09214272, 0.02429825, 0.003583715, 0.03795948, 0.09239236, 0.1761976, 
    0.191503, 0.2177886, 0.1612483, 0.1101699, 0.04667274,
  0.04285882, 0.01761669, 0.0007546554, 0.002075333, -5.619351e-08, 
    -1.734957e-05, 0.0005882705, 0, 0, 0, 0, 0, 0.0002653324, 0.009711266, 
    0.03378781, 0.03603423, 0.05946385, 0.0361988, 0.04779297, 0.009500693, 
    0.002750952, 0.001194595, 0.003522683, 0.004511564, 0.04379909, 
    0.0956583, 0.1451271, 0.1511967, 0.1007479,
  0.02335908, 0.01328696, 0.001526146, 9.256212e-05, -3.520213e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 3.317553e-05, 0.003953528, 0.005401731, 0.01209604, 
    0.02737483, 0.009307571, 0.0003975576, 0.002625287, 8.094181e-05, 0, 0, 
    0.00392315, 0.0153655, 0.03308312, 0.05288875, 0.04580673,
  0.001942917, 0.002149774, 6.953394e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004399241, 0.001295436, -1.259191e-05, 0.001232654, 0.002151835, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0009378723, 0.002012277,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.467837e-09, 0, 0, 0, 0, 
    0, 0, -5.446688e-05, 0.003498308, -0.00115229, 0.001070663, 0, 0,
  0, 0, 0, -1.624977e-05, -1.055032e-10, 0.001449337, 0.01361339, 
    -0.0001166103, 0, 0, 0, 0, 0.004483502, 0.011634, 0.01654984, 0.02289681, 
    0.02577501, 0.0191281, 0.01023054, 0.005409189, 0.003959998, 
    0.0001392156, 1.906472e-05, 0.000180211, 0.01496248, 0.01647783, 
    0.004854428, 0.0003091106, 0.0002498972,
  0.03451947, 0.02554355, 0.01650727, 0.02304205, 0.03237609, 0.05667613, 
    0.06690219, 0.05058987, 0.06581777, 0.02655706, 0.02369065, 0.02575162, 
    0.03844099, 0.06602067, 0.08697314, 0.09967668, 0.1289421, 0.08567755, 
    0.07007782, 0.04287773, 0.03492109, 0.03396852, 0.03159874, 0.05614011, 
    0.07627203, 0.07677788, 0.04966911, 0.04979283, 0.02730669,
  0.1411104, 0.1232616, 0.1456885, 0.1871317, 0.1716211, 0.1694373, 0.163015, 
    0.1794639, 0.1883657, 0.1673494, 0.1355747, 0.119853, 0.1809921, 
    0.1506521, 0.1871196, 0.1738068, 0.1693045, 0.1333354, 0.1670296, 
    0.1571336, 0.14121, 0.1583971, 0.1784602, 0.0696129, 0.104412, 0.1434266, 
    0.1491373, 0.1410009, 0.1439308,
  0.08407659, 0.05158908, 0.03137034, 0.06951948, 0.1059725, 0.09309609, 
    0.1159597, 0.1034388, 0.0723177, 0.05597819, 0.08998042, 0.07978186, 
    0.07748471, 0.1403565, 0.1229701, 0.128943, 0.1355079, 0.09492287, 
    0.1184244, 0.1901052, 0.1659807, 0.1440208, 0.05605847, 0.05871817, 
    0.08834973, 0.1106111, 0.2073437, 0.1560737, 0.1149462,
  0.002810022, -5.774238e-06, 0.09322457, 0.102816, 0.0863924, 0.1059052, 
    0.1182084, 0.05695974, 0.02981001, 0.01575828, 0.07447982, 0.1415006, 
    0.1058693, 0.07116461, 0.1038615, 0.1650189, 0.1164795, 0.177875, 
    0.3076754, 0.1836062, 0.05954456, 0.01670146, 3.255995e-05, 0.004065651, 
    0.06025748, 0.1099513, 0.1279808, 0.0375886, 0.007490214,
  6.965661e-05, 0.05165463, 0.2157961, 0.026643, 0.03761292, 0.05815585, 
    0.05910648, 0.01953595, 0.0004794008, 7.641331e-06, 0.0744795, 
    0.05571415, 0.02945684, 0.03375794, 0.1196913, 0.1291556, 0.06256416, 
    0.170044, 0.02621371, 0.01332355, 0.003219558, -5.014245e-05, 
    0.009236759, 0.05605778, 0.09225383, 0.2173971, 0.05187484, 0.001328099, 
    0.00655791,
  0.0003582751, 0.0710242, 0.215561, 0.06445397, 0.1129495, 0.1162692, 
    0.1136431, 0.114404, 0.02302564, 0.02376671, 0.0125765, 0.07853024, 
    0.06034913, 0.09338348, 0.09272414, 0.05422458, 0.02510301, 0.01130068, 
    0.000743445, 5.273725e-07, 1.300393e-06, 5.335434e-07, 0.0005668327, 
    0.1987059, 0.2545188, 0.1680418, 0.04384318, -0.000189272, 9.144915e-07,
  0.002913132, 0.05608222, 0.03971796, 0.01368779, 0.02373037, 0.06336217, 
    0.1029145, 0.0564969, 0.07881233, 0.2353591, 0.04890198, 0.03473025, 
    0.08661416, 0.08099366, 0.02426808, 0.002738845, 0.005560479, 
    -2.737069e-05, 4.916608e-05, 0.000185344, 7.087779e-08, -2.498002e-05, 
    0.03438892, 0.1400117, 0.1405093, 0.09454386, 0.08341885, 0.0008828131, 
    0.00720413,
  4.333716e-05, 2.764667e-05, -8.778807e-08, 0.003614387, 0.02111419, 
    0.01372042, 4.166416e-05, 0.01896775, 0.04602636, 0.06631747, 0.08979216, 
    0.08228821, 0.05985368, 0.05082164, 0.04356233, 0.05584019, 0.04756181, 
    0.08654366, 0.07106268, 0.09603961, 0.1560131, 0.01451895, 0.00384964, 
    0.001518385, 0.007843751, 0.03809094, 0.07255311, 0.07821851, 0.006520974,
  0.06425375, 0.002647151, 1.992863e-06, 9.494215e-06, 6.042648e-05, 
    0.004252234, 0.01000837, 0.003857174, 0.02204879, 0.03252324, 0.06865, 
    0.029881, 0.000647108, 0.01122318, 0.009282632, 0.04054723, 0.07337666, 
    0.1125642, 0.1347877, 0.05157137, 0.07842731, 0.02087495, 0.009570999, 
    0.001503203, 0.03512932, 0.02781956, 0.03388219, 0.05925785, 0.1707766,
  0.05477848, 0.0295745, 0.02916688, 0.01743283, 0.02742118, 0.09044589, 
    0.07175653, -0.0001687758, -5.788807e-05, 0.04638796, 0.07197537, 
    0.08001187, 0.06256431, 0.04823288, 0.1295914, 0.151538, 0.111037, 
    0.1009641, 0.1230712, 0.08675618, 0.0919942, 0.148761, 0.09540828, 
    0.06274233, 0.09692962, 0.1047252, 0.07965886, 0.04312956, 0.04769505,
  0.07285754, 0.02839781, 0.04182817, 0.02319792, 0.05274028, 0.04766411, 
    0.005379675, 0.003298692, 0.0003831302, 0.0003605649, 0.01748925, 
    0.07670498, 0.04617503, 0.1084151, 0.141211, 0.1935171, 0.2340124, 
    0.1690349, 0.1047527, 0.07172204, 0.01603089, 0.05420621, 0.1465964, 
    0.1879941, 0.1706807, 0.2230231, 0.1748503, 0.1159869, 0.101058,
  0.1189694, 0.0590029, 0.02570025, 0.01592317, 0.01873058, -4.877828e-05, 
    0.001579188, 0, 0, 0, 0, -1.069781e-06, 0.005002121, 0.03138918, 
    0.1067244, 0.130244, 0.1344661, 0.07015729, 0.09899765, 0.02102973, 
    0.01304759, 0.0251677, 0.02114379, 0.01956548, 0.06318868, 0.1325369, 
    0.200126, 0.23149, 0.1785893,
  0.1199522, 0.04872388, 0.02470122, 0.001621331, 0.0002255649, 0.0003844807, 
    0, 0, 0, 0, 0, 0, 0, 0.003571381, 0.03768324, 0.07129361, 0.03656944, 
    0.06822889, 0.01422924, 0.005181214, 0.005385761, 0.0007024998, 
    -1.682362e-05, -3.504657e-06, 0.005050923, 0.02598385, 0.06886405, 
    0.1028592, 0.1331896,
  0.01099299, 0.008602149, 0.0003175009, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.074067e-05, 0.003918753, 0.005001369, 0.008213895, 0.003837466, 
    0.003679107, 0.002831075, 0, 0, 0, 0, 0, 0, -6.396401e-05, 0.008239624, 
    0.009254813,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.070428e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001486104, 0.006757068, 
    0.008204924, 0.006336131, 0.001754138, 2.588391e-06, 0, 0, 0, 0.00081019, 
    0.03166109, 0.03970593, 0.03671905, 0.03618967, 0.001071986, 0,
  0.01335769, 0.02001988, 5.930586e-05, 0.006915661, -0.0001817893, 
    0.003511234, 0.06841635, 0.0008894233, -0.0003387404, -4.991514e-10, 0, 
    -3.938823e-05, 0.004898896, 0.04870825, 0.05901415, 0.06858298, 
    0.05148195, 0.04345125, 0.03924312, 0.02509703, 0.02043322, 0.03148777, 
    0.02775165, 0.03362382, 0.03432866, 0.0324273, 0.08902562, 0.04551059, 
    0.02106396,
  0.07216278, 0.08254018, 0.08685338, 0.08384556, 0.108498, 0.09082753, 
    0.1061834, 0.09092027, 0.1073617, 0.07178079, 0.07979779, 0.07281536, 
    0.108338, 0.1438218, 0.1319123, 0.1365263, 0.1725419, 0.1442015, 
    0.149794, 0.1276392, 0.1263508, 0.109773, 0.1179538, 0.1121898, 
    0.1587987, 0.1391356, 0.1176117, 0.08370082, 0.08316629,
  0.1596713, 0.1440036, 0.1638536, 0.2085089, 0.1808154, 0.172104, 0.1637661, 
    0.179717, 0.1791456, 0.156001, 0.1511702, 0.1189908, 0.1808185, 
    0.1610818, 0.1861868, 0.1599407, 0.1581688, 0.1266644, 0.1621673, 
    0.1538911, 0.1651012, 0.1749179, 0.2082976, 0.1105791, 0.1103695, 
    0.1592189, 0.1691673, 0.1616049, 0.1578754,
  0.07288844, 0.04562609, 0.03027998, 0.06640097, 0.0998354, 0.07912087, 
    0.1102462, 0.09417918, 0.05999531, 0.05664751, 0.07645027, 0.06880871, 
    0.0676277, 0.1108408, 0.1054343, 0.1191614, 0.1258427, 0.08325502, 
    0.1057843, 0.1716901, 0.154188, 0.1404102, 0.04754354, 0.05833555, 
    0.07444968, 0.09781367, 0.1991473, 0.150521, 0.1143143,
  0.001846518, -4.656794e-05, 0.1002736, 0.09212652, 0.09083409, 0.08973283, 
    0.1060564, 0.05267524, 0.02536027, 0.00666474, 0.06303134, 0.1378393, 
    0.09167293, 0.05610478, 0.08565224, 0.1287986, 0.1080096, 0.1869254, 
    0.3112947, 0.1687823, 0.06861044, 0.01536571, 0.0001046255, 0.002908884, 
    0.0466674, 0.1150772, 0.1114114, 0.02344936, 0.005219054,
  1.522445e-06, 0.05260897, 0.1817386, 0.02248937, 0.03326673, 0.04129592, 
    0.04781305, 0.02431662, 0.003221571, 8.27551e-06, 0.04893336, 0.0366227, 
    0.02326586, 0.01904855, 0.1019436, 0.1127986, 0.0470489, 0.1440068, 
    0.01536313, 0.009715729, 0.0005111788, -1.981852e-05, 0.003852261, 
    0.04738818, 0.06578799, 0.1997105, 0.03807003, 0.0007285004, 0.002701598,
  3.468835e-05, 0.04318276, 0.171202, 0.0474897, 0.09931017, 0.1065769, 
    0.08957312, 0.1032923, 0.01571852, 0.01718995, 0.008450924, 0.05688481, 
    0.04799576, 0.07801726, 0.06924084, 0.04964735, 0.03005759, 0.01026037, 
    0.00010561, 1.737208e-07, 2.497374e-07, 3.125737e-07, 9.455244e-05, 
    0.1481724, 0.2276834, 0.1348373, 0.02571253, -0.000164015, 2.668522e-06,
  0.005658051, 0.04188277, 0.04074626, 0.009333577, 0.01406583, 0.05149562, 
    0.08879407, 0.04126465, 0.04525078, 0.1861027, 0.03396779, 0.0230179, 
    0.0637397, 0.07182679, 0.01696664, 0.001588698, 0.004546312, 
    -4.718682e-05, 3.152848e-05, 0.0005010103, -4.906024e-08, 5.943009e-05, 
    0.03114364, 0.1057586, 0.1175179, 0.09690581, 0.07303104, 0.003412752, 
    0.01749402,
  0.003434515, 1.632484e-05, 8.975331e-05, 0.004463329, 0.01632647, 
    0.008819697, 7.624679e-05, 0.02025617, 0.04468178, 0.05546097, 0.0686537, 
    0.0770989, 0.05351172, 0.04794865, 0.04620758, 0.05195569, 0.05232985, 
    0.0713041, 0.06978543, 0.100888, 0.1369588, 0.01049877, 0.00354785, 
    0.001529534, 0.009656813, 0.03845484, 0.06845943, 0.07674877, 0.003472465,
  0.0572687, 0.002367403, 1.223706e-07, 7.027639e-06, 0.0001032755, 
    0.0005898887, 0.01020287, 0.002807675, 0.03124683, 0.04220373, 
    0.07209865, 0.0252735, 0.0002999361, 0.0058338, 0.007920913, 0.04033747, 
    0.06243845, 0.1111476, 0.1183601, 0.03986479, 0.07174627, 0.0172017, 
    0.008126889, 0.001489678, 0.03639701, 0.02510899, 0.02834122, 0.04687447, 
    0.1378524,
  0.05658533, 0.02950646, 0.03002135, 0.01316667, 0.03011755, 0.08815386, 
    0.06555603, 0.0009092344, -0.0001023293, 0.04148865, 0.07144466, 
    0.08373158, 0.06643696, 0.05931555, 0.1164438, 0.1216156, 0.09985982, 
    0.0966268, 0.114075, 0.06674999, 0.08473867, 0.1328699, 0.06784515, 
    0.04437164, 0.05628845, 0.08953272, 0.0657424, 0.03951368, 0.05183242,
  0.1021233, 0.04634897, 0.08739001, 0.0588932, 0.1444274, 0.1318102, 
    0.01134543, 0.05182633, 0.006874719, 0.003193637, 0.06192483, 0.0979692, 
    0.07126743, 0.1358015, 0.1637109, 0.1959749, 0.2339618, 0.1528408, 
    0.09920739, 0.1041168, 0.06338966, 0.08364082, 0.1660935, 0.1849274, 
    0.177778, 0.2141944, 0.1516932, 0.1005314, 0.08928581,
  0.1631796, 0.1065836, 0.118149, 0.09947201, 0.1210093, 0.07624427, 
    0.004025731, -4.430207e-06, 0, 0, 0.0002384544, 0.0005026961, 0.02168173, 
    0.04866095, 0.1723051, 0.1755019, 0.1510863, 0.0935948, 0.1231018, 
    0.05518397, 0.04049968, 0.05437884, 0.06668611, 0.04694899, 0.09491245, 
    0.1505471, 0.2147853, 0.2343148, 0.1693209,
  0.1824799, 0.1315704, 0.08861396, 0.04401589, 0.04296082, 0.03461118, 
    0.02088223, 0.0002368814, 6.722397e-06, 0, 0, 0, -0.0003810252, 
    0.007886437, 0.1228671, 0.1204738, 0.1136596, 0.1156287, 0.03331492, 
    0.02869375, 0.03262921, 0.02846406, 0.01786341, 9.307227e-05, 
    0.008895128, 0.04120976, 0.0981997, 0.1478381, 0.195239,
  0.04953388, 0.03895507, 0.006716755, 0.001583541, 4.56027e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 4.710575e-05, 0.02964405, 0.05323632, 0.0651831, 0.05532537, 
    0.04338941, 0.01255819, 1.572192e-05, 0, 0, 0, -1.002592e-06, 
    -9.44462e-07, -0.000194247, 0.04355773, 0.04368203,
  0, 0, -6.017022e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.140412e-05, 
    0.00146104, 0.003487555, 0.002370222, 0.0003735115, -1.669923e-06, 
    -1.892155e-07, 0, 0, -1.625763e-05, -1.853923e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01924953, 0.02761934, 0.04051899, 
    0.04152514, 0.02213501, 0.002837522, 1.502839e-05, 0, 0, 0.009812121, 
    0.08823121, 0.09230056, 0.07244903, 0.08345064, 0.005690359, 0,
  0.03283707, 0.09913377, 0.09139871, 0.08993211, -0.001815754, 0.01418564, 
    0.1243455, 0.0181777, 4.96119e-05, -0.00108316, -4.085093e-05, 
    -0.0002399377, 0.01297281, 0.08081236, 0.1004608, 0.1044383, 0.09110803, 
    0.1033016, 0.06705803, 0.08466625, 0.0636954, 0.1056404, 0.1110199, 
    0.1106498, 0.1165825, 0.1356301, 0.2221872, 0.1176035, 0.04730289,
  0.1266666, 0.1624339, 0.145604, 0.1538482, 0.1447724, 0.1359067, 0.1529684, 
    0.1347029, 0.1529604, 0.1252805, 0.1201804, 0.145649, 0.1691518, 
    0.1799927, 0.1650087, 0.1704342, 0.1888848, 0.1731847, 0.1780548, 
    0.1555448, 0.1734348, 0.1686649, 0.1878261, 0.1679282, 0.2198816, 
    0.2094349, 0.1702272, 0.1257115, 0.14463,
  0.1690199, 0.1523404, 0.1689814, 0.2253616, 0.1910657, 0.1557521, 
    0.1626239, 0.1692153, 0.1635725, 0.1369542, 0.1462528, 0.1130581, 
    0.1792957, 0.1572556, 0.1850577, 0.1447813, 0.1455272, 0.1242875, 
    0.1502607, 0.1379573, 0.1540699, 0.172406, 0.1992676, 0.1349032, 
    0.1042586, 0.1500006, 0.1585206, 0.1506863, 0.168023,
  0.06318891, 0.03962888, 0.03237881, 0.06776309, 0.08443043, 0.06254461, 
    0.09691215, 0.08096591, 0.05227219, 0.04746388, 0.07635542, 0.06338772, 
    0.06733461, 0.09679739, 0.1018689, 0.1140035, 0.1197098, 0.07531959, 
    0.08380592, 0.1406311, 0.1468665, 0.1378815, 0.04185813, 0.03913537, 
    0.0643796, 0.09659892, 0.1862767, 0.1371065, 0.1036701,
  0.0001880282, -2.026508e-05, 0.09703793, 0.08660243, 0.09115097, 
    0.07905056, 0.09461193, 0.04400467, 0.02060458, 0.005123953, 0.05677773, 
    0.1255144, 0.07378876, 0.04696892, 0.06711686, 0.09806096, 0.09608762, 
    0.196729, 0.3157541, 0.1566371, 0.06284388, 0.01049943, 0.0003140569, 
    0.004793807, 0.03999047, 0.1051763, 0.09400901, 0.0208329, 0.003550772,
  9.843477e-07, 0.04962671, 0.1465875, 0.01836431, 0.02997393, 0.02568709, 
    0.03943368, 0.01471258, 9.944099e-05, 1.79137e-06, 0.02916491, 
    0.02481256, 0.0175307, 0.01434922, 0.09103239, 0.09433784, 0.04471269, 
    0.11754, 0.009777999, 0.00402612, 0.0004023621, -5.299367e-06, 
    0.00131334, 0.04036013, 0.0610432, 0.1894068, 0.03802495, 0.0001303475, 
    0.0001765739,
  3.602952e-05, 0.03227277, 0.125274, 0.03519953, 0.1016697, 0.1018803, 
    0.0810356, 0.09997909, 0.01019469, 0.01413355, 0.007227413, 0.04886735, 
    0.03328228, 0.06961048, 0.05789527, 0.03603339, 0.03726184, 0.007431779, 
    0.0001221359, 1.121135e-07, 1.010974e-07, -2.137012e-06, 0.0001911096, 
    0.104745, 0.2098254, 0.1121304, 0.01088118, -1.087022e-05, 3.846038e-06,
  0.02509576, 0.02658845, 0.03711123, 0.007450075, 0.01033702, 0.04396711, 
    0.074095, 0.03664608, 0.03617699, 0.1520799, 0.0295591, 0.0177827, 
    0.04768928, 0.06396671, 0.01571048, 0.006159123, 0.004925576, 
    0.0003961633, 8.825435e-06, 0.0009822664, -2.728239e-05, 0.002777972, 
    0.03330301, 0.0864855, 0.09528533, 0.0948648, 0.06637035, 0.02569721, 
    0.03005639,
  0.008374808, 7.534219e-06, 3.103648e-05, 0.008821724, 0.01706205, 
    0.007819545, 0.0002025684, 0.02321178, 0.0430197, 0.04404478, 0.06385206, 
    0.0708451, 0.04653854, 0.04933768, 0.04978567, 0.05740107, 0.05613679, 
    0.06885779, 0.07697713, 0.1094959, 0.1284775, 0.01102285, 0.003084144, 
    0.001416653, 0.01225677, 0.04060016, 0.04360003, 0.06277023, 0.008475938,
  0.04560955, 0.00319807, 8.242639e-09, 7.952664e-06, 7.751215e-05, 
    -7.919353e-06, 0.01030306, 0.001297693, 0.01623515, 0.04442427, 
    0.07376874, 0.02372437, 0.0009334472, 0.003591971, 0.004841754, 
    0.03664082, 0.05130174, 0.1033616, 0.1006391, 0.03178453, 0.06181046, 
    0.0136566, 0.005959762, 0.001232771, 0.03532562, 0.01499936, 0.01706041, 
    0.03777019, 0.1188603,
  0.04953596, 0.01883388, 0.02562675, 0.01294268, 0.02760287, 0.08326412, 
    0.06333938, 0.006967714, 0.0005641907, 0.04823517, 0.06579809, 
    0.06585859, 0.07317034, 0.07049223, 0.08876448, 0.1122593, 0.09423246, 
    0.09431105, 0.1054593, 0.05187761, 0.07884219, 0.1192474, 0.04140086, 
    0.04059184, 0.04154769, 0.07532968, 0.04206583, 0.02165754, 0.06114525,
  0.09389096, 0.04245793, 0.1110352, 0.1181621, 0.1769894, 0.1780862, 
    0.02006864, 0.1148531, 0.05674043, 0.04348072, 0.09504926, 0.1144955, 
    0.09040864, 0.1573475, 0.1732301, 0.1973639, 0.2316413, 0.1460086, 
    0.0874354, 0.1150012, 0.08457173, 0.08794986, 0.1612881, 0.1868745, 
    0.1784137, 0.207964, 0.1401823, 0.09669344, 0.07818868,
  0.1723911, 0.1431717, 0.1631129, 0.2122525, 0.2166955, 0.2050152, 
    0.1549071, -0.0001068722, -3.940617e-06, 0.006022076, 0.01058659, 
    0.00470856, 0.05532295, 0.0714828, 0.2053028, 0.2113321, 0.155096, 
    0.1002474, 0.1432075, 0.08234932, 0.06535639, 0.1057457, 0.1273161, 
    0.08874302, 0.1436212, 0.181901, 0.2476819, 0.2290772, 0.1825581,
  0.2418374, 0.1831244, 0.1409888, 0.1296381, 0.144287, 0.1333147, 0.117397, 
    0.08380207, 0.0412746, -3.675589e-05, -6.970007e-05, -0.0002508326, 
    0.006123879, 0.01767632, 0.1427591, 0.1606503, 0.1308243, 0.1530404, 
    0.07506789, 0.08526, 0.09860846, 0.1017747, 0.04478428, 0.01790043, 
    0.05248766, 0.07078214, 0.1347391, 0.1742996, 0.2227441,
  0.08902169, 0.101133, 0.03052997, 0.0288197, 0.0103762, 0.01152418, 
    0.01088604, -0.0003281774, 0, 0, 0, 0, -0.0002954505, 0.01816963, 
    0.09083308, 0.116903, 0.1158097, 0.102884, 0.1071334, 0.076447, 
    0.01881651, 0.01149687, -0.0002780611, -0.0004620315, 0.01148379, 
    -3.092151e-05, 0.0002458392, 0.09771901, 0.08503556,
  0.02182166, 0.01986232, 0.002522497, 0.000195617, 0.002432476, 2.77207e-05, 
    1.058589e-05, 4.370222e-08, 0, 0, 0, 0, -0.0001111508, 0.001844744, 
    0.006205137, 0.02444014, 0.0318449, 0.03114494, 0.02223484, 0.01907382, 
    0.004114291, -0.0001210365, -6.875007e-05, 0.0006429329, -7.058584e-05, 
    -1.795663e-05, -1.630605e-07, -0.0009970221, 0.0189334,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.191458e-10, 0.000144143, 0.0381065, 
    0.07655363, 0.09496227, 0.1306055, 0.08195886, 0.02109666, 0.002479618, 
    0.001062409, 0.0002563911, 0.03287535, 0.1514163, 0.133615, 0.1424442, 
    0.1161311, 0.03969336, 0.0007628592,
  0.1119955, 0.2412429, 0.1983351, 0.2309939, 0.00290539, 0.05482649, 
    0.1775567, 0.05496857, -0.002000117, 6.916723e-05, -0.000300171, 
    0.01092866, 0.03080491, 0.1786266, 0.1650116, 0.1670819, 0.165362, 
    0.1860173, 0.1360839, 0.190516, 0.1147162, 0.1899824, 0.1904894, 
    0.2187937, 0.2513046, 0.2244865, 0.2626209, 0.1295643, 0.07835224,
  0.140783, 0.250443, 0.212257, 0.2148856, 0.183395, 0.175984, 0.1644543, 
    0.1572541, 0.1873082, 0.1614972, 0.1920861, 0.2119612, 0.2317643, 0.2217, 
    0.1968873, 0.1864787, 0.1817507, 0.1736839, 0.1896552, 0.1984797, 
    0.2415353, 0.2511509, 0.2667217, 0.2142392, 0.2375217, 0.2182433, 
    0.225406, 0.1424828, 0.1855266,
  0.1626392, 0.1546, 0.1649909, 0.2115016, 0.1806432, 0.1602703, 0.1706389, 
    0.1644427, 0.1511654, 0.127235, 0.1474591, 0.1367211, 0.1730538, 
    0.1533871, 0.1724979, 0.1331322, 0.1244637, 0.1202491, 0.1377858, 
    0.1272096, 0.146936, 0.1595516, 0.1988005, 0.1403247, 0.09489694, 
    0.1408585, 0.1463263, 0.1489356, 0.1748766,
  0.05877829, 0.03429618, 0.02715174, 0.06928115, 0.07779835, 0.05441508, 
    0.09908908, 0.08285339, 0.04614004, 0.02741913, 0.06881213, 0.05376121, 
    0.0647317, 0.08806327, 0.0911157, 0.09347621, 0.1044933, 0.06543497, 
    0.06891322, 0.1326863, 0.1144433, 0.1330142, 0.03982224, 0.02641198, 
    0.05799062, 0.09316954, 0.1664235, 0.1344288, 0.08967453,
  0.001777561, -8.434855e-06, 0.08392034, 0.08229704, 0.09353831, 0.07682839, 
    0.09011358, 0.02457925, 0.01526335, 0.003441559, 0.05368855, 0.1131826, 
    0.0566991, 0.04219973, 0.05245822, 0.08174276, 0.0985461, 0.1929908, 
    0.3224248, 0.09314846, 0.06547794, 0.007372981, 0.0009301889, 
    0.002589328, 0.03524413, 0.09388237, 0.09343118, 0.02908401, 0.004051059,
  6.575382e-07, 0.04440415, 0.1211388, 0.01624833, 0.03083352, 0.01642129, 
    0.04824055, 0.01086706, -1.44921e-05, -1.038606e-06, 0.02307168, 
    0.01708105, 0.01602471, 0.007454041, 0.08040531, 0.07128063, 0.05142576, 
    0.1060857, 0.006644255, 0.001950068, 6.714086e-05, 3.858119e-08, 
    5.585002e-05, 0.03050933, 0.05830047, 0.1842144, 0.03457935, 
    4.149691e-05, 1.817404e-06,
  6.56136e-05, 0.03417415, 0.09865661, 0.02884164, 0.09800833, 0.09984805, 
    0.07604694, 0.101345, 0.008060447, 0.01116305, 0.009151381, 0.04051331, 
    0.02541598, 0.07130098, 0.04997373, 0.03160567, 0.03633163, 0.007140521, 
    0.0001844991, 4.211102e-08, 1.772748e-08, 8.559056e-08, 0.001240132, 
    0.08743767, 0.2033892, 0.102043, 0.005955402, -1.794009e-05, 5.076439e-06,
  0.06834232, 0.01640469, 0.04375285, 0.00610608, 0.01472589, 0.04594702, 
    0.05769844, 0.03588954, 0.02301729, 0.1435407, 0.03051521, 0.01652686, 
    0.0371244, 0.05134532, 0.01510788, 0.002666082, 0.004590208, 
    -3.770547e-05, 6.768166e-05, 0.0005864107, 0.0001772578, 0.0009052714, 
    0.03832268, 0.07538125, 0.07870129, 0.09496729, 0.07594395, 0.03298282, 
    0.0354716,
  0.01467595, 3.333487e-06, 0.0001701444, 0.008282918, 0.01515916, 
    0.008202914, 8.283103e-05, 0.01635981, 0.0374711, 0.04813511, 0.06548985, 
    0.06746837, 0.04461465, 0.05064368, 0.05104145, 0.07027861, 0.06683193, 
    0.06433317, 0.07530156, 0.1183624, 0.1213578, 0.01469119, 0.003954835, 
    0.002275848, 0.01806617, 0.02980182, 0.02460451, 0.03284794, 0.01158264,
  0.04277709, 0.003294793, 2.436623e-08, 7.239853e-06, 8.95679e-05, 
    0.001677378, 0.01084035, 0.001978054, 0.00543938, 0.040242, 0.07396766, 
    0.01576318, 0.0004531507, 0.002643454, 0.002596564, 0.03159572, 
    0.04950359, 0.0844666, 0.1014825, 0.02444641, 0.05360316, 0.008678405, 
    0.003599373, 0.001061649, 0.03444958, 0.005716563, 0.0149236, 0.01944226, 
    0.07493869,
  0.03323724, 0.02358486, 0.02394869, 0.01562651, 0.02361425, 0.08636599, 
    0.06832998, 0.007930619, 0.01128951, 0.05536789, 0.06438064, 0.05310483, 
    0.08471388, 0.07755098, 0.06905298, 0.1061442, 0.08680011, 0.09031999, 
    0.09414311, 0.04038706, 0.07866929, 0.09157667, 0.03690964, 0.02280109, 
    0.02863519, 0.07972495, 0.02862168, 0.008908518, 0.06009137,
  0.07144253, 0.04113689, 0.1058731, 0.1859435, 0.1615618, 0.1639944, 
    0.03954103, 0.143629, 0.0733581, 0.1034194, 0.1061559, 0.1102038, 
    0.1007474, 0.1601902, 0.1794887, 0.1961532, 0.215966, 0.1373169, 
    0.09191242, 0.1365838, 0.09272847, 0.0816626, 0.1622135, 0.1899357, 
    0.1762515, 0.1836238, 0.1254055, 0.08553918, 0.085756,
  0.1794772, 0.1592681, 0.1978521, 0.2445813, 0.233002, 0.2348356, 0.2523173, 
    0.001695492, 0.005974972, 0.01968702, 0.04325933, 0.01705661, 0.1530455, 
    0.1346353, 0.2331427, 0.2335541, 0.1435818, 0.1127523, 0.1439597, 
    0.0882697, 0.09298012, 0.1415444, 0.180983, 0.1474351, 0.1558554, 
    0.203304, 0.2585275, 0.228488, 0.1824998,
  0.2852822, 0.2303226, 0.1824537, 0.2123126, 0.1967542, 0.1876305, 
    0.1740521, 0.1604437, 0.1361508, 0.08038145, 0.02119329, 0.01011835, 
    0.01495165, 0.05268668, 0.2063591, 0.1897944, 0.1888466, 0.2169858, 
    0.1282345, 0.1523603, 0.187654, 0.1517196, 0.1084916, 0.0909391, 
    0.1035084, 0.1227957, 0.1832381, 0.2395676, 0.2825073,
  0.1698501, 0.1803829, 0.1184604, 0.09484975, 0.06761898, 0.0722101, 
    0.07675787, 0.04233209, 0.006728672, 0.004332801, -3.174357e-05, 
    -0.0001454055, 0.01108024, 0.06806467, 0.1392784, 0.1532303, 0.1753857, 
    0.1659954, 0.1739347, 0.1433635, 0.08202851, 0.03183627, 0.0423323, 
    0.006803819, 0.05287673, 9.601997e-05, 0.004468851, 0.154225, 0.1626633,
  0.100546, 0.0840772, 0.05258947, 0.03710751, 0.03635971, 0.01700902, 
    0.0125946, 0.006722001, 0.01726584, 0.01445547, 0.009819349, 0.009111786, 
    0.01758008, 0.02987616, 0.05563468, 0.05300866, 0.05405152, 0.05628113, 
    0.05283535, 0.04999239, 0.04900397, 0.03857485, 0.006317989, 
    0.0002345467, 0.001305579, 7.822777e-05, -0.0007914932, 0.003700451, 
    0.07137547,
  0.00199512, 0.001180082, 0.0003650437, -0.0004499943, -0.001265032, 
    -0.00208007, -0.002895108, -0.0001259678, -5.676929e-05, 1.242922e-05, 
    8.162773e-05, 0.0001508263, 0.0002200248, 0.0002892233, 0.001695169, 
    0.001706385, 0.001717602, 0.001728818, 0.001740034, 0.001751251, 
    0.001762467, -0.003456842, -0.002722219, -0.001987596, -0.001252973, 
    -0.0005183503, 0.0002162727, 0.0009508957, 0.00264715,
  -0.001071631, -1.023944e-05, -3.364077e-07, 0, 0, -0.0003379439, 0, 0, 0, 
    0, 0, -1.199864e-05, 0.001197911, 0.08303577, 0.08382231, 0.1195551, 
    0.1716282, 0.2319879, 0.06345523, 0.01641236, 0.009571344, 0.01935981, 
    0.1065082, 0.1294063, 0.1229238, 0.1319026, 0.1421696, 0.07377426, 
    0.01950472,
  0.1188314, 0.2479757, 0.2058359, 0.2775636, 0.04990463, 0.1268362, 
    0.2363921, 0.08815551, 0.02552782, 0.04883801, 0.01336061, 0.01860156, 
    0.09381153, 0.199522, 0.19119, 0.1989687, 0.1818029, 0.2156038, 
    0.1504031, 0.2017125, 0.1226794, 0.1948742, 0.2326193, 0.2912613, 
    0.2868286, 0.2178687, 0.2588639, 0.1247487, 0.1035636,
  0.135907, 0.2594708, 0.2357305, 0.2357229, 0.1995023, 0.1813658, 0.171894, 
    0.150637, 0.1998728, 0.1751167, 0.2289829, 0.2557692, 0.2398265, 
    0.2297834, 0.2025941, 0.1994161, 0.1789585, 0.1729018, 0.2048507, 
    0.2226323, 0.2823609, 0.2780979, 0.2740352, 0.2250172, 0.2519158, 
    0.2307572, 0.2128927, 0.1364872, 0.1862306,
  0.1661991, 0.1519042, 0.1634004, 0.1965236, 0.1646418, 0.1646097, 
    0.1684517, 0.1768365, 0.1678018, 0.1456398, 0.144399, 0.1548205, 
    0.1717381, 0.1504501, 0.1608113, 0.112231, 0.09880535, 0.1093411, 
    0.1138857, 0.1181863, 0.1417476, 0.1549909, 0.1831324, 0.1464659, 
    0.08562981, 0.1367165, 0.1459142, 0.1538581, 0.1739076,
  0.06122247, 0.02820023, 0.02259443, 0.0783257, 0.07129028, 0.04706212, 
    0.09031315, 0.07320944, 0.0368409, 0.02516529, 0.0711538, 0.05089185, 
    0.05940305, 0.08043861, 0.08133058, 0.08902851, 0.09278198, 0.05212544, 
    0.05679541, 0.1173812, 0.1177205, 0.1140492, 0.03611009, 0.02186296, 
    0.0542464, 0.09454854, 0.1510446, 0.1314984, 0.09751739,
  0.0005691197, 4.802282e-06, 0.07656613, 0.05939741, 0.08311, 0.07653989, 
    0.07920226, 0.01937685, 0.006444084, 0.0005049577, 0.06955708, 0.1007248, 
    0.05427265, 0.03754685, 0.03964511, 0.06659729, 0.07469692, 0.181814, 
    0.2840505, 0.06703363, 0.05757184, 0.004777981, 0.0008106609, 
    0.001916429, 0.03781623, 0.08692604, 0.09765926, 0.03328981, 0.00755854,
  5.717746e-07, 0.04346459, 0.1078017, 0.02175134, 0.0311016, 0.01102005, 
    0.05659946, 0.01422293, -3.16861e-06, 6.440809e-06, 0.02102832, 
    0.01357003, 0.01378604, 0.01123347, 0.07247727, 0.05964053, 0.06385587, 
    0.09002912, 0.007623084, 0.001821596, 7.623377e-05, 4.874347e-08, 
    3.9362e-06, 0.02135059, 0.06574681, 0.1741082, 0.02808059, 0.000113999, 
    4.697571e-07,
  0.0006426761, 0.03479379, 0.08448824, 0.03991914, 0.1036127, 0.09513313, 
    0.07726991, 0.09554186, 0.006360458, 0.01182075, 0.01022563, 0.03698822, 
    0.02103085, 0.06460451, 0.04726163, 0.03493506, 0.03508166, 0.006297072, 
    0.0005546008, 1.704956e-08, 5.705978e-10, 9.389026e-09, 0.003652286, 
    0.07771946, 0.2005899, 0.09065502, 0.005389958, -1.897707e-05, 7.99188e-05,
  0.1412203, 0.01116368, 0.05243955, 0.008632407, 0.01330547, 0.03707797, 
    0.04697758, 0.03332437, 0.02379155, 0.1365096, 0.03264445, 0.01391203, 
    0.02948627, 0.04433684, 0.01569331, 0.001929558, 0.004740998, 
    5.739045e-05, 0.0003520227, 0.0004671293, 0.002830032, 0.002393644, 
    0.05512226, 0.08627547, 0.07168564, 0.08776799, 0.06632235, 0.03584831, 
    0.05744115,
  0.01500039, 1.790578e-06, 0.005592717, 0.00618095, 0.01489189, 0.00739858, 
    0.0001092192, 0.00875731, 0.03467575, 0.04639836, 0.07422581, 0.07196963, 
    0.04408362, 0.04750038, 0.04864477, 0.07029827, 0.07800458, 0.05573519, 
    0.08327202, 0.1189815, 0.1107939, 0.01447771, 0.005036104, 0.004081184, 
    0.02558118, 0.02078836, 0.01337125, 0.008003333, 0.02718119,
  0.0444502, 3.83257e-05, 1.764702e-08, 7.42124e-06, 0.0001895388, 
    0.0007571302, 0.008378018, 0.0002738293, 0.001745633, 0.03990498, 
    0.08075822, 0.01574859, 0.000557256, 0.003096485, 0.0006255193, 
    0.03056607, 0.04560564, 0.06646988, 0.08467829, 0.01800315, 0.04609302, 
    0.005616843, 0.0030218, 0.001152048, 0.03325091, 0.002210761, 0.01543514, 
    0.00743096, 0.06407666,
  0.03038519, 0.02265434, 0.02241856, 0.02197961, 0.02340929, 0.08825028, 
    0.0718143, 0.007629205, 0.03530459, 0.05139229, 0.06523541, 0.05558607, 
    0.0800522, 0.08088072, 0.0454291, 0.1045307, 0.06956662, 0.08825435, 
    0.0840239, 0.04185311, 0.0754854, 0.07548785, 0.03575267, 0.01913684, 
    0.02930617, 0.05552754, 0.02518844, 0.006417735, 0.04686006,
  0.06297662, 0.042674, 0.1038202, 0.2094994, 0.1457736, 0.1432613, 
    0.0982418, 0.1371643, 0.08657152, 0.1117445, 0.09596275, 0.1006396, 
    0.1067922, 0.1703915, 0.1694557, 0.1927353, 0.1975854, 0.1305166, 
    0.09978116, 0.1518196, 0.1001143, 0.07113086, 0.1688034, 0.1881225, 
    0.1815977, 0.1785145, 0.107537, 0.07934728, 0.08645,
  0.1625134, 0.1705161, 0.225058, 0.2503828, 0.2338606, 0.2467301, 0.2515372, 
    0.06476719, 0.04434038, 0.07005429, 0.09595221, 0.05372814, 0.2133309, 
    0.218562, 0.248574, 0.2525377, 0.1661364, 0.1323622, 0.1607739, 
    0.1171976, 0.1147974, 0.1711667, 0.195069, 0.1729886, 0.1661741, 
    0.2104489, 0.2748462, 0.2228723, 0.1809387,
  0.3095551, 0.2716222, 0.2402635, 0.2617798, 0.2466015, 0.2679252, 
    0.2461734, 0.2491911, 0.219979, 0.1916351, 0.07536478, 0.01303758, 
    0.02443356, 0.1360324, 0.2558465, 0.217745, 0.2384927, 0.2842652, 
    0.2000197, 0.2148186, 0.2446418, 0.2014869, 0.1457148, 0.2068474, 
    0.1475438, 0.1940892, 0.2103136, 0.2592018, 0.2975146,
  0.1857825, 0.2660897, 0.2208358, 0.1646728, 0.1356653, 0.1636865, 
    0.2141788, 0.153035, 0.07582139, 0.05372889, 0.0100806, 0.04602616, 
    0.07428918, 0.1834537, 0.1920547, 0.2143423, 0.2374734, 0.2433916, 
    0.2617857, 0.2084552, 0.1346556, 0.06585616, 0.1077874, 0.04972088, 
    0.07733772, 0.005188059, 0.0171868, 0.2064397, 0.1850082,
  0.1478756, 0.1485455, 0.1223013, 0.09603535, 0.07827938, 0.03854437, 
    0.04711851, 0.03969545, 0.04877608, 0.04531954, 0.0586066, 0.07641357, 
    0.06823592, 0.08011211, 0.08936605, 0.07589464, 0.07254719, 0.06874425, 
    0.0985167, 0.1129046, 0.09031455, 0.08013616, 0.02056379, -0.000944298, 
    0.001091632, 0.0005679057, -0.002553786, 0.04067416, 0.1279624,
  0.03363658, 0.03295411, 0.03227164, 0.03158918, 0.03090671, 0.03022424, 
    0.02954177, 0.03203926, 0.03053847, 0.02903768, 0.02753688, 0.02603609, 
    0.0245353, 0.02303451, 0.01235709, 0.01413985, 0.01592262, 0.01770539, 
    0.01948815, 0.02127092, 0.02305368, 0.03557501, 0.03597551, 0.036376, 
    0.03677649, 0.03717699, 0.03757748, 0.03797798, 0.03418255,
  0.04353306, -0.001942705, -0.0001087095, -1.421287e-06, 0.0007895736, 
    0.001255522, -0.0004001631, -0.0001742851, 0.0001129594, 0.001718368, 
    -0.0005737437, 0.001473686, 0.01025894, 0.109887, 0.08347093, 0.1141766, 
    0.165893, 0.2487676, 0.1363018, 0.07135682, 0.05921858, 0.07909531, 
    0.1617391, 0.1188131, 0.1115666, 0.1223384, 0.1401954, 0.1032801, 
    0.08173196,
  0.1118095, 0.2230526, 0.1922932, 0.2736115, 0.2036462, 0.1918257, 
    0.2715183, 0.1263255, 0.08511254, 0.1138575, 0.07060471, 0.03067521, 
    0.1418826, 0.193625, 0.1930756, 0.2076878, 0.1899706, 0.223374, 
    0.1562788, 0.1986868, 0.1272879, 0.1846446, 0.2290244, 0.2854922, 
    0.2747309, 0.1945561, 0.2504193, 0.1130016, 0.1028495,
  0.137342, 0.2646297, 0.2655407, 0.242714, 0.2124978, 0.1889829, 0.1833118, 
    0.151854, 0.2047289, 0.182855, 0.2636514, 0.265269, 0.2452645, 0.2312654, 
    0.2250436, 0.2087154, 0.1773269, 0.1954042, 0.2302025, 0.2404876, 
    0.2876644, 0.2863988, 0.2778973, 0.2293976, 0.240999, 0.2480243, 
    0.2165641, 0.1419282, 0.1844597,
  0.1668722, 0.1512783, 0.1619757, 0.1885982, 0.1623866, 0.1559981, 0.161421, 
    0.1806671, 0.1728686, 0.1495451, 0.1447585, 0.1294478, 0.1502405, 
    0.1512503, 0.1491197, 0.09920132, 0.09343481, 0.0988972, 0.1138152, 
    0.1108685, 0.1477236, 0.1478429, 0.1772044, 0.1425272, 0.07912253, 
    0.1350079, 0.141172, 0.1529332, 0.1736863,
  0.05602697, 0.02468768, 0.01973573, 0.08876577, 0.06753649, 0.04378296, 
    0.09496931, 0.06630701, 0.02995245, 0.02808292, 0.07344745, 0.04840928, 
    0.05746939, 0.07803845, 0.07206331, 0.08492369, 0.07771927, 0.04230842, 
    0.04561918, 0.1184175, 0.1025578, 0.1033993, 0.032405, 0.01756562, 
    0.06082851, 0.09029961, 0.1393111, 0.1149016, 0.08205135,
  0.002421481, 2.195312e-05, 0.07228725, 0.04535956, 0.07907934, 0.08205575, 
    0.07165285, 0.01212835, 0.003936179, 0.0006204359, 0.0776606, 0.08199738, 
    0.04985123, 0.0331741, 0.03211745, 0.05982034, 0.05106352, 0.1757829, 
    0.2359233, 0.05351212, 0.05992549, 0.003258978, 0.001263581, 0.00146562, 
    0.04177821, 0.07707951, 0.1091983, 0.03248404, 0.008876191,
  1.15474e-05, 0.05223736, 0.0987138, 0.02669993, 0.03238383, 0.01007485, 
    0.05881615, 0.02516294, 9.692926e-07, 0.0001005652, 0.03109757, 
    0.01819148, 0.01275298, 0.01077701, 0.07025546, 0.0640789, 0.07190333, 
    0.08617587, 0.00858635, 0.001873283, 0.0006348405, 7.438044e-08, 
    5.352204e-06, 0.01681964, 0.08338514, 0.1894286, 0.02311413, 9.44792e-06, 
    3.569856e-07,
  0.004869028, 0.04840045, 0.0837332, 0.04802062, 0.1085879, 0.09616701, 
    0.0844699, 0.0969286, 0.006837221, 0.01434475, 0.01056318, 0.0402465, 
    0.02198591, 0.06930859, 0.04965456, 0.03900536, 0.03382459, 0.008430085, 
    0.0009769404, 2.122831e-07, 7.050049e-09, -7.910498e-07, 0.003456753, 
    0.07552385, 0.2240333, 0.08435486, 0.00443603, 0.0001098079, 0.003511293,
  0.2480674, 0.01313526, 0.06744503, 0.01554635, 0.02540125, 0.02989199, 
    0.0485343, 0.04071046, 0.02743827, 0.1357941, 0.03379023, 0.009381545, 
    0.02679294, 0.04305075, 0.01604929, 0.003585077, 0.001702867, 
    0.0004170978, 5.409856e-05, 4.697813e-05, 0.007091617, 6.550246e-05, 
    0.08273438, 0.1026977, 0.07479313, 0.07934874, 0.06713813, 0.03800419, 
    0.1127603,
  0.00194528, 1.236564e-06, 0.008538604, 0.005048009, 0.01334613, 
    0.006461184, 0.0001588339, 0.00507451, 0.03494419, 0.04159208, 
    0.09026483, 0.07332911, 0.0445478, 0.04743335, 0.04764133, 0.0725053, 
    0.09116995, 0.05374051, 0.08758406, 0.1183025, 0.1070922, 0.0171124, 
    0.005698054, 0.00578062, 0.03006302, 0.01227276, 0.008690288, 
    0.004679522, 0.00871657,
  0.04086183, 3.20671e-06, 1.532292e-08, 6.957397e-06, 0.0001523044, 
    0.0001602398, 0.007054846, 9.992784e-05, 0.0001016633, 0.04876573, 
    0.09601976, 0.01663933, 0.0009191048, 0.006569764, 0.000725801, 
    0.02594903, 0.04117937, 0.06197276, 0.06829023, 0.01246951, 0.03227685, 
    0.004694864, 0.00236013, 0.001846312, 0.03274629, 0.002816819, 
    0.02235671, 0.004799562, 0.04564817,
  0.02125488, 0.01869385, 0.0225142, 0.02404622, 0.02268121, 0.07847902, 
    0.06556811, 0.01113767, 0.08469579, 0.06069965, 0.0692069, 0.06589488, 
    0.08729284, 0.08419021, 0.04424241, 0.1013563, 0.0626998, 0.07620255, 
    0.07058403, 0.03002348, 0.07282413, 0.06577595, 0.03479708, 0.01645662, 
    0.02558516, 0.04512878, 0.02354692, 0.005818384, 0.03648585,
  0.05422007, 0.04079774, 0.09950456, 0.2104632, 0.1413433, 0.134341, 
    0.1322735, 0.1277575, 0.08624507, 0.1015763, 0.09029378, 0.09424827, 
    0.1035244, 0.164135, 0.1625641, 0.1844197, 0.1869489, 0.1129293, 
    0.088385, 0.1559579, 0.1049166, 0.06056635, 0.16028, 0.1741488, 0.170986, 
    0.1769219, 0.1035169, 0.0705381, 0.08539619,
  0.1550706, 0.17102, 0.1962659, 0.2517684, 0.2374434, 0.2408913, 0.2557583, 
    0.1527941, 0.08936866, 0.106371, 0.1183904, 0.09642985, 0.2353431, 
    0.2338847, 0.2644387, 0.2466882, 0.1717454, 0.1306368, 0.1729965, 
    0.1761341, 0.1277774, 0.1889131, 0.1913272, 0.1804239, 0.1804093, 
    0.2111473, 0.2756198, 0.2161311, 0.164975,
  0.2924396, 0.2902431, 0.2395903, 0.279888, 0.2873879, 0.3140104, 0.2614961, 
    0.2907968, 0.2508754, 0.2479896, 0.1569293, 0.01578703, 0.08073275, 
    0.1654402, 0.2840966, 0.2383517, 0.2460516, 0.3194532, 0.267639, 
    0.2424098, 0.2710357, 0.2169665, 0.1748251, 0.3007566, 0.1633528, 
    0.2177546, 0.22434, 0.2697715, 0.3001938,
  0.2132617, 0.2866074, 0.2815832, 0.2037793, 0.1937135, 0.2533509, 
    0.2794863, 0.2585777, 0.1762118, 0.1806992, 0.1055057, 0.1343027, 
    0.1779084, 0.2486546, 0.2571127, 0.2436191, 0.2534943, 0.2726222, 
    0.284305, 0.2333089, 0.1632058, 0.09270714, 0.1887731, 0.09122071, 
    0.09943171, 0.01603426, 0.02829282, 0.2052819, 0.1991989,
  0.2305958, 0.2314201, 0.215621, 0.1205551, 0.1032749, 0.077084, 0.1145639, 
    0.1159396, 0.1388528, 0.1399179, 0.1396872, 0.1466113, 0.1546081, 
    0.1542875, 0.1648948, 0.1428477, 0.1471769, 0.1503471, 0.1723146, 
    0.1917742, 0.1532626, 0.117373, 0.0572279, 0.01102954, 0.03714646, 
    0.008668871, 0.005100203, 0.06035037, 0.2242374,
  0.05202241, 0.05113681, 0.0502512, 0.04936559, 0.04847999, 0.04759439, 
    0.04670878, 0.0450895, 0.04469497, 0.04430044, 0.04390591, 0.04351138, 
    0.04311685, 0.04272232, 0.03942934, 0.04096131, 0.04249327, 0.04402523, 
    0.04555719, 0.04708915, 0.04862111, 0.05664004, 0.05638822, 0.05613639, 
    0.05588456, 0.05563273, 0.0553809, 0.05512908, 0.05273089,
  0.0896319, 0.01383123, 0.004113882, 0.01051191, 0.01843416, 0.005131719, 
    0.004677486, 0.0136809, 0.01354466, 0.009104768, 0.008707389, 0.02513546, 
    0.02983131, 0.1047356, 0.09730595, 0.1253494, 0.1552811, 0.2266136, 
    0.1611217, 0.1260798, 0.1206093, 0.1985443, 0.1955254, 0.110818, 
    0.09960767, 0.1173046, 0.1350081, 0.09759755, 0.087403,
  0.1103884, 0.2073278, 0.1834799, 0.2684265, 0.3240561, 0.2489357, 
    0.2723385, 0.2073739, 0.1428839, 0.1391465, 0.1159426, 0.0529201, 
    0.1791119, 0.1885383, 0.1987719, 0.201726, 0.1925406, 0.2280621, 
    0.1718644, 0.1973012, 0.1305914, 0.1837972, 0.2256116, 0.2896323, 
    0.2719988, 0.1830854, 0.2319497, 0.1009439, 0.09452356,
  0.143424, 0.2489844, 0.2778798, 0.2592641, 0.2196683, 0.199668, 0.2019007, 
    0.1671656, 0.2198004, 0.1772395, 0.2752507, 0.2790239, 0.2512833, 
    0.240906, 0.2376815, 0.2138429, 0.2004079, 0.2070907, 0.2484346, 
    0.2496036, 0.2988601, 0.2819123, 0.2746187, 0.2482415, 0.2491328, 
    0.2503997, 0.226647, 0.1502321, 0.1838883,
  0.1802093, 0.1618665, 0.1598629, 0.1868719, 0.163869, 0.1562766, 0.1557568, 
    0.1812011, 0.1634038, 0.166063, 0.1469018, 0.1429773, 0.1510561, 
    0.1512851, 0.1408442, 0.1027261, 0.08488442, 0.1047534, 0.11352, 
    0.1162902, 0.1274653, 0.1381024, 0.1591547, 0.134801, 0.08586608, 
    0.143337, 0.1391984, 0.1584706, 0.1719425,
  0.05793864, 0.026328, 0.02331553, 0.08865713, 0.06864595, 0.04319875, 
    0.09483044, 0.06801292, 0.04017957, 0.0240931, 0.07316657, 0.04143486, 
    0.05705836, 0.07539877, 0.06910647, 0.0879712, 0.06574313, 0.03751466, 
    0.0411251, 0.1141641, 0.09643625, 0.09093674, 0.03203597, 0.01530791, 
    0.07337285, 0.08584008, 0.1276088, 0.1040985, 0.07339151,
  0.005030812, -1.068436e-05, 0.08422144, 0.04229784, 0.07924078, 0.08091646, 
    0.07000431, 0.01068178, 0.0003179773, 0.002775666, 0.06271061, 
    0.07411035, 0.05559305, 0.03075848, 0.03302047, 0.04760781, 0.04575812, 
    0.1816523, 0.2076227, 0.04550786, 0.06531119, 0.002026092, 0.001307578, 
    0.001757464, 0.06155663, 0.07685291, 0.1196454, 0.02778672, 0.007456501,
  0.006311927, 0.08485681, 0.1067479, 0.02879847, 0.03552597, 0.01511426, 
    0.06758307, 0.02512265, 5.898027e-06, 7.573212e-05, 0.05027891, 
    0.03329977, 0.0140474, 0.01360062, 0.08088832, 0.07544515, 0.07309815, 
    0.08757947, 0.01148518, 0.002264379, 0.0002893113, 9.708852e-08, 
    9.395481e-06, 0.01494858, 0.1095213, 0.2202756, 0.02446294, 1.038589e-05, 
    1.218911e-06,
  0.007492094, 0.09328964, 0.1100602, 0.07175348, 0.1205796, 0.1096634, 
    0.09079599, 0.1022072, 0.01049612, 0.01922503, 0.0144099, 0.04521457, 
    0.03533911, 0.07731794, 0.06134417, 0.0459605, 0.03355204, 0.01354156, 
    0.001780644, 3.759857e-06, 3.350794e-08, -1.056127e-07, 0.003969118, 
    0.08830438, 0.2671681, 0.09579947, 0.003054157, 0.0003847973, 0.003824077,
  0.2652103, 0.02766384, 0.08778892, 0.0189515, 0.02619492, 0.03244006, 
    0.05516891, 0.05873241, 0.0401712, 0.1490613, 0.03886459, 0.01138798, 
    0.03647434, 0.04659229, 0.01702937, 0.004468503, 0.001160737, 
    0.001642843, -3.146155e-05, 9.615481e-05, 0.00879874, 0.01486236, 
    0.1189835, 0.1357732, 0.09658787, 0.0715574, 0.06993898, 0.04041082, 
    0.1065784,
  -3.085546e-05, 1.026763e-06, 0.009939821, 0.003663422, 0.01619558, 
    0.01065694, 0.000445744, 0.00436922, 0.04041878, 0.04667119, 0.1094118, 
    0.08619279, 0.04954384, 0.05296955, 0.05471691, 0.08358878, 0.09409252, 
    0.05558729, 0.09379669, 0.1272585, 0.108052, 0.01881271, 0.009807127, 
    0.009241159, 0.03290169, 0.0156328, 0.02061455, 0.007380946, 0.009750454,
  0.03296608, 6.198246e-06, 3.345053e-08, 2.660903e-05, 0.0008520944, 
    0.0008023478, 0.009434198, 0.001872485, 5.635793e-06, 0.05470793, 
    0.1093494, 0.02514372, 0.001214859, 0.007296773, 0.0008992929, 
    0.02774435, 0.03812168, 0.06360318, 0.05611075, 0.01151179, 0.0242243, 
    0.005057229, 0.002675479, 0.002739865, 0.03217356, 0.003329009, 
    0.01941889, 0.001305412, 0.03404712,
  0.01410047, 0.01896798, 0.01136929, 0.01876088, 0.02478525, 0.07697549, 
    0.05917059, 0.02707093, 0.112355, 0.06430026, 0.07761533, 0.07184797, 
    0.08927776, 0.07899322, 0.04442886, 0.1009887, 0.05829217, 0.06864797, 
    0.05515605, 0.0298335, 0.07089791, 0.06138469, 0.0425358, 0.02684358, 
    0.02301189, 0.04560613, 0.02650316, 0.005257635, 0.03281203,
  0.04607297, 0.03670185, 0.09839987, 0.2120256, 0.1355205, 0.1233737, 
    0.1653912, 0.1108199, 0.0735895, 0.1000697, 0.07710446, 0.08902455, 
    0.1018864, 0.1594482, 0.1529908, 0.1788377, 0.173573, 0.09450174, 
    0.07778372, 0.156929, 0.1135539, 0.05222449, 0.1532299, 0.1712398, 
    0.1675274, 0.1703038, 0.09856495, 0.07738936, 0.08336515,
  0.1486386, 0.1710545, 0.1963999, 0.2583089, 0.2237988, 0.2356993, 
    0.2480709, 0.1741744, 0.114071, 0.1076402, 0.1326614, 0.1071395, 
    0.2546281, 0.2327448, 0.2505825, 0.2404826, 0.1652093, 0.1290061, 
    0.1571536, 0.2215602, 0.1301441, 0.1898708, 0.1787624, 0.2054047, 
    0.186612, 0.2033423, 0.2803343, 0.1968771, 0.1592075,
  0.285901, 0.2861962, 0.2587053, 0.2627306, 0.2992354, 0.3235341, 0.2424728, 
    0.2707398, 0.2729607, 0.275875, 0.1994355, 0.05577573, 0.1457865, 
    0.2085029, 0.282252, 0.2366631, 0.2506242, 0.3174235, 0.3204538, 
    0.2329701, 0.2642885, 0.2143763, 0.1959174, 0.3374748, 0.1863086, 
    0.227716, 0.2171843, 0.265689, 0.3041822,
  0.2224069, 0.2709071, 0.2918666, 0.2157281, 0.223376, 0.2827719, 0.3433364, 
    0.3192428, 0.2272625, 0.2446802, 0.203889, 0.1925375, 0.2102292, 
    0.2709162, 0.2868707, 0.2443282, 0.2562021, 0.2848972, 0.2876065, 
    0.2327485, 0.1745087, 0.1123453, 0.2278863, 0.1170316, 0.1996114, 
    0.07746415, 0.07238957, 0.199349, 0.2137085,
  0.2243578, 0.2403536, 0.2034404, 0.1169093, 0.09729359, 0.09809584, 
    0.1311161, 0.1290706, 0.1495904, 0.2001931, 0.2117679, 0.2168602, 
    0.2173575, 0.2024235, 0.2013935, 0.157725, 0.1695813, 0.2015327, 
    0.2193725, 0.2072138, 0.172399, 0.1586723, 0.1213575, 0.05799027, 
    0.11503, 0.04196151, 0.05406696, 0.1670705, 0.2332881,
  0.07996757, 0.07746294, 0.0749583, 0.07245366, 0.06994903, 0.06744439, 
    0.06493975, 0.07823532, 0.07940403, 0.08057274, 0.08174144, 0.08291015, 
    0.08407885, 0.08524755, 0.07485828, 0.07748713, 0.08011597, 0.08274482, 
    0.08537368, 0.08800253, 0.09063137, 0.1082379, 0.106945, 0.105652, 
    0.1043591, 0.1030662, 0.1017733, 0.1004804, 0.08197128,
  0.1021045, 0.05916663, 0.00576089, 0.01868637, 0.0254067, 0.003920977, 
    0.01684357, 0.01990358, 0.0221001, 0.02707297, 0.04254844, 0.07109256, 
    0.06761558, 0.1038662, 0.09007208, 0.147043, 0.168467, 0.1999505, 
    0.1305292, 0.1504114, 0.1365414, 0.2732118, 0.1920688, 0.110048, 
    0.09351767, 0.1132975, 0.1301228, 0.09606848, 0.0828481,
  0.13229, 0.2295905, 0.1952304, 0.2898545, 0.4008349, 0.3038997, 0.2692415, 
    0.2569956, 0.1638721, 0.174246, 0.1555878, 0.09258564, 0.1878516, 
    0.1924974, 0.2024601, 0.2070361, 0.2004121, 0.24996, 0.2029093, 
    0.2000097, 0.1486722, 0.2226393, 0.2752452, 0.3317894, 0.2929282, 
    0.1795204, 0.2071424, 0.09090567, 0.09378716,
  0.1517107, 0.2404334, 0.3182174, 0.2687549, 0.2533996, 0.2005118, 
    0.2108878, 0.1679883, 0.229954, 0.1868152, 0.2992448, 0.2927257, 
    0.2640434, 0.2585982, 0.2177015, 0.2433335, 0.209631, 0.2142067, 
    0.2655134, 0.2724759, 0.3329093, 0.308691, 0.2985182, 0.2438515, 
    0.2669614, 0.2599841, 0.2428495, 0.1671633, 0.1927077,
  0.1984231, 0.1656151, 0.1513917, 0.1860236, 0.1709116, 0.1726259, 
    0.1591217, 0.1849777, 0.1597787, 0.181718, 0.1504808, 0.1486093, 
    0.150427, 0.1511066, 0.137077, 0.1058238, 0.08312081, 0.0955001, 
    0.107896, 0.1280377, 0.157885, 0.1513768, 0.150844, 0.1301519, 0.1017277, 
    0.1532013, 0.1362079, 0.1542386, 0.1754844,
  0.04755066, 0.02942427, 0.02066531, 0.08754008, 0.07410038, 0.04279719, 
    0.09540837, 0.08136454, 0.04124938, 0.02538908, 0.06043248, 0.03828467, 
    0.05732557, 0.07627353, 0.07206279, 0.08261512, 0.06779024, 0.03024525, 
    0.0389962, 0.1114423, 0.1003097, 0.07965424, 0.03284817, 0.01461582, 
    0.0864979, 0.08912463, 0.1295395, 0.1025138, 0.07342324,
  0.004153931, -2.975165e-07, 0.1074947, 0.04388633, 0.07854534, 0.07978171, 
    0.07168156, 0.006016521, 8.378006e-06, 0.006323192, 0.04118054, 
    0.06289808, 0.06984804, 0.0302888, 0.03987459, 0.03794644, 0.04069728, 
    0.1862931, 0.2168033, 0.04360082, 0.06794456, 0.0009508683, 0.0008861895, 
    0.002171997, 0.07557093, 0.08723409, 0.1148388, 0.02559377, 0.01169764,
  0.004198059, 0.1149352, 0.1304028, 0.03423661, 0.0364648, 0.02353999, 
    0.07281311, 0.02736684, 6.533959e-06, 0.001051999, 0.05934609, 
    0.04797768, 0.01639698, 0.01895581, 0.08556789, 0.09832616, 0.07338153, 
    0.09525534, 0.01833133, 0.003705619, 8.870784e-07, 4.755922e-08, 
    6.231588e-06, 0.01344662, 0.1356272, 0.2472993, 0.02681347, 4.295437e-05, 
    5.110556e-06,
  0.009995899, 0.1187449, 0.147599, 0.09391537, 0.1351723, 0.1125923, 
    0.1068646, 0.1163397, 0.01468183, 0.02522548, 0.0199863, 0.05248763, 
    0.04028841, 0.08633596, 0.07809041, 0.04799552, 0.031425, 0.02414637, 
    0.005276897, 0.0001287015, 2.460614e-08, -1.033132e-05, 0.00472215, 
    0.123479, 0.3082662, 0.1064265, 0.004036723, 3.113734e-05, 0.005559793,
  0.2760472, 0.04783653, 0.1049939, 0.02069074, 0.03084143, 0.03584553, 
    0.06748916, 0.08112587, 0.07284396, 0.1786143, 0.04294339, 0.0141942, 
    0.04607331, 0.05411356, 0.02065408, 0.006663921, -5.925449e-06, 
    0.0003932733, -1.593966e-05, 0.002795651, 0.01018943, 0.02266061, 
    0.1586471, 0.1727753, 0.1273535, 0.07460482, 0.07151433, 0.04286378, 
    0.08377077,
  6.21761e-07, 3.531462e-06, 0.002475312, 0.003830701, 0.01774282, 
    0.01546919, 0.001334052, 0.007662349, 0.04637385, 0.05271303, 0.1298278, 
    0.09371148, 0.0548867, 0.05340465, 0.06668077, 0.08833167, 0.08780798, 
    0.06798415, 0.09853339, 0.1265064, 0.1202315, 0.02082481, 0.01659164, 
    0.01269056, 0.0433368, 0.0149812, 0.01681756, 0.003798683, 0.004246241,
  0.01399366, 3.515794e-06, 7.944354e-08, 0.0003817661, 0.005828904, 
    0.003509276, 0.0118076, 0.004119661, 1.473412e-05, 0.06343936, 0.1315159, 
    0.0345204, 0.00229717, 0.008629272, 0.001459378, 0.02940474, 0.03985943, 
    0.06922439, 0.05032333, 0.009245766, 0.02667009, 0.009762606, 
    0.002859761, 0.004714926, 0.03309329, 0.005815024, 0.01796422, 
    -1.486716e-05, 0.02542982,
  0.003016517, 0.01432791, 0.005897151, 0.01902824, 0.0276363, 0.08176103, 
    0.0500591, 0.03698158, 0.1378449, 0.09230497, 0.07857495, 0.06763607, 
    0.08513542, 0.08383138, 0.05385324, 0.1036661, 0.0612575, 0.06370325, 
    0.05230324, 0.03026888, 0.07237552, 0.06372529, 0.04546839, 0.02357028, 
    0.03101247, 0.05111456, 0.03157304, 0.01015544, 0.04172119,
  0.04158445, 0.03658312, 0.1134687, 0.2195894, 0.1304494, 0.1168947, 
    0.1818815, 0.09375724, 0.05586861, 0.0954885, 0.05821756, 0.08562459, 
    0.1103191, 0.1510748, 0.1545761, 0.1637918, 0.1635611, 0.08307672, 
    0.0842756, 0.1580349, 0.1312592, 0.05238733, 0.1460269, 0.1721534, 
    0.1664878, 0.1744801, 0.1022813, 0.08107179, 0.08796108,
  0.1511599, 0.1804313, 0.1868457, 0.2488975, 0.2062905, 0.2206209, 
    0.2433213, 0.1735228, 0.1296514, 0.1015805, 0.1275919, 0.1084589, 
    0.2489233, 0.2229171, 0.246044, 0.2188057, 0.1637707, 0.1227466, 
    0.1652166, 0.2523707, 0.1390363, 0.1803087, 0.1760506, 0.2016958, 
    0.1816932, 0.2001111, 0.2888671, 0.1997177, 0.1661954,
  0.2910074, 0.2879516, 0.2697839, 0.2642909, 0.2777781, 0.3094718, 
    0.2282511, 0.2994052, 0.2638968, 0.3065528, 0.2259195, 0.09638341, 
    0.1882304, 0.2230956, 0.2752076, 0.2541508, 0.222775, 0.3208058, 
    0.3090172, 0.2349665, 0.2680833, 0.2070225, 0.2238944, 0.3656813, 
    0.2087186, 0.2177947, 0.2132773, 0.2510383, 0.2930214,
  0.2198241, 0.2713992, 0.2850045, 0.2348088, 0.2554233, 0.3052373, 
    0.3619282, 0.3897554, 0.2410403, 0.2533687, 0.2647057, 0.201519, 
    0.2705941, 0.3171684, 0.3041767, 0.2371103, 0.2579052, 0.2934829, 
    0.3136047, 0.2383481, 0.2039842, 0.1570156, 0.2376382, 0.1552457, 
    0.2281817, 0.1519483, 0.1444417, 0.1920563, 0.2092749,
  0.2220993, 0.2412587, 0.1847185, 0.1147025, 0.09307003, 0.1041139, 
    0.1348143, 0.1327731, 0.1579361, 0.1976014, 0.2068326, 0.2388927, 
    0.214684, 0.2217858, 0.2019719, 0.1649378, 0.1612062, 0.2243488, 
    0.2986585, 0.2807831, 0.2133139, 0.2151776, 0.2027711, 0.06675321, 
    0.1576611, 0.07719992, 0.06905661, 0.1888265, 0.2451775,
  0.1135352, 0.1123481, 0.111161, 0.1099739, 0.1087869, 0.1075998, 0.1064127, 
    0.1131338, 0.1135091, 0.1138845, 0.1142598, 0.1146351, 0.1150105, 
    0.1153858, 0.1135336, 0.1160699, 0.1186062, 0.1211425, 0.1236788, 
    0.1262151, 0.1287514, 0.125526, 0.1238015, 0.1220769, 0.1203524, 
    0.1186278, 0.1169033, 0.1151787, 0.1144848,
  0.102823, 0.1120222, 0.06667099, 0.04531994, 0.04236373, 0.02070287, 
    0.02597528, 0.03218425, 0.04691374, 0.07471089, 0.08852618, 0.1258591, 
    0.1323013, 0.09063335, 0.1007977, 0.1564705, 0.1734187, 0.1798961, 
    0.1099793, 0.1328618, 0.1310686, 0.2766935, 0.197015, 0.1084002, 
    0.07985306, 0.1227804, 0.1309883, 0.09179486, 0.08626509,
  0.1430512, 0.2496369, 0.2144826, 0.333984, 0.4276903, 0.3266804, 0.2738039, 
    0.2643484, 0.2071888, 0.1844725, 0.1349015, 0.1179581, 0.1979062, 
    0.1810127, 0.2077946, 0.2124669, 0.2471948, 0.2428064, 0.2039865, 
    0.191693, 0.1970096, 0.2052798, 0.2580823, 0.352354, 0.2803565, 
    0.1894286, 0.1809594, 0.0924364, 0.0671266,
  0.2130675, 0.2620663, 0.3237104, 0.3063333, 0.2981721, 0.2801088, 
    0.2811581, 0.2243336, 0.2263201, 0.213021, 0.2793505, 0.2911205, 
    0.2608035, 0.2621133, 0.2174358, 0.2402544, 0.2054034, 0.205797, 
    0.2660796, 0.277676, 0.3427637, 0.2760949, 0.2995754, 0.2660683, 0.27872, 
    0.2665493, 0.2421195, 0.2109281, 0.2395201,
  0.1968859, 0.1812232, 0.1582789, 0.1911618, 0.1639667, 0.1639098, 
    0.1575194, 0.1929953, 0.1794094, 0.1676928, 0.1543157, 0.156789, 
    0.1595085, 0.1472861, 0.1300212, 0.1046135, 0.09060346, 0.09948061, 
    0.1173778, 0.1427119, 0.1644647, 0.1568745, 0.1419149, 0.1275564, 
    0.1280057, 0.1495375, 0.1316039, 0.16059, 0.1884558,
  0.05736528, 0.03219049, 0.02262028, 0.07962858, 0.08696249, 0.04111934, 
    0.09487511, 0.08962619, 0.04353996, 0.02783517, 0.04879014, 0.04018822, 
    0.06302053, 0.08454549, 0.08097959, 0.08744002, 0.07749409, 0.03354433, 
    0.05116227, 0.120219, 0.1049216, 0.0880377, 0.04154506, 0.01673681, 
    0.09562515, 0.08445998, 0.1243222, 0.1024581, 0.07110429,
  0.006357502, -2.333633e-07, 0.1153083, 0.04625076, 0.08097682, 0.08100717, 
    0.07200796, 0.00223129, 9.19747e-06, 0.004063797, 0.02027717, 0.05559409, 
    0.07813521, 0.03240718, 0.0523502, 0.04414261, 0.0364456, 0.1899311, 
    0.2153247, 0.04074766, 0.08000983, 0.001236714, 6.656578e-05, 
    0.002448865, 0.07977502, 0.09237968, 0.1198272, 0.02691658, 0.02045601,
  0.002278791, 0.1132966, 0.1675693, 0.02879961, 0.03855978, 0.02042634, 
    0.07415236, 0.02370608, 5.267225e-06, 0.001384519, 0.06459872, 
    0.06312152, 0.01282668, 0.02445879, 0.0841196, 0.07508221, 0.06083532, 
    0.09586722, 0.01738817, 0.009120161, 0.000242071, 1.797536e-08, 
    5.827426e-06, 0.004758306, 0.1211527, 0.2795925, 0.02201543, 
    0.0002688828, 1.25632e-05,
  0.00930338, 0.08132183, 0.2012596, 0.1039124, 0.1145093, 0.1069652, 
    0.1002109, 0.1051365, 0.01348763, 0.01730881, 0.02839526, 0.03400696, 
    0.03354173, 0.0629085, 0.0607643, 0.04522218, 0.0329981, 0.03666566, 
    0.004950424, 0.0004876681, 9.682034e-08, 7.371732e-08, 0.002209799, 
    0.1230809, 0.3032324, 0.1206473, 0.006294453, 3.330408e-06, 0.001757854,
  0.2606178, 0.08248673, 0.1228299, 0.03453203, 0.03628677, 0.03448205, 
    0.07244516, 0.07394356, 0.10077, 0.1979713, 0.04198349, 0.01111551, 
    0.02842363, 0.04527463, 0.01800377, 0.002940462, 0.00048041, 
    0.0001593728, 2.311532e-05, -8.143703e-06, 0.008895466, 0.0168603, 
    0.1836429, 0.1954134, 0.1318937, 0.07308062, 0.07041534, 0.04740591, 
    0.07887094,
  -4.912373e-06, 2.052305e-06, 0.006693279, 0.01253769, 0.0198486, 
    0.01848175, 0.001864818, 0.004175345, 0.05014866, 0.04666035, 0.1288228, 
    0.08090162, 0.0505322, 0.05341823, 0.06110891, 0.07633179, 0.07733556, 
    0.08037211, 0.1115784, 0.1247417, 0.1166462, 0.02298116, 0.02862331, 
    0.01398504, 0.04642902, 0.01453979, 0.01156595, 0.0024975, 0.0002147976,
  0.0004169498, 1.038017e-06, 5.288978e-07, 0.00203746, 0.01381033, 
    0.004107946, 0.01437659, 0.01280883, 9.427132e-05, 0.06090039, 0.1425822, 
    0.0342454, 0.003375279, 0.007967692, 0.002984334, 0.03328883, 0.04610756, 
    0.07158005, 0.05635455, 0.01417575, 0.02797718, 0.01456833, 0.005478282, 
    0.008696175, 0.04066056, 0.0141374, 0.01884069, 0.001069739, 0.01756652,
  0.0001313892, 0.008948341, 0.006548323, 0.02871636, 0.03967436, 0.0858627, 
    0.05287339, 0.05553148, 0.1560115, 0.116811, 0.08755977, 0.06393977, 
    0.07828106, 0.08785239, 0.06422544, 0.1202758, 0.0692883, 0.06121256, 
    0.05581817, 0.03044086, 0.08524119, 0.06970774, 0.05043534, 0.02290254, 
    0.04053485, 0.05547934, 0.03822371, 0.01257577, 0.03139399,
  0.03887664, 0.03742961, 0.1429914, 0.231395, 0.1350789, 0.1204159, 
    0.188907, 0.07102241, 0.04614074, 0.08707847, 0.05090333, 0.08521684, 
    0.1124011, 0.1527724, 0.1477078, 0.1645592, 0.1566605, 0.07701097, 
    0.08148063, 0.1682077, 0.1466674, 0.05683257, 0.1492283, 0.1751626, 
    0.1819895, 0.1735955, 0.1056523, 0.07845414, 0.09371363,
  0.156656, 0.1843572, 0.1887293, 0.2468752, 0.1943362, 0.2064265, 0.2153072, 
    0.1745421, 0.1406034, 0.08727883, 0.1227092, 0.105904, 0.2427937, 
    0.207105, 0.2481918, 0.2343695, 0.1713206, 0.1300689, 0.1836339, 
    0.2659957, 0.137954, 0.1740205, 0.1891442, 0.2226631, 0.1932081, 
    0.2024075, 0.2889818, 0.1985024, 0.173874,
  0.2922944, 0.3140968, 0.2981221, 0.2613392, 0.3089532, 0.3064989, 
    0.2375608, 0.2988857, 0.2606692, 0.3274217, 0.2889604, 0.1025744, 
    0.2319453, 0.2183447, 0.2679912, 0.2562439, 0.2316171, 0.3188311, 
    0.3032886, 0.2640678, 0.272788, 0.2169302, 0.2122884, 0.3488674, 
    0.2180075, 0.2212807, 0.224992, 0.2596409, 0.3079671,
  0.242507, 0.2765839, 0.2977994, 0.2517418, 0.2526733, 0.3357027, 0.3731539, 
    0.4051069, 0.2681862, 0.2812075, 0.2810463, 0.2316427, 0.2805614, 
    0.329214, 0.3362851, 0.2306263, 0.2388722, 0.3036882, 0.3210658, 
    0.2622127, 0.2318171, 0.1799745, 0.2710753, 0.1753382, 0.2177761, 
    0.2103171, 0.2241004, 0.2135311, 0.2204047,
  0.229394, 0.2441579, 0.1590965, 0.1181538, 0.1066085, 0.1215079, 0.1433099, 
    0.1660378, 0.165099, 0.2253454, 0.2171169, 0.2356302, 0.209301, 
    0.2352708, 0.2273723, 0.1745018, 0.1635926, 0.2276265, 0.3054597, 
    0.2922004, 0.2655995, 0.2854491, 0.2340063, 0.07071179, 0.1591621, 
    0.09122045, 0.1074945, 0.2136999, 0.2598097,
  0.1220157, 0.123149, 0.1242823, 0.1254156, 0.1265488, 0.1276821, 0.1288154, 
    0.1366473, 0.1380062, 0.1393651, 0.140724, 0.142083, 0.1434419, 
    0.1448008, 0.1518269, 0.1542243, 0.1566217, 0.1590191, 0.1614165, 
    0.1638139, 0.1662112, 0.1522934, 0.1474038, 0.1425142, 0.1376246, 
    0.132735, 0.1278454, 0.1229558, 0.1211091,
  0.09415144, 0.1177171, 0.10244, 0.08981159, 0.0782023, 0.0632189, 
    0.04258578, 0.03779361, 0.1035128, 0.143777, 0.1213166, 0.1470095, 
    0.1541415, 0.08250547, 0.09326877, 0.1091531, 0.1475337, 0.1729719, 
    0.1028805, 0.1205637, 0.1274486, 0.2822462, 0.1916169, 0.1030907, 
    0.07607668, 0.1092646, 0.1279252, 0.09156474, 0.09450655,
  0.1388752, 0.2556554, 0.2467628, 0.3478662, 0.4342235, 0.3384295, 0.258496, 
    0.287752, 0.2037182, 0.1679353, 0.1230584, 0.1193908, 0.2095343, 
    0.1923589, 0.2358227, 0.2297501, 0.2578981, 0.3086796, 0.2385341, 
    0.2906092, 0.1827538, 0.2483689, 0.287578, 0.3968781, 0.2703846, 
    0.2593747, 0.1699851, 0.1476559, 0.07615348,
  0.3340821, 0.3494673, 0.4357777, 0.3843141, 0.3424838, 0.298653, 0.3118936, 
    0.2264276, 0.2667732, 0.2370181, 0.3540885, 0.2866892, 0.2859738, 
    0.2558481, 0.2223389, 0.2271254, 0.2144456, 0.2247354, 0.3004345, 
    0.284684, 0.3189643, 0.2725639, 0.3040286, 0.2419872, 0.2774742, 
    0.2686346, 0.270042, 0.2365783, 0.2971174,
  0.2082125, 0.1923781, 0.1561375, 0.1938199, 0.1737733, 0.1637562, 
    0.1605007, 0.2077878, 0.1935665, 0.1881624, 0.1693514, 0.1484567, 
    0.1644247, 0.1394046, 0.1263116, 0.1155343, 0.09387951, 0.1026022, 
    0.1161204, 0.1480971, 0.166463, 0.1508823, 0.1356805, 0.1281471, 
    0.1172737, 0.1401679, 0.1259116, 0.1459154, 0.1715237,
  0.0691057, 0.03225962, 0.02422489, 0.06563377, 0.0888799, 0.04689825, 
    0.101616, 0.095565, 0.05822147, 0.0278487, 0.03792583, 0.04120694, 
    0.05550603, 0.1074084, 0.09171103, 0.0901407, 0.08257578, 0.04289475, 
    0.05851223, 0.1314062, 0.1134486, 0.09998351, 0.05698406, 0.02112678, 
    0.07548963, 0.088562, 0.1192697, 0.1098156, 0.07798579,
  0.007046002, -1.623598e-08, 0.1206408, 0.04773967, 0.09052394, 0.08201282, 
    0.06579033, 0.001123758, 4.468822e-06, 0.001272452, 0.006050777, 
    0.0301989, 0.08300671, 0.0360605, 0.07308406, 0.05093765, 0.03740682, 
    0.2036672, 0.2104195, 0.03483327, 0.09724182, 0.003127841, 8.861191e-06, 
    0.001965172, 0.05373757, 0.09753315, 0.1326365, 0.03575578, 0.01353379,
  0.0005876971, 0.07566146, 0.1702534, 0.0222586, 0.04135582, 0.02107871, 
    0.0697374, 0.01741275, 2.439982e-06, 0.0009531783, 0.05044565, 
    0.04943997, 0.01426755, 0.02970313, 0.09166443, 0.05367639, 0.0530863, 
    0.07087004, 0.02463047, 0.01764917, 0.003065023, 1.180505e-08, 
    3.687876e-06, 0.001582142, 0.1113286, 0.2964025, 0.0141807, 0.0001256033, 
    1.288899e-05,
  0.003062131, 0.02865521, 0.2246763, 0.09017271, 0.1014153, 0.09457511, 
    0.09045848, 0.0940506, 0.0130767, 0.01359136, 0.0255018, 0.0266524, 
    0.03074221, 0.05627289, 0.05009475, 0.04640614, 0.03065828, 0.04455366, 
    0.007012675, 0.0002549264, -1.346547e-07, -6.290048e-07, 0.001054846, 
    0.08485707, 0.2036391, 0.1021864, 0.007026669, -2.15337e-06, 5.185686e-05,
  0.2290493, 0.08596136, 0.1081889, 0.04799325, 0.03954861, 0.0316697, 
    0.06628233, 0.06829118, 0.1003394, 0.1729403, 0.03953752, 0.009727955, 
    0.01936293, 0.04071323, 0.01520882, 0.002050069, 0.004949414, 
    -4.211512e-06, 7.344112e-05, 0.0005948232, 0.006755047, 0.01085672, 
    0.159821, 0.1703814, 0.1222095, 0.05626482, 0.07602772, 0.03962241, 
    0.06940441,
  2.425276e-06, 1.599345e-05, 0.001842805, 0.05196567, 0.02585456, 
    0.01584472, 0.004479466, 0.005045491, 0.05164043, 0.04311696, 0.1308843, 
    0.07196615, 0.04873833, 0.05517481, 0.05909187, 0.06135004, 0.07319873, 
    0.09150362, 0.1067085, 0.1178891, 0.1066386, 0.02649408, 0.04669414, 
    0.0196955, 0.05449152, 0.01187065, 0.004790875, 0.0003394786, 0.0004257692,
  3.763994e-05, 5.283166e-07, 4.606623e-07, 0.004715206, 0.01794248, 
    8.346033e-05, 0.01471584, 0.01882847, 0.004405664, 0.04420684, 0.1517157, 
    0.0351745, 0.004105476, 0.007311225, 0.005809018, 0.03506906, 0.04453801, 
    0.08459004, 0.06309673, 0.01699547, 0.01403849, 0.0256134, 0.01007419, 
    0.01993893, 0.04921551, 0.01878493, 0.01105755, 0.001096909, 0.006426232,
  5.559642e-05, 0.00738477, 0.005383072, 0.03098631, 0.05896833, 0.09053439, 
    0.05292591, 0.06306869, 0.1616442, 0.1289503, 0.08424981, 0.05657173, 
    0.0786934, 0.09832767, 0.08101774, 0.1466107, 0.07766716, 0.06707792, 
    0.06951318, 0.03804163, 0.09846811, 0.0823964, 0.04245772, 0.02784098, 
    0.05199951, 0.06043315, 0.04293662, 0.01508413, 0.02118126,
  0.03832944, 0.0431568, 0.1381391, 0.2589929, 0.1389283, 0.1179526, 
    0.2025231, 0.05628118, 0.04058872, 0.07838254, 0.04786517, 0.08477259, 
    0.1222797, 0.1495046, 0.1550238, 0.166311, 0.1615097, 0.08417921, 
    0.08675767, 0.1876919, 0.1569436, 0.06334237, 0.1466191, 0.1700962, 
    0.1911383, 0.1908723, 0.1176385, 0.09050511, 0.09921796,
  0.1557533, 0.1920927, 0.1747932, 0.2185557, 0.2053659, 0.2255927, 
    0.2196009, 0.1809159, 0.1350964, 0.07908393, 0.1142763, 0.09761357, 
    0.2446243, 0.2260876, 0.2534407, 0.233218, 0.1722056, 0.1341338, 
    0.1801905, 0.2778729, 0.170005, 0.1591656, 0.1949281, 0.2632232, 
    0.1948853, 0.2108211, 0.3087671, 0.1935273, 0.1746751,
  0.275535, 0.3132443, 0.2768418, 0.2811409, 0.3451913, 0.3482946, 0.2567362, 
    0.2920557, 0.2448523, 0.3292714, 0.3109531, 0.1040014, 0.2431035, 
    0.234102, 0.2684922, 0.2625882, 0.226034, 0.3316302, 0.2903723, 
    0.2567622, 0.2837917, 0.2081273, 0.2667325, 0.3756181, 0.2244785, 
    0.2324778, 0.2388587, 0.2712067, 0.3090302,
  0.2538099, 0.2992533, 0.3034419, 0.3173853, 0.2858189, 0.4502052, 
    0.4875557, 0.4352327, 0.2967914, 0.2781447, 0.3132464, 0.2356792, 
    0.3030206, 0.338316, 0.3626186, 0.2401051, 0.2362326, 0.3221212, 
    0.3217902, 0.2931057, 0.2516125, 0.1735103, 0.2971298, 0.2200188, 
    0.2100882, 0.2455848, 0.3078702, 0.2917272, 0.2356943,
  0.2667305, 0.2469459, 0.1885528, 0.1563557, 0.1389084, 0.1537825, 
    0.1927572, 0.2416805, 0.2203338, 0.2888941, 0.2423442, 0.267682, 
    0.2697406, 0.2617334, 0.2646441, 0.2222066, 0.1747004, 0.2435014, 
    0.3208488, 0.302557, 0.2623088, 0.3140917, 0.2550669, 0.08343881, 
    0.136379, 0.1193822, 0.1341889, 0.2300212, 0.3041426,
  0.1189404, 0.1198753, 0.1208104, 0.1217453, 0.1226803, 0.1236153, 
    0.1245503, 0.1252275, 0.128934, 0.1326406, 0.1363471, 0.1400537, 
    0.1437603, 0.1474668, 0.1512745, 0.1519526, 0.1526307, 0.1533089, 
    0.153987, 0.1546651, 0.1553432, 0.1469314, 0.1416117, 0.136292, 
    0.1309724, 0.1256527, 0.120333, 0.1150133, 0.1181924,
  0.08492156, 0.1122582, 0.1114361, 0.1113092, 0.1160421, 0.1100642, 
    0.07581764, 0.08755634, 0.1491563, 0.1479659, 0.130733, 0.1485797, 
    0.1455348, 0.08015651, 0.06387258, 0.06316884, 0.1139313, 0.1509567, 
    0.09299931, 0.1343951, 0.1325087, 0.270849, 0.1922048, 0.09229319, 
    0.1141075, 0.1587389, 0.1420092, 0.09798084, 0.09445705,
  0.1290541, 0.3145441, 0.2607027, 0.3406586, 0.4268564, 0.3669813, 
    0.2746546, 0.2848851, 0.2018326, 0.1668989, 0.1192349, 0.1235267, 
    0.2340865, 0.2156444, 0.2495823, 0.2670701, 0.35059, 0.3450212, 0.300344, 
    0.339098, 0.30075, 0.3487028, 0.3265274, 0.4249795, 0.2803861, 0.2168597, 
    0.1557431, 0.1383934, 0.09500982,
  0.3870786, 0.4165187, 0.4691623, 0.4370539, 0.3715401, 0.3336242, 
    0.3562184, 0.2743087, 0.3156264, 0.2867795, 0.3648339, 0.3051772, 
    0.3044747, 0.274963, 0.250815, 0.2547928, 0.2472707, 0.2609102, 
    0.3237536, 0.3356509, 0.3809217, 0.2800554, 0.2840756, 0.2722637, 
    0.2832419, 0.2677409, 0.2512708, 0.2351231, 0.3601154,
  0.2324295, 0.1862596, 0.1584001, 0.2060567, 0.1689345, 0.1740709, 
    0.1695652, 0.2029552, 0.1905355, 0.2096764, 0.1899692, 0.1693796, 
    0.1776612, 0.1399053, 0.1316367, 0.1403259, 0.09824872, 0.119394, 
    0.1430497, 0.1538012, 0.1799114, 0.1514849, 0.1500927, 0.1466404, 
    0.108026, 0.1325526, 0.1284076, 0.1535482, 0.191621,
  0.07509089, 0.03933702, 0.03064833, 0.06818454, 0.1046761, 0.06241624, 
    0.1237796, 0.1125402, 0.06905465, 0.03532956, 0.03401376, 0.04149918, 
    0.05158112, 0.1053467, 0.1069886, 0.09605863, 0.09786636, 0.05268907, 
    0.0703532, 0.1400521, 0.1124054, 0.1164295, 0.07404412, 0.02482382, 
    0.05255486, 0.09612852, 0.1217112, 0.1162266, 0.08496988,
  0.01403332, -1.508322e-08, 0.1133653, 0.04414619, 0.06479126, 0.08294917, 
    0.06391466, 0.00804179, 2.036654e-05, 0.0001162122, 0.00121705, 
    0.01592956, 0.06577142, 0.03825834, 0.06629109, 0.05894121, 0.04186286, 
    0.2032156, 0.1555892, 0.02946536, 0.1030296, 0.006704913, 2.432674e-06, 
    0.001160683, 0.03542321, 0.09488906, 0.1190451, 0.03842711, 0.01359189,
  2.555802e-05, 0.04625008, 0.1316879, 0.02017222, 0.04787158, 0.02749971, 
    0.07225845, 0.01538955, 2.686191e-05, 3.102078e-05, 0.03767795, 
    0.03538137, 0.02416999, 0.02965811, 0.09248346, 0.04838046, 0.04930773, 
    0.05464914, 0.03420283, 0.0432438, 0.01062068, -1.469101e-07, 
    2.474081e-06, 0.0009412831, 0.1056641, 0.2656969, 0.0143909, 
    0.0005857837, 1.502566e-05,
  0.000512588, 0.01304471, 0.1773134, 0.08478554, 0.09248947, 0.09028076, 
    0.09106456, 0.08765925, 0.01205753, 0.01031169, 0.0233939, 0.02324967, 
    0.02945927, 0.05441834, 0.04502124, 0.04928406, 0.03401481, 0.05714311, 
    0.01688144, 0.001210741, 1.110453e-06, 6.471108e-08, 0.0005926398, 
    0.07953729, 0.1644732, 0.08667653, 0.008565385, 2.286689e-07, 0.000506852,
  0.1958107, 0.07438495, 0.1041615, 0.06576359, 0.04912435, 0.0335015, 
    0.06350272, 0.06152027, 0.11437, 0.1604048, 0.0371989, 0.008703196, 
    0.01918576, 0.03637619, 0.0182666, 0.002238571, 0.002774062, 
    -0.0002009158, 0.0004013002, 0.0009935441, 0.004811567, 0.01267039, 
    0.1244286, 0.1613882, 0.1245526, 0.04381843, 0.08490573, 0.03867565, 
    0.06810389,
  5.54271e-07, 0.0002401902, 0.01194645, 0.0986663, 0.03174265, 0.0152997, 
    0.005734987, 0.007099208, 0.05468767, 0.04773306, 0.1414853, 0.07068709, 
    0.05337945, 0.06026788, 0.06745329, 0.05421554, 0.06723636, 0.09577392, 
    0.1036692, 0.1113568, 0.0938888, 0.03451492, 0.05827925, 0.02616805, 
    0.06020886, 0.01319822, 0.002540431, 1.634868e-05, 0.0003369678,
  4.487333e-05, 4.261783e-07, 2.214787e-07, 0.01053821, 0.03529958, 
    0.001654464, 0.01075504, 0.02703233, 0.009621418, 0.07124387, 0.1446671, 
    0.03720326, 0.006483301, 0.009385394, 0.01520583, 0.02986773, 0.04017594, 
    0.09607439, 0.0614457, 0.01836149, 0.01258867, 0.05433779, 0.0181373, 
    0.03238915, 0.05190799, 0.02975055, 0.01518364, 0.003760847, 0.0003078097,
  4.658693e-06, 0.007933155, 0.0127966, 0.03617868, 0.07557368, 0.09489997, 
    0.05504513, 0.06581461, 0.161073, 0.1414708, 0.08306114, 0.05591298, 
    0.08786422, 0.1035632, 0.09677751, 0.1576439, 0.1012998, 0.07442206, 
    0.09646138, 0.0520911, 0.1147228, 0.07994102, 0.04101294, 0.03280967, 
    0.05640477, 0.06268853, 0.04769929, 0.02853772, 0.01856867,
  0.04669127, 0.05628585, 0.1534762, 0.3017461, 0.1611173, 0.09374978, 
    0.1970937, 0.04267405, 0.03639629, 0.07989009, 0.04659234, 0.09548488, 
    0.1500729, 0.1594875, 0.1560568, 0.1688343, 0.1701041, 0.111563, 
    0.09685929, 0.2047144, 0.1605635, 0.05054573, 0.1442842, 0.1828776, 
    0.212317, 0.2102177, 0.1379101, 0.1097467, 0.1099997,
  0.1674795, 0.1949005, 0.1809479, 0.2288086, 0.222767, 0.2414875, 0.2183861, 
    0.1884522, 0.1270819, 0.07579827, 0.1087874, 0.08973318, 0.2590826, 
    0.2605551, 0.2648423, 0.2380079, 0.1931895, 0.1454595, 0.1827571, 
    0.2954588, 0.177588, 0.1491974, 0.2109793, 0.2584655, 0.1806597, 
    0.2143024, 0.3223979, 0.204293, 0.1872823,
  0.2550057, 0.3269963, 0.2901822, 0.290859, 0.3564136, 0.3856699, 0.2809117, 
    0.299304, 0.2612195, 0.3327388, 0.3367639, 0.1139021, 0.2577187, 
    0.2299798, 0.2636248, 0.2738945, 0.2318805, 0.3400606, 0.2937517, 
    0.2930277, 0.2742483, 0.2091509, 0.3011014, 0.3801563, 0.2116252, 
    0.2457366, 0.2609195, 0.2789935, 0.3109347,
  0.2758795, 0.2792723, 0.3735774, 0.3433291, 0.3054576, 0.4513979, 
    0.4704512, 0.4808969, 0.2870031, 0.2864527, 0.3180132, 0.2444232, 
    0.3137886, 0.3425819, 0.3750326, 0.22583, 0.2199937, 0.3375669, 
    0.3002081, 0.2924207, 0.2679374, 0.1905701, 0.3001891, 0.2340868, 
    0.2064658, 0.2653002, 0.3512689, 0.3382618, 0.2576896,
  0.2536831, 0.2769891, 0.2416009, 0.2247754, 0.2069513, 0.1911867, 
    0.2005134, 0.2528077, 0.2271621, 0.2758196, 0.2957827, 0.3223587, 
    0.3320413, 0.2817203, 0.2663787, 0.2285904, 0.185654, 0.239763, 
    0.3328605, 0.3292444, 0.2790435, 0.3118004, 0.2735959, 0.09288199, 
    0.1355984, 0.1249086, 0.1560699, 0.2395742, 0.3185809,
  0.1143611, 0.1148742, 0.1153872, 0.1159003, 0.1164133, 0.1169264, 
    0.1174395, 0.1231092, 0.1272012, 0.1312932, 0.1353851, 0.1394771, 
    0.1435691, 0.1476611, 0.146203, 0.1462979, 0.1463929, 0.1464878, 
    0.1465828, 0.1466777, 0.1467726, 0.1341445, 0.1294445, 0.1247445, 
    0.1200445, 0.1153446, 0.1106446, 0.1059446, 0.1139506,
  0.07593368, 0.1018048, 0.120947, 0.1194392, 0.1506791, 0.1264719, 
    0.1100621, 0.127224, 0.1687818, 0.1361468, 0.1323675, 0.1418378, 
    0.1417232, 0.05248929, 0.045249, 0.08368562, 0.07741837, 0.1328715, 
    0.09574699, 0.1176519, 0.1322275, 0.2817344, 0.2158348, 0.1190223, 
    0.1127118, 0.1691098, 0.1532954, 0.09896622, 0.09176733,
  0.1090299, 0.2039505, 0.2277321, 0.3073503, 0.4252549, 0.37173, 0.2707313, 
    0.2664508, 0.1839017, 0.1697568, 0.1241011, 0.1232597, 0.2379615, 
    0.1525552, 0.2499114, 0.2650569, 0.3066334, 0.3030117, 0.2856907, 
    0.3099935, 0.2215513, 0.2778295, 0.3787466, 0.4259702, 0.2581702, 
    0.203916, 0.1609926, 0.1590795, 0.1055036,
  0.270828, 0.3544426, 0.3790031, 0.4356322, 0.358297, 0.3344193, 0.3537982, 
    0.2937078, 0.3288524, 0.293328, 0.3609815, 0.3122864, 0.3237416, 
    0.3054899, 0.2555099, 0.258821, 0.2557542, 0.3089901, 0.3335215, 
    0.3336875, 0.35098, 0.2834837, 0.2856985, 0.2624374, 0.2972386, 
    0.2449889, 0.2401205, 0.2511316, 0.2811359,
  0.2390148, 0.1979231, 0.184368, 0.1948736, 0.1708179, 0.1856803, 0.1727777, 
    0.2165849, 0.2300598, 0.2368319, 0.2066507, 0.1792509, 0.1970149, 
    0.149496, 0.1467199, 0.1548964, 0.1407434, 0.1376638, 0.1613447, 
    0.1538185, 0.2009016, 0.1684394, 0.1631654, 0.1642779, 0.09542604, 
    0.1118182, 0.117833, 0.1621785, 0.1916783,
  0.0901182, 0.0495133, 0.04172066, 0.07363967, 0.09594294, 0.07528663, 
    0.132764, 0.1233638, 0.07475225, 0.04742546, 0.04142422, 0.04668747, 
    0.05194539, 0.09400333, 0.1262354, 0.09162708, 0.1154856, 0.05859611, 
    0.06978163, 0.1242192, 0.1095237, 0.1289378, 0.0766578, 0.02246651, 
    0.04502613, 0.1016786, 0.1204828, 0.1145072, 0.09519473,
  0.01796061, -3.54265e-08, 0.09166102, 0.04868394, 0.05061346, 0.07520358, 
    0.06400955, 0.008980299, 0.0007406129, 8.176237e-05, 0.0005457688, 
    0.008982117, 0.04696491, 0.03947283, 0.06920539, 0.07390913, 0.0487653, 
    0.2099158, 0.1296762, 0.02472854, 0.1068057, 0.006928614, 9.392471e-05, 
    0.0006511885, 0.02659219, 0.1059486, 0.1169164, 0.05057508, 0.01916279,
  1.301762e-05, 0.02912147, 0.1235663, 0.01940195, 0.05555641, 0.03513233, 
    0.07171214, 0.01563541, 0.0008878402, 7.26458e-07, 0.02745895, 
    0.02003834, 0.03659749, 0.02726978, 0.09010037, 0.05131627, 0.04941842, 
    0.04554771, 0.03260151, 0.06181838, 0.02823651, 0.0002523073, 
    7.526649e-07, 0.001006307, 0.09743543, 0.2360284, 0.02313361, 
    0.006140349, -1.085485e-05,
  1.472607e-05, 0.0093995, 0.1690493, 0.0779922, 0.08286683, 0.08565921, 
    0.08623088, 0.08129434, 0.01386248, 0.008920139, 0.02462648, 0.02127288, 
    0.03091099, 0.05316876, 0.04026168, 0.04897968, 0.04216658, 0.05702654, 
    0.02091389, 0.004165265, 0.0004413994, 7.340191e-08, 3.655945e-05, 
    0.08118956, 0.1406999, 0.07336636, 0.01505245, -4.190842e-06, 0.0006986241,
  0.1710014, 0.06244583, 0.09904772, 0.07886697, 0.05194259, 0.03281483, 
    0.06114356, 0.05400343, 0.1410966, 0.160897, 0.03474566, 0.008593411, 
    0.01964511, 0.0315293, 0.02136039, 0.003897536, 0.001228814, 
    0.0004285749, 0.0007381053, 0.00102364, 0.0009935214, 0.009455139, 
    0.1059709, 0.147053, 0.133309, 0.03589031, 0.08694184, 0.05253605, 
    0.0663498,
  1.933763e-07, 1.699493e-05, 0.001247197, 0.1206552, 0.04046773, 0.02048311, 
    0.009563209, 0.01099243, 0.06107424, 0.05331794, 0.1455171, 0.07388568, 
    0.0604971, 0.06856432, 0.07799703, 0.05669229, 0.06443354, 0.1007713, 
    0.1121408, 0.1070449, 0.08516464, 0.03887609, 0.0751912, 0.03196416, 
    0.05476848, 0.01599551, 0.002139581, 5.424412e-05, 2.161688e-05,
  3.955995e-06, 3.969191e-07, 6.170106e-08, 0.01701281, 0.01592631, 
    0.006021274, 0.01317945, 0.03088192, 0.01626685, 0.09013452, 0.1447556, 
    0.04377168, 0.02219289, 0.01638212, 0.02696678, 0.03089151, 0.03883692, 
    0.09062666, 0.0566972, 0.02262526, 0.0130064, 0.08916283, 0.02241542, 
    0.03863925, 0.05023741, 0.05159805, 0.03873414, 0.003319308, 3.652862e-06,
  9.214617e-07, 0.01357866, 0.02375185, 0.05249574, 0.09217778, 0.09814166, 
    0.03541661, 0.05927435, 0.1441057, 0.1437551, 0.08187389, 0.05566051, 
    0.1004255, 0.1105386, 0.103809, 0.1653166, 0.102858, 0.0834633, 
    0.1104819, 0.05191616, 0.1197164, 0.07911576, 0.04648071, 0.04115613, 
    0.06216614, 0.06888341, 0.05734746, 0.03883176, 0.02786284,
  0.04231985, 0.07063805, 0.1672777, 0.3288777, 0.161584, 0.09980188, 
    0.1941873, 0.03455691, 0.03081164, 0.06992639, 0.04249346, 0.1228669, 
    0.1823638, 0.1707045, 0.1766337, 0.1806918, 0.1984479, 0.1229551, 
    0.1086803, 0.2082493, 0.1674883, 0.04074561, 0.142404, 0.1905755, 
    0.2313417, 0.2251116, 0.1476281, 0.1199438, 0.128113,
  0.169028, 0.2038916, 0.1822917, 0.2134987, 0.2022682, 0.2304319, 0.202087, 
    0.194172, 0.1239261, 0.07473738, 0.1006694, 0.08464783, 0.3026631, 
    0.2812147, 0.2831467, 0.2443578, 0.2231237, 0.151388, 0.1936015, 
    0.2935551, 0.1697381, 0.142358, 0.2020803, 0.2180237, 0.1783534, 
    0.2479283, 0.3263509, 0.2180822, 0.1869547,
  0.2389809, 0.2757828, 0.2953955, 0.2850278, 0.3016933, 0.3642989, 
    0.2767923, 0.3271946, 0.245466, 0.346061, 0.3586792, 0.1232771, 
    0.2933669, 0.2506842, 0.2591337, 0.2581393, 0.2618117, 0.3484352, 
    0.2848814, 0.266303, 0.2713893, 0.2148635, 0.2577625, 0.3447477, 
    0.2432895, 0.2550273, 0.2657035, 0.2857158, 0.3139495,
  0.2997543, 0.2759053, 0.3038136, 0.3185047, 0.3310145, 0.4506502, 0.42994, 
    0.5037727, 0.2995675, 0.3111279, 0.32438, 0.242464, 0.3137933, 0.3324341, 
    0.3558428, 0.1996301, 0.217796, 0.3255884, 0.2739874, 0.2958875, 
    0.2824672, 0.1608849, 0.3125622, 0.2058478, 0.1769161, 0.2966393, 
    0.373757, 0.3208496, 0.2513947,
  0.3115776, 0.3600999, 0.2740449, 0.2365963, 0.1811656, 0.2026027, 
    0.2005776, 0.2275554, 0.2333355, 0.2567258, 0.2791578, 0.2839116, 
    0.3022136, 0.2929434, 0.2495607, 0.2395222, 0.18877, 0.2344729, 
    0.3202801, 0.3234491, 0.2744213, 0.2926537, 0.2656816, 0.1014704, 
    0.1272829, 0.1071435, 0.158508, 0.2566864, 0.3581836,
  0.1126131, 0.1129964, 0.1133796, 0.1137629, 0.1141462, 0.1145295, 
    0.1149127, 0.1283027, 0.1325124, 0.1367221, 0.1409318, 0.1451415, 
    0.1493512, 0.1535608, 0.1403224, 0.1405729, 0.1408234, 0.1410739, 
    0.1413244, 0.1415749, 0.1418254, 0.1423439, 0.1375005, 0.132657, 
    0.1278136, 0.1229701, 0.1181267, 0.1132832, 0.1123065,
  0.07554144, 0.09154752, 0.1181739, 0.1282488, 0.1566981, 0.1354903, 
    0.1320864, 0.1692553, 0.1895902, 0.1441776, 0.1410839, 0.1381882, 
    0.1730897, 0.03923268, 0.06554391, 0.08096785, 0.09819856, 0.1189745, 
    0.0742617, 0.1084191, 0.1518268, 0.2846119, 0.2593702, 0.1975571, 
    0.1181715, 0.1776073, 0.1384605, 0.1174655, 0.09289001,
  0.096287, 0.1528442, 0.195635, 0.2669113, 0.4246679, 0.3803342, 0.2474702, 
    0.2639824, 0.1796465, 0.179609, 0.1285436, 0.136351, 0.2234058, 0.122752, 
    0.2445261, 0.2533129, 0.2765942, 0.2620559, 0.2155128, 0.2532935, 
    0.1663148, 0.2489541, 0.2812181, 0.3982885, 0.2118898, 0.1612231, 
    0.234822, 0.1912221, 0.09353691,
  0.1997764, 0.2747806, 0.4205329, 0.3491489, 0.3231285, 0.3085198, 
    0.2973859, 0.2863433, 0.3219309, 0.2819504, 0.3379868, 0.2852058, 
    0.2965276, 0.2956534, 0.2599444, 0.266314, 0.2434666, 0.2783409, 
    0.2984483, 0.3001729, 0.3216425, 0.3089954, 0.308234, 0.2515568, 
    0.2863613, 0.2339566, 0.2666306, 0.2454852, 0.24806,
  0.2522683, 0.2109383, 0.2029551, 0.2020996, 0.1887877, 0.1866927, 
    0.1831997, 0.2235582, 0.236034, 0.2588345, 0.2335547, 0.2119329, 
    0.2198503, 0.181518, 0.1565226, 0.1583081, 0.1489495, 0.1508963, 
    0.1864142, 0.1660876, 0.2109363, 0.1922645, 0.1856846, 0.1723938, 
    0.07562187, 0.1064966, 0.1164142, 0.1729141, 0.200081,
  0.09732233, 0.06380136, 0.06119025, 0.09243813, 0.09960485, 0.0789689, 
    0.1361766, 0.1202824, 0.08753989, 0.05716033, 0.04658181, 0.04950647, 
    0.05291653, 0.1002986, 0.1585442, 0.09720675, 0.1067214, 0.07095312, 
    0.08181604, 0.1287904, 0.1158002, 0.1245805, 0.08680987, 0.02589306, 
    0.03732052, 0.099922, 0.1211215, 0.1118533, 0.105072,
  0.02672347, -1.136879e-06, 0.07574608, 0.04071176, 0.06690807, 0.06563441, 
    0.0815932, 0.02329525, 0.004338006, 0.0005521849, 0.0002062601, 
    0.003167263, 0.0348797, 0.0389412, 0.07761218, 0.08628245, 0.05699302, 
    0.2051224, 0.1168239, 0.02828248, 0.1073714, 0.01705591, 0.002089205, 
    0.0004535852, 0.01835028, 0.1051606, 0.1327119, 0.06429026, 0.03678597,
  3.166036e-06, 0.01712986, 0.1181853, 0.01821409, 0.05983013, 0.03970517, 
    0.07442461, 0.02220147, 0.003599874, -2.087996e-07, 0.02267184, 
    0.01409921, 0.0432165, 0.02901806, 0.09054545, 0.05554155, 0.05146421, 
    0.03604782, 0.02860845, 0.04968365, 0.06692571, 0.01270349, 5.577505e-07, 
    0.0005817012, 0.09339722, 0.2127803, 0.02562683, 0.02281852, 0.001225926,
  6.929851e-06, 0.008739237, 0.1601932, 0.06828108, 0.06754516, 0.08378628, 
    0.07566966, 0.08071961, 0.01888373, 0.009582818, 0.0306677, 0.01844084, 
    0.0317998, 0.04685783, 0.03132769, 0.04715515, 0.03813347, 0.04849172, 
    0.02286078, 0.01027338, 0.003508026, 2.239751e-07, 1.331103e-05, 
    0.07864634, 0.1163637, 0.05170017, 0.03300028, 0.0002574659, 0.003449704,
  0.1448976, 0.06293375, 0.1028497, 0.1009478, 0.0500979, 0.02902856, 
    0.05612881, 0.04597095, 0.1532075, 0.163794, 0.03379252, 0.008918889, 
    0.02006057, 0.02491579, 0.02183485, 0.008839791, 0.002584099, 
    0.003300223, 0.002827391, 0.0003354373, 0.001383681, 0.01919836, 
    0.09048815, 0.1397698, 0.1126508, 0.03154002, 0.08423132, 0.06027211, 
    0.06845702,
  1.116233e-07, 7.934034e-07, -1.110061e-05, 0.1038557, 0.0584056, 
    0.02637398, 0.02011538, 0.01754855, 0.06306379, 0.05501856, 0.1388825, 
    0.06704903, 0.05911291, 0.06508562, 0.08166461, 0.0596152, 0.06081042, 
    0.1001789, 0.1215768, 0.1066419, 0.07823037, 0.03566343, 0.08263139, 
    0.03284384, 0.04693575, 0.01976946, 0.002990718, 1.032351e-05, 
    -1.526555e-06,
  2.106086e-06, 2.360441e-07, 2.628044e-08, 0.032224, 0.002880538, 
    0.01566702, 0.02132769, 0.03348876, 0.01849521, 0.1049305, 0.1417638, 
    0.07470002, 0.03580683, 0.03054747, 0.04204245, 0.04283793, 0.04023058, 
    0.09530647, 0.05552588, 0.03838602, 0.01482072, 0.1155686, 0.03062513, 
    0.0395832, 0.04147246, 0.0374805, 0.04384762, 0.00377555, 2.973883e-06,
  -2.372216e-05, 0.02928837, 0.03548177, 0.06283194, 0.09970613, 0.09540825, 
    0.01717197, 0.04908762, 0.1174112, 0.1244443, 0.08231422, 0.08037291, 
    0.1034691, 0.11721, 0.1074179, 0.1716046, 0.1129879, 0.08926739, 
    0.1196641, 0.05092578, 0.1113897, 0.08780985, 0.05908745, 0.0504322, 
    0.06937934, 0.07422452, 0.06203964, 0.04689464, 0.03174864,
  0.03554358, 0.07756211, 0.1646479, 0.3368262, 0.1571487, 0.09494399, 
    0.1925711, 0.0326109, 0.02590879, 0.06211689, 0.0435406, 0.1831948, 
    0.2204961, 0.2057365, 0.2120521, 0.2031052, 0.2200281, 0.1538077, 
    0.1623811, 0.1998732, 0.1859729, 0.03569997, 0.1357936, 0.1873498, 
    0.2611971, 0.2279298, 0.1624312, 0.1187843, 0.1462273,
  0.1646594, 0.216081, 0.1789949, 0.2329933, 0.1671087, 0.2157212, 0.184734, 
    0.1964676, 0.1206359, 0.07413487, 0.1011143, 0.08382249, 0.3746097, 
    0.3157439, 0.2981971, 0.2596879, 0.2127705, 0.1592643, 0.213116, 
    0.2908261, 0.1730361, 0.1512225, 0.200808, 0.2615108, 0.2108799, 
    0.2946455, 0.3393834, 0.2225068, 0.1854309,
  0.2511216, 0.2737166, 0.2940059, 0.3682483, 0.2974014, 0.3273462, 0.260429, 
    0.2920901, 0.2419668, 0.3670232, 0.3778372, 0.1113356, 0.318347, 
    0.2579281, 0.2819872, 0.2809184, 0.2625296, 0.3486211, 0.2759026, 
    0.228617, 0.2549717, 0.1932663, 0.2286129, 0.3024264, 0.288664, 
    0.2614822, 0.2832493, 0.2881439, 0.3199629,
  0.2805528, 0.2805932, 0.2959405, 0.3273813, 0.2637883, 0.4112598, 
    0.4173697, 0.497143, 0.3185772, 0.3643106, 0.3343181, 0.2451239, 
    0.3235707, 0.34276, 0.4035161, 0.2191198, 0.2280629, 0.3315245, 
    0.2602917, 0.2791273, 0.2936524, 0.1557414, 0.3220114, 0.2040598, 
    0.167181, 0.3095252, 0.3857812, 0.3487843, 0.2680289,
  0.3288362, 0.3033644, 0.2770615, 0.2344454, 0.1944855, 0.1740441, 
    0.1809111, 0.2243474, 0.2365101, 0.2605263, 0.2857203, 0.2909243, 
    0.2940048, 0.2857775, 0.2475837, 0.2505185, 0.2266006, 0.2555901, 
    0.3267885, 0.3682477, 0.3135426, 0.3211068, 0.2641093, 0.090027, 
    0.1160425, 0.09030773, 0.1639813, 0.2511837, 0.3682004,
  0.113094, 0.1137209, 0.1143478, 0.1149748, 0.1156017, 0.1162286, 0.1168555, 
    0.1192766, 0.1226823, 0.126088, 0.1294938, 0.1328995, 0.1363052, 
    0.139711, 0.128202, 0.128973, 0.1297439, 0.1305149, 0.1312859, 0.1320568, 
    0.1328278, 0.141878, 0.1370744, 0.1322708, 0.1274671, 0.1226635, 
    0.1178599, 0.1130563, 0.1125925,
  0.08581737, 0.09398684, 0.1116374, 0.1240097, 0.1512266, 0.1416471, 
    0.1637827, 0.1847922, 0.189481, 0.1659279, 0.1539198, 0.133872, 
    0.1906596, 0.03428087, 0.08616813, 0.1175682, 0.1004451, 0.1165331, 
    0.07479464, 0.1027798, 0.1886309, 0.3080893, 0.2969446, 0.2467573, 
    0.2150048, 0.2082281, 0.1797132, 0.105015, 0.1135013,
  0.09206925, 0.1495731, 0.2223769, 0.214843, 0.3995388, 0.3956397, 
    0.2160938, 0.2449472, 0.1768048, 0.1969155, 0.1458248, 0.1348378, 
    0.1978072, 0.161362, 0.2239443, 0.2530184, 0.3300113, 0.350386, 
    0.2434135, 0.2712787, 0.2038741, 0.2644199, 0.2856452, 0.3877648, 
    0.2212636, 0.2029565, 0.1775981, 0.1669325, 0.08966388,
  0.2476416, 0.2944619, 0.4687362, 0.3472112, 0.3405331, 0.2948208, 
    0.3376975, 0.2933979, 0.343524, 0.3233147, 0.3457831, 0.2969372, 
    0.3198741, 0.3170647, 0.2942399, 0.2763929, 0.2415978, 0.269193, 
    0.3177681, 0.3413348, 0.3469772, 0.3460582, 0.3354903, 0.2858802, 
    0.3117145, 0.2678693, 0.2891714, 0.3171458, 0.3290843,
  0.2785926, 0.2448344, 0.239803, 0.2409029, 0.217289, 0.2061158, 0.1984593, 
    0.2430596, 0.2785601, 0.2962881, 0.2868265, 0.2607017, 0.2570905, 
    0.2113853, 0.1514837, 0.1665757, 0.1686035, 0.2070614, 0.2236279, 
    0.1996584, 0.2410897, 0.223373, 0.2186156, 0.1762713, 0.05956984, 
    0.1057827, 0.1387853, 0.1978599, 0.2343011,
  0.13011, 0.1130033, 0.1150802, 0.1380193, 0.1188324, 0.1115465, 0.1520041, 
    0.1347982, 0.116317, 0.0904253, 0.06069099, 0.06603862, 0.06735072, 
    0.1269275, 0.1953781, 0.09948842, 0.1149805, 0.09873079, 0.1130795, 
    0.1437812, 0.1668368, 0.1530592, 0.1185535, 0.03006049, 0.02679922, 
    0.1224481, 0.1544297, 0.1298004, 0.1144689,
  0.0433757, 3.002965e-05, 0.06879886, 0.04606442, 0.07301884, 0.07004113, 
    0.1072572, 0.04797989, 0.02351842, 0.003382348, 8.173261e-05, 
    0.001025569, 0.0308526, 0.0490649, 0.08935632, 0.1067576, 0.07042995, 
    0.2269565, 0.1135049, 0.0289388, 0.1221752, 0.04407679, 0.01502126, 
    0.0002330828, 0.01375435, 0.11098, 0.1259626, 0.07725057, 0.05443327,
  0.0001515142, 0.008831807, 0.1049564, 0.01912493, 0.06204163, 0.04184352, 
    0.07708412, 0.02920018, 0.01644396, 3.623064e-08, 0.0197196, 0.01154714, 
    0.04116888, 0.02714868, 0.09076442, 0.05282991, 0.05265491, 0.02998906, 
    0.02675628, 0.04751769, 0.09025282, 0.04405684, 1.678387e-05, 
    0.0004731846, 0.09422661, 0.2011237, 0.03308977, 0.06429434, 0.01357232,
  1.574942e-05, 0.009489536, 0.1561059, 0.06007573, 0.0546611, 0.07153513, 
    0.06305182, 0.07730392, 0.02623168, 0.01329328, 0.03653339, 0.0164208, 
    0.03097216, 0.03837272, 0.02552751, 0.04418484, 0.03377096, 0.04215904, 
    0.02444233, 0.01825538, 0.01002601, 0.0006133163, 3.974668e-06, 
    0.07256564, 0.09685783, 0.04235662, 0.05282965, 0.008587044, 0.002691348,
  0.1233028, 0.0707617, 0.1167454, 0.107302, 0.04643179, 0.0269494, 
    0.05117627, 0.0389549, 0.163206, 0.1698912, 0.03238843, 0.01028941, 
    0.01998155, 0.019533, 0.02435125, 0.01179716, 0.007414828, 0.008516619, 
    0.008908058, 0.005028707, 0.006346682, 0.01855062, 0.06783153, 0.1254096, 
    0.09053396, 0.0303239, 0.0747225, 0.04945516, 0.05620122,
  2.508901e-08, 6.233785e-08, -3.983791e-06, 0.06982305, 0.0951957, 
    0.03415574, 0.01901057, 0.02575753, 0.07072592, 0.0490229, 0.1246706, 
    0.051601, 0.05719981, 0.05612837, 0.07635011, 0.05886859, 0.05557268, 
    0.09184089, 0.120963, 0.1018611, 0.07333186, 0.02928966, 0.09496987, 
    0.03521895, 0.0421828, 0.02802076, 0.007983935, -3.788207e-05, 
    -1.303918e-06,
  6.635206e-07, 1.499056e-07, 1.643198e-08, 0.07012333, 0.001068705, 
    0.03982551, 0.02822965, 0.03503155, 0.04102427, 0.1402707, 0.1638826, 
    0.0848615, 0.0425104, 0.04981838, 0.04795887, 0.04716074, 0.05168023, 
    0.1050189, 0.06607492, 0.05846131, 0.01706215, 0.1573729, 0.03608298, 
    0.03643317, 0.03819539, 0.03249672, 0.04677888, 0.005729879, -3.010928e-07,
  0.001261446, 0.03037603, 0.076571, 0.06388404, 0.104204, 0.07980721, 
    0.009919186, 0.03304609, 0.09535152, 0.1302015, 0.1073878, 0.1502181, 
    0.151879, 0.1635481, 0.1318896, 0.1755932, 0.1265405, 0.0973951, 
    0.162185, 0.08392316, 0.1214117, 0.1213864, 0.07220469, 0.09350792, 
    0.09499654, 0.1014142, 0.07232894, 0.07581948, 0.02307351,
  0.03504742, 0.08470716, 0.1579697, 0.3503429, 0.1532789, 0.1081632, 
    0.1780629, 0.02948672, 0.02127465, 0.06022415, 0.0517076, 0.2496386, 
    0.2460494, 0.2475928, 0.2486047, 0.2330047, 0.2568528, 0.2172078, 
    0.2440292, 0.2223968, 0.1912567, 0.03787653, 0.1459573, 0.2010659, 
    0.30011, 0.2383655, 0.1782947, 0.1328508, 0.1638298,
  0.1931472, 0.2431703, 0.2609789, 0.2694505, 0.1793317, 0.2408008, 
    0.1861522, 0.207991, 0.09507453, 0.08038871, 0.1130754, 0.09031875, 
    0.3913478, 0.352598, 0.3145947, 0.258113, 0.2082852, 0.1915933, 
    0.2551993, 0.3166927, 0.1722674, 0.1839606, 0.2147045, 0.2837723, 
    0.2261925, 0.3279154, 0.3345275, 0.2280618, 0.2241393,
  0.2565327, 0.2841974, 0.3298981, 0.343254, 0.3487402, 0.3199569, 0.3073173, 
    0.2866125, 0.3106673, 0.3803807, 0.4158956, 0.1138087, 0.3460466, 
    0.2660992, 0.3590564, 0.3241928, 0.2755606, 0.3565023, 0.2777309, 
    0.2421381, 0.2674998, 0.2063638, 0.2565737, 0.3218057, 0.4122498, 
    0.2426735, 0.3066605, 0.2917108, 0.3307928,
  0.2998419, 0.3046346, 0.2672946, 0.3952773, 0.3277723, 0.4332521, 
    0.4312292, 0.4584246, 0.3176785, 0.4204403, 0.3488512, 0.2619641, 
    0.3528018, 0.3847989, 0.4403774, 0.2167323, 0.2458684, 0.3590681, 
    0.2520832, 0.3016031, 0.305509, 0.2159357, 0.3357064, 0.2146366, 
    0.1627463, 0.3213697, 0.3954623, 0.3698355, 0.3134937,
  0.3522784, 0.2214972, 0.2323063, 0.2150175, 0.2020038, 0.1781582, 0.192181, 
    0.2448318, 0.2386845, 0.2564821, 0.2759685, 0.3115349, 0.3114588, 
    0.312039, 0.2556178, 0.250888, 0.2528839, 0.2768164, 0.335424, 0.3937374, 
    0.3109262, 0.3718469, 0.2614812, 0.08910921, 0.1181068, 0.08146249, 
    0.1617019, 0.2615437, 0.3927392,
  0.1226261, 0.1232454, 0.1238647, 0.124484, 0.1251033, 0.1257226, 0.126342, 
    0.1270058, 0.1289541, 0.1309023, 0.1328506, 0.1347989, 0.1367471, 
    0.1386954, 0.1474949, 0.150392, 0.1532891, 0.1561862, 0.1590833, 
    0.1619804, 0.1648775, 0.1746237, 0.169159, 0.1636943, 0.1582297, 
    0.152765, 0.1473003, 0.1418357, 0.1221307,
  0.1051437, 0.1115251, 0.1182359, 0.1476565, 0.1592335, 0.1459581, 
    0.1616252, 0.2020019, 0.2369596, 0.2299709, 0.2151545, 0.1609956, 
    0.202596, 0.01169765, 0.1718276, 0.1315004, 0.1652597, 0.1247865, 
    0.1015629, 0.1197347, 0.1944944, 0.3354771, 0.3241403, 0.1588499, 
    0.1871342, 0.2202113, 0.1468284, 0.1288993, 0.1324211,
  0.1241931, 0.1384515, 0.1895987, 0.1669322, 0.3563578, 0.3997914, 
    0.2040201, 0.2387346, 0.1814069, 0.1947643, 0.179302, 0.1435601, 
    0.1712222, 0.1544786, 0.2746759, 0.3277738, 0.4278421, 0.4109155, 
    0.3045588, 0.3300714, 0.2476293, 0.2765225, 0.2862962, 0.3987597, 
    0.2452795, 0.3095316, 0.2277587, 0.2065029, 0.1223884,
  0.3394618, 0.3569775, 0.5076181, 0.3981164, 0.3988395, 0.4281894, 
    0.4130723, 0.3843864, 0.3644777, 0.3756144, 0.3919399, 0.3623891, 
    0.3608139, 0.3662627, 0.328702, 0.3200574, 0.3207819, 0.3352005, 0.36725, 
    0.4049906, 0.4125206, 0.4188184, 0.4172985, 0.3374067, 0.3697147, 
    0.3297793, 0.337388, 0.3719183, 0.4728894,
  0.320365, 0.2946296, 0.2794088, 0.2990818, 0.2600116, 0.24597, 0.2506378, 
    0.3040012, 0.3377131, 0.3580728, 0.364604, 0.3072175, 0.2865312, 
    0.2512764, 0.1666216, 0.1988308, 0.205491, 0.2520942, 0.2835531, 
    0.2816142, 0.2994291, 0.2600868, 0.2500468, 0.1699775, 0.05221035, 
    0.1231243, 0.1967108, 0.2603061, 0.2761981,
  0.1780704, 0.1962809, 0.1839221, 0.1741315, 0.1716968, 0.1734798, 
    0.2268838, 0.2158638, 0.1888274, 0.1673486, 0.1207148, 0.08886229, 
    0.08666572, 0.1411945, 0.1971621, 0.1438031, 0.1563223, 0.1562234, 
    0.1653658, 0.1792016, 0.2361036, 0.2159606, 0.2010069, 0.03286039, 
    0.02868314, 0.1561555, 0.1953126, 0.186344, 0.1589445,
  0.07879235, 0.0109452, 0.05569835, 0.05452327, 0.1013424, 0.1036046, 
    0.1323051, 0.09314251, 0.09052393, 0.02324874, 0.0001309664, 
    0.0004542181, 0.0197361, 0.08576038, 0.1055507, 0.1329121, 0.09123448, 
    0.2333288, 0.1141065, 0.04911078, 0.1365683, 0.1046347, 0.09217985, 
    9.188957e-05, 0.01265582, 0.120911, 0.1337819, 0.08811412, 0.09021973,
  0.006258553, 0.003873421, 0.08298141, 0.02079308, 0.07462095, 0.04294163, 
    0.08210953, 0.05702374, 0.04346395, 1.472568e-08, 0.01376587, 0.00981853, 
    0.04630575, 0.0268659, 0.08976747, 0.0587021, 0.05252635, 0.0276651, 
    0.03001648, 0.04554687, 0.08359935, 0.1639622, 0.005216357, 0.0006036759, 
    0.08951771, 0.1856378, 0.04618029, 0.1052636, 0.09398514,
  0.001819881, 0.01720994, 0.1432088, 0.05459798, 0.04707535, 0.06610455, 
    0.05447955, 0.06461835, 0.03497504, 0.0230839, 0.0354034, 0.02006021, 
    0.03376672, 0.03388753, 0.0264072, 0.04261941, 0.03874461, 0.04109055, 
    0.02856729, 0.03694148, 0.05746745, 0.01759528, 0.001051525, 0.06663517, 
    0.08118069, 0.03475441, 0.06327263, 0.04550156, 0.01679066,
  0.09941579, 0.05736061, 0.09336594, 0.1025864, 0.04584096, 0.0254375, 
    0.04790431, 0.0352748, 0.1576834, 0.1772638, 0.03609701, 0.01436548, 
    0.02204776, 0.02137765, 0.02876984, 0.01427551, 0.009492531, 0.009847693, 
    0.0140952, 0.01740746, 0.02527544, 0.02333803, 0.05340526, 0.1049073, 
    0.080259, 0.03118018, 0.06304155, 0.03860103, 0.05216676,
  2.83699e-09, 1.193968e-08, -2.674671e-07, 0.03686435, 0.1338428, 
    0.03441051, 0.01437542, 0.06665659, 0.1130324, 0.05032605, 0.116342, 
    0.04609139, 0.0509723, 0.05122222, 0.06889641, 0.0603689, 0.05182169, 
    0.08860181, 0.1193465, 0.09309676, 0.06672099, 0.02970137, 0.1035793, 
    0.03939175, 0.04365024, 0.03701206, 0.03502341, -5.767228e-05, 
    -6.815347e-07,
  2.189386e-07, 8.526481e-08, -1.999454e-07, 0.07118299, 0.002741263, 
    0.09525175, 0.01974559, 0.05829558, 0.05572617, 0.2602965, 0.2402782, 
    0.1177895, 0.07204107, 0.07920235, 0.05490628, 0.06439891, 0.09232843, 
    0.1032767, 0.1046555, 0.1107639, 0.01647679, 0.2144988, 0.07137179, 
    0.04224781, 0.04135922, 0.04059215, 0.06486315, 0.009886424, -3.57871e-06,
  0.01211696, 0.06891073, 0.113214, 0.08256453, 0.1149769, 0.06542969, 
    0.006278899, 0.02278812, 0.07614428, 0.1566719, 0.2254921, 0.2105252, 
    0.1354688, 0.1643006, 0.1709829, 0.1907382, 0.1886506, 0.125242, 
    0.2201507, 0.1166006, 0.1308212, 0.1674089, 0.1073158, 0.1975609, 
    0.1497374, 0.15372, 0.1292776, 0.115438, 0.02255645,
  0.04233995, 0.07984757, 0.1746231, 0.358973, 0.1376388, 0.1090367, 
    0.1593264, 0.01942672, 0.0154082, 0.04927351, 0.08623925, 0.3263974, 
    0.271111, 0.2637552, 0.2557187, 0.2501011, 0.2939026, 0.3000591, 
    0.2295706, 0.256878, 0.1881238, 0.04213278, 0.1813633, 0.2201223, 
    0.3110339, 0.2296413, 0.1938856, 0.1792438, 0.1924029,
  0.2053848, 0.2671627, 0.3084328, 0.2821442, 0.2450278, 0.2485584, 
    0.2067412, 0.2234566, 0.07296452, 0.07846621, 0.1296442, 0.1061062, 
    0.3965392, 0.3016483, 0.2683572, 0.2435628, 0.2263136, 0.1993731, 
    0.2770166, 0.3511339, 0.1626091, 0.1749208, 0.272813, 0.3385542, 
    0.2528604, 0.3090227, 0.3049469, 0.2243833, 0.2321629,
  0.2720269, 0.2951477, 0.3792521, 0.3873374, 0.3807761, 0.3772147, 
    0.3268171, 0.3323255, 0.3238468, 0.4205864, 0.4769795, 0.1245606, 
    0.3616401, 0.2457205, 0.4898619, 0.3705582, 0.2965955, 0.3607772, 
    0.2907591, 0.2591792, 0.3085119, 0.2062327, 0.2967191, 0.3480355, 
    0.6041601, 0.2060216, 0.2973315, 0.2744359, 0.3218362,
  0.3369908, 0.3439181, 0.2554846, 0.4113486, 0.4356875, 0.4694301, 
    0.4810949, 0.4520474, 0.3274906, 0.4662637, 0.3898277, 0.2985258, 
    0.401219, 0.421599, 0.4710777, 0.210538, 0.2813314, 0.3743457, 0.2709427, 
    0.3471565, 0.3019601, 0.2943759, 0.3589969, 0.2045522, 0.1497468, 
    0.3196737, 0.4155067, 0.3610743, 0.3629419,
  0.2993615, 0.2233081, 0.2098701, 0.1800268, 0.1723134, 0.1647017, 
    0.2146794, 0.2516764, 0.2229398, 0.2708862, 0.3008965, 0.3332725, 
    0.3523552, 0.3757376, 0.2777583, 0.2850986, 0.2824523, 0.3219937, 
    0.3768717, 0.3979776, 0.3284889, 0.3973721, 0.2939101, 0.09990277, 
    0.1198522, 0.06891748, 0.1697714, 0.2882376, 0.4284298,
  0.1653553, 0.1671763, 0.1689973, 0.1708183, 0.1726393, 0.1744602, 
    0.1762812, 0.1621766, 0.1617954, 0.1614142, 0.161033, 0.1606518, 
    0.1602706, 0.1598894, 0.1927365, 0.1977093, 0.202682, 0.2076547, 
    0.2126275, 0.2176002, 0.222573, 0.2013042, 0.1948917, 0.1884792, 
    0.1820666, 0.1756541, 0.1692415, 0.162829, 0.1638985,
  0.1387183, 0.1345223, 0.1427954, 0.1648795, 0.1784588, 0.1467242, 
    0.1626769, 0.207771, 0.25485, 0.2465972, 0.2257434, 0.1944188, 0.2094576, 
    0.002149967, 0.2072491, 0.1402115, 0.1739654, 0.1528266, 0.1443453, 
    0.1487909, 0.2549737, 0.3324545, 0.3330535, 0.1559997, 0.1927004, 
    0.2392442, 0.1674635, 0.1244796, 0.125464,
  0.1463785, 0.1731229, 0.1706184, 0.1482019, 0.3101055, 0.4262487, 
    0.1933132, 0.2224003, 0.1926602, 0.1950345, 0.2214523, 0.2009906, 
    0.141133, 0.1673881, 0.2907704, 0.4410949, 0.4095158, 0.4370131, 
    0.4031802, 0.389918, 0.29767, 0.3087154, 0.3674972, 0.4216775, 0.22425, 
    0.3294351, 0.3814708, 0.3026316, 0.1268516,
  0.4285945, 0.4326926, 0.5530019, 0.4751195, 0.4854752, 0.477138, 0.4442275, 
    0.4166247, 0.3935868, 0.3956057, 0.426673, 0.4116273, 0.4260438, 
    0.4172183, 0.3450477, 0.3644277, 0.3823044, 0.385708, 0.4216381, 
    0.4161938, 0.4456761, 0.4225684, 0.4289947, 0.402414, 0.4610229, 
    0.381475, 0.4199159, 0.4297175, 0.5192846,
  0.3932921, 0.3770272, 0.3333309, 0.3622199, 0.3476776, 0.3528219, 0.309022, 
    0.377739, 0.3812312, 0.3898709, 0.382365, 0.3283253, 0.3265517, 
    0.2910063, 0.1922737, 0.2191732, 0.251891, 0.3213498, 0.315491, 
    0.3402412, 0.3306908, 0.2995131, 0.3140086, 0.1707568, 0.04891495, 
    0.1526531, 0.2475365, 0.3413163, 0.3551182,
  0.2726926, 0.2330998, 0.2190404, 0.2238344, 0.2490768, 0.2484003, 
    0.3014719, 0.2760085, 0.3024806, 0.2630273, 0.1682088, 0.124314, 
    0.1181167, 0.2224083, 0.2129402, 0.2343373, 0.2201664, 0.2330683, 
    0.270476, 0.2702699, 0.2865839, 0.2451769, 0.2303122, 0.04292249, 
    0.04228411, 0.178542, 0.2648297, 0.2443222, 0.2122635,
  0.2414674, 0.06435917, 0.0445862, 0.1146452, 0.1427701, 0.1567983, 
    0.1478154, 0.1853189, 0.2208624, 0.06912844, 0.0008430105, 0.0007319528, 
    0.009263653, 0.1068752, 0.160903, 0.1336112, 0.1269249, 0.2512142, 
    0.1463727, 0.08362401, 0.139355, 0.1364503, 0.2508084, 9.403231e-05, 
    0.01140863, 0.1486611, 0.1422359, 0.1336958, 0.1986531,
  0.1476114, 0.004358052, 0.06020284, 0.02725966, 0.0953019, 0.06053934, 
    0.08020077, 0.1034155, 0.1829972, -0.0001127032, 0.008682271, 
    0.005778498, 0.05901545, 0.03743571, 0.09746324, 0.06758144, 0.07869984, 
    0.03007734, 0.04017177, 0.05261343, 0.07804179, 0.2557671, 0.1413541, 
    0.001244416, 0.06689803, 0.1605458, 0.05357426, 0.1409583, 0.2589565,
  0.02909852, 0.02972895, 0.1129941, 0.04702085, 0.04979395, 0.06781822, 
    0.05202203, 0.06438579, 0.04483233, 0.03533613, 0.04001472, 0.03282616, 
    0.04405419, 0.03842658, 0.04140685, 0.06096872, 0.03967138, 0.05206322, 
    0.04465749, 0.0794201, 0.1207438, 0.1290131, 0.01051889, 0.05002622, 
    0.06475203, 0.02413997, 0.0874407, 0.09004957, 0.07065262,
  0.08528028, 0.02725872, 0.05768447, 0.09413695, 0.05073429, 0.02958864, 
    0.05146733, 0.04068763, 0.15927, 0.1851494, 0.04269221, 0.02143659, 
    0.02777871, 0.0360681, 0.05210807, 0.04911472, 0.01112832, 0.008891195, 
    0.02475269, 0.02304517, 0.05706368, 0.04205009, 0.04957572, 0.07451545, 
    0.06662478, 0.03811863, 0.05910827, 0.03417698, 0.03909274,
  8.267824e-10, 4.12571e-09, 9.396017e-08, 0.01907453, 0.1480235, 0.0990902, 
    0.004035046, 0.1199026, 0.1586999, 0.06983887, 0.1101512, 0.05006585, 
    0.05422188, 0.0765473, 0.08150305, 0.0738865, 0.05627602, 0.0917221, 
    0.1141896, 0.08448733, 0.06522877, 0.03701597, 0.1413256, 0.05410492, 
    0.0559772, 0.0559614, 0.1958621, 0.004984154, -6.357009e-07,
  7.059227e-08, -5.119429e-06, 3.828707e-05, 0.03962206, 0.002457118, 
    0.1882458, 0.01681845, 0.08652712, 0.03896189, 0.3403634, 0.248624, 
    0.1661801, 0.08976337, 0.08397415, 0.09072185, 0.08150337, 0.1159676, 
    0.1062197, 0.1891819, 0.1990702, 0.0167481, 0.2329034, 0.08784683, 
    0.0505115, 0.05028085, 0.05532356, 0.07880958, 0.005622896, -2.430742e-06,
  0.005612458, 0.1415764, 0.06535186, 0.1135, 0.1188009, 0.06637497, 
    0.00202144, 0.01566028, 0.05590075, 0.1631046, 0.3626416, 0.1081203, 
    0.1075304, 0.1201279, 0.1504541, 0.2173226, 0.2089792, 0.1566286, 
    0.1872324, 0.1109796, 0.1390314, 0.1927211, 0.1358082, 0.1935217, 
    0.1314645, 0.1298346, 0.1354588, 0.1561169, 0.01852664,
  0.05256736, 0.1075041, 0.2079007, 0.3620382, 0.1212547, 0.1124615, 
    0.1486848, 0.008455135, 0.01263629, 0.05839601, 0.1474139, 0.2570318, 
    0.2187466, 0.1788302, 0.2227325, 0.2269864, 0.3369936, 0.3303475, 
    0.1897755, 0.2963074, 0.1861446, 0.04790388, 0.2312569, 0.2735494, 
    0.2743006, 0.2068449, 0.1692387, 0.1921652, 0.2438561,
  0.2256212, 0.3304263, 0.311599, 0.3572366, 0.306192, 0.2619096, 0.2114083, 
    0.2486253, 0.06412072, 0.1029782, 0.1502227, 0.1222478, 0.2959221, 
    0.2304933, 0.2224919, 0.2525158, 0.2974799, 0.1816798, 0.2425891, 
    0.3694446, 0.1570004, 0.1961472, 0.3006339, 0.4194237, 0.2784868, 
    0.2725765, 0.2635091, 0.2040991, 0.2260955,
  0.2518343, 0.293414, 0.401081, 0.3973569, 0.44669, 0.4044086, 0.345155, 
    0.387677, 0.3903682, 0.4744697, 0.5333937, 0.167227, 0.3869064, 
    0.2469931, 0.5673884, 0.3545514, 0.3376904, 0.3576148, 0.350325, 
    0.264945, 0.3714727, 0.2650383, 0.3106015, 0.3765036, 0.5412265, 
    0.1536571, 0.2235648, 0.2460954, 0.3016621,
  0.3340352, 0.3025256, 0.2875224, 0.3622339, 0.4801183, 0.5240726, 
    0.4789495, 0.4763003, 0.3566769, 0.4866805, 0.3895482, 0.3374949, 
    0.446397, 0.4482927, 0.5257137, 0.2310227, 0.3154622, 0.3831929, 
    0.2921502, 0.4095571, 0.3461302, 0.326927, 0.3903233, 0.2148618, 
    0.1148987, 0.3119341, 0.4406972, 0.3197502, 0.4553026,
  0.2840788, 0.2278108, 0.233747, 0.2107543, 0.1852548, 0.160905, 0.2609142, 
    0.3099751, 0.2327131, 0.3173156, 0.3832473, 0.3572424, 0.3841019, 
    0.4272171, 0.3271127, 0.34759, 0.3204873, 0.3680107, 0.3988027, 
    0.4078806, 0.3341835, 0.4084966, 0.2983834, 0.1106246, 0.1135287, 
    0.06479272, 0.1652857, 0.2960909, 0.4269479,
  0.2382834, 0.2375309, 0.2367784, 0.2360258, 0.2352733, 0.2345208, 
    0.2337683, 0.25374, 0.2546552, 0.2555704, 0.2564856, 0.2574008, 0.258316, 
    0.2592312, 0.282976, 0.288834, 0.294692, 0.30055, 0.3064079, 0.3122659, 
    0.3181239, 0.297878, 0.2918573, 0.2858366, 0.2798159, 0.2737953, 
    0.2677746, 0.2617539, 0.2388854,
  0.146882, 0.1620955, 0.1760684, 0.1526761, 0.1935666, 0.1438102, 0.1527439, 
    0.2113294, 0.3079911, 0.262823, 0.2512779, 0.2611479, 0.2726252, 
    0.003268171, 0.1840685, 0.2138869, 0.1753237, 0.1963033, 0.1474188, 
    0.1580467, 0.3387406, 0.3489028, 0.3595943, 0.1503464, 0.2252631, 
    0.2455303, 0.1445988, 0.131261, 0.1487895,
  0.1229725, 0.2245556, 0.2415134, 0.1318981, 0.2053193, 0.442587, 0.1656075, 
    0.1669647, 0.1563004, 0.1549023, 0.2173715, 0.2324759, 0.1083674, 
    0.1811827, 0.3131576, 0.4518912, 0.4390567, 0.3864364, 0.3835449, 
    0.3895632, 0.3252754, 0.3306349, 0.4126445, 0.4141846, 0.2164842, 
    0.2734095, 0.3755873, 0.3491801, 0.1516569,
  0.4842794, 0.4486013, 0.5730792, 0.4923525, 0.5728986, 0.5175681, 0.490569, 
    0.4106775, 0.4119141, 0.4093986, 0.4149584, 0.4075355, 0.4838687, 
    0.4417683, 0.3604919, 0.3873191, 0.4389988, 0.4289201, 0.4772248, 
    0.4061236, 0.439904, 0.4205523, 0.4062446, 0.4161057, 0.4685494, 
    0.4496431, 0.4976797, 0.4638588, 0.5398334,
  0.4266534, 0.4111103, 0.4019305, 0.4251258, 0.3967867, 0.4122356, 
    0.3954104, 0.42835, 0.4285546, 0.4189277, 0.3698909, 0.3153616, 0.299964, 
    0.264895, 0.1779609, 0.247272, 0.3412099, 0.3772144, 0.3173444, 
    0.3292457, 0.3146979, 0.3125345, 0.3249079, 0.1714495, 0.04135902, 
    0.1554118, 0.2824091, 0.4012809, 0.3954898,
  0.2728779, 0.2272301, 0.1498329, 0.2018718, 0.2347503, 0.2616348, 
    0.3470039, 0.3220066, 0.3498021, 0.2609524, 0.2472048, 0.1116897, 
    0.1223984, 0.3179083, 0.2047844, 0.2844049, 0.3321007, 0.3544291, 
    0.3351257, 0.2630228, 0.2618421, 0.2361425, 0.1919905, 0.05049343, 
    0.03552131, 0.1793904, 0.2884995, 0.2532478, 0.2162875,
  0.3284234, 0.08146772, 0.03697054, 0.1423119, 0.1413813, 0.1539175, 
    0.1951138, 0.2552006, 0.3480718, 0.04088899, 0.01020441, 5.049053e-05, 
    0.003264658, 0.1138903, 0.1383817, 0.1615141, 0.1204322, 0.2577193, 
    0.1353694, 0.1116586, 0.1706493, 0.1804689, 0.3009252, 0.0002129876, 
    0.01256881, 0.2049572, 0.1545265, 0.1466115, 0.2379277,
  0.5245249, 0.006734914, 0.04606709, 0.0589585, 0.09695746, 0.07734715, 
    0.09550564, 0.09774719, 0.2584319, 0.001745233, 0.006237237, 0.001922124, 
    0.09270118, 0.09131561, 0.1045496, 0.07184459, 0.07667383, 0.04498089, 
    0.04891261, 0.05863995, 0.04447808, 0.1900744, 0.6189395, 0.003796131, 
    0.04517576, 0.1488353, 0.07064891, 0.1062761, 0.3102489,
  0.1703579, 0.06477525, 0.08249591, 0.04439333, 0.06507792, 0.07303056, 
    0.0622524, 0.08780168, 0.1056761, 0.1307877, 0.05880536, 0.08824956, 
    0.06952731, 0.07511806, 0.07376219, 0.06214872, 0.03797778, 0.0467108, 
    0.05336957, 0.05866091, 0.1599933, 0.2893178, 0.115475, 0.03069731, 
    0.04745368, 0.01363528, 0.1095029, 0.1094109, 0.1985691,
  0.05331714, 0.01022557, 0.03350843, 0.0944972, 0.07519346, 0.05543255, 
    0.1004004, 0.09546488, 0.1656577, 0.1657267, 0.07568122, 0.1585592, 
    0.0883006, 0.1307969, 0.08514987, 0.09609042, 0.03096795, 0.01730529, 
    0.0305221, 0.05872228, 0.08309336, 0.09385274, 0.05751324, 0.04402096, 
    0.04440111, 0.05145338, 0.05643681, 0.04693136, 0.03173163,
  4.83455e-10, 1.820294e-09, -4.920086e-08, 0.00694516, 0.18962, 0.1119063, 
    0.0004034677, 0.07465848, 0.1640455, 0.07817236, 0.1080939, 0.04909299, 
    0.04422503, 0.06348839, 0.1048696, 0.0924545, 0.06882021, 0.09853785, 
    0.1083944, 0.09100019, 0.06450238, 0.06431234, 0.2801751, 0.09163656, 
    0.04722457, 0.0275523, 0.09126001, 0.0002689366, -9.841834e-07,
  2.320619e-08, -8.558602e-06, 0.0008394858, 0.0134398, 5.471995e-05, 
    0.05471959, 0.00666531, 0.03805688, 0.03371166, 0.3516038, 0.202147, 
    0.133819, 0.05571898, 0.05565389, 0.06026091, 0.05451833, 0.06554653, 
    0.08430831, 0.1406826, 0.2003403, 0.04392945, 0.2452836, 0.08705884, 
    0.04215289, 0.0324022, 0.02816313, 0.05115698, 0.001092484, -2.191599e-07,
  0.001346745, 0.1033804, 0.0578994, 0.1049289, 0.1103205, 0.07834876, 
    -0.0007790694, 0.01015322, 0.03944318, 0.1629409, 0.2214832, 0.06013142, 
    0.08003972, 0.08703128, 0.117271, 0.2016551, 0.1628957, 0.1537488, 
    0.1733555, 0.1710847, 0.1430083, 0.2351288, 0.1487957, 0.1529619, 
    0.1183737, 0.1093354, 0.08027285, 0.1697861, 0.0110988,
  0.04540534, 0.1341115, 0.2332556, 0.3672571, 0.088314, 0.1277584, 
    0.1523926, 0.002855492, 0.009372668, 0.07193296, 0.2059951, 0.1402712, 
    0.1393084, 0.1190484, 0.2157654, 0.2660365, 0.3759128, 0.2808665, 
    0.1378562, 0.3243479, 0.1715001, 0.04370994, 0.2751694, 0.2662638, 
    0.2295005, 0.1849425, 0.1869819, 0.1782841, 0.2454304,
  0.2797062, 0.3834051, 0.3767775, 0.4740157, 0.360032, 0.3034341, 0.2291215, 
    0.2627288, 0.05748344, 0.1430493, 0.1695995, 0.138932, 0.1721395, 
    0.1510118, 0.20768, 0.2729808, 0.3122781, 0.297151, 0.225253, 0.3824476, 
    0.1519451, 0.2237045, 0.3149571, 0.4741083, 0.2880172, 0.2147115, 
    0.2336303, 0.2068075, 0.2580906,
  0.2452595, 0.2975456, 0.4681497, 0.4494029, 0.5328205, 0.4489366, 
    0.3993375, 0.4318928, 0.4528023, 0.5401641, 0.5965649, 0.2177, 0.3737427, 
    0.2218963, 0.5187092, 0.3564168, 0.3717414, 0.356522, 0.3790037, 
    0.2611632, 0.4508604, 0.3268018, 0.3445675, 0.3821262, 0.3678584, 
    0.08631584, 0.1808617, 0.2318282, 0.2884257,
  0.2961735, 0.2588138, 0.2684998, 0.2977663, 0.4791748, 0.583486, 0.5030707, 
    0.4860266, 0.3582149, 0.5223743, 0.3968601, 0.3746507, 0.4545007, 
    0.4883402, 0.5424464, 0.2390613, 0.3329897, 0.3917136, 0.3167944, 
    0.4694608, 0.3750538, 0.3821275, 0.3837019, 0.2022646, 0.1380083, 
    0.3073516, 0.4563164, 0.2693843, 0.4040635,
  0.3263873, 0.1878324, 0.205175, 0.1931436, 0.1828369, 0.2082339, 0.3448905, 
    0.3886201, 0.3448356, 0.3636495, 0.4024149, 0.3753285, 0.4317653, 
    0.4647708, 0.360778, 0.3809266, 0.365273, 0.4068554, 0.474411, 0.4643713, 
    0.3929923, 0.4173492, 0.3188583, 0.1403706, 0.1225271, 0.05813175, 
    0.16363, 0.2961144, 0.4562216,
  0.2741393, 0.2766001, 0.2790609, 0.2815217, 0.2839826, 0.2864434, 
    0.2889042, 0.2735557, 0.2764733, 0.279391, 0.2823086, 0.2852263, 
    0.2881439, 0.2910616, 0.3499761, 0.3539867, 0.3579974, 0.362008, 
    0.3660186, 0.3700293, 0.3740399, 0.330589, 0.3212, 0.3118109, 0.3024217, 
    0.2930326, 0.2836435, 0.2742544, 0.2721707,
  0.1964493, 0.1756134, 0.1737436, 0.1551869, 0.2062864, 0.1197627, 
    0.1401079, 0.2184672, 0.3470233, 0.2580734, 0.2495293, 0.2743657, 
    0.2972261, 0.00603998, 0.2183052, 0.2074268, 0.1699719, 0.2055443, 
    0.1330387, 0.1270458, 0.2681663, 0.3320297, 0.3425656, 0.1603213, 
    0.2127147, 0.2550266, 0.1799087, 0.1250565, 0.1086068,
  0.197596, 0.1791641, 0.2260954, 0.1320316, 0.123101, 0.4099134, 0.1306313, 
    0.1091583, 0.09675519, 0.09835004, 0.1582346, 0.2258942, 0.08772098, 
    0.153844, 0.3383674, 0.3961423, 0.416913, 0.3761594, 0.4099033, 
    0.3996839, 0.3200346, 0.3915974, 0.403811, 0.4475645, 0.2259504, 
    0.268731, 0.3118015, 0.3128733, 0.2785081,
  0.4581928, 0.4460363, 0.5508847, 0.5463504, 0.5692773, 0.5505208, 
    0.5439765, 0.4162225, 0.4563618, 0.4062298, 0.4153448, 0.351794, 
    0.4919997, 0.4596576, 0.3283384, 0.380347, 0.4602388, 0.4928917, 
    0.4736689, 0.3683442, 0.3967929, 0.4075424, 0.4022471, 0.4317117, 
    0.4435695, 0.4576415, 0.5505866, 0.487666, 0.5234565,
  0.4075976, 0.3899068, 0.4219845, 0.3830773, 0.3724872, 0.4004592, 
    0.4161372, 0.4665379, 0.4423231, 0.4062849, 0.3307438, 0.2909624, 
    0.2602085, 0.2326851, 0.1483667, 0.2693353, 0.3566533, 0.3845947, 
    0.3321277, 0.2854934, 0.2864546, 0.3124329, 0.3191974, 0.1635506, 
    0.03524635, 0.1391837, 0.3270832, 0.4066546, 0.4066773,
  0.2571834, 0.1798055, 0.09653927, 0.2020923, 0.1887957, 0.1558152, 
    0.3071239, 0.2601099, 0.3342882, 0.2404045, 0.2316049, 0.07362498, 
    0.1294946, 0.2393827, 0.2161218, 0.2560845, 0.2504494, 0.2840708, 
    0.3351364, 0.2385806, 0.2236355, 0.244974, 0.147094, 0.0642966, 
    0.03934761, 0.1657092, 0.21167, 0.2184488, 0.216515,
  0.21393, 0.08351663, 0.02670708, 0.1621048, 0.1528331, 0.1244919, 
    0.1833587, 0.1818387, 0.1703848, 0.03143262, 0.01207446, -1.399732e-05, 
    -0.0001159163, 0.09252068, 0.1140106, 0.1230037, 0.06201962, 0.2424715, 
    0.1275369, 0.1575428, 0.1712434, 0.09803787, 0.2099349, 0.008881229, 
    0.01130893, 0.1523885, 0.1673234, 0.09103586, 0.127769,
  0.3722882, 0.01836088, 0.03535307, 0.1307974, 0.03427689, 0.06807066, 
    0.04617714, 0.02524696, 0.1477365, 0.03429144, 0.006069863, 0.0006093311, 
    0.05371297, 0.0450711, 0.08141471, 0.0551208, 0.07602146, 0.04256748, 
    0.02925964, 0.01280172, 0.006619047, 0.0649052, 0.3920956, 0.07913975, 
    0.032482, 0.1379584, 0.02607588, 0.05423534, 0.1411983,
  0.4363245, 0.1473371, 0.05825635, 0.05795556, 0.04455276, 0.0720264, 
    0.05079872, 0.04676757, 0.06840076, 0.1376252, 0.03037629, 0.02575971, 
    0.03783448, 0.02831896, 0.02788622, 0.02016061, 0.01725836, 0.01840636, 
    0.01032263, 0.01130059, 0.04072812, 0.1766147, 0.5169018, 0.01788408, 
    0.03200629, 0.008775471, 0.03482284, 0.04895151, 0.2130336,
  0.04624635, 0.004920914, 0.02211605, 0.09212609, 0.07998607, 0.09355316, 
    0.08795955, 0.05236669, 0.1057342, 0.134315, 0.02499255, 0.08106548, 
    0.02089713, 0.02880002, 0.03535151, 0.03760265, 0.05141114, 0.03240042, 
    0.03537063, 0.04447453, 0.1296999, 0.2027588, 0.1042227, 0.02507394, 
    0.02193318, 0.02774651, 0.04991836, 0.09383617, 0.04212734,
  4.09572e-10, 1.034295e-09, -2.805502e-08, 0.005427914, 0.1930454, 
    0.03169128, -0.001145792, 0.01495105, 0.06746684, 0.05252821, 0.09346981, 
    0.03021235, 0.01852742, 0.02775089, 0.0441549, 0.06782319, 0.04005977, 
    0.06553692, 0.08826501, 0.1135195, 0.06810488, 0.04173541, 0.4205637, 
    0.1450957, 0.01772045, 0.00812762, 0.02491725, 5.090487e-06, -1.303167e-06,
  1.126464e-08, -2.659465e-05, 0.0004927964, 0.0027013, 0.001969294, 
    0.01381158, 0.002556146, 0.02065788, 0.03126235, 0.3033126, 0.1154836, 
    0.06005026, 0.0146198, 0.0203584, 0.02276226, 0.02734466, 0.03445225, 
    0.06256136, 0.07450696, 0.1992554, 0.06664219, 0.2244584, 0.02303253, 
    0.01321496, 0.01327114, 0.009438941, 0.01086589, 0.0004574653, 
    -8.978851e-09,
  8.637906e-05, 0.05226808, 0.02067994, 0.06583545, 0.1103708, 0.06262574, 
    -0.0009021438, 0.006110949, 0.02736166, 0.1596211, 0.1296614, 0.03834147, 
    0.06070448, 0.06510638, 0.08592469, 0.1843604, 0.1615981, 0.1095094, 
    0.1347496, 0.1129832, 0.1366145, 0.2606097, 0.1403811, 0.1330064, 
    0.09620684, 0.06043583, 0.0376974, 0.0923048, 0.005190954,
  0.05017851, 0.1009011, 0.1835128, 0.3705602, 0.04882539, 0.1307899, 
    0.1536792, 0.0007238423, 0.009251376, 0.07429299, 0.2129013, 0.08452237, 
    0.09781707, 0.09047, 0.1945298, 0.2416101, 0.3450738, 0.183194, 
    0.0957031, 0.3422162, 0.1611566, 0.04886898, 0.269301, 0.224121, 
    0.1766248, 0.1864671, 0.1659223, 0.1335766, 0.2065572,
  0.3619078, 0.4153703, 0.3943273, 0.5304432, 0.4067038, 0.322957, 0.2649857, 
    0.2579347, 0.05137523, 0.1677629, 0.1800849, 0.1637965, 0.1134132, 
    0.09881163, 0.1880346, 0.2953367, 0.284372, 0.2770315, 0.1894528, 
    0.4242797, 0.1720562, 0.2191162, 0.2869387, 0.4809535, 0.2844897, 
    0.1777771, 0.2032677, 0.224797, 0.2861321,
  0.2336543, 0.317663, 0.5358354, 0.5366155, 0.5830162, 0.5041826, 0.4476376, 
    0.5183805, 0.5183352, 0.6126224, 0.6579976, 0.2885141, 0.3474219, 
    0.1953798, 0.4451929, 0.3561056, 0.4273041, 0.3362721, 0.3656333, 
    0.2583143, 0.5569189, 0.3384106, 0.3682376, 0.3748274, 0.2652303, 
    0.05669947, 0.1571781, 0.2038139, 0.2704638,
  0.2252824, 0.2064605, 0.2656462, 0.2199684, 0.419539, 0.6019177, 0.5509326, 
    0.5183907, 0.3774772, 0.5196317, 0.4223189, 0.4139326, 0.4650736, 
    0.5511872, 0.5458893, 0.2584654, 0.3302149, 0.3690054, 0.3484801, 
    0.4953603, 0.3590274, 0.3838963, 0.4039947, 0.227838, 0.1351471, 
    0.3177533, 0.4594823, 0.2461729, 0.3720357,
  0.3383981, 0.184031, 0.2186393, 0.1916893, 0.1994989, 0.3000315, 0.3922906, 
    0.4276121, 0.3975418, 0.3884285, 0.4440207, 0.4455808, 0.5020079, 
    0.5175169, 0.4126327, 0.432014, 0.4153073, 0.420986, 0.4917266, 
    0.4836208, 0.4725073, 0.4249388, 0.3316502, 0.1701059, 0.1343814, 
    0.05599986, 0.1601379, 0.2994287, 0.4899018,
  0.2599322, 0.264559, 0.2691857, 0.2738124, 0.2784392, 0.2830659, 0.2876926, 
    0.2731214, 0.2747599, 0.2763983, 0.2780368, 0.2796752, 0.2813137, 
    0.2829521, 0.3402653, 0.3416567, 0.3430483, 0.3444397, 0.3458312, 
    0.3472227, 0.3486142, 0.3029023, 0.2952456, 0.287589, 0.2799323, 
    0.2722757, 0.264619, 0.2569624, 0.2562309,
  0.1671591, 0.1593369, 0.1360452, 0.1417333, 0.1844812, 0.08276465, 
    0.1266507, 0.2420115, 0.3100587, 0.2396021, 0.2025111, 0.1996066, 
    0.2288903, 0.001341635, 0.1830088, 0.1939959, 0.1669385, 0.1975007, 
    0.09991462, 0.09133568, 0.169359, 0.2576498, 0.2779302, 0.158544, 
    0.1355303, 0.2048219, 0.1419754, 0.09872133, 0.09485691,
  0.1776437, 0.1482819, 0.2215777, 0.1242268, 0.06395059, 0.3406869, 
    0.1200564, 0.07653565, 0.0600371, 0.05637943, 0.1001936, 0.1712, 
    0.0532107, 0.1661133, 0.3377734, 0.3611616, 0.3888896, 0.3430797, 
    0.3836075, 0.4263121, 0.3322978, 0.4152088, 0.389869, 0.4578272, 
    0.247113, 0.3166126, 0.2729517, 0.2739686, 0.342815,
  0.4030043, 0.436365, 0.5220006, 0.5256032, 0.5364774, 0.5178574, 0.5351601, 
    0.3977533, 0.4644591, 0.3990282, 0.3697013, 0.304113, 0.483178, 
    0.4100053, 0.3162047, 0.3758873, 0.4345201, 0.5029411, 0.4511426, 
    0.3227057, 0.3710312, 0.3680167, 0.3866054, 0.3975464, 0.3962184, 
    0.4452865, 0.5339922, 0.4680285, 0.4835688,
  0.3968134, 0.3662696, 0.3866777, 0.3421084, 0.3518145, 0.387586, 0.3923908, 
    0.3967181, 0.4278628, 0.376427, 0.2870823, 0.2712697, 0.2260848, 
    0.2153994, 0.1621054, 0.281576, 0.3201092, 0.3429743, 0.2845443, 
    0.2499757, 0.2465542, 0.2857747, 0.3073004, 0.1464439, 0.03258263, 
    0.1381867, 0.3425344, 0.3917302, 0.3875696,
  0.2220544, 0.124406, 0.06395772, 0.1839254, 0.1753564, 0.1244187, 
    0.2521741, 0.2550948, 0.2341715, 0.2131329, 0.1579732, 0.06893048, 
    0.09236006, 0.1839923, 0.2224606, 0.1994811, 0.1700125, 0.181686, 
    0.2847351, 0.2160982, 0.2213181, 0.2315282, 0.1148573, 0.076865, 
    0.05583912, 0.1435631, 0.206002, 0.1860574, 0.1984505,
  0.1188089, 0.06028087, 0.02142491, 0.1292897, 0.1227154, 0.05971668, 
    0.1456863, 0.06809344, 0.06338602, 0.009494971, 0.01068085, 0.0001236767, 
    -0.001257197, 0.04511423, 0.08699343, 0.08531652, 0.04192407, 0.2158051, 
    0.1594928, 0.1174516, 0.07898919, 0.03038072, 0.08685091, 0.03362761, 
    0.009505811, 0.1087546, 0.1495125, 0.04196894, 0.08333527,
  0.1285941, 0.05469676, 0.02626099, 0.05446833, 0.007281716, 0.02318974, 
    0.01472314, 0.005316012, 0.0678887, 0.01091304, 0.004589128, 
    0.0002867484, 0.01184485, 0.01746948, 0.0560234, 0.02975718, 0.03615301, 
    0.01831684, 0.003950658, 0.001572914, 0.0004349705, 0.01950586, 
    0.1457282, 0.2572041, 0.02738607, 0.1342291, 0.003379353, 0.01505051, 
    0.04027975,
  0.1569877, 0.1102583, 0.04560438, 0.07862423, 0.01289032, 0.03518826, 
    0.01943249, 0.01940366, 0.02194725, 0.02609684, 0.01187463, 0.006386783, 
    0.01322275, 0.008358669, 0.005092793, 0.007953777, 0.003373591, 
    0.003325397, 0.001034662, 0.001543077, 0.01001035, 0.05199187, 0.3044199, 
    0.0130975, 0.02276292, 0.006638455, 0.001392147, 0.007416672, 0.06598905,
  0.04813514, 0.003774765, 0.01580145, 0.08488618, 0.03811067, 0.02230849, 
    0.02590121, 0.01498063, 0.07408676, 0.1021432, 0.01061875, 0.01378495, 
    0.005236939, 0.005831265, 0.006911149, 0.005442104, 0.009587845, 
    0.01515065, 0.01054326, 0.01615387, 0.07356109, 0.3360127, 0.3372579, 
    0.01961549, 0.01099315, 0.007630254, 0.03192146, 0.05064021, 0.03956069,
  3.766392e-10, 8.029873e-10, 1.904602e-09, 0.007742939, 0.1558467, 
    0.0102294, -0.002431551, 0.003622717, 0.02377915, 0.01829637, 0.05179852, 
    0.007622321, 0.007354917, 0.009200797, 0.01845127, 0.03708182, 
    0.02453663, 0.03584428, 0.05749102, 0.08169331, 0.02894446, 0.01007245, 
    0.4058078, 0.1240037, 0.00620123, 0.0009797951, 0.00774981, 
    -6.679772e-06, -7.005731e-07,
  6.626438e-09, -3.910705e-05, 0.0001140897, 0.000284827, 0.002299913, 
    0.00447365, 0.008099901, 0.01355613, 0.02707965, 0.2117262, 0.06826657, 
    0.02423951, 0.004185457, 0.003114124, 0.008047477, 0.008870535, 
    0.0172129, 0.04018059, 0.04036919, 0.1504436, 0.03301287, 0.2014328, 
    0.004350158, -0.002150709, 0.006115498, 0.002359413, 0.002947934, 
    0.0001255274, 1.448459e-08,
  -2.246221e-05, 0.03393717, 0.0107317, 0.03156473, 0.1023173, 0.04291854, 
    -0.001191007, 0.004616911, 0.01840592, 0.1493467, 0.08682495, 0.0215985, 
    0.04498138, 0.04697155, 0.06758024, 0.1700984, 0.142736, 0.05391541, 
    0.07723895, 0.08758091, 0.1310548, 0.2434424, 0.1276856, 0.08675961, 
    0.06498419, 0.04325981, 0.01629069, 0.03123349, 0.003162462,
  0.03096344, 0.05561654, 0.1265428, 0.3698063, 0.02977142, 0.1123425, 
    0.1546203, -9.245434e-05, 0.003510519, 0.0762303, 0.2004361, 0.05830546, 
    0.07191716, 0.06912187, 0.1686492, 0.1938049, 0.2980057, 0.1437848, 
    0.07826014, 0.3445069, 0.1386903, 0.04936612, 0.2458054, 0.2051386, 
    0.1384647, 0.1572585, 0.1410133, 0.1002294, 0.1834565,
  0.3600582, 0.4234369, 0.4311052, 0.5406201, 0.4055424, 0.334417, 0.2121654, 
    0.2359436, 0.04927637, 0.1722136, 0.1709463, 0.1891276, 0.07940711, 
    0.06910095, 0.1692906, 0.2920748, 0.2748877, 0.202992, 0.1458549, 
    0.4502234, 0.1562345, 0.1980024, 0.2577779, 0.5099761, 0.2808039, 
    0.1553794, 0.1775564, 0.2019573, 0.2895324,
  0.1958151, 0.3519508, 0.5332105, 0.5871629, 0.6243297, 0.5597308, 
    0.4885854, 0.5742685, 0.5785697, 0.6629868, 0.6935546, 0.3966273, 
    0.3052331, 0.1690506, 0.380237, 0.3714654, 0.4802704, 0.3052568, 
    0.3704222, 0.2633045, 0.6620691, 0.3655066, 0.4119791, 0.3352437, 
    0.2089813, 0.03586392, 0.1338143, 0.1671967, 0.2204611,
  0.1686864, 0.1580749, 0.2827533, 0.1438487, 0.3352218, 0.5711241, 
    0.6001523, 0.4977697, 0.40953, 0.5290152, 0.466361, 0.4463482, 0.4971228, 
    0.6053718, 0.5455436, 0.2806357, 0.3514681, 0.3303025, 0.3631196, 
    0.4766502, 0.3384381, 0.4162162, 0.4427432, 0.2559977, 0.1602009, 
    0.3239726, 0.4669967, 0.2130135, 0.309241,
  0.3934458, 0.2410979, 0.2465289, 0.2164482, 0.279902, 0.3980811, 0.4350488, 
    0.4352747, 0.4096978, 0.4613177, 0.5200741, 0.5338762, 0.5966712, 
    0.5874131, 0.4848062, 0.4813237, 0.4510918, 0.4499626, 0.5524045, 
    0.5134574, 0.5454012, 0.4358484, 0.3668313, 0.1967689, 0.1276935, 
    0.05514599, 0.156884, 0.2867319, 0.5299937,
  0.2413553, 0.2457491, 0.2501429, 0.2545367, 0.2589305, 0.2633243, 
    0.2677181, 0.2374328, 0.2388137, 0.2401946, 0.2415756, 0.2429565, 
    0.2443374, 0.2457184, 0.3123495, 0.3110401, 0.3097307, 0.3084214, 
    0.307112, 0.3058026, 0.3044932, 0.2628917, 0.2584263, 0.253961, 
    0.2494956, 0.2450303, 0.2405649, 0.2360995, 0.2378402,
  0.1237733, 0.119131, 0.09746015, 0.1178758, 0.1302703, 0.05724706, 
    0.1054259, 0.2042444, 0.2355677, 0.1630632, 0.134599, 0.109778, 0.127433, 
    -0.001275278, 0.1213762, 0.192555, 0.15519, 0.1494461, 0.07709563, 
    0.06003442, 0.1090377, 0.1783567, 0.2241002, 0.1345991, 0.07876511, 
    0.1239592, 0.09744263, 0.06238403, 0.07726856,
  0.1615579, 0.1208284, 0.1679824, 0.09368762, 0.03324252, 0.2874543, 
    0.1115851, 0.05145468, 0.03758857, 0.03577257, 0.05808907, 0.1148174, 
    0.03782226, 0.1683619, 0.3290116, 0.3082732, 0.3498842, 0.3160433, 
    0.3331759, 0.4029674, 0.3091701, 0.3980691, 0.3854993, 0.4144874, 
    0.2442507, 0.3315334, 0.2349494, 0.2307649, 0.2512008,
  0.3418134, 0.3984022, 0.4613515, 0.428656, 0.4712443, 0.4671543, 0.5017993, 
    0.3297498, 0.4188972, 0.3692061, 0.3235656, 0.2648485, 0.4329116, 
    0.3594311, 0.2786577, 0.3583169, 0.4032779, 0.4736501, 0.4150547, 
    0.2722552, 0.3266056, 0.3227701, 0.3344747, 0.326654, 0.3483474, 
    0.4362102, 0.4759639, 0.4087969, 0.442836,
  0.3536896, 0.3156689, 0.3467739, 0.319431, 0.3445944, 0.3486541, 0.3589221, 
    0.332779, 0.3912367, 0.3301038, 0.2455429, 0.2265404, 0.1851157, 
    0.1838138, 0.1728801, 0.2678811, 0.2713386, 0.2932153, 0.2329772, 
    0.2088121, 0.20927, 0.2537006, 0.2618719, 0.1200911, 0.03247079, 
    0.1451021, 0.3209433, 0.3665716, 0.3629497,
  0.1770683, 0.08972584, 0.04178031, 0.1552711, 0.1484438, 0.1039577, 
    0.2175051, 0.2023375, 0.1539004, 0.1297781, 0.09073787, 0.04964337, 
    0.07493901, 0.161166, 0.2142111, 0.1534773, 0.1138162, 0.1270104, 
    0.2321728, 0.2018552, 0.2062384, 0.1914811, 0.1022443, 0.09224037, 
    0.05851471, 0.1200767, 0.1890777, 0.1714785, 0.173014,
  0.06111779, 0.02925526, 0.01673814, 0.06830132, 0.07818629, 0.03440337, 
    0.09776272, 0.03473271, 0.02782741, 0.007121762, 0.006066083, 
    0.0001583579, -0.0002513955, 0.02190304, 0.06808715, 0.05209108, 
    0.02970091, 0.1832049, 0.1788364, 0.07253838, 0.03808013, 0.01249322, 
    0.03392202, 0.02954341, 0.00558423, 0.08053851, 0.1083483, 0.0212618, 
    0.04387847,
  0.04658407, 0.06908114, 0.01612704, 0.01623482, 0.0002687576, 0.004235826, 
    0.005147396, 0.002028056, 0.03113133, 0.01306324, 0.003351977, 
    4.317342e-05, 0.003818206, 0.005680013, 0.03223083, 0.00839876, 
    0.01023147, 0.003630346, 0.000427075, 0.0003368612, 0.0001676328, 
    0.007374894, 0.05317847, 0.1357072, 0.02277612, 0.1288387, 0.0007862365, 
    0.005626977, 0.01311534,
  0.05535349, 0.02728834, 0.03699637, 0.07639773, 0.006394776, 0.01397339, 
    0.007677992, 0.007602585, 0.003780813, 0.005697615, 0.005697483, 
    0.001926943, 0.003240335, 0.002100912, 0.0009030497, 0.003518493, 
    0.00127009, 0.001068797, 0.0003951291, 0.0006793612, 0.004129925, 
    0.01904822, 0.1056022, 0.01313779, 0.02228859, 0.006246326, 
    -0.0005353654, 0.002284283, 0.01994056,
  0.03197328, 0.003296343, 0.01327315, 0.07757155, 0.007554688, 0.003741932, 
    0.01385672, 0.003821486, 0.06038788, 0.08784147, 0.00647895, 0.004997042, 
    0.0007584339, 0.001867543, 0.003212937, 0.001664098, 0.00202236, 
    0.002527213, 0.002115459, 0.002324461, 0.02216112, 0.1570764, 0.1537751, 
    0.01989183, 0.006939453, 0.002887809, 0.01955502, 0.009572187, 0.005489462,
  3.608751e-10, 7.396477e-10, 5.586846e-09, 0.009561745, 0.1030544, 
    0.002692633, -0.002984795, 0.001605222, 0.01101797, 0.003677285, 
    0.02133772, 0.002116511, 0.003934096, 0.001652918, 0.005764663, 
    0.01433888, 0.01146827, 0.01290602, 0.02469222, 0.0287823, 0.01251694, 
    0.001981381, 0.3110171, 0.08583355, 0.002537632, 0.0001491538, 
    0.003751416, -5.933977e-06, -2.98222e-07,
  5.39517e-09, -3.132542e-05, 4.147915e-05, -7.07883e-06, 0.0006229257, 
    0.002258472, 0.01442311, 0.006111373, 0.02586442, 0.1212824, 0.03451226, 
    0.008126339, 0.0009268412, 0.0007896933, 0.001646352, 0.003713895, 
    0.008661322, 0.02243654, 0.0218191, 0.09838861, 0.01376934, 0.1480551, 
    0.00150987, -0.002759791, 0.00524537, 0.0004059855, 0.001395832, 
    6.541501e-05, 2.072997e-08,
  -1.696758e-05, 0.02561901, 0.00630288, 0.01766403, 0.09584299, 0.03698951, 
    -0.001172002, 0.004858378, 0.01697341, 0.1368215, 0.0637808, 0.01175204, 
    0.03021056, 0.03131335, 0.06146929, 0.1314895, 0.08707878, 0.02506959, 
    0.04484317, 0.05599006, 0.1205262, 0.2112171, 0.1096554, 0.05980613, 
    0.04152729, 0.02622521, 0.006449992, 0.01315726, 0.002184697,
  0.01912138, 0.02653987, 0.08524503, 0.3549975, 0.0168048, 0.07854553, 
    0.1507193, -0.0002525654, 0.001894266, 0.06075474, 0.1887159, 0.0448736, 
    0.05433477, 0.05273613, 0.14476, 0.143303, 0.2392555, 0.115489, 
    0.05841941, 0.3284098, 0.1199277, 0.04448791, 0.2488956, 0.1928835, 
    0.1053391, 0.114163, 0.1054946, 0.06740226, 0.1385257,
  0.2971573, 0.4119613, 0.4229056, 0.5013359, 0.3871063, 0.3210599, 
    0.1464355, 0.2097721, 0.05525351, 0.1585408, 0.1515709, 0.2151684, 
    0.05198925, 0.05358978, 0.1556377, 0.2568977, 0.2312133, 0.1557195, 
    0.1115982, 0.4506868, 0.1265436, 0.1578457, 0.2281803, 0.5288466, 
    0.2195338, 0.1301432, 0.1453134, 0.1605709, 0.2509402,
  0.1536723, 0.3660243, 0.5095025, 0.6114314, 0.6573802, 0.5698332, 
    0.5520449, 0.5845751, 0.6214714, 0.6726038, 0.6915962, 0.4657184, 
    0.2718857, 0.1685933, 0.326215, 0.3579521, 0.5119966, 0.2672507, 
    0.3761796, 0.2709508, 0.7253869, 0.3804417, 0.423663, 0.3190041, 
    0.1700479, 0.02714604, 0.1115354, 0.1293882, 0.1661793,
  0.1387348, 0.1228657, 0.2896219, 0.08774991, 0.2676393, 0.5114137, 
    0.6078016, 0.4774889, 0.4289094, 0.5388077, 0.5275605, 0.5241186, 
    0.564795, 0.6326849, 0.5336748, 0.3279937, 0.3686315, 0.3033898, 
    0.3598619, 0.4162211, 0.4016982, 0.494203, 0.5172101, 0.3035484, 
    0.2678699, 0.2725253, 0.4748433, 0.154365, 0.2641606,
  0.4304306, 0.2409367, 0.2774612, 0.2693211, 0.3568773, 0.4671021, 
    0.4896742, 0.5049108, 0.4643847, 0.5430439, 0.5995696, 0.6239447, 
    0.68503, 0.6438861, 0.5661306, 0.5798475, 0.5156832, 0.526096, 0.6121191, 
    0.5602554, 0.5984119, 0.4215716, 0.4059725, 0.2810981, 0.1168975, 
    0.05906913, 0.141194, 0.2542899, 0.5496026,
  0.1919879, 0.1961426, 0.2002974, 0.2044521, 0.2086068, 0.2127616, 
    0.2169163, 0.1806251, 0.182458, 0.1842909, 0.1861238, 0.1879567, 
    0.1897896, 0.1916225, 0.262481, 0.2593888, 0.2562965, 0.2532043, 
    0.250112, 0.2470197, 0.2439275, 0.2013459, 0.1984505, 0.1955552, 
    0.1926598, 0.1897644, 0.186869, 0.1839736, 0.1886641,
  0.08977295, 0.08338043, 0.07232963, 0.09202436, 0.08973078, 0.03988553, 
    0.08316505, 0.1516247, 0.1687796, 0.1089627, 0.08059882, 0.05953251, 
    0.06714882, -0.001117963, 0.08721436, 0.1570205, 0.1402488, 0.103773, 
    0.05320831, 0.04734855, 0.0690937, 0.125675, 0.1757948, 0.09918596, 
    0.05058496, 0.08598279, 0.07333684, 0.04195526, 0.0482372,
  0.1519589, 0.0872019, 0.1092668, 0.0699826, 0.01913559, 0.2372788, 
    0.1000145, 0.0341235, 0.02583854, 0.02623501, 0.03777967, 0.07547255, 
    0.02485518, 0.1528166, 0.3034903, 0.2492948, 0.3124862, 0.2699305, 
    0.2720036, 0.3386228, 0.2643999, 0.3596608, 0.3763759, 0.3579673, 
    0.2220209, 0.3182829, 0.204912, 0.1907671, 0.1790772,
  0.2815298, 0.3278972, 0.3669724, 0.3304256, 0.3923923, 0.3882229, 
    0.4248041, 0.2485741, 0.3444009, 0.3191365, 0.2583166, 0.2308176, 
    0.351993, 0.3092364, 0.2237822, 0.3076864, 0.357013, 0.4097916, 
    0.3438573, 0.2237006, 0.2727647, 0.2535635, 0.2661563, 0.232512, 
    0.3064843, 0.410523, 0.3991661, 0.326373, 0.3575052,
  0.2871912, 0.2465631, 0.2771, 0.2696935, 0.301932, 0.2947983, 0.2949452, 
    0.2670682, 0.3352093, 0.2643281, 0.1939913, 0.169336, 0.1435664, 
    0.1338331, 0.1536001, 0.2190838, 0.2088449, 0.2227002, 0.1751873, 
    0.1601952, 0.1577122, 0.2025118, 0.1907632, 0.09321326, 0.02875728, 
    0.1226655, 0.2699602, 0.3047794, 0.3015577,
  0.1386926, 0.06490013, 0.02699516, 0.1304068, 0.1154565, 0.07777353, 
    0.1781797, 0.142907, 0.1014797, 0.07499395, 0.06665036, 0.03147579, 
    0.05284481, 0.134371, 0.1890482, 0.109502, 0.08198481, 0.09150238, 
    0.1903406, 0.1766773, 0.1621757, 0.1471285, 0.07704201, 0.09222872, 
    0.0569813, 0.0956036, 0.1518291, 0.1349722, 0.1377561,
  0.03863729, 0.01508103, 0.01314734, 0.03776464, 0.04225764, 0.01757729, 
    0.06675944, 0.023601, 0.01598536, 0.007684845, 0.002955228, 0.0001636026, 
    -0.0002770052, 0.007566546, 0.05293655, 0.02917614, 0.02006173, 0.160818, 
    0.1416086, 0.04200594, 0.01728609, 0.006379275, 0.01714339, 0.01642729, 
    0.003302263, 0.05002736, 0.07974781, 0.01271326, 0.02806161,
  0.02235764, 0.05900142, 0.009841526, 0.007681513, -0.001475594, 
    0.001146712, 0.001804297, 0.001114804, 0.01740567, 0.004025547, 
    0.003017236, -9.732441e-06, 0.001677334, 0.002512185, 0.009545406, 
    0.002202187, 0.002819524, 0.0006782649, 0.0001796866, 0.0001008257, 
    9.093282e-05, 0.003791743, 0.02388521, 0.07487309, 0.01771392, 0.110423, 
    0.0004198321, 0.003050014, 0.005958654,
  0.02775498, 0.008887235, 0.03518863, 0.06641645, 0.003902785, 0.006078506, 
    0.002724115, 0.002935897, 0.001534339, 0.002843217, 0.002709416, 
    0.001084418, 0.0004603384, 0.000651343, 0.0004637411, 0.001129158, 
    0.0004927611, 0.0004233939, 0.0002238004, 0.0003877663, 0.002296613, 
    0.009381765, 0.05242557, 0.01141411, 0.02513922, 0.006070057, 
    -8.902788e-05, 0.001173304, 0.009224196,
  0.01367496, 0.001891338, 0.02405174, 0.06498244, 0.002227729, 0.001405851, 
    0.008066555, 0.001874525, 0.04547701, 0.08102824, 0.003913964, 
    0.002682846, 0.0002864359, 0.0009621439, 0.001738595, 0.0008295776, 
    0.0009509445, 0.0006873034, 0.0009624609, 0.0009377984, 0.005574091, 
    0.05078271, 0.06708875, 0.01802217, 0.006097042, 0.000969499, 
    0.008696512, 0.003518502, 0.001749801,
  3.641636e-10, 7.216023e-10, 5.451312e-09, 0.00908844, 0.06331576, 
    0.001210301, -0.002944595, 0.0009804657, 0.005207689, 0.001400318, 
    0.009045843, 0.000672636, 0.001739838, 0.0002744297, 0.0013594, 
    0.009838272, 0.006315158, 0.004322939, 0.007722219, 0.01179121, 
    0.007231158, 0.0006540162, 0.2304986, 0.06480266, 0.001032271, 
    4.909309e-05, 0.002242594, -4.772451e-06, -1.027048e-07,
  5.049552e-09, -1.40952e-05, 2.163189e-05, 6.576569e-05, 0.0002570072, 
    0.001477626, 0.01539491, 0.002847709, 0.02655007, 0.06407181, 0.01378958, 
    0.003358876, 0.0004426814, 0.0003901225, 0.0007447689, 0.001550713, 
    0.003783095, 0.0110214, 0.01529071, 0.04724915, 0.006249434, 0.09917301, 
    0.0008321489, -0.002113747, 0.003421244, 0.0001605928, 0.0008444406, 
    4.153812e-05, 2.222372e-08,
  -1.730525e-05, 0.02305232, 0.004401125, 0.01198461, 0.08654986, 0.03544855, 
    0.0005813308, 0.004737566, 0.01604476, 0.1053998, 0.0507196, 0.006858109, 
    0.01792331, 0.01939917, 0.0296834, 0.08083848, 0.04224104, 0.01299159, 
    0.0261595, 0.03369237, 0.1027746, 0.1910182, 0.09598775, 0.036673, 
    0.02787093, 0.01022911, 0.003020856, 0.007109602, 0.0008017233,
  0.01214695, 0.01621523, 0.05731766, 0.3380861, 0.008564504, 0.0562239, 
    0.1369373, 0.0003444396, 0.0010118, 0.0540707, 0.170327, 0.03564075, 
    0.04299188, 0.03763031, 0.1139317, 0.1064159, 0.1858602, 0.07756843, 
    0.04032495, 0.3100922, 0.09885097, 0.03727061, 0.2162181, 0.1698429, 
    0.07481931, 0.07468598, 0.06843626, 0.04718074, 0.103306,
  0.2330069, 0.3800283, 0.3675947, 0.4320961, 0.3210758, 0.2642105, 
    0.1061969, 0.1793963, 0.06451605, 0.1586529, 0.13426, 0.2291507, 
    0.0311833, 0.04180558, 0.1355289, 0.202644, 0.1892008, 0.1165281, 
    0.08203766, 0.4215051, 0.09172265, 0.1119141, 0.2036948, 0.5101409, 
    0.1654953, 0.1077462, 0.1121237, 0.1134587, 0.1828556,
  0.1051572, 0.3708309, 0.4426489, 0.5956678, 0.6492205, 0.5229904, 
    0.5627642, 0.5858094, 0.6372809, 0.6647757, 0.6760023, 0.5068935, 
    0.2493069, 0.1924542, 0.273247, 0.3100196, 0.5334129, 0.233243, 0.350093, 
    0.2894395, 0.7506665, 0.3524593, 0.3896574, 0.3239651, 0.1440587, 
    0.02076077, 0.09521865, 0.0964536, 0.1157709,
  0.1132278, 0.09411722, 0.310203, 0.05283054, 0.211038, 0.4283941, 
    0.5518106, 0.4367782, 0.4400615, 0.5394977, 0.6499047, 0.5611554, 
    0.7330179, 0.542016, 0.4972473, 0.3821548, 0.3428927, 0.2606349, 0.35322, 
    0.353485, 0.4339337, 0.5935428, 0.6201833, 0.3650418, 0.3842383, 
    0.2241543, 0.4677894, 0.1083072, 0.2290492,
  0.4457555, 0.2085423, 0.3132439, 0.3799205, 0.475102, 0.5175037, 0.521511, 
    0.5493459, 0.5172008, 0.5649617, 0.626256, 0.6793005, 0.6963999, 
    0.6999096, 0.6231527, 0.6270577, 0.5905939, 0.5848845, 0.6311926, 
    0.6197386, 0.6390648, 0.3764116, 0.4345294, 0.3754008, 0.09107185, 
    0.05795079, 0.1307508, 0.2034852, 0.5505656,
  0.1269742, 0.130211, 0.1334478, 0.1366846, 0.1399213, 0.1431581, 0.1463949, 
    0.1144344, 0.1161147, 0.1177951, 0.1194754, 0.1211557, 0.1228361, 
    0.1245164, 0.1693905, 0.1664011, 0.1634117, 0.1604223, 0.1574329, 
    0.1544436, 0.1514542, 0.1264253, 0.1244975, 0.1225698, 0.1206421, 
    0.1187143, 0.1167866, 0.1148588, 0.1243847,
  0.06768899, 0.05846855, 0.05410823, 0.07840906, 0.06202214, 0.02741074, 
    0.06036767, 0.1042019, 0.1170595, 0.07437953, 0.05270241, 0.03547117, 
    0.04347681, -0.0005314479, 0.06500989, 0.1267511, 0.1230155, 0.08233829, 
    0.03789707, 0.03520057, 0.04265017, 0.08969368, 0.1426076, 0.071623, 
    0.03519639, 0.06548126, 0.04962974, 0.03006, 0.0313027,
  0.1313293, 0.06566186, 0.07762128, 0.05353642, 0.01167398, 0.1947785, 
    0.09400997, 0.02452366, 0.01918153, 0.01903822, 0.02517938, 0.05224482, 
    0.01670252, 0.1345188, 0.2474739, 0.1867009, 0.2416871, 0.2144691, 
    0.2050009, 0.2579368, 0.2058363, 0.2886556, 0.3111693, 0.2937823, 
    0.2102606, 0.2692879, 0.1663629, 0.1449865, 0.1408409,
  0.2096028, 0.2271037, 0.2594799, 0.2342924, 0.2892938, 0.293272, 0.3333547, 
    0.1789786, 0.2684715, 0.2418715, 0.1892656, 0.1834091, 0.2762231, 
    0.2478845, 0.1638538, 0.2289662, 0.2853892, 0.3312563, 0.2657174, 
    0.1706268, 0.2025252, 0.1655312, 0.1795718, 0.1517191, 0.2449867, 
    0.3506757, 0.3203267, 0.2474867, 0.260444,
  0.2155466, 0.1871351, 0.2116191, 0.2138367, 0.2372231, 0.2385119, 
    0.2231439, 0.1881965, 0.2528364, 0.1911125, 0.1331717, 0.1133911, 
    0.09609929, 0.08965279, 0.1342054, 0.1541915, 0.1386002, 0.1473169, 
    0.1167429, 0.111218, 0.1063333, 0.1471206, 0.1355733, 0.07119741, 
    0.0204811, 0.09428672, 0.205855, 0.2301118, 0.2312735,
  0.1012098, 0.03981368, 0.01966465, 0.0979614, 0.07152138, 0.05235949, 
    0.1242238, 0.09790744, 0.06561363, 0.04324797, 0.04418512, 0.02251602, 
    0.03504166, 0.1031515, 0.1606084, 0.06913503, 0.0565342, 0.06457677, 
    0.1346282, 0.1224664, 0.1075814, 0.09767147, 0.04885868, 0.09014456, 
    0.04898335, 0.0632998, 0.1071083, 0.08701587, 0.09225206,
  0.02575662, 0.00917195, 0.008459713, 0.0181332, 0.0233482, 0.009677289, 
    0.04395099, 0.01841972, 0.0110576, 0.005954644, 0.001675791, 
    6.564273e-05, -0.0005200225, 0.003429961, 0.03500534, 0.01456276, 
    0.01214923, 0.1198855, 0.08096528, 0.02190838, 0.007724198, 0.004174773, 
    0.01101665, 0.01019682, 0.001924445, 0.02612434, 0.05121789, 0.005714073, 
    0.01417549,
  0.01341294, 0.04012731, 0.004788083, 0.004331099, -0.001492656, 
    0.0006635155, 0.0006633734, 0.0007311994, 0.0112161, 0.002264672, 
    0.002462705, 1.610875e-05, 0.0009786966, 0.0008121135, 0.003674502, 
    0.001091953, 0.001225895, 0.0002353644, 0.0001106133, 4.977048e-05, 
    5.890991e-05, 0.002371266, 0.01363152, 0.04904034, 0.01231891, 
    0.08894722, 0.0002813716, 0.002018926, 0.003516652,
  0.0176484, 0.003281124, 0.03341789, 0.05224038, 0.001991973, 0.002411236, 
    0.0009167496, 0.001137357, 0.0009486104, 0.00213296, 0.0008533529, 
    0.0006006806, 0.0001694093, 0.0002518781, 0.0002666835, 0.000383076, 
    0.0002072983, 0.0002013185, 0.0001485703, 0.000259533, 0.001504515, 
    0.005778768, 0.03326415, 0.01017443, 0.02379522, 0.004705191, 
    0.0001115052, 0.000748139, 0.005715812,
  0.005953155, 0.003341896, 0.02141246, 0.05345943, 0.001078754, 
    0.0007256725, 0.003861549, 0.0009115067, 0.03898346, 0.07927722, 
    0.001907741, 0.001711945, 0.0001694878, 0.0005824803, 0.0008406078, 
    0.0005072162, 0.0005691446, 0.0003720178, 0.0005939347, 0.0005533276, 
    0.003043436, 0.02567954, 0.03374838, 0.01517233, 0.004721889, 
    0.0003950671, 0.003300996, 0.001819686, 0.0008577746,
  3.662507e-10, 7.179639e-10, 5.197238e-09, 0.01225816, 0.03417275, 
    0.0007818632, -0.002456997, 0.0006857647, 0.002633881, 0.0008349462, 
    0.004049969, 0.0002753199, 0.0007169443, 7.35414e-05, 0.0004997913, 
    0.005875626, 0.002995814, 0.001561141, 0.002739308, 0.00548012, 
    0.003305343, 0.0004228088, 0.1865592, 0.04963256, 0.0003538309, 
    2.686611e-05, 0.001531067, -3.842205e-06, -2.509623e-08,
  4.97982e-09, -8.036515e-06, 1.39231e-05, 9.632119e-05, 0.000149906, 
    0.001099016, 0.01052408, 0.00162239, 0.02490756, 0.03441767, 0.005497428, 
    0.001498915, 0.0003005996, 0.0002558602, 0.0004895109, 0.0007882583, 
    0.001729581, 0.004822026, 0.008301984, 0.02133331, 0.003479553, 
    0.06962442, 0.0005609595, -0.001736611, 0.001831955, 0.0001027785, 
    0.0005861325, 2.985856e-05, 2.226574e-08,
  -1.865054e-05, 0.01715528, 0.003334602, 0.008297524, 0.07250834, 
    0.03260745, 0.004489292, 0.006306563, 0.01808571, 0.07434664, 0.03927541, 
    0.004244138, 0.008616135, 0.01000255, 0.01406352, 0.04885665, 0.0244862, 
    0.00650225, 0.01619771, 0.0203553, 0.0847083, 0.1600287, 0.08039992, 
    0.02307357, 0.01611412, 0.004281273, 0.001799969, 0.004820894, 
    0.0002662688,
  0.009673987, 0.0107502, 0.04213531, 0.314823, 0.005044912, 0.04089393, 
    0.1186429, 0.001131749, 0.0004905806, 0.04603474, 0.1494428, 0.02693705, 
    0.03126364, 0.02581424, 0.08228093, 0.07223514, 0.1299468, 0.05464566, 
    0.02451449, 0.2852357, 0.08158814, 0.03107214, 0.1793024, 0.1430683, 
    0.04947473, 0.04097518, 0.04048054, 0.03018273, 0.06865123,
  0.1650739, 0.3244714, 0.3066755, 0.3524467, 0.2525296, 0.2113803, 
    0.07996403, 0.1617051, 0.08788125, 0.1521554, 0.1197328, 0.2447168, 
    0.02029783, 0.03298118, 0.1068923, 0.1565464, 0.1414523, 0.08700427, 
    0.05592097, 0.3995564, 0.07097086, 0.08017437, 0.1697365, 0.4682165, 
    0.1369422, 0.08854397, 0.07905908, 0.07472271, 0.1194555,
  0.06768575, 0.3776715, 0.3754892, 0.5329574, 0.5912884, 0.44122, 0.5287393, 
    0.5267615, 0.5877048, 0.6184772, 0.6485788, 0.5648176, 0.2552349, 
    0.2196965, 0.2288025, 0.2616693, 0.5454652, 0.205078, 0.314016, 
    0.2882389, 0.7471532, 0.3169783, 0.2853097, 0.3742566, 0.1293488, 
    0.01574215, 0.07291498, 0.06660661, 0.07754184,
  0.08847167, 0.06727027, 0.3347591, 0.03753805, 0.1668736, 0.3247738, 
    0.488885, 0.4462537, 0.4650187, 0.5856463, 0.701874, 0.5166007, 0.800616, 
    0.4076243, 0.4214421, 0.3552061, 0.3183624, 0.1888989, 0.3264188, 
    0.2882925, 0.4288936, 0.6497742, 0.5767107, 0.4818686, 0.3648832, 
    0.1716761, 0.4456332, 0.08145972, 0.1888998,
  0.4279202, 0.1857562, 0.3572384, 0.4229821, 0.5147824, 0.5345687, 
    0.5068419, 0.5333613, 0.5340725, 0.510841, 0.5961705, 0.5866437, 
    0.626574, 0.6472, 0.6047645, 0.5739014, 0.5491754, 0.5297946, 0.5424982, 
    0.5136518, 0.5594766, 0.3271902, 0.4226868, 0.462023, 0.07689729, 
    0.04725762, 0.1071445, 0.1721952, 0.516846,
  0.09840515, 0.1005122, 0.1026192, 0.1047263, 0.1068333, 0.1089403, 
    0.1110474, 0.08068121, 0.08075473, 0.08082823, 0.08090176, 0.08097526, 
    0.08104879, 0.08112229, 0.1060644, 0.1049133, 0.1037623, 0.1026113, 
    0.1014603, 0.1003092, 0.09915821, 0.08842559, 0.08739607, 0.08636655, 
    0.08533703, 0.08430751, 0.08327799, 0.08224846, 0.09671953,
  0.05667485, 0.04202874, 0.0433706, 0.07041144, 0.04071259, 0.01936425, 
    0.04098346, 0.07632983, 0.07411613, 0.05364798, 0.03419692, 0.02575869, 
    0.0310476, 3.918639e-05, 0.05238031, 0.1038105, 0.1122577, 0.06782953, 
    0.03059717, 0.02964253, 0.02965957, 0.06763597, 0.121735, 0.05536554, 
    0.02468683, 0.05435775, 0.03965605, 0.02317897, 0.02041086,
  0.1228089, 0.05396422, 0.06521551, 0.0450487, 0.008885532, 0.1609713, 
    0.08174303, 0.02034547, 0.01462736, 0.01588092, 0.018833, 0.04394822, 
    0.01195049, 0.1195679, 0.2029461, 0.1454916, 0.1851989, 0.1726687, 
    0.1568782, 0.1957763, 0.1694094, 0.2275925, 0.252049, 0.2422239, 
    0.1797607, 0.2210702, 0.1332668, 0.1153344, 0.1187776,
  0.1593211, 0.1703401, 0.1941697, 0.1800316, 0.2246806, 0.231949, 0.2613764, 
    0.1388403, 0.2094117, 0.1901027, 0.1495738, 0.146989, 0.221009, 
    0.1993908, 0.1282706, 0.1817324, 0.2339387, 0.2726277, 0.2118192, 
    0.1324553, 0.151918, 0.1146128, 0.1282959, 0.1052936, 0.1978664, 
    0.279315, 0.247666, 0.1982503, 0.2038424,
  0.1706828, 0.1497984, 0.1680786, 0.1752513, 0.1935101, 0.2023994, 
    0.1792529, 0.1385578, 0.1972075, 0.1456667, 0.09783545, 0.07920501, 
    0.06395819, 0.06526186, 0.09938455, 0.1093426, 0.09326816, 0.09838268, 
    0.07721239, 0.07783086, 0.07246864, 0.1081241, 0.1003934, 0.05957946, 
    0.01188786, 0.07409872, 0.159373, 0.1864384, 0.1858487,
  0.0695938, 0.02470567, 0.0135781, 0.0683205, 0.04126729, 0.0352729, 
    0.0826607, 0.06415582, 0.04576315, 0.02861951, 0.02750839, 0.01734858, 
    0.02291241, 0.07456382, 0.1383511, 0.04175532, 0.03437546, 0.04550235, 
    0.08943933, 0.08120526, 0.06726125, 0.0648248, 0.03087409, 0.08645368, 
    0.03987816, 0.04020949, 0.0716356, 0.0573908, 0.06274737,
  0.01686935, 0.006600005, 0.005206696, 0.00992653, 0.01361458, 0.006329053, 
    0.02892753, 0.01106155, 0.008560766, 0.004526999, 0.001076699, 
    3.119409e-05, 0.0001128912, 0.002105004, 0.01917945, 0.008433532, 
    0.007777318, 0.08120228, 0.04804402, 0.01151458, 0.003880847, 
    0.003160649, 0.008154622, 0.007569592, 0.001368398, 0.01440801, 
    0.02975674, 0.00287538, 0.007572799,
  0.009435287, 0.02899729, 0.002267063, 0.002895874, -0.001079794, 
    0.0004778217, 0.0004308239, 0.0005444821, 0.008241249, 0.001577739, 
    0.001153533, 1.371771e-06, 0.000685096, 0.0003950566, 0.001657323, 
    0.0007064746, 0.0007471313, 0.0001359978, 8.027978e-05, 4.056264e-05, 
    4.368107e-05, 0.001705402, 0.009291615, 0.03702465, 0.009385752, 
    0.07026194, 0.0002110771, 0.001506527, 0.002435787,
  0.0129444, 0.001507243, 0.03333521, 0.05426198, 0.001056349, 0.001237841, 
    0.0004146459, 0.000567837, 0.0006904132, 0.001711274, 0.0003912462, 
    0.0003900821, 0.0001801819, 0.000159381, 0.0001976602, 0.0001936861, 
    0.0001177129, 0.0001109973, 0.0001108402, 0.0001957168, 0.001120829, 
    0.004138824, 0.02425764, 0.01152224, 0.01818074, 0.003328026, 
    0.0001424087, 0.0005457322, 0.004122335,
  0.002756159, 0.008461501, 0.01536751, 0.04714412, 0.0007197451, 
    0.0004666301, 0.002023143, 0.0005112838, 0.03966322, 0.09037088, 
    0.0008546307, 0.001243483, 0.0001191793, 0.0004146119, 0.0005339228, 
    0.0003586899, 0.000396228, 0.0002507681, 0.0004251252, 0.0003833045, 
    0.002138414, 0.01698959, 0.02149071, 0.01084836, 0.004131462, 
    0.0002039155, 0.001276705, 0.001134863, 0.0005362692,
  3.754832e-10, 7.237322e-10, 4.989368e-09, 0.0144083, 0.02087096, 
    0.0005710383, -0.001764914, 0.0005318669, 0.001647628, 0.0006188205, 
    0.002202725, 0.0001572416, 0.0003280442, 7.585045e-05, 0.0003203214, 
    0.002925557, 0.001389048, 0.0007466438, 0.001218513, 0.002729423, 
    0.00157423, 0.0003257373, 0.1393635, 0.03554709, 0.0001152559, 
    1.910229e-05, 0.001162504, -3.267681e-06, 6.269609e-09,
  4.986267e-09, -4.838311e-06, 1.021142e-05, 9.66194e-05, 9.96126e-05, 
    0.0008824719, 0.007501468, 0.00115113, 0.02218432, 0.02110713, 
    0.00292663, 0.0008318051, 0.0002323572, 0.0001918272, 0.000372493, 
    0.0005014973, 0.0009679826, 0.002305519, 0.003996457, 0.01196473, 
    0.002396144, 0.05241917, 0.0004261688, -0.001365912, 0.0009842925, 
    7.586682e-05, 0.000452792, 2.368264e-05, 2.206647e-08,
  -1.834128e-05, 0.01237447, 0.00233068, 0.006334816, 0.06215977, 0.02825592, 
    0.008635798, 0.01121418, 0.02314657, 0.05754227, 0.02876091, 0.002898563, 
    0.00449626, 0.004464339, 0.007741408, 0.02984248, 0.01491241, 
    0.003815778, 0.01007917, 0.01385002, 0.07132258, 0.130651, 0.06910994, 
    0.01451687, 0.0093311, 0.002377577, 0.001279506, 0.003716073, 0.0001832674,
  0.009168297, 0.008380586, 0.03446306, 0.2942001, 0.003498746, 0.03083541, 
    0.1061925, 0.002161821, 0.0003310961, 0.04314224, 0.1336956, 0.02017933, 
    0.02391481, 0.01838695, 0.06360137, 0.05128681, 0.09344932, 0.03827647, 
    0.01456014, 0.2648799, 0.07207473, 0.02934657, 0.1564972, 0.1206844, 
    0.03339605, 0.02439331, 0.02453467, 0.019655, 0.0471858,
  0.1242271, 0.2968806, 0.2717316, 0.3045884, 0.2104511, 0.1768987, 
    0.06618927, 0.1650511, 0.159399, 0.141939, 0.1121387, 0.2571747, 
    0.01554833, 0.02709331, 0.0853224, 0.1265815, 0.1093176, 0.06641416, 
    0.04045173, 0.3835755, 0.05941735, 0.06420982, 0.149618, 0.4353599, 
    0.1198511, 0.07453446, 0.05698052, 0.04932791, 0.08121195,
  0.04869505, 0.4127176, 0.3361591, 0.4841756, 0.5368558, 0.3676068, 
    0.4526632, 0.4375543, 0.5139212, 0.5285117, 0.5847479, 0.6218214, 
    0.2915917, 0.2862759, 0.1968865, 0.231612, 0.5183554, 0.1975663, 
    0.2945881, 0.294272, 0.6942753, 0.3183545, 0.2315393, 0.3751965, 
    0.1213105, 0.01421641, 0.05710275, 0.04865097, 0.0543849,
  0.07101393, 0.0515347, 0.3489541, 0.0300264, 0.1418237, 0.2640459, 
    0.4777649, 0.4622568, 0.515626, 0.6322424, 0.7094619, 0.4610062, 
    0.7454165, 0.2948744, 0.3407652, 0.2921231, 0.322072, 0.1456741, 
    0.2797319, 0.2164681, 0.3661087, 0.579343, 0.4847225, 0.5285913, 
    0.3480188, 0.1178346, 0.4897313, 0.0663736, 0.1590601,
  0.4112927, 0.1754772, 0.3517069, 0.3945239, 0.4480289, 0.4782487, 
    0.4213721, 0.4279156, 0.413173, 0.3615327, 0.4568487, 0.4358368, 
    0.4592795, 0.4814524, 0.4260479, 0.418286, 0.4141584, 0.3857674, 0.40616, 
    0.3857582, 0.4416783, 0.29815, 0.4024321, 0.572209, 0.0762053, 0.0198255, 
    0.09300555, 0.1746335, 0.4675114,
  0.0724664, 0.07403128, 0.07559615, 0.07716101, 0.07872589, 0.08029076, 
    0.08185564, 0.06631727, 0.06627509, 0.0662329, 0.06619073, 0.06614855, 
    0.06610636, 0.06606418, 0.0820141, 0.08157755, 0.08114102, 0.08070449, 
    0.08026795, 0.07983141, 0.07939488, 0.07328109, 0.07219493, 0.07110879, 
    0.07002264, 0.06893648, 0.06785032, 0.06676418, 0.07121451,
  0.05374101, 0.03470445, 0.04313329, 0.07593192, 0.03789479, 0.01640716, 
    0.033712, 0.06568468, 0.05630128, 0.05131031, 0.02664379, 0.02062297, 
    0.02581946, 0.0004428828, 0.0521825, 0.09185749, 0.1092377, 0.06058774, 
    0.02675473, 0.03494858, 0.02393295, 0.05583933, 0.1082134, 0.04779716, 
    0.02082738, 0.04859213, 0.03547468, 0.01985042, 0.0192467,
  0.1180319, 0.04878757, 0.06504662, 0.04120249, 0.008899781, 0.1459998, 
    0.07357186, 0.01755421, 0.01307898, 0.01662142, 0.01826113, 0.04127519, 
    0.007768424, 0.1153938, 0.1807854, 0.1215414, 0.1564393, 0.1491205, 
    0.1324575, 0.1669834, 0.1475317, 0.1948921, 0.2212661, 0.211611, 
    0.163078, 0.1895244, 0.1168843, 0.09858508, 0.1091778,
  0.1352407, 0.1484789, 0.1616381, 0.1558759, 0.1943518, 0.2002059, 
    0.2197984, 0.1180421, 0.174861, 0.1617829, 0.1269317, 0.1226769, 
    0.1876405, 0.1649409, 0.1068936, 0.1505872, 0.1998395, 0.2339228, 
    0.1809607, 0.1100266, 0.1202867, 0.09036317, 0.1000776, 0.08319907, 
    0.1617538, 0.2314951, 0.2134318, 0.1716732, 0.1740363,
  0.1452323, 0.1283354, 0.1437639, 0.1399502, 0.1598507, 0.1703137, 
    0.1457448, 0.1105647, 0.1592567, 0.1200539, 0.07605769, 0.06161509, 
    0.04884394, 0.05070851, 0.07461356, 0.08407139, 0.07026585, 0.07042968, 
    0.05442331, 0.05654625, 0.05414843, 0.08365415, 0.07890654, 0.06038857, 
    0.008991154, 0.05963462, 0.1287495, 0.1571011, 0.158265,
  0.05092769, 0.01719355, 0.008922894, 0.05079488, 0.02745297, 0.02569964, 
    0.06098176, 0.04429662, 0.03200191, 0.02243126, 0.01982824, 0.01338942, 
    0.01342016, 0.0541282, 0.1370881, 0.02650217, 0.02290499, 0.03316092, 
    0.06476688, 0.05662708, 0.04527656, 0.04674584, 0.02136448, 0.08620415, 
    0.03243963, 0.02837668, 0.05352814, 0.04250113, 0.04673337,
  0.01127667, 0.005368831, 0.004808124, 0.006578302, 0.008282457, 
    0.004662342, 0.01863915, 0.007698109, 0.007286865, 0.004008672, 
    0.0007587444, 2.012156e-05, 0.007068196, 0.001624485, 0.01222223, 
    0.005130152, 0.005226634, 0.0512685, 0.03126651, 0.006988412, 
    0.002737759, 0.002633812, 0.006786472, 0.006236731, 0.006624863, 
    0.008700056, 0.0166749, 0.00191277, 0.00534787,
  0.007646146, 0.02236615, 0.001039297, 0.002283808, -0.000997026, 
    0.000362008, 0.0003361239, 0.0004570312, 0.006809176, 0.001266665, 
    0.000658677, 1.94953e-06, 0.0005531278, 0.0002787141, 0.001101572, 
    0.000534996, 0.0005691109, 0.0001077399, 6.581791e-05, 3.633379e-05, 
    3.652634e-05, 0.001403739, 0.00740525, 0.03085161, 0.02146246, 0.1463911, 
    0.0001754604, 0.001247462, 0.001963096,
  0.0105922, 0.0006134944, 0.0950999, 0.1458278, 0.0007287647, 0.0008328243, 
    0.0002714025, 0.0003975164, 0.0005608721, 0.001260864, 0.000275032, 
    0.0003052912, 0.000154676, 0.0001219638, 0.0001621196, 0.0001402533, 
    8.574247e-05, 8.069997e-05, 9.164352e-05, 0.0001652632, 0.0009385254, 
    0.003373837, 0.01983827, 0.0802182, 0.0453693, 0.01008691, 0.0001302289, 
    0.0004524282, 0.003360636,
  0.001815771, 0.01361968, 0.01504741, 0.05295727, 0.0004423162, 
    0.0003618172, 0.001396261, 0.0003697316, 0.07420488, 0.1415353, 
    0.0005189807, 0.001015888, 9.467179e-05, 0.0003258122, 0.000410019, 
    0.0002925288, 0.0003164909, 0.00020102, 0.0003466586, 0.0003087253, 
    0.001728073, 0.01318595, 0.01645918, 0.06350949, 0.0432175, 0.0001426577, 
    0.0007581802, 0.0008672399, 0.0004115305,
  3.962579e-10, 7.34778e-10, 4.752717e-09, 0.02271144, 0.01554928, 
    0.0004757438, -0.001213771, 0.0004563229, 0.0009223949, 0.0005219636, 
    0.001510426, 0.0001146995, 0.0001951916, 7.743206e-05, 0.0002660664, 
    0.001653375, 0.0008393885, 0.0004956484, 0.0007881028, 0.001771369, 
    0.0009793375, 0.0001718437, 0.1774268, 0.03300691, 6.956433e-05, 
    1.621114e-05, 0.0009987038, -2.818136e-06, 2.168475e-08,
  5.043109e-09, -3.156171e-06, 7.903089e-06, 9.518083e-05, 7.411707e-05, 
    0.0007616424, 0.008534116, 0.0008309274, 0.02418033, 0.01565736, 
    0.002081895, 0.0006408289, 0.0002019417, 0.0001623138, 0.000315233, 
    0.0003966545, 0.0007029894, 0.001437597, 0.002557107, 0.008144515, 
    0.001899208, 0.04397907, 0.0003615773, -0.001497738, 0.0006624849, 
    6.312491e-05, 0.0003889489, 2.093407e-05, 2.206773e-08,
  -2.031972e-05, 0.01032215, 0.001770844, 0.005806352, 0.05835856, 
    0.02528676, 0.01720681, 0.03595109, 0.04573704, 0.05577793, 0.02273129, 
    0.002313372, 0.00287588, 0.002611046, 0.005234917, 0.01961306, 
    0.009381648, 0.002829052, 0.007055376, 0.01035007, 0.06182091, 0.1197334, 
    0.07363937, 0.01037096, 0.005995658, 0.001835238, 0.001073738, 
    0.003152688, 0.0005254619,
  0.01266974, 0.00685681, 0.03055678, 0.2890388, 0.002788278, 0.0258194, 
    0.1066817, 0.00279365, 0.0002550701, 0.04527283, 0.1417086, 0.01601903, 
    0.02097998, 0.01427917, 0.05400928, 0.04012164, 0.07165416, 0.02952601, 
    0.01055211, 0.2596259, 0.07078246, 0.03272794, 0.1549675, 0.1000464, 
    0.0261244, 0.01695417, 0.01618416, 0.01331461, 0.03923728,
  0.1039308, 0.2936234, 0.2627546, 0.2960447, 0.1915541, 0.1603783, 
    0.06190936, 0.2463085, 0.2692175, 0.1518053, 0.1274555, 0.2897893, 
    0.01340526, 0.02363774, 0.07058586, 0.1074914, 0.09136268, 0.05482646, 
    0.03220914, 0.3929007, 0.06125284, 0.06319314, 0.175141, 0.4377422, 
    0.1176793, 0.06631864, 0.04525603, 0.03753328, 0.06109177,
  0.03945691, 0.5135787, 0.3399109, 0.4635801, 0.5205984, 0.3771578, 
    0.447062, 0.4405097, 0.5089597, 0.5070896, 0.5576035, 0.6000118, 
    0.3516074, 0.3564245, 0.1820877, 0.2194174, 0.5535332, 0.2080815, 
    0.3206457, 0.3725866, 0.658527, 0.3279846, 0.2052102, 0.3765762, 
    0.1188163, 0.01642504, 0.04999758, 0.04060066, 0.04310827,
  0.06058336, 0.04411628, 0.4171079, 0.02569881, 0.1298467, 0.2158926, 
    0.4485125, 0.4716138, 0.5697477, 0.6122737, 0.6926557, 0.5268344, 
    0.6291879, 0.2437807, 0.2996838, 0.2598727, 0.3415389, 0.1370672, 
    0.2618245, 0.1887634, 0.3367308, 0.5243326, 0.4523367, 0.555617, 
    0.3845113, 0.107663, 0.4956807, 0.06364949, 0.1422456,
  0.3957975, 0.1760375, 0.3294809, 0.3394448, 0.3753548, 0.4186321, 
    0.3400738, 0.3346105, 0.335862, 0.2902879, 0.3638584, 0.3305224, 
    0.3431205, 0.3843691, 0.3437188, 0.3263881, 0.3157547, 0.3017714, 
    0.3044128, 0.3043474, 0.3257819, 0.2719927, 0.4169219, 0.6409438, 
    0.07584643, 0.009650025, 0.0918745, 0.2145067, 0.4339011 ;

 average_DT = 730 ;

 average_T1 = 350.5 ;

 average_T2 = 1080.5 ;

 climatology_bounds =
  350.5, 1080.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
