netcdf atmos.1980-1981.aliq.05 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	pfull = 65 ;
	lat = 18 ;
	lon = 29 ;
	bnds = 2 ;
variables:
	float aliq(time, pfull, lat, lon) ;
		aliq:long_name = "Cloud fraction for large-scale liquid clouds" ;
		aliq:units = "dimensionless" ;
		aliq:_FillValue = -999.f ;
		aliq:missing_value = -999.f ;
		aliq:interp_method = "conserve_order2" ;
		aliq:cell_methods = "time: mean within months time: mean over years" ;
		aliq:time_avg_info = "average_T1,average_T2,average_DT" ;
	double average_DT(time) ;
		average_DT:long_name = "Length of average period" ;
		average_DT:units = "days" ;
	double average_T1(time) ;
		average_T1:long_name = "Start time for average period" ;
		average_T1:units = "days since 1979-01-01 00:00:00" ;
	double average_T2(time) ;
		average_T2:long_name = "End time for average period" ;
		average_T2:units = "days since 1979-01-01 00:00:00" ;
	double climatology_bounds(time, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double pfull(pfull) ;
		pfull:standard_name = "air_pressure" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:units = "mb" ;
		pfull:positive = "down" ;
		pfull:axis = "Z" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:climatology = "climatology_bounds" ;
		time:units = "days since 1979-01-01 00:00:00" ;
		time:calendar = "standard" ;
		time:axis = "T" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.4.4 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f9d8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2024.05" ;
		:git_hash = "5d306c05d9fe755cab04eedc8fd3de0d3c8355a0" ;
		:creationtime = "Mon Aug 25 14:09:46 2025" ;
		:hostname = "pp050" ;
		:history = "Mon Aug 25 13:32:18 2025: ncks -d lat,,,10 -d lon,,,10 atmos.1980-1981.aliq.05.nc reduced/atmos.1980-1981.aliq.05.nc\n",
			"Mon Aug 25 14:40:39 2025: cdo -O -s -select,month=5 merged_output.nc monthly_nc_files/all_years.5.nc\n",
			"Mon Aug 25 14:40:11 2025: cdo -O -s -mergetime /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198001-198012.aliq.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/shards/ts/regrid-xy/180_288.conserve_order2/atmos_month/P1M/P1Y/atmos_month.198101-198112.aliq.nc merged_output.nc\n",
			"Mon Aug 25 14:12:17 2025: cdo --history splitname 19800101.atmos_month.nc /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/split/regrid-xy/180_288.conserve_order2/19800101.atmos_month.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_month --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f10d9r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/run2/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field (**please see the field list in this file**) --output_file 19800101.atmos_month.nc" ;
		:CDO = "Climate Data Operators version 2.4.4 (https://mpimet.mpg.de/cdo)" ;
		:comment = "FMS time averaging, version 3.0, precision=double" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 aliq =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.931458e-06, 0, 0, 0.0004217719, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001464731, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -1.000506e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -7.22403e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, -3.795297e-06, -1.562435e-05, 0.0002832587, 0, 
    0.0009912022, 0, 4.627312e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, -1.152206e-05, 0, 0, -1.3172e-10, 0, 0, 0, 0.0006554348, 0, 
    -7.091822e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -2.465902e-06, 0.0009058582, 0, -4.796604e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0001297366, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.392871e-05, 0, 4.888447e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0007294652, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, -1.672548e-05, -6.532519e-05, -5.189622e-05, 
    -1.633792e-05, 0.0004248859, 0, 0.00254446, 0, 0.0004856471, 0, 0, 0, 
    -8.640995e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0001351755, -4.505384e-05, 0, 0, 0.0006141434, 0, 0, 1.060849e-06, 
    0.0006958305, 9.376515e-05, 6.605856e-06, 0, 0, -8.942249e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.515256e-06, -2.011133e-05, 0.001095627, -1.56103e-06, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -3.842625e-06, 0, -1.672076e-05, 0.0023941, 
    -1.294166e-05, -2.113139e-05, 0.0007239438, -1.497403e-05, 0, 
    0.0004383897, 0, 0, 0, 0, 0.0005600438, 0.0006745072, 5.323235e-05, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -6.978162e-05, 0, 0.0005574608, 2.043964e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -1.67956e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.578687e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.003270302, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.0006518459, -1.051628e-05, 0.001452566, 0.0005115222, 
    -0.000162939, -3.087936e-05, 0.001501128, 0, 0.006435539, 0.0001911041, 
    0.001580561, 0, 0, 0.0001802597, 0.0004319295, 0, 0, 0, 0, 0.0001089035, 
    0, 0, 0, 0, 0,
  0, 0.0009749716, -8.548899e-06, 0, 0, 0.003087224, 0.001222309, 0, 
    1.381448e-06, 0.002625988, 0.000593749, 9.908818e-06, 0, 0, 2.390758e-05, 
    -7.522971e-07, 0, 0, 0, 0, 0, 0, 0, 0.0006986505, 0.0001146364, 
    0.002605401, -1.239167e-06, 0, -2.616027e-06,
  0, 0, 0, -1.347393e-05, 0, 0, 0, 0.0001703137, 0, -2.042109e-05, 
    0.004856185, -3.459854e-05, 0.0008178277, 0.00129677, -8.981859e-05, 
    -1.157316e-05, 0.001023011, -1.379753e-05, -4.456248e-05, 3.749007e-05, 
    -2.587019e-06, 0.002853111, 0.001091944, 7.097646e-05, 0, 0, 0, 0, 
    -3.019034e-05,
  0, 0, 0, 0, 0, 0, 0, -0.0001382719, 0, 0.00143389, 0.0002033284, 0, 
    -9.283653e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.315791e-05, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, -8.904625e-06, 0, 0, -2.720448e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -7.834731e-06, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.67826e-05, 0, 0, 0, 0, 
    0, 0, 0.0002534864, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.929174e-05, 0, 0, 0, 
    0.0003010255, 0, 0, 0, 0, 0, -2.011013e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, -4.832841e-05, -4.787767e-06, -5.596027e-06, 0.004261035, 0, 
    0, 0, 0, 0, 0, 0, 0, -1.65371e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -7.685328e-06, -1.089744e-05, 0.0007483457, 0.001808396, -1.682604e-05, 
    0.003364738, 0.001198417, -0.0003427539, 7.006159e-05, 0.002992623, 
    0.0008550304, 0.01444678, 0.000630553, 0.002915886, 3.162509e-05, 
    -1.944466e-05, 0.001516827, 0.002542111, 0, 0, 0, 0, 0.0006075018, 0, 0, 
    0, 0, 0,
  0, 0.001418193, 0.001345851, 0, 0, 0.003935997, 0.0022998, 0, 
    -4.928847e-08, 0.006055068, 0.001534214, 3.949881e-06, 0, 7.600853e-08, 
    0.0009906676, -4.052117e-06, 0, 0, 0, 0, 0, 0, -9.82668e-09, 0.002223721, 
    0.0002576975, 0.006735558, 0.001336975, 0, 1.546308e-06,
  0.0002200004, 0, 0, -4.596807e-05, 0, 0, 0, 0.0003339257, -2.500871e-06, 
    0.0004067128, 0.007235026, -6.343191e-05, 0.002971411, 0.003140795, 
    -8.937294e-05, -0.0001055581, 0.001779027, -1.020555e-05, 0.0002410554, 
    0.000574308, -2.847727e-05, 0.005903941, 0.001781755, 7.809616e-05, 0, 0, 
    0, -1.271654e-06, -4.405013e-05,
  0, 0, 0, 0, 0, 0, 0, 0.0005831743, 0, 0.005583041, 0.0007467261, 
    9.761417e-06, 0.0004197596, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.053587e-05, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, -1.450251e-05, -3.266134e-07, 0.0004000245, 0, 0, 
    1.627542e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001451634, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.92756e-06, 0, 0.0002185175, 
    0, 8.445352e-05, 0, 0, 0, 0, 0.0003620958, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001754618, -3.230659e-05, 
    -2.329369e-05, 0, 0.002765543, 0, 0.0001682408, 0, 0, 0, -8.042512e-06, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, -0.0001232747, -4.866593e-05, -5.167222e-05, 0.006507847, 0, 
    -4.69105e-05, 0, 0, -4.893588e-06, -4.262056e-06, 0, -2.831031e-06, 
    -9.079308e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -8.261809e-05, 4.953992e-05, 0.001847097, 0.003119288, -3.763913e-05, 
    0.006923003, 0.00577636, 0.0008123766, 0.0002625615, 0.00411155, 
    0.001532752, 0.02302158, 0.00228998, 0.003994298, 0.0002778833, 
    0.0005930269, 0.004349252, 0.007521033, 0, 0, 0, 0, 0.001279187, 0, 0, 0, 
    0, 0,
  0, 0.002360849, 0.003959097, -9.388677e-06, 0, 0.007731568, 0.00317703, 0, 
    0.000237174, 0.008047153, 0.005106866, -5.135601e-05, 2.029658e-08, 
    1.350239e-06, 0.003519978, -1.797541e-05, 3.626971e-06, 0, 0, 0, 0, 0, 
    -4.253006e-06, 0.004588048, 0.0005926063, 0.01620585, 0.003046623, 0, 
    -1.424749e-07,
  0.0006386475, 0, 0, -5.682501e-05, 0, -5.637463e-06, 0.0002557493, 
    0.0003712892, 0.0002740616, 0.0005329544, 0.01042856, 0.0004657667, 
    0.004824128, 0.009807611, 0.001011153, -0.0002124122, 0.00265365, 
    0.001030203, 0.001009707, 0.002223142, -6.51539e-05, 0.01230887, 
    0.003260375, 0.001497572, 0, 0, 0, -8.72786e-06, -9.220134e-05,
  0, 0, 0, 0, 0, 0, 0, 0.0008828237, 7.486448e-05, 0.01462178, 0.001205788, 
    9.00949e-06, 0.002058711, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001584367, 0, 0, 
    0, 0, 0, 0,
  0, 0, -1.266891e-06, 0, 0, 0, 0, -2.341668e-05, 0.0006017851, 0.001221007, 
    0.0001355232, -8.917156e-06, 8.200636e-05, 0, 0, -2.393843e-06, 0, 0, 0, 
    0, 0, 0, 0, 0.002097081, 0.0001223958, 0.0002614789, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002884301, 0.0001011387, 0.0001798022, 
    0.001297359, 0, 0, 0, 0, 0, 0, 0, 8.228622e-05, 0.0008094377, 0, 
    -1.305308e-06, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.696389e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.105186e-06, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, -5.507155e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.377338e-05, 0, 0, 0, 0, 0, -4.960617e-06, 0, 0, 0,
  0, 0, 0, -9.870622e-07, -6.814016e-06, 0.000139517, -2.690606e-05, 0, 0, 0, 
    0, 0, 0, 0, -4.427516e-06, 0.0003214221, -1.527183e-05, 0.00142323, 
    0.0006903075, 0.002547357, 0.0001590827, 0.0002925516, 0, 0, 0.001218603, 
    -2.908844e-10, 0, 0.0001860205, 0,
  0, 0, 0, 0, 0, 2.933863e-05, 0, 0, 6.396435e-05, -3.242874e-06, 0, 0, 0, 0, 
    0.005643395, 0.001606559, 0.0002311201, -3.040755e-05, 0.005201221, 
    -2.859942e-06, 0.001738496, 0, 0, 0, -8.057094e-06, 0.0001452275, 0, 0, 0,
  0, 0, 0, 0, 0, 0.0008292352, 0.0005263247, -0.0001605758, 0.01075668, 0, 
    0.0005272753, 0, -6.926212e-08, 0.0001236189, 0.0002114917, 0, 
    -4.900622e-05, 5.80966e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3.690157e-06,
  0, 0.0004624509, 0.0006487574, 0.003004132, 0.005229983, -3.576794e-05, 
    0.01124566, 0.01794947, 0.003856898, 0.001495263, 0.006733372, 
    0.001877184, 0.03238798, 0.004513183, 0.006097125, 0.0003250385, 
    0.002533772, 0.007271932, 0.01023554, 0, 0, 0, 0, 0.003727494, 0, 0, 0, 
    0, 0,
  0, 0.004163113, 0.006697887, -3.89265e-05, -7.508174e-06, 0.0203313, 
    0.005071045, -3.531083e-06, 0.0004917769, 0.01177531, 0.00967791, 
    0.000800237, -4.021126e-05, 1.876785e-05, 0.008271453, -2.450251e-05, 
    0.001742943, 0, -1.977378e-05, -3.229898e-06, 0, 0, -3.93028e-05, 
    0.008423574, 0.003429514, 0.02165291, 0.003836782, -1.056071e-05, 
    2.823322e-06,
  0.001610722, 0, -6.207634e-07, -4.400915e-05, 0, -7.079389e-06, 
    0.001090333, 0.001322135, 0.0009001691, 0.003441112, 0.01713064, 
    0.001269444, 0.01031006, 0.01788332, 0.007929162, 0.002079983, 
    0.004258029, 0.005705659, 0.004978967, 0.006749169, -0.0001536718, 
    0.02786263, 0.006002946, 0.002370498, 1.509126e-06, -7.767677e-07, 
    8.303438e-05, -6.447262e-06, 7.599997e-05,
  0, 0, 0, 0, 0, 0, 0, 0.00320539, 0.0006983045, 0.02989193, 0.004345196, 
    3.10132e-05, 0.004465709, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0002523029, 
    -1.061371e-05, 0, 0, 0, 0, 0,
  0, 0, 0.0005889809, -1.551584e-07, 0, 0, 0, -6.127553e-05, 0.001739229, 
    0.003170017, 0.003561696, 0.002297898, 0.001325859, 0, 0, 0.0003686511, 
    0, 0, 0, 0, 0, 0, 0, 0.003443677, 0.002582382, 0.003095291, 0, 0, 0,
  0, 0, 0, 0, 0.000211446, 6.013811e-05, 0, 0, 0, -1.205991e-05, 0.001232142, 
    0.0004588784, 0.001355965, 0.004506717, 0, 0, 0, 0, 0, 0, 0, 
    0.0007147809, 0.004571886, 0.002031224, -9.773903e-06, 0.001097385, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.317971e-05, 0.0004867511, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0009870816, 0, 0, 0, -4.100635e-08, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0.0007756878, 0, -3.648337e-06, -1.275005e-05, -7.869753e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001984724, 0.0009291113, 0.00024674, 
    0.0004952084, 0, 0, -3.367645e-05, 0, 0, 0,
  -2.532302e-05, 0, 0, 0.0001167051, 0.0004118886, 0.0003509431, 
    -4.406045e-05, 0, 0, 0, 0, 0, 0, 0, 8.300721e-05, 0.0009994671, 
    0.002874453, 0.004111587, 0.002756568, 0.009172041, 0.003454119, 
    0.00192821, 0.0003719774, 0, 0.008258888, -1.884708e-05, 8.470852e-05, 
    0.002536427, 0.002283558,
  0, 0, 0, 7.545619e-05, -1.364022e-05, 0.0004475828, -1.293669e-05, 0, 
    0.001092252, 7.823759e-05, 0, -3.537763e-09, 0, 0.002947352, 0.01111683, 
    0.007046032, 0.001183839, 0.002324201, 0.009756302, -2.521927e-05, 
    0.003476018, 0, 0, 0, -3.2777e-05, 0.002947938, -1.174435e-05, 
    -4.708702e-08, 0,
  0, 0, 0, 0.0003392454, 0.0001004524, 0.002774376, 0.003188243, 
    -0.0003574878, 0.01753849, 0, 0.002048902, -1.722601e-08, -4.341906e-06, 
    0.001135674, 0.0006681791, 0, 0.0003139534, 0.000186363, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, -3.922547e-06,
  0, 0.0009479094, 0.002766274, 0.003916116, 0.009213631, -2.286122e-05, 
    0.0192393, 0.03262218, 0.009430562, 0.005929054, 0.01595593, 0.003368223, 
    0.05071411, 0.01173052, 0.01138955, 0.001719212, 0.003473327, 0.01044587, 
    0.01523348, -2.171265e-05, 0, 0, 0, 0.007115236, -3.03508e-05, 0, 
    -8.127403e-07, -1.085819e-07, 0,
  0.0004822912, 0.0102293, 0.009438099, 0.0005317004, -5.809327e-05, 
    0.03179464, 0.009499637, 3.539005e-07, 0.001761037, 0.01813821, 
    0.02268226, 0.004477268, 0.0002410842, 0.0002342579, 0.0274243, 
    -3.803485e-05, 0.003872406, -1.155194e-05, -0.0001049776, -3.45911e-05, 
    0, -1.613064e-05, 0.0002042639, 0.01954544, 0.007235221, 0.02984523, 
    0.008950971, 0.0001318791, 0.002878682,
  0.002657374, -3.034713e-05, 0.0002194347, -0.0001646279, 4.54003e-05, 
    -1.577155e-05, 0.002884612, 0.005737952, 0.004147401, 0.01210816, 
    0.02999531, 0.003725366, 0.02268514, 0.02839344, 0.03036369, 0.01054854, 
    0.007653302, 0.01066164, 0.01181801, 0.01361805, 0.000230382, 0.05109303, 
    0.02225078, 0.006036574, 0.000334342, -4.733394e-05, 0.0005006853, 
    0.0003145549, 0.0001581689,
  0, 0, 0, 0, 0, 0, 0, 0.009532969, 0.005058317, 0.04888959, 0.00582332, 
    0.001035479, 0.01089428, -5.084943e-06, 0, -1.439893e-05, 5.665509e-05, 
    7.666832e-05, -4.850528e-05, -3.337639e-06, 0, 0.0001158398, 0.000427134, 
    5.473106e-05, 0, 0, 0, 0, 0,
  0, -1.66396e-05, 0.001497456, 3.345532e-05, -1.208187e-05, 0, 0, 
    -0.0001045613, 0.003768049, 0.008647558, 0.009692214, 0.0140473, 
    0.01022658, 6.630804e-06, 0, 0.002242771, 0, 0, 0, 0, 0, -4.643384e-06, 
    6.935582e-05, 0.007834665, 0.006652053, 0.004537304, 0, 0, 0,
  0, 0, 0, 0, 0.001786981, 0.001967748, 0.0004459114, 0, 0, 2.7454e-05, 
    0.004019842, 0.004143251, 0.006184311, 0.009328702, 1.290384e-07, 
    0.000310222, -9.590163e-06, -6.724109e-06, 0, 0, 0, 0.008032285, 
    0.01041007, 0.003278008, 0.0005794803, 0.002655575, 0, 0, 0,
  0, 0, 0, -2.752565e-05, 0, -7.882581e-06, 0, -1.8771e-06, 0, 0, 
    3.742468e-05, 0.002002493, -5.026823e-05, 0, -3.859574e-07, 0, 0, 0, 0, 
    0, 0, 0.00157244, -4.503684e-05, 0, 0, -6.216187e-05, 0, 0, 0,
  0, 2.575562e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, -5.257683e-06, 0, 4.585094e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -1.764971e-05, 0, 0, 0, 0, 0,
  0.0003960162, -9.414861e-07, 4.14672e-05, 0.0003210897, 0.002930389, 0, 
    -1.215352e-05, 0.0002289963, -2.359817e-05, 3.008866e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 9.268535e-05, 0.003577892, 0.002408821, 0.002026846, 
    0.001160445, 0, 0, -9.182678e-05, 0.0007013725, 3.743633e-05, 0.0006143294,
  0.0009894897, 0, -3.759267e-06, 0.002032161, 0.003909652, 0.002203049, 
    0.001430778, 0.0003739042, 5.191189e-06, 0, 0, 0, 0, -6.261067e-06, 
    0.0007732882, 0.004411926, 0.01131372, 0.006917406, 0.01192913, 
    0.01672057, 0.01488594, 0.002698166, 0.003066474, -1.119021e-05, 
    0.0123454, -2.124641e-05, 0.001498542, 0.004439256, 0.004958468,
  0, 0, 0, 0.001827703, 0.002009425, 0.004283194, 0.0001027755, 0, 
    0.00469079, 0.001638266, -3.90299e-10, 0.0001473914, -9.608672e-06, 
    0.007814287, 0.02821572, 0.01896144, 0.007846607, 0.01458183, 0.02719152, 
    0.0008785454, 0.005442978, -3.699619e-05, 0, 0, -8.951152e-05, 0.0113244, 
    2.968739e-05, -6.07097e-05, 8.458977e-05,
  5.012976e-10, 0, 0, 0.005416007, 0.001057501, 0.005758014, 0.01335213, 
    -9.997138e-05, 0.02452498, 2.095786e-05, 0.003589678, -7.490272e-06, 
    -1.656091e-05, 0.004947674, 0.005525218, 0.001500996, 0.005760043, 
    0.004675243, 6.543159e-05, -1.565931e-07, -1.96325e-06, 0, 0, 0, 0, 
    -2.255907e-08, 2.364794e-05, 0, -1.027357e-05,
  0, 0.002634413, 0.003966549, 0.004145352, 0.01559956, 0.0004806066, 
    0.03398456, 0.04891604, 0.03260555, 0.02102558, 0.03140022, 0.009821318, 
    0.06446159, 0.03681591, 0.01819405, 0.01016074, 0.007129788, 0.01279492, 
    0.01982703, -4.256075e-05, 0, 0, 3.194674e-11, 0.0134421, 0.002157792, 
    -3.695423e-07, 0.0001048171, 0.0001904481, 0,
  0.004382317, 0.02606909, 0.02156611, 0.003772516, 0.0003296061, 0.06060515, 
    0.01815601, 0.0004542809, 0.0236972, 0.04471096, 0.04369313, 0.01612407, 
    0.006083823, 0.009553416, 0.04605227, 0.003202534, 0.006433118, 
    1.924005e-05, 0.0006677774, -7.406105e-05, 3.838469e-08, -4.36044e-05, 
    0.003997124, 0.06530188, 0.01660183, 0.04055624, 0.01902887, 0.005252049, 
    0.00736545,
  0.0111771, -7.361638e-05, 0.001933482, 0.002320808, 4.357264e-05, 
    0.0002788665, 0.01245176, 0.02415342, 0.01632394, 0.03646146, 0.05741679, 
    0.02890933, 0.07602035, 0.06335384, 0.05894679, 0.03097776, 0.01049638, 
    0.02047131, 0.0213944, 0.02892594, 0.00752838, 0.08518626, 0.06623567, 
    0.02530545, 0.001405773, 0.000235202, 0.0004485531, 0.0009156307, 
    0.007520046,
  -4.817646e-10, -3.716874e-07, 0, -1.04757e-06, 0, 0, 0, 0.02133761, 
    0.02766275, 0.0738842, 0.008208273, 0.003645631, 0.0269907, 
    -1.384247e-05, 7.281025e-05, 0.001343456, 7.283443e-07, 0.002581616, 
    0.0005686281, 0.0004926994, 1.055893e-07, 0.0006720031, 0.002459628, 
    0.0008829512, 0.0001132579, 1.512121e-05, 5.227636e-08, 0, 0.0001959493,
  0, -4.314432e-05, 0.002708255, 0.0007763099, 0.0002574047, 0, 0, 
    8.339204e-05, 0.01091461, 0.02226798, 0.02040898, 0.03109236, 0.02740478, 
    0.000487219, -8.479987e-06, 0.004351371, -8.822726e-05, -9.290664e-06, 0, 
    0, 0, 0.000615406, 0.0002797791, 0.01564377, 0.01665263, 0.004936429, 
    0.000550781, 0, 0,
  0, -1.128937e-07, 0.0006834548, -8.479584e-06, 0.006077639, 0.004256128, 
    0.003730318, 0.000260305, -9.796815e-06, 0.00117345, 0.009786545, 
    0.01357523, 0.0265069, 0.02170976, 0.00129237, 0.002065827, 0.000291691, 
    0.001197492, 0, 8.567058e-06, -1.018233e-05, 0.01546188, 0.02026878, 
    0.008318071, 0.00794838, 0.005568815, 4.353031e-06, 0.0004476227, 0,
  0, 0, -2.054751e-06, 0.0004001279, -6.73257e-06, -5.701203e-05, 0, 
    -3.769499e-05, 0, 0, 0.0003356008, 0.003489876, 0.002461804, 0.001497818, 
    0.0005827273, -1.696216e-05, 9.758508e-05, 0, 0, 0, -2.108404e-05, 
    0.003603063, 0.001683513, -3.913312e-05, 0, 0.0004056987, -9.827605e-06, 
    0, 3.31341e-05,
  -6.260596e-05, 3.018613e-05, 0.0009019166, 0, 0.003254998, -1.058905e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2.432631e-06, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000851453, 
    0, -3.721102e-06, 0, 0, 0, 0, 0,
  0, -3.826501e-06, 0, 6.540021e-05, 0, 0.0007164631, 0.0006150104, 
    9.523023e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000615862, 
    0, 0, 0, 0, 0,
  0.001964078, 0.0009422193, 0.001742256, 0.001199956, 0.01173552, 
    0.0001280295, -5.423606e-05, 0.0009073021, -6.677469e-05, 0.0002839538, 
    0, 0.001379252, 0, 0.0001033693, 0, 0.0009538566, 0, 3.425548e-05, 
    0.001548276, 0.004078331, 0.006634839, 0.004623994, 0.002548607, 
    -5.390757e-06, 0, 7.966592e-07, 0.004875324, 0.001147779, 0.004717439,
  0.01168442, 0.001168698, 0.0002143955, 0.00560889, 0.01340679, 0.006786221, 
    0.006269074, 0.001607523, 0.002286077, 0.0002759011, -8.76433e-06, 0, 
    -2.727133e-06, 0.0008563575, 0.002513079, 0.02342721, 0.01975447, 
    0.01928565, 0.02817741, 0.0524648, 0.02870387, 0.0123057, 0.008673381, 
    0.0009361359, 0.01799763, 0.002451298, 0.003868079, 0.01523513, 
    0.009555856,
  3.02773e-06, -2.436597e-06, 0, 0.008592485, 0.01315417, 0.01217197, 
    0.001004369, 0.0004357525, 0.02088728, 0.01291521, 0.002030458, 
    0.0008461868, -8.245556e-05, 0.01619563, 0.05266272, 0.05128671, 
    0.02995235, 0.04716518, 0.05651502, 0.009207361, 0.02192744, 0.004687204, 
    0.002447906, 0.0005891083, -0.0001759655, 0.02156194, 0.002052154, 
    0.001334454, 0.0003083366,
  2.46411e-05, -2.012207e-06, 0, 0.01480783, 0.006237368, 0.007370987, 
    0.0215311, 0.003144844, 0.02846515, 0.01637958, 0.004669885, 
    8.687971e-05, 0.003141525, 0.0140998, 0.0327247, 0.0112138, 0.01282181, 
    0.0165459, 0.001429455, 0.0007482986, -2.540846e-05, 0.0003720771, 
    -1.036928e-06, 4.132264e-06, 0.0002432289, -9.979649e-06, 0.0008616226, 
    0.000603169, 9.356641e-05,
  -1.023523e-05, 0.0176381, 0.006287547, 0.004848538, 0.04029765, 0.03334127, 
    0.05977606, 0.09149531, 0.1284881, 0.1158388, 0.08018632, 0.04614487, 
    0.1071867, 0.1963012, 0.08785263, 0.06431323, 0.01494213, 0.01651463, 
    0.02502227, 0.0003463529, 2.331296e-07, -4.035502e-08, -1.201646e-06, 
    0.02483754, 0.02093459, 0.0001381549, 6.350756e-05, 0.0005582244, 
    1.755859e-06,
  0.05811811, 0.05787885, 0.08470906, 0.00798232, 0.005427241, 0.1183341, 
    0.09727756, 0.07583601, 0.1805751, 0.1699767, 0.1629425, 0.09436248, 
    0.09842747, 0.05002961, 0.128001, 0.06597102, 0.02749452, 0.01279567, 
    0.004768308, 0.007355877, -3.919394e-05, 0.002561842, 0.03138319, 
    0.2048112, 0.1050447, 0.08236351, 0.06440189, 0.03388169, 0.025126,
  0.06605768, 0.01326944, 0.005364755, 0.002578902, -1.705317e-05, 0.0215888, 
    0.1174791, 0.2062919, 0.2067982, 0.1746719, 0.142283, 0.1512951, 
    0.2734661, 0.2091446, 0.1975717, 0.1769679, 0.03680296, 0.03887586, 
    0.03495193, 0.05830466, 0.04288733, 0.1479053, 0.1583551, 0.1585017, 
    0.01117954, 0.02179492, 0.0007919116, 0.02886228, 0.05120285,
  1.617296e-05, -1.482798e-05, -6.79013e-08, 0.0006314865, -2.577514e-05, 
    -4.997965e-06, 2.566582e-05, 0.03715745, 0.1272144, 0.1896755, 
    0.04253804, 0.04664381, 0.1233769, 0.002235826, 0.003667179, 0.00716948, 
    0.002102934, 0.009269066, 0.01303804, 0.004989831, 0.0006823697, 
    0.002732964, 0.005976755, 0.0370176, 0.001116146, 0.002367076, 
    0.003167692, 2.356947e-06, 2.499672e-05,
  -2.110375e-09, 0.001824551, 0.00334496, 0.003849721, 0.0001457856, 
    1.73625e-05, 5.814938e-05, 0.0002046456, 0.02701908, 0.05823918, 
    0.0693711, 0.0675756, 0.07234914, 0.007542071, 1.117337e-05, 0.007080278, 
    0.002628946, -4.201082e-05, 2.153913e-07, 0, 0, 0.002815647, 0.002722228, 
    0.02932599, 0.02446185, 0.005275617, 0.003866661, -1.124934e-06, 
    -8.838962e-11,
  0.0002031231, 0.001722552, 0.002319872, 0.0003670377, 0.01196793, 
    0.007846713, 0.005906883, 0.0007733342, -1.046899e-05, 0.00377841, 
    0.01427661, 0.02932192, 0.05747892, 0.04271168, 0.009609488, 0.01042777, 
    0.0017171, 0.004462, 0, 0.0007010059, 3.811334e-05, 0.02881174, 
    0.04071614, 0.02069575, 0.02826286, 0.0142871, 0.001882426, 0.001396672, 0,
  0.003192171, 0.0008181183, 0.0001256204, 0.000933414, 0.0003624817, 
    0.0003652859, 0.000134225, -4.642938e-05, 0, -5.991858e-06, 0.001756069, 
    0.00664061, 0.005452281, 0.002506973, 0.006316662, 0.001841267, 
    0.0001476428, 0.0004097113, 0, 0, -9.32748e-05, 0.004873151, 0.004847817, 
    0.0003716619, 0.001655397, 0.003847223, 0.00442408, 0.001308806, 
    0.002794062,
  4.895186e-05, 5.986193e-05, 0.001897249, 1.982741e-05, 0.006207857, 
    -2.073521e-05, 8.921781e-05, -1.318452e-05, -8.989588e-06, 0, 0, 0, 0, 0, 
    0, 0, 0, -3.209202e-05, 0, 0, -3.143456e-05, -2.054828e-05, 0, 
    0.001624582, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.1334e-06, 0.0001690591, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002686299, 
    -5.618872e-06, 7.031783e-05, 9.428334e-05, 0, 0, 0, 0,
  -2.15186e-06, -2.93982e-05, -2.704203e-06, 0.001614009, 0.0002198569, 
    0.001093762, 0.002022254, 2.592289e-05, -7.866701e-06, 0, 0, 
    -1.933912e-06, 0, 0, 3.912799e-06, 0, 0, 0, 0.0001751063, 8.650933e-06, 
    0.0001073958, 9.85732e-05, 0.0005038619, 0.001888136, -8.064687e-05, 
    0.0001528188, 0, 0, -1.435328e-05,
  0.01183025, 0.00414825, 0.003269948, 0.00806048, 0.0225221, 0.002269404, 
    0.003070049, 0.002666739, 0.0007210669, 0.001357687, 0, 0.003195382, 
    -2.21173e-06, 0.001375405, 7.115286e-05, 0.0009530399, 0.001701164, 
    0.001098887, 0.004747258, 0.009390553, 0.01373856, 0.01113853, 
    0.01157141, 0.001954725, 0.00433508, 0.002262429, 0.01143697, 
    0.008041618, 0.01031019,
  0.0202383, 0.004108567, 0.0009765058, 0.01269607, 0.02395172, 0.01335999, 
    0.01338424, 0.00521988, 0.005980561, 0.0009912425, 0.003526817, 
    -5.142336e-05, 0.0005358262, 0.003933838, 0.01115803, 0.04363623, 
    0.03499422, 0.04235392, 0.05465516, 0.09742413, 0.0579119, 0.03616167, 
    0.01380179, 0.007196809, 0.02270782, 0.009197511, 0.008086927, 
    0.03079301, 0.01675574,
  0.0009411698, 0.0005884903, -9.108546e-06, 0.02069898, 0.03208735, 
    0.02427442, 0.007256697, 0.005054265, 0.03058759, 0.0214558, 0.008887588, 
    0.0106565, 0.0008385707, 0.0273843, 0.09464209, 0.1446086, 0.09206061, 
    0.09944437, 0.1232825, 0.0702849, 0.05056475, 0.03525247, 0.01114319, 
    0.008777598, 0.0008092515, 0.04385082, 0.01592184, 0.005724174, 
    0.003505923,
  0.003029862, 0.0002160132, 0.0001249268, 0.05064426, 0.05768396, 
    0.04871878, 0.05626502, 0.02579885, 0.03754277, 0.04502567, 0.01394858, 
    0.0007433483, 0.002626693, 0.04111702, 0.1041197, 0.05058818, 0.05378107, 
    0.1053517, 0.1240586, 0.02090189, 0.002898311, 0.003336355, 0.0001815005, 
    0.002922755, 0.01685697, 0.002671427, 0.01916809, 0.01867976, 0.002017497,
  0.0008445301, 0.04606196, 0.01940602, 0.007039751, 0.06977004, 0.06625128, 
    0.08371919, 0.0967901, 0.1000297, 0.08239633, 0.08393638, 0.03021263, 
    0.09744571, 0.1567904, 0.07780939, 0.07094651, 0.02812071, 0.03010242, 
    0.0405071, 0.00144006, 1.960844e-06, 1.475512e-05, 0.005884382, 
    0.1783972, 0.1127812, 0.05237522, 0.001750162, 0.001077135, 0.0002722572,
  0.1341842, 0.3091594, 0.3211286, 0.03052654, 0.02916066, 0.1422819, 
    0.09438218, 0.08354311, 0.3173068, 0.3482069, 0.1350092, 0.07329914, 
    0.06797423, 0.03933283, 0.1177368, 0.04331613, 0.02971365, 0.01359411, 
    0.00323323, 0.007525878, 0.001869595, 0.00181072, 0.1055849, 0.3620977, 
    0.1606051, 0.1065236, 0.0799937, 0.05496503, 0.04201382,
  0.1745875, 0.08147734, 0.05759223, 0.004558799, 0.001562403, 0.03009169, 
    0.09579609, 0.15806, 0.1635042, 0.1339763, 0.1180185, 0.1081891, 
    0.2175025, 0.1855874, 0.2049972, 0.235685, 0.120797, 0.09164768, 
    0.09729324, 0.1023507, 0.08044037, 0.180507, 0.2712829, 0.3015443, 
    0.02725486, 0.04637188, 0.02335136, 0.02299177, 0.2797704,
  0.04180923, 0.004622896, 1.9617e-06, 0.03568023, 0.02629406, 1.506079e-06, 
    0.009401107, 0.0302083, 0.2073298, 0.170619, 0.09177762, 0.05791997, 
    0.1362292, 0.05448698, 0.02351342, 0.07399677, 0.05995495, 0.1055008, 
    0.1395094, 0.09104348, 0.04041518, 0.007641326, 0.03518074, 0.1947708, 
    0.1796941, 0.08549183, 0.02942289, 0.02345563, 0.06222314,
  0.002658651, 0.005517377, 0.006622932, 0.01169336, 0.006363641, 
    0.0007589583, 0.002226989, 0.001216307, 0.0647386, 0.2240138, 0.2009273, 
    0.2089192, 0.1658574, 0.06987638, 0.02981498, 0.01944641, 0.01488833, 
    0.001539044, 0.003250165, -8.585702e-06, 0.001322519, 0.01170999, 
    0.01975693, 0.06018054, 0.08434532, 0.01783325, 0.01693359, 0.003955805, 
    -6.850401e-05,
  0.001404494, 0.004277295, 0.006002094, 0.003471501, 0.02266888, 0.01427502, 
    0.01169082, 0.00283891, 0.000382505, 0.009935601, 0.03466776, 0.06289283, 
    0.150727, 0.1505167, 0.06787477, 0.03596479, 0.0153604, 0.01599516, 
    0.001995286, 0.001770929, 0.0001740456, 0.04215157, 0.06203474, 
    0.04098748, 0.05244109, 0.03232792, 0.005114105, 0.003243855, 0.0002871123,
  0.01040563, 0.001422447, 0.001034656, 0.001449507, 0.00153505, 0.004745448, 
    0.003262052, 2.25568e-05, 0, -4.104155e-05, 0.005777903, 0.01377976, 
    0.01497164, 0.01718523, 0.0203166, 0.004676496, 0.002638942, 0.01112948, 
    -8.039822e-08, 0, 0.0008017922, 0.01007358, 0.0101705, 0.001807757, 
    0.005510918, 0.00852439, 0.007344872, 0.001409184, 0.008444987,
  0.001019191, 0.0005418799, 0.002394808, 0.003549975, 0.01251254, 
    0.001585297, 0.001180208, -2.295133e-05, -3.856835e-05, 0, 4.981212e-07, 
    -4.95821e-06, 0.0002404821, -1.206861e-06, -4.587008e-05, 1.326188e-06, 
    -7.57385e-10, -3.20927e-05, 0, 0, 0.000337588, 0.00160053, -1.576638e-06, 
    0.003603541, -8.115183e-06, -2.884033e-05, 0, 0, -8.672306e-06,
  0, 0, 0, 1.954716e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0004028437, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.393453e-06, -5.136636e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    -2.1334e-06, 0.0001690591, -2.257666e-05, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -9.975085e-06, 
    -5.29112e-06, 0.003424906, 0.004589954, 4.781629e-05, 0.0006171091, 0, 0, 
    0, 0,
  0.0006765334, 0.002097253, 0.0006220159, 0.006575354, 0.0006460593, 
    0.003834603, 0.004466647, 0.0003987826, 0.0001299485, -2.946355e-05, 
    0.001068015, 5.415304e-05, 2.412722e-06, -2.804049e-06, 0.0005471886, 
    -4.140163e-06, 0, 0, 0.0008972179, 0.001012345, 0.003922225, 0.00707191, 
    0.004820946, 0.00750128, 0.003103409, 0.001212548, -0.0001696185, 
    -3.275751e-08, -6.217464e-05,
  0.03218257, 0.01312917, 0.006384327, 0.01775395, 0.03382286, 0.01118389, 
    0.009360569, 0.009493073, 0.00803232, 0.006452621, 0.002309944, 
    0.006582222, 0.001768287, 0.002896749, 0.002960386, 0.00118563, 
    0.006195836, 0.006839838, 0.008185854, 0.02159569, 0.02858977, 
    0.02579788, 0.03862736, 0.01947125, 0.01982798, 0.007872472, 0.0205582, 
    0.01746441, 0.02341088,
  0.03356952, 0.009763952, 0.00840284, 0.02281011, 0.05640676, 0.03433834, 
    0.02862389, 0.01577076, 0.01863511, 0.01001904, 0.01700288, 0.00282293, 
    0.00379179, 0.01257223, 0.03685857, 0.06790301, 0.05160438, 0.06684314, 
    0.09414053, 0.178324, 0.136861, 0.09033558, 0.03666376, 0.0319235, 
    0.03842106, 0.03684471, 0.04400265, 0.06702486, 0.04164068,
  0.03336008, 0.01118509, 0.006864028, 0.03285127, 0.0857139, 0.0582207, 
    0.04115191, 0.02125619, 0.07402429, 0.07140694, 0.04962639, 0.03108983, 
    0.00483699, 0.05051637, 0.1301737, 0.2054919, 0.1607575, 0.1647791, 
    0.2475288, 0.1990014, 0.1199269, 0.07229413, 0.03114512, 0.03683032, 
    0.02246653, 0.09031247, 0.06947767, 0.0439119, 0.02633333,
  0.0002463651, 0.003638173, 0.0004914881, 0.06306381, 0.06032694, 
    0.04481776, 0.04908039, 0.02775048, 0.04060014, 0.04768519, 0.01370011, 
    0.0005058197, 0.004493975, 0.04590176, 0.1005111, 0.04476448, 0.0552638, 
    0.1023598, 0.07262778, 0.01249132, 0.001647928, 0.001565276, 
    3.603275e-05, 0.0005982987, 0.007180006, 0.005030564, 0.01003761, 
    0.01683371, -0.0001044787,
  0.00057021, 0.04294917, 0.01463495, 0.007924105, 0.05468028, 0.03572847, 
    0.06930591, 0.07299693, 0.0815459, 0.06314945, 0.07283963, 0.01943407, 
    0.08302896, 0.1236719, 0.06063305, 0.05391848, 0.02014993, 0.0263281, 
    0.03387934, -2.1239e-05, 1.797009e-06, 2.538248e-06, 0.01147986, 
    0.1179935, 0.06747674, 0.03040287, 0.000930063, 6.203815e-05, 2.226964e-05,
  0.09955934, 0.2806593, 0.2421535, 0.02033596, 0.01629018, 0.1089133, 
    0.07677004, 0.03742041, 0.2323178, 0.276117, 0.1176445, 0.0588792, 
    0.04499932, 0.03208981, 0.09712392, 0.02990135, 0.02527518, 0.02350719, 
    0.009237677, 0.004843215, 0.0007737276, 6.356544e-05, 0.06340831, 
    0.3196102, 0.1139515, 0.08506133, 0.06448511, 0.03564873, 0.02310148,
  0.1468823, 0.06100188, 0.05494639, 0.07044331, 0.001177677, 0.01708472, 
    0.06477712, 0.1237943, 0.1374921, 0.1079888, 0.1077219, 0.0789957, 
    0.1773156, 0.1577719, 0.1538978, 0.1861505, 0.08622912, 0.07909267, 
    0.05407715, 0.08230051, 0.05895973, 0.1507248, 0.2278699, 0.2549978, 
    0.01943243, 0.03115397, 0.01361147, 0.01804966, 0.2351726,
  0.04723215, 0.01231259, 0.01543286, 0.034008, 0.05096134, 0.01952024, 
    0.01273489, 0.02262891, 0.1485017, 0.1466295, 0.08333052, 0.0403427, 
    0.103721, 0.03964629, 0.009542055, 0.06979895, 0.06891631, 0.1020608, 
    0.1575246, 0.06278956, 0.02581846, 0.01124732, 0.03204018, 0.1605981, 
    0.1783949, 0.08157295, 0.03972489, 0.04292145, 0.06654246,
  0.03349723, 0.05927019, 0.03007278, 0.04263953, 0.05993164, 0.02663273, 
    0.03257477, 0.002976368, 0.1102267, 0.1997381, 0.1903038, 0.2154922, 
    0.1741601, 0.08610193, 0.04286034, 0.1006039, 0.1083341, 0.05914468, 
    0.04709779, 0.02342501, 0.0113675, 0.1000913, 0.06902924, 0.1277423, 
    0.1393257, 0.1306426, 0.1017457, 0.05208836, 0.02245202,
  0.01110637, 0.00887601, 0.0152226, 0.01092413, 0.04436275, 0.06871562, 
    0.018657, 0.03714303, 0.0248754, 0.04007938, 0.07191674, 0.106108, 
    0.2337644, 0.2540165, 0.1657996, 0.1315945, 0.1105942, 0.09312019, 
    0.02441782, 0.007855231, 0.0007794785, 0.05776951, 0.09611725, 
    0.09524546, 0.1349119, 0.08827896, 0.05136937, 0.02535916, 0.0123962,
  0.02035536, 0.003656063, 0.004595268, 0.006148776, 0.00645261, 0.01495025, 
    0.01066782, 0.001750535, 2.836925e-05, 0.0006636821, 0.01824046, 
    0.02446193, 0.05003853, 0.06110447, 0.08807674, 0.05786606, 0.03261521, 
    0.03427329, 0.006786749, -4.782041e-10, 0.002297967, 0.01997656, 
    0.02020389, 0.005651198, 0.01509974, 0.02539193, 0.03599836, 0.01426609, 
    0.02002593,
  0.004853519, 0.0034707, 0.006233886, 0.008783766, 0.01698051, 0.007908915, 
    0.002031218, 0.0006291957, 0.0001278894, 8.256061e-05, 0.0001148564, 
    0.002091073, 0.002003743, 0.001595046, 0.003834847, 0.0026961, 
    5.384618e-05, 0.0006774247, 0.0004723782, -1.630589e-06, 0.00094001, 
    0.004788341, -7.043845e-05, 0.007164919, 0.0004197746, 0.004923885, 
    -1.175925e-05, 0, -0.0001308259,
  0, 0, 0, -7.418493e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.849632e-05, 
    6.556978e-05, 0, 0, -9.194177e-05, 0.005098426, -9.182073e-07, 0, 
    -0.0001833894, 0.0002139655, 1.523805e-05, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.885814e-06, 0.0002791039, 
    0.001320244, 0.0004751557, 9.791765e-05, 3.138692e-10, 7.413558e-10, 
    -2.185443e-07, -2.430605e-06, 0.0003728437, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001544959, -2.834877e-05, 0.0002071966, -0.000116082, -1.537285e-05, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.293647e-05, 0, -7.235091e-05, 
    2.00126e-05, 0, 0, 0, 0.0005967339, 2.643361e-05, 0.005176361, 
    0.006718998, 0.00148391, 0.005525313, -3.757672e-05, 0, 0, 0,
  0.003997725, 0.009915698, 0.005466089, 0.01488982, 0.00275123, 0.005403784, 
    0.006279323, 0.002398605, 0.0006583925, 0.001524008, 0.001911468, 
    0.002315218, 0.002266477, 0.0001012243, 0.001310442, 0.001403501, 
    0.000932765, 7.743095e-05, 0.004379264, 0.005299206, 0.008674573, 
    0.01217584, 0.01935153, 0.01926379, 0.01063958, 0.005540519, 0.001587222, 
    -5.808456e-05, 0.0009030345,
  0.05619432, 0.05501853, 0.03539766, 0.04305145, 0.08185543, 0.06462079, 
    0.04267138, 0.03199598, 0.02012949, 0.0287449, 0.01830653, 0.03101971, 
    0.006247136, 0.008227002, 0.01262236, 0.01708243, 0.01743662, 0.02836078, 
    0.02678947, 0.04010009, 0.07394849, 0.07823154, 0.1272055, 0.05951186, 
    0.05213836, 0.04403932, 0.05937076, 0.04430328, 0.05596556,
  0.1144942, 0.1077542, 0.09322108, 0.1146901, 0.1471963, 0.08500378, 
    0.07561576, 0.06639144, 0.05609326, 0.06430069, 0.06919697, 0.05114827, 
    0.02338762, 0.02626881, 0.06749962, 0.1130307, 0.08669673, 0.09055835, 
    0.1410798, 0.2510309, 0.1978051, 0.1931255, 0.1410623, 0.08754058, 
    0.1132199, 0.08729317, 0.09624903, 0.1299124, 0.1328444,
  0.03690279, 0.0269228, 0.01580799, 0.05993424, 0.112383, 0.0706308, 
    0.0692538, 0.05355239, 0.0959351, 0.08715247, 0.07915489, 0.04080141, 
    0.02193115, 0.06143779, 0.1589273, 0.1687292, 0.1657959, 0.148066, 
    0.2305251, 0.1588278, 0.1226621, 0.06131144, 0.02085524, 0.04217444, 
    0.02698647, 0.09439054, 0.07471325, 0.05753905, 0.03698755,
  5.216787e-06, 0.001796721, 0.0006044683, 0.0654528, 0.0699798, 0.04437169, 
    0.04579027, 0.02932241, 0.04151158, 0.03432881, 0.01759051, 0.001367466, 
    0.006305457, 0.04360818, 0.09172708, 0.03356931, 0.05642302, 0.07896499, 
    0.03544625, 0.004840555, 0.0002394218, -2.414131e-05, 1.615849e-06, 
    4.727276e-05, 0.00403647, 0.002717398, 0.01114257, 0.003956873, 
    0.0008345835,
  0.0003660303, 0.04298322, 0.0129319, 0.0131876, 0.05049635, 0.02590795, 
    0.06427021, 0.06644835, 0.07813742, 0.05576222, 0.06914958, 0.01920661, 
    0.07861429, 0.1077471, 0.05443343, 0.04455632, 0.02180643, 0.02631779, 
    0.03111926, -9.8677e-05, 7.748986e-07, 1.414927e-06, 0.009712161, 
    0.07562634, 0.04189783, 0.02096582, 0.0008138314, -2.49521e-06, 
    6.938417e-06,
  0.07498789, 0.2828153, 0.2020343, 0.01937066, 0.01407288, 0.09443571, 
    0.07160901, 0.02670899, 0.1887448, 0.2395171, 0.106418, 0.0483449, 
    0.04301675, 0.03326505, 0.08666904, 0.024039, 0.01812623, 0.01965568, 
    0.01018961, 0.002193, 0.0001836591, 2.48975e-06, 0.03229491, 0.2795177, 
    0.1034104, 0.0805912, 0.05826472, 0.03069075, 0.01784003,
  0.1359403, 0.05561632, 0.0578684, 0.05532727, 0.001576376, 0.01369618, 
    0.05875974, 0.0997598, 0.1195927, 0.08967948, 0.09976936, 0.05942647, 
    0.1512441, 0.1448137, 0.1312813, 0.1589815, 0.06500274, 0.07481059, 
    0.03850045, 0.06618664, 0.0488765, 0.1416523, 0.1810087, 0.2304352, 
    0.0187626, 0.02810571, 0.006858276, 0.0146389, 0.2134601,
  0.05112947, 0.008582365, 0.01402752, 0.02893921, 0.05261605, 0.00505546, 
    0.019161, 0.01388404, 0.1158325, 0.1329992, 0.07201395, 0.03283497, 
    0.09155645, 0.02259063, 0.003245052, 0.04489434, 0.06024016, 0.07792938, 
    0.1493904, 0.04825904, 0.01934507, 0.01087306, 0.03008252, 0.1385121, 
    0.1548495, 0.07137886, 0.03489377, 0.03566172, 0.04784176,
  0.05662701, 0.1061042, 0.08927202, 0.1065958, 0.07822442, 0.0496839, 
    0.03368127, 0.005474616, 0.177165, 0.1655826, 0.1728514, 0.2034699, 
    0.1659143, 0.07692385, 0.03694008, 0.09632416, 0.09139241, 0.06628891, 
    0.04373198, 0.01837121, 0.07570978, 0.07005006, 0.05883143, 0.1174355, 
    0.1251768, 0.1082373, 0.09968983, 0.04331895, 0.04536942,
  0.08855677, 0.07531138, 0.06426765, 0.03326606, 0.1229508, 0.143527, 
    0.0338352, 0.1241297, 0.1261194, 0.1018194, 0.1258846, 0.1419197, 
    0.2269815, 0.2566087, 0.1923058, 0.210989, 0.1707551, 0.1888103, 
    0.07801279, 0.05402521, 0.01443074, 0.148185, 0.1458327, 0.182753, 
    0.2010057, 0.140006, 0.1067035, 0.09216349, 0.08278656,
  0.06223563, 0.02522948, 0.03069006, 0.04368018, 0.04464149, 0.07972296, 
    0.05850025, 0.006538372, 0.0005169577, 0.007537469, 0.05293614, 
    0.07315122, 0.08000197, 0.09679464, 0.1325627, 0.1215537, 0.09126483, 
    0.1125701, 0.1079144, 0.001155746, 0.02232771, 0.07005029, 0.04056733, 
    0.02725744, 0.08212758, 0.08655277, 0.04850201, 0.04961778, 0.04663033,
  0.02254395, 0.005215181, 0.0119719, 0.02502278, 0.02866095, 0.0227018, 
    0.01429456, 0.008375495, 3.798574e-05, 0.001419294, 0.006249664, 
    0.009366196, 0.01754651, 0.03543769, 0.03624972, 0.02422942, 0.002256208, 
    0.00814078, 0.0006012337, 0.005553891, 0.003482208, 0.01914334, 
    0.002047999, 0.02181228, 0.02041066, 0.01785968, 0.01020426, 0.002864988, 
    0.02125805,
  0, -7.400727e-09, 0, 0.001689558, 3.638442e-05, 2.307538e-05, 0, 0, 0, 0, 
    0.004708277, 0.006002005, 0.017693, 0.01629623, 0.02020674, 0.009960721, 
    0.001350645, 0.003742282, 0.0003657295, 0.006573922, -8.825174e-05, 
    8.925776e-06, 0.0003103166, 0.0006413762, 0.006981873, -4.601686e-06, 0, 
    0.000525116, -0.0002328086,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -6.028308e-10, 3.878883e-06, 0.0001855813, 
    0.002155571, 0.01373469, 0.01521569, 0.008512678, 0.008420585, 
    0.008174748, 0.005538237, 0.0004476388, 0.00126439, 0.0001694057, 
    -8.213001e-07, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -5.910725e-05, 
    0.0003173416, 0, 0, 0, 0.001018368, 0.002345759, 0.002901543, 
    0.0004425396, 0.0001242175, -3.998135e-05, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001748857, 0, 0, -4.690863e-05, 
    -9.975398e-05, 0.001069571, 0.0001094566, 1.000893e-05, 0.0003304867, 0, 
    0.002936603, 0.01691212, 0.02000928, 0.02718218, 0.02001865, 0.01216953, 
    -0.0001140918, 0.0005581736, -6.525718e-07, -6.334082e-07,
  0.01818406, 0.02575357, 0.02426001, 0.0446986, 0.03698783, 0.0274259, 
    0.02395547, 0.007175019, 0.005208346, 0.005713494, 0.007350715, 
    0.0108497, 0.02266853, 0.02031462, 0.01788196, 0.02120329, 0.01831216, 
    0.007746987, 0.01491706, 0.01593589, 0.02898238, 0.03007414, 0.04568348, 
    0.04439809, 0.03255279, 0.02264971, 0.02108121, 0.007216216, 0.007808686,
  0.1288457, 0.1333676, 0.1222303, 0.1213922, 0.1714187, 0.1622557, 
    0.1216991, 0.1108135, 0.1103857, 0.1060619, 0.09154554, 0.1197176, 
    0.06346523, 0.07787237, 0.09501318, 0.06898458, 0.1063662, 0.1098108, 
    0.0838832, 0.07504702, 0.118914, 0.1223955, 0.1945294, 0.1235396, 
    0.122823, 0.1346388, 0.1193584, 0.08377609, 0.1153952,
  0.1560559, 0.1407297, 0.1386954, 0.1764387, 0.1638733, 0.1002672, 
    0.08367825, 0.08613005, 0.1091467, 0.1174253, 0.1414058, 0.1323926, 
    0.09597345, 0.09329673, 0.09535937, 0.1500688, 0.1181368, 0.1117562, 
    0.1667377, 0.2628042, 0.1908102, 0.1883565, 0.1497183, 0.1433971, 
    0.1379448, 0.08962649, 0.1287204, 0.1545969, 0.1534538,
  0.03146768, 0.0195561, 0.01909806, 0.04395532, 0.09237741, 0.05930037, 
    0.06856973, 0.03221143, 0.1088201, 0.07487217, 0.08268453, 0.03507082, 
    0.02230932, 0.05771921, 0.1448523, 0.1575484, 0.1380451, 0.1354983, 
    0.2056504, 0.1339812, 0.107868, 0.05211147, 0.02061611, 0.03723666, 
    0.0189431, 0.09247954, 0.06515134, 0.05086383, 0.04673744,
  6.871177e-06, 5.481387e-05, 0.0001835781, 0.05194446, 0.06131246, 
    0.03607757, 0.0388137, 0.03111048, 0.05382728, 0.03152531, 0.02540269, 
    0.005441454, 0.01632948, 0.05560483, 0.09062052, 0.03478478, 0.0536247, 
    0.06098917, 0.02271872, 0.007912494, 9.629909e-05, 1.848247e-05, 
    8.432986e-08, 0.0001820157, 0.004139642, 0.002325418, 0.01309461, 
    0.000857644, 5.158981e-05,
  0.0001092488, 0.02965502, 0.01213438, 0.02023306, 0.05235775, 0.01937647, 
    0.06087449, 0.06066529, 0.07111926, 0.04116669, 0.06631669, 0.01959337, 
    0.08283328, 0.07736212, 0.0440265, 0.03017501, 0.02119046, 0.02291008, 
    0.02983197, -0.0001212353, 5.913885e-07, 1.134475e-06, 0.0003690973, 
    0.0551172, 0.02758193, 0.008408741, 0.004712424, 9.770427e-06, 
    7.729633e-06,
  0.0522188, 0.2365279, 0.1625522, 0.02598847, 0.01064491, 0.08136608, 
    0.06117986, 0.02094429, 0.1362242, 0.1880029, 0.09573967, 0.04195862, 
    0.03574325, 0.02987337, 0.07214198, 0.02431158, 0.01645996, 0.01846882, 
    0.009485703, 0.00302284, 3.285167e-05, 4.019995e-06, 0.01565887, 
    0.2472625, 0.09744217, 0.08516654, 0.05309222, 0.02560291, 0.01439648,
  0.133429, 0.0373817, 0.04419945, 0.0410049, 0.001281985, 0.01073744, 
    0.04547013, 0.07394404, 0.0972349, 0.07155196, 0.09660413, 0.04423886, 
    0.133479, 0.1396524, 0.1238482, 0.1359269, 0.05222026, 0.07255464, 
    0.0491451, 0.05232754, 0.03384784, 0.1326378, 0.1340823, 0.1715384, 
    0.02011145, 0.0183849, 0.003113457, 0.01206149, 0.1745108,
  0.04726122, 0.005267596, 0.01685796, 0.01552002, 0.03603525, 2.422058e-05, 
    0.02301532, 0.01186229, 0.08659124, 0.1322455, 0.06718774, 0.02351336, 
    0.08212301, 0.009884492, 0.003260448, 0.03197537, 0.03757418, 0.05073303, 
    0.1184059, 0.02695853, 0.02393759, 0.01130031, 0.03144703, 0.1191688, 
    0.1194951, 0.07261981, 0.03238802, 0.02488128, 0.03434123,
  0.05253949, 0.09262948, 0.08386858, 0.09712787, 0.05353174, 0.03451903, 
    0.02828675, 0.01192749, 0.3049695, 0.1430473, 0.1573088, 0.2032367, 
    0.1651214, 0.0551603, 0.0305652, 0.07689022, 0.06616618, 0.05091303, 
    0.03512537, 0.01470575, 0.06211053, 0.05429175, 0.0507969, 0.1103709, 
    0.1221326, 0.08657736, 0.07757506, 0.03229424, 0.0371832,
  0.143877, 0.0982419, 0.09506894, 0.07880313, 0.1076897, 0.1220512, 
    0.06760293, 0.1381353, 0.130649, 0.1466263, 0.1315426, 0.1415825, 
    0.2029746, 0.2505188, 0.1989526, 0.1866342, 0.172729, 0.1877466, 
    0.07283399, 0.09303793, 0.06135166, 0.1453034, 0.1424652, 0.1874706, 
    0.2027863, 0.1605624, 0.11581, 0.1055675, 0.1009224,
  0.188743, 0.0710831, 0.1054186, 0.1004544, 0.09625365, 0.1195656, 
    0.1284828, 0.02367866, 0.01771903, 0.05894008, 0.1103714, 0.1185893, 
    0.1480847, 0.1311669, 0.14891, 0.1589285, 0.1542036, 0.175698, 0.1645169, 
    0.03497531, 0.1103316, 0.1261596, 0.07834855, 0.06732658, 0.1324333, 
    0.1243594, 0.0876075, 0.119672, 0.165378,
  0.1003978, 0.0558469, 0.07838932, 0.07553129, 0.07590602, 0.06908557, 
    0.05477463, 0.07228486, 0.02049383, 0.005566957, 0.02365372, 0.02728486, 
    0.04902764, 0.1281706, 0.0655177, 0.04877621, 0.03146023, 0.04889194, 
    0.0295424, 0.05150001, 0.04400908, 0.05187279, 0.04204677, 0.05068749, 
    0.05690331, 0.128529, 0.0618431, 0.1006383, 0.1089534,
  0.03501239, 0.02203855, 0.000462591, 0.006144471, 0.00957031, 0.01385699, 
    0.02297824, 0.01066023, 0.009352716, 0.002055772, 0.01162833, 0.01030984, 
    0.01742781, 0.02216892, 0.04024642, 0.0335935, 0.02245224, 0.03740627, 
    0.03969246, 0.07605492, 0.04215219, 0.02767166, 0.05732528, 0.04009459, 
    0.03074053, 6.842914e-06, -1.283141e-06, 0.02428612, 0.04854867,
  -9.941949e-06, 3.703076e-05, 0.0036381, 0.004653781, 0.00357483, 
    2.653622e-05, 0, -2.997465e-07, -2.210508e-05, 0.0004402148, 0.00178198, 
    0.004065124, 0.01529561, 0.01714066, 0.02568115, 0.02901613, 0.02892338, 
    0.01016219, 0.00997488, 0.01097139, 0.01535221, 0.01031402, 0.004509998, 
    0.0003869825, 0.0002107889, -1.658705e-06, -2.382641e-07, -0.0001669621, 
    6.290605e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.000138759, 
    0.003218802, -4.61808e-05, -1.687132e-05, -1.358219e-05, 0.005757904, 
    0.01857581, 0.01667231, 0.0185855, 0.01963034, -0.0008959009, 0,
  0, 0.0001292234, -1.238942e-05, 8.395118e-05, 0, 0, 0, 0, 0, 0.0006851953, 
    0, -1.420797e-05, 0.0002015892, 0.008204882, 0.01111833, 0.01136381, 
    0.008527477, 0.002298265, -3.029967e-05, 0.01056821, 0.04506465, 
    0.064767, 0.04574759, 0.03726546, 0.02848391, 0.01081867, 0.005922784, 
    0.004649544, 0.0004245199,
  0.04363853, 0.05207733, 0.06255685, 0.09827253, 0.107747, 0.08509701, 
    0.06173994, 0.04444014, 0.04354368, 0.03565697, 0.05578038, 0.08638102, 
    0.1658738, 0.1711398, 0.1149906, 0.1071744, 0.09604746, 0.04130907, 
    0.05347458, 0.08537493, 0.0739715, 0.09349109, 0.11365, 0.1125386, 
    0.09480514, 0.06461077, 0.0636586, 0.07119234, 0.03181868,
  0.1750047, 0.1909881, 0.1838431, 0.2165461, 0.2045976, 0.2122972, 
    0.1620147, 0.1679386, 0.1508296, 0.1818458, 0.1825821, 0.1967463, 
    0.1901998, 0.1301696, 0.1412681, 0.1341645, 0.140417, 0.139204, 
    0.1333267, 0.1089501, 0.1416726, 0.1489135, 0.2407218, 0.1779265, 
    0.1831797, 0.2022215, 0.178634, 0.1564098, 0.1749866,
  0.1521084, 0.1248972, 0.1372435, 0.157632, 0.1457797, 0.08115289, 
    0.08085127, 0.07942105, 0.1079429, 0.1120385, 0.14662, 0.1514475, 
    0.1259994, 0.09156185, 0.1199619, 0.1883565, 0.1268306, 0.1054131, 
    0.1787778, 0.2439336, 0.1885464, 0.1765378, 0.1574573, 0.1623528, 
    0.1382902, 0.08937185, 0.1242876, 0.1627833, 0.1535121,
  0.01768802, 0.006641335, 0.01353817, 0.03344186, 0.07824306, 0.0468462, 
    0.06607138, 0.02381522, 0.09925746, 0.06320966, 0.05996126, 0.02673952, 
    0.02023497, 0.05351948, 0.1224397, 0.1446834, 0.1187237, 0.1269296, 
    0.1913668, 0.1130129, 0.1120361, 0.0667284, 0.01420355, 0.03670931, 
    0.01685543, 0.07865186, 0.05064478, 0.04395083, 0.03631604,
  2.249318e-06, 4.726417e-06, 9.029372e-05, 0.03689016, 0.04788518, 
    0.02587455, 0.03392771, 0.02326288, 0.05041755, 0.03930168, 0.02853899, 
    0.004958905, 0.01276682, 0.07376119, 0.08676486, 0.02419223, 0.05071909, 
    0.05952591, 0.01713213, 0.01019406, 0.000336728, 1.412054e-05, 
    3.960085e-09, 0.003234475, 0.005283413, 0.00263599, 0.01539826, 
    0.0004211765, 3.213957e-06,
  2.835827e-05, 0.02306312, 0.008997773, 0.03029291, 0.05194626, 0.01914012, 
    0.05350335, 0.05662923, 0.06477219, 0.03091294, 0.07068137, 0.02140402, 
    0.08550192, 0.05043622, 0.03452147, 0.01919118, 0.0211046, 0.02090444, 
    0.02879648, -5.16291e-05, 2.93129e-07, 3.752054e-07, -3.397152e-05, 
    0.04235831, 0.01596453, 0.002306046, 0.009451807, 2.73326e-05, 
    5.983551e-06,
  0.03745591, 0.2125756, 0.1421635, 0.02819255, 0.008674851, 0.06639657, 
    0.04999226, 0.01794621, 0.09125171, 0.1469229, 0.08535878, 0.03497559, 
    0.02348669, 0.0201783, 0.05576022, 0.02034293, 0.01571511, 0.01268608, 
    0.002123937, 0.005797111, 8.445321e-05, 0.0006625769, 0.01304883, 
    0.2039539, 0.09537423, 0.08826383, 0.05157178, 0.02235057, 0.01171958,
  0.0871607, 0.02247819, 0.02976846, 0.03850636, 0.002274449, 0.007545243, 
    0.03268864, 0.04944956, 0.07453968, 0.05655912, 0.09420282, 0.03368896, 
    0.1096465, 0.1267359, 0.1218262, 0.09450696, 0.04333116, 0.06147262, 
    0.0682402, 0.0417098, 0.01971719, 0.1135426, 0.1037634, 0.1183893, 
    0.01449449, 0.01262262, 0.001549075, 0.008103106, 0.1417022,
  0.0342611, 0.002873079, 0.01584625, 0.005754086, 0.02362821, 4.831554e-06, 
    0.01973391, 0.01422383, 0.06601086, 0.1374127, 0.05735235, 0.01920045, 
    0.06780145, 0.006606648, 0.002726734, 0.02555659, 0.02426215, 0.04516026, 
    0.06525875, 0.009099177, 0.01334294, 0.01134732, 0.0248853, 0.1081533, 
    0.114696, 0.07756671, 0.01165934, 0.01116862, 0.03226351,
  0.0431052, 0.06598423, 0.07316034, 0.07471649, 0.03515749, 0.02830223, 
    0.03139006, 0.04098184, 0.3354831, 0.1345993, 0.1448773, 0.2065648, 
    0.1719164, 0.04615342, 0.0301298, 0.06049022, 0.04938695, 0.0364049, 
    0.02899254, 0.01250346, 0.05052857, 0.04063779, 0.04422963, 0.09223759, 
    0.1049232, 0.07031647, 0.05605527, 0.02205811, 0.02845173,
  0.1371652, 0.09534305, 0.09147483, 0.1304242, 0.09721787, 0.1041136, 
    0.1080315, 0.1088349, 0.1155146, 0.1415342, 0.1262595, 0.1285341, 
    0.1856554, 0.2470115, 0.2025302, 0.1779284, 0.1424496, 0.1745571, 
    0.05992018, 0.1044867, 0.09596057, 0.1305935, 0.1315221, 0.1750757, 
    0.1877739, 0.152299, 0.1068592, 0.09568466, 0.09017453,
  0.206755, 0.143065, 0.1291221, 0.149226, 0.1092378, 0.1164565, 0.1293598, 
    0.06930287, 0.07153456, 0.1401427, 0.1766805, 0.1845046, 0.1718206, 
    0.1444865, 0.159418, 0.1834435, 0.1824483, 0.1943681, 0.1757964, 
    0.1169283, 0.1780272, 0.1282952, 0.1113906, 0.1292619, 0.1631665, 
    0.1319761, 0.1341705, 0.1613974, 0.2062467,
  0.1703484, 0.1111083, 0.1141199, 0.1502897, 0.1585872, 0.1178252, 
    0.1222689, 0.1170185, 0.08564885, 0.0643425, 0.09894879, 0.07019306, 
    0.0964268, 0.1592193, 0.1059998, 0.08411831, 0.09057344, 0.1047094, 
    0.07442623, 0.07988302, 0.07603465, 0.1077941, 0.06377053, 0.08617926, 
    0.169426, 0.2027968, 0.1312117, 0.233476, 0.1585837,
  0.135195, 0.08063396, 0.03839853, 0.03664285, 0.02628991, 0.028153, 
    0.05295287, 0.01643012, 0.01736088, 0.02196338, 0.01652339, 0.01775747, 
    0.03959464, 0.08081127, 0.07417437, 0.05479404, 0.07814112, 0.08703791, 
    0.1038343, 0.1276566, 0.06812782, 0.07587484, 0.09845524, 0.06990417, 
    0.05528706, 0.001447187, -7.100006e-05, 0.1488747, 0.1825164,
  0.002114012, 0.006083157, 0.008438936, 0.005825175, 0.01091905, 
    0.005050242, 0.02016718, 0.03054606, 0.02767782, 0.03235868, 0.02922668, 
    0.02418167, 0.03142793, 0.03124107, 0.03851391, 0.05499523, 0.0719415, 
    0.08088359, 0.06927461, 0.07345548, 0.0761857, 0.06806575, 0.02244257, 
    0.008097559, 0.00903579, 0.001493451, -0.0008081649, 0.003628771, 
    0.008591644,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1.327729e-08, 0, 
    0.0004856891, 0.004371252, -7.309947e-05, -0.0003383333, -0.0002163427, 
    0.01728766, 0.06871218, 0.06191072, 0.02481723, 0.03304776, 0.01613803, 
    0.0001156818,
  0.004225461, 0.02460781, 0.02075418, 0.004445989, -8.588632e-05, 0, 
    -6.332803e-05, 0, -5.753645e-05, 0.001170465, -2.641887e-05, 
    -0.000320504, 0.009855953, 0.07002956, 0.0793936, 0.06313273, 0.04416296, 
    0.02427321, 0.01443726, 0.04532505, 0.1063231, 0.1643349, 0.1404934, 
    0.09365225, 0.08305161, 0.04809386, 0.05059417, 0.03357939, 0.01361759,
  0.08997391, 0.118604, 0.1243244, 0.1382787, 0.1522415, 0.1374856, 
    0.09474743, 0.1083496, 0.1201804, 0.1038786, 0.1529263, 0.2215577, 
    0.2798959, 0.2566527, 0.1810105, 0.2105678, 0.2126949, 0.1500986, 
    0.181307, 0.1726265, 0.1429867, 0.1470718, 0.1704943, 0.1891566, 
    0.1967122, 0.1689614, 0.1314285, 0.1502848, 0.06847596,
  0.2093402, 0.2116615, 0.200803, 0.2249211, 0.2109125, 0.1924913, 0.1694107, 
    0.1773654, 0.177306, 0.1931894, 0.2175878, 0.2486188, 0.1803167, 
    0.1317434, 0.1263703, 0.1294903, 0.1450284, 0.1489287, 0.1637087, 
    0.138822, 0.1694965, 0.1989474, 0.2769651, 0.2292518, 0.1918206, 
    0.2170715, 0.1889774, 0.1749575, 0.2034654,
  0.1582822, 0.1232094, 0.1186311, 0.1350224, 0.1282254, 0.07764661, 
    0.06788865, 0.07523967, 0.09036138, 0.105989, 0.1322725, 0.1431944, 
    0.1261349, 0.07528478, 0.1300698, 0.1931465, 0.1276488, 0.09164543, 
    0.1622966, 0.2232529, 0.1753571, 0.1743806, 0.1530882, 0.1579256, 
    0.1246447, 0.08924389, 0.1226024, 0.1516294, 0.1469908,
  0.007612949, 0.0006217818, 0.005970215, 0.02394534, 0.06952184, 0.03771272, 
    0.06504212, 0.02408666, 0.08748389, 0.04841975, 0.03541277, 0.0258451, 
    0.02338752, 0.04521501, 0.1046987, 0.1387793, 0.1250203, 0.1293937, 
    0.1754083, 0.09411679, 0.1063004, 0.05618303, 0.0111239, 0.04007566, 
    0.01577302, 0.06779738, 0.04693437, 0.04851528, 0.03105341,
  4.797918e-07, 9.974124e-06, 0.0001721443, 0.02857909, 0.03998687, 
    0.02652694, 0.02965895, 0.01382289, 0.05129877, 0.02978276, 0.02511604, 
    0.01200448, 0.01450551, 0.07652392, 0.08167, 0.01958686, 0.04750214, 
    0.05122207, 0.0112699, 0.00593783, 0.0003186033, 9.123586e-06, 
    2.828522e-08, 0.01008742, 0.006980394, 0.001805008, 0.01493123, 
    0.002598282, 5.62729e-07,
  -6.683709e-06, 0.01833029, 0.007905155, 0.04033486, 0.06057452, 0.01621127, 
    0.04832428, 0.05427726, 0.06437374, 0.02418825, 0.06666171, 0.01455996, 
    0.09390147, 0.03372705, 0.02926087, 0.01252155, 0.0211725, 0.01940657, 
    0.02953353, 0.004064463, -2.652887e-07, 1.893725e-07, 0.001043396, 
    0.04176223, 0.006830772, 0.001340318, 0.0166498, 0.001060599, 5.891759e-07,
  0.02910872, 0.1755204, 0.1348988, 0.03454013, 0.008072911, 0.06160332, 
    0.04678268, 0.01452541, 0.06912811, 0.1331652, 0.08079885, 0.03105841, 
    0.01548097, 0.0152356, 0.04491485, 0.01757986, 0.01477657, 0.008743405, 
    0.0002891214, 0.006782011, 0.0006790033, 0.0006506843, 0.01982832, 
    0.1776919, 0.0905749, 0.09655324, 0.0579137, 0.02661209, 0.01468141,
  0.05961092, 0.01604277, 0.02701863, 0.03123279, 0.002063937, 0.005981598, 
    0.02406823, 0.04485483, 0.06039925, 0.04969947, 0.09620316, 0.02687718, 
    0.09862123, 0.1140207, 0.1175417, 0.08490245, 0.04192095, 0.03666753, 
    0.06911866, 0.03301342, 0.01300262, 0.09836277, 0.07601964, 0.08793603, 
    0.01545801, 0.007269735, 0.003786453, 0.005017472, 0.1143792,
  0.0241145, 0.005120781, 0.01696684, 0.003180757, 0.009536515, 3.868518e-06, 
    0.01153946, 0.01571587, 0.05221817, 0.1400542, 0.03926379, 0.01599293, 
    0.06297375, 0.005143708, 0.001989012, 0.02193479, 0.01374982, 0.03989256, 
    0.02846296, 0.0003466124, 0.007143185, 0.01280154, 0.01905455, 
    0.09573583, 0.08363932, 0.04319055, 0.005383682, 0.007056362, 0.02430687,
  0.02739264, 0.05505599, 0.07153133, 0.06652042, 0.02865012, 0.02403294, 
    0.03442209, 0.08369327, 0.3307353, 0.1213258, 0.1251207, 0.1934994, 
    0.1505077, 0.02921944, 0.01486291, 0.04824011, 0.03898469, 0.03087716, 
    0.01863253, 0.006114581, 0.03903832, 0.0297616, 0.03487148, 0.07997031, 
    0.08799802, 0.04372882, 0.0346392, 0.007724171, 0.01848205,
  0.1237356, 0.08454184, 0.07866176, 0.1241861, 0.09097911, 0.0958514, 
    0.1317906, 0.09045386, 0.1002626, 0.1193871, 0.1190048, 0.1188921, 
    0.1781969, 0.2359981, 0.1756734, 0.1602051, 0.1227501, 0.1713124, 
    0.05666135, 0.09754729, 0.1207363, 0.1286312, 0.1098422, 0.1570928, 
    0.1853515, 0.1521582, 0.1110023, 0.09174366, 0.07742798,
  0.1753337, 0.1431251, 0.1254295, 0.1265583, 0.1018539, 0.1126686, 
    0.1268202, 0.09679917, 0.1389815, 0.1590221, 0.2304129, 0.2121212, 
    0.1787874, 0.1485851, 0.1554713, 0.1885513, 0.1979363, 0.1909559, 
    0.1653676, 0.1225353, 0.16691, 0.1186892, 0.1188063, 0.1540417, 
    0.1813325, 0.1313208, 0.1450771, 0.156372, 0.1916608,
  0.1521825, 0.1266461, 0.1059881, 0.160816, 0.1734429, 0.1799188, 0.1912708, 
    0.1989564, 0.143946, 0.1487282, 0.1371257, 0.09562336, 0.125823, 
    0.2514105, 0.1403002, 0.09808964, 0.1450748, 0.1618558, 0.1519714, 
    0.1366082, 0.109761, 0.1615287, 0.09803247, 0.1192788, 0.2189626, 
    0.2326901, 0.1290997, 0.2364883, 0.1485724,
  0.223938, 0.1319623, 0.06845511, 0.07811537, 0.06800622, 0.05737085, 
    0.08573413, 0.06757804, 0.05810715, 0.08103427, 0.0569163, 0.09138384, 
    0.1037003, 0.139495, 0.1050436, 0.1284903, 0.119665, 0.1465263, 
    0.1366032, 0.1062816, 0.08250576, 0.07360556, 0.1253585, 0.08062942, 
    0.10005, 0.007532703, -5.435139e-05, 0.2608021, 0.255885,
  0.0653544, 0.07062615, 0.06599375, 0.05776398, 0.08306511, 0.07508402, 
    0.07335383, 0.1028542, 0.08091582, 0.07560299, 0.0726496, 0.1289927, 
    0.1746808, 0.1990409, 0.1910635, 0.1659848, 0.1527306, 0.1290225, 
    0.1097335, 0.09456103, 0.09798031, 0.1090092, 0.06097235, 0.03440639, 
    0.02507661, 0.01017021, 0.006906386, 0.0176214, 0.08398272,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  -8.729692e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.40283e-06, 
    0.0001619727, 0.0001712284, 0.002318701, 0.001593886, 0.008189383, 
    -0.0001706173, 0.0001186324, 0.0008216398, 0.04498947, 0.1288703, 
    0.1189732, 0.06089605, 0.06251755, 0.0327487, 0.0008003354,
  0.07026052, 0.09900336, 0.09351543, 0.03730379, -0.0007394229, 
    -3.073357e-05, 0.02060524, -3.825761e-05, -0.0001663084, 0.0008355228, 
    0.001632127, 0.003894861, 0.04253659, 0.1283818, 0.1592246, 0.1253159, 
    0.09397197, 0.06553752, 0.0466105, 0.07468355, 0.2070518, 0.2135803, 
    0.2248166, 0.1865823, 0.1681264, 0.1290627, 0.1631036, 0.1175378, 
    0.09641469,
  0.1614549, 0.1494795, 0.1684567, 0.1565143, 0.1818948, 0.1712233, 
    0.1496681, 0.1399887, 0.1664484, 0.1519273, 0.2167917, 0.2731895, 
    0.2897078, 0.283015, 0.1920926, 0.2225299, 0.2256209, 0.1710156, 
    0.2215778, 0.244481, 0.2148665, 0.2215721, 0.2325063, 0.2428778, 
    0.2639461, 0.2397419, 0.1766133, 0.2104605, 0.1563216,
  0.2049771, 0.2173902, 0.193373, 0.2110705, 0.1978832, 0.1928123, 0.1643015, 
    0.1658311, 0.1805904, 0.1950776, 0.2424009, 0.2524194, 0.1672022, 
    0.1236551, 0.1231603, 0.1286811, 0.1487834, 0.149525, 0.1585615, 
    0.1477727, 0.1790886, 0.2164305, 0.2693334, 0.2323412, 0.1904394, 
    0.2075162, 0.1897368, 0.1904385, 0.2009348,
  0.1661019, 0.1165822, 0.1123427, 0.1148582, 0.1139908, 0.07207163, 
    0.07186186, 0.07429545, 0.08428044, 0.08433241, 0.1132232, 0.1256245, 
    0.1153613, 0.06931159, 0.1212231, 0.186801, 0.1209833, 0.08723743, 
    0.1546387, 0.2006201, 0.1589274, 0.1857319, 0.1335707, 0.1542115, 
    0.1208061, 0.07844787, 0.1149316, 0.1395887, 0.1364763,
  0.006315259, 0.003817461, 0.006582005, 0.02223582, 0.06301215, 0.03463406, 
    0.05652194, 0.01327956, 0.07481578, 0.04210972, 0.02875892, 0.02474975, 
    0.02434767, 0.04425864, 0.09777009, 0.1425111, 0.1201778, 0.1212308, 
    0.1611838, 0.07472288, 0.09630811, 0.05734251, 0.01572582, 0.0499124, 
    0.01801002, 0.06248706, 0.04563566, 0.05212552, 0.03627761,
  1.035913e-07, 6.300197e-06, 0.0004076972, 0.02028364, 0.0362868, 
    0.02724751, 0.03735238, 0.01329119, 0.04486821, 0.02055818, 0.02888003, 
    0.01079397, 0.0174634, 0.07963672, 0.05889866, 0.01343388, 0.05208421, 
    0.04091264, 0.01146993, 0.001030103, 0.0003197714, 7.589343e-06, 
    8.001653e-09, 0.01252186, 0.007433295, 0.0005869732, 0.01376675, 
    0.002698876, 2.435216e-07,
  -2.661085e-05, 0.02652466, 0.003513853, 0.04676463, 0.05672977, 0.01675378, 
    0.04557173, 0.0539514, 0.0634746, 0.02818542, 0.06165162, 0.01571694, 
    0.09818278, 0.02596746, 0.02463668, 0.01180789, 0.02067122, 0.01967707, 
    0.03103442, 0.009558755, -8.660287e-05, 9.645167e-07, 0.0001343127, 
    0.03307893, 0.004430126, 0.001112652, 0.01771123, 0.0002695258, 
    2.298215e-06,
  0.02536505, 0.1722901, 0.132791, 0.0450703, 0.009550233, 0.05775253, 
    0.05027578, 0.01207118, 0.05828988, 0.1208951, 0.07520759, 0.02871766, 
    0.01255992, 0.01220034, 0.04053855, 0.0182987, 0.01471687, 0.01148136, 
    0.008642917, 0.003418369, 3.223359e-05, 0.002470068, 0.03886015, 
    0.1565458, 0.09279254, 0.1058472, 0.07255585, 0.02441172, 0.0175862,
  0.03553765, 0.01782301, 0.03908102, 0.03298614, 0.002465405, 0.005654934, 
    0.01793717, 0.03563318, 0.05321604, 0.04736538, 0.09693927, 0.02611562, 
    0.08346177, 0.09716623, 0.1164248, 0.09530966, 0.04371808, 0.01933521, 
    0.0764986, 0.02868042, 0.009612277, 0.08936106, 0.06083427, 0.07486589, 
    0.01577434, 0.006868919, 0.006062623, 0.01058826, 0.08973152,
  0.02508003, 0.01447009, 0.01658164, 0.005608308, 0.00170007, 1.647668e-06, 
    0.004308256, 0.01635274, 0.06035107, 0.1369661, 0.02685686, 0.01593204, 
    0.05631229, 0.003437575, 0.006148007, 0.02215733, 0.01694926, 0.02996982, 
    0.01568351, 0.0002087476, 0.008603926, 0.01550547, 0.01646885, 
    0.09863082, 0.06706572, 0.03109255, 0.001284688, 0.01502379, 0.01619883,
  0.01956161, 0.05588796, 0.06264237, 0.06135697, 0.02585901, 0.02145306, 
    0.05403228, 0.1364942, 0.327924, 0.1136276, 0.1132728, 0.1850789, 
    0.1545752, 0.02436262, 0.00830307, 0.03849946, 0.03091594, 0.01875128, 
    0.01430349, 0.004007497, 0.01956985, 0.02488934, 0.03490626, 0.07317829, 
    0.07677396, 0.04660394, 0.02113155, 0.002162912, 0.009545047,
  0.1142907, 0.08214319, 0.07574331, 0.1090772, 0.08017318, 0.08660536, 
    0.1266313, 0.08381279, 0.09022179, 0.1085307, 0.1213645, 0.1154826, 
    0.1664377, 0.231483, 0.1554795, 0.1538255, 0.1171055, 0.1577527, 
    0.05518486, 0.0944422, 0.114213, 0.1328546, 0.09229583, 0.1507751, 
    0.1842541, 0.1367177, 0.09426446, 0.08855657, 0.08303396,
  0.1475929, 0.1305182, 0.1153651, 0.1144314, 0.09717099, 0.1045466, 
    0.1162527, 0.1146586, 0.1589431, 0.1623419, 0.247476, 0.2210001, 
    0.1758688, 0.134897, 0.1562941, 0.1836482, 0.2114355, 0.1744927, 
    0.1618643, 0.1216625, 0.1488247, 0.1234597, 0.1159962, 0.1611355, 
    0.1909561, 0.1297661, 0.1330535, 0.1386005, 0.1839278,
  0.1390402, 0.116316, 0.1012097, 0.1605594, 0.1714787, 0.1961094, 0.2135435, 
    0.2194071, 0.2089784, 0.2042871, 0.1887414, 0.1163949, 0.15204, 
    0.2697514, 0.1398859, 0.114251, 0.1938737, 0.2207029, 0.182758, 
    0.1446038, 0.1450519, 0.1563462, 0.09784829, 0.1447138, 0.2184665, 
    0.2292045, 0.1171352, 0.2155184, 0.1267589,
  0.2026566, 0.129527, 0.08788808, 0.09405126, 0.09261382, 0.1591227, 
    0.1420494, 0.1333107, 0.1091973, 0.1687859, 0.1054837, 0.1768061, 
    0.1653472, 0.1776705, 0.1094523, 0.1355949, 0.1193867, 0.1548544, 
    0.1566909, 0.1054868, 0.08799273, 0.08276992, 0.1378677, 0.09943384, 
    0.1130559, 0.05256018, 0.007384133, 0.2445559, 0.2260497,
  0.09865055, 0.1206002, 0.1419972, 0.15664, 0.1776008, 0.1686013, 0.113525, 
    0.1361365, 0.1145522, 0.09969313, 0.09787691, 0.1677004, 0.1987576, 
    0.1876644, 0.1892873, 0.167843, 0.1510677, 0.1299496, 0.1061883, 
    0.1084776, 0.115689, 0.1236419, 0.09827814, 0.06051537, 0.04839323, 
    0.01869207, 0.01805485, 0.07263459, 0.1183787,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -8.567094e-06, -8.567094e-06, 
    -8.567094e-06, -8.567094e-06, -8.567094e-06, -8.567094e-06, 
    -8.567094e-06, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.001276528, -3.079629e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.352359e-05, 
    0.01607454, 0.02853291, 0.05103444, 0.05321425, 0.0225978, 0.02049845, 
    0.002041974, 0.005294694, 0.005682768, 0.1125339, 0.2722842, 0.2372203, 
    0.1263725, 0.1079871, 0.03912003, 0.01196019,
  0.1187394, 0.1988253, 0.1632598, 0.09210269, -0.002279156, -0.001447365, 
    0.05750371, -0.0002063174, 8.936937e-05, 0.002681567, 0.005382586, 
    0.007561855, 0.1018383, 0.1759874, 0.1785498, 0.1560848, 0.1316365, 
    0.1250591, 0.1333343, 0.206064, 0.3451073, 0.2757475, 0.2918426, 
    0.2956462, 0.2991337, 0.2186264, 0.2283148, 0.2228284, 0.1989979,
  0.2056546, 0.1723068, 0.2108631, 0.1868759, 0.2363029, 0.1937266, 
    0.1942917, 0.1919569, 0.2097248, 0.2362911, 0.290791, 0.305731, 
    0.3157519, 0.2827299, 0.1892679, 0.221862, 0.2274004, 0.192491, 
    0.2639942, 0.290666, 0.2754177, 0.2803817, 0.2534514, 0.2670432, 
    0.2741165, 0.2562634, 0.2106757, 0.2358553, 0.1946304,
  0.2071559, 0.2229504, 0.2095599, 0.2102239, 0.1860817, 0.1905095, 0.165477, 
    0.1527401, 0.2003649, 0.2062527, 0.2568902, 0.2460349, 0.1651786, 0.1032, 
    0.1063164, 0.1122238, 0.1457453, 0.1384587, 0.1573789, 0.1451616, 
    0.1733595, 0.2213473, 0.2579405, 0.2235118, 0.1896866, 0.2086056, 
    0.1771989, 0.1942415, 0.2034761,
  0.1561638, 0.09632041, 0.09893758, 0.0985698, 0.102321, 0.06431597, 
    0.07524879, 0.07416026, 0.06972036, 0.08525608, 0.1133309, 0.117131, 
    0.1086681, 0.06482504, 0.1127646, 0.1757366, 0.1169387, 0.08746672, 
    0.1415957, 0.1917196, 0.1374276, 0.1647143, 0.1251567, 0.1522639, 
    0.09561375, 0.07690656, 0.105351, 0.1393152, 0.1519988,
  0.004131509, 0.002420249, 0.006398007, 0.02560425, 0.05569452, 0.03029865, 
    0.04633667, 0.005939695, 0.06670322, 0.02864723, 0.02562628, 0.02363081, 
    0.02550945, 0.04295884, 0.08760275, 0.1390027, 0.136601, 0.1111877, 
    0.1440507, 0.07082454, 0.08170288, 0.0544972, 0.007927209, 0.05412804, 
    0.01850986, 0.05271631, 0.04123767, 0.0496231, 0.03119109,
  -1.192569e-07, 2.82458e-06, 0.002552709, 0.01580932, 0.02887483, 
    0.03458691, 0.03531703, 0.01244289, 0.05317133, 0.0042613, 0.03635002, 
    0.01091915, 0.01794936, 0.1041951, 0.03990645, 0.009658814, 0.04606532, 
    0.0351253, 0.009769898, 0.0004263902, 0.000313845, 9.892334e-07, 
    -2.888703e-10, 0.006781992, 0.008528277, 0.0001797757, 0.01313212, 
    0.0001239131, 1.636448e-07,
  7.73847e-06, 0.02859878, 0.002695038, 0.05199493, 0.05720839, 0.01935071, 
    0.04617397, 0.05387438, 0.06106322, 0.02806536, 0.05180513, 0.01805284, 
    0.09653567, 0.02656729, 0.02202667, 0.01157181, 0.01876644, 0.02048627, 
    0.0318759, 0.0138006, 0.0009338805, 1.989521e-07, 0.0007787185, 
    0.03164793, 0.003286306, 0.002661107, 0.00671948, -4.302701e-05, 
    7.261211e-06,
  0.01815371, 0.1568973, 0.1299466, 0.0463383, 0.01282642, 0.06521638, 
    0.04904239, 0.01061487, 0.05223478, 0.1100437, 0.07074033, 0.02748274, 
    0.009973944, 0.01159655, 0.03789972, 0.02209084, 0.01642479, 0.01311729, 
    0.00522568, 0.009020009, 0.001184116, 0.0130065, 0.03837562, 0.1571553, 
    0.08668478, 0.1097039, 0.07699273, 0.02363056, 0.0131116,
  0.02999317, 0.02072869, 0.04727383, 0.03249457, 0.002885046, 0.005134924, 
    0.01383615, 0.03673307, 0.04965592, 0.04640397, 0.1018445, 0.02581776, 
    0.07639208, 0.08979472, 0.1154541, 0.1111006, 0.03744132, 0.01721593, 
    0.06974164, 0.04160381, 0.01028785, 0.084012, 0.06026495, 0.06660547, 
    0.01214482, 0.009296704, 0.005527988, 0.01098983, 0.08168017,
  0.01034824, 0.02223164, 0.01573533, 0.008247753, 7.853614e-05, 
    6.825798e-07, 0.002218022, 0.01986298, 0.0552121, 0.1488822, 0.02241944, 
    0.0183387, 0.05730441, 0.002089832, 0.002303645, 0.02193914, 0.01634826, 
    0.02722099, 0.009220219, 0.0002084167, 0.0005920202, 0.01856917, 
    0.01976728, 0.09594177, 0.04256842, 0.02421814, 0.00188055, 0.02366582, 
    0.009027326,
  0.02758036, 0.04574963, 0.04864137, 0.05575497, 0.0241129, 0.01880401, 
    0.03353275, 0.146821, 0.3228942, 0.103818, 0.106383, 0.171684, 0.1482425, 
    0.02232411, 0.00230023, 0.04165347, 0.03150481, 0.01276588, 0.008051652, 
    0.0007145457, 0.008170085, 0.01897163, 0.0323376, 0.06650425, 0.06480202, 
    0.04234862, 0.01742001, 0.0002984374, 0.003347341,
  0.1010102, 0.07278647, 0.07202805, 0.1008856, 0.06779735, 0.08144645, 
    0.1225037, 0.07733263, 0.08195397, 0.1060598, 0.1172133, 0.1093676, 
    0.1512088, 0.2190119, 0.1356819, 0.1392951, 0.1004516, 0.137819, 
    0.04468597, 0.08572792, 0.1212958, 0.1332703, 0.08329265, 0.1434073, 
    0.178857, 0.1372901, 0.09541361, 0.08250902, 0.08061615,
  0.1291044, 0.1208543, 0.1094458, 0.1092866, 0.09706187, 0.09790929, 
    0.1103403, 0.1251676, 0.1753782, 0.1550937, 0.2541178, 0.2123, 0.1716444, 
    0.1183306, 0.1551181, 0.1763536, 0.22521, 0.1693407, 0.1503285, 
    0.1242537, 0.1351258, 0.127671, 0.1129557, 0.1660194, 0.1904823, 
    0.1236465, 0.1175328, 0.1324625, 0.1741108,
  0.1405777, 0.1115907, 0.09320911, 0.1647123, 0.1655853, 0.2020662, 
    0.2371529, 0.2270081, 0.2219625, 0.2311696, 0.1920723, 0.1762283, 
    0.167056, 0.2717232, 0.1436147, 0.1166638, 0.2047103, 0.2524397, 
    0.2100317, 0.1663733, 0.1451584, 0.1669463, 0.09606415, 0.1416302, 
    0.206819, 0.2205429, 0.1140403, 0.2043952, 0.121024,
  0.1879147, 0.1243757, 0.09258482, 0.0921725, 0.1080045, 0.1934521, 
    0.1782513, 0.1578705, 0.122258, 0.1843904, 0.1167355, 0.2386246, 
    0.1751787, 0.1779928, 0.107233, 0.1418634, 0.1032685, 0.156031, 
    0.1618937, 0.1178654, 0.09287629, 0.07595506, 0.1432872, 0.1083731, 
    0.1132452, 0.1049879, 0.01952367, 0.2354969, 0.2139011,
  0.08703257, 0.1155177, 0.1427638, 0.1896021, 0.1741597, 0.169672, 
    0.1060097, 0.1308922, 0.1155832, 0.08946197, 0.09488997, 0.1373305, 
    0.18258, 0.1731016, 0.1906799, 0.1729528, 0.1606848, 0.1667579, 
    0.1062446, 0.1034312, 0.1047695, 0.1172811, 0.09942363, 0.07282728, 
    0.07709436, 0.05152435, 0.04650746, 0.08282714, 0.1071225,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -0.0001441262, -0.0001394953, 
    -0.0001348644, -0.0001302336, -0.0001256027, -0.0001209719, -0.000116341, 
    -2.585292e-05, -3.048377e-05, -3.511462e-05, -3.974548e-05, 
    -4.437633e-05, -4.900718e-05, -5.363803e-05, 0,
  0.008009796, -9.111826e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009796174, 
    0.0904834, 0.1165313, 0.09938537, 0.1218199, 0.07755123, 0.07272796, 
    0.02306053, 0.03133618, 0.02971501, 0.1976772, 0.354188, 0.311519, 
    0.2182751, 0.1465946, 0.07392316, 0.03265179,
  0.1868178, 0.2358858, 0.2970845, 0.1769426, -0.001179858, -0.001803121, 
    0.1146846, 0.0006190812, 0.001764904, 0.0203154, 0.03127801, 0.0379033, 
    0.15898, 0.1781628, 0.2196744, 0.2049108, 0.1730529, 0.2163911, 
    0.2593075, 0.3099043, 0.4108098, 0.3126442, 0.316227, 0.3673037, 
    0.3623501, 0.2370464, 0.2306869, 0.259761, 0.2747834,
  0.2134607, 0.2094831, 0.2355635, 0.241221, 0.2864522, 0.2200398, 0.2158699, 
    0.2131001, 0.2294989, 0.25408, 0.301404, 0.3052649, 0.3204169, 0.2837278, 
    0.1900034, 0.2204904, 0.2393278, 0.2027483, 0.2926323, 0.306422, 
    0.3034055, 0.2841061, 0.2797787, 0.2638188, 0.262816, 0.2639825, 
    0.2215727, 0.2601963, 0.180902,
  0.2096837, 0.2169833, 0.2051582, 0.2049134, 0.1815062, 0.1813211, 
    0.1614474, 0.1543686, 0.2192007, 0.2150947, 0.2522209, 0.2511019, 
    0.1531865, 0.1098914, 0.1043395, 0.09839561, 0.1276296, 0.1239888, 
    0.145147, 0.1346501, 0.1834648, 0.2010148, 0.2365121, 0.2057831, 
    0.166928, 0.1930621, 0.168621, 0.1770466, 0.2090851,
  0.1436226, 0.07980472, 0.09148085, 0.08918628, 0.09633245, 0.0501233, 
    0.07376366, 0.06237562, 0.06312833, 0.08030757, 0.09653622, 0.1039752, 
    0.08566979, 0.06493121, 0.1027837, 0.1603037, 0.1136502, 0.0884769, 
    0.1224336, 0.1915787, 0.1266017, 0.1635749, 0.1135344, 0.1485212, 
    0.08268704, 0.07479377, 0.1077888, 0.1292045, 0.1445885,
  0.005295753, 0.0009258099, 0.006244812, 0.0332913, 0.05691277, 0.02967276, 
    0.03481207, 0.004146306, 0.05643018, 0.02392315, 0.01156417, 0.01564391, 
    0.03347024, 0.04210933, 0.08868128, 0.132319, 0.1200385, 0.1056287, 
    0.136481, 0.06408241, 0.07343423, 0.05367856, 0.005715435, 0.05138448, 
    0.01803268, 0.04908487, 0.04211237, 0.04475256, 0.02791658,
  -1.585866e-06, -1.976657e-05, 0.003807247, 0.007192179, 0.03470908, 
    0.04089189, 0.02448379, 0.01899043, 0.05273365, 0.004135271, 0.05039239, 
    0.005322209, 0.01984761, 0.1270097, 0.03541248, 0.008008955, 0.03548619, 
    0.029892, 0.008352518, 0.0004062757, 0.0001863592, -1.740281e-06, 
    -2.615995e-07, 0.0008461324, 0.01362127, 0.0001647025, 0.01325351, 
    0.0001762109, 1.505236e-07,
  6.467228e-05, 0.01837507, 0.003466161, 0.05434192, 0.06774458, 0.03425531, 
    0.04757136, 0.05670661, 0.06004568, 0.03358455, 0.05624687, 0.02455319, 
    0.1129223, 0.03019755, 0.02437605, 0.01107709, 0.01663735, 0.0218636, 
    0.02974589, 0.01360136, 0.0009914478, 2.083972e-06, 0.007684, 0.02554274, 
    0.003270376, 0.00127632, 0.009182854, 1.316824e-05, 2.379353e-05,
  0.02166911, 0.1509427, 0.1410538, 0.04665092, 0.009596983, 0.06653614, 
    0.04961738, 0.01032995, 0.05715548, 0.1100002, 0.06627865, 0.02527162, 
    0.009242661, 0.01126334, 0.03562093, 0.02025086, 0.01504091, 0.01661672, 
    0.003821112, 0.01353215, 0.01064656, 0.01455176, 0.0468679, 0.1802517, 
    0.09877198, 0.1105895, 0.07423922, 0.0346923, 0.01814062,
  0.03477755, 0.02888712, 0.04289548, 0.03691272, 0.00332446, 0.004325763, 
    0.01410591, 0.04110396, 0.05178158, 0.05922215, 0.1065566, 0.02752101, 
    0.08600052, 0.09391514, 0.1269968, 0.1287861, 0.04186669, 0.01558945, 
    0.06914059, 0.05144259, 0.01157615, 0.07854237, 0.06726512, 0.06733898, 
    0.01044678, 0.01003476, 0.007723781, 0.01041035, 0.089255,
  0.005281173, 0.01767338, 0.01810945, 0.0109337, 0.001326111, 4.261808e-07, 
    0.004698022, 0.0181895, 0.06558335, 0.154868, 0.02786627, 0.02201462, 
    0.05973264, 0.002471809, 0.00188709, 0.02557797, 0.01490926, 0.01248501, 
    0.004037917, 0.0002268405, 0.0002021109, 0.01717192, 0.02299834, 
    0.1057375, 0.02490469, 0.01636073, 0.000121737, 0.02145023, 0.009162155,
  0.02599345, 0.03040252, 0.03449715, 0.04353701, 0.028229, 0.02006955, 
    0.01449168, 0.1658344, 0.3250797, 0.1058871, 0.09593183, 0.1579477, 
    0.1425918, 0.02878264, 0.002001588, 0.0336701, 0.02279479, 0.01277658, 
    0.001961506, -1.102284e-05, 0.006210294, 0.01645342, 0.02339035, 
    0.06139649, 0.05765156, 0.02880967, 0.01263054, 0.0003836309, 0.001318763,
  0.08769862, 0.05373585, 0.07031687, 0.09797263, 0.0600928, 0.07693771, 
    0.1158426, 0.06578128, 0.06976368, 0.1080462, 0.112422, 0.09406546, 
    0.1473849, 0.2110366, 0.1314328, 0.1354905, 0.08532216, 0.1222971, 
    0.04432809, 0.07541757, 0.1351407, 0.115832, 0.08779758, 0.1421234, 
    0.1756108, 0.114672, 0.08945061, 0.07446559, 0.07225073,
  0.1198812, 0.1133439, 0.1108687, 0.1036838, 0.101541, 0.1032801, 0.1072116, 
    0.1439312, 0.1808478, 0.1480029, 0.256374, 0.2041023, 0.1633349, 
    0.1069865, 0.1552596, 0.1765074, 0.2099816, 0.1714022, 0.1408255, 
    0.1148634, 0.1314569, 0.1245949, 0.1057814, 0.1727603, 0.1881907, 
    0.1241662, 0.1157058, 0.1191948, 0.1499292,
  0.1402656, 0.1164454, 0.07968428, 0.1696435, 0.1584673, 0.2067651, 
    0.2331454, 0.2229459, 0.2170114, 0.2200291, 0.1913825, 0.1903082, 
    0.1766999, 0.2746298, 0.1568079, 0.1159745, 0.2151598, 0.25862, 
    0.2248797, 0.1705999, 0.1442472, 0.1799295, 0.1003147, 0.1389659, 
    0.2002045, 0.2205945, 0.1219452, 0.1992252, 0.1129106,
  0.1796992, 0.1246919, 0.0915487, 0.0922304, 0.1160766, 0.1906712, 
    0.1931856, 0.1884482, 0.1449581, 0.2083659, 0.1563304, 0.2145359, 
    0.1636007, 0.1631375, 0.1019677, 0.1432004, 0.09595014, 0.1566112, 
    0.1619712, 0.1252926, 0.09800757, 0.07822157, 0.1394413, 0.1176763, 
    0.1074984, 0.1900412, 0.07120575, 0.2242594, 0.1932238,
  0.07120363, 0.0964487, 0.1372612, 0.1888374, 0.1714948, 0.1515456, 
    0.0871889, 0.1039756, 0.1005687, 0.07896999, 0.09745757, 0.1245271, 
    0.1665267, 0.1737029, 0.1842495, 0.175168, 0.1551221, 0.1650929, 
    0.1023507, 0.08493169, 0.09528409, 0.1126762, 0.09723996, 0.06109638, 
    0.06836373, 0.0688207, 0.1043412, 0.07545099, 0.09847473,
  6.52957e-05, 4.926872e-05, 3.324173e-05, 1.721474e-05, 1.187758e-06, 
    -1.483923e-05, -3.086621e-05, -0.0010673, -0.0007091003, -0.0003509005, 
    7.299242e-06, 0.000365499, 0.0007236988, 0.001081899, 5.648239e-06, 
    -0.000173974, -0.0003535962, -0.0005332184, -0.0007128406, -0.0008924628, 
    -0.001072085, 0.0001488842, -1.366635e-05, -0.0001762169, -0.0003387675, 
    -0.0005013181, -0.0006638687, -0.0008264192, 7.811729e-05,
  0.02334857, 0.0001115556, -5.166032e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.691316e-06, 0.008811889, 0.1466924, 0.1438964, 0.1592477, 0.2079227, 
    0.1509933, 0.1208889, 0.07307152, 0.08384346, 0.08836538, 0.2908672, 
    0.3764693, 0.3143412, 0.2244782, 0.1512392, 0.1202112, 0.04085785,
  0.2009714, 0.235838, 0.3480419, 0.2700863, 0.008494233, 0.01921362, 
    0.1598847, 0.0222514, 0.02293374, 0.05457223, 0.07996358, 0.08355178, 
    0.189281, 0.1884012, 0.231678, 0.2110604, 0.206401, 0.2367446, 0.2931616, 
    0.3137462, 0.4087012, 0.3268038, 0.3355904, 0.3715817, 0.3539891, 
    0.2474716, 0.2273853, 0.2674981, 0.2863148,
  0.2157131, 0.2135443, 0.2427123, 0.2517355, 0.2903173, 0.2387062, 
    0.2470163, 0.2379645, 0.2782263, 0.2642144, 0.3144155, 0.32201, 
    0.3241283, 0.2748288, 0.1947787, 0.2196064, 0.248276, 0.2114173, 
    0.3099749, 0.2985733, 0.2863946, 0.2582867, 0.261185, 0.2486844, 
    0.2531053, 0.2671439, 0.217847, 0.2543554, 0.1902148,
  0.2064208, 0.2099213, 0.2089302, 0.2046133, 0.1684601, 0.1797157, 
    0.1590274, 0.1596447, 0.2146405, 0.222849, 0.2416048, 0.2414874, 
    0.1471584, 0.09147161, 0.1004165, 0.09756134, 0.125612, 0.1068241, 
    0.1486392, 0.1426386, 0.1878556, 0.195404, 0.2277459, 0.1917391, 
    0.1612372, 0.177597, 0.1739263, 0.1939669, 0.2059762,
  0.1330518, 0.06471484, 0.08933085, 0.08808579, 0.08868722, 0.05516358, 
    0.06625839, 0.05889655, 0.05663809, 0.07035444, 0.0944993, 0.09378165, 
    0.08369074, 0.06097197, 0.1012874, 0.1522155, 0.1032421, 0.09354714, 
    0.1257015, 0.1683414, 0.1149958, 0.1596876, 0.09936017, 0.1473757, 
    0.08353013, 0.07450511, 0.1059187, 0.1266132, 0.1483817,
  0.002697796, 0.001234669, 0.004768396, 0.03725293, 0.05152164, 0.03497491, 
    0.02233876, 0.006602108, 0.05911974, 0.02740846, 0.01623875, 0.01248042, 
    0.03427143, 0.04870953, 0.09371668, 0.1347544, 0.113248, 0.09965377, 
    0.1339549, 0.07008521, 0.07136273, 0.05630222, 0.009757886, 0.0404207, 
    0.02268255, 0.04659355, 0.03993734, 0.04678866, 0.02487706,
  9.036764e-08, -1.708649e-05, 0.005490124, 0.00253504, 0.04286761, 
    0.04686335, 0.01472403, 0.01377513, 0.05777621, 0.003780503, 0.05218294, 
    0.001891941, 0.02169592, 0.1342848, 0.03631286, 0.007292789, 0.03361902, 
    0.02799852, 0.01097484, 0.0004844062, 0.0002030313, -3.075142e-07, 
    1.828049e-08, 1.169919e-05, 0.01798724, 0.0003052197, 0.01407471, 
    0.001006223, 2.211124e-07,
  0.0002700266, 0.01882944, 0.005586914, 0.06396497, 0.07568538, 0.04765807, 
    0.06458318, 0.06628938, 0.06658584, 0.04960854, 0.06735987, 0.0267701, 
    0.1364059, 0.04218969, 0.02999399, 0.01534072, 0.02013534, 0.02335253, 
    0.02528903, 0.01647594, 0.0007422434, 2.167866e-07, 0.001733073, 
    0.03032413, 0.005018781, 0.001393493, 0.016946, 0.0001589377, 0.0008309478,
  0.03372872, 0.1840121, 0.1770884, 0.03405701, 0.01315189, 0.07705092, 
    0.05197034, 0.01310005, 0.07868806, 0.1248977, 0.08019707, 0.0296321, 
    0.01367287, 0.01250289, 0.03455161, 0.02030008, 0.01459969, 0.01670755, 
    0.01350501, 0.01524465, 0.01609007, 0.01518294, 0.05882774, 0.2040172, 
    0.1112729, 0.1154923, 0.07957737, 0.03175058, 0.0222158,
  0.03420123, 0.0413617, 0.03492671, 0.1023254, 0.004318727, 0.005185806, 
    0.01653423, 0.05783089, 0.06374102, 0.0748182, 0.1220367, 0.03340371, 
    0.1085611, 0.1162607, 0.1503729, 0.1453848, 0.04952538, 0.01962885, 
    0.06844341, 0.05099265, 0.01837563, 0.0901888, 0.09143345, 0.08228828, 
    0.01045835, 0.01467478, 0.01021602, 0.01554837, 0.09924614,
  0.008321711, 0.006953743, 0.0097115, 0.007149704, 0.01120094, 1.874445e-06, 
    0.004992444, 0.01838586, 0.08860323, 0.1793115, 0.03914911, 0.02667638, 
    0.06705926, 0.003672724, 0.003334477, 0.03785487, 0.01188572, 0.01232122, 
    0.002014966, 0.000413083, 0.002132731, 0.01706839, 0.03063182, 0.1218054, 
    0.01656298, 0.01312027, -0.0001294284, 0.02009537, 0.006000501,
  0.01724306, 0.02241955, 0.01726653, 0.02389773, 0.03284139, 0.01153149, 
    0.009173066, 0.1810004, 0.3226717, 0.1068981, 0.1022808, 0.149341, 
    0.1363407, 0.03379802, 0.002812983, 0.03184489, 0.02761255, 0.01436313, 
    2.443572e-05, 8.803095e-07, 0.01155652, 0.01337754, 0.02165311, 
    0.05730437, 0.05889632, 0.02252681, 0.01371757, 2.337342e-05, 0.0006339037,
  0.06829014, 0.03832566, 0.06282698, 0.09683277, 0.06312686, 0.06189199, 
    0.1155683, 0.06129131, 0.0573955, 0.1140089, 0.1112738, 0.08695267, 
    0.1430015, 0.1928653, 0.1211756, 0.1307145, 0.08743896, 0.1097833, 
    0.04499052, 0.07007258, 0.1539564, 0.1052452, 0.09040841, 0.1368376, 
    0.1733131, 0.1127998, 0.08774999, 0.06116759, 0.07901993,
  0.1132372, 0.104714, 0.1094106, 0.1033014, 0.1102386, 0.1111827, 0.1082228, 
    0.1583098, 0.1841713, 0.1365894, 0.2471866, 0.1961295, 0.1659352, 
    0.1011535, 0.1569365, 0.169504, 0.2283682, 0.1720097, 0.1366985, 
    0.1107343, 0.1229259, 0.1280847, 0.1009032, 0.1898379, 0.1976682, 
    0.1248148, 0.1074154, 0.1277328, 0.1541498,
  0.1211351, 0.1397921, 0.07231463, 0.1789788, 0.177765, 0.2186488, 
    0.2280026, 0.2341927, 0.2291057, 0.2029724, 0.1964781, 0.1889322, 
    0.1857248, 0.2805448, 0.1560174, 0.1275676, 0.2118295, 0.2769764, 
    0.2141718, 0.1643153, 0.1593425, 0.1978051, 0.1015114, 0.1475829, 
    0.1686561, 0.2369264, 0.1433546, 0.1831737, 0.1068321,
  0.1829485, 0.1185308, 0.10218, 0.09615314, 0.1096707, 0.1865377, 0.1972036, 
    0.2003736, 0.1590724, 0.2121976, 0.1557691, 0.1798522, 0.1592267, 
    0.1479307, 0.09321235, 0.1426715, 0.09265608, 0.1589438, 0.1581734, 
    0.1282973, 0.10767, 0.1033051, 0.1297171, 0.1204584, 0.1033155, 
    0.2010688, 0.1362475, 0.2186284, 0.1739152,
  0.06194233, 0.07873435, 0.1313688, 0.1759599, 0.1630021, 0.1421383, 
    0.08647881, 0.1048809, 0.1168215, 0.09805055, 0.1014984, 0.1267218, 
    0.1567647, 0.18249, 0.1774251, 0.1638361, 0.1508572, 0.1641408, 
    0.0920864, 0.07277111, 0.08091252, 0.102354, 0.0964558, 0.05303152, 
    0.06389637, 0.07481822, 0.1115744, 0.06739566, 0.08927189,
  0.004230002, 0.002867249, 0.001504497, 0.0001417447, -0.001221008, 
    -0.00258376, -0.003946512, -0.001343762, -0.0005570342, 0.0002296934, 
    0.001016421, 0.001803149, 0.002589876, 0.003376604, 0.003793053, 
    0.005028098, 0.006263143, 0.007498189, 0.008733234, 0.009968279, 
    0.01120332, 0.005385799, 0.004726779, 0.004067758, 0.003408738, 
    0.002749717, 0.002090696, 0.001431676, 0.005320204,
  0.03142602, 0.01095541, 0.0008659515, 0, 0, 0, 0, 0, 0, 0, -3.884251e-07, 
    0.0004651452, 0.02622327, 0.19685, 0.1553226, 0.1720049, 0.2179136, 
    0.2094412, 0.1594434, 0.1210286, 0.1634025, 0.1790543, 0.3581836, 
    0.3941707, 0.319911, 0.2190632, 0.1533986, 0.1392674, 0.05624439,
  0.1990715, 0.2560518, 0.3483913, 0.2882801, 0.05144458, 0.03940358, 
    0.2093809, 0.05265058, 0.06683214, 0.1592014, 0.1349352, 0.1497375, 
    0.1927363, 0.1652677, 0.2382192, 0.2139451, 0.2185247, 0.2501839, 
    0.3117875, 0.2958906, 0.4334219, 0.3342757, 0.3384317, 0.3686987, 
    0.3366917, 0.2360073, 0.2189599, 0.2666523, 0.2910756,
  0.2327767, 0.2236247, 0.2452262, 0.2686123, 0.3112789, 0.2518973, 0.2406, 
    0.248604, 0.2846162, 0.3007126, 0.3129351, 0.3089986, 0.3246629, 
    0.2775015, 0.1962135, 0.2104469, 0.2377211, 0.2237935, 0.3069664, 
    0.291227, 0.2874702, 0.2318996, 0.2529128, 0.2582335, 0.2430423, 
    0.2495876, 0.2250076, 0.2247528, 0.1917977,
  0.2198438, 0.2005266, 0.1934708, 0.1977012, 0.1638543, 0.1757765, 
    0.1525478, 0.1637854, 0.2216964, 0.2116995, 0.2540183, 0.2290653, 
    0.1393129, 0.1084878, 0.09895633, 0.09294038, 0.1184207, 0.1098115, 
    0.1527266, 0.1524304, 0.2000425, 0.1879915, 0.2104133, 0.180337, 
    0.1447944, 0.1788197, 0.1676601, 0.1842587, 0.2180152,
  0.1341986, 0.0684288, 0.09125923, 0.09072568, 0.09305908, 0.05801483, 
    0.0775474, 0.05702636, 0.05863332, 0.09147216, 0.0935894, 0.07989328, 
    0.08327859, 0.06580766, 0.1133977, 0.1409691, 0.1057601, 0.09266159, 
    0.1242092, 0.1609597, 0.119527, 0.1594926, 0.09403171, 0.1469555, 
    0.07217491, 0.08186784, 0.1095878, 0.1244339, 0.151098,
  0.005413592, 0.001301282, 0.00549577, 0.0384367, 0.04908489, 0.04308266, 
    0.01680125, 0.008840236, 0.0647966, 0.03210104, 0.02989426, 0.01472305, 
    0.03596507, 0.05142388, 0.09061201, 0.1436592, 0.1127076, 0.1063397, 
    0.1308469, 0.08266141, 0.07438301, 0.06124403, 0.01633799, 0.02878932, 
    0.0286851, 0.04299476, 0.04160802, 0.05051782, 0.02825719,
  -3.700422e-06, 2.8247e-05, 0.01100211, 0.001901256, 0.0643646, 0.07021437, 
    0.01509332, 0.009744673, 0.05841091, 0.007766676, 0.04184884, 
    0.0009893976, 0.02163487, 0.1314826, 0.03805987, 0.006906379, 0.03639828, 
    0.02874878, 0.02046958, 0.001660803, 0.0004666382, -1.159539e-06, 
    -3.175855e-07, 1.578467e-05, 0.03486857, 0.001237841, 0.01479134, 
    0.001842003, 2.952863e-07,
  0.0008911518, 0.02003944, 0.004051568, 0.07429896, 0.08481891, 0.06002451, 
    0.07882051, 0.07218786, 0.07725001, 0.05280338, 0.08050971, 0.02929998, 
    0.1458784, 0.04851585, 0.02561457, 0.01775866, 0.02045553, 0.02293963, 
    0.02676248, 0.01468924, 0.0004211195, -1.248948e-06, 0.005046248, 
    0.04985212, 0.005906126, 0.002627216, 0.0198509, 0.0002051201, 
    0.0007440593,
  0.04998916, 0.2369868, 0.219861, 0.02099367, 0.01249319, 0.07994705, 
    0.04966506, 0.01391812, 0.09518694, 0.1675826, 0.0863104, 0.03547345, 
    0.01882102, 0.01254849, 0.03598404, 0.01911863, 0.01704968, 0.0164922, 
    0.01707401, 0.02245234, 0.01877642, 0.01585288, 0.07265939, 0.2548578, 
    0.1399077, 0.1213851, 0.08504983, 0.03361971, 0.03373134,
  0.04487265, 0.05203471, 0.03243079, 0.1675358, 0.004263878, 0.004634834, 
    0.01532732, 0.07535621, 0.06713695, 0.07823213, 0.1446914, 0.04186814, 
    0.1283483, 0.1243007, 0.163446, 0.1549478, 0.0556185, 0.02492951, 
    0.06449393, 0.04841705, 0.02180058, 0.09140851, 0.1121209, 0.1032209, 
    0.01175335, 0.01955378, 0.01205327, 0.01880724, 0.1165246,
  0.004619641, 0.006983843, 0.002001359, 0.004471296, 0.02472027, 
    2.538969e-06, 0.002253709, 0.0144355, 0.1271659, 0.2001456, 0.05513991, 
    0.03004823, 0.06910967, 0.004997849, 0.005295989, 0.03715483, 0.01692487, 
    0.01859122, 0.0007296444, 0.000724073, 0.0006098803, 0.01881891, 
    0.03310779, 0.1633265, 0.01789109, 0.01009678, -0.0002638836, 0.00521831, 
    0.002272351,
  0.009256422, 0.0124355, 0.005475228, 0.01229308, 0.04110677, 0.005600166, 
    0.001474368, 0.1674026, 0.2995818, 0.1122044, 0.1143405, 0.1568131, 
    0.1428663, 0.03737119, 0.005776297, 0.03055809, 0.03380048, 0.01550592, 
    -8.432551e-07, 4.383914e-06, 0.003582774, 0.01187974, 0.02082954, 
    0.05691436, 0.06289373, 0.02335479, 0.0167229, 8.963742e-05, 0.0005421813,
  0.06371468, 0.03300344, 0.06320485, 0.08998182, 0.06805372, 0.04712857, 
    0.1189533, 0.04697148, 0.03348263, 0.1048634, 0.1124095, 0.07997606, 
    0.1401476, 0.1818486, 0.1266708, 0.1303383, 0.09971158, 0.1115017, 
    0.04143988, 0.0683658, 0.1374649, 0.09457015, 0.0856682, 0.136722, 
    0.1732767, 0.109798, 0.08926166, 0.06127353, 0.08742836,
  0.1283265, 0.108019, 0.1133273, 0.1001662, 0.1147121, 0.1241492, 0.1201046, 
    0.1605225, 0.1845826, 0.1219761, 0.225302, 0.1942385, 0.1689906, 
    0.1035318, 0.1509749, 0.1621037, 0.2405451, 0.1914911, 0.1399124, 
    0.1197083, 0.1247503, 0.1260979, 0.1066162, 0.2183035, 0.2155932, 
    0.1403075, 0.1290186, 0.1365064, 0.1539725,
  0.1132095, 0.1438583, 0.08329646, 0.1855241, 0.2050386, 0.2216501, 
    0.2195514, 0.2471401, 0.2316465, 0.1999976, 0.1948542, 0.196028, 
    0.1849215, 0.2672128, 0.1524558, 0.1603025, 0.2256548, 0.3006641, 
    0.2065778, 0.1718892, 0.1694078, 0.1969913, 0.1257757, 0.1648817, 
    0.1780867, 0.2427835, 0.1475468, 0.1644975, 0.09675471,
  0.177134, 0.1152235, 0.1299935, 0.1044853, 0.1159865, 0.182154, 0.1997522, 
    0.2037087, 0.1572632, 0.2088669, 0.1574315, 0.1545755, 0.1500218, 
    0.1247666, 0.0815192, 0.1352833, 0.0976107, 0.156996, 0.1516946, 
    0.1470352, 0.1060979, 0.1042794, 0.1225808, 0.136824, 0.1060172, 
    0.2211247, 0.1683879, 0.2118627, 0.1744148,
  0.05917882, 0.0868201, 0.126195, 0.1800769, 0.1588779, 0.1459468, 
    0.08705056, 0.1014915, 0.1210765, 0.1060596, 0.117242, 0.1242844, 
    0.1653087, 0.1950055, 0.1815883, 0.1729419, 0.1816755, 0.1723624, 
    0.08239314, 0.06749887, 0.07280389, 0.1029157, 0.1090276, 0.05367895, 
    0.06749973, 0.07033747, 0.1010141, 0.07182793, 0.08942987,
  0.06572561, 0.05981055, 0.05389548, 0.04798042, 0.04206536, 0.03615029, 
    0.03023523, 0.03598479, 0.03719855, 0.03841231, 0.03962608, 0.04083984, 
    0.0420536, 0.04326737, 0.03548228, 0.04152265, 0.04756302, 0.0536034, 
    0.05964378, 0.06568415, 0.07172453, 0.1000932, 0.09875412, 0.09741504, 
    0.09607597, 0.09473689, 0.09339782, 0.09205874, 0.07045767,
  0.0436606, 0.02214793, 0.002353843, -3.367959e-05, 0, 0, 0, 0, 0, 0, 
    0.004096909, 0.0149184, 0.04253996, 0.2329344, 0.1602621, 0.1880937, 
    0.2228167, 0.2256079, 0.2278727, 0.1978418, 0.279196, 0.3185133, 
    0.399758, 0.4058975, 0.3156697, 0.2117778, 0.1574415, 0.1328637, 0.0975958,
  0.1898288, 0.2593458, 0.3474382, 0.2816035, 0.1088319, 0.05175987, 
    0.2479191, 0.1159111, 0.1532771, 0.2506883, 0.2235948, 0.2384036, 
    0.1918022, 0.1767632, 0.2403624, 0.2132183, 0.2375415, 0.2766654, 
    0.3426173, 0.3038521, 0.4209725, 0.3335153, 0.3409488, 0.3732019, 
    0.3486392, 0.2374865, 0.2008104, 0.2624596, 0.3003038,
  0.2583494, 0.2573953, 0.2454711, 0.2768168, 0.3168347, 0.2526786, 
    0.2818611, 0.2554681, 0.3159486, 0.2679435, 0.3062223, 0.2956095, 
    0.3068845, 0.2959664, 0.1990569, 0.207087, 0.2292368, 0.2220043, 
    0.285355, 0.2840708, 0.2990121, 0.2430963, 0.2526584, 0.2387195, 
    0.2268544, 0.2526885, 0.2410733, 0.2406399, 0.2112512,
  0.2430473, 0.2037869, 0.2139814, 0.1965252, 0.1743349, 0.1730547, 
    0.1528508, 0.1879334, 0.2319504, 0.2219568, 0.25972, 0.2340174, 
    0.1355943, 0.1018867, 0.09519842, 0.08807936, 0.1229258, 0.1248826, 
    0.1675164, 0.1638525, 0.193267, 0.1713371, 0.1919254, 0.1766189, 0.1364, 
    0.1720037, 0.161769, 0.1935004, 0.2087648,
  0.1386333, 0.07910579, 0.08896445, 0.1037906, 0.09902801, 0.06075897, 
    0.08248261, 0.05919609, 0.06840142, 0.08014773, 0.09218551, 0.08940673, 
    0.09338111, 0.06482621, 0.1112107, 0.1419703, 0.1131629, 0.0951336, 
    0.1153221, 0.1463974, 0.1219873, 0.1595535, 0.1030688, 0.1446086, 
    0.07918029, 0.09296374, 0.1116457, 0.1298182, 0.1742313,
  0.008206678, 0.001178781, 0.008441969, 0.03748263, 0.04466426, 0.05016441, 
    0.01511766, 0.01388121, 0.06705409, 0.04235655, 0.02222021, 0.01158328, 
    0.04929937, 0.05443085, 0.09789264, 0.1471318, 0.1131324, 0.1088176, 
    0.1285745, 0.1094806, 0.08403382, 0.06411319, 0.02090685, 0.0189869, 
    0.03580868, 0.04032668, 0.0450416, 0.05037761, 0.03271952,
  1.845972e-07, 5.406846e-05, 0.01818946, 0.005991194, 0.07853891, 
    0.07813718, 0.0170977, 0.009701504, 0.05494488, 0.01142315, 0.03419981, 
    0.0001140146, 0.02388539, 0.1236425, 0.03206826, 0.006541506, 0.03972236, 
    0.03309684, 0.0309936, 0.005486303, 0.001170079, -3.478351e-06, 
    1.08284e-07, 1.934939e-05, 0.04780629, 0.001931689, 0.01901341, 
    0.004642066, 3.244181e-07,
  0.00122491, 0.01644779, 0.006322719, 0.07844169, 0.08537854, 0.0625904, 
    0.07518516, 0.07620562, 0.07050335, 0.039582, 0.07505849, 0.02475862, 
    0.1430135, 0.04225968, 0.02302807, 0.01748398, 0.01923504, 0.02372296, 
    0.02647852, 0.0107076, 0.001637338, 1.799131e-05, 0.002503529, 
    0.05909895, 0.007080282, 0.004950821, 0.02490257, 5.604921e-05, 
    8.782527e-05,
  0.03310848, 0.2638064, 0.2411829, 0.02706906, 0.011759, 0.06226876, 
    0.03760039, 0.01067849, 0.09872727, 0.1872353, 0.06428427, 0.02604393, 
    0.01760571, 0.01050989, 0.0335725, 0.0172951, 0.01737597, 0.01487468, 
    0.01091003, 0.01476606, 0.01068925, 0.00946291, 0.05566707, 0.2647652, 
    0.1678616, 0.1166805, 0.09302963, 0.02795499, 0.0186469,
  0.03824555, 0.03413826, 0.02829494, 0.1747459, 0.007295368, 0.003997361, 
    0.01113191, 0.04426127, 0.04737665, 0.05173706, 0.1279035, 0.03178802, 
    0.09391309, 0.1023787, 0.1403337, 0.1219213, 0.05963466, 0.02948894, 
    0.04663802, 0.04014508, 0.01869248, 0.0748914, 0.1159662, 0.1083734, 
    0.01017387, 0.01842453, 0.009638262, 0.009818978, 0.1179318,
  0.002323444, 0.002799733, 0.0001731563, 0.001071534, 0.008605635, 
    4.652255e-06, 0.002547414, 0.006440082, 0.1502077, 0.1645008, 0.05284272, 
    0.02323487, 0.05843607, 0.005433276, 0.008635765, 0.03196658, 0.01798473, 
    0.0126589, 0.0003851327, 0.0007142274, 1.965483e-05, 0.02161084, 
    0.02994851, 0.141343, 0.02319349, 0.00732253, -0.0001951961, 
    5.841933e-05, 0.0004857857,
  0.003300357, 0.003616557, 0.002984935, 0.008085577, 0.04356356, 
    0.002193162, -0.0001102499, 0.1503057, 0.3052925, 0.109096, 0.1192541, 
    0.1453823, 0.1404091, 0.03530839, 0.01089675, 0.02884619, 0.03820888, 
    0.014653, -1.249138e-05, 2.886085e-06, 0.0008916973, 0.01010585, 
    0.02074955, 0.05904614, 0.07308441, 0.02810437, 0.01969507, 0.003182095, 
    3.725707e-05,
  0.0668259, 0.03481656, 0.0611446, 0.09084563, 0.06979096, 0.03268464, 
    0.1191662, 0.0360905, 0.02152364, 0.08531304, 0.112969, 0.07487933, 
    0.1407362, 0.175059, 0.1311512, 0.139108, 0.1048116, 0.1210968, 
    0.04593414, 0.07315842, 0.1142374, 0.08772765, 0.09216645, 0.1397429, 
    0.177276, 0.1153429, 0.09830311, 0.06661068, 0.08898084,
  0.1333247, 0.1013167, 0.1184989, 0.09593613, 0.1140975, 0.1221382, 
    0.1188657, 0.1706148, 0.1755663, 0.1115174, 0.2170991, 0.1982163, 
    0.1661834, 0.0995737, 0.1508158, 0.1753244, 0.2469194, 0.1926921, 
    0.1252692, 0.129513, 0.126398, 0.1372126, 0.1333427, 0.230068, 0.2313869, 
    0.151844, 0.1342228, 0.1322085, 0.1597383,
  0.1131917, 0.149497, 0.09950498, 0.1913572, 0.1985007, 0.2255912, 
    0.2229035, 0.2582865, 0.232109, 0.2098707, 0.1989006, 0.1949489, 
    0.1868142, 0.2887364, 0.1406623, 0.2116556, 0.2400833, 0.3254974, 
    0.2214585, 0.1797745, 0.1774691, 0.2118591, 0.1227196, 0.1813613, 
    0.1764133, 0.248735, 0.1576585, 0.1846303, 0.1060358,
  0.1816796, 0.1141624, 0.1496017, 0.1034861, 0.1262657, 0.1660863, 
    0.1943297, 0.2016688, 0.1610095, 0.2138234, 0.1530399, 0.147818, 
    0.1347611, 0.107522, 0.07314051, 0.1326401, 0.107703, 0.1594963, 
    0.1461745, 0.1439022, 0.1211398, 0.1010042, 0.1199584, 0.1378045, 
    0.1281893, 0.2351094, 0.1680214, 0.1986909, 0.1759388,
  0.06310795, 0.08198303, 0.1287955, 0.1833242, 0.1632617, 0.1503275, 
    0.1031175, 0.1204839, 0.1402202, 0.1386996, 0.1482078, 0.1468632, 
    0.1845204, 0.1989316, 0.1886532, 0.1993354, 0.215725, 0.1749407, 
    0.08492997, 0.06224028, 0.07064615, 0.1135318, 0.1143962, 0.06200384, 
    0.06538338, 0.07003875, 0.09802215, 0.1027048, 0.100368,
  0.1359361, 0.1318708, 0.1278054, 0.1237401, 0.1196747, 0.1156094, 0.111544, 
    0.1078686, 0.1087525, 0.1096364, 0.1105203, 0.1114043, 0.1122882, 
    0.1131721, 0.1053518, 0.1105959, 0.1158399, 0.121084, 0.1263281, 
    0.1315722, 0.1368163, 0.1555406, 0.1534779, 0.1514153, 0.1493526, 
    0.1472899, 0.1452273, 0.1431646, 0.1391884,
  0.07189687, 0.03782665, 0.01496918, -4.53254e-05, 0, -1.188653e-05, 
    -4.59965e-05, 0, 7.44241e-05, 0.009674239, 0.02296196, 0.0440363, 
    0.0986148, 0.2499039, 0.1640401, 0.1820634, 0.2126874, 0.2024539, 
    0.2304769, 0.2515954, 0.3428336, 0.4294159, 0.4421365, 0.41052, 0.328613, 
    0.218581, 0.1725458, 0.1365626, 0.1280428,
  0.2199726, 0.2756709, 0.3390658, 0.3042094, 0.1629285, 0.06101842, 
    0.2338894, 0.2005055, 0.244453, 0.3116538, 0.2789276, 0.2727072, 
    0.1990348, 0.1912619, 0.281255, 0.228277, 0.2639596, 0.297958, 0.3729036, 
    0.3513744, 0.4174449, 0.3553227, 0.3468001, 0.4249246, 0.3516116, 
    0.2317734, 0.2850351, 0.2810656, 0.3137059,
  0.2642743, 0.2960206, 0.2670361, 0.2984355, 0.299738, 0.2597443, 0.268216, 
    0.2770608, 0.3286772, 0.309657, 0.319982, 0.2812456, 0.2738119, 0.268755, 
    0.1970074, 0.2277088, 0.2365715, 0.2361248, 0.298505, 0.3173967, 
    0.3106625, 0.2519997, 0.260165, 0.2385058, 0.2494024, 0.2707533, 
    0.2223155, 0.2475112, 0.2548068,
  0.256797, 0.228831, 0.2241202, 0.1981096, 0.1848683, 0.1741973, 0.1534939, 
    0.1970746, 0.2359926, 0.2343642, 0.2485335, 0.2303771, 0.1393178, 
    0.1154003, 0.1022667, 0.09620818, 0.1307216, 0.1193212, 0.1696917, 
    0.1789641, 0.2061929, 0.1709235, 0.175085, 0.1745863, 0.1266335, 
    0.1676815, 0.1614361, 0.1971664, 0.2230101,
  0.1481444, 0.08763586, 0.08956071, 0.1110736, 0.1090677, 0.07052454, 
    0.09228881, 0.05766003, 0.08009854, 0.0884548, 0.1035645, 0.09260482, 
    0.09734272, 0.07006647, 0.1353517, 0.1394577, 0.1145243, 0.106068, 
    0.1208723, 0.1425759, 0.1301413, 0.1597068, 0.1102282, 0.1461639, 
    0.08669832, 0.09728426, 0.1182517, 0.1312366, 0.1682296,
  0.01010988, 0.002372826, 0.01992293, 0.03175661, 0.04917569, 0.06330656, 
    0.01735501, 0.01935216, 0.06392627, 0.04433045, 0.02034192, 0.01329938, 
    0.05928215, 0.0613963, 0.1042239, 0.15675, 0.1261895, 0.1152318, 
    0.123991, 0.1229183, 0.09354463, 0.0723999, 0.02908125, 0.01169969, 
    0.04609432, 0.04435177, 0.05330447, 0.05665076, 0.03682309,
  1.882536e-07, 4.065042e-05, 0.03027965, 0.01490012, 0.09658799, 0.07952201, 
    0.03888667, 0.009964317, 0.04342232, 0.007723869, 0.03103696, 
    1.917858e-05, 0.02429124, 0.1150847, 0.02828144, 0.01292352, 0.04754779, 
    0.03726571, 0.04065485, 0.01232413, 0.002404994, -2.289426e-05, 
    -8.009501e-07, 1.944853e-05, 0.04441857, 0.003213514, 0.02903058, 
    0.006457723, 6.178431e-07,
  0.001778149, 0.01683294, 0.01204307, 0.08482544, 0.08276677, 0.05761711, 
    0.07202071, 0.07696055, 0.06480586, 0.03747316, 0.0658821, 0.02389602, 
    0.1432223, 0.03673296, 0.02341846, 0.01924447, 0.01982393, 0.02495856, 
    0.02428592, 0.008709713, 0.002064739, 0.0002054136, 0.0004933528, 
    0.05306634, 0.007980289, 0.006118203, 0.03493823, 7.719497e-05, 
    1.192353e-06,
  0.01603461, 0.1853428, 0.186951, 0.03736353, 0.01075726, 0.05112112, 
    0.0352665, 0.008977399, 0.08742512, 0.1686716, 0.05506057, 0.02207394, 
    0.01645446, 0.01040561, 0.030906, 0.01816437, 0.01737412, 0.01409986, 
    0.009255506, 0.01150667, 0.0141144, 0.00476955, 0.05234104, 0.2425241, 
    0.160665, 0.1078718, 0.09931543, 0.02679297, 0.0105623,
  0.02386468, 0.01623515, 0.01765732, 0.1666928, 0.006135951, 0.00337528, 
    0.007163989, 0.01237497, 0.03760972, 0.03718273, 0.1095762, 0.02461177, 
    0.07528456, 0.09495509, 0.1258639, 0.09977584, 0.06081492, 0.02683933, 
    0.03744135, 0.03450634, 0.01090489, 0.06507934, 0.1129022, 0.08035008, 
    0.0111389, 0.01899904, 0.008681634, 0.003515359, 0.06203979,
  6.741587e-06, 0.0007759502, 9.229252e-06, 1.784644e-05, 0.0007143979, 
    6.034985e-06, 0.001237043, 0.004091586, 0.1315197, 0.14194, 0.05244282, 
    0.01838768, 0.05085126, 0.009749774, 0.01426328, 0.03056967, 0.01862034, 
    0.01052585, 0.0001101165, 6.884558e-05, 5.010725e-06, 0.02284454, 
    0.02342998, 0.09062371, 0.01893928, 0.006464486, 6.637964e-05, 
    1.100819e-05, 0.0004323737,
  0.0006739138, 0.001816544, 0.002033798, 0.008063621, 0.03757434, 
    0.0007474663, -0.0008188308, 0.109442, 0.3191345, 0.09267497, 0.1076458, 
    0.1337336, 0.138833, 0.04119041, 0.01842612, 0.03577173, 0.0586372, 
    0.01694161, -2.157129e-05, 2.027963e-06, 0.0001207932, 0.009589653, 
    0.02164285, 0.06288727, 0.08479343, 0.02948771, 0.02405755, 0.003415584, 
    5.441244e-05,
  0.06395328, 0.03778345, 0.06708182, 0.09840729, 0.06923448, 0.02868619, 
    0.117984, 0.03102896, 0.01200707, 0.07089006, 0.1138914, 0.08185202, 
    0.1450023, 0.1810591, 0.1382813, 0.1438438, 0.1141287, 0.1297015, 
    0.04533983, 0.08321899, 0.1072747, 0.08736114, 0.119413, 0.1484854, 
    0.1820386, 0.1177442, 0.1128742, 0.07905765, 0.09424029,
  0.1253869, 0.1083597, 0.1177568, 0.1097001, 0.13696, 0.1268228, 0.1258869, 
    0.1820767, 0.1607025, 0.1103818, 0.2280808, 0.2070757, 0.184889, 
    0.102437, 0.1525317, 0.2064289, 0.2380563, 0.2082859, 0.1431173, 
    0.1347991, 0.1354241, 0.1251755, 0.1571314, 0.2669472, 0.2254962, 
    0.1497482, 0.1187404, 0.1411736, 0.1749511,
  0.120141, 0.1727039, 0.1058024, 0.2130907, 0.2284594, 0.2484306, 0.2238455, 
    0.271119, 0.2414633, 0.2379669, 0.2499404, 0.2378335, 0.1770358, 
    0.2854428, 0.2012057, 0.2563615, 0.2548354, 0.3701916, 0.2737221, 0.1857, 
    0.1751403, 0.2065097, 0.1103811, 0.1974796, 0.1783809, 0.2339433, 
    0.163533, 0.1710679, 0.1112369,
  0.1922964, 0.1275938, 0.1490835, 0.1175277, 0.1309146, 0.1794949, 
    0.1824105, 0.2007383, 0.1723242, 0.2450103, 0.1583296, 0.1464485, 
    0.1280215, 0.1035287, 0.07259297, 0.1447004, 0.1525038, 0.1637398, 
    0.1200238, 0.1520161, 0.1397328, 0.1326278, 0.1353112, 0.1456446, 
    0.09642549, 0.2673782, 0.1647736, 0.1866155, 0.1891844,
  0.09074096, 0.1342686, 0.1618451, 0.1856012, 0.1744635, 0.1759849, 
    0.1424347, 0.1604055, 0.1907421, 0.1735719, 0.1748532, 0.1867345, 
    0.2461377, 0.2369416, 0.2106977, 0.1866719, 0.2204916, 0.1534927, 
    0.09787276, 0.05952841, 0.08153126, 0.1390397, 0.1408622, 0.07799758, 
    0.09263597, 0.07799697, 0.1108747, 0.1336042, 0.1299473,
  0.1962645, 0.1933652, 0.190466, 0.1875667, 0.1846674, 0.1817682, 0.1788689, 
    0.1820375, 0.1838476, 0.1856577, 0.1874678, 0.1892779, 0.191088, 
    0.1928981, 0.1798722, 0.1850745, 0.1902769, 0.1954793, 0.2006817, 
    0.2058841, 0.2110865, 0.2184877, 0.2143745, 0.2102612, 0.206148, 
    0.2020348, 0.1979216, 0.1938083, 0.1985839,
  0.1115852, 0.04744579, 0.0417692, 0.002957344, -6.539147e-05, 
    -1.154467e-05, -0.0007750007, -0.0004998766, 0.010074, 0.02724497, 
    0.0383468, 0.117197, 0.1474262, 0.2644911, 0.1593934, 0.1630869, 
    0.1713648, 0.1892504, 0.2166235, 0.2498091, 0.3980239, 0.5272629, 
    0.4612612, 0.4132044, 0.3050309, 0.2052878, 0.1678158, 0.1435291, 
    0.1480346,
  0.1993278, 0.2652215, 0.3634049, 0.3176698, 0.1929783, 0.07748894, 
    0.2424291, 0.2686095, 0.2797357, 0.356903, 0.3518107, 0.2798096, 
    0.1954316, 0.1780936, 0.2979337, 0.2486345, 0.2890971, 0.3116155, 
    0.3624731, 0.3364178, 0.3707075, 0.4021704, 0.3795768, 0.4509201, 
    0.3528187, 0.2368357, 0.2582472, 0.2555401, 0.3096227,
  0.2594282, 0.2982405, 0.2906772, 0.3039551, 0.2977101, 0.2845965, 
    0.2954087, 0.3129117, 0.357611, 0.3373135, 0.3675162, 0.2826971, 
    0.2915546, 0.2924908, 0.2170146, 0.2343144, 0.2420374, 0.2707619, 
    0.3508324, 0.3371339, 0.3346137, 0.2849966, 0.2754092, 0.2939281, 
    0.3001323, 0.3228556, 0.2763693, 0.2425735, 0.2434536,
  0.2632818, 0.2382236, 0.2333573, 0.2089973, 0.1945833, 0.1839269, 
    0.1582564, 0.2341396, 0.2479774, 0.2502541, 0.261056, 0.2330913, 
    0.1514134, 0.1210509, 0.1087613, 0.1177225, 0.1421085, 0.1436529, 
    0.1813935, 0.1984635, 0.2209206, 0.1793292, 0.1754396, 0.1754619, 
    0.1163317, 0.1668806, 0.1718817, 0.2067969, 0.2395289,
  0.1751709, 0.09320115, 0.09721012, 0.1139751, 0.1309525, 0.086309, 
    0.1123953, 0.08321275, 0.09953517, 0.1070944, 0.1082912, 0.1062414, 
    0.112457, 0.1001199, 0.1636509, 0.1523028, 0.1146734, 0.1186686, 
    0.1265524, 0.1521038, 0.1361223, 0.1778418, 0.1286106, 0.1500074, 
    0.09925506, 0.1088987, 0.1333466, 0.1396986, 0.1726048,
  0.01728458, 0.00363392, 0.06617348, 0.0273096, 0.04860796, 0.07094968, 
    0.02187944, 0.02490497, 0.06422353, 0.03888042, 0.00833222, 0.01841089, 
    0.07168265, 0.06148662, 0.1136742, 0.1666485, 0.1447329, 0.1244538, 
    0.1310647, 0.1140018, 0.09396619, 0.07458717, 0.03497674, 0.009699358, 
    0.05654509, 0.0541289, 0.05963688, 0.06324083, 0.04550353,
  5.947126e-07, 0.007162381, 0.03334911, 0.01726227, 0.1136577, 0.08807684, 
    0.04988485, 0.01513552, 0.0389946, 0.00169983, 0.01306057, 0.0004440042, 
    0.02583359, 0.1078391, 0.02732238, 0.02250783, 0.04485699, 0.04349447, 
    0.06240236, 0.03830107, 0.01372257, 0.0007640306, -0.000108134, 
    1.102699e-05, 0.04901625, 0.004267707, 0.03708768, 0.01193858, 
    9.086954e-05,
  0.003625157, 0.02596592, 0.01513308, 0.09442816, 0.08004176, 0.0563008, 
    0.06622197, 0.07693964, 0.07390195, 0.03634543, 0.07020189, 0.03034448, 
    0.1428589, 0.03982259, 0.02602556, 0.02239681, 0.02598127, 0.02870841, 
    0.01802941, 0.01021922, 0.000859727, 1.929282e-06, 7.223536e-05, 
    0.05609839, 0.01259798, 0.04663759, 0.05258046, 0.000308778, 3.739792e-07,
  0.009889469, 0.151402, 0.1665273, 0.04966827, 0.009201623, 0.0498374, 
    0.03247013, 0.009344406, 0.08826771, 0.1633494, 0.05340168, 0.02098909, 
    0.01698934, 0.01335268, 0.03719096, 0.02188025, 0.01739007, 0.01475301, 
    0.009518119, 0.005745417, 0.008363528, 0.002628662, 0.03765043, 
    0.2361507, 0.1649285, 0.09616436, 0.1017161, 0.02825643, 0.009692546,
  0.01693724, 0.008167331, 0.01208969, 0.1410955, 0.01099484, 0.00329867, 
    0.004918316, 0.00707901, 0.03121249, 0.03056839, 0.09609032, 0.02308628, 
    0.06646039, 0.09393692, 0.1156204, 0.08570436, 0.07057732, 0.03007216, 
    0.04104822, 0.03526847, 0.01065136, 0.0572623, 0.1123218, 0.06833367, 
    0.01510066, 0.02015886, 0.009813365, 0.0009690913, 0.04333215,
  2.96627e-06, 0.0001339607, 2.672091e-06, -1.196819e-05, 8.67605e-05, 
    4.818268e-06, 0.0006561354, 0.00241371, 0.1259125, 0.1410307, 0.05412088, 
    0.01665184, 0.04500087, 0.01669468, 0.02816225, 0.03438091, 0.02568947, 
    0.01454358, 1.846625e-05, 7.7885e-06, 2.682493e-06, 0.02566536, 
    0.02157337, 0.06810618, 0.02202973, 0.01336545, 0.001472512, 
    3.907488e-06, -2.899001e-05,
  2.951492e-05, 0.0006928386, 0.001037092, 0.003251225, 0.02559444, 
    0.000132749, -0.0007089342, 0.0722838, 0.3138472, 0.08925644, 0.0961131, 
    0.1405347, 0.1336336, 0.04715722, 0.02500615, 0.04091962, 0.07659284, 
    0.0229268, 0.002663711, 2.305814e-06, 0.0003369198, 0.01654033, 
    0.02038612, 0.05470964, 0.08234049, 0.02969605, 0.02345621, 0.003110833, 
    0.001160708,
  0.0568528, 0.04196354, 0.07459483, 0.1133727, 0.06827548, 0.02017269, 
    0.1157631, 0.02288847, 0.005244507, 0.05673474, 0.1213192, 0.09042954, 
    0.1469492, 0.1908183, 0.1377899, 0.1502412, 0.1249552, 0.1298367, 
    0.05855138, 0.09612826, 0.09650487, 0.08696458, 0.1503783, 0.1564827, 
    0.1867441, 0.1287408, 0.125003, 0.1022325, 0.1102786,
  0.1486244, 0.1146098, 0.1388146, 0.1209728, 0.1350376, 0.1392207, 
    0.1289965, 0.2011289, 0.1458068, 0.1114661, 0.2462942, 0.2337006, 
    0.2028549, 0.1161566, 0.151096, 0.2152607, 0.2542684, 0.2202921, 
    0.1376088, 0.1411848, 0.1257104, 0.1212373, 0.1514827, 0.283202, 
    0.2412478, 0.1912505, 0.1333393, 0.1456853, 0.1975151,
  0.1552686, 0.2240079, 0.1672772, 0.2342992, 0.2586102, 0.2908748, 
    0.2502863, 0.2894327, 0.2734696, 0.2792358, 0.322604, 0.2702112, 
    0.174025, 0.3179716, 0.2484211, 0.3440259, 0.3352399, 0.4040547, 
    0.2643767, 0.1993687, 0.1685861, 0.2357504, 0.1252421, 0.2211435, 
    0.2010066, 0.2268585, 0.1741023, 0.1952683, 0.1456903,
  0.2472602, 0.1437318, 0.1911857, 0.1228359, 0.1661474, 0.2144619, 
    0.1707553, 0.1891457, 0.1842394, 0.2873424, 0.2128831, 0.1854776, 
    0.1446096, 0.1146344, 0.0938274, 0.2091474, 0.194889, 0.1736594, 
    0.1264036, 0.1585632, 0.1541165, 0.141484, 0.1492553, 0.156043, 
    0.1348794, 0.2861634, 0.1714253, 0.1635822, 0.2432742,
  0.1224733, 0.1527926, 0.1424735, 0.1896822, 0.1738542, 0.1791872, 0.152513, 
    0.1681544, 0.209016, 0.2365278, 0.1941612, 0.1811451, 0.2672428, 
    0.2901689, 0.2782412, 0.2397122, 0.2203676, 0.1508005, 0.08861633, 
    0.0615793, 0.1096232, 0.1440036, 0.1393749, 0.1059738, 0.1146402, 
    0.08538945, 0.1268241, 0.175872, 0.1714005,
  0.2259708, 0.2242051, 0.2224393, 0.2206737, 0.218908, 0.2171422, 0.2153765, 
    0.2254842, 0.2279491, 0.230414, 0.232879, 0.2353439, 0.2378088, 
    0.2402737, 0.2235445, 0.2315668, 0.239589, 0.2476112, 0.2556334, 
    0.2636557, 0.2716779, 0.2997056, 0.2909842, 0.2822627, 0.2735412, 
    0.2648198, 0.2560983, 0.2473769, 0.2273833,
  0.12984, 0.07503171, 0.05628926, 0.01508932, 0.004746191, 0.0006605799, 
    0.005707429, 0.01272894, 0.01559494, 0.0328312, 0.08828212, 0.132546, 
    0.1888553, 0.2584682, 0.107243, 0.128102, 0.1608912, 0.1601499, 
    0.1839708, 0.2341401, 0.425161, 0.5820104, 0.4808364, 0.4019754, 
    0.2674259, 0.1744868, 0.1508418, 0.160127, 0.1497009,
  0.1791263, 0.2521143, 0.3326881, 0.3040444, 0.2137899, 0.08853081, 
    0.2586436, 0.2910402, 0.3323717, 0.3932332, 0.3875007, 0.2791491, 
    0.1772753, 0.187025, 0.292883, 0.2701001, 0.2413646, 0.2652479, 
    0.3172379, 0.2715402, 0.3582346, 0.3376886, 0.335619, 0.433136, 
    0.3280893, 0.215755, 0.2065772, 0.2068002, 0.3233219,
  0.2738732, 0.2882005, 0.2941148, 0.2949238, 0.2765698, 0.2916687, 
    0.2895531, 0.2851551, 0.3555679, 0.3457502, 0.3510929, 0.3029307, 
    0.2783095, 0.2945981, 0.2415748, 0.2645686, 0.2672922, 0.2924598, 
    0.3766162, 0.3522442, 0.3247793, 0.2843174, 0.2879471, 0.2754183, 
    0.2831998, 0.2884744, 0.2606109, 0.2473814, 0.2640342,
  0.2604384, 0.2340078, 0.2437032, 0.2126952, 0.2021292, 0.2065791, 
    0.1876095, 0.2492343, 0.2624526, 0.2711208, 0.278777, 0.2484102, 
    0.1723825, 0.1197241, 0.153204, 0.1334436, 0.1644128, 0.182481, 0.225071, 
    0.2134182, 0.2442057, 0.1760101, 0.2050158, 0.1879386, 0.113798, 
    0.1785971, 0.1752283, 0.2260617, 0.2549147,
  0.1975204, 0.1083957, 0.1132452, 0.1162853, 0.1568835, 0.09663975, 
    0.1164653, 0.1049642, 0.1318709, 0.1422801, 0.1328098, 0.1208983, 
    0.1241325, 0.1099502, 0.1948919, 0.1867084, 0.1366832, 0.1269096, 
    0.1421673, 0.1659127, 0.1571997, 0.1785539, 0.1536749, 0.1591095, 
    0.1218934, 0.1266719, 0.1466886, 0.1572703, 0.187442,
  0.0276621, 0.00728789, 0.05719937, 0.03610712, 0.04882285, 0.07478698, 
    0.02917353, 0.03739069, 0.07104781, 0.0355235, 0.005433739, 0.007450803, 
    0.07645866, 0.06864993, 0.1105329, 0.1562407, 0.1301401, 0.1398201, 
    0.1408017, 0.1141963, 0.09755015, 0.09247583, 0.04127581, 0.009242764, 
    0.07105644, 0.06330486, 0.06658865, 0.0679937, 0.05184519,
  2.035262e-06, 0.0003807879, 0.05417228, 0.02245061, 0.1176683, 0.102609, 
    0.05920117, 0.03017643, 0.03950949, 0.001394284, 0.005220056, 
    0.0005164176, 0.02529697, 0.1033516, 0.02660649, 0.032501, 0.04647373, 
    0.04955352, 0.06976195, 0.06735092, 0.03549863, 0.01265104, 0.004544248, 
    5.892502e-06, 0.05350197, 0.007802249, 0.04650421, 0.03046868, 0.003104865,
  0.001704255, 0.02965737, 0.01736956, 0.101154, 0.07715721, 0.05667589, 
    0.06351615, 0.08097161, 0.08332521, 0.04028587, 0.08325864, 0.04209556, 
    0.1536365, 0.04199702, 0.0292857, 0.02691039, 0.03026262, 0.03323307, 
    0.01872033, 0.01107057, 0.0005020349, 9.677806e-05, 6.060042e-06, 
    0.05791686, 0.01821298, 0.1248221, 0.07953915, 0.0009377948, 7.29316e-07,
  0.008793825, 0.1359823, 0.1416281, 0.07583898, 0.007783527, 0.04724173, 
    0.03084822, 0.01046773, 0.09724977, 0.172764, 0.04812717, 0.02112015, 
    0.01749132, 0.01554951, 0.03797266, 0.02648583, 0.02080108, 0.01855426, 
    0.01527848, 0.006058794, 0.003332344, 0.001488602, 0.02733566, 0.2449441, 
    0.163901, 0.08472803, 0.1007162, 0.03502683, 0.01081788,
  0.0123872, 0.005134309, 0.005411816, 0.105506, 0.007852947, 0.003218165, 
    0.004981498, 0.006359485, 0.02503353, 0.0252767, 0.08493029, 0.02495809, 
    0.05943868, 0.0877941, 0.1011136, 0.0823051, 0.07263552, 0.03644585, 
    0.054751, 0.04049091, 0.01412879, 0.05520061, 0.1138628, 0.06788477, 
    0.01987555, 0.02214378, 0.01265543, 0.0002407761, 0.03170309,
  1.430675e-06, 1.368507e-05, 1.362787e-06, -9.429282e-06, 1.45978e-05, 
    3.069298e-06, 0.0002532325, 0.0008879333, 0.1461151, 0.1372585, 
    0.05287756, 0.01748656, 0.0457158, 0.02718567, 0.03346977, 0.03729862, 
    0.02879447, 0.01856824, 7.85412e-06, 3.121568e-06, 1.111349e-06, 
    0.02940963, 0.02366944, 0.05565792, 0.0232526, 0.02398462, 0.005998613, 
    1.737724e-06, -5.673165e-07,
  2.684986e-06, 0.0004031745, 0.0002914751, 0.003145456, 0.01643068, 
    1.174039e-05, -0.0005127934, 0.05050778, 0.2944826, 0.09403872, 
    0.08615258, 0.1373597, 0.1372886, 0.05398812, 0.028699, 0.03904259, 
    0.08462389, 0.02319116, 0.002643753, 1.250326e-05, -4.163563e-06, 
    0.01253492, 0.01621744, 0.06142328, 0.09365951, 0.02906973, 0.02474809, 
    0.006203974, 0.002922692,
  0.0446559, 0.03408159, 0.07760318, 0.1270597, 0.03653535, 0.007347913, 
    0.1052781, 0.01806113, 0.002323457, 0.046596, 0.1288294, 0.08810918, 
    0.149061, 0.1891453, 0.1374271, 0.1458647, 0.1255304, 0.1367202, 
    0.07397632, 0.1068541, 0.07924715, 0.08332693, 0.1753083, 0.1455291, 
    0.1872405, 0.1378971, 0.1288013, 0.1113278, 0.1304666,
  0.1799352, 0.1283534, 0.1496084, 0.1461624, 0.1105146, 0.1128773, 
    0.1089447, 0.2149355, 0.1305323, 0.1070961, 0.2382697, 0.2648622, 
    0.2046665, 0.120002, 0.1606075, 0.2210982, 0.2652382, 0.2323978, 
    0.1477069, 0.1514494, 0.1156554, 0.09887699, 0.1681358, 0.3034424, 
    0.2294902, 0.2075252, 0.179832, 0.1622134, 0.2197834,
  0.2137544, 0.2691747, 0.195283, 0.2574696, 0.2938146, 0.3185051, 0.2600594, 
    0.2734485, 0.2521198, 0.2790407, 0.3119013, 0.2866902, 0.1896453, 
    0.3321643, 0.2076784, 0.2966473, 0.3740581, 0.4130673, 0.2420491, 
    0.2035509, 0.1508849, 0.2168059, 0.1324704, 0.2143905, 0.160724, 
    0.2081408, 0.1806738, 0.2295529, 0.2173755,
  0.2331191, 0.1481878, 0.2095201, 0.1461437, 0.1520866, 0.2088403, 
    0.1733959, 0.1909272, 0.2121332, 0.2819601, 0.2153199, 0.1909332, 
    0.1028032, 0.1385741, 0.08494452, 0.1539701, 0.1630242, 0.1475845, 
    0.1464478, 0.1686212, 0.1439987, 0.13298, 0.168345, 0.200449, 0.1244741, 
    0.2974606, 0.1687573, 0.1383276, 0.2421342,
  0.09776148, 0.1256928, 0.1485206, 0.1437949, 0.1173408, 0.1385437, 
    0.1289453, 0.1309311, 0.1737698, 0.1557058, 0.1484117, 0.1611666, 
    0.2300446, 0.2546947, 0.1701456, 0.1913578, 0.1693095, 0.1080872, 
    0.05367651, 0.06139779, 0.09681235, 0.1650744, 0.1604827, 0.1497047, 
    0.1505133, 0.1038332, 0.13224, 0.1736139, 0.1648958,
  0.2770053, 0.2761574, 0.2753096, 0.2744618, 0.273614, 0.2727662, 0.2719183, 
    0.2932001, 0.2991897, 0.3051793, 0.311169, 0.3171586, 0.3231482, 
    0.3291378, 0.3190279, 0.3254445, 0.331861, 0.3382775, 0.344694, 
    0.3511106, 0.3575271, 0.3509845, 0.3394262, 0.3278678, 0.3163095, 
    0.3047512, 0.2931929, 0.2816345, 0.2776836,
  0.1438477, 0.1168844, 0.06975776, 0.04554823, 0.007694853, 0.01006032, 
    0.01144549, 0.01684831, 0.01853047, 0.05623386, 0.1431179, 0.1563847, 
    0.2077501, 0.2302064, 0.1771487, 0.1578804, 0.1623338, 0.1648134, 
    0.1628945, 0.2378272, 0.4751809, 0.6154671, 0.4753808, 0.365766, 
    0.2794907, 0.1676157, 0.1471592, 0.169692, 0.1628861,
  0.2121533, 0.2510179, 0.2953836, 0.306083, 0.2340574, 0.09835997, 
    0.2636034, 0.3244305, 0.3815091, 0.408085, 0.4152149, 0.2805778, 
    0.1709858, 0.2178568, 0.3120364, 0.2931889, 0.2499276, 0.2717166, 
    0.3167315, 0.2409956, 0.3377338, 0.3021457, 0.3096271, 0.4108259, 
    0.3008711, 0.2069297, 0.2267315, 0.2161614, 0.3231961,
  0.2922839, 0.2908428, 0.2925196, 0.2869889, 0.2801016, 0.2905238, 
    0.2621083, 0.3036816, 0.3421097, 0.338962, 0.314231, 0.3156224, 
    0.2933347, 0.3079734, 0.271993, 0.2688741, 0.2755435, 0.2915845, 
    0.3531387, 0.3469748, 0.3317966, 0.2893437, 0.2901541, 0.2522008, 
    0.2554367, 0.2480843, 0.2285898, 0.2182977, 0.2695228,
  0.2459928, 0.2674642, 0.2459926, 0.2218109, 0.2119396, 0.2138451, 
    0.2079717, 0.2792442, 0.27448, 0.2773516, 0.2967541, 0.2652087, 
    0.1768573, 0.1303907, 0.1912009, 0.1536017, 0.1995149, 0.20992, 
    0.2603381, 0.2225363, 0.2595172, 0.1927813, 0.2019192, 0.1963195, 
    0.1263275, 0.2056043, 0.1792059, 0.2385761, 0.2412237,
  0.2138578, 0.1214943, 0.1230762, 0.1206641, 0.1725377, 0.107628, 0.1185565, 
    0.1127886, 0.1683283, 0.1871959, 0.167938, 0.1302341, 0.1271603, 
    0.1255192, 0.1721172, 0.2171201, 0.1552038, 0.1558934, 0.168058, 
    0.1769575, 0.1714004, 0.1844315, 0.1668997, 0.17508, 0.1335822, 
    0.1524467, 0.1616095, 0.188402, 0.197694,
  0.04599378, 0.01150916, 0.03476778, 0.0491659, 0.05272247, 0.08936845, 
    0.03980618, 0.05897503, 0.1012863, 0.0465446, 0.01666086, 0.003461328, 
    0.05345234, 0.07540802, 0.1064477, 0.1404211, 0.1281662, 0.1477053, 
    0.1597794, 0.106674, 0.09243743, 0.09788249, 0.05386029, 0.01070411, 
    0.06890644, 0.07147948, 0.08457762, 0.0817655, 0.05639587,
  -1.187838e-05, -2.660403e-05, 0.0566796, 0.02388495, 0.1014664, 0.0896218, 
    0.05747379, 0.04225949, 0.04314895, 0.01742191, 0.0009383807, 
    0.002570196, 0.03101748, 0.09299652, 0.02413865, 0.03994576, 0.04629407, 
    0.05387219, 0.06876377, 0.064787, 0.05210441, 0.04974219, 0.005579168, 
    2.161598e-05, 0.0612871, 0.01431883, 0.05015367, 0.0519859, 0.02959092,
  6.826406e-05, 0.02479009, 0.0191216, 0.1045498, 0.07003354, 0.05828189, 
    0.06138289, 0.0830943, 0.0837786, 0.05072014, 0.108307, 0.05952192, 
    0.1621222, 0.04004472, 0.03027596, 0.02641299, 0.02711796, 0.03411593, 
    0.02210605, 0.01228875, 0.001985092, 0.001261553, 1.434169e-06, 
    0.05748276, 0.02179369, 0.08035061, 0.08596303, 0.00278859, 1.514693e-05,
  0.01327745, 0.122223, 0.1201757, 0.08269271, 0.008803335, 0.04529358, 
    0.02817055, 0.0116671, 0.1016043, 0.1778418, 0.04399167, 0.02030255, 
    0.01710334, 0.01632585, 0.03470735, 0.02586515, 0.02516934, 0.02224447, 
    0.01874881, 0.01068335, 0.003104134, 0.003070996, 0.01703313, 0.2510242, 
    0.1625384, 0.0718774, 0.09525412, 0.0425585, 0.01180647,
  0.009745003, 0.003588913, 0.002100454, 0.07161526, 0.006344882, 
    0.004066777, 0.01173681, 0.00695375, 0.02164438, 0.02195878, 0.07161459, 
    0.02439059, 0.05588617, 0.07843129, 0.08864387, 0.07958621, 0.078938, 
    0.04421278, 0.07077511, 0.04100329, 0.01711513, 0.05188164, 0.1178376, 
    0.07643038, 0.02414402, 0.02556715, 0.01601493, -1.477583e-05, 0.02171495,
  7.349893e-07, 8.998538e-07, 9.250876e-07, -5.683178e-06, 2.076589e-06, 
    1.524584e-06, 7.703452e-05, 0.0001207739, 0.1521417, 0.147837, 
    0.05021019, 0.02238284, 0.04307541, 0.03296172, 0.03993204, 0.03315533, 
    0.03319416, 0.03808801, 0.0002035248, 1.673493e-06, 9.029993e-07, 
    0.03727808, 0.02580708, 0.04668446, 0.02040434, 0.02808516, 0.01459066, 
    -5.550951e-06, 3.306039e-07,
  -1.826457e-05, 9.104107e-05, 1.677562e-05, 0.00181849, 0.007649081, 
    3.450604e-06, -0.0003553045, 0.03423596, 0.2790563, 0.106596, 0.07842317, 
    0.1539837, 0.1310595, 0.05904222, 0.03407995, 0.05574527, 0.09011775, 
    0.03630018, 0.003083458, 0.000182851, -4.491242e-06, 0.01356705, 
    0.01756977, 0.05769157, 0.1078009, 0.0327751, 0.0302741, 0.00718522, 
    0.004874684,
  0.03492361, 0.02877826, 0.07025127, 0.1366529, 0.01611779, 0.004193014, 
    0.1010223, 0.01482866, 0.003831476, 0.03697105, 0.12788, 0.08614558, 
    0.1621474, 0.1875843, 0.146708, 0.1483836, 0.1319868, 0.1520126, 
    0.07161679, 0.1041648, 0.07088228, 0.08530038, 0.1716645, 0.143806, 
    0.1729608, 0.1317462, 0.1156217, 0.1249181, 0.1322106,
  0.1773265, 0.1364717, 0.1624144, 0.1620456, 0.06482575, 0.08461502, 
    0.08735292, 0.2120411, 0.1080343, 0.09240149, 0.2290097, 0.2818586, 
    0.2056192, 0.1177542, 0.1551885, 0.2119619, 0.2688003, 0.2432151, 
    0.148765, 0.1745486, 0.1024806, 0.08028617, 0.1823149, 0.3225889, 
    0.2323366, 0.2049474, 0.2298704, 0.1991931, 0.2313372,
  0.2149365, 0.2839115, 0.154104, 0.2843093, 0.2840427, 0.2963117, 0.2634024, 
    0.250289, 0.231531, 0.2821481, 0.2485368, 0.3014072, 0.190022, 0.2990382, 
    0.2065647, 0.2239114, 0.3501805, 0.4303951, 0.2306862, 0.1761538, 
    0.1478227, 0.1799398, 0.1313984, 0.1942593, 0.1367981, 0.1934764, 
    0.1753108, 0.2433035, 0.2279245,
  0.2235727, 0.1792168, 0.2250103, 0.2049688, 0.1254141, 0.1719735, 
    0.2323035, 0.2194069, 0.2139928, 0.2122918, 0.1686254, 0.1743977, 
    0.07807278, 0.09874361, 0.06629872, 0.08619963, 0.1036586, 0.1108948, 
    0.1331509, 0.1322982, 0.1725039, 0.1457355, 0.1610582, 0.1832464, 
    0.1118545, 0.3136006, 0.1671352, 0.1270406, 0.1912124,
  0.06817689, 0.06891356, 0.1019941, 0.1033546, 0.09302896, 0.1456605, 
    0.1176855, 0.111932, 0.1322099, 0.1182209, 0.1269037, 0.1211736, 
    0.1723026, 0.1992604, 0.1165151, 0.1430813, 0.1492599, 0.06841089, 
    0.05086159, 0.0581663, 0.08029602, 0.1668836, 0.1700979, 0.1116252, 
    0.1199793, 0.1262426, 0.1639706, 0.1888337, 0.175515,
  0.3025506, 0.3013915, 0.3002325, 0.2990735, 0.2979144, 0.2967554, 
    0.2955964, 0.3117726, 0.3200956, 0.3284187, 0.3367417, 0.3450648, 
    0.3533878, 0.3617108, 0.3674465, 0.3735814, 0.3797163, 0.3858511, 
    0.391986, 0.3981209, 0.4042557, 0.3989966, 0.3856977, 0.3723988, 
    0.3590999, 0.345801, 0.3325021, 0.3192032, 0.3034778,
  0.1535209, 0.1742658, 0.08341175, 0.07075365, 0.01263932, 0.03320207, 
    0.03347347, 0.03364523, 0.03486944, 0.08543412, 0.1671085, 0.1786588, 
    0.2525329, 0.2036541, 0.1965069, 0.1778733, 0.1796962, 0.1593739, 
    0.1560298, 0.2243377, 0.5180898, 0.6279365, 0.4722584, 0.3478956, 
    0.2538938, 0.1731175, 0.1658931, 0.1619767, 0.1624776,
  0.2127236, 0.2736658, 0.2956337, 0.272526, 0.2486499, 0.1163927, 0.2425735, 
    0.3492854, 0.4172835, 0.4201741, 0.4279332, 0.2807233, 0.1731205, 
    0.2199446, 0.3073354, 0.3024274, 0.2459001, 0.3026696, 0.3245597, 
    0.2847402, 0.3521271, 0.3207855, 0.3472444, 0.4325285, 0.2782924, 
    0.2157511, 0.2030912, 0.229324, 0.3195395,
  0.3737319, 0.3591658, 0.3515649, 0.3109627, 0.2918615, 0.3174306, 
    0.3271149, 0.3547166, 0.3782665, 0.3586899, 0.3181272, 0.3646518, 
    0.3341119, 0.3580295, 0.2957038, 0.3126181, 0.3218675, 0.3296468, 
    0.3605502, 0.36591, 0.3430405, 0.313068, 0.3256264, 0.2700782, 0.2848535, 
    0.2627026, 0.2237662, 0.242058, 0.3288796,
  0.2601272, 0.2950532, 0.2771167, 0.2458887, 0.245068, 0.2313849, 0.2492502, 
    0.3159884, 0.2988727, 0.3082166, 0.3282966, 0.2867448, 0.2066395, 
    0.1687884, 0.191533, 0.1748893, 0.2505355, 0.2609761, 0.3179325, 
    0.2641214, 0.2704461, 0.2047922, 0.2156447, 0.2104486, 0.164882, 
    0.2430646, 0.2175332, 0.2783317, 0.2613997,
  0.2265431, 0.1447571, 0.1339438, 0.1341213, 0.1684897, 0.1187632, 
    0.1403054, 0.1398357, 0.2131201, 0.2152727, 0.1788467, 0.1413759, 
    0.1559363, 0.1458606, 0.2001992, 0.2135209, 0.1773736, 0.188993, 
    0.1985514, 0.1954775, 0.1725871, 0.2002115, 0.1717956, 0.1947493, 
    0.1313502, 0.1738363, 0.1871804, 0.2030374, 0.2102083,
  0.08853032, 0.02218634, 0.02219514, 0.05999291, 0.05298747, 0.1002382, 
    0.05422952, 0.08704633, 0.1252305, 0.07767828, 0.01600831, 0.005370596, 
    0.04061969, 0.09815954, 0.09454829, 0.1424138, 0.1432446, 0.1723921, 
    0.1752725, 0.1077007, 0.09076588, 0.1053909, 0.06466077, 0.01102507, 
    0.05331655, 0.09687513, 0.09816077, 0.1114776, 0.09738605,
  0.003916902, -1.656337e-06, 0.01513433, 0.02817432, 0.09329682, 0.0801233, 
    0.05819526, 0.05087344, 0.06324095, 0.04021201, 5.395234e-05, 
    2.468758e-06, 0.05777772, 0.09918278, 0.0282619, 0.06101902, 0.05795704, 
    0.05347407, 0.06689244, 0.04733004, 0.09423913, 0.07561369, 0.02843489, 
    4.495776e-05, 0.08529817, 0.02135795, 0.04428212, 0.06318317, 0.05528867,
  7.949244e-05, 0.02011206, 0.01835075, 0.1107316, 0.06281266, 0.04952503, 
    0.05518489, 0.06909262, 0.07542103, 0.05500444, 0.1098612, 0.06928614, 
    0.1635133, 0.03329422, 0.0276497, 0.02685336, 0.02429893, 0.03112407, 
    0.02050847, 0.01580289, 0.01096703, 0.007002574, -7.466018e-06, 
    0.05477616, 0.02458017, 0.01664105, 0.08306246, 0.0120383, 0.0009216096,
  0.02021592, 0.1149304, 0.09788676, 0.07186849, 0.01092675, 0.03934155, 
    0.02583819, 0.01438964, 0.09575422, 0.1820842, 0.03783482, 0.01852456, 
    0.0167515, 0.01646265, 0.02814503, 0.02423987, 0.02472681, 0.01908361, 
    0.01891307, 0.01214187, 0.00612892, 0.003587003, 0.008559494, 0.255423, 
    0.1590101, 0.05997811, 0.0816901, 0.03426198, 0.01663687,
  0.007663342, 0.002493642, 0.000930725, 0.04573829, 0.00342366, 0.006796619, 
    0.024644, 0.01059571, 0.02114371, 0.02329848, 0.05930733, 0.02670243, 
    0.04737527, 0.06669401, 0.07470252, 0.07166878, 0.08196309, 0.05449403, 
    0.08750023, 0.04283005, 0.02152521, 0.04709348, 0.1144102, 0.08406171, 
    0.03212371, 0.03834757, 0.02305972, 0.0004941156, 0.01580641,
  4.996726e-07, 7.324572e-07, 6.35018e-07, -3.394245e-06, 9.669363e-07, 
    4.949082e-07, 3.299136e-05, -3.239286e-05, 0.1533174, 0.1574079, 
    0.04585357, 0.03304876, 0.03792129, 0.02885292, 0.03421405, 0.03151507, 
    0.03007509, 0.04830059, 0.005092766, 1.552857e-06, 6.143196e-07, 
    0.0438774, 0.02564246, 0.03786258, 0.01959867, 0.03080805, 0.0273755, 
    -2.591788e-05, 2.803061e-07,
  4.217773e-07, 1.998642e-05, 2.921893e-05, 0.001038028, 0.003316686, 
    1.155966e-06, -0.0002396151, 0.02347438, 0.2768011, 0.1052143, 
    0.08155626, 0.1651835, 0.1326566, 0.07208198, 0.04592168, 0.08804326, 
    0.09911006, 0.06312346, 0.02155113, 0.003613481, 7.497393e-06, 
    0.02670154, 0.02010223, 0.07666278, 0.1075097, 0.04750945, 0.03780902, 
    0.02207249, 0.004856003,
  0.02341741, 0.0181106, 0.04979708, 0.1400277, 0.00738913, 0.001515337, 
    0.09776164, 0.008504336, 0.002135755, 0.03133811, 0.1228514, 0.09105752, 
    0.1690328, 0.194716, 0.1616, 0.1927204, 0.173132, 0.1818019, 0.07557975, 
    0.09613833, 0.06730792, 0.09730678, 0.189331, 0.1245768, 0.2062905, 
    0.1498487, 0.132806, 0.1465012, 0.1365287,
  0.1529537, 0.1650804, 0.213441, 0.1629155, 0.03854699, 0.05869397, 
    0.07257526, 0.2127682, 0.09545559, 0.07442676, 0.2265438, 0.2696289, 
    0.2085928, 0.1274069, 0.1832854, 0.2459409, 0.3231786, 0.2695065, 
    0.1692338, 0.1695236, 0.09624325, 0.0832001, 0.18354, 0.3059592, 
    0.2542887, 0.2106485, 0.2606445, 0.2344404, 0.2385471,
  0.2125372, 0.2816765, 0.1601855, 0.2671905, 0.2614617, 0.2548887, 
    0.2366889, 0.2634761, 0.2332796, 0.2716549, 0.2026111, 0.2640696, 
    0.2009431, 0.2790104, 0.229158, 0.2151526, 0.3593035, 0.4407064, 
    0.2373746, 0.1547095, 0.1160233, 0.1569912, 0.1314836, 0.2144777, 
    0.151232, 0.1840814, 0.2712154, 0.278762, 0.2376054,
  0.2856195, 0.1985361, 0.274906, 0.2207989, 0.1882588, 0.178604, 0.1966299, 
    0.2301763, 0.1910614, 0.1968628, 0.1870806, 0.1512777, 0.07070434, 
    0.08195032, 0.05888919, 0.0884237, 0.09476513, 0.09928242, 0.1015722, 
    0.1271674, 0.2005387, 0.1335971, 0.1550767, 0.1447068, 0.1113108, 
    0.3217733, 0.166153, 0.1300122, 0.2162289,
  0.1045602, 0.06458829, 0.1041237, 0.1343806, 0.1026134, 0.1606231, 
    0.1701933, 0.1612847, 0.2046529, 0.1342039, 0.1066526, 0.1709473, 
    0.197338, 0.1971682, 0.1615054, 0.1330318, 0.1375177, 0.1057565, 
    0.07019305, 0.05288886, 0.1285284, 0.1218959, 0.1603106, 0.1107033, 
    0.1165336, 0.1618003, 0.1741261, 0.1993201, 0.1877059,
  0.3362897, 0.3356628, 0.335036, 0.3344091, 0.3337823, 0.3331554, 0.3325286, 
    0.3463939, 0.3563682, 0.3663425, 0.3763168, 0.386291, 0.3962653, 
    0.4062396, 0.4195336, 0.423407, 0.4272803, 0.4311537, 0.435027, 
    0.4389004, 0.4427736, 0.413549, 0.4003283, 0.3871075, 0.3738867, 
    0.360666, 0.3474452, 0.3342244, 0.3367912,
  0.1653518, 0.2117149, 0.126521, 0.08462457, 0.02130192, 0.05801668, 0.0793, 
    0.05488686, 0.04220772, 0.1260584, 0.1809644, 0.2256775, 0.2667392, 
    0.168494, 0.1604874, 0.1817194, 0.1497132, 0.132061, 0.1622501, 
    0.2233225, 0.5614271, 0.6504167, 0.4997382, 0.2904592, 0.2491727, 
    0.1711416, 0.1895262, 0.1540053, 0.1653687,
  0.2021289, 0.3017311, 0.284004, 0.2399973, 0.2491353, 0.1334888, 0.2403716, 
    0.3706887, 0.4168551, 0.4321867, 0.4297124, 0.2724537, 0.1737691, 
    0.2315516, 0.3159154, 0.3230978, 0.264718, 0.333574, 0.4107288, 
    0.3100138, 0.3663964, 0.356085, 0.3686354, 0.470831, 0.2614612, 
    0.2050677, 0.2410031, 0.2520548, 0.3208672,
  0.4359707, 0.3914927, 0.3499933, 0.3191914, 0.3151113, 0.3671514, 
    0.4196478, 0.4420066, 0.4640023, 0.4403768, 0.3417019, 0.3867099, 
    0.389366, 0.4072123, 0.3419009, 0.3468174, 0.3638788, 0.3568336, 
    0.3520116, 0.3565667, 0.3394281, 0.2985206, 0.3665431, 0.3564574, 
    0.341965, 0.3081727, 0.2806045, 0.3192068, 0.4147999,
  0.3235206, 0.2809046, 0.2904833, 0.2792703, 0.2798081, 0.2944011, 
    0.2780232, 0.3478543, 0.3196779, 0.3020557, 0.3256744, 0.3099264, 
    0.2251529, 0.2408386, 0.2205782, 0.2045891, 0.282034, 0.2926368, 
    0.3440151, 0.298926, 0.2658238, 0.2302033, 0.2382713, 0.221697, 
    0.2232586, 0.326534, 0.3222013, 0.3119438, 0.3163546,
  0.2523655, 0.1742315, 0.1329099, 0.1466964, 0.1670532, 0.1500513, 
    0.1908425, 0.2068657, 0.2308703, 0.2013637, 0.1368522, 0.1199823, 
    0.1539685, 0.1680152, 0.2197109, 0.2038638, 0.2018918, 0.2249095, 
    0.229315, 0.2277622, 0.2220354, 0.2342887, 0.1838647, 0.2183696, 
    0.1258552, 0.1921513, 0.2001345, 0.1850633, 0.2063197,
  0.1590021, 0.0489716, 0.01453112, 0.08432746, 0.08199698, 0.09096222, 
    0.1177123, 0.1397312, 0.1624395, 0.09434295, 0.004661882, 0.0005611867, 
    0.02961093, 0.1274144, 0.1030585, 0.1394952, 0.154182, 0.1755033, 
    0.1800688, 0.1389953, 0.1051312, 0.1317683, 0.1014986, 0.01152711, 
    0.06800596, 0.09119227, 0.1240719, 0.1203711, 0.1240218,
  0.09029236, 2.646986e-06, 0.006808193, 0.05234352, 0.09284352, 0.07722756, 
    0.07367908, 0.05815577, 0.06760907, 0.01573145, 1.075369e-05, 
    -9.595559e-07, 0.09494691, 0.1288107, 0.04361446, 0.07972564, 0.08583851, 
    0.05771368, 0.06520708, 0.04929315, 0.09126653, 0.1218811, 0.07387157, 
    0.0003628356, 0.09252874, 0.03497842, 0.0475559, 0.07892481, 0.09406024,
  6.485241e-05, 0.02444771, 0.04071491, 0.1283582, 0.05903935, 0.04269954, 
    0.04852257, 0.06330789, 0.06814975, 0.06160372, 0.113581, 0.07732502, 
    0.1554841, 0.02886932, 0.02833349, 0.02954893, 0.02497707, 0.03136139, 
    0.02294141, 0.02014235, 0.02853226, 0.02995789, 0.0009959325, 0.05518969, 
    0.02554958, 0.005466547, 0.08078101, 0.03088857, 0.01449819,
  0.02899153, 0.109021, 0.07972949, 0.05279934, 0.01504008, 0.03323814, 
    0.02576046, 0.01992821, 0.08381845, 0.1862179, 0.03733977, 0.0181916, 
    0.01887066, 0.01930296, 0.02747887, 0.0253759, 0.02452645, 0.01709181, 
    0.01868472, 0.01552489, 0.01065599, 0.00481593, 0.005448057, 0.2426685, 
    0.1514572, 0.05189002, 0.0690652, 0.03024339, 0.02404036,
  0.006278763, 0.002048181, 0.0003864812, 0.02958175, 0.006800702, 
    0.01502766, 0.0391115, 0.01929042, 0.02120016, 0.02642336, 0.04854019, 
    0.02724361, 0.04111828, 0.05545125, 0.06149893, 0.06457339, 0.07370874, 
    0.07249389, 0.09653783, 0.04747533, 0.02848193, 0.04392055, 0.109678, 
    0.07377233, 0.03470962, 0.05207796, 0.03434032, 0.0008920659, 0.01092697,
  3.574939e-07, 6.593395e-07, 4.328151e-07, -2.475682e-06, 6.53122e-07, 
    2.305456e-07, 6.811752e-06, 0.0006301113, 0.1638021, 0.1474022, 
    0.04234097, 0.04383878, 0.03731784, 0.03225528, 0.03706761, 0.03785021, 
    0.03545204, 0.05621106, 0.03387845, 8.402233e-05, 3.726983e-07, 
    0.04973437, 0.02751369, 0.03212621, 0.02628414, 0.03903222, 0.08772817, 
    0.0005981917, 1.669392e-07,
  1.100558e-06, 6.054787e-06, -1.11444e-05, 0.0006955095, 0.001485973, 
    7.154177e-07, -0.0001635277, 0.01369217, 0.278374, 0.09058234, 
    0.08388871, 0.170736, 0.1644132, 0.09619598, 0.08383967, 0.1141773, 
    0.1311155, 0.1137091, 0.07215474, 0.03232944, 2.901089e-07, 0.0295884, 
    0.02609659, 0.08743177, 0.1169231, 0.06229194, 0.0674509, 0.08277396, 
    0.00589832,
  0.01555125, 0.01161043, 0.02904633, 0.1315761, 0.001604901, 0.0009513355, 
    0.0954596, 0.004838466, 0.0007957704, 0.02672811, 0.1276911, 0.08958116, 
    0.1881398, 0.2275631, 0.2270964, 0.2502074, 0.2688501, 0.3096369, 
    0.1536076, 0.09085795, 0.0594621, 0.1025475, 0.1639402, 0.1186493, 
    0.228218, 0.204801, 0.1658692, 0.1648734, 0.1487887,
  0.1241497, 0.1982812, 0.1664782, 0.1042946, 0.03022227, 0.04960015, 
    0.06082437, 0.202107, 0.07376148, 0.06585976, 0.211579, 0.2855963, 
    0.232794, 0.1334894, 0.2627811, 0.3092992, 0.3625894, 0.3559316, 
    0.2030792, 0.1520489, 0.09162265, 0.07990626, 0.1472896, 0.2944594, 
    0.2569318, 0.2592248, 0.2871308, 0.2718197, 0.2679244,
  0.2228751, 0.2288067, 0.1464995, 0.2606842, 0.2121979, 0.2066267, 
    0.2050165, 0.2219713, 0.2218451, 0.2231638, 0.1922143, 0.2129979, 
    0.2104395, 0.2921191, 0.2517257, 0.2136591, 0.3678934, 0.4216664, 
    0.2415549, 0.1654219, 0.08538993, 0.172427, 0.126214, 0.225783, 
    0.1609506, 0.1988928, 0.3493535, 0.3327849, 0.243146,
  0.3789464, 0.2176984, 0.3069472, 0.2914568, 0.1915256, 0.2309824, 
    0.2620011, 0.1911485, 0.1588878, 0.1535212, 0.1584113, 0.1431368, 
    0.06903698, 0.09880845, 0.03931059, 0.1241881, 0.08448353, 0.1058601, 
    0.09330378, 0.1315082, 0.240758, 0.124993, 0.1648771, 0.1508304, 
    0.1580992, 0.3465635, 0.1560614, 0.1824156, 0.3374754,
  0.1702892, 0.1335386, 0.1136938, 0.139648, 0.1196091, 0.1762217, 0.1773023, 
    0.1980608, 0.2130238, 0.1672751, 0.1333978, 0.1757391, 0.2187107, 
    0.2202811, 0.205553, 0.1904519, 0.1692062, 0.1025396, 0.07123417, 
    0.1007976, 0.1108362, 0.129358, 0.1487314, 0.1406192, 0.1252172, 
    0.1621804, 0.1577565, 0.233146, 0.2507443,
  0.3623399, 0.3620615, 0.3617831, 0.3615047, 0.3612263, 0.3609478, 
    0.3606694, 0.3496498, 0.3594642, 0.3692785, 0.3790928, 0.3889071, 
    0.3987215, 0.4085358, 0.4250911, 0.4279544, 0.4308177, 0.4336809, 
    0.4365441, 0.4394074, 0.4422706, 0.4352508, 0.4228516, 0.4104525, 
    0.3980533, 0.3856542, 0.373255, 0.3608558, 0.3625627,
  0.1810529, 0.2505689, 0.1743746, 0.09480494, 0.0242652, 0.1203957, 
    0.1101033, 0.09409536, 0.04577707, 0.1468216, 0.1953538, 0.2382947, 
    0.2758759, 0.1371466, 0.1489694, 0.1608461, 0.1362694, 0.09762583, 
    0.1441085, 0.2368381, 0.5922039, 0.6787593, 0.5234381, 0.2527782, 
    0.2425988, 0.1801183, 0.1968823, 0.1612372, 0.1771862,
  0.2328368, 0.2823833, 0.2969319, 0.2118889, 0.2588106, 0.1597873, 
    0.2221043, 0.3901331, 0.402122, 0.4410021, 0.4255069, 0.2514833, 
    0.177404, 0.233601, 0.3202543, 0.2977307, 0.315792, 0.4083854, 0.4387991, 
    0.3232592, 0.381012, 0.3815604, 0.3853688, 0.4913224, 0.2503444, 
    0.216653, 0.3345788, 0.302948, 0.333894,
  0.3914198, 0.3678914, 0.3089019, 0.3286017, 0.3351138, 0.3891657, 
    0.5034772, 0.4475719, 0.4330395, 0.4429295, 0.4220954, 0.3750971, 
    0.3977422, 0.4076929, 0.3681312, 0.3794245, 0.3989081, 0.3728327, 
    0.3479087, 0.325515, 0.3198358, 0.2964817, 0.3649921, 0.3750189, 
    0.3860238, 0.3814958, 0.3346981, 0.4057979, 0.4675803,
  0.3140795, 0.2619048, 0.2784237, 0.2921402, 0.3098351, 0.3353259, 0.304971, 
    0.3419878, 0.3039933, 0.2898926, 0.2835149, 0.3275084, 0.2662632, 
    0.2743536, 0.2566068, 0.2576675, 0.2840544, 0.2961862, 0.2952303, 
    0.2848421, 0.2474006, 0.2469964, 0.3043084, 0.2262, 0.2228652, 0.4019587, 
    0.403459, 0.3771179, 0.2914404,
  0.2761429, 0.225657, 0.1285725, 0.1729298, 0.1828249, 0.1698157, 0.222465, 
    0.2652383, 0.2750724, 0.1878829, 0.1392856, 0.1043116, 0.1500365, 
    0.1651212, 0.2484529, 0.1859443, 0.2541191, 0.2706059, 0.2735267, 
    0.2152937, 0.2530886, 0.2678561, 0.2245912, 0.2568258, 0.1117008, 
    0.163122, 0.1731947, 0.1798293, 0.224232,
  0.162755, 0.03775622, 0.01204962, 0.08092186, 0.1057174, 0.09287213, 
    0.1213878, 0.1507301, 0.1931814, 0.09904993, 0.0009394538, 6.210037e-05, 
    0.02355625, 0.08160421, 0.0911324, 0.117678, 0.1371583, 0.1694229, 
    0.1951349, 0.1426022, 0.1272417, 0.1718238, 0.1906083, 0.0119247, 
    0.07872084, 0.08029141, 0.09306988, 0.1041425, 0.1539257,
  0.1548238, -5.234224e-05, 0.002835715, 0.06866328, 0.1007637, 0.08028548, 
    0.06772606, 0.08610471, 0.07355501, 0.008991765, 1.438564e-06, 
    1.154287e-07, 0.07547763, 0.1303483, 0.05342288, 0.08467077, 0.1041347, 
    0.09133597, 0.08107477, 0.06457832, 0.07716817, 0.1632384, 0.2661243, 
    0.0005846971, 0.1230271, 0.05550702, 0.07094898, 0.1047429, 0.1175259,
  0.004889708, 0.02825769, 0.02160628, 0.151388, 0.05792617, 0.05013514, 
    0.05733917, 0.07918007, 0.08271629, 0.07853255, 0.1187033, 0.1094952, 
    0.1503606, 0.03238966, 0.03970498, 0.04460898, 0.0418022, 0.04744793, 
    0.04848146, 0.05646892, 0.05942839, 0.1128206, 0.02100732, 0.06004681, 
    0.03463182, 0.00142967, 0.0887854, 0.0879072, 0.1214772,
  0.04057983, 0.09045475, 0.06145316, 0.0368583, 0.02565672, 0.0379574, 
    0.03908702, 0.03996933, 0.07607619, 0.173022, 0.04073192, 0.02200149, 
    0.02718583, 0.026696, 0.03912052, 0.03417033, 0.02626893, 0.01862625, 
    0.02193794, 0.01680646, 0.01694864, 0.01829131, 0.004708872, 0.2159578, 
    0.1299762, 0.05087827, 0.06223091, 0.03321998, 0.03186603,
  0.004767521, 0.001236169, 0.0001520428, 0.01876737, 0.004785328, 
    0.03508504, 0.05041081, 0.04339053, 0.01510799, 0.04043948, 0.04949981, 
    0.03209525, 0.04027793, 0.05237138, 0.05827358, 0.06286001, 0.06689149, 
    0.09305759, 0.1200553, 0.06240478, 0.04884461, 0.06985121, 0.1064323, 
    0.06838926, 0.03927415, 0.06220839, 0.06736903, 0.002822251, 0.00727672,
  2.853892e-07, 5.867959e-07, 2.822896e-07, -7.54793e-07, 5.116401e-07, 
    1.039812e-07, -3.253429e-06, 0.004537447, 0.1619475, 0.1375445, 
    0.06810857, 0.04962159, 0.05451686, 0.04417955, 0.05033127, 0.06319448, 
    0.0562534, 0.108011, 0.174554, 0.01417597, 2.01759e-07, 0.05328729, 
    0.02873775, 0.03266357, 0.04986039, 0.06392723, 0.1346194, 0.03165057, 
    1.061263e-07,
  5.674372e-07, 3.217098e-06, -0.0001158103, 0.0004215884, 0.0008259129, 
    4.802877e-07, -0.0001234988, 0.006069368, 0.2833455, 0.07305764, 
    0.1166769, 0.211092, 0.2169641, 0.1097806, 0.1684074, 0.199742, 0.199268, 
    0.1746996, 0.2230969, 0.07415006, -9.310689e-05, 0.03596706, 0.03108624, 
    0.1274765, 0.1316195, 0.0886941, 0.09738632, 0.1833013, 0.005167867,
  0.01200847, 0.006488853, 0.0240332, 0.1270851, 0.0008660613, 0.0002497919, 
    0.0994698, 0.005147266, 0.0004340524, 0.02451533, 0.1310928, 0.08816689, 
    0.1891212, 0.2648246, 0.2775527, 0.337289, 0.3406333, 0.4132297, 
    0.2514555, 0.08200379, 0.05538312, 0.1487613, 0.1564898, 0.1198712, 
    0.2516996, 0.2669248, 0.2096283, 0.1874834, 0.1861949,
  0.1211953, 0.1455705, 0.1393929, 0.07668994, 0.03397945, 0.03312592, 
    0.05408777, 0.1883261, 0.06149395, 0.06189102, 0.198456, 0.2909119, 
    0.250509, 0.2200362, 0.3440017, 0.4240794, 0.4464203, 0.3864282, 
    0.2630942, 0.1439284, 0.0840198, 0.06576502, 0.1179811, 0.2768508, 
    0.2625909, 0.3738726, 0.3051845, 0.2472008, 0.2609464,
  0.1885116, 0.1910832, 0.1229549, 0.2280564, 0.1872908, 0.1999227, 0.178091, 
    0.1858961, 0.2039416, 0.1805338, 0.177189, 0.1844177, 0.1964616, 
    0.269646, 0.3488092, 0.3403307, 0.3393773, 0.4195346, 0.2239069, 
    0.1371948, 0.07088464, 0.1696718, 0.1460261, 0.2552113, 0.184644, 
    0.2213863, 0.4650924, 0.407349, 0.2817191,
  0.4600766, 0.2952213, 0.3220631, 0.367368, 0.32617, 0.2530378, 0.2013181, 
    0.1611587, 0.188988, 0.1910695, 0.1271351, 0.1370879, 0.08529525, 
    0.09791821, 0.07909954, 0.1992702, 0.1019965, 0.1272163, 0.08722796, 
    0.1279548, 0.2541797, 0.1727079, 0.2041332, 0.1768872, 0.2639953, 
    0.3860361, 0.1599491, 0.2758216, 0.5197068,
  0.197535, 0.1961311, 0.1553714, 0.1689681, 0.1548965, 0.2282469, 0.2108965, 
    0.231951, 0.2822363, 0.2441784, 0.2623671, 0.2524472, 0.3295755, 
    0.3082457, 0.2591316, 0.2418572, 0.2184328, 0.1377927, 0.1554883, 
    0.1558675, 0.1305378, 0.1400651, 0.1506277, 0.2183537, 0.1785714, 
    0.1825835, 0.1527245, 0.2856535, 0.2832906,
  0.3798408, 0.3795196, 0.3791983, 0.378877, 0.3785558, 0.3782345, 0.3779133, 
    0.3589508, 0.3685895, 0.3782282, 0.387867, 0.3975057, 0.4071445, 
    0.4167832, 0.4300366, 0.4308299, 0.4316232, 0.4324164, 0.4332097, 
    0.4340029, 0.4347962, 0.437171, 0.4270603, 0.4169496, 0.4068388, 
    0.3967281, 0.3866174, 0.3765066, 0.3800978,
  0.2040619, 0.2825764, 0.1987241, 0.1072611, 0.03371281, 0.1604678, 
    0.1426752, 0.1066482, 0.04836977, 0.1486048, 0.2095659, 0.2549365, 
    0.2884701, 0.09152184, 0.1308934, 0.1542603, 0.1459768, 0.08580069, 
    0.1380332, 0.2777025, 0.636893, 0.7029637, 0.5165385, 0.2570741, 
    0.2392237, 0.1962797, 0.2188468, 0.1819362, 0.2287169,
  0.2266801, 0.2585464, 0.2885095, 0.1709921, 0.2497152, 0.1599244, 
    0.1881363, 0.4023437, 0.396526, 0.4406243, 0.4078517, 0.2289501, 
    0.1755593, 0.2301385, 0.3286856, 0.3282795, 0.3826213, 0.4438367, 
    0.3804839, 0.3154149, 0.3940237, 0.4145626, 0.402876, 0.4966351, 
    0.2617747, 0.2392752, 0.3636707, 0.3600864, 0.3240496,
  0.3042472, 0.3030013, 0.2585568, 0.3279122, 0.33293, 0.3442342, 0.46193, 
    0.3758256, 0.3591864, 0.3773775, 0.4053087, 0.357739, 0.4233639, 
    0.3873091, 0.3575493, 0.3773405, 0.3912607, 0.3604647, 0.3431802, 
    0.2919836, 0.332689, 0.3029689, 0.3722863, 0.370328, 0.4571048, 
    0.4636298, 0.3914213, 0.4146654, 0.3799291,
  0.3401344, 0.3099948, 0.3152383, 0.3137268, 0.3348618, 0.3048146, 
    0.3133211, 0.3241002, 0.2902774, 0.2673696, 0.2942773, 0.3350693, 
    0.273589, 0.2470363, 0.2903665, 0.2839313, 0.2727061, 0.3178095, 
    0.2623847, 0.2258847, 0.2261681, 0.2414367, 0.2902979, 0.2390264, 
    0.2068132, 0.3776731, 0.3349453, 0.3562075, 0.3136507,
  0.2787699, 0.2241118, 0.1025158, 0.1678126, 0.1747414, 0.1754702, 
    0.2403629, 0.2238184, 0.2211604, 0.151027, 0.1294731, 0.08893836, 
    0.07870303, 0.1552774, 0.3074418, 0.1711316, 0.2260824, 0.2888275, 
    0.1856032, 0.1807976, 0.1977362, 0.2436438, 0.1919852, 0.2850726, 
    0.1043277, 0.1307718, 0.1542429, 0.1577541, 0.2442098,
  0.207918, 0.05460002, 0.01640501, 0.07716789, 0.07413012, 0.1044244, 
    0.07354444, 0.1425781, 0.163533, 0.03531128, 0.001357174, -8.640588e-06, 
    0.01824489, 0.05183222, 0.08481133, 0.1029387, 0.1081844, 0.1400388, 
    0.1881723, 0.1251115, 0.1401881, 0.1441938, 0.229267, 0.01609038, 
    0.06866805, 0.07196289, 0.0582222, 0.1027887, 0.1085998,
  0.300754, -0.0001135459, 0.002654249, 0.05329287, 0.0887097, 0.06616716, 
    0.06463671, 0.06948734, 0.07107569, 0.02280768, 5.657935e-07, 
    4.829274e-08, 0.04526759, 0.1410969, 0.09373475, 0.08020955, 0.1039982, 
    0.08695713, 0.0956066, 0.05425375, 0.06537104, 0.1061502, 0.3387725, 
    -4.176213e-05, 0.1099671, 0.0485049, 0.1002087, 0.07740262, 0.1503849,
  0.153695, 0.0284344, 0.005045002, 0.1282549, 0.07542907, 0.07778801, 
    0.07380419, 0.08068819, 0.07139063, 0.05281152, 0.07408118, 0.08068836, 
    0.1474463, 0.05020032, 0.04228795, 0.06972712, 0.04590929, 0.05451079, 
    0.0487663, 0.04573834, 0.1012078, 0.21324, 0.2491579, 0.05623967, 
    0.01110391, 0.0003412948, 0.1004939, 0.09302132, 0.2756756,
  0.08795372, 0.0610077, 0.04477797, 0.03714012, 0.2079891, 0.1251216, 
    0.1499722, 0.122418, 0.05092017, 0.1525458, 0.07163309, 0.07052581, 
    0.0449979, 0.1206253, 0.05807041, 0.04706245, 0.04650457, 0.03320278, 
    0.04222581, 0.02579475, 0.03991816, 0.0514629, 0.006769293, 0.1678012, 
    0.0834021, 0.0528133, 0.08477093, 0.1016866, 0.07575449,
  0.002886615, 0.0006756201, 3.566547e-05, 0.01319554, 0.008205894, 
    0.2185903, 0.05885524, 0.1211012, 0.02829746, 0.1556576, 0.07903263, 
    0.0896458, 0.05486159, 0.07000446, 0.06740498, 0.06842485, 0.07424578, 
    0.1316091, 0.1325909, 0.1538793, 0.1834972, 0.09480076, 0.1017939, 
    0.05311028, 0.04690621, 0.1000994, 0.229963, 0.009145275, 0.004068226,
  2.432397e-07, 5.332724e-07, 2.143805e-07, 2.776259e-06, 4.629178e-07, 
    -1.474597e-06, -1.591384e-05, 0.01774743, 0.139314, 0.1527339, 
    0.08665895, 0.06120199, 0.06743886, 0.06377555, 0.05044458, 0.05702233, 
    0.08559398, 0.1059421, 0.3201288, 0.1922459, -1.589371e-06, 0.06592454, 
    0.05408135, 0.04513284, 0.07040302, 0.09464115, 0.1217091, 0.08369658, 
    7.858578e-08,
  6.709521e-08, 2.383837e-06, -0.0001411469, 0.0001371516, 0.000513632, 
    3.639505e-07, -8.82793e-05, 0.003262515, 0.2942212, 0.06789001, 
    0.1325293, 0.2572862, 0.2469603, 0.1719006, 0.2006572, 0.2260167, 
    0.2098432, 0.2392756, 0.3307734, 0.1020378, -0.0001290489, 0.0398988, 
    0.0214014, 0.1358382, 0.1730956, 0.1780815, 0.1871096, 0.2821085, 
    0.01021685,
  0.009951514, 0.004283897, 0.01908925, 0.1312314, 0.007301631, 0.0001397777, 
    0.1047513, 0.005809071, 0.0002588163, 0.02209543, 0.1354905, 0.0763588, 
    0.2116325, 0.3459876, 0.3716905, 0.360629, 0.3612437, 0.4339793, 
    0.304537, 0.07701456, 0.04896237, 0.1555686, 0.1439279, 0.1244561, 
    0.26139, 0.2952208, 0.2254862, 0.2203814, 0.193559,
  0.1171261, 0.1329532, 0.1185306, 0.06590244, 0.02976413, 0.02373808, 
    0.05132895, 0.174213, 0.04829635, 0.05566863, 0.1811071, 0.2964784, 
    0.276609, 0.3499155, 0.3559692, 0.4322359, 0.4493514, 0.3687897, 
    0.2817547, 0.1337777, 0.07368419, 0.05410825, 0.1044114, 0.2707486, 
    0.2535365, 0.4741904, 0.3197492, 0.2698925, 0.2805266,
  0.1470501, 0.141624, 0.1075833, 0.2061044, 0.171673, 0.1811845, 0.1657645, 
    0.1762098, 0.1866087, 0.1609316, 0.1522387, 0.1705514, 0.1839262, 
    0.2432033, 0.4243119, 0.4016638, 0.3244317, 0.418204, 0.2322625, 
    0.1151956, 0.06142962, 0.1660322, 0.2130325, 0.267235, 0.2472418, 
    0.2078512, 0.5523242, 0.4474627, 0.2917944,
  0.4052126, 0.2391044, 0.2705216, 0.2725698, 0.2982529, 0.2496174, 
    0.1362706, 0.1743018, 0.1288242, 0.1355001, 0.1184286, 0.1174465, 
    0.116212, 0.1487089, 0.1595407, 0.3195084, 0.1227641, 0.1249963, 
    0.09641737, 0.1315474, 0.2387611, 0.1851477, 0.2150806, 0.2713867, 
    0.3803972, 0.4005506, 0.1514362, 0.2549102, 0.5534717,
  0.2955596, 0.2059937, 0.2093392, 0.2020268, 0.2528807, 0.2461692, 
    0.2542327, 0.2656008, 0.3234531, 0.3160686, 0.2625702, 0.2568749, 
    0.3503032, 0.4069273, 0.3428665, 0.2745413, 0.2651544, 0.2185709, 
    0.2452708, 0.1616459, 0.1361796, 0.1729668, 0.1644799, 0.277069, 
    0.2184969, 0.2258037, 0.1800567, 0.3276621, 0.2832253,
  0.3730154, 0.372845, 0.3726746, 0.3725042, 0.3723338, 0.3721634, 0.3719929, 
    0.3549257, 0.3643996, 0.3738734, 0.3833473, 0.3928211, 0.402295, 
    0.4117689, 0.4230528, 0.4224039, 0.4217551, 0.4211063, 0.4204574, 
    0.4198086, 0.4191598, 0.4263871, 0.4177325, 0.4090779, 0.4004233, 
    0.3917686, 0.383114, 0.3744594, 0.3731517,
  0.2311891, 0.301556, 0.2280954, 0.1141848, 0.04765359, 0.1688073, 
    0.1629676, 0.1126656, 0.03688885, 0.1409665, 0.2111811, 0.2718334, 
    0.3521349, 0.05264354, 0.1153534, 0.1696465, 0.1909421, 0.1031531, 
    0.1419903, 0.3170437, 0.6633224, 0.7189903, 0.5130656, 0.2653324, 
    0.2269559, 0.2052813, 0.2004249, 0.1997057, 0.2488762,
  0.1930612, 0.1974071, 0.2459425, 0.1362745, 0.2201867, 0.1488863, 
    0.1398872, 0.4032339, 0.3855876, 0.4360341, 0.3977141, 0.2113133, 
    0.1697873, 0.2228418, 0.3220121, 0.3676302, 0.3954241, 0.4091939, 
    0.3184894, 0.307536, 0.4053347, 0.4394558, 0.4128098, 0.508818, 
    0.2829807, 0.2926447, 0.3605841, 0.4371891, 0.3279265,
  0.2638399, 0.254979, 0.2260211, 0.3096826, 0.3412247, 0.3320373, 0.370533, 
    0.2864888, 0.2808525, 0.3059258, 0.3426712, 0.3602332, 0.4250937, 
    0.3963993, 0.3687752, 0.3982102, 0.371233, 0.3502638, 0.32318, 0.2569222, 
    0.3122532, 0.3201427, 0.3737855, 0.3433443, 0.4957082, 0.4954433, 
    0.3973898, 0.3535399, 0.2883936,
  0.3284917, 0.3089097, 0.3532382, 0.3288268, 0.3340808, 0.3191799, 
    0.3262782, 0.3164402, 0.2799503, 0.2478116, 0.2733039, 0.3130749, 
    0.2556817, 0.2796659, 0.2858481, 0.2355313, 0.2603121, 0.2811336, 
    0.2161084, 0.1908888, 0.1862105, 0.2049331, 0.2553115, 0.2569063, 
    0.1919952, 0.3250154, 0.2840593, 0.2960095, 0.3375425,
  0.2312364, 0.1560568, 0.06130946, 0.1298001, 0.1757455, 0.1863265, 
    0.267391, 0.2112139, 0.2040326, 0.1123524, 0.0919247, 0.05612306, 
    0.036228, 0.1326676, 0.3707112, 0.1473341, 0.1536614, 0.1847947, 
    0.1297128, 0.168772, 0.1916417, 0.2165549, 0.175634, 0.3131422, 
    0.07680684, 0.1121372, 0.1289866, 0.124763, 0.2306148,
  0.1164096, 0.07278267, 0.01431877, 0.0392498, 0.03475918, 0.09002496, 
    0.0601499, 0.0620066, 0.1040998, 0.01849917, 0.001079206, -1.95696e-05, 
    0.0158518, 0.02628824, 0.0596591, 0.08587149, 0.1032135, 0.1301109, 
    0.1571654, 0.1053631, 0.1102841, 0.07404044, 0.1088087, 0.01710283, 
    0.0577581, 0.0382335, 0.04024678, 0.05928217, 0.08245976,
  0.1999938, -0.0004601637, 0.003180985, 0.03571893, 0.04110105, 0.04538476, 
    0.02297528, 0.02575861, 0.04505972, 0.004220376, 2.894373e-07, 
    2.624737e-08, 0.01760307, 0.0830187, 0.06740273, 0.08516529, 0.1127127, 
    0.05301594, 0.03985516, 0.01367999, 0.03015605, 0.03762734, 0.1885883, 
    0.01379538, 0.09737369, 0.03698992, 0.02590191, 0.02709172, 0.1575381,
  0.325985, 0.02403264, 0.00135453, 0.08284892, 0.04650853, 0.06092534, 
    0.0392758, 0.04580494, 0.03834186, 0.04573495, 0.04522265, 0.02136524, 
    0.1154307, 0.05709027, 0.02228369, 0.02228079, 0.01928713, 0.02175603, 
    0.01853073, 0.01078347, 0.03097032, 0.07205534, 0.4272352, 0.03263649, 
    0.002115126, 8.309803e-05, 0.03668651, 0.02076061, 0.1052531,
  0.1704859, 0.03707239, 0.03487948, 0.04054663, 0.0575561, 0.03639722, 
    0.0519487, 0.03095623, 0.04054055, 0.1042304, 0.0476632, 0.1284523, 
    0.02000487, 0.02970562, 0.03055224, 0.03372023, 0.04113616, 0.05242693, 
    0.04006233, 0.03861356, 0.06416768, 0.1783877, 0.08398081, 0.1306933, 
    0.05055114, 0.04850129, 0.07760516, 0.1244801, 0.1532952,
  0.001246027, 0.0003929458, -1.714751e-05, 0.007833902, 0.008587605, 
    0.04066445, 0.06643357, 0.02231611, 0.006105795, 0.03167628, 0.05164663, 
    0.03965209, 0.03858393, 0.04755621, 0.04786868, 0.05369198, 0.05170368, 
    0.08047222, 0.08981435, 0.1262704, 0.09436119, 0.06463292, 0.1423444, 
    0.0447414, 0.02043374, 0.03608771, 0.1264029, 0.2097217, 0.001083826,
  2.172901e-07, 4.911602e-07, 1.859795e-07, 2.911748e-05, 4.319431e-07, 
    -0.0004375012, 2.275517e-05, 0.06524246, 0.0985388, 0.1806812, 
    0.09903783, 0.1008984, 0.02714011, 0.01836657, 0.01797365, 0.0239488, 
    0.04364144, 0.03172246, 0.2331413, 0.3769247, 0.005562902, 0.05716251, 
    0.01926751, 0.02955633, 0.05819772, 0.04411821, 0.09073392, 0.0815462, 
    6.709364e-08,
  -2.487266e-07, -6.520115e-06, -3.950026e-05, -1.171165e-06, 0.0005905065, 
    3.008677e-07, -7.218136e-05, 0.002602045, 0.306637, 0.06264273, 
    0.1512048, 0.2459454, 0.3008449, 0.1584116, 0.225942, 0.2112896, 
    0.1832036, 0.1649681, 0.2566249, 0.177543, 0.001125959, 0.03669732, 
    0.01904181, 0.1819319, 0.1858133, 0.1629184, 0.1753842, 0.1622426, 
    0.01164864,
  0.01148669, 0.003990273, 0.01778675, 0.1400304, 0.02452951, -6.987279e-06, 
    0.1050437, 0.004639428, 9.951724e-05, 0.01898391, 0.1381246, 0.08340324, 
    0.2220274, 0.3694928, 0.4326601, 0.370084, 0.3529086, 0.3824839, 
    0.3176866, 0.08258081, 0.04480081, 0.12438, 0.1219364, 0.1325105, 
    0.2392715, 0.2869477, 0.2296469, 0.186594, 0.1866528,
  0.1025036, 0.1146302, 0.1059038, 0.0574754, 0.02695533, 0.02127446, 
    0.04548752, 0.1546868, 0.03673257, 0.05109513, 0.1725818, 0.3008204, 
    0.2971662, 0.3441861, 0.3347303, 0.3801541, 0.4277687, 0.3425698, 
    0.2588744, 0.1338867, 0.0653307, 0.04165341, 0.09121044, 0.2483947, 
    0.2423712, 0.4222372, 0.2996158, 0.2363259, 0.2664132,
  0.1086275, 0.1170722, 0.0940161, 0.1797429, 0.1510832, 0.1655331, 
    0.1518494, 0.1614491, 0.1798465, 0.1517626, 0.1325362, 0.1364681, 
    0.1607595, 0.227098, 0.3773515, 0.4841387, 0.3117784, 0.396991, 
    0.2068862, 0.1035365, 0.06225655, 0.1661563, 0.2059743, 0.293249, 
    0.3155078, 0.194172, 0.4916167, 0.353005, 0.2559473,
  0.2805226, 0.1469658, 0.2005762, 0.1494789, 0.2276229, 0.2162162, 
    0.1159869, 0.1307645, 0.07519541, 0.1113464, 0.1226483, 0.1110979, 
    0.08434124, 0.1585651, 0.2103959, 0.4201249, 0.2018173, 0.1284512, 
    0.1095713, 0.1421271, 0.224871, 0.2079709, 0.1919188, 0.3417934, 
    0.394846, 0.3755098, 0.1576369, 0.1988331, 0.4891531,
  0.3470479, 0.271021, 0.2878663, 0.2441986, 0.3081033, 0.3054601, 0.3084269, 
    0.3284323, 0.3658629, 0.3514266, 0.3235126, 0.3281587, 0.378563, 
    0.4402669, 0.4059241, 0.3159695, 0.332849, 0.2626358, 0.240341, 
    0.2213222, 0.1441397, 0.2136463, 0.183085, 0.2930537, 0.1879374, 
    0.1893575, 0.1781304, 0.3019512, 0.2496251,
  0.3340692, 0.3351592, 0.3362491, 0.3373391, 0.3384291, 0.339519, 0.340609, 
    0.3093495, 0.319352, 0.3293546, 0.3393572, 0.3493598, 0.3593623, 
    0.3693649, 0.4027661, 0.4004191, 0.3980721, 0.3957251, 0.3933781, 
    0.3910311, 0.3886842, 0.382759, 0.3740135, 0.3652679, 0.3565224, 
    0.3477769, 0.3390313, 0.3302858, 0.3331972,
  0.2627349, 0.3079674, 0.2155036, 0.1149828, 0.04114729, 0.1520845, 
    0.1549583, 0.1101031, 0.01963943, 0.1007874, 0.1765297, 0.2552302, 
    0.4046982, 0.02383611, 0.1194876, 0.2181254, 0.2421676, 0.1323698, 
    0.148904, 0.3378007, 0.6690458, 0.7343356, 0.4951044, 0.246162, 
    0.2156939, 0.2203016, 0.2051748, 0.2276311, 0.2607036,
  0.1667297, 0.1416431, 0.2027941, 0.09983222, 0.1861992, 0.1374949, 
    0.09386273, 0.3767676, 0.383365, 0.4302758, 0.3867601, 0.2135496, 
    0.163554, 0.192253, 0.314841, 0.394655, 0.4073116, 0.3865919, 0.2711076, 
    0.3089578, 0.4085333, 0.4703528, 0.4538525, 0.5239679, 0.2834959, 
    0.3259793, 0.4192112, 0.4289521, 0.3135345,
  0.2253702, 0.2223858, 0.2055723, 0.2849768, 0.3173923, 0.309385, 0.2858221, 
    0.2116542, 0.2153833, 0.2436486, 0.2925734, 0.3265886, 0.4119625, 
    0.4169846, 0.3683668, 0.4100313, 0.3534819, 0.3324964, 0.2926229, 
    0.2357949, 0.2673954, 0.2951644, 0.3464898, 0.3031575, 0.4581729, 
    0.5102944, 0.4253587, 0.2847905, 0.2453011,
  0.2969509, 0.3100463, 0.3373066, 0.3264196, 0.3405832, 0.3379547, 
    0.3317357, 0.2988635, 0.2802441, 0.2286423, 0.2458881, 0.2956634, 
    0.2197046, 0.2343351, 0.2605768, 0.2235432, 0.2403529, 0.2441839, 
    0.1814516, 0.169291, 0.161979, 0.1863314, 0.2268174, 0.2482358, 
    0.1619092, 0.2874573, 0.2503356, 0.2592882, 0.3199458,
  0.2136684, 0.1009424, 0.04101109, 0.1003843, 0.150277, 0.1529574, 
    0.2159317, 0.167218, 0.1660982, 0.07781267, 0.0575355, 0.02592826, 
    0.01164141, 0.09579834, 0.3760022, 0.1099985, 0.1143689, 0.1315635, 
    0.1010269, 0.1527276, 0.162028, 0.1891122, 0.1373056, 0.3287169, 
    0.07278661, 0.1179231, 0.1051747, 0.1107347, 0.2252157,
  0.04638365, 0.0377817, 0.01084172, 0.01978261, 0.01677789, 0.05251039, 
    0.02548657, 0.03764819, 0.0551989, 0.009898629, 0.0003372215, 
    -1.931919e-05, 0.01369558, 0.01443354, 0.04740338, 0.06990048, 0.1089224, 
    0.09457122, 0.1235866, 0.1027362, 0.0628216, 0.04213334, 0.05279624, 
    0.02445898, 0.04515398, 0.02245212, 0.0401295, 0.03425995, 0.02717166,
  0.09326653, 0.001891699, 0.002450758, 0.00548801, 0.02121621, 0.02245032, 
    0.006760301, 0.007681002, 0.03683659, 0.0008788565, 2.874519e-06, 
    1.583434e-08, 0.003949803, 0.05189488, 0.03137442, 0.05632719, 
    0.04319393, 0.02235935, 0.01626771, 0.001385631, 0.008515493, 
    0.008925566, 0.06907804, 0.01852216, 0.07336329, 0.03914188, 0.00547659, 
    0.007269457, 0.05724731,
  0.169625, 0.02008847, 0.0004764426, 0.06788631, 0.0152742, 0.01652851, 
    0.01407374, 0.02132487, 0.01007604, 0.006987282, 0.03111051, 0.003041308, 
    0.09380442, 0.01366031, 0.004813104, 0.003988793, 0.003533024, 
    0.01064952, 0.00646951, 0.001586111, 0.007778558, 0.02168303, 0.1813785, 
    0.01535146, 0.0005760876, 2.426769e-05, 0.008039061, 0.004420348, 
    0.03447588,
  0.06318625, 0.02830392, 0.03033051, 0.03601044, 0.009876056, 0.01475722, 
    0.01445327, 0.005937165, 0.04965086, 0.06725009, 0.02381264, 0.02253259, 
    0.002932914, 0.005024309, 0.01346256, 0.005038181, 0.009493677, 
    0.01389607, 0.01008884, 0.01912242, 0.03318408, 0.1038969, 0.4150904, 
    0.1098179, 0.03443381, 0.03236358, 0.04531169, 0.02522554, 0.05925553,
  0.0006031158, 0.0002742112, -1.872424e-05, 0.003988255, 0.01017915, 
    0.01013961, 0.04132213, 0.007951127, 0.00126739, 0.006843484, 0.02492619, 
    0.01460856, 0.01511057, 0.01970076, 0.02382834, 0.02850476, 0.02468325, 
    0.03253243, 0.03761686, 0.03888813, 0.02500747, 0.02298868, 0.1877641, 
    0.03820767, 0.003341276, 0.01171891, 0.03576175, 0.1506656, -0.0001462807,
  1.950206e-07, 4.55306e-07, 1.741589e-07, 0.001578836, 4.102028e-07, 
    0.001091549, -9.628724e-05, 0.05920521, 0.06810133, 0.1629288, 
    0.03486986, 0.02047881, 0.004909382, 0.00270615, 0.005091768, 
    0.007765233, 0.01157655, 0.007625916, 0.1053012, 0.230278, 0.002073157, 
    0.05352626, 0.006073736, 0.01541125, 0.01252643, 0.04109614, 0.02837062, 
    0.02277437, 6.177206e-08,
  4.301637e-08, -4.093354e-05, -2.21931e-05, 9.435344e-06, 0.0006679932, 
    2.683794e-07, -6.754343e-05, 0.002002309, 0.3115065, 0.05591328, 
    0.1369434, 0.2599685, 0.2843179, 0.1688577, 0.2211227, 0.1896366, 
    0.1410972, 0.07235508, 0.1509978, 0.1611702, 0.0009588695, 0.0394106, 
    0.02929407, 0.1291891, 0.1251192, 0.07917552, 0.08210876, 0.06192294, 
    0.01569616,
  0.01116785, 0.002094352, 0.01349082, 0.1417413, 0.03262713, -9.855736e-07, 
    0.1002656, 0.003572582, 5.581311e-05, 0.01552266, 0.1496145, 0.09418302, 
    0.2216578, 0.3585701, 0.39441, 0.3021405, 0.3045806, 0.3465387, 
    0.2534556, 0.0834482, 0.03798599, 0.09791021, 0.1079843, 0.1395483, 
    0.2056976, 0.2577433, 0.1987091, 0.1433101, 0.1598951,
  0.1057804, 0.1002954, 0.08824283, 0.05334679, 0.02178161, 0.02097234, 
    0.03611058, 0.136422, 0.0308971, 0.04460048, 0.1575341, 0.2903131, 
    0.3237509, 0.295884, 0.2887488, 0.3425724, 0.3955859, 0.3155169, 
    0.2082773, 0.1288846, 0.04931153, 0.03138702, 0.08127019, 0.2251427, 
    0.2195086, 0.3816715, 0.2484783, 0.200578, 0.2581798,
  0.09397313, 0.1012561, 0.08300039, 0.1588695, 0.1341315, 0.1487279, 
    0.1344613, 0.134737, 0.1675135, 0.1443722, 0.1181206, 0.1096622, 
    0.1422207, 0.1875652, 0.3011887, 0.5129168, 0.2782457, 0.3783295, 
    0.1791824, 0.09094903, 0.06096104, 0.1350095, 0.1862063, 0.288081, 
    0.4070252, 0.19416, 0.3737712, 0.2854568, 0.2206873,
  0.2386242, 0.09952997, 0.1575676, 0.1005812, 0.1589472, 0.2450584, 
    0.109587, 0.08437596, 0.04015052, 0.08320813, 0.09993691, 0.09188708, 
    0.06495167, 0.140725, 0.1850709, 0.4102504, 0.2261767, 0.1316632, 
    0.1323449, 0.151594, 0.2891768, 0.2470464, 0.1897342, 0.3790484, 
    0.3707055, 0.3308297, 0.1562591, 0.1604372, 0.4112853,
  0.2704151, 0.2389363, 0.2487957, 0.2243779, 0.3383769, 0.3897291, 
    0.3523037, 0.3716567, 0.408494, 0.3739957, 0.337217, 0.4051063, 
    0.4098835, 0.4451255, 0.4692094, 0.3800277, 0.361383, 0.337771, 
    0.2082432, 0.2141788, 0.2135897, 0.2312396, 0.1714023, 0.2529784, 
    0.1511201, 0.1598543, 0.1592796, 0.2784618, 0.2361904,
  0.269727, 0.2678617, 0.2659963, 0.264131, 0.2622657, 0.2604004, 0.258535, 
    0.2173166, 0.2270998, 0.236883, 0.2466662, 0.2564493, 0.2662325, 
    0.2760157, 0.3307649, 0.3312949, 0.3318249, 0.3323549, 0.3328849, 
    0.3334149, 0.3339449, 0.3283283, 0.3198805, 0.3114326, 0.3029848, 
    0.2945369, 0.2860891, 0.2776412, 0.2712193,
  0.2779807, 0.2936892, 0.1647304, 0.09858744, 0.03431733, 0.119722, 
    0.1227179, 0.1085627, 0.004388134, 0.05172193, 0.1392638, 0.2309882, 
    0.4374457, 0.007079394, 0.174623, 0.281587, 0.3307256, 0.1804325, 
    0.1517076, 0.3593632, 0.6636971, 0.7346855, 0.455348, 0.2307338, 
    0.2492245, 0.2470163, 0.2257747, 0.2179341, 0.2598907,
  0.1519185, 0.1005883, 0.1658015, 0.07088399, 0.1591001, 0.1260321, 
    0.0564223, 0.3410923, 0.3739903, 0.4070966, 0.3639779, 0.2239356, 
    0.1522004, 0.1579417, 0.3257662, 0.422531, 0.4191136, 0.3653811, 
    0.225678, 0.3090386, 0.4011759, 0.4842057, 0.4458318, 0.5375938, 
    0.281722, 0.4053477, 0.4695219, 0.4367228, 0.3066171,
  0.1822703, 0.1919954, 0.1803324, 0.233904, 0.2494388, 0.2573938, 0.2265337, 
    0.1579571, 0.1651151, 0.1919702, 0.242468, 0.2816055, 0.3746362, 0.40786, 
    0.3340793, 0.3807902, 0.3204809, 0.3019152, 0.2470949, 0.2057666, 
    0.2336817, 0.2509097, 0.2998625, 0.2610346, 0.4203501, 0.485523, 
    0.4239709, 0.2305593, 0.2015317,
  0.2687706, 0.3132318, 0.2989353, 0.3001419, 0.3381104, 0.3457313, 
    0.3152602, 0.2633377, 0.2445222, 0.2012821, 0.2077619, 0.2480915, 
    0.174545, 0.1700607, 0.2328278, 0.2006776, 0.1883132, 0.2077698, 
    0.1486193, 0.1479173, 0.1355941, 0.1635386, 0.1955344, 0.2160705, 
    0.1393587, 0.2317484, 0.2138253, 0.2241056, 0.2777413,
  0.1860841, 0.06914164, 0.02885323, 0.06774567, 0.1268257, 0.110412, 
    0.1489339, 0.114324, 0.1070664, 0.05052472, 0.03555439, 0.01146295, 
    0.00486521, 0.0554044, 0.3516848, 0.07614519, 0.09266879, 0.1100056, 
    0.08156594, 0.1266094, 0.134438, 0.1531249, 0.09985037, 0.3173459, 
    0.05420449, 0.09440199, 0.0822774, 0.09540978, 0.2075095,
  0.01952348, 0.01289853, 0.01353472, 0.009876384, 0.007359867, 0.02497312, 
    0.01295252, 0.0174705, 0.02958027, 0.005959211, 0.0001476921, 
    -1.984239e-05, 0.01163984, 0.008151384, 0.03225437, 0.0520521, 
    0.08272523, 0.06082856, 0.09200613, 0.06566405, 0.03315877, 0.02411019, 
    0.02970583, 0.03064888, 0.03606711, 0.01349835, 0.01978295, 0.01877588, 
    0.01104465,
  0.03552853, 0.004113724, 0.001742236, 0.002118337, 0.008398074, 
    0.008870874, 0.001262276, 0.002484587, 0.02113475, 0.0003815647, 
    8.033709e-05, 1.387881e-08, 0.001297872, 0.02673372, 0.007379517, 
    0.01091315, 0.01453456, 0.007437529, 0.007373953, 0.0003678364, 
    0.003270275, 0.002394994, 0.02737075, 0.02768327, 0.05431616, 0.04647011, 
    0.001849434, 0.001693759, 0.01870839,
  0.07536823, 0.02184438, 0.0001820106, 0.06106354, 0.004538988, 0.004218709, 
    0.003886228, 0.005722144, 0.003226341, 0.0002762103, 0.02266128, 
    0.0005513885, 0.06178984, 0.002043606, 0.001337345, 0.0006825379, 
    0.0007189033, 0.006968539, 0.003421059, 0.0005976522, 0.003044986, 
    0.007469088, 0.07640364, 0.005002988, 0.0001643804, 8.49705e-06, 
    0.00377298, 0.001638953, 0.01381041,
  0.01388732, 0.02407586, 0.03188578, 0.0331552, 0.003038351, 0.007559459, 
    0.008062718, 0.001932039, 0.05138109, 0.05134358, 0.007869437, 
    0.007731696, 0.0003295796, 0.001475611, 0.006053485, 0.0006309723, 
    0.001433591, 0.002222224, 0.001162663, 0.001619317, 0.006591442, 
    0.02421663, 0.3069577, 0.1021335, 0.02986728, 0.02720157, 0.02016417, 
    0.006286534, 0.01106976,
  0.0002159197, 0.0001236387, -1.457026e-05, 0.004033772, 0.004370985, 
    0.004404346, 0.01223704, 0.001943704, 0.0001805121, 0.002553967, 
    0.01154125, 0.00361344, 0.003241438, 0.005738284, 0.007648483, 
    0.01130627, 0.00983611, 0.01209978, 0.01324638, 0.01254144, 0.008882202, 
    0.00874836, 0.1861893, 0.03381988, 0.0002641724, 0.004040881, 0.01179034, 
    0.05365168, -0.0006727428,
  1.798571e-07, 4.318673e-07, 1.691721e-07, 0.002025053, 4.010924e-07, 
    3.917693e-05, -0.0001782404, 0.02001781, 0.05326743, 0.07832873, 
    0.007897235, 0.005409287, 0.001049131, 0.0005879696, 0.0005713706, 
    0.002178922, 0.003615452, 0.002550036, 0.04626162, 0.1220535, 
    0.0009004621, 0.04320209, 0.002584767, 0.002499395, 0.003230644, 
    0.01469374, 0.01078923, 0.00898277, 5.871368e-08,
  3.905454e-07, -9.408644e-05, -6.976752e-06, 6.155567e-05, 0.000646921, 
    2.506131e-07, -6.483614e-05, 0.002841411, 0.3067303, 0.04789783, 
    0.1290874, 0.2338565, 0.2364895, 0.1490642, 0.1528026, 0.161012, 
    0.08924365, 0.02955352, 0.06764559, 0.09414802, 0.0006793608, 0.03961566, 
    0.01994711, 0.0882215, 0.08760352, 0.03747164, 0.03809878, 0.02299787, 
    0.01499474,
  0.008589418, 0.002296958, 0.00870177, 0.1450014, 0.01433906, 5.186571e-07, 
    0.09128317, 0.002238699, 1.086728e-05, 0.01249592, 0.1587316, 0.08421137, 
    0.2192987, 0.3491518, 0.3428954, 0.2438079, 0.2429947, 0.3254488, 
    0.1755538, 0.07880569, 0.03112904, 0.08967546, 0.08654836, 0.1283178, 
    0.1498397, 0.2088957, 0.1515894, 0.1039694, 0.1431207,
  0.08153722, 0.09319679, 0.07273378, 0.04630043, 0.016172, 0.01879473, 
    0.02792358, 0.1180634, 0.02769298, 0.03659207, 0.1415363, 0.2656816, 
    0.3626618, 0.2605751, 0.2376372, 0.2862542, 0.3503559, 0.2709472, 
    0.1745274, 0.1144993, 0.03843826, 0.02270592, 0.06879652, 0.2021001, 
    0.1942308, 0.3466552, 0.1893706, 0.1654398, 0.2376266,
  0.09470075, 0.09113316, 0.07186304, 0.1352277, 0.1177935, 0.1319976, 
    0.120783, 0.1152073, 0.1477166, 0.1344308, 0.1104679, 0.07713379, 
    0.1159295, 0.1527064, 0.2445853, 0.482989, 0.2379192, 0.3177558, 
    0.1628486, 0.08408211, 0.05354588, 0.09734264, 0.1532891, 0.2499557, 
    0.3386994, 0.1876827, 0.2950248, 0.2672107, 0.1903391,
  0.2250146, 0.07573631, 0.133077, 0.07507849, 0.1058888, 0.2399558, 
    0.1010648, 0.04434606, 0.02457005, 0.06193744, 0.08575084, 0.07194317, 
    0.05224561, 0.1480456, 0.1896376, 0.3602756, 0.2447697, 0.1240316, 
    0.1594896, 0.1571013, 0.3295569, 0.2788182, 0.1639443, 0.3885888, 
    0.3712265, 0.2631809, 0.1384086, 0.1339628, 0.3896211,
  0.1973828, 0.1833856, 0.2389228, 0.2784152, 0.331571, 0.4017274, 0.4238787, 
    0.3946783, 0.3830667, 0.3708397, 0.3529024, 0.4081219, 0.4488592, 
    0.4625134, 0.450613, 0.3939782, 0.3776679, 0.3385588, 0.201537, 
    0.2274413, 0.2304058, 0.2235584, 0.1759518, 0.2127557, 0.1303395, 
    0.1369874, 0.1327182, 0.2703646, 0.2188207,
  0.1937702, 0.1893401, 0.18491, 0.18048, 0.1760499, 0.1716198, 0.1671897, 
    0.1445824, 0.1541828, 0.1637832, 0.1733837, 0.1829841, 0.1925845, 
    0.2021849, 0.2602311, 0.2638725, 0.267514, 0.2711554, 0.2747969, 
    0.2784383, 0.2820798, 0.2688134, 0.2600017, 0.2511898, 0.2423781, 
    0.2335663, 0.2247545, 0.2159427, 0.1973142,
  0.2899847, 0.2459759, 0.100277, 0.0699413, 0.03598092, 0.05457942, 
    0.04136691, 0.05410485, 0.00174866, 0.01125463, 0.07031695, 0.2290469, 
    0.4371204, -0.002162075, 0.2722279, 0.3588991, 0.4374511, 0.2297787, 
    0.1558752, 0.3565221, 0.6437883, 0.7497617, 0.413639, 0.2155996, 
    0.2672789, 0.3060068, 0.2321831, 0.1839024, 0.259967,
  0.1399397, 0.07938947, 0.1303977, 0.05135413, 0.1451602, 0.1138749, 
    0.03412378, 0.2966538, 0.3371167, 0.3552366, 0.3292114, 0.2261099, 
    0.1344534, 0.1282182, 0.3347101, 0.4325889, 0.4092266, 0.3265488, 
    0.1867711, 0.2691478, 0.3695211, 0.4398546, 0.4060463, 0.5261022, 
    0.2758866, 0.4607513, 0.5066816, 0.4111784, 0.284734,
  0.1338301, 0.1576791, 0.1446915, 0.1779169, 0.1894721, 0.1982071, 
    0.1801949, 0.1179802, 0.1260128, 0.1454532, 0.1991207, 0.2330649, 
    0.3294688, 0.3621873, 0.2686037, 0.3033446, 0.2610906, 0.2473687, 
    0.1991614, 0.1672951, 0.1959708, 0.1895571, 0.2381061, 0.2124048, 
    0.3711678, 0.4330053, 0.3502973, 0.1805343, 0.1504595,
  0.2448751, 0.2842701, 0.2546759, 0.2630242, 0.3125976, 0.3099469, 
    0.2788169, 0.214782, 0.1946597, 0.1547756, 0.1540642, 0.1695523, 
    0.1220121, 0.1167471, 0.2013703, 0.1574286, 0.1412964, 0.1530035, 
    0.1123592, 0.1210162, 0.1042516, 0.1317841, 0.1502825, 0.1848676, 
    0.1223472, 0.1865366, 0.1695773, 0.1790848, 0.2377634,
  0.1445189, 0.04537892, 0.01485994, 0.04266858, 0.08700831, 0.07058004, 
    0.09355239, 0.07480562, 0.06487478, 0.03270939, 0.02346306, 0.006541719, 
    0.002608317, 0.03014703, 0.3083272, 0.0544411, 0.06766847, 0.08735996, 
    0.06519904, 0.09245818, 0.1024327, 0.1139699, 0.06737273, 0.297585, 
    0.0383663, 0.05669734, 0.05884984, 0.06756289, 0.1759372,
  0.01092873, 0.005838503, 0.01261766, 0.004511687, 0.002846345, 0.01229667, 
    0.008339122, 0.00998964, 0.0171713, 0.003894222, 0.0001493039, 
    -6.877113e-06, 0.009622602, 0.002590135, 0.0182804, 0.03247941, 
    0.04863145, 0.03524394, 0.06312966, 0.03238949, 0.01614759, 0.01511059, 
    0.01548286, 0.02680314, 0.03052599, 0.008226849, 0.009391443, 
    0.008263926, 0.005126242,
  0.01961251, 0.002959465, 0.0009011542, 0.001169809, 0.003177443, 
    0.003569324, 0.0005226929, 0.0005481719, 0.008554641, 0.0002258444, 
    0.0001763236, 1.149049e-08, 0.0006141556, 0.01233425, 0.002050438, 
    0.003913958, 0.005156402, 0.00276343, 0.003228631, 0.0002011279, 
    0.001502106, 0.001205513, 0.01444742, 0.01901058, 0.03847291, 0.05185806, 
    0.0009472317, 0.0008254625, 0.009225909,
  0.03949796, 0.01840835, -0.0001357516, 0.03833824, 0.001277709, 
    0.001741304, 0.001550824, 0.0008581662, 0.001023826, -0.0006436521, 
    0.01555707, 0.0002999328, 0.03255673, 0.000480487, 0.000421213, 
    0.0002826263, 0.000290189, 0.00346351, 0.001114031, 0.0002606395, 
    0.001614974, 0.00364016, 0.03996351, 0.002805491, 9.439669e-05, 
    4.923653e-06, 0.0010731, 0.0008568577, 0.007359795,
  0.006050503, 0.04016817, 0.03671936, 0.02376613, 0.001576785, 0.003660932, 
    0.004483307, 0.0009874764, 0.03964202, 0.05733457, 0.003616174, 
    0.004332344, 0.0001301762, 0.0007819121, 0.003132169, 0.0002425768, 
    0.0005156043, 0.0009258767, 0.0004045248, 0.0003976519, 0.001644503, 
    0.008355968, 0.1387556, 0.1021274, 0.02973298, 0.01848828, 0.01072645, 
    0.003320335, 0.004128674,
  8.418523e-05, 5.84863e-05, -1.026393e-05, 0.005350275, 0.002807668, 
    0.002546566, 0.002788186, 0.001005763, -0.0001850332, 0.001336088, 
    0.004663371, 0.001601079, 0.0007142867, 0.001679503, 0.002005538, 
    0.003368262, 0.004154881, 0.005424926, 0.003107662, 0.005698712, 
    0.004764598, 0.004032881, 0.1603817, 0.03348145, 2.527601e-05, 
    0.001384246, 0.005082155, 0.02669789, -0.001055671,
  1.727491e-07, 4.167512e-07, 1.667417e-07, 0.00137087, 3.944212e-07, 
    -1.574575e-05, -0.0001897431, 0.003497991, 0.04043855, 0.03706471, 
    0.003271461, 0.002118076, 0.0003490794, 0.0002709606, 0.0002445856, 
    0.0006977638, 0.001131029, 0.001322239, 0.02470041, 0.07654004, 
    0.0005110546, 0.03619023, 0.0008838618, -0.0004885808, 0.001579786, 
    0.006785536, 0.00551111, 0.005074367, 5.692476e-08,
  4.586416e-07, -8.468363e-05, -1.974745e-06, -4.195246e-06, 0.0004396511, 
    2.404643e-07, -6.65367e-05, 0.003784262, 0.2910758, 0.0361941, 0.1302636, 
    0.1810088, 0.1753827, 0.0985461, 0.08540814, 0.1032526, 0.05616387, 
    0.01415934, 0.03847037, 0.05452189, 0.0004220424, 0.0339755, 0.009684531, 
    0.0457353, 0.06722927, 0.01586781, 0.02387864, 0.01165677, 0.01278564,
  0.006492148, 0.001685921, 0.005225513, 0.1402552, 0.007357035, 
    5.818043e-07, 0.07888268, 0.00133642, -1.114965e-05, 0.009142576, 
    0.151923, 0.07998477, 0.2035693, 0.3255699, 0.2914612, 0.1928105, 
    0.1830707, 0.2892051, 0.1266657, 0.07305746, 0.02468702, 0.07489362, 
    0.06604808, 0.1071724, 0.09947193, 0.1511906, 0.09604678, 0.06261467, 
    0.1120656,
  0.05210443, 0.07687646, 0.05556874, 0.03658255, 0.01080598, 0.01311054, 
    0.02103849, 0.1002263, 0.0222978, 0.03176674, 0.125402, 0.2391797, 
    0.3420089, 0.2094219, 0.196494, 0.2304345, 0.2833413, 0.2206259, 
    0.1601485, 0.09602565, 0.02871138, 0.01607638, 0.05617414, 0.1790573, 
    0.1666162, 0.3089216, 0.1322321, 0.11382, 0.1893282,
  0.09983874, 0.07887918, 0.06270251, 0.1157486, 0.09957602, 0.1128477, 
    0.1077219, 0.09621243, 0.1263317, 0.1181663, 0.1014588, 0.05469505, 
    0.09177711, 0.1196176, 0.2014738, 0.4248693, 0.1986649, 0.2494708, 
    0.1347296, 0.07585205, 0.04224434, 0.06783995, 0.1515812, 0.2305165, 
    0.2692623, 0.1569088, 0.2508176, 0.228339, 0.1512201,
  0.196859, 0.05699415, 0.1118063, 0.05798038, 0.0857635, 0.2083172, 
    0.08462825, 0.02628907, 0.01652995, 0.05420629, 0.06801474, 0.0530345, 
    0.06193221, 0.1307201, 0.192185, 0.3089204, 0.2576816, 0.1254367, 
    0.165962, 0.1503833, 0.2986465, 0.3225805, 0.1327007, 0.3513932, 
    0.3300155, 0.2081249, 0.129637, 0.1110444, 0.3605428,
  0.1491402, 0.1497275, 0.2291996, 0.2693309, 0.286638, 0.3364089, 0.4008914, 
    0.3512461, 0.3351924, 0.3515457, 0.3534642, 0.3875744, 0.4174218, 
    0.4367317, 0.3964764, 0.3721691, 0.3512034, 0.320384, 0.2051929, 
    0.2431926, 0.2200673, 0.2060824, 0.1450625, 0.1743998, 0.1123369, 
    0.101979, 0.1084658, 0.2401986, 0.1778636,
  0.1462742, 0.1407825, 0.1352908, 0.1297992, 0.1243075, 0.1188158, 
    0.1133242, 0.08199498, 0.09186076, 0.1017265, 0.1115923, 0.1214581, 
    0.1313239, 0.1411897, 0.1992767, 0.2045269, 0.2097771, 0.2150273, 
    0.2202775, 0.2255278, 0.230778, 0.2149098, 0.2052855, 0.1956612, 
    0.1860368, 0.1764125, 0.1667881, 0.1571638, 0.1506675,
  0.3304689, 0.1834798, 0.06160196, 0.02255329, 0.0005017065, 0.01926953, 
    0.004518808, 0.004412643, 0.02670772, 0.03165247, 0.04894365, 0.1946773, 
    0.3725669, -0.005143736, 0.3516735, 0.4154928, 0.4359503, 0.2270657, 
    0.1408601, 0.3687312, 0.6355458, 0.7751976, 0.366315, 0.1772678, 
    0.2578128, 0.352997, 0.2515163, 0.1561028, 0.2518289,
  0.1242167, 0.06541348, 0.1062608, 0.0387149, 0.1336343, 0.09971581, 
    0.02331001, 0.2408825, 0.2999845, 0.3008761, 0.2889091, 0.2462569, 
    0.1155789, 0.1115659, 0.3284927, 0.3861216, 0.3857138, 0.2717731, 
    0.1482976, 0.2377025, 0.3252071, 0.3749214, 0.3527329, 0.4782834, 
    0.2750124, 0.477469, 0.48125, 0.3476762, 0.2657404,
  0.09482427, 0.1181061, 0.1097476, 0.1321058, 0.141104, 0.1483208, 0.136469, 
    0.08727843, 0.09460313, 0.1045911, 0.1564827, 0.1831401, 0.2809058, 
    0.2856423, 0.2015244, 0.2208483, 0.2004151, 0.1902593, 0.1570164, 
    0.1320913, 0.1520933, 0.1323906, 0.1742681, 0.1628079, 0.3023154, 
    0.3665198, 0.2796182, 0.1379347, 0.1040944,
  0.2023884, 0.2377794, 0.202052, 0.2159561, 0.2677096, 0.257968, 0.2377888, 
    0.1660151, 0.1453021, 0.1098049, 0.1055689, 0.1084657, 0.07503631, 
    0.07331982, 0.1607887, 0.1127048, 0.1024721, 0.1059192, 0.07284403, 
    0.08907539, 0.07512117, 0.09166136, 0.1050341, 0.1609374, 0.1008531, 
    0.142924, 0.1278721, 0.1365723, 0.1996204,
  0.1011218, 0.02948123, 0.007810225, 0.02478304, 0.05196978, 0.04110048, 
    0.05563627, 0.04476041, 0.03647638, 0.02251949, 0.01374017, 0.00348653, 
    0.001763291, 0.01623368, 0.2691101, 0.03525952, 0.04537344, 0.05959553, 
    0.04357101, 0.059759, 0.06724034, 0.08019878, 0.03901651, 0.27641, 
    0.02640338, 0.03537545, 0.03546137, 0.04015039, 0.1307465,
  0.006733176, 0.003702874, 0.01310778, 0.002273035, 0.001431063, 
    0.005346412, 0.005562979, 0.006040662, 0.009599907, 0.002569158, 
    2.247615e-05, -8.165048e-06, 0.00733707, 0.001081675, 0.00920139, 
    0.0174957, 0.02855095, 0.016892, 0.03692898, 0.01481687, 0.006782393, 
    0.008640874, 0.008864156, 0.01881944, 0.02617393, 0.004427645, 
    0.004721012, 0.004077758, 0.003072261,
  0.01304174, 0.002051522, 0.0003231316, 0.0007820253, 0.0005298565, 
    0.00143771, 0.0003412355, 0.0003121094, 0.00310674, 0.0001622229, 
    9.409495e-05, 9.990398e-09, 0.0004324884, 0.005601684, 0.0008556077, 
    0.002112254, 0.002520576, 0.001249024, 0.001491062, 0.0001352587, 
    0.0008076387, 0.0007659924, 0.009312393, 0.01527362, 0.02689075, 
    0.05362687, 0.0006367485, 0.0005423193, 0.005905533,
  0.02491136, 0.01374176, -0.0002235801, 0.02151816, 0.0005031365, 
    0.001020011, 0.0006634454, 0.00021749, 0.0005230883, -0.0004252813, 
    0.009777043, 0.0001869418, 0.01641966, 0.0002462821, 0.0001440854, 
    0.000184984, 0.000149721, 0.001490427, 0.0003960575, 0.0001531305, 
    0.001038817, 0.002235293, 0.02545114, 0.004224671, 0.0005075334, 
    2.865745e-06, 0.0001291146, 0.0005397493, 0.00478295,
  0.003663389, 0.04885117, 0.03427605, 0.01685287, 0.0009946314, 0.001691306, 
    0.002345475, 0.0006349572, 0.03174495, 0.062866, 0.001676211, 
    0.002498045, 7.665021e-05, 0.0004978739, 0.00159522, 0.0001458781, 
    0.0002956903, 0.0005431665, 0.0002266214, 0.0002198275, 0.0008884478, 
    0.004781041, 0.08091378, 0.08680288, 0.02781325, 0.009115203, 
    0.005155533, 0.001680255, 0.002416198,
  4.405259e-05, 3.387679e-05, -6.709904e-06, 0.005688572, 0.001385428, 
    0.001710063, -0.0002559217, 0.0006604768, -0.0001212028, 0.0008491554, 
    0.001904881, 0.0009752783, 0.0002631845, 0.0005758031, 0.0005618234, 
    0.001151274, 0.001915593, 0.002403254, 0.001066072, 0.003273125, 
    0.003204475, 0.001879334, 0.1301302, 0.03574711, 1.435316e-05, 
    0.0006736838, 0.00292481, 0.0166493, -0.000670578,
  1.689965e-07, 4.064436e-07, 1.654086e-07, 0.0007376375, 3.896103e-07, 
    -1.082514e-05, -0.0001223413, 0.001539344, 0.03367971, 0.01511119, 
    0.001867115, 0.001213082, 0.0001988308, 0.0001687532, 0.0001515666, 
    0.0004218727, 0.0006401027, 0.0008430281, 0.01597964, 0.0547186, 
    0.0003572169, 0.02982017, 0.0003619775, -0.0009890932, 0.0009991259, 
    0.004146075, 0.003468852, 0.003349286, 5.633758e-08,
  4.714725e-07, -3.611207e-05, -1.20834e-06, -1.439061e-05, 0.000347307, 
    2.33086e-07, -6.783921e-05, 0.004516033, 0.2678495, 0.02259899, 
    0.1110482, 0.1211755, 0.1145259, 0.05336025, 0.06275417, 0.06134724, 
    0.03141008, 0.007653979, 0.02565777, 0.03662314, 0.0002748393, 
    0.02652366, 0.005502537, 0.02302127, 0.04069708, 0.007612601, 0.01616875, 
    0.006719242, 0.01216898,
  0.004289412, 0.0008320828, 0.003110904, 0.1240937, 0.004453436, 
    5.681286e-07, 0.06737007, 0.000942678, -1.801431e-05, 0.00671899, 
    0.1362039, 0.08016715, 0.1818867, 0.288494, 0.2303053, 0.1431556, 
    0.1269852, 0.2314677, 0.09455702, 0.06442872, 0.01951681, 0.06039879, 
    0.05005092, 0.08539814, 0.06235923, 0.09354073, 0.05270094, 0.03244343, 
    0.07713536,
  0.03922995, 0.06220531, 0.03950124, 0.02908793, 0.007530469, 0.008742749, 
    0.01590627, 0.0866413, 0.01867861, 0.02618572, 0.1083837, 0.2140237, 
    0.3036124, 0.1638954, 0.1616992, 0.1867992, 0.2083022, 0.1638728, 
    0.1265448, 0.08047258, 0.01914725, 0.01269291, 0.0438513, 0.1555053, 
    0.1415845, 0.2621658, 0.08243045, 0.07355689, 0.1318927,
  0.07890879, 0.06482005, 0.05237758, 0.0913678, 0.08129345, 0.09303258, 
    0.09180814, 0.07762586, 0.106475, 0.09808336, 0.09071408, 0.04150432, 
    0.07242849, 0.08842395, 0.1545391, 0.3333669, 0.1635095, 0.1962112, 
    0.1069184, 0.06813048, 0.03265116, 0.05223632, 0.170649, 0.2084064, 
    0.2116611, 0.1334197, 0.1864982, 0.1527713, 0.1116224,
  0.1665758, 0.04134724, 0.09572209, 0.0482766, 0.0655861, 0.151223, 
    0.07573912, 0.01930038, 0.01611603, 0.04915005, 0.05940194, 0.04478534, 
    0.07569204, 0.1142197, 0.159623, 0.2305576, 0.2355172, 0.1151857, 
    0.1679451, 0.1538374, 0.2821087, 0.319925, 0.1100109, 0.3062239, 
    0.2734919, 0.1743582, 0.1241599, 0.09543462, 0.3115404,
  0.129896, 0.1379464, 0.1715848, 0.2284486, 0.213659, 0.2597406, 0.3126835, 
    0.2857605, 0.3003886, 0.3118231, 0.3051127, 0.3359166, 0.3220584, 
    0.347244, 0.3257059, 0.317171, 0.3006217, 0.2749778, 0.2001778, 
    0.2270057, 0.2147511, 0.1753487, 0.115841, 0.1556038, 0.09101921, 
    0.07802007, 0.08736924, 0.2170002, 0.1374757,
  0.1197918, 0.1161266, 0.1124615, 0.1087963, 0.1051311, 0.101466, 
    0.09780082, 0.08549565, 0.09245449, 0.09941332, 0.1063721, 0.113331, 
    0.1202898, 0.1272486, 0.1451044, 0.1494392, 0.1537741, 0.158109, 
    0.1624439, 0.1667788, 0.1711137, 0.1698356, 0.1622071, 0.1545785, 
    0.1469499, 0.1393214, 0.1316928, 0.1240643, 0.1227239,
  0.410231, 0.1421735, 0.04915243, 0.005355892, 0.001461716, 0.007364472, 
    0.005779859, 0.002883017, 0.001127333, 0.02280847, 0.04359207, 0.152953, 
    0.3197132, -0.005523743, 0.4191004, 0.4295393, 0.4483228, 0.2291664, 
    0.1177048, 0.4207714, 0.6230697, 0.8041072, 0.3391725, 0.1538457, 
    0.2506306, 0.371922, 0.2658703, 0.1429361, 0.2514217,
  0.1174764, 0.05860229, 0.09575931, 0.03279164, 0.1210454, 0.0893051, 
    0.01848899, 0.2021348, 0.272985, 0.2562057, 0.2870382, 0.2633195, 
    0.1025919, 0.1029805, 0.3329908, 0.3509404, 0.3568208, 0.2308595, 
    0.12803, 0.2154501, 0.2973355, 0.3317519, 0.3160951, 0.419288, 0.2684858, 
    0.4377095, 0.4224223, 0.2898988, 0.2476724,
  0.0745652, 0.09313749, 0.08677237, 0.1059555, 0.1129993, 0.1194781, 
    0.1097174, 0.06778081, 0.07390582, 0.08170044, 0.1266601, 0.1481169, 
    0.2396162, 0.2306857, 0.156357, 0.1706003, 0.1603072, 0.156368, 
    0.1270758, 0.1060041, 0.1203455, 0.09979207, 0.1349225, 0.1239832, 
    0.249214, 0.3049037, 0.2319649, 0.1103938, 0.07935882,
  0.1675702, 0.2027237, 0.1707785, 0.1807466, 0.2320476, 0.2199537, 
    0.2079689, 0.1323484, 0.1141863, 0.08307271, 0.07505955, 0.07715206, 
    0.04999999, 0.04884909, 0.1295095, 0.08212683, 0.07478913, 0.07207632, 
    0.04945961, 0.06636485, 0.05470432, 0.06732819, 0.0774994, 0.1546981, 
    0.07665386, 0.1052344, 0.09966749, 0.109466, 0.1712564,
  0.06727849, 0.01802988, 0.005013593, 0.01461522, 0.03200659, 0.02341601, 
    0.03474426, 0.02945028, 0.02131227, 0.01531739, 0.00764606, 0.00191552, 
    0.00138625, 0.009364655, 0.2391494, 0.0211546, 0.03005017, 0.04128304, 
    0.02819502, 0.03808356, 0.04416689, 0.05475762, 0.0243719, 0.2533767, 
    0.01957989, 0.02126494, 0.0210414, 0.02346067, 0.09200875,
  0.004701577, 0.002752617, 0.01328629, 0.001379674, 0.001006707, 
    0.003076911, 0.003080645, 0.004134602, 0.006256131, 0.001702041, 
    -4.89544e-05, -5.567462e-06, 0.008290159, 0.0006939308, 0.004604252, 
    0.008319368, 0.01679809, 0.008906643, 0.02152146, 0.008034956, 
    0.003592851, 0.00480297, 0.006232313, 0.01467766, 0.0228576, 0.002376074, 
    0.002722945, 0.002348029, 0.002224676,
  0.009788642, 0.001576613, 6.534132e-05, 0.000581654, -0.0004053485, 
    0.0007187881, 0.0002582191, 0.0002243142, 0.001725444, 0.0001262856, 
    4.123746e-05, 9.090988e-09, 0.0003387138, 0.002843978, 0.0005378451, 
    0.001449775, 0.001553998, 0.0006960951, 0.0007479681, 0.0001024158, 
    0.0005227982, 0.0005596846, 0.006849858, 0.01280857, 0.02218732, 
    0.05126622, 0.0004668954, 0.0004055398, 0.004322661,
  0.01793147, 0.008373125, 4.539412e-06, 0.01558974, 0.0003255113, 
    0.0007309064, 0.0003829534, 0.0001133183, 0.0003038681, -0.0002949244, 
    0.00671999, 0.0001369063, 0.008628101, 0.0001456927, 9.416827e-05, 
    0.0001371703, 0.0001002239, 0.0006814961, 0.0002364841, 0.0001084763, 
    0.0007636073, 0.001596726, 0.01853726, 0.008749587, 0.001571283, 
    1.109918e-05, -3.086446e-05, 0.0003912018, 0.003550243,
  0.002539128, 0.04890571, 0.02559245, 0.01198973, 0.0007163339, 
    0.0008272298, 0.001362666, 0.0004638752, 0.0253759, 0.0640178, 
    0.000845247, 0.001658327, 5.404881e-05, 0.0003592921, 0.0008240399, 
    0.0001054267, 0.0002133506, 0.0003795285, 0.0001540544, 0.0001521805, 
    0.0006038825, 0.003298027, 0.05545429, 0.06057039, 0.02358664, 
    0.00420313, 0.002528788, 0.001060044, 0.001695805,
  9.259042e-05, 9.14534e-06, -3.775364e-06, 0.004981176, 0.0007399899, 
    0.001277807, -0.0009439036, 0.0004778351, -7.205363e-05, 0.0006288578, 
    0.001046427, 0.0006342512, 0.0001471826, 0.000295237, 0.0002244694, 
    0.0004473378, 0.0009160445, 0.001241316, 0.0006144481, 0.002258654, 
    0.002426309, 0.001056514, 0.1183067, 0.03762747, 8.965466e-06, 
    0.0004203088, 0.00202609, 0.01202528, -5.529728e-08,
  1.66167e-07, 3.997932e-07, 1.644625e-07, 0.0005038213, 3.848644e-07, 
    -7.933277e-06, -8.024747e-05, 0.001012627, 0.03799513, 0.007792893, 
    0.00132883, 0.0008470141, 0.0001398596, 0.000121607, 0.0001105987, 
    0.0003066258, 0.0004841499, 0.0006156524, 0.01175762, 0.04281007, 
    0.00027613, 0.02447257, 0.0002252449, -0.001189379, 0.0007220671, 
    0.002995744, 0.002511066, 0.00249864, 5.620898e-08,
  4.746905e-07, -2.132203e-05, -8.384883e-07, -1.080127e-05, 0.0002796464, 
    2.263784e-07, -6.752484e-05, 0.004940654, 0.2513947, 0.01403912, 
    0.09380762, 0.07205494, 0.07282572, 0.03402773, 0.0457516, 0.03942901, 
    0.01814773, 0.005270619, 0.01941115, 0.02757099, 0.0001967694, 
    0.02146294, 0.006092828, 0.01306651, 0.02055342, 0.004606459, 0.01132909, 
    0.004663455, 0.009276293,
  0.002521374, 0.0001851708, 0.002115446, 0.1127723, 0.003233293, 
    5.550078e-07, 0.05785393, 0.0007510652, -2.064229e-05, 0.005204744, 
    0.1212792, 0.07321854, 0.1539777, 0.2444218, 0.1755536, 0.1067269, 
    0.08928382, 0.1666579, 0.06571702, 0.05927439, 0.01648991, 0.04994763, 
    0.03722135, 0.06830851, 0.04306471, 0.05853575, 0.03087704, 0.01782413, 
    0.05342956,
  0.03775577, 0.05028107, 0.02796565, 0.02298506, 0.005593771, 0.00660208, 
    0.01275145, 0.07727006, 0.01723571, 0.02286697, 0.0927895, 0.1947663, 
    0.2345589, 0.1334131, 0.1356975, 0.153739, 0.1544455, 0.1179044, 
    0.0936238, 0.07156202, 0.01488241, 0.01043758, 0.03545759, 0.1383037, 
    0.1210701, 0.2075282, 0.05322155, 0.04715764, 0.09015889,
  0.06108536, 0.05164299, 0.04494303, 0.07558755, 0.07057117, 0.07777545, 
    0.08313259, 0.06683808, 0.09589258, 0.08542025, 0.07997166, 0.03848201, 
    0.0654024, 0.07565261, 0.1218895, 0.2634851, 0.1382339, 0.1621819, 
    0.1041214, 0.05983789, 0.02876444, 0.04947371, 0.1603163, 0.194478, 
    0.165103, 0.1138845, 0.1327371, 0.09557332, 0.07887936,
  0.1240706, 0.0299798, 0.08515544, 0.03973584, 0.05706757, 0.1137932, 
    0.07990948, 0.02500645, 0.02494761, 0.04820039, 0.05580901, 0.04325904, 
    0.1034492, 0.1088709, 0.1362557, 0.1947653, 0.2357806, 0.1046646, 
    0.1586388, 0.1599505, 0.261, 0.3011975, 0.1140359, 0.2797294, 0.2493033, 
    0.148607, 0.1399529, 0.08741114, 0.2596238,
  0.1167684, 0.1369655, 0.1352786, 0.1609226, 0.1558578, 0.1870763, 
    0.2154951, 0.2000725, 0.2427379, 0.2481516, 0.2390487, 0.2653415, 
    0.2408133, 0.2610517, 0.2590349, 0.2585779, 0.229154, 0.2247697, 
    0.1725202, 0.1944431, 0.2020529, 0.152022, 0.09918277, 0.1414777, 
    0.0767578, 0.063508, 0.0740408, 0.2030188, 0.1264487,
  0.1088978, 0.1052621, 0.1016263, 0.09799059, 0.09435487, 0.09071913, 
    0.08708341, 0.08453381, 0.09120835, 0.09788288, 0.1045574, 0.111232, 
    0.1179065, 0.124581, 0.135769, 0.1400553, 0.1443415, 0.1486277, 0.152914, 
    0.1572002, 0.1614864, 0.1606748, 0.1533497, 0.1460246, 0.1386996, 
    0.1313746, 0.1240495, 0.1167245, 0.1118064,
  0.3479094, 0.08747892, 0.03145437, 0.004625401, 0.00090971, 0.005764563, 
    0.005314622, 0.002729503, 0.0007736965, 0.01685616, 0.03768448, 
    0.1344914, 0.3018792, -0.005269331, 0.4924117, 0.4288682, 0.4122508, 
    0.2611133, 0.1235106, 0.4538516, 0.5901955, 0.8000121, 0.3425182, 
    0.1544909, 0.2389031, 0.3702553, 0.285054, 0.1448143, 0.2534832,
  0.115358, 0.06448407, 0.08918658, 0.0328666, 0.1374305, 0.07674992, 
    0.01662032, 0.1895307, 0.2641983, 0.2481522, 0.2713484, 0.2698165, 
    0.09870444, 0.09804, 0.3348456, 0.3364098, 0.3466166, 0.2095964, 
    0.1168638, 0.1976461, 0.276958, 0.3165303, 0.2994844, 0.3826464, 
    0.2586446, 0.4031601, 0.379237, 0.254922, 0.2262785,
  0.06422618, 0.07894117, 0.07440189, 0.09280749, 0.09893908, 0.1040844, 
    0.0951653, 0.05702818, 0.06201496, 0.07005948, 0.1112915, 0.1286961, 
    0.2072291, 0.197561, 0.1328624, 0.1448863, 0.1398515, 0.1400174, 
    0.1102702, 0.08998187, 0.1012813, 0.08295554, 0.1129945, 0.09953722, 
    0.2124103, 0.2645453, 0.2066714, 0.09552166, 0.06745651,
  0.1423388, 0.1704457, 0.1434567, 0.1477014, 0.2018704, 0.1850079, 
    0.1785757, 0.1114706, 0.0980981, 0.06931037, 0.06035944, 0.06208653, 
    0.03887695, 0.03706317, 0.1016631, 0.06161184, 0.05844025, 0.05166269, 
    0.03761396, 0.05449015, 0.04437681, 0.05309168, 0.06152035, 0.1806472, 
    0.05833243, 0.0809534, 0.08498507, 0.09312093, 0.1462788,
  0.05141096, 0.01233065, 0.003811886, 0.01023927, 0.02198764, 0.01624577, 
    0.02547654, 0.02183837, 0.01498112, 0.01083323, 0.004700731, 0.001489864, 
    0.001196826, 0.006808206, 0.2534348, 0.01339228, 0.02059165, 0.03102488, 
    0.02041513, 0.02772908, 0.03060313, 0.03683125, 0.01706091, 0.2586418, 
    0.01546469, 0.01438574, 0.01347661, 0.01525334, 0.06804878,
  0.003791938, 0.002287904, 0.01628807, 0.001017676, 0.0008409099, 
    0.00225829, 0.002168352, 0.003127658, 0.004728028, 0.001286572, 
    -6.704092e-05, -2.992828e-06, 0.01494902, 0.0005559899, 0.002751822, 
    0.004949208, 0.009630371, 0.005887434, 0.01383621, 0.005090538, 
    0.002576437, 0.003241861, 0.005025278, 0.01295151, 0.03815763, 
    0.001541987, 0.002018618, 0.001735732, 0.001839563,
  0.008185137, 0.001358004, -8.264672e-05, 0.0004815701, -0.0008016769, 
    0.0004833466, 0.0002179888, 0.0001871159, 0.001073815, 0.0001070776, 
    2.992881e-05, 8.552901e-09, 0.0002889616, 0.001796207, 0.0004220185, 
    0.001126361, 0.00118481, 0.0005141764, 0.0005064863, 8.607771e-05, 
    0.0003975373, 0.0004607117, 0.005661463, 0.01132718, 0.03652582, 
    0.05473954, 0.0003866748, 0.0003373511, 0.003539531,
  0.01455102, 0.004393557, 0.002343675, 0.02543116, 0.0002563074, 
    0.0005868917, 0.0002868273, 8.813512e-05, 0.0002274979, -0.0003374457, 
    0.005297855, 0.0001156218, 0.005344696, 0.000114005, 8.110856e-05, 
    0.0001129894, 7.953036e-05, 0.0004241203, 0.0001829997, 8.832872e-05, 
    0.0006344282, 0.00130902, 0.01519684, 0.04702835, 0.02740595, 
    0.0005302813, -7.701854e-05, 0.0003235881, 0.002961419,
  0.002033298, 0.07519222, 0.02787553, 0.01221732, 0.0005718645, 
    0.0005481961, 0.0009373817, 0.0003800793, 0.0306624, 0.09010632, 
    0.0005786021, 0.001275536, 4.339924e-05, 0.0002892578, 0.0005216555, 
    8.653769e-05, 0.0001737464, 0.000302414, 0.0001221, 0.0001203791, 
    0.0004858258, 0.002624937, 0.04326499, 0.07154274, 0.06005062, 
    0.002576614, 0.001646729, 0.0008164098, 0.001358659,
  0.003302969, -1.967686e-05, -6.658551e-06, 0.006431667, 0.0004700738, 
    0.001057587, -0.002667031, 0.000391031, -0.001006569, 0.000524026, 
    0.0007659678, 0.000498404, 0.0001071747, 0.0002244718, 0.0001585509, 
    0.0002827691, 0.0005426314, 0.0008662035, 0.0004943078, 0.001815693, 
    0.00201451, 0.0007422449, 0.1764326, 0.05031925, 6.920263e-06, 
    0.0003349346, 0.00163457, 0.009735073, 0.02492581,
  1.649037e-07, 3.951908e-07, 1.639882e-07, 0.0003943831, 3.825284e-07, 
    -6.322065e-06, -5.784749e-05, 0.0007045197, 0.08527806, 0.004370415, 
    0.001069375, 0.0006744012, 0.0001151838, 0.000101005, 9.03815e-05, 
    0.0002531322, 0.0004107667, 0.0005138821, 0.009736948, 0.03652167, 
    0.0002335262, 0.02237607, 0.0001765587, -0.001716491, 0.000589327, 
    0.002431182, 0.002059206, 0.002106312, 5.657296e-08,
  4.770579e-07, -1.141839e-05, -6.216649e-07, -6.780853e-06, 0.0002366246, 
    2.234629e-07, -7.134914e-05, 0.006298909, 0.2606399, 0.01754331, 
    0.06853798, 0.0435464, 0.0472948, 0.02275769, 0.03492851, 0.02420533, 
    0.01168873, 0.004028746, 0.01623386, 0.02277736, 0.0001501877, 
    0.04392941, 0.02204186, 0.008466698, 0.01124471, 0.003389052, 
    0.008553892, 0.003777343, 0.007021805,
  0.001832371, 3.497204e-05, 0.001716356, 0.1101237, 0.002610593, 
    5.499814e-07, 0.05168576, 0.0006550947, -2.194866e-05, 0.004335882, 
    0.1178119, 0.05959539, 0.1236374, 0.1853947, 0.1391423, 0.08267471, 
    0.06672084, 0.1227982, 0.04979489, 0.05989117, 0.01505261, 0.04895478, 
    0.03288665, 0.05616724, 0.03410737, 0.03852377, 0.02084914, 0.01179201, 
    0.0415223,
  0.03061105, 0.04734638, 0.02374201, 0.02012147, 0.004586069, 0.005562736, 
    0.01123286, 0.07505868, 0.01920985, 0.02427668, 0.09787756, 0.1997297, 
    0.1763098, 0.1124834, 0.1114964, 0.1321877, 0.1235004, 0.09040302, 
    0.07370927, 0.0757294, 0.01291653, 0.009928863, 0.03962031, 0.1546592, 
    0.1106259, 0.1654046, 0.04010786, 0.03344389, 0.06560022,
  0.0444948, 0.05166754, 0.0421403, 0.07451779, 0.07528158, 0.08288585, 
    0.08958472, 0.08019984, 0.1060776, 0.09127635, 0.08247021, 0.05563495, 
    0.09528668, 0.08126977, 0.1030338, 0.2238031, 0.1325893, 0.1464607, 
    0.1307088, 0.06290074, 0.030573, 0.07051999, 0.1563045, 0.1950839, 
    0.1420081, 0.09920099, 0.103431, 0.0714671, 0.06364074,
  0.09629168, 0.021074, 0.08224464, 0.03470103, 0.06532987, 0.09819545, 
    0.1041342, 0.05390827, 0.05093174, 0.07666779, 0.07715678, 0.05231095, 
    0.1607953, 0.1145555, 0.1402056, 0.1714372, 0.254434, 0.1071318, 
    0.1618293, 0.1531865, 0.2415819, 0.2913605, 0.1586809, 0.2779827, 
    0.2236658, 0.1329602, 0.1906721, 0.0841836, 0.2150545,
  0.1327226, 0.1301705, 0.1259818, 0.1313576, 0.1293601, 0.156966, 0.1769489, 
    0.1634416, 0.1991432, 0.2067314, 0.2016762, 0.2105934, 0.1997329, 
    0.2206492, 0.2224358, 0.223944, 0.1923757, 0.1961853, 0.1553807, 
    0.1731807, 0.187161, 0.1393626, 0.09249684, 0.1341716, 0.06965475, 
    0.0549037, 0.06714649, 0.1900134, 0.1460582 ;

 average_DT = 730 ;

 average_T1 = 136.5 ;

 average_T2 = 866.5 ;

 climatology_bounds =
  136.5, 866.5 ;

 lat = -89.5, -79.5, -69.5, -59.5, -49.5, -39.5, -29.5, -19.5, -9.5, 0.5, 
    10.5, 20.5, 30.5, 40.5, 50.5, 60.5, 70.5, 80.5 ;

 lat_bnds =
  -90, -89,
  -80, -79,
  -70, -69,
  -60, -59,
  -50, -49,
  -40, -39,
  -30, -29,
  -20, -19,
  -10, -9,
  0, 1,
  10, 11,
  20, 21,
  30, 31,
  40, 41,
  50, 51,
  60, 61,
  70, 71,
  80, 81 ;

 lon = 0.625, 13.125, 25.625, 38.125, 50.625, 63.125, 75.625, 88.125, 
    100.625, 113.125, 125.625, 138.125, 150.625, 163.125, 175.625, 188.125, 
    200.625, 213.125, 225.625, 238.125, 250.625, 263.125, 275.625, 288.125, 
    300.625, 313.125, 325.625, 338.125, 350.625 ;

 lon_bnds =
  0, 1.25,
  12.5, 13.75,
  25, 26.25,
  37.5, 38.75,
  50, 51.25,
  62.5, 63.75,
  75, 76.25,
  87.5, 88.75,
  100, 101.25,
  112.5, 113.75,
  125, 126.25,
  137.5, 138.75,
  150, 151.25,
  162.5, 163.75,
  175, 176.25,
  187.5, 188.75,
  200, 201.25,
  212.5, 213.75,
  225, 226.25,
  237.5, 238.75,
  250, 251.25,
  262.5, 263.75,
  275, 276.25,
  287.5, 288.75,
  300, 301.25,
  312.5, 313.75,
  325, 326.25,
  337.5, 338.75,
  350, 351.25 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 time = 0 ;
}
