netcdf \00010101.ocean_static.deptho {
dimensions:
	time = UNLIMITED ; // (1 currently)
	yh = 10 ;
	xh = 15 ;
	xq = 15 ;
	yq = 10 ;
variables:
	float deptho(yh, xh) ;
		deptho:_FillValue = 1.e+20f ;
		deptho:missing_value = 1.e+20f ;
		deptho:units = "m" ;
		deptho:long_name = "Sea Floor Depth" ;
		deptho:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		deptho:cell_measures = "area: areacello" ;
		deptho:standard_name = "sea_floor_depth_below_geoid" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Jun 13 14:06:58 2025: ncks -d xh,532,546 -d yh,526,535 -d xq,532,546 -d yq,526,535 /home/cew/Code/cmip7-sprint/testfiles/input/00010101.ocean_static.nc -O /home/cew/Code/cmip7-sprint/testfiles/00010101.ocean_static.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 deptho =
  5459.581, 5518.351, 5471.555, 5464.517, 5493.351, 5443.992, 5481.438, 
    5399.232, 5437.585, 5564.116, 5508.024, 5278.302, 5339.634, 5338.516, 
    5362.45,
  5444.997, 5526.517, 5558.977, 5506.794, 5539.163, 5464.714, 5371.029, 
    5283.403, 5344.632, 5276.831, 5453.903, 5460.983, 5401.993, 5373.839, 
    5222.505,
  5469.43, 5485.55, 5484.331, 5534.783, 5515.036, 5381.512, 5379.43, 
    5436.272, 5353.861, 5308.952, 5356.044, 5565.796, 5455.912, 5291.331, 
    5030.697,
  5377.339, 5432.107, 5414.18, 5474.686, 5430.449, 5403.279, 5411.458, 
    5495.017, 5410.293, 5379.038, 5393.203, 5604.945, 5393.119, 4742.138, 
    4438.138,
  5412.795, 5426.14, 5400.57, 5435.193, 5439.468, 5473.852, 5430.786, 
    5391.758, 5547.167, 5492.971, 5509.514, 5286.06, 4352.004, 4455.662, 
    3532.009,
  5441.89, 5533.067, 5532.043, 5451.808, 5465.8, 5563.95, 5503.784, 5289.503, 
    5447.585, 5495.046, 5438.338, 5136.738, 4889.081, 4330.568, 3322.158,
  5367.564, 5623.584, 5646.252, 5546.898, 5537.195, 5522.411, 4901.873, 
    5396.403, 5512.202, 5424.177, 5183.489, 5008.471, 5015.458, 3874.39, 
    3237.326,
  5536.536, 5390.403, 5186.029, 5572.206, 5660.611, 5683.173, 5679.197, 
    5480.841, 5338.633, 5219.022, 5189.761, 4972.972, 4596.265, 3853.92, 3078,
  5527.949, 5094.13, 4281.74, 5565.208, 5684.5, 5743.412, 5613.496, 5286.793, 
    5167.222, 5019.19, 4948.869, 4768.419, 4239.951, 3896.296, 3292.449,
  5542.585, 5490.353, 5468.412, 5531.694, 5649.889, 5580.06, 5496.899, 
    4881.083, 4591.047, 4642.272, 4266.763, 3973.73, 3807.69, 3853.071, 
    3504.758 ;

 time = 0 ;

 xh = -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 xq = -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 yh = -14.3476556382336, -14.1053228834302, -13.862732304759, 
    -13.6198879813569, -13.3767940148509, -13.1334545290505, 
    -12.889873669635, -12.6460556038367, -12.4020045201193, -12.1577246278516 ;

 yq = -14.4687240631789, -14.2265217428746, -13.9840595676627, 
    -13.7413416053212, -13.4983719462701, -13.2551547032665, 
    -13.011694011094, -12.7679940262485, -12.5240589266184, -12.279892911161 ;
}
